module basic_5000_50000_5000_25_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
or U0 (N_0,In_2939,In_4403);
nand U1 (N_1,In_3518,In_409);
nor U2 (N_2,In_268,In_4052);
xor U3 (N_3,In_192,In_844);
and U4 (N_4,In_3295,In_4066);
nor U5 (N_5,In_4554,In_801);
and U6 (N_6,In_3565,In_4630);
and U7 (N_7,In_2112,In_184);
nand U8 (N_8,In_2142,In_4875);
nand U9 (N_9,In_669,In_2318);
nor U10 (N_10,In_2342,In_3659);
xor U11 (N_11,In_4786,In_2212);
nor U12 (N_12,In_1544,In_3523);
nor U13 (N_13,In_4046,In_4252);
nand U14 (N_14,In_3081,In_222);
and U15 (N_15,In_4010,In_1507);
nor U16 (N_16,In_2160,In_1153);
xor U17 (N_17,In_3801,In_3242);
nor U18 (N_18,In_2822,In_3316);
or U19 (N_19,In_3310,In_749);
and U20 (N_20,In_2666,In_1754);
and U21 (N_21,In_4412,In_657);
xor U22 (N_22,In_2698,In_4043);
and U23 (N_23,In_1430,In_322);
nor U24 (N_24,In_355,In_1368);
nand U25 (N_25,In_3756,In_3172);
nor U26 (N_26,In_893,In_2231);
nor U27 (N_27,In_1637,In_3581);
nand U28 (N_28,In_4406,In_599);
or U29 (N_29,In_1003,In_3837);
nand U30 (N_30,In_983,In_2158);
nor U31 (N_31,In_3309,In_2128);
and U32 (N_32,In_284,In_2030);
nand U33 (N_33,In_3326,In_4433);
and U34 (N_34,In_3584,In_3588);
xor U35 (N_35,In_4131,In_4409);
or U36 (N_36,In_3069,In_2347);
nor U37 (N_37,In_3270,In_2750);
nor U38 (N_38,In_1363,In_3332);
or U39 (N_39,In_1574,In_1538);
or U40 (N_40,In_1858,In_3506);
nand U41 (N_41,In_3184,In_579);
and U42 (N_42,In_122,In_802);
nand U43 (N_43,In_4949,In_3196);
and U44 (N_44,In_2528,In_4099);
nand U45 (N_45,In_1839,In_2092);
nand U46 (N_46,In_3449,In_3509);
xnor U47 (N_47,In_1037,In_4021);
and U48 (N_48,In_787,In_2287);
xnor U49 (N_49,In_4737,In_2174);
or U50 (N_50,In_1552,In_2751);
nand U51 (N_51,In_2619,In_2562);
nand U52 (N_52,In_1567,In_3194);
and U53 (N_53,In_1540,In_4995);
or U54 (N_54,In_1585,In_2912);
and U55 (N_55,In_2625,In_4226);
nor U56 (N_56,In_794,In_803);
nand U57 (N_57,In_2982,In_1974);
nor U58 (N_58,In_2059,In_508);
xnor U59 (N_59,In_3403,In_2977);
or U60 (N_60,In_3789,In_4727);
nand U61 (N_61,In_4149,In_4808);
or U62 (N_62,In_373,In_9);
nor U63 (N_63,In_3397,In_1164);
xnor U64 (N_64,In_4474,In_4861);
xnor U65 (N_65,In_1563,In_3420);
nor U66 (N_66,In_82,In_890);
nand U67 (N_67,In_4680,In_3535);
or U68 (N_68,In_2271,In_2333);
or U69 (N_69,In_2875,In_540);
nand U70 (N_70,In_1799,In_208);
and U71 (N_71,In_4364,In_3440);
xnor U72 (N_72,In_4061,In_554);
or U73 (N_73,In_1231,In_4651);
nor U74 (N_74,In_1741,In_1838);
nand U75 (N_75,In_2456,In_1206);
nand U76 (N_76,In_443,In_2466);
nand U77 (N_77,In_2246,In_2644);
or U78 (N_78,In_2087,In_851);
nor U79 (N_79,In_3505,In_2754);
xnor U80 (N_80,In_814,In_45);
nand U81 (N_81,In_3973,In_1715);
nor U82 (N_82,In_2260,In_4846);
and U83 (N_83,In_2501,In_2366);
or U84 (N_84,In_1590,In_992);
or U85 (N_85,In_569,In_245);
nor U86 (N_86,In_1528,In_3849);
nor U87 (N_87,In_3266,In_3923);
nor U88 (N_88,In_2304,In_1808);
and U89 (N_89,In_1644,In_1381);
and U90 (N_90,In_4877,In_3094);
and U91 (N_91,In_4550,In_4038);
xnor U92 (N_92,In_2392,In_1142);
and U93 (N_93,In_22,In_3103);
nor U94 (N_94,In_435,In_3753);
and U95 (N_95,In_4289,In_832);
nand U96 (N_96,In_4696,In_3624);
xor U97 (N_97,In_1539,In_4481);
nand U98 (N_98,In_2767,In_3180);
nand U99 (N_99,In_3394,In_954);
and U100 (N_100,In_1118,In_2129);
nand U101 (N_101,In_3031,In_3819);
and U102 (N_102,In_2435,In_1559);
nand U103 (N_103,In_1271,In_4055);
and U104 (N_104,In_1289,In_2487);
nor U105 (N_105,In_3878,In_3743);
xnor U106 (N_106,In_1401,In_155);
or U107 (N_107,In_2937,In_4675);
nand U108 (N_108,In_532,In_2821);
xor U109 (N_109,In_3437,In_4771);
nor U110 (N_110,In_734,In_156);
and U111 (N_111,In_4411,In_1583);
or U112 (N_112,In_4785,In_1944);
xnor U113 (N_113,In_3728,In_417);
nor U114 (N_114,In_2918,In_3919);
and U115 (N_115,In_4393,In_1143);
nor U116 (N_116,In_1973,In_2150);
or U117 (N_117,In_4421,In_4624);
nor U118 (N_118,In_791,In_3223);
or U119 (N_119,In_1367,In_610);
or U120 (N_120,In_4767,In_2125);
xor U121 (N_121,In_3576,In_1155);
xnor U122 (N_122,In_4265,In_2868);
nor U123 (N_123,In_1092,In_2100);
nor U124 (N_124,In_312,In_1774);
and U125 (N_125,In_4320,In_2393);
nand U126 (N_126,In_4606,In_2682);
and U127 (N_127,In_2293,In_1285);
and U128 (N_128,In_3469,In_4078);
nor U129 (N_129,In_1776,In_464);
nand U130 (N_130,In_2034,In_2403);
and U131 (N_131,In_4479,In_2075);
or U132 (N_132,In_1679,In_3977);
or U133 (N_133,In_478,In_3820);
or U134 (N_134,In_2014,In_4962);
and U135 (N_135,In_416,In_473);
or U136 (N_136,In_4672,In_3736);
and U137 (N_137,In_3544,In_3924);
nand U138 (N_138,In_2406,In_2820);
or U139 (N_139,In_3818,In_658);
and U140 (N_140,In_1959,In_1803);
and U141 (N_141,In_2976,In_399);
nand U142 (N_142,In_2131,In_2355);
xnor U143 (N_143,In_1364,In_446);
nor U144 (N_144,In_4908,In_793);
nor U145 (N_145,In_3459,In_4015);
xnor U146 (N_146,In_1110,In_4080);
or U147 (N_147,In_4519,In_2575);
xor U148 (N_148,In_4148,In_1758);
and U149 (N_149,In_199,In_4313);
and U150 (N_150,In_1900,In_2923);
xor U151 (N_151,In_2073,In_2770);
and U152 (N_152,In_4595,In_1829);
nand U153 (N_153,In_1467,In_58);
nand U154 (N_154,In_574,In_2949);
and U155 (N_155,In_424,In_2864);
nor U156 (N_156,In_1094,In_1470);
or U157 (N_157,In_3467,In_2235);
nor U158 (N_158,In_412,In_936);
nor U159 (N_159,In_1211,In_915);
nand U160 (N_160,In_1713,In_1300);
or U161 (N_161,In_2119,In_518);
nor U162 (N_162,In_4490,In_1924);
nand U163 (N_163,In_2683,In_2654);
nor U164 (N_164,In_700,In_3807);
nor U165 (N_165,In_2773,In_4706);
or U166 (N_166,In_1055,In_3873);
xnor U167 (N_167,In_3298,In_2900);
and U168 (N_168,In_1498,In_976);
and U169 (N_169,In_4452,In_2757);
or U170 (N_170,In_1920,In_829);
nor U171 (N_171,In_3043,In_3092);
nand U172 (N_172,In_105,In_1443);
nand U173 (N_173,In_3626,In_1454);
nor U174 (N_174,In_4203,In_4363);
xnor U175 (N_175,In_2993,In_3828);
or U176 (N_176,In_2680,In_4016);
or U177 (N_177,In_2960,In_54);
xnor U178 (N_178,In_3466,In_1531);
or U179 (N_179,In_4954,In_3607);
nor U180 (N_180,In_2455,In_1852);
xor U181 (N_181,In_3610,In_2673);
or U182 (N_182,In_987,In_3978);
nor U183 (N_183,In_4604,In_62);
and U184 (N_184,In_2672,In_2249);
and U185 (N_185,In_4821,In_4563);
or U186 (N_186,In_4612,In_4723);
or U187 (N_187,In_2042,In_789);
nor U188 (N_188,In_2892,In_3646);
and U189 (N_189,In_3,In_1685);
nor U190 (N_190,In_432,In_581);
nor U191 (N_191,In_1221,In_3453);
nor U192 (N_192,In_1301,In_1500);
and U193 (N_193,In_3246,In_948);
nor U194 (N_194,In_2439,In_583);
or U195 (N_195,In_349,In_3686);
xor U196 (N_196,In_782,In_1875);
nand U197 (N_197,In_390,In_938);
and U198 (N_198,In_2447,In_2274);
nand U199 (N_199,In_4151,In_4269);
and U200 (N_200,In_3300,In_2186);
xor U201 (N_201,In_1566,In_203);
nand U202 (N_202,In_3853,In_838);
nor U203 (N_203,In_14,In_3110);
or U204 (N_204,In_1186,In_535);
xnor U205 (N_205,In_605,In_1691);
and U206 (N_206,In_1114,In_391);
xnor U207 (N_207,In_546,In_524);
nor U208 (N_208,In_152,In_1284);
and U209 (N_209,In_1948,In_2958);
nor U210 (N_210,In_4556,In_1485);
and U211 (N_211,In_2047,In_4611);
or U212 (N_212,In_3579,In_1358);
nor U213 (N_213,In_4152,In_848);
nor U214 (N_214,In_4516,In_217);
or U215 (N_215,In_32,In_3770);
and U216 (N_216,In_3158,In_2675);
and U217 (N_217,In_3694,In_4960);
nand U218 (N_218,In_1650,In_151);
xnor U219 (N_219,In_2394,In_3857);
nand U220 (N_220,In_698,In_258);
or U221 (N_221,In_1343,In_2259);
nand U222 (N_222,In_650,In_1756);
and U223 (N_223,In_709,In_1747);
nor U224 (N_224,In_4841,In_1684);
and U225 (N_225,In_4378,In_41);
nand U226 (N_226,In_3755,In_1322);
or U227 (N_227,In_163,In_3815);
and U228 (N_228,In_4537,In_3229);
nand U229 (N_229,In_447,In_1910);
nand U230 (N_230,In_4157,In_2498);
nor U231 (N_231,In_2825,In_4872);
xor U232 (N_232,In_4628,In_1380);
nand U233 (N_233,In_1148,In_4141);
nor U234 (N_234,In_1666,In_2718);
nor U235 (N_235,In_4386,In_897);
nand U236 (N_236,In_1617,In_950);
nand U237 (N_237,In_3665,In_4114);
or U238 (N_238,In_3721,In_2413);
nand U239 (N_239,In_2307,In_598);
xnor U240 (N_240,In_4329,In_840);
xnor U241 (N_241,In_2827,In_3008);
xnor U242 (N_242,In_1259,In_3143);
or U243 (N_243,In_1082,In_1378);
nor U244 (N_244,In_2512,In_4986);
xnor U245 (N_245,In_2678,In_364);
and U246 (N_246,In_2152,In_1336);
nor U247 (N_247,In_1714,In_4561);
or U248 (N_248,In_2987,In_4530);
or U249 (N_249,In_604,In_23);
and U250 (N_250,In_188,In_1266);
nor U251 (N_251,In_295,In_3577);
and U252 (N_252,In_1763,In_2179);
or U253 (N_253,In_2148,In_288);
xor U254 (N_254,In_2370,In_2584);
and U255 (N_255,In_1993,In_2273);
and U256 (N_256,In_633,In_3943);
nor U257 (N_257,In_1668,In_1742);
nand U258 (N_258,In_4056,In_1111);
and U259 (N_259,In_2414,In_1177);
nand U260 (N_260,In_4221,In_4577);
nand U261 (N_261,In_2572,In_4643);
or U262 (N_262,In_4301,In_2991);
nor U263 (N_263,In_2348,In_3843);
xnor U264 (N_264,In_1136,In_1862);
nand U265 (N_265,In_1333,In_3503);
nand U266 (N_266,In_3429,In_3240);
and U267 (N_267,In_4180,In_2634);
nand U268 (N_268,In_2614,In_4116);
and U269 (N_269,In_568,In_566);
and U270 (N_270,In_3785,In_3946);
xnor U271 (N_271,In_1699,In_760);
nand U272 (N_272,In_4568,In_3017);
and U273 (N_273,In_1984,In_1176);
or U274 (N_274,In_310,In_495);
nor U275 (N_275,In_1847,In_2922);
and U276 (N_276,In_1365,In_3417);
xnor U277 (N_277,In_1295,In_4354);
and U278 (N_278,In_4002,In_3809);
nor U279 (N_279,In_1441,In_110);
and U280 (N_280,In_3638,In_1116);
xnor U281 (N_281,In_2289,In_1703);
nand U282 (N_282,In_2668,In_1814);
nor U283 (N_283,In_1825,In_396);
nor U284 (N_284,In_3934,In_2190);
nor U285 (N_285,In_3104,In_3513);
or U286 (N_286,In_2856,In_3562);
nor U287 (N_287,In_2924,In_1410);
xnor U288 (N_288,In_393,In_2409);
or U289 (N_289,In_2037,In_3254);
or U290 (N_290,In_4473,In_3619);
or U291 (N_291,In_2758,In_4136);
xnor U292 (N_292,In_15,In_2566);
and U293 (N_293,In_2805,In_4968);
or U294 (N_294,In_3292,In_3838);
xor U295 (N_295,In_1234,In_528);
xor U296 (N_296,In_644,In_2464);
nand U297 (N_297,In_2156,In_1282);
and U298 (N_298,In_4186,In_2188);
and U299 (N_299,In_1936,In_1866);
or U300 (N_300,In_1844,In_1070);
xor U301 (N_301,In_4396,In_4208);
and U302 (N_302,In_2839,In_4984);
and U303 (N_303,In_663,In_3552);
nor U304 (N_304,In_2296,In_382);
and U305 (N_305,In_692,In_229);
nand U306 (N_306,In_1989,In_4246);
and U307 (N_307,In_1612,In_2986);
or U308 (N_308,In_3937,In_1375);
nor U309 (N_309,In_1723,In_1901);
and U310 (N_310,In_3011,In_296);
or U311 (N_311,In_1298,In_3117);
xor U312 (N_312,In_4772,In_3333);
nand U313 (N_313,In_193,In_1853);
nor U314 (N_314,In_4024,In_1731);
xor U315 (N_315,In_4076,In_3542);
nor U316 (N_316,In_1571,In_218);
nand U317 (N_317,In_150,In_525);
and U318 (N_318,In_4688,In_3091);
nor U319 (N_319,In_3426,In_2191);
and U320 (N_320,In_406,In_2791);
nor U321 (N_321,In_71,In_3670);
or U322 (N_322,In_2649,In_503);
or U323 (N_323,In_211,In_2007);
xor U324 (N_324,In_3222,In_1213);
nand U325 (N_325,In_640,In_1214);
nand U326 (N_326,In_2185,In_4726);
or U327 (N_327,In_2914,In_781);
and U328 (N_328,In_690,In_1857);
or U329 (N_329,In_4679,In_255);
and U330 (N_330,In_2226,In_1694);
or U331 (N_331,In_3026,In_2570);
or U332 (N_332,In_265,In_3001);
xnor U333 (N_333,In_3307,In_687);
nor U334 (N_334,In_2266,In_3649);
and U335 (N_335,In_2207,In_4096);
nand U336 (N_336,In_65,In_3205);
xor U337 (N_337,In_2078,In_1690);
or U338 (N_338,In_2748,In_3377);
or U339 (N_339,In_4491,In_4695);
xor U340 (N_340,In_2039,In_4361);
xor U341 (N_341,In_2421,In_2703);
nor U342 (N_342,In_4918,In_4093);
nand U343 (N_343,In_11,In_1011);
xnor U344 (N_344,In_3095,In_1426);
nand U345 (N_345,In_4860,In_4536);
nand U346 (N_346,In_1260,In_1504);
and U347 (N_347,In_142,In_4719);
or U348 (N_348,In_2390,In_3428);
and U349 (N_349,In_3217,In_4333);
nor U350 (N_350,In_750,In_3048);
xor U351 (N_351,In_127,In_3303);
nand U352 (N_352,In_543,In_2088);
nand U353 (N_353,In_4807,In_816);
xor U354 (N_354,In_1874,In_3102);
and U355 (N_355,In_526,In_632);
and U356 (N_356,In_3623,In_3707);
and U357 (N_357,In_4047,In_974);
nand U358 (N_358,In_4236,In_3971);
xor U359 (N_359,In_4826,In_3167);
and U360 (N_360,In_3145,In_2558);
nand U361 (N_361,In_4032,In_2520);
or U362 (N_362,In_2133,In_666);
nor U363 (N_363,In_3073,In_3149);
xnor U364 (N_364,In_1772,In_4738);
nand U365 (N_365,In_4469,In_3522);
nor U366 (N_366,In_738,In_631);
or U367 (N_367,In_2015,In_2070);
nor U368 (N_368,In_1501,In_3765);
or U369 (N_369,In_1914,In_710);
nand U370 (N_370,In_2609,In_4763);
and U371 (N_371,In_261,In_1074);
xor U372 (N_372,In_4322,In_1352);
and U373 (N_373,In_2033,In_2084);
and U374 (N_374,In_3047,In_1089);
or U375 (N_375,In_3633,In_1979);
and U376 (N_376,In_1005,In_2488);
and U377 (N_377,In_1876,In_2103);
or U378 (N_378,In_1387,In_3913);
xnor U379 (N_379,In_3134,In_178);
xor U380 (N_380,In_3286,In_86);
and U381 (N_381,In_4553,In_1670);
nor U382 (N_382,In_3359,In_2899);
and U383 (N_383,In_665,In_1591);
nand U384 (N_384,In_4258,In_1344);
xnor U385 (N_385,In_111,In_4929);
nor U386 (N_386,In_3261,In_2517);
or U387 (N_387,In_708,In_2658);
or U388 (N_388,In_370,In_1311);
nand U389 (N_389,In_3601,In_3364);
nand U390 (N_390,In_3460,In_2154);
or U391 (N_391,In_3639,In_1191);
nor U392 (N_392,In_4665,In_1242);
or U393 (N_393,In_1614,In_2518);
and U394 (N_394,In_1218,In_759);
nand U395 (N_395,In_3808,In_4829);
xnor U396 (N_396,In_2146,In_4887);
nor U397 (N_397,In_4483,In_3587);
nand U398 (N_398,In_3448,In_3224);
nor U399 (N_399,In_1908,In_2239);
xnor U400 (N_400,In_891,In_2021);
or U401 (N_401,In_1072,In_4725);
and U402 (N_402,In_4071,In_2012);
and U403 (N_403,In_2963,In_3508);
or U404 (N_404,In_2589,In_1643);
and U405 (N_405,In_1719,In_4220);
or U406 (N_406,In_4040,In_719);
or U407 (N_407,In_4343,In_2324);
or U408 (N_408,In_36,In_4605);
nand U409 (N_409,In_2854,In_995);
and U410 (N_410,In_910,In_3101);
xnor U411 (N_411,In_2699,In_4617);
and U412 (N_412,In_981,In_1315);
and U413 (N_413,In_3836,In_1930);
xor U414 (N_414,In_1257,In_1593);
or U415 (N_415,In_4276,In_1018);
and U416 (N_416,In_4170,In_394);
xnor U417 (N_417,In_648,In_3390);
or U418 (N_418,In_2928,In_1325);
xor U419 (N_419,In_1717,In_269);
or U420 (N_420,In_2327,In_3991);
nand U421 (N_421,In_298,In_805);
nand U422 (N_422,In_757,In_2247);
nand U423 (N_423,In_2395,In_130);
nand U424 (N_424,In_1299,In_701);
or U425 (N_425,In_3621,In_1098);
or U426 (N_426,In_788,In_3336);
nor U427 (N_427,In_4121,In_2026);
nand U428 (N_428,In_2879,In_4891);
xnor U429 (N_429,In_3410,In_3966);
and U430 (N_430,In_426,In_2136);
nand U431 (N_431,In_4117,In_3250);
xnor U432 (N_432,In_4060,In_2588);
and U433 (N_433,In_884,In_360);
nand U434 (N_434,In_4710,In_161);
nor U435 (N_435,In_213,In_3965);
nand U436 (N_436,In_2916,In_1199);
xor U437 (N_437,In_4224,In_4685);
nand U438 (N_438,In_2617,In_3931);
nor U439 (N_439,In_2338,In_3214);
nor U440 (N_440,In_4797,In_4341);
xnor U441 (N_441,In_351,In_593);
and U442 (N_442,In_4230,In_4248);
xnor U443 (N_443,In_323,In_3539);
nor U444 (N_444,In_227,In_3140);
and U445 (N_445,In_1709,In_1052);
or U446 (N_446,In_3122,In_2140);
and U447 (N_447,In_922,In_2743);
xnor U448 (N_448,In_3635,In_1499);
or U449 (N_449,In_3471,In_4042);
nor U450 (N_450,In_12,In_1706);
nand U451 (N_451,In_1716,In_3572);
and U452 (N_452,In_4172,In_1562);
and U453 (N_453,In_3760,In_1794);
nand U454 (N_454,In_3450,In_3941);
xnor U455 (N_455,In_548,In_1558);
or U456 (N_456,In_1041,In_2031);
xor U457 (N_457,In_2897,In_1798);
nor U458 (N_458,In_1941,In_1466);
nand U459 (N_459,In_2647,In_1887);
nand U460 (N_460,In_654,In_3510);
nor U461 (N_461,In_462,In_154);
nor U462 (N_462,In_4026,In_2244);
xor U463 (N_463,In_3846,In_4440);
xnor U464 (N_464,In_754,In_2571);
or U465 (N_465,In_4247,In_2123);
xor U466 (N_466,In_3540,In_455);
and U467 (N_467,In_3276,In_1506);
xnor U468 (N_468,In_4708,In_868);
nor U469 (N_469,In_4123,In_3538);
nor U470 (N_470,In_1681,In_3960);
nand U471 (N_471,In_2947,In_2432);
nand U472 (N_472,In_588,In_2543);
and U473 (N_473,In_3352,In_240);
xnor U474 (N_474,In_2894,In_216);
xor U475 (N_475,In_3500,In_1113);
or U476 (N_476,In_3938,In_3338);
or U477 (N_477,In_169,In_1764);
or U478 (N_478,In_4880,In_1028);
xnor U479 (N_479,In_2515,In_1580);
nand U480 (N_480,In_1320,In_4864);
xor U481 (N_481,In_4511,In_877);
and U482 (N_482,In_10,In_4165);
nor U483 (N_483,In_250,In_1149);
nand U484 (N_484,In_3614,In_3514);
xnor U485 (N_485,In_4755,In_2412);
and U486 (N_486,In_1296,In_2760);
and U487 (N_487,In_1252,In_2643);
nor U488 (N_488,In_1620,In_4823);
nor U489 (N_489,In_479,In_3065);
or U490 (N_490,In_2232,In_4994);
nor U491 (N_491,In_2277,In_3676);
xnor U492 (N_492,In_3763,In_3715);
nand U493 (N_493,In_3906,In_3021);
nor U494 (N_494,In_3629,In_2374);
nand U495 (N_495,In_1475,In_4260);
or U496 (N_496,In_1280,In_1788);
nand U497 (N_497,In_3136,In_2869);
nor U498 (N_498,In_328,In_1452);
and U499 (N_499,In_2491,In_2779);
or U500 (N_500,In_1837,In_2745);
xor U501 (N_501,In_3443,In_2422);
xnor U502 (N_502,In_78,In_1753);
or U503 (N_503,In_1130,In_2215);
xor U504 (N_504,In_401,In_1128);
nor U505 (N_505,In_244,In_817);
and U506 (N_506,In_3957,In_3348);
or U507 (N_507,In_4657,In_55);
xor U508 (N_508,In_712,In_906);
and U509 (N_509,In_1196,In_1511);
nor U510 (N_510,In_626,In_57);
and U511 (N_511,In_3634,In_3221);
nor U512 (N_512,In_2314,In_2263);
and U513 (N_513,In_1276,In_3220);
or U514 (N_514,In_4906,In_3648);
nand U515 (N_515,In_3474,In_1548);
xor U516 (N_516,In_1613,In_4307);
and U517 (N_517,In_1739,In_4415);
nand U518 (N_518,In_2706,In_1929);
nand U519 (N_519,In_3035,In_2648);
xnor U520 (N_520,In_1459,In_1261);
nor U521 (N_521,In_980,In_3653);
nand U522 (N_522,In_1437,In_4735);
xnor U523 (N_523,In_4145,In_4133);
xnor U524 (N_524,In_902,In_2019);
and U525 (N_525,In_1351,In_2241);
nand U526 (N_526,In_4642,In_2983);
xor U527 (N_527,In_3392,In_4018);
or U528 (N_528,In_3419,In_1255);
and U529 (N_529,In_3880,In_1881);
and U530 (N_530,In_1262,In_1581);
nand U531 (N_531,In_901,In_4896);
xor U532 (N_532,In_489,In_1610);
or U533 (N_533,In_716,In_134);
or U534 (N_534,In_4128,In_3285);
nand U535 (N_535,In_3150,In_1222);
and U536 (N_536,In_1088,In_3383);
nand U537 (N_537,In_4989,In_1103);
nor U538 (N_538,In_3144,In_1649);
nor U539 (N_539,In_187,In_1425);
nand U540 (N_540,In_3495,In_4990);
nand U541 (N_541,In_779,In_4477);
nor U542 (N_542,In_3688,In_2707);
or U543 (N_543,In_1561,In_3989);
xnor U544 (N_544,In_3959,In_205);
nor U545 (N_545,In_4594,In_1968);
xor U546 (N_546,In_3375,In_3687);
nor U547 (N_547,In_4204,In_1856);
or U548 (N_548,In_622,In_3100);
xnor U549 (N_549,In_4009,In_4634);
xor U550 (N_550,In_1870,In_88);
nand U551 (N_551,In_1241,In_859);
xor U552 (N_552,In_3473,In_645);
nand U553 (N_553,In_1292,In_2067);
xor U554 (N_554,In_3729,In_1460);
or U555 (N_555,In_2620,In_4251);
and U556 (N_556,In_4054,In_1060);
or U557 (N_557,In_267,In_536);
or U558 (N_558,In_2514,In_1646);
xnor U559 (N_559,In_985,In_852);
or U560 (N_560,In_2062,In_600);
or U561 (N_561,In_338,In_4788);
nor U562 (N_562,In_4713,In_1270);
and U563 (N_563,In_474,In_1992);
nor U564 (N_564,In_3015,In_1995);
or U565 (N_565,In_234,In_601);
or U566 (N_566,In_407,In_2199);
nand U567 (N_567,In_2002,In_387);
and U568 (N_568,In_1013,In_3032);
nand U569 (N_569,In_1748,In_1616);
and U570 (N_570,In_1471,In_2974);
xnor U571 (N_571,In_3598,In_2253);
xor U572 (N_572,In_4843,In_2218);
nor U573 (N_573,In_3115,In_3054);
xor U574 (N_574,In_215,In_2214);
and U575 (N_575,In_4413,In_2857);
nor U576 (N_576,In_3232,In_874);
xnor U577 (N_577,In_400,In_3613);
nor U578 (N_578,In_1383,In_4715);
nor U579 (N_579,In_3086,In_3181);
or U580 (N_580,In_2637,In_4504);
nor U581 (N_581,In_3373,In_4351);
or U582 (N_582,In_3325,In_4274);
or U583 (N_583,In_4712,In_634);
nor U584 (N_584,In_2684,In_4671);
nor U585 (N_585,In_3877,In_3125);
or U586 (N_586,In_748,In_1084);
nand U587 (N_587,In_3833,In_892);
nor U588 (N_588,In_2623,In_2426);
and U589 (N_589,In_682,In_3247);
or U590 (N_590,In_232,In_118);
nand U591 (N_591,In_2752,In_2474);
xnor U592 (N_592,In_1537,In_3121);
nor U593 (N_593,In_3457,In_3166);
nand U594 (N_594,In_475,In_3477);
and U595 (N_595,In_1890,In_4105);
nand U596 (N_596,In_1955,In_1135);
xor U597 (N_597,In_3288,In_272);
nand U598 (N_598,In_3447,In_3832);
and U599 (N_599,In_2870,In_1834);
xor U600 (N_600,In_4743,In_2952);
xnor U601 (N_601,In_1031,In_3810);
or U602 (N_602,In_375,In_2704);
nor U603 (N_603,In_2813,In_4721);
xor U604 (N_604,In_4104,In_228);
nand U605 (N_605,In_705,In_4164);
and U606 (N_606,In_680,In_4268);
nor U607 (N_607,In_1445,In_429);
and U608 (N_608,In_1399,In_4531);
and U609 (N_609,In_4559,In_1768);
nand U610 (N_610,In_372,In_1288);
and U611 (N_611,In_4597,In_2890);
nor U612 (N_612,In_4836,In_1030);
xor U613 (N_613,In_3899,In_4280);
or U614 (N_614,In_4178,In_2339);
or U615 (N_615,In_3675,In_900);
nand U616 (N_616,In_3967,In_2826);
xor U617 (N_617,In_3424,In_369);
and U618 (N_618,In_1810,In_1319);
nor U619 (N_619,In_2664,In_1146);
or U620 (N_620,In_3408,In_2990);
nor U621 (N_621,In_551,In_4119);
or U622 (N_622,In_3068,In_1317);
xnor U623 (N_623,In_3814,In_3725);
and U624 (N_624,In_3560,In_1240);
and U625 (N_625,In_2130,In_18);
nor U626 (N_626,In_4648,In_3131);
xor U627 (N_627,In_2669,In_1604);
and U628 (N_628,In_1369,In_3396);
xor U629 (N_629,In_867,In_3841);
and U630 (N_630,In_3439,In_4800);
nor U631 (N_631,In_3493,In_2369);
and U632 (N_632,In_2946,In_1836);
nor U633 (N_633,In_4703,In_3088);
xor U634 (N_634,In_977,In_4575);
nor U635 (N_635,In_4586,In_1554);
and U636 (N_636,In_1263,In_35);
nor U637 (N_637,In_3418,In_13);
or U638 (N_638,In_1664,In_4485);
nor U639 (N_639,In_3803,In_1569);
or U640 (N_640,In_121,In_3640);
nand U641 (N_641,In_1335,In_43);
xor U642 (N_642,In_40,In_2283);
and U643 (N_643,In_1264,In_3876);
and U644 (N_644,In_2113,In_1496);
or U645 (N_645,In_2523,In_4253);
nor U646 (N_646,In_2862,In_3273);
or U647 (N_647,In_320,In_66);
nand U648 (N_648,In_2089,In_1725);
or U649 (N_649,In_301,In_761);
xor U650 (N_650,In_2323,In_4782);
nand U651 (N_651,In_4524,In_4964);
nor U652 (N_652,In_4613,In_4905);
xnor U653 (N_653,In_4293,In_4316);
nand U654 (N_654,In_243,In_3727);
nand U655 (N_655,In_836,In_4297);
nor U656 (N_656,In_4209,In_4692);
or U657 (N_657,In_3272,In_1100);
xnor U658 (N_658,In_1708,In_1209);
or U659 (N_659,In_4885,In_2382);
and U660 (N_660,In_3255,In_2800);
xnor U661 (N_661,In_752,In_2269);
nor U662 (N_662,In_3645,In_4094);
and U663 (N_663,In_488,In_3782);
nand U664 (N_664,In_2115,In_4304);
nor U665 (N_665,In_3176,In_2043);
or U666 (N_666,In_2898,In_1534);
or U667 (N_667,In_774,In_4340);
xor U668 (N_668,In_1895,In_83);
nor U669 (N_669,In_2169,In_2689);
and U670 (N_670,In_4231,In_1778);
xor U671 (N_671,In_4423,In_570);
and U672 (N_672,In_1438,In_3147);
xor U673 (N_673,In_3984,In_345);
nand U674 (N_674,In_4127,In_436);
xor U675 (N_675,In_3337,In_294);
nor U676 (N_676,In_4866,In_4328);
and U677 (N_677,In_1912,In_1830);
nand U678 (N_678,In_3182,In_3034);
and U679 (N_679,In_3339,In_1896);
and U680 (N_680,In_186,In_2484);
nand U681 (N_681,In_1812,In_4831);
xnor U682 (N_682,In_1698,In_4532);
xnor U683 (N_683,In_1589,In_4373);
and U684 (N_684,In_1492,In_2719);
nor U685 (N_685,In_4509,In_4660);
nor U686 (N_686,In_221,In_4948);
xnor U687 (N_687,In_2828,In_2011);
nor U688 (N_688,In_4299,In_751);
nand U689 (N_689,In_2985,In_1105);
or U690 (N_690,In_4238,In_2736);
nand U691 (N_691,In_627,In_3162);
or U692 (N_692,In_3974,In_4176);
nor U693 (N_693,In_714,In_1216);
xor U694 (N_694,In_766,In_2118);
and U695 (N_695,In_4227,In_4574);
nor U696 (N_696,In_4489,In_4756);
nor U697 (N_697,In_2145,In_2832);
xnor U698 (N_698,In_2308,In_4687);
nor U699 (N_699,In_1630,In_2094);
nor U700 (N_700,In_324,In_3311);
nand U701 (N_701,In_3987,In_630);
and U702 (N_702,In_1239,In_3999);
nand U703 (N_703,In_2602,In_2303);
xnor U704 (N_704,In_1346,In_1791);
or U705 (N_705,In_1059,In_3040);
or U706 (N_706,In_1187,In_4924);
nand U707 (N_707,In_2090,In_2054);
or U708 (N_708,In_280,In_4189);
nand U709 (N_709,In_4773,In_978);
nor U710 (N_710,In_678,In_933);
nand U711 (N_711,In_2910,In_180);
nor U712 (N_712,In_42,In_2741);
nor U713 (N_713,In_3367,In_4407);
nor U714 (N_714,In_1345,In_3672);
and U715 (N_715,In_1108,In_1269);
and U716 (N_716,In_1045,In_3969);
or U717 (N_717,In_3695,In_3305);
or U718 (N_718,In_567,In_4928);
and U719 (N_719,In_4930,In_1243);
nor U720 (N_720,In_4228,In_2772);
nor U721 (N_721,In_292,In_1268);
xnor U722 (N_722,In_1245,In_33);
or U723 (N_723,In_1855,In_3208);
and U724 (N_724,In_3757,In_1570);
nand U725 (N_725,In_4259,In_3183);
and U726 (N_726,In_3593,In_2956);
and U727 (N_727,In_4927,In_2592);
nand U728 (N_728,In_4317,In_1075);
and U729 (N_729,In_2797,In_274);
nor U730 (N_730,In_4374,In_3012);
nand U731 (N_731,In_3666,In_4515);
nor U732 (N_732,In_472,In_3884);
and U733 (N_733,In_997,In_305);
or U734 (N_734,In_989,In_795);
nand U735 (N_735,In_2877,In_1131);
nand U736 (N_736,In_4272,In_2053);
nand U737 (N_737,In_943,In_656);
and U738 (N_738,In_1469,In_2726);
xnor U739 (N_739,In_2110,In_804);
or U740 (N_740,In_3543,In_1960);
nor U741 (N_741,In_2691,In_251);
or U742 (N_742,In_2749,In_2243);
and U743 (N_743,In_1781,In_1210);
xnor U744 (N_744,In_4308,In_1073);
and U745 (N_745,In_4234,In_2401);
or U746 (N_746,In_2352,In_3312);
xnor U747 (N_747,In_4132,In_2099);
and U748 (N_748,In_4678,In_4045);
xnor U749 (N_749,In_1893,In_2267);
or U750 (N_750,In_2483,In_170);
xnor U751 (N_751,In_2358,In_2265);
xor U752 (N_752,In_242,In_2845);
nand U753 (N_753,In_2117,In_3831);
and U754 (N_754,In_1693,In_3042);
and U755 (N_755,In_3747,In_1621);
and U756 (N_756,In_53,In_3004);
xnor U757 (N_757,In_2601,In_4818);
nor U758 (N_758,In_3865,In_4034);
xnor U759 (N_759,In_2375,In_2252);
xor U760 (N_760,In_869,In_3372);
nor U761 (N_761,In_1529,In_982);
or U762 (N_762,In_4089,In_968);
xor U763 (N_763,In_4443,In_453);
or U764 (N_764,In_1598,In_4035);
nor U765 (N_765,In_2763,In_2920);
and U766 (N_766,In_1721,In_4894);
xnor U767 (N_767,In_4366,In_3682);
xor U768 (N_768,In_1790,In_725);
nor U769 (N_769,In_3128,In_2220);
nand U770 (N_770,In_504,In_2859);
or U771 (N_771,In_637,In_4270);
nand U772 (N_772,In_1811,In_522);
and U773 (N_773,In_1928,In_4352);
and U774 (N_774,In_3446,In_3813);
xor U775 (N_775,In_1692,In_461);
or U776 (N_776,In_1516,In_2803);
nor U777 (N_777,In_2362,In_4130);
nand U778 (N_778,In_4919,In_2107);
nor U779 (N_779,In_2843,In_4349);
nand U780 (N_780,In_2051,In_2457);
or U781 (N_781,In_3597,In_1409);
nand U782 (N_782,In_1969,In_1039);
nand U783 (N_783,In_403,In_4000);
or U784 (N_784,In_2685,In_2387);
and U785 (N_785,In_676,In_3123);
or U786 (N_786,In_2887,In_547);
nand U787 (N_787,In_1491,In_855);
xor U788 (N_788,In_3483,In_1519);
or U789 (N_789,In_683,In_3668);
nand U790 (N_790,In_3708,In_4661);
or U791 (N_791,In_4822,In_2134);
and U792 (N_792,In_4359,In_378);
or U793 (N_793,In_4883,In_2801);
nand U794 (N_794,In_560,In_2470);
and U795 (N_795,In_1198,In_1964);
or U796 (N_796,In_4051,In_4862);
nand U797 (N_797,In_1565,In_1050);
xnor U798 (N_798,In_2594,In_3926);
nor U799 (N_799,In_4184,In_2490);
xor U800 (N_800,In_4641,In_2903);
and U801 (N_801,In_3492,In_2547);
nor U802 (N_802,In_618,In_4368);
nand U803 (N_803,In_1682,In_1783);
nand U804 (N_804,In_2837,In_289);
or U805 (N_805,In_843,In_4006);
xor U806 (N_806,In_736,In_4527);
nand U807 (N_807,In_3177,In_3616);
and U808 (N_808,In_920,In_511);
nand U809 (N_809,In_1526,In_4162);
or U810 (N_810,In_98,In_2553);
and U811 (N_811,In_76,In_1913);
nand U812 (N_812,In_4879,In_1357);
or U813 (N_813,In_1918,In_4087);
xor U814 (N_814,In_3262,In_2934);
or U815 (N_815,In_1999,In_4314);
and U816 (N_816,In_3592,In_4961);
nand U817 (N_817,In_3398,In_767);
and U818 (N_818,In_1034,In_918);
nand U819 (N_819,In_3141,In_395);
and U820 (N_820,In_4581,In_2881);
or U821 (N_821,In_1056,In_4851);
or U822 (N_822,In_4972,In_1405);
and U823 (N_823,In_2715,In_4871);
nor U824 (N_824,In_4855,In_2077);
or U825 (N_825,In_925,In_1390);
xnor U826 (N_826,In_2454,In_2230);
or U827 (N_827,In_3784,In_1642);
nand U828 (N_828,In_3320,In_3561);
or U829 (N_829,In_1606,In_2733);
nand U830 (N_830,In_4795,In_4362);
or U831 (N_831,In_177,In_4399);
nor U832 (N_832,In_1633,In_3455);
nor U833 (N_833,In_4683,In_3655);
nand U834 (N_834,In_1167,In_1773);
and U835 (N_835,In_1048,In_4750);
or U836 (N_836,In_835,In_1915);
xor U837 (N_837,In_4645,In_2453);
nor U838 (N_838,In_2389,In_1095);
nand U839 (N_839,In_823,In_2878);
and U840 (N_840,In_2627,In_2000);
or U841 (N_841,In_1087,In_4716);
or U842 (N_842,In_4370,In_3362);
and U843 (N_843,In_4012,In_3772);
xnor U844 (N_844,In_2808,In_3118);
nand U845 (N_845,In_723,In_515);
and U846 (N_846,In_1523,In_4951);
or U847 (N_847,In_1027,In_3712);
xor U848 (N_848,In_1432,In_1022);
or U849 (N_849,In_3573,In_2549);
or U850 (N_850,In_4640,In_2322);
or U851 (N_851,In_862,In_4664);
xor U852 (N_852,In_2561,In_4486);
xor U853 (N_853,In_1672,In_959);
nor U854 (N_854,In_4059,In_1180);
nor U855 (N_855,In_1328,In_4944);
nand U856 (N_856,In_477,In_201);
nor U857 (N_857,In_3992,In_4416);
and U858 (N_858,In_1156,In_659);
nor U859 (N_859,In_2652,In_4796);
or U860 (N_860,In_2628,In_784);
or U861 (N_861,In_589,In_4223);
or U862 (N_862,In_3749,In_1009);
xnor U863 (N_863,In_2438,In_912);
xnor U864 (N_864,In_1412,In_2433);
nand U865 (N_865,In_2458,In_4779);
xor U866 (N_866,In_4502,In_4144);
and U867 (N_867,In_4192,In_3218);
and U868 (N_868,In_4083,In_3402);
xnor U869 (N_869,In_4395,In_3603);
or U870 (N_870,In_385,In_3160);
or U871 (N_871,In_643,In_4603);
or U872 (N_872,In_37,In_1938);
nor U873 (N_873,In_3290,In_77);
nor U874 (N_874,In_1727,In_1977);
nand U875 (N_875,In_587,In_4633);
xor U876 (N_876,In_4463,In_4456);
nand U877 (N_877,In_2473,In_2921);
and U878 (N_878,In_3355,In_448);
xor U879 (N_879,In_2463,In_3776);
or U880 (N_880,In_2055,In_842);
or U881 (N_881,In_306,In_2563);
and U882 (N_882,In_2550,In_769);
nand U883 (N_883,In_2966,In_4385);
and U884 (N_884,In_1584,In_3702);
nand U885 (N_885,In_3775,In_4824);
xnor U886 (N_886,In_1171,In_662);
and U887 (N_887,In_2777,In_2102);
and U888 (N_888,In_492,In_2294);
or U889 (N_889,In_191,In_1305);
nor U890 (N_890,In_3874,In_4031);
xor U891 (N_891,In_2496,In_297);
nand U892 (N_892,In_4277,In_3074);
xor U893 (N_893,In_2341,In_3003);
nand U894 (N_894,In_4801,In_4741);
or U895 (N_895,In_2176,In_4988);
nor U896 (N_896,In_2240,In_2744);
or U897 (N_897,In_247,In_2807);
nor U898 (N_898,In_1869,In_4544);
and U899 (N_899,In_4210,In_4560);
xor U900 (N_900,In_185,In_4218);
and U901 (N_901,In_3112,In_3995);
xnor U902 (N_902,In_1663,In_4211);
nor U903 (N_903,In_4616,In_4008);
xor U904 (N_904,In_4909,In_4088);
or U905 (N_905,In_458,In_4878);
nand U906 (N_906,In_3927,In_1680);
and U907 (N_907,In_107,In_3591);
nor U908 (N_908,In_2925,In_2686);
or U909 (N_909,In_1448,In_758);
and U910 (N_910,In_326,In_4249);
nand U911 (N_911,In_2167,In_2838);
nor U912 (N_912,In_4206,In_381);
or U913 (N_913,In_1109,In_128);
or U914 (N_914,In_3096,In_4392);
or U915 (N_915,In_649,In_3157);
nand U916 (N_916,In_1197,In_263);
or U917 (N_917,In_413,In_1297);
or U918 (N_918,In_4580,In_2361);
and U919 (N_919,In_502,In_3226);
nor U920 (N_920,In_4939,In_2511);
nor U921 (N_921,In_207,In_2506);
nor U922 (N_922,In_3382,In_4813);
nor U923 (N_923,In_4036,In_996);
or U924 (N_924,In_945,In_1029);
nor U925 (N_925,In_318,In_1954);
nand U926 (N_926,In_3006,In_549);
nor U927 (N_927,In_553,In_3870);
and U928 (N_928,In_4195,In_97);
nor U929 (N_929,In_3507,In_3007);
nand U930 (N_930,In_2172,In_2332);
xor U931 (N_931,In_3779,In_2376);
nand U932 (N_932,In_52,In_4355);
or U933 (N_933,In_3023,In_1123);
and U934 (N_934,In_2636,In_3341);
xnor U935 (N_935,In_4079,In_3430);
xnor U936 (N_936,In_1889,In_2940);
and U937 (N_937,In_3159,In_3720);
and U938 (N_938,In_1172,In_3821);
xnor U939 (N_939,In_2535,In_2943);
and U940 (N_940,In_917,In_772);
nand U941 (N_941,In_365,In_559);
nor U942 (N_942,In_3824,In_61);
nor U943 (N_943,In_1112,In_4566);
and U944 (N_944,In_1503,In_1014);
nand U945 (N_945,In_1793,In_144);
nor U946 (N_946,In_2610,In_1165);
xnor U947 (N_947,In_2844,In_1250);
nand U948 (N_948,In_277,In_955);
nand U949 (N_949,In_941,In_1806);
nor U950 (N_950,In_4837,In_1750);
nand U951 (N_951,In_523,In_3650);
or U952 (N_952,In_4219,In_1414);
or U953 (N_953,In_3175,In_4957);
xor U954 (N_954,In_4817,In_2280);
or U955 (N_955,In_2953,In_2159);
and U956 (N_956,In_2568,In_4113);
nor U957 (N_957,In_1886,In_99);
and U958 (N_958,In_3793,In_4731);
or U959 (N_959,In_2577,In_230);
nor U960 (N_960,In_4107,In_3239);
nand U961 (N_961,In_4709,In_353);
xor U962 (N_962,In_745,In_344);
nor U963 (N_963,In_2972,In_596);
or U964 (N_964,In_3557,In_1483);
and U965 (N_965,In_4937,In_590);
and U966 (N_966,In_3050,In_4118);
nor U967 (N_967,In_1287,In_1379);
nor U968 (N_968,In_2629,In_2742);
nand U969 (N_969,In_1767,In_1374);
xnor U970 (N_970,In_1151,In_4291);
nor U971 (N_971,In_4585,In_1545);
xor U972 (N_972,In_3106,In_4492);
or U973 (N_973,In_2607,In_3152);
xor U974 (N_974,In_2460,In_4315);
nor U975 (N_975,In_498,In_2936);
xor U976 (N_976,In_293,In_946);
or U977 (N_977,In_3963,In_1550);
nor U978 (N_978,In_1556,In_520);
nor U979 (N_979,In_1867,In_4330);
and U980 (N_980,In_4081,In_3056);
and U981 (N_981,In_1487,In_4637);
or U982 (N_982,In_1509,In_3354);
nor U983 (N_983,In_3153,In_4091);
or U984 (N_984,In_3993,In_4287);
or U985 (N_985,In_3244,In_4462);
xnor U986 (N_986,In_2189,In_1431);
nor U987 (N_987,In_1971,In_1667);
nand U988 (N_988,In_1906,In_3028);
or U989 (N_989,In_377,In_2416);
and U990 (N_990,In_3918,In_4589);
and U991 (N_991,In_60,In_3942);
nor U992 (N_992,In_1450,In_792);
nand U993 (N_993,In_2978,In_4718);
nor U994 (N_994,In_471,In_3932);
nand U995 (N_995,In_1140,In_4865);
nor U996 (N_996,In_3308,In_2580);
or U997 (N_997,In_38,In_4775);
or U998 (N_998,In_2004,In_3627);
xnor U999 (N_999,In_418,In_2035);
and U1000 (N_1000,In_2661,In_1508);
nor U1001 (N_1001,In_2793,In_1872);
xnor U1002 (N_1002,In_92,In_214);
nor U1003 (N_1003,In_2492,In_3260);
nor U1004 (N_1004,In_410,In_3949);
nand U1005 (N_1005,In_4284,In_246);
or U1006 (N_1006,In_3301,In_2219);
nor U1007 (N_1007,In_3741,In_3411);
xor U1008 (N_1008,In_512,In_4840);
xnor U1009 (N_1009,In_2717,In_397);
xnor U1010 (N_1010,In_2139,In_3318);
nand U1011 (N_1011,In_290,In_3282);
nand U1012 (N_1012,In_1648,In_2049);
or U1013 (N_1013,In_3154,In_2651);
xor U1014 (N_1014,In_833,In_2415);
or U1015 (N_1015,In_677,In_762);
and U1016 (N_1016,In_2071,In_4090);
and U1017 (N_1017,In_2477,In_2527);
nor U1018 (N_1018,In_4514,In_4619);
nor U1019 (N_1019,In_3767,In_4394);
xnor U1020 (N_1020,In_1435,In_1996);
or U1021 (N_1021,In_679,In_2402);
and U1022 (N_1022,In_2806,In_4827);
or U1023 (N_1023,In_2824,In_1440);
nand U1024 (N_1024,In_1406,In_770);
xnor U1025 (N_1025,In_4694,In_470);
nand U1026 (N_1026,In_2823,In_3233);
or U1027 (N_1027,In_1711,In_1184);
nor U1028 (N_1028,In_614,In_420);
and U1029 (N_1029,In_2873,In_1724);
nand U1030 (N_1030,In_1535,In_2111);
and U1031 (N_1031,In_2804,In_3072);
nor U1032 (N_1032,In_2896,In_4902);
xnor U1033 (N_1033,In_3163,In_68);
xnor U1034 (N_1034,In_2692,In_3264);
nand U1035 (N_1035,In_2641,In_979);
or U1036 (N_1036,In_879,In_4825);
nand U1037 (N_1037,In_681,In_612);
nor U1038 (N_1038,In_3608,In_4806);
or U1039 (N_1039,In_517,In_3714);
or U1040 (N_1040,In_3537,In_1978);
nand U1041 (N_1041,In_4027,In_4139);
nand U1042 (N_1042,In_2400,In_3546);
and U1043 (N_1043,In_3678,In_3025);
xnor U1044 (N_1044,In_1592,In_4153);
nand U1045 (N_1045,In_388,In_2889);
xor U1046 (N_1046,In_871,In_3681);
and U1047 (N_1047,In_335,In_374);
or U1048 (N_1048,In_4444,In_1230);
xor U1049 (N_1049,In_1159,In_2657);
xor U1050 (N_1050,In_1396,In_2880);
and U1051 (N_1051,In_34,In_2270);
and U1052 (N_1052,In_2578,In_3041);
or U1053 (N_1053,In_2712,In_2994);
or U1054 (N_1054,In_3739,In_3342);
xnor U1055 (N_1055,In_4759,In_3586);
nor U1056 (N_1056,In_108,In_2367);
and U1057 (N_1057,In_671,In_3197);
and U1058 (N_1058,In_4517,In_2979);
nand U1059 (N_1059,In_3107,In_2256);
and U1060 (N_1060,In_3773,In_4432);
and U1061 (N_1061,In_2101,In_3433);
nor U1062 (N_1062,In_1174,In_500);
and U1063 (N_1063,In_4446,In_2573);
xnor U1064 (N_1064,In_2911,In_168);
or U1065 (N_1065,In_4649,In_4312);
and U1066 (N_1066,In_220,In_1204);
xor U1067 (N_1067,In_4834,In_3461);
and U1068 (N_1068,In_3800,In_3754);
nor U1069 (N_1069,In_3683,In_2313);
nand U1070 (N_1070,In_704,In_3531);
nand U1071 (N_1071,In_4997,In_3190);
nor U1072 (N_1072,In_1385,In_4934);
nor U1073 (N_1073,In_1926,In_4213);
or U1074 (N_1074,In_2973,In_2286);
nor U1075 (N_1075,In_1476,In_2867);
nor U1076 (N_1076,In_4436,In_2238);
and U1077 (N_1077,In_1966,In_176);
nand U1078 (N_1078,In_4744,In_30);
nor U1079 (N_1079,In_865,In_4654);
nor U1080 (N_1080,In_4233,In_1877);
xor U1081 (N_1081,In_2585,In_1673);
and U1082 (N_1082,In_592,In_2599);
xor U1083 (N_1083,In_2687,In_1809);
xnor U1084 (N_1084,In_4360,In_1386);
nor U1085 (N_1085,In_1035,In_4874);
and U1086 (N_1086,In_1017,In_3432);
nand U1087 (N_1087,In_3210,In_2396);
nand U1088 (N_1088,In_4358,In_3511);
and U1089 (N_1089,In_1596,In_3612);
or U1090 (N_1090,In_1796,In_872);
or U1091 (N_1091,In_2254,In_4319);
nand U1092 (N_1092,In_4256,In_451);
nand U1093 (N_1093,In_2482,In_3230);
or U1094 (N_1094,In_1290,In_1937);
nand U1095 (N_1095,In_3059,In_3281);
nor U1096 (N_1096,In_875,In_4762);
xor U1097 (N_1097,In_646,In_4733);
or U1098 (N_1098,In_3829,In_1162);
nand U1099 (N_1099,In_2211,In_3953);
nand U1100 (N_1100,In_3252,In_800);
nand U1101 (N_1101,In_2328,In_449);
nor U1102 (N_1102,In_3958,In_2671);
nor U1103 (N_1103,In_3093,In_1329);
and U1104 (N_1104,In_597,In_1833);
or U1105 (N_1105,In_755,In_4048);
or U1106 (N_1106,In_4484,In_4684);
nand U1107 (N_1107,In_2998,In_2597);
xor U1108 (N_1108,In_3187,In_2315);
or U1109 (N_1109,In_1323,In_3016);
or U1110 (N_1110,In_3732,In_1587);
nor U1111 (N_1111,In_3961,In_3915);
and U1112 (N_1112,In_3794,In_4019);
and U1113 (N_1113,In_3651,In_2163);
nor U1114 (N_1114,In_935,In_1777);
or U1115 (N_1115,In_3236,In_4457);
nor U1116 (N_1116,In_3049,In_2025);
and U1117 (N_1117,In_887,In_2083);
or U1118 (N_1118,In_3983,In_1376);
nor U1119 (N_1119,In_854,In_3851);
nor U1120 (N_1120,In_845,In_4588);
and U1121 (N_1121,In_3481,In_3988);
and U1122 (N_1122,In_4424,In_4576);
xnor U1123 (N_1123,In_3321,In_4915);
xnor U1124 (N_1124,In_3314,In_1586);
nor U1125 (N_1125,In_3939,In_2233);
nor U1126 (N_1126,In_2710,In_2829);
or U1127 (N_1127,In_4169,In_1976);
nor U1128 (N_1128,In_2755,In_3189);
nand U1129 (N_1129,In_3228,In_703);
or U1130 (N_1130,In_1416,In_2930);
nand U1131 (N_1131,In_3265,In_2022);
or U1132 (N_1132,In_450,In_1686);
and U1133 (N_1133,In_4528,In_4126);
xor U1134 (N_1134,In_2436,In_3271);
and U1135 (N_1135,In_2151,In_4109);
or U1136 (N_1136,In_2365,In_1020);
nor U1137 (N_1137,In_3227,In_3498);
nand U1138 (N_1138,In_674,In_2948);
or U1139 (N_1139,In_1389,In_4926);
nor U1140 (N_1140,In_1760,In_4629);
xor U1141 (N_1141,In_1998,In_3404);
nor U1142 (N_1142,In_4970,In_109);
nand U1143 (N_1143,In_405,In_806);
or U1144 (N_1144,In_2541,In_4739);
nor U1145 (N_1145,In_1819,In_2863);
and U1146 (N_1146,In_2831,In_3386);
or U1147 (N_1147,In_2346,In_939);
xor U1148 (N_1148,In_2181,In_3549);
and U1149 (N_1149,In_1536,In_898);
xnor U1150 (N_1150,In_1016,In_1008);
or U1151 (N_1151,In_270,In_4805);
or U1152 (N_1152,In_4342,In_3759);
nor U1153 (N_1153,In_3178,In_209);
nor U1154 (N_1154,In_2716,In_2245);
and U1155 (N_1155,In_3677,In_4461);
and U1156 (N_1156,In_1254,In_4017);
nor U1157 (N_1157,In_1533,In_3174);
nor U1158 (N_1158,In_3528,In_4803);
xor U1159 (N_1159,In_3038,In_3347);
and U1160 (N_1160,In_2962,In_2292);
nor U1161 (N_1161,In_4985,In_1626);
or U1162 (N_1162,In_2009,In_1482);
and U1163 (N_1163,In_4959,In_3766);
nor U1164 (N_1164,In_841,In_830);
nand U1165 (N_1165,In_1175,In_2006);
xor U1166 (N_1166,In_1951,In_3705);
xor U1167 (N_1167,In_4690,In_3871);
or U1168 (N_1168,In_1813,In_1543);
or U1169 (N_1169,In_2180,In_2068);
nor U1170 (N_1170,In_1551,In_2105);
or U1171 (N_1171,In_675,In_1408);
xnor U1172 (N_1172,In_886,In_21);
xnor U1173 (N_1173,In_2872,In_2281);
or U1174 (N_1174,In_1286,In_352);
nor U1175 (N_1175,In_2309,In_3490);
or U1176 (N_1176,In_958,In_3839);
xnor U1177 (N_1177,In_4493,In_578);
and U1178 (N_1178,In_582,In_4978);
nor U1179 (N_1179,In_3165,In_1395);
or U1180 (N_1180,In_595,In_2876);
xor U1181 (N_1181,In_4058,In_636);
or U1182 (N_1182,In_2694,In_206);
and U1183 (N_1183,In_1339,In_2907);
and U1184 (N_1184,In_813,In_2041);
and U1185 (N_1185,In_4337,In_2536);
xor U1186 (N_1186,In_357,In_3504);
or U1187 (N_1187,In_4367,In_3792);
and U1188 (N_1188,In_4858,In_3742);
nand U1189 (N_1189,In_2171,In_1494);
xor U1190 (N_1190,In_4523,In_1823);
and U1191 (N_1191,In_2098,In_4593);
xnor U1192 (N_1192,In_129,In_3060);
and U1193 (N_1193,In_1307,In_1341);
nor U1194 (N_1194,In_602,In_3164);
nand U1195 (N_1195,In_2622,In_2127);
xor U1196 (N_1196,In_2251,In_4845);
nor U1197 (N_1197,In_1086,In_1348);
or U1198 (N_1198,In_847,In_4529);
and U1199 (N_1199,In_863,In_4168);
xnor U1200 (N_1200,In_4571,In_1860);
or U1201 (N_1201,In_262,In_2871);
nor U1202 (N_1202,In_839,In_986);
or U1203 (N_1203,In_16,In_2737);
and U1204 (N_1204,In_75,In_2036);
and U1205 (N_1205,In_133,In_1192);
or U1206 (N_1206,In_860,In_1849);
nand U1207 (N_1207,In_2778,In_433);
xor U1208 (N_1208,In_1983,In_456);
xor U1209 (N_1209,In_3085,In_3487);
nor U1210 (N_1210,In_1785,In_2799);
nor U1211 (N_1211,In_2193,In_3925);
xor U1212 (N_1212,In_1010,In_4442);
and U1213 (N_1213,In_2497,In_1560);
nor U1214 (N_1214,In_2693,In_1373);
and U1215 (N_1215,In_965,In_3968);
nand U1216 (N_1216,In_1265,In_4325);
or U1217 (N_1217,In_2834,In_3737);
nand U1218 (N_1218,In_457,In_4535);
xnor U1219 (N_1219,In_2866,In_469);
and U1220 (N_1220,In_3002,In_1398);
or U1221 (N_1221,In_2255,In_3532);
xor U1222 (N_1222,In_1434,In_3771);
and U1223 (N_1223,In_991,In_237);
nand U1224 (N_1224,In_798,In_3463);
xor U1225 (N_1225,In_56,In_1980);
xor U1226 (N_1226,In_2551,In_1738);
nand U1227 (N_1227,In_1104,In_4101);
nor U1228 (N_1228,In_1154,In_3280);
and U1229 (N_1229,In_2816,In_858);
or U1230 (N_1230,In_3067,In_4023);
or U1231 (N_1231,In_2086,In_785);
or U1232 (N_1232,In_1949,In_1660);
and U1233 (N_1233,In_2326,In_1415);
nand U1234 (N_1234,In_4185,In_4541);
and U1235 (N_1235,In_4408,In_3350);
nand U1236 (N_1236,In_850,In_786);
or U1237 (N_1237,In_3636,In_337);
or U1238 (N_1238,In_286,In_223);
or U1239 (N_1239,In_2590,In_4635);
and U1240 (N_1240,In_402,In_2723);
nand U1241 (N_1241,In_2809,In_3299);
and U1242 (N_1242,In_2386,In_3948);
or U1243 (N_1243,In_2095,In_1002);
or U1244 (N_1244,In_530,In_1229);
and U1245 (N_1245,In_2331,In_3861);
and U1246 (N_1246,In_1291,In_3209);
nor U1247 (N_1247,In_4572,In_4435);
and U1248 (N_1248,In_4938,In_2320);
and U1249 (N_1249,In_1124,In_2204);
and U1250 (N_1250,In_1859,In_694);
or U1251 (N_1251,In_2448,In_4804);
and U1252 (N_1252,In_4757,In_501);
nor U1253 (N_1253,In_3484,In_4967);
xnor U1254 (N_1254,In_2177,In_3442);
and U1255 (N_1255,In_3033,In_138);
and U1256 (N_1256,In_4449,In_3405);
or U1257 (N_1257,In_2122,In_4501);
or U1258 (N_1258,In_3179,In_2399);
or U1259 (N_1259,In_1429,In_3858);
xnor U1260 (N_1260,In_287,In_1656);
nor U1261 (N_1261,In_4539,In_2003);
xor U1262 (N_1262,In_931,In_2530);
nor U1263 (N_1263,In_695,In_864);
and U1264 (N_1264,In_972,In_1982);
xnor U1265 (N_1265,In_136,In_1413);
and U1266 (N_1266,In_4138,In_2583);
xor U1267 (N_1267,In_4980,In_115);
and U1268 (N_1268,In_4670,In_2591);
nand U1269 (N_1269,In_2278,In_1391);
and U1270 (N_1270,In_3274,In_356);
and U1271 (N_1271,In_4480,In_3680);
xor U1272 (N_1272,In_3696,In_2200);
and U1273 (N_1273,In_3744,In_1083);
xnor U1274 (N_1274,In_2450,In_2264);
and U1275 (N_1275,In_3445,In_1081);
nand U1276 (N_1276,In_4387,In_2708);
and U1277 (N_1277,In_95,In_4904);
nor U1278 (N_1278,In_1141,In_3524);
xnor U1279 (N_1279,In_1274,In_3955);
nand U1280 (N_1280,In_330,In_2451);
xnor U1281 (N_1281,In_3283,In_302);
nor U1282 (N_1282,In_730,In_3910);
and U1283 (N_1283,In_619,In_4740);
and U1284 (N_1284,In_4789,In_4521);
and U1285 (N_1285,In_4669,In_3997);
and U1286 (N_1286,In_4111,In_2905);
xor U1287 (N_1287,In_1712,In_1377);
and U1288 (N_1288,In_2802,In_3127);
and U1289 (N_1289,In_3980,In_2556);
nor U1290 (N_1290,In_4124,In_4022);
and U1291 (N_1291,In_4267,In_4014);
and U1292 (N_1292,In_2057,In_1824);
nor U1293 (N_1293,In_1611,In_1647);
nor U1294 (N_1294,In_509,In_1331);
or U1295 (N_1295,In_1439,In_69);
xor U1296 (N_1296,In_3936,In_3275);
and U1297 (N_1297,In_3787,In_116);
nand U1298 (N_1298,In_2480,In_2695);
nor U1299 (N_1299,In_4979,In_2714);
and U1300 (N_1300,In_4623,In_4552);
nor U1301 (N_1301,In_125,In_3589);
nor U1302 (N_1302,In_3805,In_2028);
or U1303 (N_1303,In_4607,In_2428);
xor U1304 (N_1304,In_2407,In_1865);
nand U1305 (N_1305,In_81,In_4600);
xnor U1306 (N_1306,In_101,In_3520);
or U1307 (N_1307,In_4912,In_1659);
and U1308 (N_1308,In_4142,In_2229);
nand U1309 (N_1309,In_973,In_1729);
nand U1310 (N_1310,In_3105,In_3076);
nand U1311 (N_1311,In_190,In_2768);
nor U1312 (N_1312,In_189,In_1848);
or U1313 (N_1313,In_2941,In_2780);
xnor U1314 (N_1314,In_1121,In_1797);
nand U1315 (N_1315,In_1779,In_2702);
or U1316 (N_1316,In_309,In_2383);
xnor U1317 (N_1317,In_4041,In_1700);
nor U1318 (N_1318,In_3893,In_1683);
xor U1319 (N_1319,In_573,In_4682);
nand U1320 (N_1320,In_2384,In_2999);
nor U1321 (N_1321,In_926,In_1770);
nor U1322 (N_1322,In_2980,In_3647);
nand U1323 (N_1323,In_1318,In_2554);
nor U1324 (N_1324,In_2971,In_4472);
xnor U1325 (N_1325,In_3891,In_454);
and U1326 (N_1326,In_4644,In_3090);
or U1327 (N_1327,In_2555,In_4167);
xor U1328 (N_1328,In_2291,In_4115);
and U1329 (N_1329,In_4215,In_3409);
nor U1330 (N_1330,In_1157,In_2425);
nand U1331 (N_1331,In_607,In_2574);
and U1332 (N_1332,In_746,In_3173);
or U1333 (N_1333,In_4798,In_1444);
and U1334 (N_1334,In_2882,In_1905);
or U1335 (N_1335,In_358,In_359);
xnor U1336 (N_1336,In_442,In_661);
nor U1337 (N_1337,In_4922,In_3569);
xor U1338 (N_1338,In_4819,In_339);
nor U1339 (N_1339,In_4146,In_117);
or U1340 (N_1340,In_3748,In_3530);
nor U1341 (N_1341,In_1594,In_2722);
nand U1342 (N_1342,In_2461,In_319);
or U1343 (N_1343,In_4357,In_3361);
or U1344 (N_1344,In_1883,In_2931);
xnor U1345 (N_1345,In_4699,In_1832);
nor U1346 (N_1346,In_1780,In_3351);
nor U1347 (N_1347,In_4464,In_2301);
and U1348 (N_1348,In_4467,In_17);
or U1349 (N_1349,In_4261,In_1759);
or U1350 (N_1350,In_4379,In_2975);
or U1351 (N_1351,In_642,In_4547);
or U1352 (N_1352,In_1049,In_2048);
xor U1353 (N_1353,In_4478,In_3171);
nand U1354 (N_1354,In_2891,In_4942);
or U1355 (N_1355,In_2340,In_2135);
and U1356 (N_1356,In_3862,In_4916);
or U1357 (N_1357,In_3697,In_4549);
or U1358 (N_1358,In_2519,In_3284);
xor U1359 (N_1359,In_2096,In_4838);
nor U1360 (N_1360,In_1530,In_4921);
or U1361 (N_1361,In_4339,In_1063);
nand U1362 (N_1362,In_1669,In_2729);
xnor U1363 (N_1363,In_2182,In_3594);
nor U1364 (N_1364,In_4867,In_4886);
nor U1365 (N_1365,In_1579,In_811);
nor U1366 (N_1366,In_256,In_4179);
nand U1367 (N_1367,In_3894,In_4476);
xnor U1368 (N_1368,In_2225,In_1025);
or U1369 (N_1369,In_3456,In_3225);
nor U1370 (N_1370,In_533,In_3758);
and U1371 (N_1371,In_1161,In_2965);
xnor U1372 (N_1372,In_2356,In_771);
or U1373 (N_1373,In_2720,In_4667);
nor U1374 (N_1374,In_1354,In_2679);
nand U1375 (N_1375,In_2796,In_3422);
and U1376 (N_1376,In_1215,In_3935);
or U1377 (N_1377,In_2961,In_2531);
or U1378 (N_1378,In_2008,In_2330);
and U1379 (N_1379,In_3830,In_3387);
xnor U1380 (N_1380,In_1134,In_3019);
xor U1381 (N_1381,In_2108,In_970);
and U1382 (N_1382,In_3278,In_537);
nor U1383 (N_1383,In_379,In_39);
or U1384 (N_1384,In_591,In_1707);
xor U1385 (N_1385,In_885,In_1486);
and U1386 (N_1386,In_241,In_2586);
nand U1387 (N_1387,In_2874,In_2261);
xor U1388 (N_1388,In_4106,In_1420);
xnor U1389 (N_1389,In_1474,In_2798);
xor U1390 (N_1390,In_4011,In_4097);
or U1391 (N_1391,In_1359,In_4609);
and U1392 (N_1392,In_3907,In_1645);
nand U1393 (N_1393,In_4398,In_3356);
or U1394 (N_1394,In_1372,In_3711);
nor U1395 (N_1395,In_3990,In_252);
nand U1396 (N_1396,In_1145,In_2444);
or U1397 (N_1397,In_1568,In_3790);
and U1398 (N_1398,In_576,In_4956);
nand U1399 (N_1399,In_3192,In_4283);
or U1400 (N_1400,In_1599,In_1986);
and U1401 (N_1401,In_308,In_2545);
nand U1402 (N_1402,In_3578,In_341);
or U1403 (N_1403,In_3267,In_195);
nor U1404 (N_1404,In_143,In_3622);
or U1405 (N_1405,In_300,In_1226);
and U1406 (N_1406,In_2630,In_3855);
nand U1407 (N_1407,In_1640,In_1967);
or U1408 (N_1408,In_3920,In_3053);
nor U1409 (N_1409,In_2408,In_4068);
nor U1410 (N_1410,In_3193,In_2633);
or U1411 (N_1411,In_3058,In_2500);
or U1412 (N_1412,In_4030,In_4285);
nand U1413 (N_1413,In_84,In_4507);
xnor U1414 (N_1414,In_2524,In_4494);
xnor U1415 (N_1415,In_4857,In_336);
nor U1416 (N_1416,In_4999,In_1939);
and U1417 (N_1417,In_380,In_59);
nand U1418 (N_1418,In_3399,In_1370);
xnor U1419 (N_1419,In_1958,In_4075);
and U1420 (N_1420,In_1512,In_4526);
xnor U1421 (N_1421,In_3703,In_4437);
nor U1422 (N_1422,In_4870,In_3425);
nor U1423 (N_1423,In_668,In_4653);
xnor U1424 (N_1424,In_505,In_1484);
or U1425 (N_1425,In_3882,In_2298);
xor U1426 (N_1426,In_4650,In_1044);
xor U1427 (N_1427,In_4522,In_141);
or U1428 (N_1428,In_4419,In_1355);
nand U1429 (N_1429,In_3881,In_2045);
xor U1430 (N_1430,In_3039,In_3722);
nor U1431 (N_1431,In_585,In_4102);
nor U1432 (N_1432,In_930,In_2072);
and U1433 (N_1433,In_4190,In_4013);
xnor U1434 (N_1434,In_1472,In_4601);
or U1435 (N_1435,In_2173,In_1054);
and U1436 (N_1436,In_1635,In_3036);
or U1437 (N_1437,In_4202,In_1916);
nor U1438 (N_1438,In_827,In_4422);
nand U1439 (N_1439,In_660,In_856);
or U1440 (N_1440,In_3662,In_275);
and U1441 (N_1441,In_2852,In_3947);
or U1442 (N_1442,In_1628,In_1481);
nand U1443 (N_1443,In_1687,In_3840);
nor U1444 (N_1444,In_2917,In_1705);
xor U1445 (N_1445,In_4086,In_2093);
nor U1446 (N_1446,In_2833,In_2792);
xnor U1447 (N_1447,In_1840,In_2184);
nand U1448 (N_1448,In_2893,In_3628);
nand U1449 (N_1449,In_1688,In_1106);
xor U1450 (N_1450,In_2613,In_4278);
xnor U1451 (N_1451,In_1479,In_4794);
xor U1452 (N_1452,In_3596,In_4397);
or U1453 (N_1453,In_3024,In_2785);
nand U1454 (N_1454,In_2769,In_1981);
or U1455 (N_1455,In_940,In_2840);
nor U1456 (N_1456,In_3717,In_2539);
nor U1457 (N_1457,In_4525,In_1934);
nor U1458 (N_1458,In_624,In_1864);
or U1459 (N_1459,In_3704,In_889);
or U1460 (N_1460,In_1127,In_4599);
nor U1461 (N_1461,In_3071,In_325);
nand U1462 (N_1462,In_3366,In_2149);
nor U1463 (N_1463,In_3502,In_1600);
xor U1464 (N_1464,In_3109,In_652);
or U1465 (N_1465,In_2268,In_1388);
nand U1466 (N_1466,In_279,In_3982);
xor U1467 (N_1467,In_4958,In_4029);
nand U1468 (N_1468,In_4698,In_2841);
and U1469 (N_1469,In_1085,In_1223);
xnor U1470 (N_1470,In_3259,In_2932);
xor U1471 (N_1471,In_239,In_2279);
xnor U1472 (N_1472,In_1907,In_123);
nor U1473 (N_1473,In_4205,In_3719);
nor U1474 (N_1474,In_613,In_212);
nand U1475 (N_1475,In_2775,In_732);
nor U1476 (N_1476,In_428,In_1093);
or U1477 (N_1477,In_3037,In_3258);
xnor U1478 (N_1478,In_4371,In_2942);
nand U1479 (N_1479,In_2540,In_4778);
and U1480 (N_1480,In_2109,In_3964);
xnor U1481 (N_1481,In_577,In_4175);
nand U1482 (N_1482,In_4508,In_4636);
and U1483 (N_1483,In_2606,In_3952);
nand U1484 (N_1484,In_1061,In_3435);
xnor U1485 (N_1485,In_4229,In_3970);
or U1486 (N_1486,In_2164,In_2237);
nor U1487 (N_1487,In_2659,In_4306);
nand U1488 (N_1488,In_4888,In_3774);
or U1489 (N_1489,In_1737,In_2771);
nor U1490 (N_1490,In_3609,In_1024);
or U1491 (N_1491,In_3661,In_929);
nand U1492 (N_1492,In_3368,In_3761);
and U1493 (N_1493,In_742,In_2631);
and U1494 (N_1494,In_445,In_4540);
xnor U1495 (N_1495,In_966,In_3575);
and U1496 (N_1496,In_1404,In_1189);
nand U1497 (N_1497,In_4776,In_198);
xnor U1498 (N_1498,In_4615,In_4263);
nand U1499 (N_1499,In_4488,In_4701);
and U1500 (N_1500,In_4760,In_4856);
xnor U1501 (N_1501,In_4940,In_3064);
nand U1502 (N_1502,In_3674,In_4946);
or U1503 (N_1503,In_894,In_4720);
nand U1504 (N_1504,In_1190,In_307);
xor U1505 (N_1505,In_2650,In_735);
xor U1506 (N_1506,In_4335,In_2065);
xor U1507 (N_1507,In_3916,In_1513);
or U1508 (N_1508,In_4331,In_124);
and U1509 (N_1509,In_2810,In_3020);
and U1510 (N_1510,In_1588,In_2593);
nand U1511 (N_1511,In_3658,In_1745);
nand U1512 (N_1512,In_4626,In_1456);
xor U1513 (N_1513,In_964,In_4383);
or U1514 (N_1514,In_2794,In_3464);
and U1515 (N_1515,In_4873,In_1067);
nand U1516 (N_1516,In_1202,In_2202);
and U1517 (N_1517,In_3777,In_4691);
nand U1518 (N_1518,In_2016,In_2063);
nor U1519 (N_1519,In_4567,In_3547);
nand U1520 (N_1520,In_519,In_3868);
nand U1521 (N_1521,In_3485,In_1782);
or U1522 (N_1522,In_4402,In_4177);
nor U1523 (N_1523,In_182,In_2368);
nand U1524 (N_1524,In_1816,In_235);
and U1525 (N_1525,In_825,In_3850);
and U1526 (N_1526,In_3692,In_1880);
or U1527 (N_1527,In_4618,In_857);
nand U1528 (N_1528,In_3497,In_3287);
and U1529 (N_1529,In_4810,In_3986);
nand U1530 (N_1530,In_2064,In_2538);
nand U1531 (N_1531,In_2559,In_2242);
or U1532 (N_1532,In_684,In_4722);
nand U1533 (N_1533,In_2765,In_3238);
nor U1534 (N_1534,In_2639,In_3022);
or U1535 (N_1535,In_2349,In_3371);
and U1536 (N_1536,In_571,In_4711);
or U1537 (N_1537,In_4729,In_3709);
or U1538 (N_1538,In_148,In_1878);
nand U1539 (N_1539,In_2449,In_3185);
nor U1540 (N_1540,In_1991,In_1304);
nor U1541 (N_1541,In_4573,In_1805);
xnor U1542 (N_1542,In_3657,In_4241);
or U1543 (N_1543,In_20,In_3905);
and U1544 (N_1544,In_3207,In_2336);
and U1545 (N_1545,In_4950,In_1312);
nor U1546 (N_1546,In_4758,In_1332);
and U1547 (N_1547,In_3216,In_482);
or U1548 (N_1548,In_3486,In_908);
xor U1549 (N_1549,In_4704,In_916);
nor U1550 (N_1550,In_3234,In_4543);
and U1551 (N_1551,In_1302,In_594);
xnor U1552 (N_1552,In_4850,In_799);
nor U1553 (N_1553,In_4854,In_4913);
nand U1554 (N_1554,In_4869,In_2761);
xor U1555 (N_1555,In_3571,In_969);
xnor U1556 (N_1556,In_3731,In_541);
or U1557 (N_1557,In_3890,In_1898);
xnor U1558 (N_1558,In_3346,In_4787);
nor U1559 (N_1559,In_2485,In_4792);
or U1560 (N_1560,In_1382,In_2305);
and U1561 (N_1561,In_1522,In_2901);
nor U1562 (N_1562,In_2419,In_3294);
and U1563 (N_1563,In_3806,In_3231);
and U1564 (N_1564,In_4973,In_928);
xor U1565 (N_1565,In_2850,In_74);
and U1566 (N_1566,In_87,In_529);
nand U1567 (N_1567,In_3903,In_1371);
nand U1568 (N_1568,In_4300,In_2343);
xnor U1569 (N_1569,In_3548,In_4863);
xnor U1570 (N_1570,In_3516,In_3536);
or U1571 (N_1571,In_4381,In_2104);
and U1572 (N_1572,In_2441,In_3826);
nand U1573 (N_1573,In_3901,In_181);
and U1574 (N_1574,In_3740,In_414);
or U1575 (N_1575,In_1309,In_333);
and U1576 (N_1576,In_3219,In_2909);
nand U1577 (N_1577,In_2915,In_3212);
nand U1578 (N_1578,In_149,In_173);
nand U1579 (N_1579,In_4816,In_2372);
xor U1580 (N_1580,In_4482,In_4652);
xor U1581 (N_1581,In_1940,In_2730);
nand U1582 (N_1582,In_460,In_2560);
and U1583 (N_1583,In_3353,In_4941);
and U1584 (N_1584,In_1337,In_1752);
or U1585 (N_1585,In_408,In_722);
nand U1586 (N_1586,In_1678,In_3940);
nand U1587 (N_1587,In_3126,In_3480);
or U1588 (N_1588,In_2904,In_4793);
nor U1589 (N_1589,In_1120,In_563);
nand U1590 (N_1590,In_1316,In_4639);
xnor U1591 (N_1591,In_2724,In_112);
or U1592 (N_1592,In_994,In_1542);
nand U1593 (N_1593,In_3945,In_2417);
nand U1594 (N_1594,In_430,In_4137);
nor U1595 (N_1595,In_4182,In_1662);
xnor U1596 (N_1596,In_3567,In_4037);
nor U1597 (N_1597,In_2981,In_2502);
xor U1598 (N_1598,In_2618,In_2137);
and U1599 (N_1599,In_4842,In_2);
nand U1600 (N_1600,In_809,In_2984);
xnor U1601 (N_1601,In_383,In_1578);
xor U1602 (N_1602,In_2746,In_4375);
xnor U1603 (N_1603,In_2581,In_1004);
and U1604 (N_1604,In_1525,In_3618);
xor U1605 (N_1605,In_866,In_558);
nand U1606 (N_1606,In_3764,In_3406);
nor U1607 (N_1607,In_3010,In_1549);
nand U1608 (N_1608,In_4656,In_2132);
or U1609 (N_1609,In_485,In_4007);
or U1610 (N_1610,In_689,In_4475);
and U1611 (N_1611,In_1702,In_3693);
nand U1612 (N_1612,In_2624,In_119);
nor U1613 (N_1613,In_635,In_4882);
and U1614 (N_1614,In_4584,In_140);
and U1615 (N_1615,In_4296,In_73);
nand U1616 (N_1616,In_686,In_2766);
xor U1617 (N_1617,In_713,In_2153);
nand U1618 (N_1618,In_4487,In_2774);
nor U1619 (N_1619,In_1158,In_3735);
nor U1620 (N_1620,In_2895,In_2027);
and U1621 (N_1621,In_4222,In_1710);
and U1622 (N_1622,In_166,In_1625);
or U1623 (N_1623,In_1899,In_3879);
or U1624 (N_1624,In_4592,In_3804);
and U1625 (N_1625,In_1942,In_881);
xnor U1626 (N_1626,In_2951,In_1956);
xor U1627 (N_1627,In_3898,In_1064);
nor U1628 (N_1628,In_2964,In_828);
nor U1629 (N_1629,In_1330,In_3313);
nor U1630 (N_1630,In_510,In_4311);
nor U1631 (N_1631,In_231,In_46);
and U1632 (N_1632,In_1970,In_1572);
nor U1633 (N_1633,In_1841,In_4125);
xnor U1634 (N_1634,In_3421,In_1671);
and U1635 (N_1635,In_947,In_3656);
and U1636 (N_1636,In_693,In_4892);
and U1637 (N_1637,In_949,In_2440);
nor U1638 (N_1638,In_556,In_2363);
or U1639 (N_1639,In_702,In_132);
nor U1640 (N_1640,In_4214,In_2677);
xor U1641 (N_1641,In_146,In_4271);
or U1642 (N_1642,In_1220,In_3241);
and U1643 (N_1643,In_4468,In_2997);
and U1644 (N_1644,In_2957,In_1827);
xnor U1645 (N_1645,In_4450,In_691);
nand U1646 (N_1646,In_3525,In_2954);
and U1647 (N_1647,In_1828,In_4557);
and U1648 (N_1648,In_2359,In_1273);
and U1649 (N_1649,In_744,In_1757);
and U1650 (N_1650,In_499,In_158);
xor U1651 (N_1651,In_4057,In_2865);
nand U1652 (N_1652,In_1076,In_4188);
xor U1653 (N_1653,In_4859,In_4914);
nand U1654 (N_1654,In_496,In_3723);
xor U1655 (N_1655,In_4844,In_463);
and U1656 (N_1656,In_3327,In_1194);
nand U1657 (N_1657,In_3393,In_3797);
nand U1658 (N_1658,In_3902,In_2494);
xor U1659 (N_1659,In_3752,In_1267);
or U1660 (N_1660,In_3673,In_3663);
and U1661 (N_1661,In_3120,In_4232);
xnor U1662 (N_1662,In_3852,In_990);
nor U1663 (N_1663,In_3358,In_2884);
and U1664 (N_1664,In_4327,In_3370);
nor U1665 (N_1665,In_1101,In_4591);
and U1666 (N_1666,In_4073,In_4971);
or U1667 (N_1667,In_834,In_2377);
nand U1668 (N_1668,In_2091,In_3574);
nor U1669 (N_1669,In_1854,In_1170);
and U1670 (N_1670,In_724,In_507);
nand U1671 (N_1671,In_1546,In_1015);
nor U1672 (N_1672,In_638,In_1179);
or U1673 (N_1673,In_1233,In_4200);
xor U1674 (N_1674,In_999,In_685);
or U1675 (N_1675,In_3554,In_4852);
nand U1676 (N_1676,In_1053,In_1227);
xor U1677 (N_1677,In_1417,In_2935);
and U1678 (N_1678,In_3482,In_1947);
nor U1679 (N_1679,In_4199,In_3416);
and U1680 (N_1680,In_1766,In_331);
and U1681 (N_1681,In_343,In_3796);
and U1682 (N_1682,In_1356,In_47);
xor U1683 (N_1683,In_4790,In_2205);
or U1684 (N_1684,In_1884,In_4598);
nor U1685 (N_1685,In_4752,In_4666);
and U1686 (N_1686,In_4303,In_2478);
and U1687 (N_1687,In_4753,In_2295);
nor U1688 (N_1688,In_2886,In_153);
and U1689 (N_1689,In_4935,In_4910);
xnor U1690 (N_1690,In_2275,In_346);
xnor U1691 (N_1691,In_2290,In_2969);
nor U1692 (N_1692,In_1001,In_2919);
nor U1693 (N_1693,In_1478,In_3378);
nor U1694 (N_1694,In_1801,In_812);
xnor U1695 (N_1695,In_904,In_1818);
or U1696 (N_1696,In_4216,In_3005);
xor U1697 (N_1697,In_4646,In_3137);
nor U1698 (N_1698,In_2532,In_1919);
and U1699 (N_1699,In_4512,In_740);
and U1700 (N_1700,In_4345,In_4534);
xnor U1701 (N_1701,In_3734,In_3044);
and U1702 (N_1702,In_545,In_4579);
or U1703 (N_1703,In_3489,In_3834);
nand U1704 (N_1704,In_4376,In_2812);
nor U1705 (N_1705,In_4438,In_4901);
and U1706 (N_1706,In_967,In_4420);
nand U1707 (N_1707,In_998,In_4417);
nor U1708 (N_1708,In_2319,In_3087);
nand U1709 (N_1709,In_3322,In_2410);
nand U1710 (N_1710,In_861,In_2228);
or U1711 (N_1711,In_1674,In_4932);
or U1712 (N_1712,In_1495,In_1733);
or U1713 (N_1713,In_1384,In_4310);
nor U1714 (N_1714,In_3706,In_487);
or U1715 (N_1715,In_2534,In_3781);
xnor U1716 (N_1716,In_362,In_4520);
nand U1717 (N_1717,In_2206,In_1602);
xor U1718 (N_1718,In_3343,In_4533);
or U1719 (N_1719,In_2300,In_3602);
xnor U1720 (N_1720,In_1502,In_3256);
or U1721 (N_1721,In_1677,In_266);
and U1722 (N_1722,In_468,In_1879);
nor U1723 (N_1723,In_4069,In_2124);
and U1724 (N_1724,In_1279,In_3684);
nand U1725 (N_1725,In_2819,In_422);
or U1726 (N_1726,In_3599,In_3710);
and U1727 (N_1727,In_4266,In_1446);
or U1728 (N_1728,In_4174,In_4955);
or U1729 (N_1729,In_3494,In_1892);
xnor U1730 (N_1730,In_2544,In_1873);
xor U1731 (N_1731,In_1277,In_2709);
and U1732 (N_1732,In_3835,In_3872);
nand U1733 (N_1733,In_3243,In_2731);
nand U1734 (N_1734,In_3954,In_1160);
xnor U1735 (N_1735,In_3045,In_2166);
or U1736 (N_1736,In_1922,In_1624);
or U1737 (N_1737,In_4899,In_4791);
or U1738 (N_1738,In_616,In_4693);
or U1739 (N_1739,In_1310,In_3892);
and U1740 (N_1740,In_3730,In_1573);
and U1741 (N_1741,In_878,In_2471);
and U1742 (N_1742,In_486,In_1340);
nand U1743 (N_1743,In_4134,In_1527);
or U1744 (N_1744,In_1327,In_3615);
or U1745 (N_1745,In_3385,In_2927);
and U1746 (N_1746,In_200,In_1972);
nand U1747 (N_1747,In_2345,In_1043);
nor U1748 (N_1748,In_2424,In_4497);
nand U1749 (N_1749,In_4996,In_2611);
or U1750 (N_1750,In_580,In_1126);
nor U1751 (N_1751,In_2546,In_2431);
and U1752 (N_1752,In_2288,In_4730);
nor U1753 (N_1753,In_1096,In_2735);
or U1754 (N_1754,In_4039,In_3129);
or U1755 (N_1755,In_3786,In_1789);
or U1756 (N_1756,In_1462,In_3476);
xor U1757 (N_1757,In_2632,In_914);
xor U1758 (N_1758,In_4884,In_611);
and U1759 (N_1759,In_3690,In_3534);
xnor U1760 (N_1760,In_1987,In_3200);
nand U1761 (N_1761,In_1458,In_2603);
and U1762 (N_1762,In_2753,In_3191);
nand U1763 (N_1763,In_2740,In_2955);
nand U1764 (N_1764,In_363,In_4781);
and U1765 (N_1765,In_4049,In_276);
xnor U1766 (N_1766,In_3155,In_4429);
or U1767 (N_1767,In_4945,In_984);
nor U1768 (N_1768,In_905,In_2835);
xnor U1769 (N_1769,In_70,In_233);
or U1770 (N_1770,In_4098,In_224);
nand U1771 (N_1771,In_2811,In_1457);
and U1772 (N_1772,In_137,In_4295);
or U1773 (N_1773,In_1032,In_1497);
or U1774 (N_1774,In_1615,In_2944);
nor U1775 (N_1775,In_2989,In_1068);
nand U1776 (N_1776,In_4815,In_1755);
nand U1777 (N_1777,In_1200,In_1603);
and U1778 (N_1778,In_4499,In_4647);
nand U1779 (N_1779,In_1946,In_4434);
xor U1780 (N_1780,In_3778,In_4150);
nor U1781 (N_1781,In_4832,In_3454);
or U1782 (N_1782,In_4587,In_4135);
nand U1783 (N_1783,In_2222,In_575);
and U1784 (N_1784,In_1314,In_737);
or U1785 (N_1785,In_4965,In_623);
nand U1786 (N_1786,In_2697,In_2522);
or U1787 (N_1787,In_1152,In_3323);
and U1788 (N_1788,In_3130,In_1769);
or U1789 (N_1789,In_1697,In_4936);
and U1790 (N_1790,In_4298,In_183);
xor U1791 (N_1791,In_3585,In_4156);
nand U1792 (N_1792,In_3563,In_1453);
or U1793 (N_1793,In_2116,In_316);
nor U1794 (N_1794,In_1735,In_1338);
xnor U1795 (N_1795,In_953,In_4074);
or U1796 (N_1796,In_3802,In_304);
nor U1797 (N_1797,In_1362,In_226);
and U1798 (N_1798,In_765,In_4369);
nand U1799 (N_1799,In_2795,In_1718);
nand U1800 (N_1800,In_3431,In_1122);
or U1801 (N_1801,In_4255,In_4471);
nor U1802 (N_1802,In_4095,In_1518);
and U1803 (N_1803,In_2079,In_160);
nor U1804 (N_1804,In_3854,In_3376);
nand U1805 (N_1805,In_1166,In_4288);
nand U1806 (N_1806,In_565,In_361);
or U1807 (N_1807,In_1489,In_1107);
or U1808 (N_1808,In_1749,In_1817);
nor U1809 (N_1809,In_2223,In_2379);
nor U1810 (N_1810,In_4992,In_620);
xnor U1811 (N_1811,In_4835,In_2851);
xor U1812 (N_1812,In_3349,In_4470);
nand U1813 (N_1813,In_1185,In_3051);
nand U1814 (N_1814,In_1403,In_3499);
nand U1815 (N_1815,In_1193,In_4225);
xor U1816 (N_1816,In_3856,In_4614);
and U1817 (N_1817,In_4876,In_1547);
or U1818 (N_1818,In_1463,In_572);
nand U1819 (N_1819,In_3738,In_1195);
or U1820 (N_1820,In_4065,In_3062);
nand U1821 (N_1821,In_4243,In_1182);
nand U1822 (N_1822,In_4751,In_1366);
nor U1823 (N_1823,In_2126,In_2542);
or U1824 (N_1824,In_3606,In_2836);
and U1825 (N_1825,In_4677,In_2213);
or U1826 (N_1826,In_1392,In_1488);
or U1827 (N_1827,In_773,In_3860);
or U1828 (N_1828,In_103,In_4191);
xor U1829 (N_1829,In_2023,In_513);
and U1830 (N_1830,In_1800,In_2397);
xor U1831 (N_1831,In_1077,In_79);
nor U1832 (N_1832,In_4163,In_4505);
and U1833 (N_1833,In_157,In_431);
and U1834 (N_1834,In_2690,In_1360);
xor U1835 (N_1835,In_726,In_1751);
xor U1836 (N_1836,In_1807,In_459);
nor U1837 (N_1837,In_3746,In_4676);
nor U1838 (N_1838,In_4305,In_51);
nor U1839 (N_1839,In_2509,In_2418);
nor U1840 (N_1840,In_1278,In_1207);
nor U1841 (N_1841,In_2060,In_4853);
nand U1842 (N_1842,In_1334,In_3079);
nand U1843 (N_1843,In_4987,In_673);
and U1844 (N_1844,In_2038,In_28);
or U1845 (N_1845,In_2526,In_4705);
xnor U1846 (N_1846,In_2734,In_1726);
nor U1847 (N_1847,In_3204,In_3488);
or U1848 (N_1848,In_3811,In_197);
xor U1849 (N_1849,In_2705,In_2830);
xnor U1850 (N_1850,In_1097,In_4496);
or U1851 (N_1851,In_1147,In_4621);
and U1852 (N_1852,In_2143,In_3956);
nor U1853 (N_1853,In_3559,In_273);
xnor U1854 (N_1854,In_3168,In_4769);
or U1855 (N_1855,In_846,In_1564);
nand U1856 (N_1856,In_1675,In_24);
nand U1857 (N_1857,In_423,In_3950);
nand U1858 (N_1858,In_3660,In_1477);
nor U1859 (N_1859,In_204,In_1350);
and U1860 (N_1860,In_3827,In_3517);
xnor U1861 (N_1861,In_4920,In_219);
and U1862 (N_1862,In_2782,In_1418);
and U1863 (N_1863,In_1520,In_1845);
nor U1864 (N_1864,In_670,In_4466);
and U1865 (N_1865,In_4332,In_1258);
and U1866 (N_1866,In_2312,In_2046);
nor U1867 (N_1867,In_3533,In_3975);
and U1868 (N_1868,In_2248,In_4766);
xor U1869 (N_1869,In_2967,In_4943);
nor U1870 (N_1870,In_1217,In_1303);
or U1871 (N_1871,In_3380,In_826);
nor U1872 (N_1872,In_3066,In_777);
and U1873 (N_1873,In_1582,In_3859);
nand U1874 (N_1874,In_332,In_2434);
or U1875 (N_1875,In_1846,In_810);
or U1876 (N_1876,In_1510,In_3521);
or U1877 (N_1877,In_1421,In_291);
nand U1878 (N_1878,In_909,In_2996);
or U1879 (N_1879,In_4895,In_1517);
or U1880 (N_1880,In_1894,In_2405);
nand U1881 (N_1881,In_3630,In_3889);
or U1882 (N_1882,In_1294,In_2713);
and U1883 (N_1883,In_1654,In_3689);
xor U1884 (N_1884,In_697,In_3848);
nor U1885 (N_1885,In_3415,In_2445);
nand U1886 (N_1886,In_1897,In_3625);
xnor U1887 (N_1887,In_254,In_4510);
xor U1888 (N_1888,In_483,In_4974);
or U1889 (N_1889,In_2076,In_883);
and U1890 (N_1890,In_3795,In_3319);
and U1891 (N_1891,In_4103,In_3642);
or U1892 (N_1892,In_2612,In_3917);
nand U1893 (N_1893,In_465,In_2790);
xor U1894 (N_1894,In_4746,In_4707);
and U1895 (N_1895,In_4981,In_4050);
nand U1896 (N_1896,In_1765,In_988);
and U1897 (N_1897,In_4262,In_1424);
or U1898 (N_1898,In_1891,In_4453);
nor U1899 (N_1899,In_3930,In_3195);
and U1900 (N_1900,In_1627,In_3762);
nor U1901 (N_1901,In_384,In_4201);
and U1902 (N_1902,In_3363,In_2913);
nand U1903 (N_1903,In_4765,In_2050);
xor U1904 (N_1904,In_1658,In_3558);
xor U1905 (N_1905,In_4235,In_1042);
and U1906 (N_1906,In_531,In_4627);
nor U1907 (N_1907,In_3501,In_1119);
nor U1908 (N_1908,In_3641,In_48);
xor U1909 (N_1909,In_2711,In_491);
nor U1910 (N_1910,In_516,In_2344);
or U1911 (N_1911,In_94,In_2784);
xnor U1912 (N_1912,In_1775,In_4625);
nand U1913 (N_1913,In_3138,In_1342);
xor U1914 (N_1914,In_1168,In_664);
or U1915 (N_1915,In_1208,In_3018);
nand U1916 (N_1916,In_4728,In_4275);
xor U1917 (N_1917,In_807,In_4564);
and U1918 (N_1918,In_4513,In_19);
xor U1919 (N_1919,In_1657,In_26);
nor U1920 (N_1920,In_4389,In_3395);
and U1921 (N_1921,In_2197,In_3527);
nor U1922 (N_1922,In_4761,In_3541);
or U1923 (N_1923,In_2216,In_4005);
nor U1924 (N_1924,In_4673,In_2600);
nor U1925 (N_1925,In_3604,In_299);
xnor U1926 (N_1926,In_4334,In_2789);
nor U1927 (N_1927,In_903,In_4181);
xor U1928 (N_1928,In_1169,In_3027);
xor U1929 (N_1929,In_1040,In_2380);
and U1930 (N_1930,In_3671,In_4003);
nor U1931 (N_1931,In_1079,In_4154);
xnor U1932 (N_1932,In_2529,In_2861);
or U1933 (N_1933,In_2056,In_2210);
nor U1934 (N_1934,In_764,In_2423);
xor U1935 (N_1935,In_797,In_4053);
and U1936 (N_1936,In_753,In_1831);
nand U1937 (N_1937,In_2642,In_494);
or U1938 (N_1938,In_2660,In_1173);
nor U1939 (N_1939,In_2476,In_367);
and U1940 (N_1940,In_3170,In_4702);
nand U1941 (N_1941,In_4717,In_4207);
or U1942 (N_1942,In_497,In_259);
xnor U1943 (N_1943,In_4993,In_1746);
nor U1944 (N_1944,In_747,In_4062);
and U1945 (N_1945,In_717,In_2443);
nor U1946 (N_1946,In_2325,In_4538);
and U1947 (N_1947,In_2681,In_1326);
xor U1948 (N_1948,In_615,In_3257);
xnor U1949 (N_1949,In_1236,In_348);
or U1950 (N_1950,In_1090,In_3268);
and U1951 (N_1951,In_1455,In_2847);
xnor U1952 (N_1952,In_3414,In_3188);
nand U1953 (N_1953,In_3089,In_733);
and U1954 (N_1954,In_3391,In_4551);
nor U1955 (N_1955,In_131,In_775);
nand U1956 (N_1956,In_1019,In_3904);
nand U1957 (N_1957,In_1137,In_89);
and U1958 (N_1958,In_72,In_2351);
nor U1959 (N_1959,In_538,In_780);
nor U1960 (N_1960,In_1722,In_3847);
nand U1961 (N_1961,In_3324,In_4562);
and U1962 (N_1962,In_376,In_4064);
xor U1963 (N_1963,In_4264,In_2364);
nand U1964 (N_1964,In_3379,In_3306);
nand U1965 (N_1965,In_1012,In_2378);
nand U1966 (N_1966,In_3381,In_437);
nor U1967 (N_1967,In_1428,In_2508);
or U1968 (N_1968,In_1427,In_2786);
nor U1969 (N_1969,In_2842,In_3863);
nand U1970 (N_1970,In_3976,In_2306);
or U1971 (N_1971,In_1990,In_1524);
or U1972 (N_1972,In_4662,In_3279);
or U1973 (N_1973,In_3669,In_3718);
nor U1974 (N_1974,In_2195,In_1704);
nand U1975 (N_1975,In_2970,In_815);
nor U1976 (N_1976,In_3479,In_1078);
xor U1977 (N_1977,In_4,In_3245);
and U1978 (N_1978,In_932,In_557);
nand U1979 (N_1979,In_4686,In_1201);
nor U1980 (N_1980,In_3389,In_4294);
xor U1981 (N_1981,In_2203,In_164);
and U1982 (N_1982,In_3962,In_3124);
and U1983 (N_1983,In_4555,In_3816);
and U1984 (N_1984,In_2329,In_4674);
or U1985 (N_1985,In_3401,In_3215);
nor U1986 (N_1986,In_3357,In_2335);
xor U1987 (N_1987,In_3825,In_3075);
nand U1988 (N_1988,In_2513,In_2645);
nor U1989 (N_1989,In_4004,In_238);
or U1990 (N_1990,In_4969,In_3933);
and U1991 (N_1991,In_4590,In_1411);
xor U1992 (N_1992,In_2557,In_1349);
xnor U1993 (N_1993,In_1117,In_386);
xor U1994 (N_1994,In_3478,In_4390);
nand U1995 (N_1995,In_1021,In_542);
and U1996 (N_1996,In_2756,In_4405);
nand U1997 (N_1997,In_1046,In_539);
and U1998 (N_1998,In_2317,In_389);
or U1999 (N_1999,In_1863,In_1868);
nand U2000 (N_2000,N_1438,N_195);
nor U2001 (N_2001,N_1154,In_927);
nand U2002 (N_2002,In_4465,N_1681);
and U2003 (N_2003,N_966,In_2725);
and U2004 (N_2004,In_3595,N_1259);
and U2005 (N_2005,N_169,N_780);
or U2006 (N_2006,N_16,N_128);
nor U2007 (N_2007,N_216,In_3202);
and U2008 (N_2008,N_60,N_641);
or U2009 (N_2009,In_1634,In_3297);
nor U2010 (N_2010,N_1521,N_1662);
nand U2011 (N_2011,N_1588,N_1785);
xor U2012 (N_2012,In_2262,In_1734);
nand U2013 (N_2013,N_204,N_1227);
or U2014 (N_2014,N_1968,In_4724);
nor U2015 (N_2015,N_34,N_1889);
or U2016 (N_2016,N_1641,In_4282);
and U2017 (N_2017,In_2052,N_1740);
or U2018 (N_2018,In_4596,N_1043);
nand U2019 (N_2019,N_442,In_3413);
xnor U2020 (N_2020,N_1480,N_86);
xor U2021 (N_2021,N_1042,In_822);
and U2022 (N_2022,In_609,N_625);
xnor U2023 (N_2023,In_4377,In_2738);
nand U2024 (N_2024,N_1821,N_636);
nor U2025 (N_2025,N_663,N_245);
xor U2026 (N_2026,N_1879,N_720);
nor U2027 (N_2027,N_1387,In_4430);
nand U2028 (N_2028,N_462,N_423);
or U2029 (N_2029,N_1411,N_401);
or U2030 (N_2030,N_998,In_2371);
or U2031 (N_2031,N_1554,In_93);
or U2032 (N_2032,In_2670,N_1519);
and U2033 (N_2033,N_644,N_1903);
nand U2034 (N_2034,In_4548,N_1338);
and U2035 (N_2035,In_4923,N_38);
nand U2036 (N_2036,In_3780,N_916);
and U2037 (N_2037,N_1256,In_1281);
nand U2038 (N_2038,N_1196,N_1505);
nand U2039 (N_2039,In_145,N_1478);
and U2040 (N_2040,N_384,N_1192);
or U2041 (N_2041,N_209,N_1344);
nor U2042 (N_2042,In_3545,N_1242);
xor U2043 (N_2043,N_262,N_1914);
or U2044 (N_2044,N_1436,N_967);
xnor U2045 (N_2045,N_1346,N_393);
or U2046 (N_2046,N_297,N_123);
xor U2047 (N_2047,In_4140,N_781);
xnor U2048 (N_2048,N_515,N_1516);
and U2049 (N_2049,N_170,In_514);
and U2050 (N_2050,N_1947,In_2667);
nand U2051 (N_2051,In_4982,N_880);
nor U2052 (N_2052,N_1324,In_4365);
nand U2053 (N_2053,N_469,N_311);
nand U2054 (N_2054,In_4147,N_1823);
or U2055 (N_2055,N_1674,In_3345);
and U2056 (N_2056,N_968,In_819);
or U2057 (N_2057,In_2427,In_3553);
nor U2058 (N_2058,N_609,In_2385);
and U2059 (N_2059,In_3512,N_1584);
nor U2060 (N_2060,N_706,In_1272);
nor U2061 (N_2061,N_1663,N_1393);
xnor U2062 (N_2062,In_3713,N_1099);
and U2063 (N_2063,N_776,N_1226);
nand U2064 (N_2064,N_35,N_1090);
nand U2065 (N_2065,In_347,N_1445);
or U2066 (N_2066,N_660,N_573);
and U2067 (N_2067,In_3331,N_755);
xnor U2068 (N_2068,N_794,N_1919);
or U2069 (N_2069,N_714,N_273);
and U2070 (N_2070,N_1389,N_1190);
and U2071 (N_2071,N_414,N_783);
nor U2072 (N_2072,N_657,N_917);
or U2073 (N_2073,N_555,N_1743);
and U2074 (N_2074,N_1343,In_3979);
nor U2075 (N_2075,N_1850,N_1683);
and U2076 (N_2076,N_1132,N_649);
nand U2077 (N_2077,N_980,N_1044);
xor U2078 (N_2078,N_1945,N_1738);
or U2079 (N_2079,N_118,In_3994);
nor U2080 (N_2080,In_4281,N_1960);
nand U2081 (N_2081,N_786,N_1579);
or U2082 (N_2082,N_557,N_1397);
and U2083 (N_2083,In_452,N_418);
and U2084 (N_2084,N_1027,N_1517);
nor U2085 (N_2085,In_135,In_1720);
xor U2086 (N_2086,N_10,N_78);
or U2087 (N_2087,N_107,N_868);
or U2088 (N_2088,N_749,N_433);
nor U2089 (N_2089,In_2537,In_2507);
or U2090 (N_2090,In_4404,N_1668);
nor U2091 (N_2091,N_550,N_973);
nand U2092 (N_2092,N_1704,N_1727);
nand U2093 (N_2093,N_457,N_836);
and U2094 (N_2094,N_590,In_2663);
nor U2095 (N_2095,N_361,N_264);
or U2096 (N_2096,In_1730,N_1468);
and U2097 (N_2097,N_934,N_1509);
nand U2098 (N_2098,N_1184,In_2860);
or U2099 (N_2099,N_499,In_434);
nor U2100 (N_2100,N_1199,N_633);
or U2101 (N_2101,N_1978,N_626);
nand U2102 (N_2102,N_1975,In_1347);
xnor U2103 (N_2103,In_4356,In_1771);
and U2104 (N_2104,N_650,N_1959);
or U2105 (N_2105,N_788,N_1898);
and U2106 (N_2106,N_322,N_984);
xnor U2107 (N_2107,N_1014,N_1680);
xor U2108 (N_2108,N_106,In_2665);
xnor U2109 (N_2109,N_547,N_922);
nor U2110 (N_2110,In_1248,N_1580);
xnor U2111 (N_2111,N_1007,N_452);
nor U2112 (N_2112,In_3515,In_1952);
nor U2113 (N_2113,N_812,N_424);
and U2114 (N_2114,N_298,In_67);
nor U2115 (N_2115,In_3340,In_1843);
and U2116 (N_2116,N_1283,N_862);
nor U2117 (N_2117,N_1800,In_2696);
and U2118 (N_2118,In_2121,N_1529);
nand U2119 (N_2119,N_1363,N_632);
and U2120 (N_2120,N_772,N_347);
or U2121 (N_2121,In_1422,N_761);
nor U2122 (N_2122,N_511,N_620);
and U2123 (N_2123,In_1514,N_859);
nand U2124 (N_2124,In_167,N_743);
nor U2125 (N_2125,N_726,N_1498);
nor U2126 (N_2126,N_1459,In_4811);
nor U2127 (N_2127,N_655,In_1133);
xor U2128 (N_2128,N_1682,N_3);
and U2129 (N_2129,N_1130,N_274);
nor U2130 (N_2130,N_39,N_408);
xnor U2131 (N_2131,N_1065,In_4768);
xor U2132 (N_2132,N_882,In_586);
xnor U2133 (N_2133,N_528,In_4410);
xor U2134 (N_2134,In_3888,In_3929);
xor U2135 (N_2135,N_1334,N_68);
or U2136 (N_2136,N_380,In_476);
and U2137 (N_2137,N_841,N_1816);
nor U2138 (N_2138,N_1449,N_1345);
xnor U2139 (N_2139,N_168,N_416);
or U2140 (N_2140,N_855,N_1114);
and U2141 (N_2141,N_1031,N_472);
or U2142 (N_2142,N_1954,N_314);
or U2143 (N_2143,N_315,N_753);
and U2144 (N_2144,N_1170,N_1286);
xnor U2145 (N_2145,N_125,N_1070);
nand U2146 (N_2146,N_1780,In_350);
nor U2147 (N_2147,In_1595,N_1531);
nand U2148 (N_2148,N_1365,N_1967);
or U2149 (N_2149,N_1431,In_2069);
and U2150 (N_2150,N_825,N_1744);
and U2151 (N_2151,In_102,N_1572);
or U2152 (N_2152,N_614,N_7);
nand U2153 (N_2153,In_4425,N_1167);
or U2154 (N_2154,N_1722,N_618);
xor U2155 (N_2155,N_599,In_1631);
nand U2156 (N_2156,N_1008,In_4814);
xnor U2157 (N_2157,N_1137,N_1822);
xor U2158 (N_2158,In_1676,N_1185);
xnor U2159 (N_2159,N_71,N_1403);
nor U2160 (N_2160,N_845,In_743);
and U2161 (N_2161,N_1587,N_1485);
and U2162 (N_2162,N_854,N_1694);
or U2163 (N_2163,In_366,In_2968);
and U2164 (N_2164,N_782,In_278);
nand U2165 (N_2165,N_1054,In_225);
or U2166 (N_2166,N_1653,N_1558);
nand U2167 (N_2167,N_112,N_489);
nor U2168 (N_2168,In_4714,In_2236);
xor U2169 (N_2169,In_1728,In_1985);
nor U2170 (N_2170,In_4250,N_1470);
nor U2171 (N_2171,N_1661,N_1963);
or U2172 (N_2172,N_358,In_3198);
xor U2173 (N_2173,N_1425,N_1883);
nand U2174 (N_2174,N_356,N_970);
or U2175 (N_2175,In_1932,N_1550);
and U2176 (N_2176,N_448,In_4736);
and U2177 (N_2177,In_4898,In_639);
nor U2178 (N_2178,In_796,N_1247);
nor U2179 (N_2179,In_1026,In_1080);
nand U2180 (N_2180,In_2272,In_2040);
or U2181 (N_2181,In_4448,In_3203);
nor U2182 (N_2182,N_563,In_4747);
nor U2183 (N_2183,In_194,N_838);
nor U2184 (N_2184,N_1069,N_1559);
xor U2185 (N_2185,In_1038,In_439);
and U2186 (N_2186,N_1094,In_2662);
nor U2187 (N_2187,N_1248,In_4194);
and U2188 (N_2188,In_768,N_167);
nor U2189 (N_2189,N_198,N_300);
or U2190 (N_2190,N_1646,N_302);
and U2191 (N_2191,N_512,N_390);
nand U2192 (N_2192,N_936,N_785);
nand U2193 (N_2193,In_562,N_191);
and U2194 (N_2194,N_974,N_260);
or U2195 (N_2195,N_809,N_1512);
xnor U2196 (N_2196,In_1784,N_186);
or U2197 (N_2197,N_477,N_1049);
xor U2198 (N_2198,In_4426,N_1020);
or U2199 (N_2199,N_1706,N_535);
nor U2200 (N_2200,N_1165,N_1560);
nand U2201 (N_2201,N_1456,In_2701);
xor U2202 (N_2202,N_758,In_2888);
or U2203 (N_2203,In_196,N_1483);
nand U2204 (N_2204,N_1322,N_1932);
nor U2205 (N_2205,N_441,In_1);
nor U2206 (N_2206,In_2234,N_956);
or U2207 (N_2207,In_3886,N_1328);
xor U2208 (N_2208,N_796,N_1987);
or U2209 (N_2209,N_194,N_1144);
nand U2210 (N_2210,N_864,N_594);
nor U2211 (N_2211,N_1570,In_4324);
nand U2212 (N_2212,N_1477,N_722);
xnor U2213 (N_2213,In_3000,N_1039);
nor U2214 (N_2214,In_2516,N_1539);
nor U2215 (N_2215,In_921,In_4780);
nand U2216 (N_2216,In_3249,N_122);
and U2217 (N_2217,In_3928,N_1759);
nand U2218 (N_2218,N_1335,In_4966);
nand U2219 (N_2219,N_1213,N_830);
and U2220 (N_2220,N_1467,In_544);
nand U2221 (N_2221,In_1762,In_4774);
or U2222 (N_2222,N_645,N_728);
nor U2223 (N_2223,N_44,N_1711);
or U2224 (N_2224,In_971,In_25);
xnor U2225 (N_2225,N_124,N_1736);
or U2226 (N_2226,In_1619,N_370);
nor U2227 (N_2227,N_1360,N_1046);
or U2228 (N_2228,In_3887,In_2001);
nor U2229 (N_2229,N_1314,N_1677);
nand U2230 (N_2230,In_4893,N_248);
and U2231 (N_2231,In_3716,N_337);
and U2232 (N_2232,N_615,N_1349);
or U2233 (N_2233,N_1002,In_1394);
nand U2234 (N_2234,N_50,N_546);
or U2235 (N_2235,N_90,N_220);
nor U2236 (N_2236,N_192,In_3654);
nor U2237 (N_2237,In_3135,N_847);
or U2238 (N_2238,N_1299,N_74);
and U2239 (N_2239,In_50,N_1916);
and U2240 (N_2240,In_4198,In_706);
nor U2241 (N_2241,N_114,N_668);
nor U2242 (N_2242,In_1423,N_1532);
or U2243 (N_2243,In_2404,In_2504);
and U2244 (N_2244,In_3151,In_2598);
or U2245 (N_2245,N_565,In_1237);
and U2246 (N_2246,N_1616,N_1979);
xnor U2247 (N_2247,N_1832,N_1203);
and U2248 (N_2248,In_2510,In_2316);
xnor U2249 (N_2249,N_1219,N_1417);
xnor U2250 (N_2250,In_1629,N_1555);
or U2251 (N_2251,In_4028,N_923);
xor U2252 (N_2252,In_2908,In_1433);
nand U2253 (N_2253,In_2337,N_246);
or U2254 (N_2254,In_790,In_4658);
and U2255 (N_2255,In_729,N_558);
nand U2256 (N_2256,N_223,N_187);
or U2257 (N_2257,N_26,In_8);
and U2258 (N_2258,N_294,In_4655);
and U2259 (N_2259,In_2885,N_1262);
or U2260 (N_2260,N_31,N_556);
and U2261 (N_2261,In_1449,N_1038);
or U2262 (N_2262,N_1061,N_1557);
nor U2263 (N_2263,In_1521,N_411);
nand U2264 (N_2264,N_1941,In_2201);
or U2265 (N_2265,N_664,In_1826);
nor U2266 (N_2266,N_937,N_1788);
or U2267 (N_2267,In_3119,N_498);
or U2268 (N_2268,In_721,In_285);
xor U2269 (N_2269,N_1924,N_1095);
nand U2270 (N_2270,N_1761,N_1866);
or U2271 (N_2271,N_1909,N_1120);
nand U2272 (N_2272,In_3900,N_1669);
or U2273 (N_2273,In_2655,N_1188);
xnor U2274 (N_2274,N_1848,N_1986);
nand U2275 (N_2275,In_1575,N_1993);
and U2276 (N_2276,N_1264,N_87);
and U2277 (N_2277,N_637,N_1421);
or U2278 (N_2278,N_1133,In_1815);
nand U2279 (N_2279,In_1804,N_737);
or U2280 (N_2280,N_593,In_2616);
xor U2281 (N_2281,In_281,N_848);
nand U2282 (N_2282,In_818,N_234);
or U2283 (N_2283,N_1958,N_58);
xnor U2284 (N_2284,N_666,N_1396);
nand U2285 (N_2285,N_1464,N_189);
or U2286 (N_2286,N_268,In_3080);
or U2287 (N_2287,N_1621,N_410);
xnor U2288 (N_2288,N_53,N_1655);
nor U2289 (N_2289,In_4353,N_1942);
or U2290 (N_2290,N_1892,In_3206);
xnor U2291 (N_2291,N_1996,N_1873);
nor U2292 (N_2292,In_4025,N_478);
or U2293 (N_2293,In_4245,N_1172);
xnor U2294 (N_2294,N_1342,In_506);
nor U2295 (N_2295,In_4578,N_461);
nand U2296 (N_2296,N_612,N_345);
xor U2297 (N_2297,N_63,N_1847);
nand U2298 (N_2298,N_221,N_1923);
nand U2299 (N_2299,N_1238,N_1724);
or U2300 (N_2300,In_4783,In_1219);
and U2301 (N_2301,N_1482,N_1920);
or U2302 (N_2302,In_608,N_1614);
or U2303 (N_2303,N_250,N_152);
or U2304 (N_2304,N_1814,In_2728);
or U2305 (N_2305,N_1552,N_676);
nand U2306 (N_2306,N_444,N_519);
or U2307 (N_2307,N_629,N_62);
and U2308 (N_2308,In_2486,N_694);
xor U2309 (N_2309,N_1072,N_1371);
xnor U2310 (N_2310,N_490,N_467);
and U2311 (N_2311,In_4254,N_1409);
nor U2312 (N_2312,N_1922,In_3529);
nor U2313 (N_2313,In_3114,N_1518);
nor U2314 (N_2314,In_1607,N_1025);
nand U2315 (N_2315,N_257,N_57);
nand U2316 (N_2316,In_1925,N_82);
nand U2317 (N_2317,In_1632,N_1511);
or U2318 (N_2318,N_1490,N_500);
nand U2319 (N_2319,N_811,N_231);
xnor U2320 (N_2320,N_1157,N_131);
or U2321 (N_2321,N_927,N_1354);
nand U2322 (N_2322,N_238,In_4458);
nor U2323 (N_2323,In_2183,N_1991);
nand U2324 (N_2324,In_317,In_923);
nand U2325 (N_2325,In_1885,N_1151);
nand U2326 (N_2326,N_1605,In_1904);
or U2327 (N_2327,N_1632,N_1194);
xnor U2328 (N_2328,N_104,N_285);
and U2329 (N_2329,In_3132,N_1657);
nand U2330 (N_2330,N_746,N_1625);
nand U2331 (N_2331,N_562,In_1608);
nor U2332 (N_2332,N_536,N_619);
nand U2333 (N_2333,N_903,In_2700);
and U2334 (N_2334,N_1854,In_4077);
xnor U2335 (N_2335,In_2302,N_1323);
nand U2336 (N_2336,In_2468,N_656);
xor U2337 (N_2337,In_3883,N_1285);
or U2338 (N_2338,N_134,N_1163);
and U2339 (N_2339,In_3611,In_490);
and U2340 (N_2340,In_3468,In_2144);
and U2341 (N_2341,In_29,In_2727);
and U2342 (N_2342,N_372,N_1811);
and U2343 (N_2343,In_4900,N_1590);
nand U2344 (N_2344,N_1430,N_413);
and U2345 (N_2345,In_957,In_3750);
or U2346 (N_2346,N_819,N_564);
and U2347 (N_2347,N_779,In_4622);
and U2348 (N_2348,N_730,N_270);
nand U2349 (N_2349,N_1983,In_3099);
nand U2350 (N_2350,N_559,N_527);
xor U2351 (N_2351,N_1925,N_1428);
or U2352 (N_2352,N_249,In_315);
and U2353 (N_2353,N_1755,N_858);
or U2354 (N_2354,N_576,N_1802);
nand U2355 (N_2355,In_1882,N_105);
nand U2356 (N_2356,N_335,N_210);
and U2357 (N_2357,N_1766,N_1944);
or U2358 (N_2358,In_3444,N_1749);
and U2359 (N_2359,N_1725,N_486);
nor U2360 (N_2360,In_1963,N_1041);
and U2361 (N_2361,In_1923,In_4802);
and U2362 (N_2362,In_3211,N_41);
nor U2363 (N_2363,N_47,N_1765);
nand U2364 (N_2364,In_3866,In_415);
xor U2365 (N_2365,In_3133,N_164);
and U2366 (N_2366,N_1352,N_1169);
nand U2367 (N_2367,N_340,In_2475);
nand U2368 (N_2368,N_1401,N_1272);
nor U2369 (N_2369,N_1469,In_2462);
nand U2370 (N_2370,N_1508,N_1280);
xnor U2371 (N_2371,N_929,N_437);
nand U2372 (N_2372,N_1015,N_1865);
nor U2373 (N_2373,N_188,In_1821);
nand U2374 (N_2374,N_957,In_1911);
or U2375 (N_2375,In_2147,N_1731);
or U2376 (N_2376,In_3620,In_3605);
and U2377 (N_2377,N_803,N_200);
and U2378 (N_2378,In_1917,In_1792);
and U2379 (N_2379,In_3590,N_1257);
nor U2380 (N_2380,N_1191,N_543);
and U2381 (N_2381,N_742,N_1260);
or U2382 (N_2382,In_63,In_1850);
nand U2383 (N_2383,N_821,N_1040);
nor U2384 (N_2384,In_1235,In_3652);
or U2385 (N_2385,N_148,In_4323);
nor U2386 (N_2386,N_560,N_93);
nand U2387 (N_2387,N_307,N_1100);
or U2388 (N_2388,N_1209,N_1206);
nand U2389 (N_2389,N_1992,N_975);
or U2390 (N_2390,N_1358,In_3921);
nand U2391 (N_2391,In_919,In_3213);
and U2392 (N_2392,N_1471,In_1605);
xnor U2393 (N_2393,N_492,N_1447);
and U2394 (N_2394,In_3329,In_4620);
xnor U2395 (N_2395,N_718,N_592);
nand U2396 (N_2396,In_4445,N_491);
nor U2397 (N_2397,N_1825,In_282);
and U2398 (N_2398,N_1770,In_1665);
and U2399 (N_2399,N_607,N_362);
or U2400 (N_2400,In_3564,N_1796);
nand U2401 (N_2401,N_25,N_1465);
nand U2402 (N_2402,N_1950,In_3875);
or U2403 (N_2403,In_175,In_4418);
xor U2404 (N_2404,In_1618,N_378);
nand U2405 (N_2405,N_1977,In_899);
or U2406 (N_2406,N_482,N_1543);
or U2407 (N_2407,N_986,In_1515);
and U2408 (N_2408,N_520,In_776);
nand U2409 (N_2409,N_301,N_1782);
xor U2410 (N_2410,In_2747,N_1990);
nor U2411 (N_2411,N_1776,N_1636);
and U2412 (N_2412,N_1079,N_1212);
and U2413 (N_2413,N_892,N_915);
xor U2414 (N_2414,In_2334,N_1597);
or U2415 (N_2415,In_481,In_3148);
nor U2416 (N_2416,N_1406,In_2170);
xnor U2417 (N_2417,In_4239,N_1147);
and U2418 (N_2418,N_1384,In_1975);
or U2419 (N_2419,N_1448,N_799);
xor U2420 (N_2420,In_2097,N_601);
xnor U2421 (N_2421,N_1548,N_1880);
nor U2422 (N_2422,In_2465,In_3289);
and U2423 (N_2423,In_3570,In_2781);
xor U2424 (N_2424,In_2596,N_88);
nor U2425 (N_2425,N_276,N_977);
xnor U2426 (N_2426,N_1348,N_43);
or U2427 (N_2427,N_385,In_3436);
xnor U2428 (N_2428,N_1101,N_622);
nor U2429 (N_2429,In_951,N_1676);
xor U2430 (N_2430,N_417,N_496);
xor U2431 (N_2431,N_1528,N_1452);
nand U2432 (N_2432,N_386,N_1660);
nor U2433 (N_2433,N_1626,N_1538);
xnor U2434 (N_2434,N_674,N_1629);
nand U2435 (N_2435,In_1701,In_104);
xnor U2436 (N_2436,N_1836,N_1949);
and U2437 (N_2437,N_348,N_1862);
nor U2438 (N_2438,In_3108,N_483);
xor U2439 (N_2439,N_1455,N_373);
or U2440 (N_2440,N_793,N_531);
nor U2441 (N_2441,In_2853,N_1582);
xor U2442 (N_2442,N_1215,N_1412);
or U2443 (N_2443,In_3335,N_75);
nor U2444 (N_2444,N_1118,In_2257);
nand U2445 (N_2445,In_4809,In_1091);
nand U2446 (N_2446,In_371,N_797);
or U2447 (N_2447,In_3235,N_996);
nor U2448 (N_2448,N_1441,N_237);
nor U2449 (N_2449,N_1961,N_309);
and U2450 (N_2450,N_1730,N_1999);
xor U2451 (N_2451,N_911,N_1381);
xnor U2452 (N_2452,N_1181,N_1066);
nor U2453 (N_2453,N_1871,N_1064);
xor U2454 (N_2454,N_1062,N_1073);
xor U2455 (N_2455,In_3293,In_1541);
and U2456 (N_2456,N_387,In_2373);
nor U2457 (N_2457,N_1152,N_954);
and U2458 (N_2458,N_960,N_283);
or U2459 (N_2459,N_1210,In_3302);
xor U2460 (N_2460,N_699,N_696);
nand U2461 (N_2461,In_4344,N_471);
and U2462 (N_2462,N_99,In_603);
or U2463 (N_2463,In_3791,In_3998);
or U2464 (N_2464,N_1443,N_365);
nand U2465 (N_2465,In_4173,N_241);
xor U2466 (N_2466,In_96,N_1726);
nor U2467 (N_2467,N_375,N_1504);
nor U2468 (N_2468,N_479,N_141);
or U2469 (N_2469,In_179,In_688);
or U2470 (N_2470,N_1826,In_3269);
nand U2471 (N_2471,In_4748,N_1427);
nor U2472 (N_2472,N_1778,N_379);
or U2473 (N_2473,In_159,N_205);
and U2474 (N_2474,In_1306,In_4998);
and U2475 (N_2475,N_814,N_1718);
nand U2476 (N_2476,N_135,In_4196);
or U2477 (N_2477,N_587,N_561);
and U2478 (N_2478,N_1177,N_303);
xnor U2479 (N_2479,N_1599,In_2061);
nor U2480 (N_2480,N_1001,In_1238);
xnor U2481 (N_2481,N_1325,N_1320);
nor U2482 (N_2482,N_939,N_1769);
and U2483 (N_2483,N_940,N_28);
nand U2484 (N_2484,In_2472,In_171);
and U2485 (N_2485,N_1868,N_218);
nor U2486 (N_2486,In_1256,In_1293);
xor U2487 (N_2487,N_1028,In_4380);
and U2488 (N_2488,N_49,N_1618);
xnor U2489 (N_2489,N_1249,In_4183);
and U2490 (N_2490,N_1442,N_1884);
nand U2491 (N_2491,N_475,N_277);
and U2492 (N_2492,N_1575,In_4193);
xnor U2493 (N_2493,In_1178,In_2081);
nor U2494 (N_2494,In_1225,In_3885);
nand U2495 (N_2495,In_3751,In_1553);
xnor U2496 (N_2496,N_1288,N_1757);
or U2497 (N_2497,N_1774,N_1450);
or U2498 (N_2498,N_1908,N_792);
nor U2499 (N_2499,In_961,N_388);
xor U2500 (N_2500,N_363,In_1071);
xor U2501 (N_2501,N_1232,N_1829);
xnor U2502 (N_2502,N_190,In_3139);
nor U2503 (N_2503,N_84,N_508);
xnor U2504 (N_2504,In_1139,In_1802);
nand U2505 (N_2505,In_4384,In_4401);
nand U2506 (N_2506,N_1234,N_391);
or U2507 (N_2507,N_484,In_3568);
or U2508 (N_2508,In_4309,In_3908);
nand U2509 (N_2509,N_1756,N_27);
and U2510 (N_2510,N_1269,N_224);
or U2511 (N_2511,N_8,N_1250);
nor U2512 (N_2512,In_1689,In_1419);
or U2513 (N_2513,In_3895,In_4063);
nor U2514 (N_2514,N_1615,N_523);
or U2515 (N_2515,N_458,N_1594);
nor U2516 (N_2516,In_4495,In_100);
nor U2517 (N_2517,N_881,In_4582);
and U2518 (N_2518,N_1472,N_944);
or U2519 (N_2519,In_2759,In_741);
nand U2520 (N_2520,In_3462,N_1651);
xnor U2521 (N_2521,N_506,N_602);
xnor U2522 (N_2522,N_45,N_113);
nor U2523 (N_2523,N_750,N_305);
or U2524 (N_2524,N_654,In_647);
or U2525 (N_2525,N_1965,N_1675);
or U2526 (N_2526,N_1098,N_1878);
nand U2527 (N_2527,N_725,In_4382);
and U2528 (N_2528,N_1601,N_1155);
and U2529 (N_2529,N_1620,N_1783);
nand U2530 (N_2530,N_137,N_978);
or U2531 (N_2531,N_589,N_1520);
or U2532 (N_2532,N_905,N_1691);
nand U2533 (N_2533,N_399,In_425);
nand U2534 (N_2534,N_162,In_2155);
nand U2535 (N_2535,N_1117,In_641);
nor U2536 (N_2536,N_752,In_438);
xnor U2537 (N_2537,N_995,N_1075);
nor U2538 (N_2538,In_2567,In_2945);
and U2539 (N_2539,N_325,N_1786);
nand U2540 (N_2540,In_2576,In_4602);
nand U2541 (N_2541,In_3077,N_700);
and U2542 (N_2542,In_2815,In_1695);
nor U2543 (N_2543,N_454,N_1377);
and U2544 (N_2544,N_1807,N_1638);
or U2545 (N_2545,N_406,N_178);
or U2546 (N_2546,N_517,N_1109);
xnor U2547 (N_2547,In_4388,N_733);
nor U2548 (N_2548,In_2479,N_976);
nand U2549 (N_2549,N_585,N_497);
or U2550 (N_2550,In_4663,N_1289);
and U2551 (N_2551,In_2282,N_904);
and U2552 (N_2552,In_1740,In_3169);
nand U2553 (N_2553,N_136,N_748);
nand U2554 (N_2554,N_1969,N_1093);
and U2555 (N_2555,N_914,N_1617);
nand U2556 (N_2556,In_2818,N_459);
nand U2557 (N_2557,N_768,N_815);
xnor U2558 (N_2558,In_106,N_1495);
xnor U2559 (N_2559,N_658,N_955);
or U2560 (N_2560,In_4085,N_357);
nand U2561 (N_2561,N_684,N_144);
nand U2562 (N_2562,N_1733,N_100);
nor U2563 (N_2563,N_1398,N_1678);
nand U2564 (N_2564,N_208,In_4754);
nor U2565 (N_2565,In_895,N_287);
or U2566 (N_2566,In_653,N_724);
or U2567 (N_2567,N_1798,N_999);
nand U2568 (N_2568,In_3842,N_893);
nand U2569 (N_2569,In_963,N_1561);
and U2570 (N_2570,N_1514,N_177);
xor U2571 (N_2571,N_1591,N_1327);
or U2572 (N_2572,In_3632,In_1047);
nand U2573 (N_2573,N_501,In_4257);
or U2574 (N_2574,In_1655,N_852);
and U2575 (N_2575,N_1578,N_1240);
or U2576 (N_2576,N_947,N_1896);
xor U2577 (N_2577,In_2906,N_202);
nand U2578 (N_2578,In_4326,N_953);
or U2579 (N_2579,N_875,In_907);
or U2580 (N_2580,N_149,N_360);
nand U2581 (N_2581,In_249,N_1563);
nand U2582 (N_2582,N_296,N_1321);
nand U2583 (N_2583,N_1915,N_1197);
nand U2584 (N_2584,N_179,N_505);
or U2585 (N_2585,In_3698,N_659);
nor U2586 (N_2586,N_407,N_1523);
and U2587 (N_2587,N_1502,N_1124);
nand U2588 (N_2588,N_1021,N_704);
nand U2589 (N_2589,N_886,N_1895);
and U2590 (N_2590,N_646,In_1473);
nand U2591 (N_2591,N_235,In_4500);
and U2592 (N_2592,N_1239,In_1945);
xor U2593 (N_2593,N_524,N_1931);
nand U2594 (N_2594,In_3951,N_708);
xor U2595 (N_2595,N_670,N_116);
and U2596 (N_2596,In_3296,In_4542);
and U2597 (N_2597,N_1491,N_1493);
or U2598 (N_2598,In_3384,N_1720);
xor U2599 (N_2599,In_2360,In_3057);
nor U2600 (N_2600,In_2157,N_1650);
and U2601 (N_2601,In_2250,N_692);
nand U2602 (N_2602,In_4120,In_1965);
xor U2603 (N_2603,N_4,N_431);
nor U2604 (N_2604,N_180,In_3679);
nand U2605 (N_2605,In_2187,N_1567);
nand U2606 (N_2606,N_138,N_1679);
xnor U2607 (N_2607,In_3896,In_2676);
xnor U2608 (N_2608,N_185,In_4569);
nand U2609 (N_2609,N_1420,N_1082);
nor U2610 (N_2610,N_930,N_1844);
xnor U2611 (N_2611,In_718,In_2141);
xor U2612 (N_2612,In_3052,In_667);
or U2613 (N_2613,N_877,N_1367);
and U2614 (N_2614,N_1458,N_1408);
nor U2615 (N_2615,In_1447,In_2080);
and U2616 (N_2616,N_604,N_290);
or U2617 (N_2617,N_703,N_1178);
xnor U2618 (N_2618,In_4784,In_2849);
nor U2619 (N_2619,N_738,In_808);
or U2620 (N_2620,N_1566,In_699);
or U2621 (N_2621,N_1767,N_804);
xnor U2622 (N_2622,In_4903,In_1203);
nor U2623 (N_2623,N_1688,N_1265);
nor U2624 (N_2624,In_4460,N_971);
nand U2625 (N_2625,N_935,N_18);
nor U2626 (N_2626,N_834,N_1026);
and U2627 (N_2627,N_1263,In_4742);
nor U2628 (N_2628,In_4033,In_3441);
nand U2629 (N_2629,N_317,In_31);
and U2630 (N_2630,N_333,In_4217);
or U2631 (N_2631,In_1436,N_1775);
xnor U2632 (N_2632,In_4732,N_534);
and U2633 (N_2633,In_4155,In_2783);
nor U2634 (N_2634,In_3644,N_1510);
nor U2635 (N_2635,N_1869,N_732);
nand U2636 (N_2636,In_4828,N_1708);
nand U2637 (N_2637,In_880,N_1574);
nand U2638 (N_2638,N_979,N_988);
and U2639 (N_2639,N_952,N_181);
nand U2640 (N_2640,N_701,N_846);
nand U2641 (N_2641,In_3996,N_1112);
xnor U2642 (N_2642,In_4890,N_610);
or U2643 (N_2643,In_2161,In_3981);
nand U2644 (N_2644,N_1623,N_1745);
or U2645 (N_2645,N_1905,N_765);
or U2646 (N_2646,In_882,N_443);
xor U2647 (N_2647,N_174,N_878);
or U2648 (N_2648,N_156,N_873);
and U2649 (N_2649,N_613,N_582);
xnor U2650 (N_2650,In_3029,In_392);
or U2651 (N_2651,In_937,N_1018);
and U2652 (N_2652,N_1697,N_635);
nand U2653 (N_2653,N_142,N_20);
or U2654 (N_2654,N_539,N_611);
and U2655 (N_2655,In_2926,N_199);
nor U2656 (N_2656,In_467,N_1053);
or U2657 (N_2657,In_3566,N_526);
xor U2658 (N_2658,N_744,In_2505);
nand U2659 (N_2659,N_709,N_1414);
or U2660 (N_2660,N_1673,N_747);
xor U2661 (N_2661,N_1233,In_2787);
and U2662 (N_2662,N_1180,In_4631);
xor U2663 (N_2663,N_1831,In_2548);
and U2664 (N_2664,N_1696,N_65);
nor U2665 (N_2665,N_1499,N_1245);
or U2666 (N_2666,N_117,N_400);
nor U2667 (N_2667,N_1361,N_1813);
nor U2668 (N_2668,N_267,N_1887);
nand U2669 (N_2669,In_90,N_263);
or U2670 (N_2670,In_3451,In_334);
nor U2671 (N_2671,N_310,In_4977);
nand U2672 (N_2672,N_51,N_1357);
or U2673 (N_2673,N_1762,In_2846);
nor U2674 (N_2674,N_1713,N_1690);
xnor U2675 (N_2675,N_292,In_3491);
nor U2676 (N_2676,N_145,N_1171);
and U2677 (N_2677,N_182,In_3691);
nor U2678 (N_2678,N_265,In_3582);
xnor U2679 (N_2679,N_1316,N_577);
nand U2680 (N_2680,N_521,In_778);
nand U2681 (N_2681,In_257,In_2120);
and U2682 (N_2682,N_1779,N_460);
xnor U2683 (N_2683,N_554,In_3526);
xor U2684 (N_2684,In_1188,In_625);
and U2685 (N_2685,N_1819,In_739);
nand U2686 (N_2686,In_3465,N_844);
and U2687 (N_2687,In_271,In_1787);
xor U2688 (N_2688,In_3317,N_569);
and U2689 (N_2689,N_247,N_1313);
nor U2690 (N_2690,N_1418,In_552);
nor U2691 (N_2691,N_72,In_911);
xor U2692 (N_2692,In_4279,N_1024);
nand U2693 (N_2693,N_1059,N_318);
or U2694 (N_2694,N_1687,In_727);
nand U2695 (N_2695,N_1108,N_1400);
xnor U2696 (N_2696,In_4350,In_4427);
xnor U2697 (N_2697,N_171,In_165);
and U2698 (N_2698,N_1773,N_1526);
nand U2699 (N_2699,N_353,N_827);
or U2700 (N_2700,N_306,N_965);
nand U2701 (N_2701,N_544,In_1000);
nor U2702 (N_2702,In_550,N_1138);
or U2703 (N_2703,N_1426,N_1698);
xnor U2704 (N_2704,N_1705,N_682);
and U2705 (N_2705,N_949,In_354);
and U2706 (N_2706,In_3098,In_1927);
nor U2707 (N_2707,N_806,In_2959);
xnor U2708 (N_2708,N_1405,N_1943);
xor U2709 (N_2709,N_15,N_1033);
nor U2710 (N_2710,In_527,N_540);
and U2711 (N_2711,In_2855,In_4889);
nand U2712 (N_2712,N_83,N_1318);
nor U2713 (N_2713,N_9,In_4001);
xnor U2714 (N_2714,In_4286,In_4318);
nor U2715 (N_2715,In_3078,In_2429);
and U2716 (N_2716,In_2388,In_4020);
nand U2717 (N_2717,In_4681,N_1104);
nand U2718 (N_2718,N_1351,In_1576);
and U2719 (N_2719,N_474,In_4431);
nor U2720 (N_2720,N_1451,N_1235);
and U2721 (N_2721,N_897,N_983);
xor U2722 (N_2722,N_1056,N_327);
nand U2723 (N_2723,N_938,In_340);
nand U2724 (N_2724,N_12,N_1984);
nor U2725 (N_2725,In_4143,In_849);
and U2726 (N_2726,N_449,N_1739);
and U2727 (N_2727,N_404,N_1378);
xor U2728 (N_2728,N_1122,In_2284);
nor U2729 (N_2729,In_327,N_958);
nand U2730 (N_2730,N_1148,N_1319);
nor U2731 (N_2731,N_1812,N_1692);
xor U2732 (N_2732,In_4100,N_1057);
nand U2733 (N_2733,N_1843,In_4983);
nor U2734 (N_2734,N_1734,N_548);
xor U2735 (N_2735,N_1340,In_3812);
or U2736 (N_2736,N_1439,In_2646);
nor U2737 (N_2737,In_876,N_1303);
nand U2738 (N_2738,N_1596,In_3434);
and U2739 (N_2739,N_1861,In_210);
nor U2740 (N_2740,In_942,N_870);
xor U2741 (N_2741,N_426,N_1074);
and U2742 (N_2742,In_4336,In_2175);
or U2743 (N_2743,N_673,N_1640);
and U2744 (N_2744,N_857,N_1994);
nor U2745 (N_2745,In_3365,N_212);
nor U2746 (N_2746,In_3334,N_1666);
nor U2747 (N_2747,N_545,N_175);
nand U2748 (N_2748,N_1060,N_1187);
nand U2749 (N_2749,N_1912,N_763);
nand U2750 (N_2750,In_1639,In_172);
nor U2751 (N_2751,N_24,In_4847);
or U2752 (N_2752,In_1651,In_3914);
nor U2753 (N_2753,N_92,N_909);
xnor U2754 (N_2754,N_1205,In_2196);
and U2755 (N_2755,N_1846,N_759);
nand U2756 (N_2756,N_214,N_89);
nor U2757 (N_2757,In_4668,N_1556);
or U2758 (N_2758,N_193,N_1833);
nor U2759 (N_2759,In_2929,In_1253);
and U2760 (N_2760,N_1751,In_162);
nor U2761 (N_2761,In_4689,In_4159);
nand U2762 (N_2762,In_1361,N_1183);
nor U2763 (N_2763,N_1433,N_228);
or U2764 (N_2764,N_121,In_1129);
nor U2765 (N_2765,N_567,N_981);
nand U2766 (N_2766,N_1193,N_271);
nand U2767 (N_2767,In_3070,N_219);
nor U2768 (N_2768,N_1976,In_4171);
xor U2769 (N_2769,N_571,N_1474);
and U2770 (N_2770,In_1820,N_1658);
and U2771 (N_2771,In_80,In_3617);
or U2772 (N_2772,N_40,N_1473);
nor U2773 (N_2773,N_638,N_810);
nor U2774 (N_2774,In_4848,N_374);
and U2775 (N_2775,N_889,N_381);
nor U2776 (N_2776,N_1175,N_1551);
xor U2777 (N_2777,In_2495,In_2739);
nand U2778 (N_2778,N_382,N_239);
nor U2779 (N_2779,In_1490,In_1994);
nor U2780 (N_2780,N_829,N_1741);
or U2781 (N_2781,N_1964,In_4820);
or U2782 (N_2782,N_1794,N_97);
and U2783 (N_2783,N_166,N_1750);
or U2784 (N_2784,In_1962,N_1952);
and U2785 (N_2785,N_1648,N_1307);
xnor U2786 (N_2786,N_1252,In_4638);
xor U2787 (N_2787,N_707,N_1153);
xnor U2788 (N_2788,In_1493,In_120);
nand U2789 (N_2789,N_871,In_2010);
nand U2790 (N_2790,In_1505,In_2058);
nand U2791 (N_2791,N_807,N_355);
nor U2792 (N_2792,In_427,N_1139);
and U2793 (N_2793,In_444,In_4570);
nand U2794 (N_2794,N_533,N_232);
nand U2795 (N_2795,N_1553,N_863);
nor U2796 (N_2796,In_2227,N_741);
nor U2797 (N_2797,N_1907,N_1851);
nor U2798 (N_2798,N_1273,N_1229);
nand U2799 (N_2799,N_945,In_4608);
nand U2800 (N_2800,N_551,N_13);
xor U2801 (N_2801,N_59,N_1781);
nand U2802 (N_2802,N_1533,N_991);
xor U2803 (N_2803,In_7,N_1953);
nor U2804 (N_2804,N_769,N_1326);
and U2805 (N_2805,In_2209,N_1547);
nor U2806 (N_2806,N_1595,In_715);
xnor U2807 (N_2807,N_1633,N_1576);
nor U2808 (N_2808,N_173,In_1283);
or U2809 (N_2809,In_2552,In_2217);
nand U2810 (N_2810,N_1536,N_1534);
or U2811 (N_2811,In_2938,N_734);
nor U2812 (N_2812,N_516,N_802);
or U2813 (N_2813,N_588,N_1141);
xnor U2814 (N_2814,In_1393,N_354);
and U2815 (N_2815,In_2029,In_2883);
or U2816 (N_2816,N_1701,N_1859);
or U2817 (N_2817,N_1935,In_1244);
and U2818 (N_2818,N_617,N_509);
xor U2819 (N_2819,N_419,N_110);
or U2820 (N_2820,In_1251,N_1630);
or U2821 (N_2821,N_316,N_1643);
xor U2822 (N_2822,N_1106,N_54);
xor U2823 (N_2823,In_3013,N_1218);
and U2824 (N_2824,N_1568,N_19);
nor U2825 (N_2825,In_1597,In_1641);
nand U2826 (N_2826,N_1789,In_4777);
nand U2827 (N_2827,N_853,N_1386);
nor U2828 (N_2828,N_1593,N_771);
nand U2829 (N_2829,In_4302,N_661);
and U2830 (N_2830,N_1267,N_816);
or U2831 (N_2831,N_1928,N_648);
nor U2832 (N_2832,N_1845,N_256);
or U2833 (N_2833,N_1855,In_2459);
nand U2834 (N_2834,N_163,N_1488);
and U2835 (N_2835,N_1266,N_822);
xor U2836 (N_2836,In_253,In_3009);
xor U2837 (N_2837,N_736,In_1313);
or U2838 (N_2838,N_906,N_1772);
nand U2839 (N_2839,In_4700,N_1050);
or U2840 (N_2840,N_207,N_1492);
nand U2841 (N_2841,N_1461,N_1067);
or U2842 (N_2842,N_1353,In_4372);
and U2843 (N_2843,N_1946,N_778);
nor U2844 (N_2844,In_2615,In_3985);
or U2845 (N_2845,N_421,In_4963);
xor U2846 (N_2846,N_1957,In_561);
and U2847 (N_2847,In_924,N_1000);
nand U2848 (N_2848,In_1480,N_1291);
nor U2849 (N_2849,In_2420,N_1111);
or U2850 (N_2850,In_4108,N_689);
nor U2851 (N_2851,N_698,N_672);
xor U2852 (N_2852,N_1951,N_1585);
nand U2853 (N_2853,N_1052,In_2082);
and U2854 (N_2854,N_6,N_1948);
and U2855 (N_2855,In_303,N_319);
nor U2856 (N_2856,N_371,N_828);
xor U2857 (N_2857,N_29,N_1746);
and U2858 (N_2858,In_4160,In_3864);
nor U2859 (N_2859,In_3745,N_1484);
or U2860 (N_2860,N_835,N_1806);
or U2861 (N_2861,N_993,N_1784);
and U2862 (N_2862,N_1347,In_313);
or U2863 (N_2863,N_1840,N_1700);
nand U2864 (N_2864,N_1763,N_150);
nor U2865 (N_2865,In_3699,N_61);
nor U2866 (N_2866,N_37,N_1737);
nor U2867 (N_2867,N_1310,N_1894);
nor U2868 (N_2868,N_1501,N_430);
nor U2869 (N_2869,In_3458,N_69);
and U2870 (N_2870,N_30,N_349);
and U2871 (N_2871,N_653,N_120);
nand U2872 (N_2872,In_1150,N_918);
nor U2873 (N_2873,N_1131,In_555);
or U2874 (N_2874,N_1004,In_3156);
nand U2875 (N_2875,N_1142,In_398);
or U2876 (N_2876,N_22,In_1144);
and U2877 (N_2877,N_1893,N_1870);
and U2878 (N_2878,N_46,N_1936);
and U2879 (N_2879,N_1809,In_2074);
or U2880 (N_2880,N_1231,N_616);
and U2881 (N_2881,N_324,In_1125);
or U2882 (N_2882,In_4749,N_1035);
nor U2883 (N_2883,N_542,In_4610);
xor U2884 (N_2884,N_1634,N_1339);
or U2885 (N_2885,N_1792,In_962);
or U2886 (N_2886,N_446,N_1435);
nor U2887 (N_2887,N_1684,N_756);
nand U2888 (N_2888,In_2653,N_1753);
and U2889 (N_2889,N_70,In_2992);
xnor U2890 (N_2890,N_96,N_1699);
xnor U2891 (N_2891,N_553,N_293);
xnor U2892 (N_2892,N_129,In_2638);
and U2893 (N_2893,N_1305,N_963);
nand U2894 (N_2894,In_4545,N_1302);
xnor U2895 (N_2895,N_229,N_818);
and U2896 (N_2896,N_1217,N_351);
or U2897 (N_2897,In_3344,In_2605);
nor U2898 (N_2898,In_1557,In_1638);
xnor U2899 (N_2899,N_510,In_3667);
nand U2900 (N_2900,N_1211,N_1168);
and U2901 (N_2901,In_3388,N_445);
or U2902 (N_2902,N_1423,In_4391);
nor U2903 (N_2903,N_1927,In_3733);
nand U2904 (N_2904,N_1317,In_1953);
nor U2905 (N_2905,In_3369,N_312);
nor U2906 (N_2906,N_1159,N_570);
or U2907 (N_2907,N_439,N_470);
xor U2908 (N_2908,N_1930,N_108);
xor U2909 (N_2909,In_1069,N_1853);
and U2910 (N_2910,N_775,N_931);
nand U2911 (N_2911,In_3583,In_3700);
or U2912 (N_2912,N_1624,N_397);
and U2913 (N_2913,In_3116,N_1707);
nor U2914 (N_2914,N_1125,N_456);
nand U2915 (N_2915,In_3199,N_1619);
or U2916 (N_2916,In_4659,N_1877);
xnor U2917 (N_2917,In_1023,In_2721);
and U2918 (N_2918,N_1716,N_1173);
nor U2919 (N_2919,N_434,N_1712);
or U2920 (N_2920,In_311,N_1906);
and U2921 (N_2921,N_652,N_1016);
xnor U2922 (N_2922,In_4122,In_606);
nand U2923 (N_2923,N_1005,N_982);
xnor U2924 (N_2924,In_2764,In_4414);
and U2925 (N_2925,N_1891,In_696);
or U2926 (N_2926,N_1956,In_3161);
and U2927 (N_2927,N_343,In_3470);
and U2928 (N_2928,N_1311,N_429);
and U2929 (N_2929,N_436,In_4244);
and U2930 (N_2930,N_1995,N_1207);
or U2931 (N_2931,In_2569,N_1670);
xor U2932 (N_2932,N_1600,N_1637);
xor U2933 (N_2933,N_902,N_376);
nand U2934 (N_2934,N_1440,N_1091);
or U2935 (N_2935,N_1355,N_1937);
or U2936 (N_2936,N_1586,In_4833);
or U2937 (N_2937,N_1258,N_66);
and U2938 (N_2938,N_1489,N_990);
xnor U2939 (N_2939,N_1275,N_790);
and U2940 (N_2940,N_1899,N_851);
nand U2941 (N_2941,In_3664,N_1399);
and U2942 (N_2942,N_1134,N_1565);
nand U2943 (N_2943,N_1116,In_3922);
xnor U2944 (N_2944,N_727,In_264);
nor U2945 (N_2945,N_919,N_729);
and U2946 (N_2946,N_1102,N_1667);
xor U2947 (N_2947,N_606,N_1081);
or U2948 (N_2948,In_4321,N_789);
nand U2949 (N_2949,In_913,N_861);
and U2950 (N_2950,In_4764,In_3061);
xnor U2951 (N_2951,N_1702,N_161);
xnor U2952 (N_2952,N_1432,In_3082);
xor U2953 (N_2953,In_2732,In_2398);
xor U2954 (N_2954,N_899,In_3909);
and U2955 (N_2955,N_329,N_713);
xnor U2956 (N_2956,N_451,N_884);
or U2957 (N_2957,N_1603,N_432);
xor U2958 (N_2958,N_1103,In_4976);
xor U2959 (N_2959,N_1723,In_1957);
nand U2960 (N_2960,N_1797,N_463);
and U2961 (N_2961,N_1372,In_4558);
nor U2962 (N_2962,N_1542,In_3055);
xor U2963 (N_2963,N_91,N_1306);
nand U2964 (N_2964,N_1110,N_1659);
and U2965 (N_2965,N_1714,N_1494);
nor U2966 (N_2966,In_1442,N_1032);
nor U2967 (N_2967,N_1747,N_1083);
nand U2968 (N_2968,In_1058,In_1353);
nor U2969 (N_2969,N_1988,N_866);
nor U2970 (N_2970,N_1282,In_731);
nand U2971 (N_2971,N_111,N_1034);
or U2972 (N_2972,N_487,In_3251);
xnor U2973 (N_2973,In_3817,N_1973);
and U2974 (N_2974,In_4799,N_396);
and U2975 (N_2975,In_4454,N_1244);
nand U2976 (N_2976,In_711,N_723);
xor U2977 (N_2977,In_4084,N_389);
and U2978 (N_2978,In_3186,In_2437);
xor U2979 (N_2979,N_336,In_728);
and U2980 (N_2980,In_2350,In_1324);
nand U2981 (N_2981,In_260,N_1237);
nand U2982 (N_2982,N_891,In_0);
and U2983 (N_2983,N_710,In_4975);
xnor U2984 (N_2984,N_215,N_1981);
nor U2985 (N_2985,N_330,N_1842);
xnor U2986 (N_2986,N_888,In_91);
and U2987 (N_2987,In_956,N_21);
nand U2988 (N_2988,In_126,N_1202);
and U2989 (N_2989,In_1464,In_4907);
xnor U2990 (N_2990,In_480,N_833);
nand U2991 (N_2991,N_1863,N_427);
nand U2992 (N_2992,N_1790,N_279);
or U2993 (N_2993,N_764,N_14);
xor U2994 (N_2994,In_4947,N_745);
nor U2995 (N_2995,N_1901,N_1760);
xor U2996 (N_2996,N_242,In_1246);
nor U2997 (N_2997,In_2258,In_4110);
xnor U2998 (N_2998,In_1062,N_1911);
nand U2999 (N_2999,In_1636,N_1271);
nand U3000 (N_3000,N_801,N_1068);
or U3001 (N_3001,N_1622,N_773);
and U3002 (N_3002,N_1902,In_2354);
xor U3003 (N_3003,N_196,In_1181);
xnor U3004 (N_3004,N_1166,N_1309);
and U3005 (N_3005,N_961,N_1818);
or U3006 (N_3006,In_2297,N_1515);
nor U3007 (N_3007,N_1980,N_574);
xor U3008 (N_3008,N_1051,In_3496);
and U3009 (N_3009,In_5,N_959);
nand U3010 (N_3010,N_1006,N_67);
nor U3011 (N_3011,In_2595,In_4451);
or U3012 (N_3012,In_756,N_805);
and U3013 (N_3013,In_3643,N_1729);
and U3014 (N_3014,N_415,N_1795);
nor U3015 (N_3015,In_2521,N_364);
and U3016 (N_3016,N_518,N_1);
and U3017 (N_3017,N_1966,In_4347);
nand U3018 (N_3018,N_1216,In_3726);
or U3019 (N_3019,N_1444,N_997);
nor U3020 (N_3020,In_975,In_1132);
nor U3021 (N_3021,N_240,N_926);
and U3022 (N_3022,In_1555,N_299);
and U3023 (N_3023,N_1872,N_1337);
nand U3024 (N_3024,In_3263,In_2381);
nand U3025 (N_3025,N_584,In_3277);
and U3026 (N_3026,N_1419,N_23);
and U3027 (N_3027,In_4447,N_140);
nand U3028 (N_3028,N_596,In_1795);
and U3029 (N_3029,In_4242,N_1496);
nor U3030 (N_3030,N_281,In_1051);
and U3031 (N_3031,N_119,In_4506);
nand U3032 (N_3032,N_1608,In_4734);
and U3033 (N_3033,N_941,In_853);
xor U3034 (N_3034,In_202,N_1063);
nand U3035 (N_3035,N_1368,In_1888);
or U3036 (N_3036,N_1087,N_1799);
nor U3037 (N_3037,In_2604,N_946);
and U3038 (N_3038,In_1950,N_735);
nand U3039 (N_3039,N_942,In_584);
or U3040 (N_3040,N_1292,In_993);
xnor U3041 (N_3041,In_3083,In_2299);
or U3042 (N_3042,In_1183,In_4583);
and U3043 (N_3043,N_465,N_1885);
xor U3044 (N_3044,N_1918,N_639);
or U3045 (N_3045,In_3798,N_1917);
xor U3046 (N_3046,N_1808,In_3291);
nand U3047 (N_3047,In_2481,N_1827);
or U3048 (N_3048,N_1955,N_1929);
and U3049 (N_3049,N_1801,In_4812);
and U3050 (N_3050,N_0,N_1278);
xor U3051 (N_3051,N_791,N_1581);
and U3052 (N_3052,N_1058,In_2198);
nor U3053 (N_3053,N_1230,N_586);
nor U3054 (N_3054,N_1838,In_248);
or U3055 (N_3055,N_715,In_2995);
nor U3056 (N_3056,N_368,N_1284);
or U3057 (N_3057,N_777,N_1577);
xnor U3058 (N_3058,N_697,N_160);
nor U3059 (N_3059,N_230,N_1715);
nand U3060 (N_3060,N_1500,In_3580);
xnor U3061 (N_3061,In_1871,In_4952);
xnor U3062 (N_3062,N_323,N_254);
nand U3063 (N_3063,N_2,N_1541);
nor U3064 (N_3064,N_468,N_1375);
nor U3065 (N_3065,N_1665,In_64);
xor U3066 (N_3066,N_369,N_1071);
or U3067 (N_3067,N_1938,In_1743);
nor U3068 (N_3068,N_1301,N_643);
xor U3069 (N_3069,In_1652,N_109);
nor U3070 (N_3070,In_1308,In_85);
or U3071 (N_3071,N_1685,In_441);
xnor U3072 (N_3072,N_1097,In_3550);
xor U3073 (N_3073,N_867,N_1270);
or U3074 (N_3074,In_672,In_1205);
nand U3075 (N_3075,N_48,N_1971);
xor U3076 (N_3076,N_1606,N_1875);
or U3077 (N_3077,N_688,In_2224);
and U3078 (N_3078,N_1198,N_1383);
or U3079 (N_3079,In_4237,N_383);
nand U3080 (N_3080,In_820,N_1803);
or U3081 (N_3081,In_4933,In_2114);
nor U3082 (N_3082,N_943,N_541);
xor U3083 (N_3083,N_987,N_1592);
nor U3084 (N_3084,In_4166,N_1308);
and U3085 (N_3085,N_675,N_1524);
nor U3086 (N_3086,N_420,N_1434);
nor U3087 (N_3087,N_1296,In_2085);
xnor U3088 (N_3088,In_321,N_1047);
xor U3089 (N_3089,N_76,In_2950);
and U3090 (N_3090,N_130,N_1241);
xor U3091 (N_3091,N_711,N_151);
xnor U3092 (N_3092,N_1395,N_272);
nand U3093 (N_3093,N_1628,In_4697);
nand U3094 (N_3094,N_502,N_1546);
or U3095 (N_3095,In_821,In_44);
and U3096 (N_3096,N_631,In_4400);
or U3097 (N_3097,N_1454,N_913);
nand U3098 (N_3098,In_1532,In_4565);
and U3099 (N_3099,N_910,In_3412);
xnor U3100 (N_3100,N_992,N_115);
xnor U3101 (N_3101,N_1415,N_1890);
nor U3102 (N_3102,N_513,N_1176);
or U3103 (N_3103,N_1145,N_969);
xor U3104 (N_3104,N_900,In_3869);
and U3105 (N_3105,N_1639,In_2208);
and U3106 (N_3106,N_1940,N_642);
nand U3107 (N_3107,In_3600,N_795);
nor U3108 (N_3108,In_3046,N_133);
and U3109 (N_3109,N_1921,N_1627);
nand U3110 (N_3110,N_591,N_1876);
xor U3111 (N_3111,N_624,N_155);
nand U3112 (N_3112,N_339,N_473);
or U3113 (N_3113,N_1728,N_1225);
nand U3114 (N_3114,N_1481,N_154);
and U3115 (N_3115,In_2017,N_1113);
and U3116 (N_3116,N_842,N_552);
or U3117 (N_3117,In_3360,N_1507);
or U3118 (N_3118,N_1497,N_1369);
xnor U3119 (N_3119,N_1635,N_678);
nand U3120 (N_3120,N_767,In_4158);
nand U3121 (N_3121,In_3248,In_3519);
and U3122 (N_3122,N_1379,In_2044);
or U3123 (N_3123,N_532,N_925);
and U3124 (N_3124,N_1631,In_4044);
nor U3125 (N_3125,N_824,N_252);
or U3126 (N_3126,In_1212,N_522);
or U3127 (N_3127,N_95,N_1121);
or U3128 (N_3128,In_1622,In_621);
nand U3129 (N_3129,N_677,N_1535);
or U3130 (N_3130,N_494,In_1997);
and U3131 (N_3131,N_1649,N_1689);
nand U3132 (N_3132,N_1341,In_2106);
and U3133 (N_3133,N_1228,In_4770);
xnor U3134 (N_3134,N_985,N_1315);
nand U3135 (N_3135,N_1852,N_1463);
nor U3136 (N_3136,N_1926,In_419);
and U3137 (N_3137,N_1029,In_896);
nor U3138 (N_3138,N_1208,N_1817);
nor U3139 (N_3139,N_1793,N_1589);
nand U3140 (N_3140,In_1744,N_1078);
xnor U3141 (N_3141,N_17,N_1156);
or U3142 (N_3142,N_840,N_1849);
and U3143 (N_3143,In_934,N_1356);
xnor U3144 (N_3144,N_1119,N_874);
and U3145 (N_3145,N_1656,N_1374);
nor U3146 (N_3146,N_608,N_438);
nand U3147 (N_3147,N_217,In_1224);
xnor U3148 (N_3148,In_1407,N_1752);
xor U3149 (N_3149,N_1214,N_403);
nand U3150 (N_3150,N_377,N_253);
nor U3151 (N_3151,N_159,N_269);
or U3152 (N_3152,N_1837,In_2762);
or U3153 (N_3153,In_3407,N_366);
xnor U3154 (N_3154,In_2321,N_1246);
nor U3155 (N_3155,N_683,N_146);
nand U3156 (N_3156,N_549,N_850);
and U3157 (N_3157,N_603,N_760);
and U3158 (N_3158,N_1297,In_3146);
xnor U3159 (N_3159,In_2353,N_739);
nand U3160 (N_3160,N_1972,In_283);
xnor U3161 (N_3161,N_495,N_1867);
xor U3162 (N_3162,N_826,N_1764);
or U3163 (N_3163,In_4745,N_227);
and U3164 (N_3164,N_537,In_2430);
xnor U3165 (N_3165,N_717,N_705);
nand U3166 (N_3166,N_879,N_1522);
nor U3167 (N_3167,In_2178,In_2018);
nand U3168 (N_3168,N_1437,In_1099);
or U3169 (N_3169,N_671,N_493);
or U3170 (N_3170,In_629,In_1933);
or U3171 (N_3171,N_455,N_1804);
or U3172 (N_3172,N_42,N_1573);
or U3173 (N_3173,N_1394,N_1391);
nand U3174 (N_3174,N_1416,In_4925);
nand U3175 (N_3175,N_1998,N_1462);
or U3176 (N_3176,N_1268,In_763);
xnor U3177 (N_3177,In_3014,N_1105);
nand U3178 (N_3178,N_890,N_972);
or U3179 (N_3179,N_774,N_282);
nor U3180 (N_3180,N_157,In_3201);
and U3181 (N_3181,N_1647,In_2858);
or U3182 (N_3182,N_712,In_2608);
nand U3183 (N_3183,In_2162,In_3844);
and U3184 (N_3184,In_1761,N_598);
nor U3185 (N_3185,In_1903,N_1333);
xor U3186 (N_3186,N_394,N_80);
nand U3187 (N_3187,N_989,In_4546);
nor U3188 (N_3188,N_36,N_255);
or U3189 (N_3189,N_226,N_64);
nand U3190 (N_3190,N_1506,N_1012);
nand U3191 (N_3191,In_4953,In_3556);
nor U3192 (N_3192,In_1228,In_1786);
xnor U3193 (N_3193,In_2013,N_435);
xor U3194 (N_3194,N_1719,In_1623);
and U3195 (N_3195,N_1609,In_2533);
xor U3196 (N_3196,In_3912,N_964);
nor U3197 (N_3197,N_1545,In_4212);
xor U3198 (N_3198,N_1904,N_165);
and U3199 (N_3199,In_174,N_1735);
xor U3200 (N_3200,N_1913,In_1057);
and U3201 (N_3201,N_1671,N_951);
xnor U3202 (N_3202,N_896,N_1404);
xnor U3203 (N_3203,N_856,N_1127);
and U3204 (N_3204,In_2446,N_1276);
and U3205 (N_3205,N_921,N_1129);
nand U3206 (N_3206,N_908,N_485);
or U3207 (N_3207,In_3475,N_1874);
or U3208 (N_3208,N_1503,In_3084);
nand U3209 (N_3209,N_1962,In_2579);
xor U3210 (N_3210,In_4459,In_2276);
nand U3211 (N_3211,In_3769,N_1446);
nor U3212 (N_3212,N_127,In_3427);
nand U3213 (N_3213,N_1422,N_690);
or U3214 (N_3214,N_1828,In_4931);
xnor U3215 (N_3215,N_1126,N_1174);
nor U3216 (N_3216,In_2688,In_314);
or U3217 (N_3217,N_1791,In_4503);
nand U3218 (N_3218,N_1236,In_3315);
nor U3219 (N_3219,N_1336,N_1709);
nand U3220 (N_3220,In_564,N_924);
nand U3221 (N_3221,N_1710,In_2988);
xnor U3222 (N_3222,N_291,N_139);
xnor U3223 (N_3223,N_1089,In_707);
nor U3224 (N_3224,In_4072,In_2621);
nand U3225 (N_3225,N_213,N_1882);
xnor U3226 (N_3226,N_1645,N_691);
or U3227 (N_3227,In_2933,N_716);
nand U3228 (N_3228,N_244,N_258);
nor U3229 (N_3229,N_326,N_566);
and U3230 (N_3230,N_1003,N_304);
xnor U3231 (N_3231,In_1851,In_2582);
or U3232 (N_3232,N_843,N_1644);
xor U3233 (N_3233,N_1150,N_1540);
nand U3234 (N_3234,N_101,N_1350);
nor U3235 (N_3235,N_85,N_288);
xor U3236 (N_3236,N_1479,N_1402);
or U3237 (N_3237,In_2452,In_888);
and U3238 (N_3238,In_2194,In_870);
or U3239 (N_3239,N_1611,In_1402);
and U3240 (N_3240,In_960,In_1115);
nor U3241 (N_3241,In_3685,In_4187);
nand U3242 (N_3242,N_1390,N_132);
nand U3243 (N_3243,N_1830,In_1007);
or U3244 (N_3244,N_1329,N_1664);
nor U3245 (N_3245,In_4498,N_1549);
nand U3246 (N_3246,N_1787,In_3374);
or U3247 (N_3247,N_1362,N_667);
nand U3248 (N_3248,In_534,In_4632);
xor U3249 (N_3249,N_102,N_1642);
or U3250 (N_3250,N_1243,In_1943);
nand U3251 (N_3251,N_1382,In_4868);
nor U3252 (N_3252,N_201,N_948);
nor U3253 (N_3253,N_1380,In_1988);
and U3254 (N_3254,N_295,N_1771);
nor U3255 (N_3255,In_3472,N_1604);
or U3256 (N_3256,In_3972,N_275);
and U3257 (N_3257,N_203,N_103);
or U3258 (N_3258,N_578,In_147);
xor U3259 (N_3259,In_1066,N_962);
and U3260 (N_3260,N_11,N_1048);
nand U3261 (N_3261,N_1881,In_2066);
and U3262 (N_3262,In_2469,N_1076);
and U3263 (N_3263,In_4991,N_1162);
xnor U3264 (N_3264,N_634,In_440);
or U3265 (N_3265,N_1839,N_1886);
or U3266 (N_3266,N_405,N_1115);
and U3267 (N_3267,In_4070,In_2499);
xor U3268 (N_3268,In_1696,N_402);
or U3269 (N_3269,In_2357,N_1939);
or U3270 (N_3270,N_1985,In_4197);
or U3271 (N_3271,In_4290,N_605);
xor U3272 (N_3272,N_1429,N_1693);
or U3273 (N_3273,In_3304,N_1453);
xnor U3274 (N_3274,N_887,In_3400);
xor U3275 (N_3275,N_1571,In_1902);
and U3276 (N_3276,In_4911,N_808);
or U3277 (N_3277,N_1304,In_1163);
and U3278 (N_3278,N_579,N_876);
nor U3279 (N_3279,In_1861,N_757);
and U3280 (N_3280,In_3845,N_412);
nor U3281 (N_3281,N_575,N_1182);
nand U3282 (N_3282,N_481,N_1274);
or U3283 (N_3283,N_332,N_1223);
nand U3284 (N_3284,N_1410,N_1602);
and U3285 (N_3285,N_352,N_1220);
nand U3286 (N_3286,N_1085,In_873);
nor U3287 (N_3287,N_932,In_720);
nand U3288 (N_3288,N_869,N_831);
and U3289 (N_3289,In_4917,In_3768);
xor U3290 (N_3290,In_49,In_2587);
nor U3291 (N_3291,In_4455,N_222);
and U3292 (N_3292,N_1457,N_1970);
nor U3293 (N_3293,N_762,N_1598);
and U3294 (N_3294,N_754,N_320);
xnor U3295 (N_3295,N_1476,In_4441);
nand U3296 (N_3296,N_1277,N_530);
or U3297 (N_3297,N_627,In_139);
and U3298 (N_3298,In_2525,N_1989);
nand U3299 (N_3299,In_3452,N_1475);
nor U3300 (N_3300,N_466,In_2020);
xnor U3301 (N_3301,N_395,N_55);
or U3302 (N_3302,N_568,N_289);
or U3303 (N_3303,N_1030,N_1293);
nor U3304 (N_3304,In_3823,N_832);
and U3305 (N_3305,N_32,N_1161);
and U3306 (N_3306,N_1080,In_952);
nand U3307 (N_3307,In_3328,N_344);
or U3308 (N_3308,N_1022,In_2902);
xnor U3309 (N_3309,N_1525,N_1019);
nand U3310 (N_3310,N_77,In_1247);
and U3311 (N_3311,N_1254,N_538);
or U3312 (N_3312,In_824,N_1366);
nand U3313 (N_3313,In_3911,In_1036);
and U3314 (N_3314,In_1468,N_1370);
xor U3315 (N_3315,N_126,In_3944);
or U3316 (N_3316,N_251,N_1934);
nand U3317 (N_3317,In_4112,In_1465);
nand U3318 (N_3318,N_1583,N_1933);
xnor U3319 (N_3319,In_6,N_1513);
nor U3320 (N_3320,N_278,N_820);
and U3321 (N_3321,N_572,In_4897);
and U3322 (N_3322,N_1856,In_1033);
or U3323 (N_3323,N_680,N_1036);
nand U3324 (N_3324,N_261,N_1300);
nor U3325 (N_3325,N_1189,In_2467);
or U3326 (N_3326,N_243,N_1754);
xnor U3327 (N_3327,In_1065,N_1017);
xnor U3328 (N_3328,N_1279,N_1128);
xnor U3329 (N_3329,In_1732,In_1601);
nor U3330 (N_3330,In_4082,N_409);
nor U3331 (N_3331,N_1835,N_331);
xor U3332 (N_3332,N_259,In_466);
and U3333 (N_3333,In_3551,In_3867);
or U3334 (N_3334,N_787,N_849);
nand U3335 (N_3335,N_1359,In_1461);
and U3336 (N_3336,N_1294,N_346);
nor U3337 (N_3337,N_1045,N_1195);
xnor U3338 (N_3338,N_313,N_1200);
and U3339 (N_3339,N_1222,N_266);
xnor U3340 (N_3340,In_3142,N_79);
xnor U3341 (N_3341,N_1011,N_1654);
nand U3342 (N_3342,N_342,N_1537);
or U3343 (N_3343,In_4129,N_1841);
xor U3344 (N_3344,In_1935,N_392);
xor U3345 (N_3345,N_286,N_507);
or U3346 (N_3346,In_831,In_1400);
or U3347 (N_3347,In_3113,In_1102);
xor U3348 (N_3348,N_662,N_1857);
and U3349 (N_3349,N_1834,N_595);
or U3350 (N_3350,N_1251,In_4849);
xor U3351 (N_3351,In_4346,N_1982);
and U3352 (N_3352,N_885,In_1609);
nor U3353 (N_3353,N_1086,In_3822);
or U3354 (N_3354,N_525,In_1138);
or U3355 (N_3355,N_1413,In_2310);
nor U3356 (N_3356,N_1974,N_1407);
and U3357 (N_3357,In_1249,N_1204);
nand U3358 (N_3358,In_2285,N_669);
xor U3359 (N_3359,N_1201,N_176);
xor U3360 (N_3360,N_1530,N_1373);
nor U3361 (N_3361,N_695,In_2656);
nor U3362 (N_3362,In_421,N_1732);
or U3363 (N_3363,In_521,N_94);
nor U3364 (N_3364,N_784,N_1721);
nor U3365 (N_3365,N_798,N_681);
and U3366 (N_3366,N_719,N_685);
nand U3367 (N_3367,N_1897,In_4428);
or U3368 (N_3368,N_236,N_5);
nand U3369 (N_3369,N_1092,In_329);
nor U3370 (N_3370,In_1577,N_1146);
nor U3371 (N_3371,N_1376,N_1820);
and U3372 (N_3372,N_1569,N_665);
nand U3373 (N_3373,N_52,N_1013);
or U3374 (N_3374,N_898,In_1822);
or U3375 (N_3375,In_3237,In_2635);
or U3376 (N_3376,In_2674,In_3438);
xor U3377 (N_3377,In_1736,In_1653);
nor U3378 (N_3378,In_3253,N_428);
and U3379 (N_3379,N_233,N_1544);
nand U3380 (N_3380,In_3631,N_1123);
or U3381 (N_3381,In_4292,In_1931);
or U3382 (N_3382,N_197,In_1661);
and U3383 (N_3383,In_2788,N_702);
xor U3384 (N_3384,In_1232,N_1037);
nand U3385 (N_3385,N_630,N_693);
nand U3386 (N_3386,N_480,N_1652);
nor U3387 (N_3387,In_4161,N_1255);
and U3388 (N_3388,In_114,In_837);
nor U3389 (N_3389,N_1312,N_81);
nor U3390 (N_3390,In_4830,N_1186);
nand U3391 (N_3391,N_1179,In_2032);
nand U3392 (N_3392,In_1835,In_404);
or U3393 (N_3393,In_2192,In_3897);
nand U3394 (N_3394,In_2489,N_1221);
nand U3395 (N_3395,In_651,N_1385);
nand U3396 (N_3396,N_628,N_1253);
nand U3397 (N_3397,N_928,In_2005);
or U3398 (N_3398,N_184,N_1810);
xnor U3399 (N_3399,N_813,In_1842);
and U3400 (N_3400,In_4092,N_865);
xor U3401 (N_3401,N_321,N_1858);
and U3402 (N_3402,In_1397,In_2814);
nand U3403 (N_3403,N_425,In_1006);
nor U3404 (N_3404,N_901,N_338);
or U3405 (N_3405,In_2493,N_225);
nor U3406 (N_3406,N_1136,N_1562);
nand U3407 (N_3407,N_860,In_4439);
and U3408 (N_3408,N_284,N_1023);
and U3409 (N_3409,N_1824,N_1290);
nand U3410 (N_3410,N_1364,N_1295);
or U3411 (N_3411,N_153,N_1815);
nor U3412 (N_3412,In_27,N_994);
nor U3413 (N_3413,N_1331,N_422);
or U3414 (N_3414,N_476,N_328);
nor U3415 (N_3415,N_687,In_4240);
nor U3416 (N_3416,In_3799,In_411);
nor U3417 (N_3417,In_3637,N_1487);
xor U3418 (N_3418,N_1742,N_1388);
nor U3419 (N_3419,N_950,N_800);
nand U3420 (N_3420,In_4348,N_823);
nor U3421 (N_3421,N_1135,N_1466);
xnor U3422 (N_3422,N_440,N_581);
xor U3423 (N_3423,N_172,N_686);
xnor U3424 (N_3424,In_2848,N_1748);
xnor U3425 (N_3425,N_600,N_1888);
nor U3426 (N_3426,N_1009,N_514);
or U3427 (N_3427,N_1424,N_453);
and U3428 (N_3428,N_1055,N_1330);
nor U3429 (N_3429,In_1451,N_1143);
xor U3430 (N_3430,N_1164,N_895);
and U3431 (N_3431,N_1261,N_751);
nor U3432 (N_3432,N_1997,N_1460);
nor U3433 (N_3433,In_2165,N_839);
and U3434 (N_3434,In_4518,N_73);
xor U3435 (N_3435,N_1717,In_2221);
nand U3436 (N_3436,In_2626,N_1096);
xor U3437 (N_3437,N_1610,In_3030);
nand U3438 (N_3438,N_1695,In_783);
and U3439 (N_3439,N_280,N_647);
xor U3440 (N_3440,N_98,N_907);
xor U3441 (N_3441,N_731,N_56);
nand U3442 (N_3442,In_2311,In_3555);
nand U3443 (N_3443,N_912,N_1612);
and U3444 (N_3444,N_580,N_464);
or U3445 (N_3445,N_621,N_158);
nor U3446 (N_3446,N_1805,N_504);
nor U3447 (N_3447,N_334,N_1864);
nor U3448 (N_3448,N_1564,In_4881);
nor U3449 (N_3449,In_342,In_1321);
nand U3450 (N_3450,In_2138,In_3330);
or U3451 (N_3451,N_1392,N_488);
or U3452 (N_3452,N_651,In_3788);
and U3453 (N_3453,N_1088,N_883);
or U3454 (N_3454,N_1224,In_1921);
and U3455 (N_3455,N_872,In_2564);
xor U3456 (N_3456,In_2640,In_3063);
xor U3457 (N_3457,N_1910,In_2391);
nand U3458 (N_3458,N_1686,N_894);
nor U3459 (N_3459,N_920,N_1160);
xor U3460 (N_3460,N_1010,In_3701);
or U3461 (N_3461,In_2168,N_367);
nand U3462 (N_3462,N_583,N_766);
nor U3463 (N_3463,In_484,In_4839);
nor U3464 (N_3464,N_1613,N_183);
nand U3465 (N_3465,In_113,N_1298);
or U3466 (N_3466,N_1672,N_206);
nor U3467 (N_3467,N_147,N_1281);
xor U3468 (N_3468,In_4338,N_450);
nor U3469 (N_3469,In_3111,N_740);
and U3470 (N_3470,N_398,N_1900);
nor U3471 (N_3471,N_933,In_236);
nand U3472 (N_3472,N_1140,N_817);
and U3473 (N_3473,N_1158,In_2817);
xor U3474 (N_3474,N_770,N_1149);
xor U3475 (N_3475,In_655,In_1961);
or U3476 (N_3476,N_143,In_2024);
nor U3477 (N_3477,N_623,N_679);
nor U3478 (N_3478,N_359,N_503);
xnor U3479 (N_3479,In_2565,In_3783);
xor U3480 (N_3480,In_3724,In_2442);
xnor U3481 (N_3481,N_33,N_1077);
and U3482 (N_3482,In_1909,N_640);
or U3483 (N_3483,N_1527,N_341);
or U3484 (N_3484,N_1287,N_1768);
and U3485 (N_3485,N_597,N_1107);
nand U3486 (N_3486,N_1703,In_493);
xor U3487 (N_3487,In_4273,N_1607);
or U3488 (N_3488,N_1860,In_628);
nor U3489 (N_3489,N_1758,In_3097);
nor U3490 (N_3490,N_211,In_944);
and U3491 (N_3491,N_308,In_2776);
and U3492 (N_3492,In_4067,In_2503);
or U3493 (N_3493,In_368,N_837);
xor U3494 (N_3494,In_3423,N_447);
xor U3495 (N_3495,N_1084,In_1275);
nand U3496 (N_3496,In_617,N_1332);
or U3497 (N_3497,N_529,N_1486);
nor U3498 (N_3498,N_721,N_350);
or U3499 (N_3499,N_1777,In_2411);
nand U3500 (N_3500,N_1663,In_4447);
or U3501 (N_3501,In_2017,N_503);
nor U3502 (N_3502,N_1475,N_1607);
xor U3503 (N_3503,N_1688,N_1908);
and U3504 (N_3504,N_1355,N_1570);
and U3505 (N_3505,N_1742,N_83);
or U3506 (N_3506,N_1704,In_2310);
xor U3507 (N_3507,N_1547,In_3413);
nand U3508 (N_3508,N_163,N_1963);
nand U3509 (N_3509,N_795,N_340);
or U3510 (N_3510,In_617,N_381);
nor U3511 (N_3511,N_1530,N_1217);
or U3512 (N_3512,N_22,N_361);
xnor U3513 (N_3513,N_514,N_1417);
or U3514 (N_3514,N_1112,N_1894);
or U3515 (N_3515,N_327,In_2357);
nand U3516 (N_3516,N_339,In_1203);
and U3517 (N_3517,N_789,N_1068);
and U3518 (N_3518,N_1804,N_1347);
or U3519 (N_3519,N_1370,N_1627);
nand U3520 (N_3520,N_936,N_1520);
nand U3521 (N_3521,N_1749,N_1086);
nor U3522 (N_3522,In_3875,In_4809);
or U3523 (N_3523,N_1620,N_1186);
nor U3524 (N_3524,N_422,N_1806);
nand U3525 (N_3525,N_1068,N_1207);
or U3526 (N_3526,In_831,N_1169);
and U3527 (N_3527,N_1361,N_19);
nor U3528 (N_3528,In_1609,N_1787);
nor U3529 (N_3529,N_1924,N_773);
nor U3530 (N_3530,N_415,N_981);
nand U3531 (N_3531,N_1727,In_739);
nor U3532 (N_3532,N_806,In_411);
nor U3533 (N_3533,In_2221,In_50);
and U3534 (N_3534,N_593,N_1721);
xor U3535 (N_3535,N_245,N_339);
or U3536 (N_3536,In_1618,N_115);
nor U3537 (N_3537,N_1400,In_3199);
xnor U3538 (N_3538,N_546,N_747);
or U3539 (N_3539,N_244,In_4318);
nand U3540 (N_3540,In_818,N_262);
nand U3541 (N_3541,In_4147,N_906);
and U3542 (N_3542,In_1256,N_905);
and U3543 (N_3543,In_2548,In_3475);
or U3544 (N_3544,In_2234,N_33);
nand U3545 (N_3545,In_1515,N_1724);
or U3546 (N_3546,N_886,N_914);
and U3547 (N_3547,In_1205,In_3000);
nor U3548 (N_3548,N_1623,In_1888);
xor U3549 (N_3549,In_3472,N_1322);
and U3550 (N_3550,N_211,N_1666);
xor U3551 (N_3551,N_455,N_648);
xor U3552 (N_3552,N_1364,N_605);
nor U3553 (N_3553,N_328,In_3289);
nand U3554 (N_3554,N_1952,N_1702);
nor U3555 (N_3555,N_71,N_517);
nor U3556 (N_3556,In_311,N_1374);
or U3557 (N_3557,N_1882,N_824);
or U3558 (N_3558,N_666,In_2032);
and U3559 (N_3559,N_1737,In_3452);
nand U3560 (N_3560,N_1342,In_1651);
and U3561 (N_3561,N_1455,N_1638);
nand U3562 (N_3562,N_309,In_3556);
xor U3563 (N_3563,In_975,N_1164);
or U3564 (N_3564,In_1423,In_4931);
nor U3565 (N_3565,N_707,In_3202);
nor U3566 (N_3566,In_1066,In_3441);
nand U3567 (N_3567,N_1368,In_1091);
nand U3568 (N_3568,N_1735,In_3344);
or U3569 (N_3569,N_318,In_880);
or U3570 (N_3570,N_1044,N_1489);
and U3571 (N_3571,N_35,N_369);
nor U3572 (N_3572,N_1847,In_2337);
and U3573 (N_3573,In_2475,N_954);
xnor U3574 (N_3574,N_1635,In_3724);
or U3575 (N_3575,N_1792,N_1853);
nand U3576 (N_3576,N_561,N_749);
xor U3577 (N_3577,N_1583,In_4418);
nand U3578 (N_3578,In_106,N_1788);
and U3579 (N_3579,In_2074,N_319);
and U3580 (N_3580,N_591,N_746);
and U3581 (N_3581,N_46,N_573);
xor U3582 (N_3582,In_2728,In_3132);
or U3583 (N_3583,N_9,In_466);
and U3584 (N_3584,In_3475,In_743);
or U3585 (N_3585,N_1834,In_4356);
or U3586 (N_3586,N_1091,In_1244);
nor U3587 (N_3587,N_1422,N_246);
xor U3588 (N_3588,In_3909,N_84);
xor U3589 (N_3589,N_1713,N_661);
and U3590 (N_3590,In_278,N_1298);
and U3591 (N_3591,N_1646,N_1502);
xnor U3592 (N_3592,In_4569,N_11);
nor U3593 (N_3593,N_314,N_1237);
xnor U3594 (N_3594,N_1790,In_3070);
nand U3595 (N_3595,N_1284,In_4348);
or U3596 (N_3596,N_1782,In_350);
xor U3597 (N_3597,N_1804,In_2595);
or U3598 (N_3598,N_644,In_1950);
or U3599 (N_3599,In_2114,In_1850);
nor U3600 (N_3600,N_31,N_801);
and U3601 (N_3601,N_1381,N_1883);
or U3602 (N_3602,N_1456,N_749);
or U3603 (N_3603,N_1828,N_1592);
xor U3604 (N_3604,N_1684,In_2815);
xnor U3605 (N_3605,N_1916,In_174);
and U3606 (N_3606,In_3427,N_1770);
and U3607 (N_3607,N_1815,In_96);
and U3608 (N_3608,N_809,N_1218);
or U3609 (N_3609,N_999,In_4212);
xnor U3610 (N_3610,N_1717,N_334);
nand U3611 (N_3611,In_3014,N_705);
nand U3612 (N_3612,In_2908,N_1537);
nor U3613 (N_3613,N_1436,N_255);
and U3614 (N_3614,In_3046,In_2638);
nor U3615 (N_3615,N_1604,N_54);
or U3616 (N_3616,N_1040,N_1048);
or U3617 (N_3617,In_2465,N_496);
nor U3618 (N_3618,N_589,N_1432);
and U3619 (N_3619,N_986,N_1634);
xnor U3620 (N_3620,N_1105,N_1824);
xor U3621 (N_3621,N_742,In_3199);
nand U3622 (N_3622,N_1628,N_1028);
and U3623 (N_3623,In_3911,N_794);
nand U3624 (N_3624,N_1216,In_4425);
and U3625 (N_3625,N_464,N_1893);
nor U3626 (N_3626,N_1258,In_3726);
xor U3627 (N_3627,N_976,N_396);
nor U3628 (N_3628,N_1243,N_1424);
xor U3629 (N_3629,N_1665,N_444);
nand U3630 (N_3630,N_177,In_2505);
xnor U3631 (N_3631,N_1970,N_745);
and U3632 (N_3632,N_1911,N_443);
xor U3633 (N_3633,In_3302,N_1119);
and U3634 (N_3634,N_1841,N_241);
and U3635 (N_3635,N_1847,In_1144);
nor U3636 (N_3636,N_356,N_911);
and U3637 (N_3637,N_1952,N_321);
xor U3638 (N_3638,In_651,N_1372);
xor U3639 (N_3639,In_837,N_1534);
xnor U3640 (N_3640,N_1848,N_1007);
xor U3641 (N_3641,N_952,N_287);
and U3642 (N_3642,N_761,N_1455);
nor U3643 (N_3643,N_1564,N_1783);
xor U3644 (N_3644,In_4638,N_818);
xnor U3645 (N_3645,N_1780,In_1629);
nor U3646 (N_3646,N_1524,N_350);
and U3647 (N_3647,N_311,N_808);
and U3648 (N_3648,In_975,In_2311);
nand U3649 (N_3649,In_1701,N_831);
nor U3650 (N_3650,N_1037,N_294);
nor U3651 (N_3651,N_651,N_626);
nand U3652 (N_3652,N_1127,N_577);
or U3653 (N_3653,N_21,N_1983);
or U3654 (N_3654,N_1226,N_1390);
or U3655 (N_3655,N_1938,In_2194);
or U3656 (N_3656,N_1837,In_3929);
xor U3657 (N_3657,N_248,In_3654);
nand U3658 (N_3658,N_283,N_947);
xnor U3659 (N_3659,N_1379,In_796);
and U3660 (N_3660,N_1402,N_994);
nand U3661 (N_3661,N_1164,N_733);
nand U3662 (N_3662,In_2674,N_671);
and U3663 (N_3663,N_6,N_1680);
and U3664 (N_3664,N_161,N_1130);
xnor U3665 (N_3665,In_2121,N_894);
and U3666 (N_3666,N_569,N_219);
nand U3667 (N_3667,In_2885,N_630);
nor U3668 (N_3668,N_419,N_1326);
nand U3669 (N_3669,N_1712,N_296);
nor U3670 (N_3670,In_4631,In_1676);
and U3671 (N_3671,N_800,N_1011);
nor U3672 (N_3672,In_3237,In_4977);
and U3673 (N_3673,In_4377,In_1961);
and U3674 (N_3674,N_403,N_217);
or U3675 (N_3675,N_379,N_1548);
and U3676 (N_3676,N_887,In_4160);
nand U3677 (N_3677,In_96,N_390);
nor U3678 (N_3678,N_173,N_526);
or U3679 (N_3679,In_1820,In_1480);
xor U3680 (N_3680,N_823,N_989);
xor U3681 (N_3681,N_1563,N_1444);
and U3682 (N_3682,N_681,In_711);
nor U3683 (N_3683,N_369,In_3161);
and U3684 (N_3684,In_4292,N_1073);
or U3685 (N_3685,N_143,N_1111);
xnor U3686 (N_3686,N_198,N_833);
xor U3687 (N_3687,In_3885,N_1820);
xnor U3688 (N_3688,N_1216,N_1625);
nand U3689 (N_3689,N_528,In_1473);
nor U3690 (N_3690,N_217,N_1339);
or U3691 (N_3691,In_2168,N_5);
xor U3692 (N_3692,N_91,N_1005);
or U3693 (N_3693,N_282,In_924);
nand U3694 (N_3694,In_2138,N_502);
and U3695 (N_3695,In_3845,N_1247);
or U3696 (N_3696,In_1480,N_969);
xnor U3697 (N_3697,N_313,In_3944);
nor U3698 (N_3698,In_1102,In_3994);
and U3699 (N_3699,N_1090,In_4898);
nor U3700 (N_3700,In_1051,N_1426);
nand U3701 (N_3701,N_779,In_1638);
nor U3702 (N_3702,N_1516,N_494);
xnor U3703 (N_3703,In_2114,In_4923);
xnor U3704 (N_3704,N_1214,In_1007);
and U3705 (N_3705,In_4346,N_1811);
or U3706 (N_3706,N_775,N_967);
nor U3707 (N_3707,In_534,In_3317);
or U3708 (N_3708,N_119,In_1313);
and U3709 (N_3709,N_1247,In_3468);
nand U3710 (N_3710,In_2888,N_680);
nor U3711 (N_3711,N_1602,In_1047);
or U3712 (N_3712,N_1334,In_1771);
nor U3713 (N_3713,In_3583,N_1732);
xor U3714 (N_3714,N_405,In_120);
and U3715 (N_3715,N_1730,In_1577);
or U3716 (N_3716,N_97,N_1313);
xnor U3717 (N_3717,N_1875,N_1163);
xnor U3718 (N_3718,N_422,N_97);
xnor U3719 (N_3719,In_64,N_1529);
nor U3720 (N_3720,In_1407,N_1170);
nor U3721 (N_3721,In_756,N_264);
or U3722 (N_3722,N_1021,N_1742);
nor U3723 (N_3723,N_1298,N_2);
or U3724 (N_3724,N_1569,N_180);
nor U3725 (N_3725,In_4622,N_1702);
and U3726 (N_3726,In_3791,N_1516);
xnor U3727 (N_3727,N_489,In_2992);
or U3728 (N_3728,N_171,In_4659);
and U3729 (N_3729,N_773,N_1165);
or U3730 (N_3730,N_548,N_1669);
nand U3731 (N_3731,N_262,N_1930);
xor U3732 (N_3732,In_4578,N_78);
or U3733 (N_3733,N_1900,N_1667);
xor U3734 (N_3734,N_46,N_1564);
xnor U3735 (N_3735,N_1082,N_398);
nand U3736 (N_3736,N_337,N_1608);
xor U3737 (N_3737,In_4975,N_712);
and U3738 (N_3738,N_64,In_3199);
or U3739 (N_3739,In_2587,N_1985);
nand U3740 (N_3740,N_1062,N_1936);
and U3741 (N_3741,N_1197,N_1926);
xor U3742 (N_3742,N_174,In_4602);
or U3743 (N_3743,In_2640,In_4350);
xor U3744 (N_3744,N_1479,N_1120);
nor U3745 (N_3745,N_1761,N_1777);
nand U3746 (N_3746,In_1026,In_4890);
and U3747 (N_3747,N_357,N_774);
nand U3748 (N_3748,N_385,N_1114);
nand U3749 (N_3749,In_2357,In_1125);
nor U3750 (N_3750,N_1828,In_783);
or U3751 (N_3751,N_1344,N_839);
and U3752 (N_3752,In_1058,N_546);
nand U3753 (N_3753,N_1829,In_822);
or U3754 (N_3754,In_3643,N_1556);
or U3755 (N_3755,N_1019,N_603);
nor U3756 (N_3756,N_599,In_3202);
nor U3757 (N_3757,N_1581,N_1278);
or U3758 (N_3758,N_935,In_1442);
and U3759 (N_3759,N_913,In_3198);
and U3760 (N_3760,N_1687,In_2764);
or U3761 (N_3761,N_1696,In_561);
or U3762 (N_3762,N_16,N_1644);
nor U3763 (N_3763,In_2120,N_281);
nand U3764 (N_3764,In_3886,N_587);
nor U3765 (N_3765,N_163,N_668);
nor U3766 (N_3766,N_952,In_2311);
nand U3767 (N_3767,N_938,N_299);
nor U3768 (N_3768,In_4122,N_424);
or U3769 (N_3769,N_1478,In_2548);
nand U3770 (N_3770,N_516,In_93);
and U3771 (N_3771,N_1364,In_4622);
xnor U3772 (N_3772,N_1354,In_4558);
and U3773 (N_3773,N_1969,N_1223);
nand U3774 (N_3774,N_1530,N_1197);
and U3775 (N_3775,In_1251,N_303);
nand U3776 (N_3776,In_1933,In_2489);
nand U3777 (N_3777,N_1532,N_1686);
or U3778 (N_3778,N_141,N_1618);
xor U3779 (N_3779,In_957,In_1815);
nand U3780 (N_3780,N_630,In_1514);
and U3781 (N_3781,N_1701,N_1089);
nand U3782 (N_3782,N_1843,N_1701);
xor U3783 (N_3783,N_1261,In_1047);
nand U3784 (N_3784,In_2815,N_249);
or U3785 (N_3785,N_396,N_1659);
nor U3786 (N_3786,N_675,N_685);
or U3787 (N_3787,N_1695,N_1371);
nor U3788 (N_3788,N_1536,In_3922);
xnor U3789 (N_3789,N_953,In_2688);
and U3790 (N_3790,N_1805,N_474);
nor U3791 (N_3791,N_1957,N_899);
and U3792 (N_3792,In_4903,N_368);
or U3793 (N_3793,N_988,N_1983);
or U3794 (N_3794,N_1176,N_1733);
nand U3795 (N_3795,N_372,In_3922);
or U3796 (N_3796,N_1866,N_852);
nand U3797 (N_3797,N_1860,N_677);
or U3798 (N_3798,In_3098,N_286);
xor U3799 (N_3799,N_1161,N_1093);
or U3800 (N_3800,In_3570,N_397);
nor U3801 (N_3801,In_2858,N_1643);
nand U3802 (N_3802,In_4326,N_725);
or U3803 (N_3803,N_1767,In_63);
nor U3804 (N_3804,In_4814,N_879);
xor U3805 (N_3805,In_3519,In_2121);
xnor U3806 (N_3806,In_3132,N_275);
nand U3807 (N_3807,N_1256,N_248);
nor U3808 (N_3808,N_1706,In_1661);
xor U3809 (N_3809,N_576,N_1883);
nor U3810 (N_3810,In_756,N_902);
nand U3811 (N_3811,N_1355,In_3654);
or U3812 (N_3812,N_869,N_810);
nor U3813 (N_3813,In_534,In_2525);
or U3814 (N_3814,N_598,N_276);
or U3815 (N_3815,In_2759,In_3600);
or U3816 (N_3816,N_1479,N_1320);
nand U3817 (N_3817,In_3698,N_292);
xor U3818 (N_3818,N_539,N_694);
xnor U3819 (N_3819,In_1784,In_4451);
or U3820 (N_3820,In_4084,In_1655);
xnor U3821 (N_3821,N_1044,N_1512);
or U3822 (N_3822,N_233,In_2727);
nand U3823 (N_3823,N_469,In_1473);
nand U3824 (N_3824,In_2081,In_2468);
xnor U3825 (N_3825,N_1814,In_4344);
nand U3826 (N_3826,N_66,N_275);
nor U3827 (N_3827,N_1817,N_1995);
xor U3828 (N_3828,In_3360,In_50);
nand U3829 (N_3829,In_4384,In_4161);
nand U3830 (N_3830,N_155,N_1513);
xnor U3831 (N_3831,In_236,N_1612);
and U3832 (N_3832,In_3716,In_1353);
or U3833 (N_3833,In_3700,N_656);
or U3834 (N_3834,N_1613,N_1327);
nor U3835 (N_3835,N_1299,N_1335);
nor U3836 (N_3836,N_864,N_1453);
or U3837 (N_3837,In_1514,N_849);
nand U3838 (N_3838,N_734,N_1197);
nand U3839 (N_3839,In_2598,In_285);
or U3840 (N_3840,N_1201,N_324);
or U3841 (N_3841,In_1888,In_3644);
nand U3842 (N_3842,In_1651,N_331);
xor U3843 (N_3843,In_2058,N_24);
and U3844 (N_3844,In_2781,In_2373);
and U3845 (N_3845,In_3911,N_1230);
or U3846 (N_3846,N_1229,In_1038);
nor U3847 (N_3847,N_869,N_1240);
nor U3848 (N_3848,In_3900,N_1306);
nor U3849 (N_3849,N_725,N_1800);
or U3850 (N_3850,In_2465,N_1935);
or U3851 (N_3851,In_2074,N_44);
or U3852 (N_3852,N_152,In_2224);
nand U3853 (N_3853,In_253,In_440);
or U3854 (N_3854,N_1931,N_1747);
nor U3855 (N_3855,N_848,N_251);
nor U3856 (N_3856,N_480,In_667);
nor U3857 (N_3857,N_1223,N_1541);
xor U3858 (N_3858,In_3277,In_3620);
nand U3859 (N_3859,In_1557,In_4063);
nor U3860 (N_3860,N_641,N_1422);
xor U3861 (N_3861,In_3099,N_1053);
and U3862 (N_3862,N_1997,N_1906);
nand U3863 (N_3863,N_508,N_66);
or U3864 (N_3864,In_4890,N_429);
xnor U3865 (N_3865,In_4020,N_559);
or U3866 (N_3866,N_1018,N_1965);
nor U3867 (N_3867,N_1240,N_1603);
nand U3868 (N_3868,N_577,N_1162);
and U3869 (N_3869,N_1528,N_1621);
or U3870 (N_3870,N_127,N_1609);
and U3871 (N_3871,N_1740,N_672);
or U3872 (N_3872,N_1873,N_778);
and U3873 (N_3873,In_3981,N_1956);
and U3874 (N_3874,N_1916,N_31);
and U3875 (N_3875,N_1395,In_1619);
nor U3876 (N_3876,N_906,In_2596);
nand U3877 (N_3877,In_90,N_1570);
nand U3878 (N_3878,N_1249,N_1089);
and U3879 (N_3879,In_2168,In_3583);
and U3880 (N_3880,N_1064,N_1786);
nand U3881 (N_3881,N_38,In_2297);
and U3882 (N_3882,N_1567,N_441);
nor U3883 (N_3883,N_32,In_311);
xnor U3884 (N_3884,N_1152,N_1694);
and U3885 (N_3885,N_1289,N_1740);
xor U3886 (N_3886,In_4100,N_1046);
and U3887 (N_3887,N_235,N_370);
xor U3888 (N_3888,N_913,N_1327);
xnor U3889 (N_3889,N_787,In_2360);
and U3890 (N_3890,In_1950,N_1381);
nand U3891 (N_3891,N_354,In_1943);
or U3892 (N_3892,N_1206,In_3788);
and U3893 (N_3893,In_4460,N_551);
xor U3894 (N_3894,N_1131,In_672);
xor U3895 (N_3895,In_4903,N_1534);
nor U3896 (N_3896,In_4044,N_1205);
and U3897 (N_3897,N_1222,In_4506);
or U3898 (N_3898,In_778,N_668);
xor U3899 (N_3899,N_1206,In_106);
nand U3900 (N_3900,In_1629,N_1706);
and U3901 (N_3901,N_1527,N_386);
or U3902 (N_3902,N_67,N_734);
xnor U3903 (N_3903,In_2262,N_1407);
or U3904 (N_3904,N_1595,N_1962);
nor U3905 (N_3905,In_1433,N_1006);
nor U3906 (N_3906,N_600,N_501);
or U3907 (N_3907,In_1945,N_518);
or U3908 (N_3908,In_2080,N_1524);
or U3909 (N_3909,N_1869,N_1326);
and U3910 (N_3910,N_1612,N_1058);
and U3911 (N_3911,N_1803,N_156);
nand U3912 (N_3912,In_2250,In_3908);
xnor U3913 (N_3913,In_2945,N_1305);
or U3914 (N_3914,N_101,In_3470);
nand U3915 (N_3915,N_254,N_1318);
nor U3916 (N_3916,N_1678,N_356);
xor U3917 (N_3917,N_811,N_1139);
or U3918 (N_3918,In_956,N_1248);
nor U3919 (N_3919,In_3315,N_1664);
or U3920 (N_3920,N_295,In_4655);
xnor U3921 (N_3921,N_1881,N_1283);
and U3922 (N_3922,N_400,In_2183);
or U3923 (N_3923,N_1939,In_1133);
xnor U3924 (N_3924,N_591,N_1268);
or U3925 (N_3925,In_313,In_2992);
xnor U3926 (N_3926,N_1889,N_1934);
or U3927 (N_3927,N_1538,N_30);
nor U3928 (N_3928,N_244,In_3685);
xnor U3929 (N_3929,N_1064,N_188);
nand U3930 (N_3930,N_506,N_915);
and U3931 (N_3931,N_1486,N_243);
nand U3932 (N_3932,N_969,N_250);
or U3933 (N_3933,N_595,N_926);
nand U3934 (N_3934,N_687,N_1916);
nand U3935 (N_3935,In_4503,N_104);
xor U3936 (N_3936,N_669,N_1790);
nor U3937 (N_3937,N_466,N_1787);
or U3938 (N_3938,N_1486,In_3823);
nor U3939 (N_3939,N_1391,N_766);
or U3940 (N_3940,N_192,N_354);
or U3941 (N_3941,N_582,N_636);
nand U3942 (N_3942,In_4745,In_1235);
or U3943 (N_3943,N_182,In_4147);
or U3944 (N_3944,N_102,In_3733);
or U3945 (N_3945,N_457,N_883);
nor U3946 (N_3946,N_956,N_465);
and U3947 (N_3947,N_1122,N_572);
and U3948 (N_3948,In_481,N_995);
xnor U3949 (N_3949,N_425,In_27);
or U3950 (N_3950,In_1306,N_1662);
or U3951 (N_3951,N_1859,N_1697);
and U3952 (N_3952,In_2781,N_925);
nand U3953 (N_3953,In_2670,N_144);
nor U3954 (N_3954,In_2537,N_1278);
or U3955 (N_3955,N_1549,N_1092);
or U3956 (N_3956,N_1625,N_298);
and U3957 (N_3957,N_307,N_327);
or U3958 (N_3958,N_164,N_523);
or U3959 (N_3959,In_4748,N_1036);
and U3960 (N_3960,N_1989,In_4663);
nand U3961 (N_3961,In_880,N_30);
nand U3962 (N_3962,In_2608,N_432);
nand U3963 (N_3963,In_4451,N_718);
and U3964 (N_3964,N_962,N_330);
xor U3965 (N_3965,N_930,In_3951);
nand U3966 (N_3966,N_459,N_340);
or U3967 (N_3967,N_865,N_928);
xor U3968 (N_3968,In_31,N_1241);
and U3969 (N_3969,N_1405,N_154);
or U3970 (N_3970,N_1829,N_621);
or U3971 (N_3971,N_941,In_3400);
nand U3972 (N_3972,In_3822,N_119);
or U3973 (N_3973,N_1628,N_757);
and U3974 (N_3974,N_816,N_958);
nand U3975 (N_3975,N_372,N_1890);
and U3976 (N_3976,In_1843,N_424);
nor U3977 (N_3977,N_1844,N_407);
and U3978 (N_3978,N_1264,N_1736);
nor U3979 (N_3979,N_1336,In_3329);
or U3980 (N_3980,N_1661,In_1283);
nor U3981 (N_3981,N_1015,In_1957);
nand U3982 (N_3982,N_1088,N_87);
nor U3983 (N_3983,N_1858,N_621);
nor U3984 (N_3984,N_201,N_533);
nand U3985 (N_3985,N_716,In_1038);
nor U3986 (N_3986,N_429,In_2276);
nor U3987 (N_3987,In_4414,N_632);
xor U3988 (N_3988,N_714,N_572);
or U3989 (N_3989,N_704,N_1092);
or U3990 (N_3990,N_278,N_1488);
nor U3991 (N_3991,N_189,N_1512);
and U3992 (N_3992,N_8,N_153);
xnor U3993 (N_3993,In_641,N_1757);
xnor U3994 (N_3994,N_1700,In_3611);
nor U3995 (N_3995,N_587,In_3198);
and U3996 (N_3996,N_259,N_924);
nor U3997 (N_3997,In_2486,N_1896);
and U3998 (N_3998,N_1104,In_4754);
and U3999 (N_3999,N_304,N_366);
nand U4000 (N_4000,N_2721,N_2002);
nor U4001 (N_4001,N_3417,N_2190);
nor U4002 (N_4002,N_2530,N_2816);
or U4003 (N_4003,N_2945,N_3238);
and U4004 (N_4004,N_3361,N_3609);
nand U4005 (N_4005,N_2381,N_3340);
or U4006 (N_4006,N_3073,N_2096);
nand U4007 (N_4007,N_3256,N_3621);
nand U4008 (N_4008,N_3865,N_2111);
or U4009 (N_4009,N_3393,N_3158);
nand U4010 (N_4010,N_2884,N_2378);
xor U4011 (N_4011,N_3444,N_2295);
nand U4012 (N_4012,N_2832,N_3831);
or U4013 (N_4013,N_2902,N_3607);
or U4014 (N_4014,N_3862,N_2586);
nor U4015 (N_4015,N_3034,N_3061);
or U4016 (N_4016,N_3431,N_3539);
nor U4017 (N_4017,N_2569,N_3412);
nor U4018 (N_4018,N_2421,N_2041);
xnor U4019 (N_4019,N_2162,N_2218);
nand U4020 (N_4020,N_3994,N_2666);
nand U4021 (N_4021,N_2213,N_2248);
or U4022 (N_4022,N_3722,N_3349);
nand U4023 (N_4023,N_2144,N_3681);
xor U4024 (N_4024,N_2799,N_2951);
or U4025 (N_4025,N_2452,N_2693);
nand U4026 (N_4026,N_2148,N_3491);
nor U4027 (N_4027,N_2632,N_2089);
and U4028 (N_4028,N_2384,N_2894);
nand U4029 (N_4029,N_3926,N_2793);
and U4030 (N_4030,N_2420,N_3072);
nand U4031 (N_4031,N_2099,N_2281);
xor U4032 (N_4032,N_2521,N_2581);
and U4033 (N_4033,N_3661,N_2734);
or U4034 (N_4034,N_3905,N_2761);
or U4035 (N_4035,N_2215,N_3744);
and U4036 (N_4036,N_3575,N_2081);
or U4037 (N_4037,N_3318,N_3648);
or U4038 (N_4038,N_2167,N_2287);
nand U4039 (N_4039,N_3578,N_3820);
or U4040 (N_4040,N_3800,N_2040);
xor U4041 (N_4041,N_3556,N_2824);
xnor U4042 (N_4042,N_2665,N_2448);
nand U4043 (N_4043,N_3778,N_2549);
nand U4044 (N_4044,N_3209,N_3967);
xor U4045 (N_4045,N_2214,N_3059);
xnor U4046 (N_4046,N_3891,N_2010);
or U4047 (N_4047,N_2819,N_3406);
nand U4048 (N_4048,N_2885,N_2102);
nor U4049 (N_4049,N_2482,N_3787);
and U4050 (N_4050,N_3021,N_3980);
xnor U4051 (N_4051,N_2490,N_2520);
nand U4052 (N_4052,N_3709,N_2327);
nand U4053 (N_4053,N_3784,N_3329);
nor U4054 (N_4054,N_2564,N_2151);
nand U4055 (N_4055,N_2636,N_3029);
nor U4056 (N_4056,N_3437,N_2686);
nand U4057 (N_4057,N_2079,N_2845);
nand U4058 (N_4058,N_2533,N_3599);
or U4059 (N_4059,N_3009,N_2515);
xnor U4060 (N_4060,N_3509,N_3813);
nand U4061 (N_4061,N_3631,N_3075);
xnor U4062 (N_4062,N_3094,N_3411);
or U4063 (N_4063,N_2787,N_2067);
nand U4064 (N_4064,N_3424,N_3514);
or U4065 (N_4065,N_3566,N_3670);
and U4066 (N_4066,N_2126,N_3789);
nand U4067 (N_4067,N_2639,N_2254);
nand U4068 (N_4068,N_3600,N_2688);
nor U4069 (N_4069,N_2472,N_2821);
nor U4070 (N_4070,N_3093,N_2669);
nor U4071 (N_4071,N_2791,N_3822);
nand U4072 (N_4072,N_3805,N_2119);
nor U4073 (N_4073,N_2414,N_2278);
or U4074 (N_4074,N_3258,N_2615);
nor U4075 (N_4075,N_2867,N_3292);
xnor U4076 (N_4076,N_2753,N_3903);
or U4077 (N_4077,N_2888,N_3794);
or U4078 (N_4078,N_2923,N_3595);
nor U4079 (N_4079,N_3137,N_2323);
nand U4080 (N_4080,N_2538,N_3825);
and U4081 (N_4081,N_3814,N_3931);
or U4082 (N_4082,N_3206,N_2455);
nand U4083 (N_4083,N_3821,N_3658);
and U4084 (N_4084,N_3022,N_2124);
nand U4085 (N_4085,N_3772,N_3752);
xor U4086 (N_4086,N_3742,N_3586);
and U4087 (N_4087,N_3512,N_2201);
and U4088 (N_4088,N_2267,N_2709);
nor U4089 (N_4089,N_2356,N_3763);
and U4090 (N_4090,N_2768,N_3558);
and U4091 (N_4091,N_2542,N_2778);
xnor U4092 (N_4092,N_3385,N_2519);
nor U4093 (N_4093,N_3957,N_3986);
and U4094 (N_4094,N_2260,N_2545);
nor U4095 (N_4095,N_3252,N_3155);
nand U4096 (N_4096,N_2018,N_2786);
nor U4097 (N_4097,N_2592,N_2765);
or U4098 (N_4098,N_3464,N_3019);
xor U4099 (N_4099,N_2391,N_2802);
nor U4100 (N_4100,N_3297,N_2350);
or U4101 (N_4101,N_3219,N_3516);
and U4102 (N_4102,N_2430,N_3795);
nand U4103 (N_4103,N_2413,N_3569);
xor U4104 (N_4104,N_2246,N_3220);
nor U4105 (N_4105,N_2337,N_2274);
xor U4106 (N_4106,N_3207,N_3978);
xnor U4107 (N_4107,N_3751,N_3223);
nand U4108 (N_4108,N_2282,N_3641);
or U4109 (N_4109,N_3462,N_3097);
nor U4110 (N_4110,N_2025,N_3843);
nand U4111 (N_4111,N_3036,N_3045);
xor U4112 (N_4112,N_3949,N_2959);
and U4113 (N_4113,N_2374,N_2966);
nor U4114 (N_4114,N_3904,N_2880);
nor U4115 (N_4115,N_3466,N_3131);
xor U4116 (N_4116,N_2322,N_2675);
or U4117 (N_4117,N_2813,N_3432);
nand U4118 (N_4118,N_2029,N_3783);
and U4119 (N_4119,N_3746,N_3878);
and U4120 (N_4120,N_3975,N_3369);
xnor U4121 (N_4121,N_2157,N_2423);
nand U4122 (N_4122,N_2409,N_3510);
xnor U4123 (N_4123,N_2974,N_2992);
xor U4124 (N_4124,N_2759,N_3737);
and U4125 (N_4125,N_3872,N_3448);
or U4126 (N_4126,N_3440,N_3495);
xnor U4127 (N_4127,N_3433,N_3506);
xor U4128 (N_4128,N_3119,N_3713);
and U4129 (N_4129,N_2840,N_2338);
nor U4130 (N_4130,N_3170,N_3705);
nand U4131 (N_4131,N_2092,N_2864);
and U4132 (N_4132,N_3798,N_2700);
nor U4133 (N_4133,N_2973,N_3912);
and U4134 (N_4134,N_3570,N_2020);
or U4135 (N_4135,N_3475,N_3511);
or U4136 (N_4136,N_2727,N_2606);
nor U4137 (N_4137,N_2780,N_3142);
nor U4138 (N_4138,N_2535,N_3041);
nand U4139 (N_4139,N_2971,N_3688);
nand U4140 (N_4140,N_2986,N_2645);
or U4141 (N_4141,N_2755,N_3345);
or U4142 (N_4142,N_2393,N_3161);
xnor U4143 (N_4143,N_2316,N_3243);
and U4144 (N_4144,N_2843,N_2475);
xnor U4145 (N_4145,N_2352,N_3567);
and U4146 (N_4146,N_3023,N_3049);
or U4147 (N_4147,N_2599,N_2294);
nor U4148 (N_4148,N_3043,N_2532);
xor U4149 (N_4149,N_3181,N_3327);
or U4150 (N_4150,N_3523,N_2345);
nor U4151 (N_4151,N_2366,N_3864);
xnor U4152 (N_4152,N_3758,N_2211);
and U4153 (N_4153,N_3754,N_2779);
nor U4154 (N_4154,N_2698,N_3188);
xor U4155 (N_4155,N_2620,N_3906);
xnor U4156 (N_4156,N_3897,N_2653);
nor U4157 (N_4157,N_2585,N_2706);
nor U4158 (N_4158,N_3973,N_2844);
and U4159 (N_4159,N_3468,N_3977);
or U4160 (N_4160,N_2596,N_2920);
xnor U4161 (N_4161,N_3502,N_2138);
or U4162 (N_4162,N_3480,N_3404);
and U4163 (N_4163,N_3262,N_3885);
xnor U4164 (N_4164,N_2749,N_2496);
nand U4165 (N_4165,N_2741,N_3900);
nor U4166 (N_4166,N_2720,N_2792);
nand U4167 (N_4167,N_3969,N_2582);
nor U4168 (N_4168,N_3067,N_2625);
nor U4169 (N_4169,N_2667,N_3488);
nor U4170 (N_4170,N_3056,N_2677);
nor U4171 (N_4171,N_2982,N_2747);
nor U4172 (N_4172,N_2663,N_3091);
xor U4173 (N_4173,N_2633,N_2271);
or U4174 (N_4174,N_2270,N_2106);
nor U4175 (N_4175,N_3372,N_2847);
and U4176 (N_4176,N_2199,N_2547);
nand U4177 (N_4177,N_2861,N_3186);
nor U4178 (N_4178,N_2371,N_3580);
nand U4179 (N_4179,N_3435,N_2283);
and U4180 (N_4180,N_3038,N_2760);
or U4181 (N_4181,N_3620,N_3302);
and U4182 (N_4182,N_2189,N_3081);
xor U4183 (N_4183,N_2155,N_2949);
nand U4184 (N_4184,N_2981,N_3453);
and U4185 (N_4185,N_3275,N_2970);
nor U4186 (N_4186,N_2094,N_3797);
xor U4187 (N_4187,N_3233,N_3529);
or U4188 (N_4188,N_2305,N_2221);
xnor U4189 (N_4189,N_2748,N_3144);
and U4190 (N_4190,N_2289,N_3637);
nor U4191 (N_4191,N_2554,N_3898);
xnor U4192 (N_4192,N_3837,N_2145);
nand U4193 (N_4193,N_2501,N_2220);
nand U4194 (N_4194,N_3070,N_3999);
xnor U4195 (N_4195,N_2480,N_2513);
and U4196 (N_4196,N_3627,N_3446);
xor U4197 (N_4197,N_3863,N_3384);
and U4198 (N_4198,N_2406,N_3652);
and U4199 (N_4199,N_2664,N_3443);
or U4200 (N_4200,N_3147,N_2397);
nor U4201 (N_4201,N_2756,N_3796);
nand U4202 (N_4202,N_2712,N_3806);
xor U4203 (N_4203,N_2197,N_3777);
xnor U4204 (N_4204,N_2929,N_2445);
or U4205 (N_4205,N_2650,N_3269);
xnor U4206 (N_4206,N_2173,N_3333);
and U4207 (N_4207,N_2196,N_2379);
and U4208 (N_4208,N_3343,N_2737);
and U4209 (N_4209,N_3151,N_2930);
xor U4210 (N_4210,N_2921,N_3968);
xnor U4211 (N_4211,N_3913,N_2723);
xor U4212 (N_4212,N_2132,N_2525);
nand U4213 (N_4213,N_2136,N_3769);
xnor U4214 (N_4214,N_3222,N_2928);
nand U4215 (N_4215,N_2955,N_3877);
nor U4216 (N_4216,N_2541,N_2178);
or U4217 (N_4217,N_2878,N_2736);
and U4218 (N_4218,N_2364,N_2691);
or U4219 (N_4219,N_3136,N_2114);
and U4220 (N_4220,N_2245,N_2516);
and U4221 (N_4221,N_3638,N_3519);
xnor U4222 (N_4222,N_2479,N_2320);
and U4223 (N_4223,N_2752,N_2926);
and U4224 (N_4224,N_2313,N_2526);
xnor U4225 (N_4225,N_2863,N_2105);
xnor U4226 (N_4226,N_3249,N_2250);
xor U4227 (N_4227,N_2838,N_3860);
and U4228 (N_4228,N_3952,N_3255);
or U4229 (N_4229,N_3571,N_3368);
and U4230 (N_4230,N_2023,N_3854);
xor U4231 (N_4231,N_3901,N_2122);
and U4232 (N_4232,N_2219,N_3234);
or U4233 (N_4233,N_3438,N_2163);
xnor U4234 (N_4234,N_2876,N_2314);
nand U4235 (N_4235,N_2217,N_2918);
xnor U4236 (N_4236,N_3665,N_3673);
xor U4237 (N_4237,N_3642,N_2623);
and U4238 (N_4238,N_3482,N_3757);
nand U4239 (N_4239,N_3392,N_3773);
and U4240 (N_4240,N_2910,N_3214);
or U4241 (N_4241,N_2093,N_2332);
xnor U4242 (N_4242,N_2416,N_2999);
nand U4243 (N_4243,N_2848,N_3005);
nand U4244 (N_4244,N_2846,N_3268);
xnor U4245 (N_4245,N_2771,N_3006);
nor U4246 (N_4246,N_2979,N_2401);
and U4247 (N_4247,N_2456,N_2470);
nor U4248 (N_4248,N_2689,N_2903);
nand U4249 (N_4249,N_2466,N_3185);
and U4250 (N_4250,N_2634,N_2643);
or U4251 (N_4251,N_3062,N_2298);
nand U4252 (N_4252,N_2039,N_3781);
nand U4253 (N_4253,N_3937,N_2830);
or U4254 (N_4254,N_2325,N_3407);
nor U4255 (N_4255,N_2508,N_3886);
xor U4256 (N_4256,N_2536,N_3166);
or U4257 (N_4257,N_2441,N_3914);
xor U4258 (N_4258,N_3715,N_2738);
nand U4259 (N_4259,N_3311,N_3313);
nor U4260 (N_4260,N_2263,N_3273);
and U4261 (N_4261,N_2383,N_2308);
or U4262 (N_4262,N_2785,N_3574);
nand U4263 (N_4263,N_2422,N_3762);
and U4264 (N_4264,N_3490,N_3321);
and U4265 (N_4265,N_3747,N_3902);
xor U4266 (N_4266,N_3749,N_2762);
xor U4267 (N_4267,N_2523,N_3615);
or U4268 (N_4268,N_3110,N_2656);
and U4269 (N_4269,N_3819,N_3471);
or U4270 (N_4270,N_2758,N_2621);
xor U4271 (N_4271,N_3373,N_2828);
nand U4272 (N_4272,N_3909,N_3092);
or U4273 (N_4273,N_2347,N_2091);
xor U4274 (N_4274,N_2563,N_3004);
or U4275 (N_4275,N_2601,N_3246);
and U4276 (N_4276,N_2499,N_2135);
and U4277 (N_4277,N_2980,N_3312);
nor U4278 (N_4278,N_3944,N_3958);
or U4279 (N_4279,N_3888,N_3871);
nand U4280 (N_4280,N_3672,N_2994);
or U4281 (N_4281,N_3013,N_3858);
xnor U4282 (N_4282,N_2370,N_3460);
nand U4283 (N_4283,N_2279,N_3071);
nor U4284 (N_4284,N_3267,N_2602);
xor U4285 (N_4285,N_3157,N_2548);
or U4286 (N_4286,N_2223,N_3782);
and U4287 (N_4287,N_3410,N_3236);
and U4288 (N_4288,N_2517,N_3786);
xnor U4289 (N_4289,N_2415,N_2154);
or U4290 (N_4290,N_3367,N_3699);
and U4291 (N_4291,N_3845,N_3533);
xnor U4292 (N_4292,N_2188,N_3046);
or U4293 (N_4293,N_3838,N_2035);
nor U4294 (N_4294,N_3643,N_3282);
and U4295 (N_4295,N_2184,N_2090);
and U4296 (N_4296,N_2403,N_3531);
or U4297 (N_4297,N_2587,N_3935);
or U4298 (N_4298,N_2382,N_3668);
or U4299 (N_4299,N_2806,N_2301);
xnor U4300 (N_4300,N_3981,N_2905);
or U4301 (N_4301,N_2005,N_2428);
and U4302 (N_4302,N_2775,N_2231);
xnor U4303 (N_4303,N_2056,N_3524);
or U4304 (N_4304,N_2065,N_2642);
or U4305 (N_4305,N_3946,N_2198);
nor U4306 (N_4306,N_3649,N_3603);
xnor U4307 (N_4307,N_3810,N_3581);
nand U4308 (N_4308,N_3577,N_3867);
nor U4309 (N_4309,N_3470,N_2690);
nand U4310 (N_4310,N_3703,N_2583);
nor U4311 (N_4311,N_2619,N_3265);
nand U4312 (N_4312,N_3010,N_2405);
nor U4313 (N_4313,N_2588,N_3505);
and U4314 (N_4314,N_3663,N_3376);
nor U4315 (N_4315,N_2553,N_3016);
nand U4316 (N_4316,N_2329,N_3254);
xor U4317 (N_4317,N_2754,N_2399);
xnor U4318 (N_4318,N_3695,N_3360);
nor U4319 (N_4319,N_3317,N_2612);
or U4320 (N_4320,N_3760,N_2075);
xnor U4321 (N_4321,N_2367,N_3096);
nor U4322 (N_4322,N_2156,N_3342);
and U4323 (N_4323,N_2942,N_3492);
nand U4324 (N_4324,N_2388,N_2941);
and U4325 (N_4325,N_3766,N_3244);
and U4326 (N_4326,N_2912,N_2509);
nand U4327 (N_4327,N_2212,N_2594);
xor U4328 (N_4328,N_3809,N_3150);
nor U4329 (N_4329,N_3889,N_2293);
or U4330 (N_4330,N_2899,N_3943);
and U4331 (N_4331,N_3674,N_3875);
or U4332 (N_4332,N_3960,N_2057);
nor U4333 (N_4333,N_2373,N_3039);
or U4334 (N_4334,N_2309,N_3543);
or U4335 (N_4335,N_3455,N_3160);
and U4336 (N_4336,N_2346,N_3149);
nor U4337 (N_4337,N_2227,N_3247);
nor U4338 (N_4338,N_3728,N_3076);
xor U4339 (N_4339,N_2365,N_2609);
and U4340 (N_4340,N_3008,N_3224);
and U4341 (N_4341,N_3759,N_2776);
and U4342 (N_4342,N_2757,N_2037);
nand U4343 (N_4343,N_2898,N_3288);
nand U4344 (N_4344,N_2872,N_2187);
nand U4345 (N_4345,N_2603,N_2299);
and U4346 (N_4346,N_2435,N_3228);
or U4347 (N_4347,N_2769,N_3442);
nor U4348 (N_4348,N_3454,N_3965);
nor U4349 (N_4349,N_3802,N_2823);
or U4350 (N_4350,N_3676,N_2070);
nand U4351 (N_4351,N_2875,N_3636);
and U4352 (N_4352,N_2186,N_3419);
nor U4353 (N_4353,N_3133,N_2084);
and U4354 (N_4354,N_2801,N_2043);
and U4355 (N_4355,N_2206,N_3387);
nor U4356 (N_4356,N_3679,N_3109);
nand U4357 (N_4357,N_2989,N_2082);
and U4358 (N_4358,N_2628,N_3537);
and U4359 (N_4359,N_3936,N_3833);
nor U4360 (N_4360,N_2476,N_2194);
xnor U4361 (N_4361,N_3741,N_3277);
xor U4362 (N_4362,N_3990,N_2534);
and U4363 (N_4363,N_2234,N_3919);
or U4364 (N_4364,N_2595,N_2465);
and U4365 (N_4365,N_3832,N_2247);
nand U4366 (N_4366,N_2764,N_2820);
nor U4367 (N_4367,N_2733,N_3353);
nand U4368 (N_4368,N_3176,N_3148);
nor U4369 (N_4369,N_2368,N_3692);
nand U4370 (N_4370,N_2210,N_3779);
nand U4371 (N_4371,N_3881,N_3196);
or U4372 (N_4372,N_2916,N_2777);
and U4373 (N_4373,N_3619,N_3316);
or U4374 (N_4374,N_3646,N_2662);
and U4375 (N_4375,N_3541,N_3325);
xor U4376 (N_4376,N_3352,N_3400);
xnor U4377 (N_4377,N_2265,N_3290);
nor U4378 (N_4378,N_2253,N_2304);
xnor U4379 (N_4379,N_2318,N_3684);
nand U4380 (N_4380,N_3130,N_2175);
nand U4381 (N_4381,N_3146,N_3685);
nor U4382 (N_4382,N_2728,N_2104);
nand U4383 (N_4383,N_3320,N_3606);
or U4384 (N_4384,N_2050,N_3476);
or U4385 (N_4385,N_3033,N_2637);
nand U4386 (N_4386,N_3211,N_3388);
nand U4387 (N_4387,N_3001,N_2209);
and U4388 (N_4388,N_2965,N_2121);
xnor U4389 (N_4389,N_3948,N_2125);
or U4390 (N_4390,N_2195,N_2681);
or U4391 (N_4391,N_3894,N_3184);
xor U4392 (N_4392,N_2788,N_2703);
xnor U4393 (N_4393,N_2975,N_2302);
nand U4394 (N_4394,N_3770,N_2054);
xnor U4395 (N_4395,N_3409,N_2931);
or U4396 (N_4396,N_3592,N_2897);
nand U4397 (N_4397,N_3811,N_3112);
nor U4398 (N_4398,N_3060,N_2351);
xnor U4399 (N_4399,N_2474,N_3610);
xnor U4400 (N_4400,N_3260,N_3927);
and U4401 (N_4401,N_3538,N_2960);
nand U4402 (N_4402,N_2537,N_2593);
nor U4403 (N_4403,N_2285,N_2730);
nor U4404 (N_4404,N_2348,N_3834);
nor U4405 (N_4405,N_3895,N_3079);
or U4406 (N_4406,N_2797,N_3295);
nand U4407 (N_4407,N_3635,N_2275);
or U4408 (N_4408,N_3044,N_3579);
nor U4409 (N_4409,N_2047,N_3378);
nand U4410 (N_4410,N_2722,N_2238);
or U4411 (N_4411,N_2837,N_2097);
or U4412 (N_4412,N_2166,N_3660);
nor U4413 (N_4413,N_3457,N_2735);
nor U4414 (N_4414,N_2454,N_3086);
nand U4415 (N_4415,N_2207,N_3874);
xor U4416 (N_4416,N_3107,N_3841);
xor U4417 (N_4417,N_3489,N_2937);
or U4418 (N_4418,N_3933,N_2419);
xnor U4419 (N_4419,N_3565,N_3594);
nor U4420 (N_4420,N_3487,N_3890);
nor U4421 (N_4421,N_3576,N_3279);
nand U4422 (N_4422,N_2746,N_3689);
xnor U4423 (N_4423,N_2203,N_3439);
nor U4424 (N_4424,N_3645,N_3322);
nand U4425 (N_4425,N_3963,N_3114);
nand U4426 (N_4426,N_2266,N_2062);
and U4427 (N_4427,N_3294,N_3711);
nor U4428 (N_4428,N_3231,N_2459);
and U4429 (N_4429,N_2064,N_3616);
nand U4430 (N_4430,N_3486,N_2176);
nand U4431 (N_4431,N_3633,N_2704);
and U4432 (N_4432,N_3750,N_3626);
nand U4433 (N_4433,N_3427,N_2659);
or U4434 (N_4434,N_2440,N_2372);
nor U4435 (N_4435,N_3467,N_3669);
xnor U4436 (N_4436,N_2944,N_3141);
nor U4437 (N_4437,N_2077,N_2361);
xnor U4438 (N_4438,N_2644,N_2386);
and U4439 (N_4439,N_2825,N_3630);
xor U4440 (N_4440,N_3377,N_3002);
or U4441 (N_4441,N_2969,N_2575);
nand U4442 (N_4442,N_3640,N_3852);
and U4443 (N_4443,N_2952,N_3598);
xor U4444 (N_4444,N_3954,N_3452);
or U4445 (N_4445,N_2240,N_2362);
and U4446 (N_4446,N_3835,N_2800);
nor U4447 (N_4447,N_2648,N_2244);
nand U4448 (N_4448,N_3479,N_3300);
xnor U4449 (N_4449,N_2953,N_3299);
nor U4450 (N_4450,N_3159,N_3793);
nand U4451 (N_4451,N_2377,N_3624);
and U4452 (N_4452,N_2657,N_2007);
and U4453 (N_4453,N_3463,N_3179);
nand U4454 (N_4454,N_3988,N_2584);
nand U4455 (N_4455,N_2781,N_2742);
nand U4456 (N_4456,N_3775,N_3680);
xor U4457 (N_4457,N_3792,N_2146);
nor U4458 (N_4458,N_3063,N_3985);
or U4459 (N_4459,N_3780,N_3966);
or U4460 (N_4460,N_3304,N_3804);
nand U4461 (N_4461,N_3162,N_3771);
and U4462 (N_4462,N_3426,N_3618);
and U4463 (N_4463,N_2672,N_2577);
or U4464 (N_4464,N_2446,N_2529);
xnor U4465 (N_4465,N_3589,N_2711);
and U4466 (N_4466,N_2006,N_3739);
nand U4467 (N_4467,N_3478,N_3920);
xnor U4468 (N_4468,N_2991,N_2607);
nor U4469 (N_4469,N_2985,N_2528);
nor U4470 (N_4470,N_3287,N_3704);
xnor U4471 (N_4471,N_3296,N_3551);
xor U4472 (N_4472,N_2336,N_3402);
xnor U4473 (N_4473,N_3164,N_2539);
and U4474 (N_4474,N_3562,N_2812);
or U4475 (N_4475,N_3723,N_2892);
nor U4476 (N_4476,N_3522,N_2164);
nand U4477 (N_4477,N_3106,N_2913);
and U4478 (N_4478,N_3706,N_2958);
nor U4479 (N_4479,N_3357,N_2964);
or U4480 (N_4480,N_3494,N_3261);
and U4481 (N_4481,N_2396,N_3899);
nand U4482 (N_4482,N_3507,N_3283);
or U4483 (N_4483,N_3216,N_2714);
nand U4484 (N_4484,N_2000,N_2012);
nand U4485 (N_4485,N_3208,N_2118);
nand U4486 (N_4486,N_2284,N_3257);
nor U4487 (N_4487,N_3213,N_2086);
and U4488 (N_4488,N_2264,N_2131);
or U4489 (N_4489,N_3917,N_3559);
nand U4490 (N_4490,N_2673,N_2193);
and U4491 (N_4491,N_2836,N_2158);
xor U4492 (N_4492,N_2321,N_2661);
xnor U4493 (N_4493,N_3582,N_2990);
xnor U4494 (N_4494,N_2058,N_2948);
xor U4495 (N_4495,N_2395,N_3032);
or U4496 (N_4496,N_3285,N_3396);
or U4497 (N_4497,N_2924,N_3712);
xnor U4498 (N_4498,N_3925,N_2502);
nor U4499 (N_4499,N_3099,N_3591);
nand U4500 (N_4500,N_3040,N_3687);
and U4501 (N_4501,N_3143,N_3276);
xor U4502 (N_4502,N_2063,N_2292);
or U4503 (N_4503,N_3694,N_2729);
nor U4504 (N_4504,N_3351,N_2032);
xnor U4505 (N_4505,N_2433,N_2022);
nand U4506 (N_4506,N_2319,N_2782);
or U4507 (N_4507,N_2552,N_2695);
nor U4508 (N_4508,N_2504,N_3116);
xor U4509 (N_4509,N_2483,N_3449);
nor U4510 (N_4510,N_2467,N_2249);
or U4511 (N_4511,N_3939,N_3953);
or U4512 (N_4512,N_3588,N_2556);
nor U4513 (N_4513,N_2555,N_3824);
or U4514 (N_4514,N_3278,N_2461);
and U4515 (N_4515,N_3028,N_3337);
nor U4516 (N_4516,N_3192,N_3259);
or U4517 (N_4517,N_3421,N_3286);
xnor U4518 (N_4518,N_2850,N_2457);
nor U4519 (N_4519,N_2597,N_3175);
and U4520 (N_4520,N_2579,N_2500);
nand U4521 (N_4521,N_2618,N_3896);
nand U4522 (N_4522,N_2795,N_2394);
and U4523 (N_4523,N_2349,N_3083);
nor U4524 (N_4524,N_2683,N_3272);
or U4525 (N_4525,N_3434,N_3270);
or U4526 (N_4526,N_2814,N_3650);
nor U4527 (N_4527,N_2524,N_3911);
or U4528 (N_4528,N_2859,N_3341);
or U4529 (N_4529,N_3550,N_2473);
or U4530 (N_4530,N_3065,N_3202);
nand U4531 (N_4531,N_3726,N_3177);
xor U4532 (N_4532,N_3271,N_2998);
or U4533 (N_4533,N_3128,N_3974);
xor U4534 (N_4534,N_2255,N_2616);
or U4535 (N_4535,N_2306,N_2315);
or U4536 (N_4536,N_2652,N_2268);
nand U4537 (N_4537,N_2589,N_2161);
xnor U4538 (N_4538,N_3035,N_3011);
xor U4539 (N_4539,N_3724,N_3493);
and U4540 (N_4540,N_2874,N_2507);
and U4541 (N_4541,N_3585,N_2076);
or U4542 (N_4542,N_2112,N_2068);
xnor U4543 (N_4543,N_3611,N_2447);
nor U4544 (N_4544,N_3846,N_2142);
and U4545 (N_4545,N_2947,N_2829);
xor U4546 (N_4546,N_2389,N_3215);
and U4547 (N_4547,N_2147,N_2463);
xnor U4548 (N_4548,N_3030,N_3861);
nor U4549 (N_4549,N_2794,N_2701);
and U4550 (N_4550,N_3557,N_2149);
nor U4551 (N_4551,N_3563,N_3774);
xor U4552 (N_4552,N_3363,N_2996);
nor U4553 (N_4553,N_2568,N_3849);
and U4554 (N_4554,N_3987,N_3517);
nor U4555 (N_4555,N_3857,N_2269);
and U4556 (N_4556,N_3623,N_2239);
nor U4557 (N_4557,N_2110,N_2572);
nand U4558 (N_4558,N_2276,N_3545);
xor U4559 (N_4559,N_2232,N_3807);
nor U4560 (N_4560,N_2494,N_2464);
nand U4561 (N_4561,N_3870,N_3066);
or U4562 (N_4562,N_3613,N_2512);
and U4563 (N_4563,N_2055,N_3102);
xnor U4564 (N_4564,N_3082,N_2716);
nand U4565 (N_4565,N_3205,N_2939);
and U4566 (N_4566,N_3138,N_2638);
xnor U4567 (N_4567,N_3441,N_3380);
nand U4568 (N_4568,N_2385,N_3000);
xnor U4569 (N_4569,N_2425,N_3907);
nor U4570 (N_4570,N_2481,N_3882);
nand U4571 (N_4571,N_3528,N_3791);
nand U4572 (N_4572,N_3513,N_3995);
nor U4573 (N_4573,N_2225,N_2439);
nand U4574 (N_4574,N_3229,N_3785);
xnor U4575 (N_4575,N_2493,N_3855);
or U4576 (N_4576,N_3942,N_2687);
nand U4577 (N_4577,N_2719,N_2976);
or U4578 (N_4578,N_2631,N_3803);
nor U4579 (N_4579,N_2886,N_2335);
nor U4580 (N_4580,N_2080,N_2855);
nand U4581 (N_4581,N_3564,N_3472);
and U4582 (N_4582,N_2339,N_2570);
and U4583 (N_4583,N_3374,N_2116);
nor U4584 (N_4584,N_2045,N_3928);
or U4585 (N_4585,N_2200,N_2139);
or U4586 (N_4586,N_3721,N_2078);
or U4587 (N_4587,N_3084,N_2497);
or U4588 (N_4588,N_3816,N_3915);
nor U4589 (N_4589,N_2604,N_3167);
and U4590 (N_4590,N_3193,N_3993);
nor U4591 (N_4591,N_3064,N_3733);
nand U4592 (N_4592,N_3548,N_3289);
xnor U4593 (N_4593,N_2817,N_2809);
nor U4594 (N_4594,N_3447,N_2137);
or U4595 (N_4595,N_3701,N_2685);
nor U4596 (N_4596,N_2877,N_3484);
xnor U4597 (N_4597,N_2444,N_3314);
or U4598 (N_4598,N_3173,N_3057);
and U4599 (N_4599,N_3568,N_2702);
or U4600 (N_4600,N_2858,N_3934);
and U4601 (N_4601,N_2103,N_2360);
and U4602 (N_4602,N_3702,N_2909);
nand U4603 (N_4603,N_3306,N_3959);
and U4604 (N_4604,N_2359,N_3540);
nor U4605 (N_4605,N_3929,N_2868);
nand U4606 (N_4606,N_3134,N_2426);
xor U4607 (N_4607,N_3430,N_2437);
or U4608 (N_4608,N_3940,N_3996);
and U4609 (N_4609,N_3250,N_3731);
nand U4610 (N_4610,N_3527,N_3127);
and U4611 (N_4611,N_3614,N_2016);
or U4612 (N_4612,N_2369,N_3251);
nand U4613 (N_4613,N_2766,N_2839);
and U4614 (N_4614,N_2561,N_3497);
and U4615 (N_4615,N_2036,N_2069);
or U4616 (N_4616,N_3239,N_2300);
nand U4617 (N_4617,N_3738,N_2705);
xor U4618 (N_4618,N_3020,N_3922);
nor U4619 (N_4619,N_3892,N_2049);
nand U4620 (N_4620,N_3970,N_3414);
xnor U4621 (N_4621,N_2804,N_2789);
and U4622 (N_4622,N_2297,N_2740);
and U4623 (N_4623,N_3827,N_2938);
or U4624 (N_4624,N_3690,N_2168);
and U4625 (N_4625,N_2066,N_3836);
nand U4626 (N_4626,N_3745,N_2376);
nand U4627 (N_4627,N_3355,N_2181);
and U4628 (N_4628,N_2849,N_3182);
nor U4629 (N_4629,N_2907,N_3686);
or U4630 (N_4630,N_3336,N_3938);
nor U4631 (N_4631,N_3263,N_2510);
or U4632 (N_4632,N_3583,N_3315);
nand U4633 (N_4633,N_2891,N_3054);
and U4634 (N_4634,N_3677,N_2123);
xnor U4635 (N_4635,N_3183,N_2143);
or U4636 (N_4636,N_3068,N_3916);
nand U4637 (N_4637,N_2591,N_2674);
nor U4638 (N_4638,N_3501,N_2291);
nand U4639 (N_4639,N_2115,N_2230);
xor U4640 (N_4640,N_3303,N_3748);
and U4641 (N_4641,N_2544,N_2498);
and U4642 (N_4642,N_3017,N_3397);
and U4643 (N_4643,N_3983,N_3436);
or U4644 (N_4644,N_2228,N_3240);
nand U4645 (N_4645,N_2358,N_3587);
or U4646 (N_4646,N_3667,N_3853);
or U4647 (N_4647,N_3651,N_2551);
xnor U4648 (N_4648,N_2262,N_2205);
or U4649 (N_4649,N_3100,N_3422);
and U4650 (N_4650,N_3590,N_3693);
nand U4651 (N_4651,N_3718,N_2908);
or U4652 (N_4652,N_2128,N_3483);
xnor U4653 (N_4653,N_3991,N_2259);
xnor U4654 (N_4654,N_3399,N_3930);
nor U4655 (N_4655,N_2208,N_2651);
and U4656 (N_4656,N_2341,N_3535);
nand U4657 (N_4657,N_2019,N_3308);
xnor U4658 (N_4658,N_2598,N_2871);
or U4659 (N_4659,N_3090,N_3753);
nand U4660 (N_4660,N_2236,N_2258);
nor U4661 (N_4661,N_2431,N_3691);
or U4662 (N_4662,N_2001,N_2251);
nand U4663 (N_4663,N_3708,N_2342);
nor U4664 (N_4664,N_2449,N_2192);
xor U4665 (N_4665,N_2424,N_2484);
nor U4666 (N_4666,N_2280,N_3601);
or U4667 (N_4667,N_2288,N_2906);
nor U4668 (N_4668,N_3235,N_3319);
nand U4669 (N_4669,N_2160,N_3174);
nand U4670 (N_4670,N_2072,N_3632);
xor U4671 (N_4671,N_3118,N_2061);
nor U4672 (N_4672,N_2531,N_3281);
nand U4673 (N_4673,N_3140,N_2344);
nor U4674 (N_4674,N_3984,N_2957);
nor U4675 (N_4675,N_3024,N_2277);
or U4676 (N_4676,N_3608,N_2172);
xnor U4677 (N_4677,N_3654,N_2943);
xnor U4678 (N_4678,N_3716,N_3815);
or U4679 (N_4679,N_2204,N_2026);
or U4680 (N_4680,N_2429,N_2805);
xor U4681 (N_4681,N_2333,N_3956);
nor U4682 (N_4682,N_3416,N_3818);
and U4683 (N_4683,N_3055,N_2404);
and U4684 (N_4684,N_2242,N_3218);
nand U4685 (N_4685,N_2546,N_2807);
or U4686 (N_4686,N_3098,N_2468);
or U4687 (N_4687,N_3335,N_2334);
xnor U4688 (N_4688,N_2127,N_2822);
xnor U4689 (N_4689,N_2357,N_2222);
and U4690 (N_4690,N_3634,N_2590);
xor U4691 (N_4691,N_3553,N_2993);
xnor U4692 (N_4692,N_2134,N_2229);
nor U4693 (N_4693,N_2629,N_3037);
xnor U4694 (N_4694,N_2558,N_3450);
nand U4695 (N_4695,N_2790,N_2995);
nor U4696 (N_4696,N_2751,N_3042);
and U4697 (N_4697,N_2834,N_3972);
and U4698 (N_4698,N_2869,N_2961);
or U4699 (N_4699,N_2453,N_2708);
nand U4700 (N_4700,N_3477,N_2518);
nand U4701 (N_4701,N_2503,N_3120);
and U4702 (N_4702,N_3089,N_3172);
or U4703 (N_4703,N_2900,N_3105);
nor U4704 (N_4704,N_3622,N_3301);
nor U4705 (N_4705,N_2492,N_3012);
nor U4706 (N_4706,N_2917,N_2073);
nor U4707 (N_4707,N_2013,N_2649);
and U4708 (N_4708,N_3659,N_2893);
nor U4709 (N_4709,N_3682,N_3765);
and U4710 (N_4710,N_2717,N_3884);
or U4711 (N_4711,N_3362,N_2811);
xor U4712 (N_4712,N_2655,N_2808);
xnor U4713 (N_4713,N_2008,N_3405);
and U4714 (N_4714,N_3375,N_3880);
nand U4715 (N_4715,N_2611,N_2640);
xor U4716 (N_4716,N_3584,N_3730);
and U4717 (N_4717,N_3573,N_3201);
and U4718 (N_4718,N_2087,N_3200);
and U4719 (N_4719,N_2956,N_3007);
and U4720 (N_4720,N_3383,N_3465);
and U4721 (N_4721,N_3625,N_2635);
nand U4722 (N_4722,N_2614,N_3428);
nor U4723 (N_4723,N_2622,N_3555);
or U4724 (N_4724,N_2380,N_2028);
xnor U4725 (N_4725,N_2522,N_3171);
xor U4726 (N_4726,N_3908,N_2605);
nor U4727 (N_4727,N_2326,N_2860);
xor U4728 (N_4728,N_3921,N_3812);
xnor U4729 (N_4729,N_2984,N_2051);
or U4730 (N_4730,N_3549,N_2744);
xnor U4731 (N_4731,N_3210,N_3152);
xnor U4732 (N_4732,N_2451,N_3203);
xnor U4733 (N_4733,N_3198,N_3883);
nor U4734 (N_4734,N_2117,N_2972);
nand U4735 (N_4735,N_3027,N_3964);
xor U4736 (N_4736,N_3237,N_3165);
nand U4737 (N_4737,N_3398,N_3532);
and U4738 (N_4738,N_2257,N_3199);
or U4739 (N_4739,N_3868,N_3178);
nand U4740 (N_4740,N_3830,N_2485);
xnor U4741 (N_4741,N_2699,N_2641);
nand U4742 (N_4742,N_3829,N_2331);
and U4743 (N_4743,N_3425,N_2678);
xor U4744 (N_4744,N_3334,N_3561);
and U4745 (N_4745,N_2713,N_3015);
xnor U4746 (N_4746,N_3113,N_3657);
xor U4747 (N_4747,N_3051,N_3391);
nand U4748 (N_4748,N_2471,N_2767);
nand U4749 (N_4749,N_3768,N_2896);
nor U4750 (N_4750,N_3379,N_3678);
nand U4751 (N_4751,N_3305,N_2743);
and U4752 (N_4752,N_3998,N_3534);
and U4753 (N_4753,N_2462,N_3291);
and U4754 (N_4754,N_2862,N_3052);
nand U4755 (N_4755,N_2477,N_3500);
nand U4756 (N_4756,N_3195,N_2578);
and U4757 (N_4757,N_2707,N_2505);
nand U4758 (N_4758,N_2034,N_3498);
or U4759 (N_4759,N_2934,N_2179);
nand U4760 (N_4760,N_3248,N_3496);
and U4761 (N_4761,N_3280,N_2987);
nand U4762 (N_4762,N_2610,N_3844);
nor U4763 (N_4763,N_2027,N_3163);
and U4764 (N_4764,N_2883,N_3346);
or U4765 (N_4765,N_2576,N_3344);
nand U4766 (N_4766,N_2489,N_3887);
nand U4767 (N_4767,N_2946,N_2977);
nor U4768 (N_4768,N_2647,N_2842);
nor U4769 (N_4769,N_2865,N_3629);
or U4770 (N_4770,N_2725,N_2460);
and U4771 (N_4771,N_3309,N_3602);
nor U4772 (N_4772,N_3401,N_3859);
nor U4773 (N_4773,N_2988,N_2646);
nand U4774 (N_4774,N_2731,N_3451);
and U4775 (N_4775,N_2031,N_2574);
or U4776 (N_4776,N_3788,N_2763);
nand U4777 (N_4777,N_3390,N_2600);
nand U4778 (N_4778,N_3204,N_3735);
and U4779 (N_4779,N_2511,N_2042);
nand U4780 (N_4780,N_3842,N_3644);
nor U4781 (N_4781,N_3696,N_2191);
nand U4782 (N_4782,N_3508,N_2671);
nor U4783 (N_4783,N_2487,N_3350);
xor U4784 (N_4784,N_3697,N_2408);
nand U4785 (N_4785,N_3026,N_2083);
xnor U4786 (N_4786,N_2887,N_3924);
xor U4787 (N_4787,N_3992,N_3503);
and U4788 (N_4788,N_3910,N_2567);
nor U4789 (N_4789,N_2954,N_2202);
or U4790 (N_4790,N_2854,N_3655);
or U4791 (N_4791,N_2922,N_2101);
or U4792 (N_4792,N_2354,N_3932);
nor U4793 (N_4793,N_2696,N_2243);
nand U4794 (N_4794,N_2895,N_3126);
nor U4795 (N_4795,N_2978,N_3683);
nor U4796 (N_4796,N_3628,N_3847);
nor U4797 (N_4797,N_2617,N_3499);
nor U4798 (N_4798,N_3828,N_3536);
nand U4799 (N_4799,N_3945,N_2566);
nand U4800 (N_4800,N_2410,N_2402);
nor U4801 (N_4801,N_2873,N_3736);
nor U4802 (N_4802,N_3025,N_3087);
or U4803 (N_4803,N_3386,N_2017);
and U4804 (N_4804,N_2307,N_2273);
and U4805 (N_4805,N_3413,N_2968);
nand U4806 (N_4806,N_3253,N_2398);
nand U4807 (N_4807,N_2033,N_2851);
and U4808 (N_4808,N_3370,N_3597);
or U4809 (N_4809,N_2458,N_2925);
nand U4810 (N_4810,N_2153,N_2491);
xnor U4811 (N_4811,N_3456,N_2296);
or U4812 (N_4812,N_2726,N_3168);
and U4813 (N_4813,N_2478,N_3951);
or U4814 (N_4814,N_3359,N_3873);
xor U4815 (N_4815,N_2684,N_2527);
xor U4816 (N_4816,N_3307,N_2272);
or U4817 (N_4817,N_2256,N_2573);
and U4818 (N_4818,N_2831,N_2732);
xor U4819 (N_4819,N_2141,N_2630);
xnor U4820 (N_4820,N_3893,N_2927);
or U4821 (N_4821,N_3115,N_3767);
xnor U4822 (N_4822,N_2739,N_3756);
or U4823 (N_4823,N_3187,N_3710);
and U4824 (N_4824,N_3338,N_2226);
and U4825 (N_4825,N_3420,N_3154);
or U4826 (N_4826,N_3266,N_3521);
nand U4827 (N_4827,N_3481,N_2469);
or U4828 (N_4828,N_3135,N_3354);
xor U4829 (N_4829,N_3546,N_2772);
nor U4830 (N_4830,N_2559,N_2095);
or U4831 (N_4831,N_2488,N_3719);
and U4832 (N_4832,N_2963,N_2940);
nor U4833 (N_4833,N_3727,N_3515);
nand U4834 (N_4834,N_2150,N_3662);
and U4835 (N_4835,N_3217,N_2053);
nand U4836 (N_4836,N_2798,N_3826);
nand U4837 (N_4837,N_3542,N_3700);
nand U4838 (N_4838,N_2495,N_3189);
and U4839 (N_4839,N_2400,N_2133);
and U4840 (N_4840,N_3947,N_2340);
and U4841 (N_4841,N_2418,N_2109);
nand U4842 (N_4842,N_3264,N_2048);
xor U4843 (N_4843,N_3525,N_3547);
or U4844 (N_4844,N_3445,N_3221);
nand U4845 (N_4845,N_2680,N_3666);
xnor U4846 (N_4846,N_3212,N_3190);
xnor U4847 (N_4847,N_2216,N_2668);
xor U4848 (N_4848,N_2827,N_2818);
nor U4849 (N_4849,N_2411,N_3078);
nand U4850 (N_4850,N_2889,N_3605);
nor U4851 (N_4851,N_3850,N_2914);
nor U4852 (N_4852,N_3232,N_3530);
nor U4853 (N_4853,N_3740,N_3518);
nor U4854 (N_4854,N_3869,N_2540);
or U4855 (N_4855,N_3018,N_2676);
nand U4856 (N_4856,N_3808,N_2170);
or U4857 (N_4857,N_2745,N_3358);
nor U4858 (N_4858,N_2543,N_2694);
or U4859 (N_4859,N_3714,N_3225);
or U4860 (N_4860,N_3941,N_3856);
nor U4861 (N_4861,N_2983,N_2915);
xor U4862 (N_4862,N_3382,N_3242);
and U4863 (N_4863,N_3197,N_2550);
or U4864 (N_4864,N_2654,N_3717);
nand U4865 (N_4865,N_3653,N_2901);
nand U4866 (N_4866,N_2235,N_2936);
nor U4867 (N_4867,N_3339,N_3764);
or U4868 (N_4868,N_2011,N_2038);
and U4869 (N_4869,N_2750,N_2180);
and U4870 (N_4870,N_3348,N_2009);
xnor U4871 (N_4871,N_3014,N_2890);
or U4872 (N_4872,N_2392,N_3031);
xor U4873 (N_4873,N_3776,N_3003);
nand U4874 (N_4874,N_2624,N_2003);
nand U4875 (N_4875,N_3732,N_2773);
xnor U4876 (N_4876,N_3104,N_2833);
nand U4877 (N_4877,N_3840,N_2626);
nor U4878 (N_4878,N_3365,N_2557);
or U4879 (N_4879,N_3982,N_3323);
or U4880 (N_4880,N_2562,N_2328);
nor U4881 (N_4881,N_3371,N_2159);
and U4882 (N_4882,N_2682,N_2071);
nor U4883 (N_4883,N_2514,N_3332);
nor U4884 (N_4884,N_2803,N_3554);
nand U4885 (N_4885,N_3156,N_3347);
and U4886 (N_4886,N_2343,N_3132);
xnor U4887 (N_4887,N_2506,N_2303);
or U4888 (N_4888,N_3298,N_2241);
or U4889 (N_4889,N_2417,N_3675);
and U4890 (N_4890,N_3664,N_2933);
xor U4891 (N_4891,N_2324,N_2074);
xor U4892 (N_4892,N_2046,N_2881);
and U4893 (N_4893,N_3129,N_3725);
and U4894 (N_4894,N_3145,N_2015);
nor U4895 (N_4895,N_3310,N_2088);
xnor U4896 (N_4896,N_2613,N_3790);
and U4897 (N_4897,N_3293,N_2438);
or U4898 (N_4898,N_2935,N_3761);
and U4899 (N_4899,N_3504,N_3799);
xor U4900 (N_4900,N_2443,N_2841);
and U4901 (N_4901,N_3572,N_3080);
xnor U4902 (N_4902,N_2442,N_2390);
nand U4903 (N_4903,N_2904,N_3997);
nand U4904 (N_4904,N_3356,N_2107);
nor U4905 (N_4905,N_3698,N_3743);
or U4906 (N_4906,N_2608,N_3473);
nor U4907 (N_4907,N_2174,N_3520);
xnor U4908 (N_4908,N_2658,N_2718);
nand U4909 (N_4909,N_3284,N_3117);
nand U4910 (N_4910,N_2856,N_2098);
xnor U4911 (N_4911,N_3415,N_2692);
nand U4912 (N_4912,N_2950,N_2434);
nor U4913 (N_4913,N_3418,N_3227);
and U4914 (N_4914,N_3560,N_2774);
nand U4915 (N_4915,N_3639,N_3458);
or U4916 (N_4916,N_2450,N_3121);
nand U4917 (N_4917,N_3593,N_3328);
and U4918 (N_4918,N_2165,N_3053);
and U4919 (N_4919,N_2962,N_2004);
nor U4920 (N_4920,N_2100,N_3389);
nand U4921 (N_4921,N_2412,N_2815);
nand U4922 (N_4922,N_2130,N_3394);
nor U4923 (N_4923,N_2835,N_2021);
nor U4924 (N_4924,N_3330,N_3950);
nor U4925 (N_4925,N_2085,N_2407);
xnor U4926 (N_4926,N_2169,N_3647);
nor U4927 (N_4927,N_2177,N_3180);
nor U4928 (N_4928,N_2363,N_3955);
xnor U4929 (N_4929,N_3552,N_3707);
nor U4930 (N_4930,N_3047,N_2014);
xor U4931 (N_4931,N_2724,N_2387);
and U4932 (N_4932,N_2152,N_2670);
or U4933 (N_4933,N_3077,N_3729);
xnor U4934 (N_4934,N_3331,N_3866);
nand U4935 (N_4935,N_3069,N_2310);
nor U4936 (N_4936,N_2796,N_2311);
and U4937 (N_4937,N_2182,N_3544);
nand U4938 (N_4938,N_3604,N_3085);
xnor U4939 (N_4939,N_2024,N_2044);
or U4940 (N_4940,N_3108,N_2783);
and U4941 (N_4941,N_2427,N_3381);
nand U4942 (N_4942,N_3088,N_2679);
nand U4943 (N_4943,N_2967,N_2932);
nand U4944 (N_4944,N_3364,N_3103);
or U4945 (N_4945,N_3961,N_3851);
nor U4946 (N_4946,N_2129,N_2140);
or U4947 (N_4947,N_2171,N_3734);
or U4948 (N_4948,N_2580,N_3122);
nand U4949 (N_4949,N_3989,N_2108);
nand U4950 (N_4950,N_3461,N_3755);
nand U4951 (N_4951,N_2052,N_3048);
or U4952 (N_4952,N_3403,N_3976);
nor U4953 (N_4953,N_2770,N_2060);
xor U4954 (N_4954,N_3245,N_3191);
xor U4955 (N_4955,N_2233,N_2030);
or U4956 (N_4956,N_3074,N_3923);
xnor U4957 (N_4957,N_2715,N_3095);
and U4958 (N_4958,N_3876,N_3879);
nor U4959 (N_4959,N_3617,N_2810);
and U4960 (N_4960,N_2826,N_3848);
xnor U4961 (N_4961,N_3979,N_2113);
nand U4962 (N_4962,N_3408,N_2660);
nor U4963 (N_4963,N_3423,N_3326);
nand U4964 (N_4964,N_2237,N_2375);
or U4965 (N_4965,N_2882,N_2317);
xnor U4966 (N_4966,N_2911,N_2290);
and U4967 (N_4967,N_2312,N_3801);
or U4968 (N_4968,N_2183,N_3123);
or U4969 (N_4969,N_3101,N_3125);
nand U4970 (N_4970,N_2120,N_2432);
and U4971 (N_4971,N_3962,N_2571);
nand U4972 (N_4972,N_2261,N_2697);
or U4973 (N_4973,N_2560,N_2353);
or U4974 (N_4974,N_3241,N_3823);
xnor U4975 (N_4975,N_3226,N_3720);
xor U4976 (N_4976,N_3111,N_2866);
and U4977 (N_4977,N_3366,N_3474);
xnor U4978 (N_4978,N_2355,N_2997);
nor U4979 (N_4979,N_2565,N_2252);
xor U4980 (N_4980,N_2436,N_2857);
nor U4981 (N_4981,N_3459,N_3429);
or U4982 (N_4982,N_2486,N_2286);
nand U4983 (N_4983,N_2879,N_2870);
nand U4984 (N_4984,N_3469,N_3058);
xor U4985 (N_4985,N_2627,N_3139);
xor U4986 (N_4986,N_2919,N_2853);
xnor U4987 (N_4987,N_2330,N_2710);
nor U4988 (N_4988,N_3324,N_3971);
nand U4989 (N_4989,N_3526,N_2784);
and U4990 (N_4990,N_3169,N_3817);
and U4991 (N_4991,N_3656,N_2185);
nor U4992 (N_4992,N_3596,N_3918);
xor U4993 (N_4993,N_3395,N_3274);
nand U4994 (N_4994,N_3124,N_3050);
nand U4995 (N_4995,N_3671,N_2852);
and U4996 (N_4996,N_3194,N_3485);
or U4997 (N_4997,N_3230,N_3612);
xor U4998 (N_4998,N_3153,N_2059);
and U4999 (N_4999,N_3839,N_2224);
nor U5000 (N_5000,N_3445,N_2533);
or U5001 (N_5001,N_2264,N_3188);
xor U5002 (N_5002,N_2880,N_2599);
and U5003 (N_5003,N_3048,N_3611);
nor U5004 (N_5004,N_2412,N_2506);
nand U5005 (N_5005,N_3468,N_3158);
or U5006 (N_5006,N_3358,N_3058);
and U5007 (N_5007,N_3733,N_3842);
and U5008 (N_5008,N_3578,N_3085);
nand U5009 (N_5009,N_3799,N_3278);
or U5010 (N_5010,N_3564,N_2192);
and U5011 (N_5011,N_2226,N_3597);
nand U5012 (N_5012,N_3491,N_3951);
xor U5013 (N_5013,N_2339,N_2730);
or U5014 (N_5014,N_2057,N_2505);
xnor U5015 (N_5015,N_3790,N_2944);
nor U5016 (N_5016,N_3348,N_2867);
xnor U5017 (N_5017,N_3059,N_3236);
or U5018 (N_5018,N_2874,N_3398);
and U5019 (N_5019,N_3209,N_3147);
and U5020 (N_5020,N_3168,N_3764);
xor U5021 (N_5021,N_2567,N_2586);
xor U5022 (N_5022,N_3145,N_3213);
and U5023 (N_5023,N_2796,N_3801);
nor U5024 (N_5024,N_2947,N_3051);
nand U5025 (N_5025,N_2806,N_2923);
nor U5026 (N_5026,N_2323,N_2947);
nand U5027 (N_5027,N_3297,N_2413);
nor U5028 (N_5028,N_3214,N_3021);
and U5029 (N_5029,N_3831,N_2353);
nor U5030 (N_5030,N_2219,N_3436);
and U5031 (N_5031,N_2194,N_3002);
or U5032 (N_5032,N_3907,N_3230);
nand U5033 (N_5033,N_2661,N_2414);
nand U5034 (N_5034,N_2713,N_2922);
nor U5035 (N_5035,N_2405,N_2786);
and U5036 (N_5036,N_2236,N_2463);
nor U5037 (N_5037,N_3797,N_2336);
or U5038 (N_5038,N_3433,N_2458);
nor U5039 (N_5039,N_2623,N_2424);
or U5040 (N_5040,N_3165,N_2268);
xnor U5041 (N_5041,N_3275,N_3521);
or U5042 (N_5042,N_3701,N_3938);
and U5043 (N_5043,N_2656,N_3435);
xnor U5044 (N_5044,N_3057,N_3833);
xor U5045 (N_5045,N_2513,N_3332);
or U5046 (N_5046,N_2535,N_3759);
xnor U5047 (N_5047,N_3790,N_2653);
and U5048 (N_5048,N_2573,N_2509);
nand U5049 (N_5049,N_3770,N_2094);
and U5050 (N_5050,N_3541,N_3918);
or U5051 (N_5051,N_2242,N_3096);
xor U5052 (N_5052,N_3610,N_2709);
nand U5053 (N_5053,N_3817,N_2976);
and U5054 (N_5054,N_3478,N_3354);
or U5055 (N_5055,N_3487,N_2235);
nand U5056 (N_5056,N_2035,N_3926);
xnor U5057 (N_5057,N_2475,N_3059);
nor U5058 (N_5058,N_2848,N_3025);
or U5059 (N_5059,N_2129,N_2436);
nor U5060 (N_5060,N_3950,N_2280);
xnor U5061 (N_5061,N_2251,N_3836);
nor U5062 (N_5062,N_2695,N_2458);
and U5063 (N_5063,N_2697,N_2307);
xnor U5064 (N_5064,N_2119,N_3007);
xor U5065 (N_5065,N_3667,N_3207);
and U5066 (N_5066,N_2189,N_2428);
xor U5067 (N_5067,N_2309,N_3721);
nor U5068 (N_5068,N_2621,N_2497);
or U5069 (N_5069,N_3906,N_3654);
and U5070 (N_5070,N_2812,N_2963);
and U5071 (N_5071,N_3587,N_3749);
nand U5072 (N_5072,N_3895,N_3038);
and U5073 (N_5073,N_3098,N_2503);
or U5074 (N_5074,N_3715,N_2727);
xor U5075 (N_5075,N_2546,N_3939);
xor U5076 (N_5076,N_2816,N_3613);
nand U5077 (N_5077,N_3371,N_3723);
nand U5078 (N_5078,N_3764,N_2465);
nand U5079 (N_5079,N_2158,N_3797);
or U5080 (N_5080,N_3938,N_3637);
nor U5081 (N_5081,N_3993,N_2777);
and U5082 (N_5082,N_2794,N_2759);
or U5083 (N_5083,N_2587,N_2433);
nor U5084 (N_5084,N_3259,N_2352);
xor U5085 (N_5085,N_2368,N_2425);
nor U5086 (N_5086,N_3315,N_2224);
nand U5087 (N_5087,N_2702,N_3812);
nor U5088 (N_5088,N_3571,N_3965);
and U5089 (N_5089,N_2481,N_3424);
or U5090 (N_5090,N_3168,N_3306);
nand U5091 (N_5091,N_3276,N_3704);
and U5092 (N_5092,N_3999,N_3487);
nor U5093 (N_5093,N_3454,N_2228);
and U5094 (N_5094,N_2825,N_3410);
or U5095 (N_5095,N_3905,N_2711);
xor U5096 (N_5096,N_2899,N_2730);
xor U5097 (N_5097,N_3726,N_3593);
and U5098 (N_5098,N_3962,N_3385);
nor U5099 (N_5099,N_3053,N_3433);
or U5100 (N_5100,N_3164,N_3264);
xnor U5101 (N_5101,N_3067,N_2830);
xnor U5102 (N_5102,N_3020,N_3149);
nand U5103 (N_5103,N_3834,N_3915);
and U5104 (N_5104,N_3461,N_2805);
nand U5105 (N_5105,N_3307,N_3857);
or U5106 (N_5106,N_2292,N_3401);
or U5107 (N_5107,N_2535,N_2377);
or U5108 (N_5108,N_2667,N_2351);
nand U5109 (N_5109,N_2196,N_2261);
nor U5110 (N_5110,N_3514,N_2770);
and U5111 (N_5111,N_3880,N_2651);
and U5112 (N_5112,N_2723,N_3542);
or U5113 (N_5113,N_3229,N_2633);
nor U5114 (N_5114,N_2537,N_3250);
nand U5115 (N_5115,N_2110,N_3510);
xor U5116 (N_5116,N_3983,N_3253);
nor U5117 (N_5117,N_3343,N_2372);
or U5118 (N_5118,N_3486,N_3326);
nor U5119 (N_5119,N_2273,N_2030);
nor U5120 (N_5120,N_2052,N_2038);
nand U5121 (N_5121,N_3662,N_3900);
xor U5122 (N_5122,N_3848,N_2774);
xnor U5123 (N_5123,N_3178,N_3596);
xor U5124 (N_5124,N_3445,N_2591);
nor U5125 (N_5125,N_2225,N_3017);
or U5126 (N_5126,N_3503,N_3829);
nand U5127 (N_5127,N_2394,N_3888);
nand U5128 (N_5128,N_3844,N_2348);
or U5129 (N_5129,N_3583,N_2023);
nand U5130 (N_5130,N_3706,N_2923);
and U5131 (N_5131,N_2311,N_2394);
xor U5132 (N_5132,N_3954,N_3038);
nor U5133 (N_5133,N_2977,N_3763);
and U5134 (N_5134,N_2748,N_3755);
and U5135 (N_5135,N_3931,N_3642);
or U5136 (N_5136,N_2214,N_2307);
nor U5137 (N_5137,N_2008,N_2025);
xor U5138 (N_5138,N_2637,N_2289);
xor U5139 (N_5139,N_3961,N_3285);
and U5140 (N_5140,N_3263,N_3543);
and U5141 (N_5141,N_3697,N_3344);
nand U5142 (N_5142,N_3686,N_2784);
nand U5143 (N_5143,N_3123,N_3640);
and U5144 (N_5144,N_2796,N_2165);
or U5145 (N_5145,N_2990,N_3701);
nor U5146 (N_5146,N_2851,N_3526);
and U5147 (N_5147,N_2229,N_3361);
xor U5148 (N_5148,N_2814,N_2513);
nor U5149 (N_5149,N_2074,N_2164);
nor U5150 (N_5150,N_3402,N_3773);
nor U5151 (N_5151,N_2588,N_3734);
xnor U5152 (N_5152,N_3388,N_2862);
and U5153 (N_5153,N_2336,N_3102);
and U5154 (N_5154,N_2691,N_2880);
or U5155 (N_5155,N_3348,N_2000);
or U5156 (N_5156,N_3278,N_3029);
xor U5157 (N_5157,N_2202,N_3829);
nand U5158 (N_5158,N_2762,N_3536);
or U5159 (N_5159,N_2723,N_2378);
and U5160 (N_5160,N_2321,N_2450);
xor U5161 (N_5161,N_2299,N_2453);
nand U5162 (N_5162,N_2833,N_3135);
or U5163 (N_5163,N_2515,N_2838);
nand U5164 (N_5164,N_3625,N_2855);
xnor U5165 (N_5165,N_3017,N_2777);
nor U5166 (N_5166,N_3641,N_2777);
nor U5167 (N_5167,N_3691,N_3422);
and U5168 (N_5168,N_3676,N_2506);
xnor U5169 (N_5169,N_3495,N_2730);
xor U5170 (N_5170,N_2559,N_2312);
and U5171 (N_5171,N_3198,N_3082);
or U5172 (N_5172,N_3644,N_3924);
nor U5173 (N_5173,N_2870,N_3243);
or U5174 (N_5174,N_3656,N_3429);
and U5175 (N_5175,N_3446,N_3635);
xor U5176 (N_5176,N_2431,N_3730);
xnor U5177 (N_5177,N_2706,N_2417);
or U5178 (N_5178,N_3516,N_2287);
xnor U5179 (N_5179,N_2247,N_3990);
nand U5180 (N_5180,N_3486,N_2736);
or U5181 (N_5181,N_3190,N_2905);
nor U5182 (N_5182,N_3160,N_2912);
and U5183 (N_5183,N_2063,N_3943);
nor U5184 (N_5184,N_3001,N_3101);
or U5185 (N_5185,N_3439,N_2795);
or U5186 (N_5186,N_2889,N_3002);
nand U5187 (N_5187,N_2114,N_2232);
nor U5188 (N_5188,N_2164,N_3694);
nor U5189 (N_5189,N_3387,N_2805);
nand U5190 (N_5190,N_2779,N_3402);
xor U5191 (N_5191,N_3555,N_2422);
nor U5192 (N_5192,N_2796,N_3727);
nand U5193 (N_5193,N_3779,N_3169);
nor U5194 (N_5194,N_3527,N_3158);
or U5195 (N_5195,N_3358,N_2118);
nand U5196 (N_5196,N_3725,N_3673);
or U5197 (N_5197,N_2526,N_2158);
nor U5198 (N_5198,N_3511,N_3911);
and U5199 (N_5199,N_2480,N_3072);
nand U5200 (N_5200,N_2562,N_2379);
nor U5201 (N_5201,N_3271,N_2263);
nor U5202 (N_5202,N_2200,N_2128);
or U5203 (N_5203,N_3758,N_3143);
or U5204 (N_5204,N_3784,N_2158);
nor U5205 (N_5205,N_3223,N_2477);
nor U5206 (N_5206,N_3391,N_2107);
and U5207 (N_5207,N_2150,N_2891);
nand U5208 (N_5208,N_3802,N_2837);
and U5209 (N_5209,N_3067,N_3813);
xor U5210 (N_5210,N_3981,N_3236);
nor U5211 (N_5211,N_2103,N_2980);
nor U5212 (N_5212,N_2451,N_2636);
nand U5213 (N_5213,N_2204,N_2160);
nand U5214 (N_5214,N_3933,N_2843);
xor U5215 (N_5215,N_3757,N_3922);
or U5216 (N_5216,N_3463,N_2387);
nor U5217 (N_5217,N_2840,N_2472);
or U5218 (N_5218,N_3884,N_2321);
xnor U5219 (N_5219,N_3493,N_3611);
nand U5220 (N_5220,N_3150,N_2064);
or U5221 (N_5221,N_3221,N_3744);
or U5222 (N_5222,N_3254,N_3255);
or U5223 (N_5223,N_3789,N_2487);
and U5224 (N_5224,N_2484,N_3806);
nor U5225 (N_5225,N_3388,N_3501);
and U5226 (N_5226,N_2391,N_3179);
nor U5227 (N_5227,N_2643,N_3458);
xnor U5228 (N_5228,N_3681,N_3623);
or U5229 (N_5229,N_3159,N_3595);
nand U5230 (N_5230,N_2465,N_3086);
xnor U5231 (N_5231,N_3819,N_2120);
and U5232 (N_5232,N_3010,N_3880);
and U5233 (N_5233,N_3416,N_3248);
or U5234 (N_5234,N_2383,N_3299);
nor U5235 (N_5235,N_3228,N_3171);
nor U5236 (N_5236,N_3773,N_3478);
xnor U5237 (N_5237,N_3934,N_2370);
or U5238 (N_5238,N_3283,N_3074);
nand U5239 (N_5239,N_3694,N_2827);
or U5240 (N_5240,N_3921,N_2682);
xor U5241 (N_5241,N_3448,N_2643);
and U5242 (N_5242,N_3560,N_3822);
xor U5243 (N_5243,N_3947,N_2366);
nand U5244 (N_5244,N_3245,N_2847);
nand U5245 (N_5245,N_3706,N_2169);
and U5246 (N_5246,N_3431,N_3861);
nand U5247 (N_5247,N_2917,N_3918);
nor U5248 (N_5248,N_3676,N_3120);
or U5249 (N_5249,N_3168,N_3193);
nand U5250 (N_5250,N_2272,N_2039);
xor U5251 (N_5251,N_3115,N_3277);
xor U5252 (N_5252,N_2230,N_2215);
nand U5253 (N_5253,N_3677,N_2349);
or U5254 (N_5254,N_3637,N_3331);
xor U5255 (N_5255,N_3181,N_2899);
and U5256 (N_5256,N_2698,N_3319);
xor U5257 (N_5257,N_2035,N_2824);
nor U5258 (N_5258,N_3739,N_2105);
or U5259 (N_5259,N_2203,N_3679);
or U5260 (N_5260,N_2111,N_2406);
xnor U5261 (N_5261,N_3705,N_2464);
nor U5262 (N_5262,N_2003,N_2499);
or U5263 (N_5263,N_2388,N_2768);
xnor U5264 (N_5264,N_2404,N_2923);
nor U5265 (N_5265,N_3332,N_2479);
xor U5266 (N_5266,N_3109,N_2028);
nor U5267 (N_5267,N_2102,N_3156);
and U5268 (N_5268,N_3908,N_2935);
xor U5269 (N_5269,N_2806,N_3832);
xor U5270 (N_5270,N_3440,N_2074);
xor U5271 (N_5271,N_3857,N_2629);
xor U5272 (N_5272,N_3065,N_3485);
nor U5273 (N_5273,N_3631,N_3512);
or U5274 (N_5274,N_2819,N_3009);
nand U5275 (N_5275,N_2053,N_3315);
xor U5276 (N_5276,N_3208,N_3689);
nand U5277 (N_5277,N_2179,N_2553);
nor U5278 (N_5278,N_2285,N_3864);
or U5279 (N_5279,N_2849,N_2890);
or U5280 (N_5280,N_3732,N_3979);
nand U5281 (N_5281,N_2663,N_2555);
nor U5282 (N_5282,N_2330,N_3303);
nand U5283 (N_5283,N_3339,N_3577);
nor U5284 (N_5284,N_2757,N_2824);
nand U5285 (N_5285,N_2709,N_3669);
nor U5286 (N_5286,N_2165,N_3856);
xnor U5287 (N_5287,N_2505,N_2616);
nor U5288 (N_5288,N_3873,N_3618);
and U5289 (N_5289,N_2157,N_2687);
nor U5290 (N_5290,N_2011,N_3294);
or U5291 (N_5291,N_2445,N_3029);
xor U5292 (N_5292,N_2386,N_3910);
nor U5293 (N_5293,N_2124,N_2852);
or U5294 (N_5294,N_3540,N_3294);
or U5295 (N_5295,N_2653,N_2629);
xor U5296 (N_5296,N_3854,N_2370);
xor U5297 (N_5297,N_2515,N_2728);
nor U5298 (N_5298,N_2147,N_3499);
and U5299 (N_5299,N_3785,N_2320);
xor U5300 (N_5300,N_2764,N_2589);
xnor U5301 (N_5301,N_3803,N_3345);
xor U5302 (N_5302,N_3369,N_3795);
nand U5303 (N_5303,N_3232,N_2935);
nor U5304 (N_5304,N_2293,N_2412);
and U5305 (N_5305,N_2644,N_3199);
or U5306 (N_5306,N_2440,N_2517);
and U5307 (N_5307,N_2915,N_2485);
and U5308 (N_5308,N_2050,N_3377);
and U5309 (N_5309,N_3266,N_3162);
xnor U5310 (N_5310,N_2766,N_3144);
xnor U5311 (N_5311,N_3785,N_3793);
or U5312 (N_5312,N_3742,N_2265);
or U5313 (N_5313,N_2300,N_3366);
and U5314 (N_5314,N_3692,N_2235);
nand U5315 (N_5315,N_2089,N_2718);
nor U5316 (N_5316,N_3603,N_3905);
or U5317 (N_5317,N_2496,N_2888);
nand U5318 (N_5318,N_3343,N_3685);
nand U5319 (N_5319,N_2002,N_2505);
nor U5320 (N_5320,N_2296,N_2471);
nor U5321 (N_5321,N_2856,N_2342);
xnor U5322 (N_5322,N_3989,N_3374);
xnor U5323 (N_5323,N_3260,N_2775);
nand U5324 (N_5324,N_2957,N_3901);
and U5325 (N_5325,N_2333,N_3341);
and U5326 (N_5326,N_3134,N_3670);
nand U5327 (N_5327,N_2589,N_2207);
or U5328 (N_5328,N_2168,N_3167);
and U5329 (N_5329,N_2810,N_2657);
nor U5330 (N_5330,N_3360,N_3154);
or U5331 (N_5331,N_2432,N_3490);
nor U5332 (N_5332,N_2334,N_2073);
nor U5333 (N_5333,N_2526,N_3070);
and U5334 (N_5334,N_3022,N_2311);
nand U5335 (N_5335,N_3547,N_2448);
and U5336 (N_5336,N_2632,N_3607);
or U5337 (N_5337,N_2384,N_3491);
or U5338 (N_5338,N_2206,N_3410);
or U5339 (N_5339,N_3182,N_3639);
and U5340 (N_5340,N_3121,N_3760);
or U5341 (N_5341,N_3453,N_2279);
nand U5342 (N_5342,N_3305,N_3299);
nor U5343 (N_5343,N_3877,N_2176);
nand U5344 (N_5344,N_3831,N_2547);
xor U5345 (N_5345,N_3686,N_3412);
and U5346 (N_5346,N_2933,N_2219);
and U5347 (N_5347,N_3088,N_3573);
and U5348 (N_5348,N_3504,N_3836);
xnor U5349 (N_5349,N_2430,N_2706);
xor U5350 (N_5350,N_2867,N_3517);
xor U5351 (N_5351,N_2855,N_2725);
and U5352 (N_5352,N_3996,N_2130);
or U5353 (N_5353,N_3588,N_2870);
nor U5354 (N_5354,N_2471,N_3059);
or U5355 (N_5355,N_3633,N_3602);
nor U5356 (N_5356,N_2176,N_3407);
nand U5357 (N_5357,N_3790,N_2108);
or U5358 (N_5358,N_3389,N_3544);
nand U5359 (N_5359,N_2103,N_2578);
or U5360 (N_5360,N_2595,N_3806);
xor U5361 (N_5361,N_3946,N_3858);
and U5362 (N_5362,N_3776,N_3320);
and U5363 (N_5363,N_3028,N_2771);
nor U5364 (N_5364,N_2273,N_3606);
nand U5365 (N_5365,N_2595,N_2730);
nand U5366 (N_5366,N_2327,N_2441);
or U5367 (N_5367,N_3703,N_2289);
or U5368 (N_5368,N_3662,N_3597);
and U5369 (N_5369,N_3006,N_3929);
nor U5370 (N_5370,N_2491,N_2781);
and U5371 (N_5371,N_3805,N_3225);
nor U5372 (N_5372,N_3027,N_3901);
nor U5373 (N_5373,N_2069,N_2490);
nand U5374 (N_5374,N_3558,N_3994);
or U5375 (N_5375,N_3462,N_3976);
and U5376 (N_5376,N_3076,N_3860);
xnor U5377 (N_5377,N_2362,N_3174);
nor U5378 (N_5378,N_3835,N_2152);
nor U5379 (N_5379,N_2158,N_2947);
nor U5380 (N_5380,N_3811,N_3204);
and U5381 (N_5381,N_2776,N_3562);
and U5382 (N_5382,N_3384,N_3248);
and U5383 (N_5383,N_3619,N_3982);
xnor U5384 (N_5384,N_2319,N_2830);
and U5385 (N_5385,N_3765,N_3159);
or U5386 (N_5386,N_2601,N_3976);
nand U5387 (N_5387,N_3862,N_2555);
and U5388 (N_5388,N_2171,N_2848);
or U5389 (N_5389,N_2412,N_3360);
and U5390 (N_5390,N_2793,N_2157);
xnor U5391 (N_5391,N_3060,N_3102);
or U5392 (N_5392,N_3263,N_3342);
nor U5393 (N_5393,N_3860,N_2111);
xnor U5394 (N_5394,N_3786,N_2028);
and U5395 (N_5395,N_3371,N_3740);
or U5396 (N_5396,N_2476,N_2828);
nor U5397 (N_5397,N_2617,N_3991);
nand U5398 (N_5398,N_3502,N_2851);
and U5399 (N_5399,N_3237,N_2011);
nor U5400 (N_5400,N_2646,N_2284);
and U5401 (N_5401,N_3766,N_2677);
nor U5402 (N_5402,N_2955,N_3203);
xnor U5403 (N_5403,N_3702,N_2156);
or U5404 (N_5404,N_3157,N_3777);
nor U5405 (N_5405,N_3345,N_2168);
nor U5406 (N_5406,N_3198,N_2744);
xnor U5407 (N_5407,N_3076,N_3968);
nand U5408 (N_5408,N_3098,N_2130);
xor U5409 (N_5409,N_2059,N_2727);
and U5410 (N_5410,N_2625,N_2030);
xnor U5411 (N_5411,N_3949,N_3544);
nor U5412 (N_5412,N_3865,N_2186);
nand U5413 (N_5413,N_2199,N_2761);
nor U5414 (N_5414,N_3559,N_3617);
and U5415 (N_5415,N_3422,N_2085);
nand U5416 (N_5416,N_2151,N_3146);
or U5417 (N_5417,N_2736,N_3895);
xnor U5418 (N_5418,N_2297,N_2519);
nor U5419 (N_5419,N_2361,N_2706);
nor U5420 (N_5420,N_2424,N_3441);
nor U5421 (N_5421,N_2935,N_3891);
and U5422 (N_5422,N_2525,N_3617);
nand U5423 (N_5423,N_3749,N_3439);
xnor U5424 (N_5424,N_2288,N_3507);
and U5425 (N_5425,N_3594,N_2210);
or U5426 (N_5426,N_3648,N_2974);
and U5427 (N_5427,N_2757,N_2120);
xnor U5428 (N_5428,N_3328,N_3544);
nor U5429 (N_5429,N_3672,N_3295);
or U5430 (N_5430,N_3845,N_2746);
nor U5431 (N_5431,N_2448,N_2957);
and U5432 (N_5432,N_3962,N_3090);
or U5433 (N_5433,N_2620,N_2831);
and U5434 (N_5434,N_3519,N_2825);
or U5435 (N_5435,N_3004,N_2858);
or U5436 (N_5436,N_2145,N_3973);
xnor U5437 (N_5437,N_2949,N_3654);
nand U5438 (N_5438,N_3129,N_3027);
xnor U5439 (N_5439,N_2875,N_3286);
or U5440 (N_5440,N_3458,N_3640);
and U5441 (N_5441,N_3829,N_2796);
and U5442 (N_5442,N_2421,N_3293);
nand U5443 (N_5443,N_3480,N_3245);
nand U5444 (N_5444,N_3279,N_2672);
nor U5445 (N_5445,N_3008,N_3757);
or U5446 (N_5446,N_3802,N_3149);
nor U5447 (N_5447,N_2707,N_3952);
xnor U5448 (N_5448,N_2691,N_2259);
and U5449 (N_5449,N_3516,N_2599);
xnor U5450 (N_5450,N_2417,N_2028);
xnor U5451 (N_5451,N_3693,N_2275);
and U5452 (N_5452,N_3283,N_2112);
xor U5453 (N_5453,N_2371,N_2407);
or U5454 (N_5454,N_2735,N_3700);
nand U5455 (N_5455,N_2794,N_3057);
xor U5456 (N_5456,N_3507,N_2641);
and U5457 (N_5457,N_3582,N_2040);
xnor U5458 (N_5458,N_3842,N_3495);
or U5459 (N_5459,N_2755,N_2495);
xnor U5460 (N_5460,N_2654,N_2983);
nand U5461 (N_5461,N_3284,N_3720);
and U5462 (N_5462,N_2679,N_2827);
or U5463 (N_5463,N_3837,N_2189);
nand U5464 (N_5464,N_3169,N_2736);
and U5465 (N_5465,N_3186,N_2974);
nand U5466 (N_5466,N_3623,N_3771);
nor U5467 (N_5467,N_3172,N_3109);
nand U5468 (N_5468,N_3972,N_3151);
nor U5469 (N_5469,N_2086,N_2074);
nor U5470 (N_5470,N_2373,N_2702);
nor U5471 (N_5471,N_2982,N_2287);
and U5472 (N_5472,N_2881,N_2547);
nor U5473 (N_5473,N_3353,N_2629);
xor U5474 (N_5474,N_2219,N_3692);
or U5475 (N_5475,N_3898,N_2978);
xnor U5476 (N_5476,N_3918,N_3925);
nand U5477 (N_5477,N_2286,N_2969);
nand U5478 (N_5478,N_3027,N_2523);
xnor U5479 (N_5479,N_2769,N_2776);
nand U5480 (N_5480,N_3780,N_3364);
and U5481 (N_5481,N_3117,N_2430);
or U5482 (N_5482,N_3501,N_2365);
xor U5483 (N_5483,N_3946,N_2338);
nand U5484 (N_5484,N_2325,N_2419);
nor U5485 (N_5485,N_2697,N_2699);
xor U5486 (N_5486,N_2308,N_3198);
nand U5487 (N_5487,N_2079,N_2267);
nor U5488 (N_5488,N_2854,N_3438);
or U5489 (N_5489,N_3079,N_3593);
or U5490 (N_5490,N_2516,N_3402);
xnor U5491 (N_5491,N_3928,N_3451);
xor U5492 (N_5492,N_3487,N_2926);
nand U5493 (N_5493,N_3233,N_3405);
or U5494 (N_5494,N_2465,N_2769);
xnor U5495 (N_5495,N_3696,N_3186);
or U5496 (N_5496,N_3922,N_3796);
or U5497 (N_5497,N_2131,N_3445);
xor U5498 (N_5498,N_3054,N_2734);
nor U5499 (N_5499,N_2952,N_3946);
nor U5500 (N_5500,N_3645,N_2557);
xor U5501 (N_5501,N_2751,N_2025);
nand U5502 (N_5502,N_3568,N_2721);
nor U5503 (N_5503,N_2406,N_3842);
nor U5504 (N_5504,N_3365,N_2920);
nor U5505 (N_5505,N_3233,N_2454);
nand U5506 (N_5506,N_2193,N_3938);
nand U5507 (N_5507,N_3019,N_2465);
and U5508 (N_5508,N_2440,N_2489);
or U5509 (N_5509,N_3298,N_3503);
nand U5510 (N_5510,N_2730,N_3964);
and U5511 (N_5511,N_3917,N_2582);
nor U5512 (N_5512,N_2659,N_2829);
nor U5513 (N_5513,N_2682,N_2944);
xor U5514 (N_5514,N_2530,N_3450);
nor U5515 (N_5515,N_3307,N_3438);
xor U5516 (N_5516,N_3040,N_2490);
xnor U5517 (N_5517,N_3942,N_3524);
nor U5518 (N_5518,N_3517,N_3853);
or U5519 (N_5519,N_3827,N_2458);
or U5520 (N_5520,N_2314,N_2392);
or U5521 (N_5521,N_2618,N_3531);
or U5522 (N_5522,N_3420,N_3615);
and U5523 (N_5523,N_3388,N_2998);
xnor U5524 (N_5524,N_2405,N_2103);
nor U5525 (N_5525,N_2366,N_3659);
nand U5526 (N_5526,N_3573,N_2428);
xor U5527 (N_5527,N_2557,N_2802);
nand U5528 (N_5528,N_3790,N_2998);
nor U5529 (N_5529,N_2312,N_3952);
xor U5530 (N_5530,N_2306,N_3659);
xnor U5531 (N_5531,N_2109,N_2743);
nand U5532 (N_5532,N_3735,N_3107);
and U5533 (N_5533,N_3319,N_2272);
xor U5534 (N_5534,N_2971,N_3683);
nor U5535 (N_5535,N_2712,N_3370);
xnor U5536 (N_5536,N_3580,N_3742);
and U5537 (N_5537,N_3043,N_2560);
xnor U5538 (N_5538,N_2007,N_3349);
or U5539 (N_5539,N_2351,N_3539);
xnor U5540 (N_5540,N_3496,N_2946);
or U5541 (N_5541,N_2181,N_2935);
nor U5542 (N_5542,N_2181,N_2946);
nand U5543 (N_5543,N_2381,N_2127);
xor U5544 (N_5544,N_2798,N_3856);
and U5545 (N_5545,N_2803,N_3379);
and U5546 (N_5546,N_3175,N_3241);
xor U5547 (N_5547,N_3771,N_3869);
or U5548 (N_5548,N_2205,N_2024);
xnor U5549 (N_5549,N_2484,N_3194);
nand U5550 (N_5550,N_2901,N_2344);
nand U5551 (N_5551,N_3488,N_2548);
or U5552 (N_5552,N_3120,N_3531);
xor U5553 (N_5553,N_2512,N_3994);
or U5554 (N_5554,N_3390,N_3673);
nor U5555 (N_5555,N_3531,N_3035);
or U5556 (N_5556,N_2954,N_2646);
nand U5557 (N_5557,N_3660,N_3927);
nor U5558 (N_5558,N_2483,N_2515);
and U5559 (N_5559,N_2433,N_3840);
nand U5560 (N_5560,N_2991,N_2025);
nand U5561 (N_5561,N_2880,N_3454);
xor U5562 (N_5562,N_2446,N_3328);
nor U5563 (N_5563,N_2231,N_2394);
xor U5564 (N_5564,N_2262,N_2141);
or U5565 (N_5565,N_2012,N_3640);
and U5566 (N_5566,N_3580,N_2994);
xor U5567 (N_5567,N_3005,N_2405);
nand U5568 (N_5568,N_3320,N_3446);
nor U5569 (N_5569,N_3512,N_3200);
and U5570 (N_5570,N_3099,N_3062);
xnor U5571 (N_5571,N_2770,N_2268);
xnor U5572 (N_5572,N_3041,N_2448);
nand U5573 (N_5573,N_3703,N_2640);
xor U5574 (N_5574,N_2616,N_3450);
nor U5575 (N_5575,N_3186,N_3483);
nand U5576 (N_5576,N_3680,N_3647);
and U5577 (N_5577,N_3046,N_2558);
nor U5578 (N_5578,N_2661,N_3898);
nand U5579 (N_5579,N_3047,N_2745);
and U5580 (N_5580,N_2969,N_3605);
and U5581 (N_5581,N_2968,N_3589);
xor U5582 (N_5582,N_3394,N_3038);
and U5583 (N_5583,N_2863,N_3030);
and U5584 (N_5584,N_2993,N_3599);
and U5585 (N_5585,N_3256,N_3598);
or U5586 (N_5586,N_2128,N_2228);
and U5587 (N_5587,N_3240,N_3794);
nand U5588 (N_5588,N_3678,N_3184);
xnor U5589 (N_5589,N_3048,N_2608);
nor U5590 (N_5590,N_3489,N_3253);
nor U5591 (N_5591,N_3083,N_2623);
and U5592 (N_5592,N_2584,N_2937);
xor U5593 (N_5593,N_2017,N_3395);
or U5594 (N_5594,N_2733,N_3373);
or U5595 (N_5595,N_2393,N_2059);
nand U5596 (N_5596,N_3497,N_3294);
or U5597 (N_5597,N_2020,N_3953);
and U5598 (N_5598,N_2739,N_2804);
nand U5599 (N_5599,N_2934,N_3685);
and U5600 (N_5600,N_3418,N_3642);
xor U5601 (N_5601,N_3473,N_3508);
nand U5602 (N_5602,N_2974,N_3834);
or U5603 (N_5603,N_2830,N_2644);
and U5604 (N_5604,N_3441,N_2562);
or U5605 (N_5605,N_3372,N_3553);
xor U5606 (N_5606,N_2063,N_2751);
and U5607 (N_5607,N_3190,N_3489);
and U5608 (N_5608,N_2331,N_3765);
xor U5609 (N_5609,N_2485,N_2384);
xor U5610 (N_5610,N_2454,N_2985);
nand U5611 (N_5611,N_2538,N_2810);
nand U5612 (N_5612,N_3792,N_3292);
or U5613 (N_5613,N_2764,N_3096);
nand U5614 (N_5614,N_3057,N_3550);
nand U5615 (N_5615,N_3136,N_2768);
and U5616 (N_5616,N_2591,N_2336);
xnor U5617 (N_5617,N_3849,N_3854);
xnor U5618 (N_5618,N_3528,N_2172);
and U5619 (N_5619,N_3382,N_3558);
nor U5620 (N_5620,N_3474,N_3340);
and U5621 (N_5621,N_2269,N_2602);
nor U5622 (N_5622,N_3023,N_3281);
or U5623 (N_5623,N_3386,N_2669);
nand U5624 (N_5624,N_3378,N_2905);
or U5625 (N_5625,N_2982,N_2200);
and U5626 (N_5626,N_3858,N_2393);
nand U5627 (N_5627,N_3259,N_2746);
nand U5628 (N_5628,N_3597,N_2337);
xnor U5629 (N_5629,N_2469,N_3051);
and U5630 (N_5630,N_3991,N_2161);
xor U5631 (N_5631,N_2968,N_2819);
xnor U5632 (N_5632,N_2571,N_2668);
xor U5633 (N_5633,N_3568,N_2744);
nand U5634 (N_5634,N_2709,N_2178);
xnor U5635 (N_5635,N_2547,N_3750);
and U5636 (N_5636,N_3499,N_3545);
or U5637 (N_5637,N_3128,N_3140);
xor U5638 (N_5638,N_3307,N_2140);
or U5639 (N_5639,N_3194,N_2135);
and U5640 (N_5640,N_3913,N_2790);
or U5641 (N_5641,N_3712,N_2595);
nor U5642 (N_5642,N_2671,N_2210);
xnor U5643 (N_5643,N_2313,N_3650);
nor U5644 (N_5644,N_2577,N_3259);
and U5645 (N_5645,N_3581,N_3656);
nor U5646 (N_5646,N_2318,N_2171);
nand U5647 (N_5647,N_2751,N_3195);
xor U5648 (N_5648,N_2504,N_2470);
nor U5649 (N_5649,N_3362,N_3035);
and U5650 (N_5650,N_3586,N_3987);
nor U5651 (N_5651,N_3635,N_3962);
nor U5652 (N_5652,N_3084,N_2872);
xnor U5653 (N_5653,N_3303,N_2519);
nand U5654 (N_5654,N_3251,N_2909);
nand U5655 (N_5655,N_3029,N_2816);
nand U5656 (N_5656,N_2164,N_2294);
and U5657 (N_5657,N_3279,N_2582);
or U5658 (N_5658,N_3976,N_3502);
or U5659 (N_5659,N_3433,N_3370);
and U5660 (N_5660,N_3394,N_3875);
or U5661 (N_5661,N_2603,N_2456);
xnor U5662 (N_5662,N_2145,N_3560);
nor U5663 (N_5663,N_2531,N_2043);
or U5664 (N_5664,N_2946,N_3612);
nand U5665 (N_5665,N_2802,N_2542);
nor U5666 (N_5666,N_3926,N_3553);
nor U5667 (N_5667,N_2045,N_2155);
nand U5668 (N_5668,N_3525,N_2301);
and U5669 (N_5669,N_3987,N_2407);
xnor U5670 (N_5670,N_3950,N_3789);
or U5671 (N_5671,N_2112,N_2127);
or U5672 (N_5672,N_3171,N_3783);
nand U5673 (N_5673,N_3301,N_2486);
nand U5674 (N_5674,N_2428,N_3093);
xor U5675 (N_5675,N_2015,N_3196);
xor U5676 (N_5676,N_3018,N_2438);
and U5677 (N_5677,N_3195,N_3130);
xnor U5678 (N_5678,N_2186,N_2869);
nand U5679 (N_5679,N_2955,N_2521);
and U5680 (N_5680,N_3384,N_2513);
xnor U5681 (N_5681,N_2474,N_3978);
or U5682 (N_5682,N_2434,N_3784);
or U5683 (N_5683,N_2370,N_3824);
or U5684 (N_5684,N_3780,N_3805);
nor U5685 (N_5685,N_2257,N_2062);
nor U5686 (N_5686,N_3322,N_3601);
and U5687 (N_5687,N_2633,N_3482);
and U5688 (N_5688,N_3197,N_3759);
nor U5689 (N_5689,N_3481,N_2735);
xor U5690 (N_5690,N_2879,N_3503);
nor U5691 (N_5691,N_2547,N_3944);
and U5692 (N_5692,N_2863,N_2317);
xor U5693 (N_5693,N_2085,N_3444);
nor U5694 (N_5694,N_3878,N_2093);
and U5695 (N_5695,N_2978,N_2430);
nor U5696 (N_5696,N_2211,N_2578);
and U5697 (N_5697,N_2720,N_2799);
xnor U5698 (N_5698,N_3767,N_3676);
nand U5699 (N_5699,N_3658,N_3276);
nand U5700 (N_5700,N_3184,N_2037);
nand U5701 (N_5701,N_2109,N_2258);
nand U5702 (N_5702,N_3276,N_2826);
or U5703 (N_5703,N_2314,N_3493);
xor U5704 (N_5704,N_2886,N_3290);
and U5705 (N_5705,N_3351,N_2614);
nor U5706 (N_5706,N_2029,N_3996);
nand U5707 (N_5707,N_2788,N_3416);
nor U5708 (N_5708,N_3791,N_3510);
or U5709 (N_5709,N_2837,N_2456);
nand U5710 (N_5710,N_2890,N_2215);
and U5711 (N_5711,N_2132,N_2905);
nor U5712 (N_5712,N_2622,N_2777);
and U5713 (N_5713,N_2465,N_2511);
xor U5714 (N_5714,N_2916,N_3426);
xnor U5715 (N_5715,N_3908,N_3076);
nand U5716 (N_5716,N_2960,N_2077);
or U5717 (N_5717,N_3715,N_2046);
and U5718 (N_5718,N_3888,N_3468);
xor U5719 (N_5719,N_3643,N_3904);
and U5720 (N_5720,N_2848,N_2288);
xnor U5721 (N_5721,N_2843,N_3346);
and U5722 (N_5722,N_3547,N_3351);
or U5723 (N_5723,N_2333,N_2155);
and U5724 (N_5724,N_2297,N_3488);
xnor U5725 (N_5725,N_2901,N_2742);
or U5726 (N_5726,N_2796,N_2547);
or U5727 (N_5727,N_2371,N_3986);
xnor U5728 (N_5728,N_2290,N_3785);
or U5729 (N_5729,N_2560,N_2202);
and U5730 (N_5730,N_2988,N_3721);
nand U5731 (N_5731,N_3273,N_3771);
xnor U5732 (N_5732,N_3633,N_2946);
xor U5733 (N_5733,N_3434,N_2929);
xor U5734 (N_5734,N_3095,N_3926);
xor U5735 (N_5735,N_2533,N_3359);
and U5736 (N_5736,N_2264,N_2161);
nor U5737 (N_5737,N_3991,N_2947);
nand U5738 (N_5738,N_2113,N_3460);
xor U5739 (N_5739,N_3884,N_2779);
nand U5740 (N_5740,N_2447,N_2587);
nand U5741 (N_5741,N_3004,N_2446);
or U5742 (N_5742,N_3692,N_2559);
nand U5743 (N_5743,N_2186,N_3383);
or U5744 (N_5744,N_3759,N_2536);
nand U5745 (N_5745,N_2593,N_2009);
xnor U5746 (N_5746,N_3512,N_3397);
nor U5747 (N_5747,N_3286,N_2434);
or U5748 (N_5748,N_3531,N_3945);
or U5749 (N_5749,N_3308,N_2651);
and U5750 (N_5750,N_3207,N_2581);
nor U5751 (N_5751,N_3083,N_3813);
nor U5752 (N_5752,N_2483,N_2160);
nand U5753 (N_5753,N_2307,N_2207);
or U5754 (N_5754,N_2142,N_2910);
nand U5755 (N_5755,N_2630,N_2153);
xnor U5756 (N_5756,N_2085,N_3831);
or U5757 (N_5757,N_2255,N_3416);
xnor U5758 (N_5758,N_2066,N_3033);
and U5759 (N_5759,N_3714,N_3987);
or U5760 (N_5760,N_3752,N_2155);
xor U5761 (N_5761,N_2882,N_2104);
nor U5762 (N_5762,N_3703,N_3028);
xnor U5763 (N_5763,N_3871,N_2633);
xor U5764 (N_5764,N_2569,N_2857);
xor U5765 (N_5765,N_2608,N_2333);
or U5766 (N_5766,N_3960,N_2864);
xor U5767 (N_5767,N_2180,N_3908);
nand U5768 (N_5768,N_2966,N_3783);
or U5769 (N_5769,N_2883,N_2555);
nor U5770 (N_5770,N_3857,N_3787);
and U5771 (N_5771,N_3095,N_3890);
and U5772 (N_5772,N_2456,N_2265);
or U5773 (N_5773,N_2295,N_3042);
xnor U5774 (N_5774,N_2564,N_3372);
xnor U5775 (N_5775,N_3167,N_3925);
and U5776 (N_5776,N_2930,N_2184);
nor U5777 (N_5777,N_3719,N_3869);
and U5778 (N_5778,N_2384,N_2865);
nand U5779 (N_5779,N_2252,N_2889);
nor U5780 (N_5780,N_2148,N_2516);
xor U5781 (N_5781,N_2361,N_3841);
xnor U5782 (N_5782,N_2538,N_2914);
and U5783 (N_5783,N_3524,N_2853);
nand U5784 (N_5784,N_2713,N_3496);
or U5785 (N_5785,N_2627,N_2997);
xor U5786 (N_5786,N_3581,N_3508);
nor U5787 (N_5787,N_3287,N_2421);
nor U5788 (N_5788,N_3974,N_3373);
or U5789 (N_5789,N_3285,N_2081);
nor U5790 (N_5790,N_3661,N_2650);
xor U5791 (N_5791,N_3665,N_3919);
and U5792 (N_5792,N_2471,N_3176);
or U5793 (N_5793,N_2521,N_2212);
xnor U5794 (N_5794,N_3866,N_3334);
and U5795 (N_5795,N_3477,N_3907);
nand U5796 (N_5796,N_2258,N_2153);
or U5797 (N_5797,N_2518,N_2329);
or U5798 (N_5798,N_2646,N_2150);
and U5799 (N_5799,N_2969,N_2347);
nand U5800 (N_5800,N_2305,N_3410);
nand U5801 (N_5801,N_2288,N_2426);
xor U5802 (N_5802,N_3142,N_2362);
and U5803 (N_5803,N_3676,N_3941);
nand U5804 (N_5804,N_3371,N_3021);
nor U5805 (N_5805,N_3956,N_3549);
or U5806 (N_5806,N_3888,N_2900);
xor U5807 (N_5807,N_2140,N_2076);
nand U5808 (N_5808,N_2610,N_3196);
or U5809 (N_5809,N_2609,N_2474);
or U5810 (N_5810,N_3192,N_2769);
or U5811 (N_5811,N_2580,N_2777);
nor U5812 (N_5812,N_3024,N_3701);
and U5813 (N_5813,N_2433,N_3586);
nand U5814 (N_5814,N_3164,N_2545);
nand U5815 (N_5815,N_2129,N_3074);
nand U5816 (N_5816,N_3040,N_2203);
and U5817 (N_5817,N_2777,N_2477);
nand U5818 (N_5818,N_2776,N_2387);
nor U5819 (N_5819,N_2966,N_2559);
or U5820 (N_5820,N_2414,N_2520);
and U5821 (N_5821,N_2279,N_2523);
nand U5822 (N_5822,N_2029,N_2267);
or U5823 (N_5823,N_3635,N_2319);
or U5824 (N_5824,N_3081,N_3011);
xor U5825 (N_5825,N_2182,N_2614);
and U5826 (N_5826,N_2362,N_2807);
nor U5827 (N_5827,N_2235,N_2934);
or U5828 (N_5828,N_3504,N_3383);
and U5829 (N_5829,N_3988,N_2004);
nand U5830 (N_5830,N_3930,N_2164);
xor U5831 (N_5831,N_2405,N_2824);
and U5832 (N_5832,N_2260,N_2321);
nor U5833 (N_5833,N_2789,N_3985);
or U5834 (N_5834,N_2612,N_2745);
xnor U5835 (N_5835,N_3944,N_2830);
nor U5836 (N_5836,N_3954,N_3019);
or U5837 (N_5837,N_3891,N_3532);
and U5838 (N_5838,N_3709,N_3674);
and U5839 (N_5839,N_2112,N_2819);
and U5840 (N_5840,N_2914,N_2564);
or U5841 (N_5841,N_2574,N_2390);
xor U5842 (N_5842,N_3438,N_2710);
nand U5843 (N_5843,N_2974,N_3661);
nand U5844 (N_5844,N_2100,N_3880);
xnor U5845 (N_5845,N_2770,N_2695);
and U5846 (N_5846,N_2384,N_2881);
and U5847 (N_5847,N_3743,N_3990);
or U5848 (N_5848,N_3495,N_2945);
and U5849 (N_5849,N_3630,N_3831);
and U5850 (N_5850,N_3088,N_3016);
or U5851 (N_5851,N_3658,N_3154);
xnor U5852 (N_5852,N_3214,N_2990);
nor U5853 (N_5853,N_3485,N_2319);
or U5854 (N_5854,N_3582,N_3940);
and U5855 (N_5855,N_3897,N_3432);
nor U5856 (N_5856,N_3279,N_2606);
nor U5857 (N_5857,N_2180,N_3031);
nor U5858 (N_5858,N_3855,N_2542);
and U5859 (N_5859,N_3281,N_2890);
xnor U5860 (N_5860,N_3058,N_2955);
nor U5861 (N_5861,N_2452,N_2634);
xnor U5862 (N_5862,N_2263,N_2425);
nor U5863 (N_5863,N_3931,N_3735);
nor U5864 (N_5864,N_3992,N_2049);
xor U5865 (N_5865,N_2853,N_2519);
nor U5866 (N_5866,N_3496,N_3789);
nor U5867 (N_5867,N_2039,N_2091);
nor U5868 (N_5868,N_3888,N_2339);
nor U5869 (N_5869,N_3771,N_3445);
nand U5870 (N_5870,N_3960,N_3588);
or U5871 (N_5871,N_3463,N_2004);
and U5872 (N_5872,N_2154,N_3073);
or U5873 (N_5873,N_3344,N_2874);
nor U5874 (N_5874,N_2054,N_2899);
nand U5875 (N_5875,N_3316,N_3895);
nand U5876 (N_5876,N_2460,N_3511);
nor U5877 (N_5877,N_3632,N_3143);
nor U5878 (N_5878,N_3118,N_2258);
and U5879 (N_5879,N_2936,N_3763);
nand U5880 (N_5880,N_3451,N_3800);
xor U5881 (N_5881,N_2467,N_2481);
nand U5882 (N_5882,N_2371,N_3582);
and U5883 (N_5883,N_3970,N_3397);
nor U5884 (N_5884,N_2143,N_2323);
and U5885 (N_5885,N_3190,N_2014);
and U5886 (N_5886,N_3150,N_2971);
xnor U5887 (N_5887,N_2130,N_3175);
xnor U5888 (N_5888,N_2730,N_2713);
or U5889 (N_5889,N_2346,N_3256);
or U5890 (N_5890,N_2381,N_2281);
and U5891 (N_5891,N_2154,N_3286);
and U5892 (N_5892,N_2153,N_3957);
and U5893 (N_5893,N_2212,N_3282);
nand U5894 (N_5894,N_2450,N_3274);
xnor U5895 (N_5895,N_3395,N_2677);
and U5896 (N_5896,N_3224,N_3294);
xor U5897 (N_5897,N_2362,N_3527);
or U5898 (N_5898,N_2091,N_3202);
or U5899 (N_5899,N_3538,N_3694);
nor U5900 (N_5900,N_3356,N_2186);
nor U5901 (N_5901,N_2712,N_2317);
nand U5902 (N_5902,N_3910,N_3336);
nand U5903 (N_5903,N_2463,N_3400);
or U5904 (N_5904,N_3216,N_3689);
nand U5905 (N_5905,N_3152,N_2896);
xnor U5906 (N_5906,N_2843,N_3275);
or U5907 (N_5907,N_3399,N_3095);
or U5908 (N_5908,N_2695,N_3590);
and U5909 (N_5909,N_2657,N_2480);
and U5910 (N_5910,N_3019,N_3343);
or U5911 (N_5911,N_3467,N_2379);
or U5912 (N_5912,N_2857,N_3289);
nor U5913 (N_5913,N_3821,N_3272);
or U5914 (N_5914,N_2901,N_2885);
nand U5915 (N_5915,N_2148,N_3035);
xor U5916 (N_5916,N_2373,N_2038);
xor U5917 (N_5917,N_3424,N_3580);
or U5918 (N_5918,N_2053,N_3199);
xor U5919 (N_5919,N_3450,N_3231);
nand U5920 (N_5920,N_3600,N_2066);
and U5921 (N_5921,N_2459,N_3880);
xnor U5922 (N_5922,N_3575,N_3140);
nand U5923 (N_5923,N_3770,N_2798);
nand U5924 (N_5924,N_2279,N_3722);
nor U5925 (N_5925,N_3091,N_3517);
nand U5926 (N_5926,N_3360,N_2717);
nand U5927 (N_5927,N_3327,N_2410);
nor U5928 (N_5928,N_2621,N_3334);
nand U5929 (N_5929,N_3365,N_3614);
or U5930 (N_5930,N_3843,N_3200);
nand U5931 (N_5931,N_3167,N_2943);
nor U5932 (N_5932,N_3164,N_2469);
nor U5933 (N_5933,N_3759,N_2797);
nand U5934 (N_5934,N_2937,N_3904);
nor U5935 (N_5935,N_2398,N_3082);
nand U5936 (N_5936,N_2659,N_3748);
xor U5937 (N_5937,N_2780,N_3857);
xor U5938 (N_5938,N_3306,N_2010);
nand U5939 (N_5939,N_2661,N_2989);
and U5940 (N_5940,N_3109,N_3199);
xor U5941 (N_5941,N_3795,N_3552);
xor U5942 (N_5942,N_2678,N_3203);
nor U5943 (N_5943,N_2054,N_3857);
nor U5944 (N_5944,N_3659,N_2866);
nand U5945 (N_5945,N_2522,N_3210);
and U5946 (N_5946,N_2660,N_3492);
nor U5947 (N_5947,N_2546,N_3108);
and U5948 (N_5948,N_3433,N_2743);
nand U5949 (N_5949,N_3790,N_2562);
and U5950 (N_5950,N_3015,N_3582);
xor U5951 (N_5951,N_2513,N_2475);
or U5952 (N_5952,N_2143,N_3786);
or U5953 (N_5953,N_3167,N_2066);
and U5954 (N_5954,N_3315,N_2112);
and U5955 (N_5955,N_3087,N_2389);
and U5956 (N_5956,N_3015,N_3269);
nand U5957 (N_5957,N_3347,N_3800);
or U5958 (N_5958,N_3325,N_3001);
nor U5959 (N_5959,N_2381,N_2961);
or U5960 (N_5960,N_2254,N_3055);
xnor U5961 (N_5961,N_2004,N_3436);
xor U5962 (N_5962,N_2322,N_2455);
and U5963 (N_5963,N_3508,N_2905);
or U5964 (N_5964,N_3815,N_3866);
nor U5965 (N_5965,N_2326,N_2137);
nor U5966 (N_5966,N_2091,N_2304);
nor U5967 (N_5967,N_3590,N_3955);
and U5968 (N_5968,N_2012,N_3745);
nand U5969 (N_5969,N_3172,N_2330);
and U5970 (N_5970,N_3941,N_2568);
xnor U5971 (N_5971,N_2863,N_3756);
xor U5972 (N_5972,N_2015,N_2458);
nor U5973 (N_5973,N_2961,N_2256);
and U5974 (N_5974,N_2472,N_3672);
and U5975 (N_5975,N_3241,N_2192);
nor U5976 (N_5976,N_3597,N_2632);
and U5977 (N_5977,N_2585,N_3048);
nand U5978 (N_5978,N_2198,N_3400);
and U5979 (N_5979,N_2558,N_3871);
nor U5980 (N_5980,N_2025,N_2194);
nor U5981 (N_5981,N_3374,N_2387);
or U5982 (N_5982,N_2038,N_3794);
or U5983 (N_5983,N_2925,N_2159);
nor U5984 (N_5984,N_2897,N_3464);
and U5985 (N_5985,N_2630,N_2582);
and U5986 (N_5986,N_2298,N_2940);
nor U5987 (N_5987,N_3034,N_2332);
nor U5988 (N_5988,N_3245,N_2724);
nand U5989 (N_5989,N_3968,N_3885);
xor U5990 (N_5990,N_3164,N_2017);
and U5991 (N_5991,N_2089,N_3243);
and U5992 (N_5992,N_3516,N_2027);
xor U5993 (N_5993,N_2339,N_3366);
nand U5994 (N_5994,N_2252,N_3980);
and U5995 (N_5995,N_2137,N_3165);
or U5996 (N_5996,N_3254,N_2067);
and U5997 (N_5997,N_2156,N_3371);
nor U5998 (N_5998,N_3051,N_3702);
or U5999 (N_5999,N_3821,N_3761);
nor U6000 (N_6000,N_4490,N_4020);
xor U6001 (N_6001,N_4353,N_4595);
and U6002 (N_6002,N_5965,N_5598);
and U6003 (N_6003,N_5955,N_5395);
or U6004 (N_6004,N_5613,N_4034);
and U6005 (N_6005,N_4513,N_5594);
nand U6006 (N_6006,N_4919,N_4845);
nand U6007 (N_6007,N_4197,N_5564);
and U6008 (N_6008,N_4665,N_5152);
or U6009 (N_6009,N_4142,N_5762);
nand U6010 (N_6010,N_4159,N_4618);
nor U6011 (N_6011,N_5056,N_4766);
nor U6012 (N_6012,N_5614,N_5209);
nand U6013 (N_6013,N_5972,N_5802);
nand U6014 (N_6014,N_5051,N_4785);
xor U6015 (N_6015,N_4322,N_5497);
nand U6016 (N_6016,N_4558,N_4327);
xor U6017 (N_6017,N_5247,N_5911);
nand U6018 (N_6018,N_5373,N_5446);
nand U6019 (N_6019,N_5898,N_5796);
nor U6020 (N_6020,N_5544,N_4896);
xnor U6021 (N_6021,N_4902,N_5007);
and U6022 (N_6022,N_4920,N_5857);
xor U6023 (N_6023,N_5738,N_4105);
xnor U6024 (N_6024,N_4072,N_4101);
and U6025 (N_6025,N_4257,N_5097);
nor U6026 (N_6026,N_5513,N_4114);
nand U6027 (N_6027,N_5824,N_5347);
and U6028 (N_6028,N_5917,N_4024);
and U6029 (N_6029,N_4841,N_5145);
or U6030 (N_6030,N_5331,N_4404);
or U6031 (N_6031,N_5945,N_4053);
xor U6032 (N_6032,N_4640,N_4723);
nand U6033 (N_6033,N_4329,N_5916);
nand U6034 (N_6034,N_5084,N_4419);
and U6035 (N_6035,N_4393,N_4437);
or U6036 (N_6036,N_5677,N_5740);
or U6037 (N_6037,N_5341,N_4097);
nor U6038 (N_6038,N_4226,N_5474);
nand U6039 (N_6039,N_4363,N_5327);
nor U6040 (N_6040,N_4647,N_5646);
or U6041 (N_6041,N_5036,N_4143);
nand U6042 (N_6042,N_4914,N_4135);
or U6043 (N_6043,N_5833,N_4435);
nand U6044 (N_6044,N_4552,N_5786);
nor U6045 (N_6045,N_4050,N_4041);
xnor U6046 (N_6046,N_5835,N_5724);
nor U6047 (N_6047,N_4499,N_5063);
xnor U6048 (N_6048,N_4645,N_4265);
or U6049 (N_6049,N_4804,N_4094);
xor U6050 (N_6050,N_4317,N_4714);
xor U6051 (N_6051,N_5683,N_5280);
nand U6052 (N_6052,N_4198,N_5383);
nand U6053 (N_6053,N_5710,N_4729);
or U6054 (N_6054,N_5132,N_4995);
or U6055 (N_6055,N_5759,N_5548);
and U6056 (N_6056,N_4667,N_5805);
xnor U6057 (N_6057,N_4290,N_4463);
nand U6058 (N_6058,N_4999,N_4140);
nor U6059 (N_6059,N_5649,N_4055);
xnor U6060 (N_6060,N_4235,N_4282);
and U6061 (N_6061,N_5340,N_5180);
and U6062 (N_6062,N_4793,N_4854);
nand U6063 (N_6063,N_4958,N_5075);
nor U6064 (N_6064,N_4959,N_5483);
or U6065 (N_6065,N_4560,N_4954);
or U6066 (N_6066,N_5828,N_4989);
xor U6067 (N_6067,N_5581,N_5905);
nor U6068 (N_6068,N_5565,N_4724);
nand U6069 (N_6069,N_5142,N_4396);
and U6070 (N_6070,N_4763,N_4040);
nand U6071 (N_6071,N_4358,N_5221);
or U6072 (N_6072,N_4448,N_4739);
or U6073 (N_6073,N_4163,N_4104);
nand U6074 (N_6074,N_4690,N_4771);
nor U6075 (N_6075,N_5733,N_4984);
and U6076 (N_6076,N_4075,N_5187);
and U6077 (N_6077,N_5692,N_4616);
nand U6078 (N_6078,N_5644,N_4337);
or U6079 (N_6079,N_5354,N_5388);
xor U6080 (N_6080,N_4885,N_4921);
nor U6081 (N_6081,N_5231,N_4009);
xor U6082 (N_6082,N_4085,N_5454);
nand U6083 (N_6083,N_4810,N_4298);
xnor U6084 (N_6084,N_4827,N_5355);
xor U6085 (N_6085,N_5700,N_4688);
and U6086 (N_6086,N_4203,N_5988);
nand U6087 (N_6087,N_5121,N_4798);
nand U6088 (N_6088,N_5682,N_5812);
nor U6089 (N_6089,N_4042,N_5936);
or U6090 (N_6090,N_5353,N_5458);
xor U6091 (N_6091,N_4023,N_5860);
and U6092 (N_6092,N_5987,N_4826);
nand U6093 (N_6093,N_5225,N_5502);
and U6094 (N_6094,N_4998,N_5727);
nand U6095 (N_6095,N_4100,N_5232);
nor U6096 (N_6096,N_4707,N_4415);
and U6097 (N_6097,N_5319,N_4225);
nand U6098 (N_6098,N_4286,N_5934);
or U6099 (N_6099,N_5204,N_4750);
nand U6100 (N_6100,N_4619,N_4658);
and U6101 (N_6101,N_4636,N_4588);
and U6102 (N_6102,N_5452,N_5848);
and U6103 (N_6103,N_4874,N_4518);
or U6104 (N_6104,N_5086,N_5018);
and U6105 (N_6105,N_5299,N_4343);
nand U6106 (N_6106,N_4745,N_5550);
nand U6107 (N_6107,N_5612,N_4234);
and U6108 (N_6108,N_4712,N_4017);
nand U6109 (N_6109,N_5892,N_5536);
and U6110 (N_6110,N_4474,N_5774);
xnor U6111 (N_6111,N_4576,N_5757);
nor U6112 (N_6112,N_4987,N_4078);
nand U6113 (N_6113,N_4746,N_4426);
xor U6114 (N_6114,N_4916,N_5694);
xnor U6115 (N_6115,N_5787,N_5509);
xor U6116 (N_6116,N_4335,N_5139);
and U6117 (N_6117,N_4506,N_5392);
xnor U6118 (N_6118,N_4856,N_4861);
xnor U6119 (N_6119,N_5306,N_4758);
nand U6120 (N_6120,N_4814,N_4735);
or U6121 (N_6121,N_5749,N_4797);
or U6122 (N_6122,N_5956,N_5432);
and U6123 (N_6123,N_5322,N_5661);
or U6124 (N_6124,N_5795,N_4007);
nand U6125 (N_6125,N_5167,N_5973);
xnor U6126 (N_6126,N_5830,N_5617);
and U6127 (N_6127,N_4162,N_5800);
and U6128 (N_6128,N_4825,N_5822);
nand U6129 (N_6129,N_4324,N_4529);
nand U6130 (N_6130,N_5950,N_5888);
and U6131 (N_6131,N_5706,N_5885);
or U6132 (N_6132,N_4439,N_4988);
and U6133 (N_6133,N_5920,N_5464);
and U6134 (N_6134,N_5198,N_4214);
xor U6135 (N_6135,N_4185,N_5140);
nor U6136 (N_6136,N_5029,N_5720);
nand U6137 (N_6137,N_4126,N_5503);
or U6138 (N_6138,N_5321,N_4220);
nor U6139 (N_6139,N_5397,N_4550);
nand U6140 (N_6140,N_4859,N_5815);
nand U6141 (N_6141,N_4939,N_4593);
nand U6142 (N_6142,N_4505,N_5393);
nor U6143 (N_6143,N_5270,N_4348);
and U6144 (N_6144,N_5557,N_4702);
xnor U6145 (N_6145,N_5978,N_5641);
nand U6146 (N_6146,N_4866,N_4720);
nor U6147 (N_6147,N_4123,N_5875);
and U6148 (N_6148,N_4212,N_4650);
nor U6149 (N_6149,N_5266,N_4762);
or U6150 (N_6150,N_4081,N_4487);
and U6151 (N_6151,N_5358,N_5348);
and U6152 (N_6152,N_4122,N_4744);
and U6153 (N_6153,N_5150,N_4389);
nor U6154 (N_6154,N_5635,N_5942);
nand U6155 (N_6155,N_4352,N_4498);
nand U6156 (N_6156,N_4218,N_5673);
xnor U6157 (N_6157,N_5567,N_5993);
nor U6158 (N_6158,N_4555,N_4124);
nand U6159 (N_6159,N_5085,N_4776);
nand U6160 (N_6160,N_5105,N_4803);
xnor U6161 (N_6161,N_4955,N_4256);
nand U6162 (N_6162,N_5357,N_4187);
nand U6163 (N_6163,N_5441,N_4992);
nor U6164 (N_6164,N_5870,N_5066);
and U6165 (N_6165,N_5074,N_4057);
xor U6166 (N_6166,N_4423,N_4013);
and U6167 (N_6167,N_4611,N_5559);
nor U6168 (N_6168,N_5017,N_4944);
nand U6169 (N_6169,N_5820,N_5995);
and U6170 (N_6170,N_5570,N_4457);
nand U6171 (N_6171,N_5171,N_5415);
nor U6172 (N_6172,N_5417,N_4003);
and U6173 (N_6173,N_5035,N_5400);
xnor U6174 (N_6174,N_5115,N_5623);
and U6175 (N_6175,N_5316,N_4131);
or U6176 (N_6176,N_5946,N_4093);
and U6177 (N_6177,N_4130,N_5494);
xnor U6178 (N_6178,N_4932,N_4682);
nand U6179 (N_6179,N_5839,N_4572);
nor U6180 (N_6180,N_4128,N_5450);
and U6181 (N_6181,N_5329,N_4546);
or U6182 (N_6182,N_4262,N_4355);
nand U6183 (N_6183,N_4508,N_5970);
xnor U6184 (N_6184,N_5268,N_4597);
nand U6185 (N_6185,N_5049,N_4068);
nor U6186 (N_6186,N_4509,N_5025);
nand U6187 (N_6187,N_4642,N_4300);
nor U6188 (N_6188,N_5194,N_5394);
or U6189 (N_6189,N_4165,N_4997);
and U6190 (N_6190,N_4086,N_4119);
and U6191 (N_6191,N_5118,N_4821);
xnor U6192 (N_6192,N_5588,N_5219);
nor U6193 (N_6193,N_4382,N_5421);
nor U6194 (N_6194,N_4191,N_4706);
or U6195 (N_6195,N_5527,N_5410);
xor U6196 (N_6196,N_5909,N_5678);
and U6197 (N_6197,N_5160,N_5052);
xnor U6198 (N_6198,N_4082,N_4301);
and U6199 (N_6199,N_5575,N_5931);
nand U6200 (N_6200,N_4943,N_5838);
or U6201 (N_6201,N_5289,N_5665);
xor U6202 (N_6202,N_4237,N_5237);
xnor U6203 (N_6203,N_4928,N_4855);
and U6204 (N_6204,N_5878,N_5591);
or U6205 (N_6205,N_4332,N_5496);
xor U6206 (N_6206,N_4133,N_5212);
and U6207 (N_6207,N_5010,N_4476);
or U6208 (N_6208,N_5825,N_4302);
and U6209 (N_6209,N_4510,N_4107);
or U6210 (N_6210,N_4087,N_5220);
nor U6211 (N_6211,N_5024,N_5624);
xnor U6212 (N_6212,N_4488,N_4189);
or U6213 (N_6213,N_5089,N_5271);
xnor U6214 (N_6214,N_4421,N_5137);
and U6215 (N_6215,N_5528,N_5420);
or U6216 (N_6216,N_5107,N_4217);
nor U6217 (N_6217,N_5182,N_4541);
or U6218 (N_6218,N_5077,N_5011);
nor U6219 (N_6219,N_5382,N_4065);
or U6220 (N_6220,N_5893,N_5255);
xor U6221 (N_6221,N_4378,N_5996);
nor U6222 (N_6222,N_4347,N_4772);
xnor U6223 (N_6223,N_5994,N_4501);
nand U6224 (N_6224,N_5076,N_4628);
and U6225 (N_6225,N_4018,N_4716);
or U6226 (N_6226,N_5504,N_4318);
xor U6227 (N_6227,N_5487,N_4395);
xor U6228 (N_6228,N_4931,N_4634);
xnor U6229 (N_6229,N_5098,N_5365);
or U6230 (N_6230,N_5758,N_5157);
xor U6231 (N_6231,N_4781,N_5293);
nand U6232 (N_6232,N_5718,N_5264);
or U6233 (N_6233,N_4076,N_5375);
or U6234 (N_6234,N_4408,N_5163);
nor U6235 (N_6235,N_4586,N_5980);
or U6236 (N_6236,N_5368,N_5267);
nand U6237 (N_6237,N_4503,N_4202);
and U6238 (N_6238,N_5478,N_5940);
nor U6239 (N_6239,N_5335,N_4346);
or U6240 (N_6240,N_4307,N_4651);
xnor U6241 (N_6241,N_5203,N_5214);
nand U6242 (N_6242,N_5574,N_5606);
nand U6243 (N_6243,N_5472,N_5073);
or U6244 (N_6244,N_5246,N_5190);
or U6245 (N_6245,N_5378,N_5431);
nand U6246 (N_6246,N_4479,N_4904);
nand U6247 (N_6247,N_4676,N_5654);
or U6248 (N_6248,N_4360,N_5957);
and U6249 (N_6249,N_5982,N_5855);
nand U6250 (N_6250,N_5999,N_5345);
nand U6251 (N_6251,N_5742,N_5664);
nand U6252 (N_6252,N_4878,N_5399);
or U6253 (N_6253,N_4548,N_5961);
and U6254 (N_6254,N_5104,N_4753);
nand U6255 (N_6255,N_5469,N_4111);
nand U6256 (N_6256,N_4542,N_5491);
and U6257 (N_6257,N_5897,N_4730);
xnor U6258 (N_6258,N_4014,N_5019);
xnor U6259 (N_6259,N_5064,N_5465);
nor U6260 (N_6260,N_5782,N_4371);
and U6261 (N_6261,N_4800,N_4264);
xnor U6262 (N_6262,N_4054,N_4258);
nand U6263 (N_6263,N_5041,N_4453);
nand U6264 (N_6264,N_5262,N_5379);
or U6265 (N_6265,N_4867,N_5261);
nand U6266 (N_6266,N_4801,N_4884);
xor U6267 (N_6267,N_5578,N_5879);
nor U6268 (N_6268,N_5638,N_4886);
xnor U6269 (N_6269,N_5989,N_4820);
nand U6270 (N_6270,N_5296,N_5881);
nand U6271 (N_6271,N_4691,N_5164);
or U6272 (N_6272,N_4917,N_4975);
nand U6273 (N_6273,N_5279,N_5585);
xor U6274 (N_6274,N_4493,N_4434);
xnor U6275 (N_6275,N_4166,N_5747);
nor U6276 (N_6276,N_5744,N_5769);
xnor U6277 (N_6277,N_4965,N_4183);
xnor U6278 (N_6278,N_5847,N_4269);
or U6279 (N_6279,N_4515,N_4227);
or U6280 (N_6280,N_5959,N_4231);
and U6281 (N_6281,N_4117,N_4045);
nor U6282 (N_6282,N_5320,N_5599);
nand U6283 (N_6283,N_5773,N_5055);
and U6284 (N_6284,N_4535,N_5087);
nand U6285 (N_6285,N_4540,N_5191);
or U6286 (N_6286,N_4146,N_5752);
nor U6287 (N_6287,N_4860,N_5236);
and U6288 (N_6288,N_5135,N_4116);
and U6289 (N_6289,N_5434,N_4005);
xnor U6290 (N_6290,N_4364,N_4000);
or U6291 (N_6291,N_4376,N_5185);
or U6292 (N_6292,N_5122,N_5584);
and U6293 (N_6293,N_4413,N_5026);
and U6294 (N_6294,N_5765,N_5113);
nand U6295 (N_6295,N_4653,N_5872);
nand U6296 (N_6296,N_5124,N_4900);
and U6297 (N_6297,N_5307,N_4551);
nand U6298 (N_6298,N_5111,N_5376);
xor U6299 (N_6299,N_4384,N_5147);
xnor U6300 (N_6300,N_4215,N_5770);
and U6301 (N_6301,N_5352,N_5736);
or U6302 (N_6302,N_5856,N_5645);
and U6303 (N_6303,N_4622,N_4794);
xor U6304 (N_6304,N_5981,N_5412);
or U6305 (N_6305,N_5958,N_4496);
xnor U6306 (N_6306,N_5159,N_4838);
or U6307 (N_6307,N_5501,N_4816);
and U6308 (N_6308,N_4211,N_4629);
nor U6309 (N_6309,N_4206,N_4848);
or U6310 (N_6310,N_5241,N_4566);
or U6311 (N_6311,N_5314,N_4134);
xor U6312 (N_6312,N_5863,N_4610);
nand U6313 (N_6313,N_4583,N_4443);
nor U6314 (N_6314,N_5760,N_5156);
and U6315 (N_6315,N_4788,N_5922);
nor U6316 (N_6316,N_5021,N_5873);
nand U6317 (N_6317,N_4177,N_4661);
or U6318 (N_6318,N_4281,N_4246);
xor U6319 (N_6319,N_5175,N_5719);
or U6320 (N_6320,N_4480,N_5748);
xor U6321 (N_6321,N_4216,N_4079);
or U6322 (N_6322,N_4406,N_4633);
xnor U6323 (N_6323,N_5633,N_4530);
and U6324 (N_6324,N_5334,N_4132);
or U6325 (N_6325,N_4233,N_5726);
or U6326 (N_6326,N_4938,N_4387);
nor U6327 (N_6327,N_4725,N_5138);
nor U6328 (N_6328,N_4339,N_5173);
nand U6329 (N_6329,N_5488,N_4747);
nand U6330 (N_6330,N_4627,N_4280);
nor U6331 (N_6331,N_4711,N_4924);
nor U6332 (N_6332,N_5510,N_4477);
nor U6333 (N_6333,N_5456,N_4314);
nor U6334 (N_6334,N_5858,N_4405);
xnor U6335 (N_6335,N_4727,N_4048);
or U6336 (N_6336,N_5523,N_5515);
or U6337 (N_6337,N_4656,N_5445);
nand U6338 (N_6338,N_5404,N_4812);
or U6339 (N_6339,N_5904,N_4492);
or U6340 (N_6340,N_4563,N_4767);
or U6341 (N_6341,N_5409,N_5034);
xor U6342 (N_6342,N_5826,N_4106);
and U6343 (N_6343,N_5014,N_4807);
nor U6344 (N_6344,N_4600,N_4775);
nor U6345 (N_6345,N_5545,N_4120);
nand U6346 (N_6346,N_5530,N_4210);
nand U6347 (N_6347,N_4674,N_4662);
or U6348 (N_6348,N_4241,N_4289);
xor U6349 (N_6349,N_4070,N_5696);
or U6350 (N_6350,N_4440,N_5439);
and U6351 (N_6351,N_4979,N_4063);
or U6352 (N_6352,N_5201,N_5475);
xnor U6353 (N_6353,N_5546,N_4313);
xnor U6354 (N_6354,N_5840,N_4209);
or U6355 (N_6355,N_4199,N_5648);
xor U6356 (N_6356,N_4580,N_5913);
xor U6357 (N_6357,N_5596,N_5846);
nor U6358 (N_6358,N_5088,N_4392);
nor U6359 (N_6359,N_5196,N_4004);
or U6360 (N_6360,N_4765,N_5324);
and U6361 (N_6361,N_5827,N_4430);
nand U6362 (N_6362,N_5100,N_4006);
and U6363 (N_6363,N_5932,N_5396);
xor U6364 (N_6364,N_5037,N_4742);
or U6365 (N_6365,N_5876,N_4125);
xnor U6366 (N_6366,N_5608,N_4303);
or U6367 (N_6367,N_4741,N_5625);
nor U6368 (N_6368,N_4685,N_5505);
nor U6369 (N_6369,N_4031,N_5803);
or U6370 (N_6370,N_4598,N_4952);
nand U6371 (N_6371,N_4178,N_4752);
nor U6372 (N_6372,N_4455,N_4088);
nand U6373 (N_6373,N_4467,N_5511);
nand U6374 (N_6374,N_4544,N_5615);
nor U6375 (N_6375,N_5914,N_5865);
nand U6376 (N_6376,N_4961,N_4773);
xnor U6377 (N_6377,N_4680,N_5667);
nor U6378 (N_6378,N_4442,N_4312);
and U6379 (N_6379,N_4584,N_5652);
or U6380 (N_6380,N_5402,N_4889);
nor U6381 (N_6381,N_4675,N_5944);
and U6382 (N_6382,N_4877,N_4468);
xor U6383 (N_6383,N_5377,N_4605);
or U6384 (N_6384,N_4731,N_4066);
or U6385 (N_6385,N_4171,N_4585);
xor U6386 (N_6386,N_5949,N_4748);
nor U6387 (N_6387,N_5659,N_5518);
nor U6388 (N_6388,N_5226,N_5778);
nor U6389 (N_6389,N_4915,N_5292);
and U6390 (N_6390,N_5535,N_4478);
nor U6391 (N_6391,N_5637,N_5701);
or U6392 (N_6392,N_5291,N_5405);
or U6393 (N_6393,N_5939,N_4843);
and U6394 (N_6394,N_4672,N_4868);
xnor U6395 (N_6395,N_4497,N_5093);
nor U6396 (N_6396,N_5133,N_5229);
xnor U6397 (N_6397,N_5886,N_4581);
nand U6398 (N_6398,N_5277,N_5273);
nand U6399 (N_6399,N_5031,N_5401);
and U6400 (N_6400,N_5123,N_4969);
or U6401 (N_6401,N_5764,N_4757);
xor U6402 (N_6402,N_5444,N_5729);
xor U6403 (N_6403,N_4922,N_4304);
xnor U6404 (N_6404,N_5583,N_5323);
or U6405 (N_6405,N_4858,N_5265);
nand U6406 (N_6406,N_4538,N_4458);
or U6407 (N_6407,N_4553,N_4657);
nor U6408 (N_6408,N_5172,N_4643);
nand U6409 (N_6409,N_5343,N_4652);
and U6410 (N_6410,N_5788,N_5941);
or U6411 (N_6411,N_4409,N_4532);
or U6412 (N_6412,N_5746,N_4981);
nor U6413 (N_6413,N_5416,N_4839);
nand U6414 (N_6414,N_4144,N_5068);
xor U6415 (N_6415,N_5880,N_5005);
and U6416 (N_6416,N_4096,N_5290);
xnor U6417 (N_6417,N_4589,N_5734);
xor U6418 (N_6418,N_5792,N_5813);
and U6419 (N_6419,N_5263,N_5679);
and U6420 (N_6420,N_4671,N_4710);
nand U6421 (N_6421,N_5466,N_5874);
and U6422 (N_6422,N_4578,N_5930);
and U6423 (N_6423,N_4913,N_4565);
or U6424 (N_6424,N_5808,N_4420);
nand U6425 (N_6425,N_4614,N_4677);
nor U6426 (N_6426,N_4470,N_5889);
or U6427 (N_6427,N_4980,N_5224);
xor U6428 (N_6428,N_5767,N_5676);
or U6429 (N_6429,N_5467,N_5038);
xnor U6430 (N_6430,N_4362,N_5817);
nor U6431 (N_6431,N_4876,N_4251);
xnor U6432 (N_6432,N_5176,N_4792);
xor U6433 (N_6433,N_4883,N_5553);
nand U6434 (N_6434,N_5604,N_4482);
xor U6435 (N_6435,N_4046,N_5042);
or U6436 (N_6436,N_4491,N_4894);
and U6437 (N_6437,N_4083,N_4181);
and U6438 (N_6438,N_5571,N_5568);
nand U6439 (N_6439,N_4447,N_4539);
or U6440 (N_6440,N_5315,N_5059);
and U6441 (N_6441,N_4986,N_4996);
xor U6442 (N_6442,N_4802,N_5109);
and U6443 (N_6443,N_5283,N_4077);
or U6444 (N_6444,N_4294,N_4719);
nor U6445 (N_6445,N_5902,N_4243);
and U6446 (N_6446,N_4974,N_4381);
or U6447 (N_6447,N_5520,N_5647);
nor U6448 (N_6448,N_4514,N_4779);
nor U6449 (N_6449,N_5883,N_5590);
and U6450 (N_6450,N_4912,N_4179);
xor U6451 (N_6451,N_5531,N_4507);
xnor U6452 (N_6452,N_4679,N_4942);
and U6453 (N_6453,N_4137,N_4032);
xor U6454 (N_6454,N_5020,N_5256);
and U6455 (N_6455,N_5754,N_5473);
nand U6456 (N_6456,N_4923,N_5816);
and U6457 (N_6457,N_4575,N_5361);
or U6458 (N_6458,N_5619,N_4722);
nand U6459 (N_6459,N_4127,N_5149);
nor U6460 (N_6460,N_4721,N_4930);
or U6461 (N_6461,N_4760,N_5609);
xnor U6462 (N_6462,N_5723,N_5630);
or U6463 (N_6463,N_4780,N_4167);
nor U6464 (N_6464,N_4273,N_5295);
xnor U6465 (N_6465,N_5338,N_5177);
or U6466 (N_6466,N_5709,N_5534);
xor U6467 (N_6467,N_4761,N_4664);
xnor U6468 (N_6468,N_4190,N_5436);
nand U6469 (N_6469,N_5065,N_4887);
and U6470 (N_6470,N_4475,N_4549);
or U6471 (N_6471,N_4905,N_4934);
xor U6472 (N_6472,N_4893,N_4242);
or U6473 (N_6473,N_5991,N_5776);
or U6474 (N_6474,N_5126,N_5387);
or U6475 (N_6475,N_4372,N_5205);
nor U6476 (N_6476,N_4279,N_5254);
nor U6477 (N_6477,N_4504,N_4051);
nor U6478 (N_6478,N_5526,N_4972);
xor U6479 (N_6479,N_5793,N_5285);
nand U6480 (N_6480,N_5811,N_5836);
nand U6481 (N_6481,N_4570,N_5882);
nand U6482 (N_6482,N_5542,N_5843);
and U6483 (N_6483,N_4873,N_5213);
or U6484 (N_6484,N_4603,N_4390);
nand U6485 (N_6485,N_4192,N_5852);
nand U6486 (N_6486,N_5197,N_5046);
or U6487 (N_6487,N_5463,N_4683);
nor U6488 (N_6488,N_4168,N_4402);
and U6489 (N_6489,N_4424,N_5114);
or U6490 (N_6490,N_5227,N_4784);
xnor U6491 (N_6491,N_4067,N_4109);
nand U6492 (N_6492,N_5566,N_4993);
nor U6493 (N_6493,N_5576,N_4933);
and U6494 (N_6494,N_4686,N_5428);
xor U6495 (N_6495,N_4840,N_5927);
or U6496 (N_6496,N_4485,N_4230);
xnor U6497 (N_6497,N_5422,N_4789);
nor U6498 (N_6498,N_4994,N_4293);
or U6499 (N_6499,N_4528,N_5351);
nand U6500 (N_6500,N_4909,N_4596);
nor U6501 (N_6501,N_5407,N_4321);
or U6502 (N_6502,N_5244,N_4407);
nand U6503 (N_6503,N_4615,N_4365);
nor U6504 (N_6504,N_5508,N_5714);
xor U6505 (N_6505,N_4521,N_5602);
and U6506 (N_6506,N_5971,N_5437);
or U6507 (N_6507,N_5771,N_5697);
or U6508 (N_6508,N_4047,N_5356);
nor U6509 (N_6509,N_4571,N_4153);
nand U6510 (N_6510,N_4935,N_5918);
or U6511 (N_6511,N_4815,N_4325);
xor U6512 (N_6512,N_5832,N_4607);
xnor U6513 (N_6513,N_4232,N_4666);
or U6514 (N_6514,N_4949,N_5006);
nor U6515 (N_6515,N_5912,N_5304);
or U6516 (N_6516,N_4222,N_4799);
nand U6517 (N_6517,N_5806,N_4774);
or U6518 (N_6518,N_5948,N_5610);
or U6519 (N_6519,N_5079,N_5082);
nand U6520 (N_6520,N_5935,N_4834);
xnor U6521 (N_6521,N_4268,N_4027);
or U6522 (N_6522,N_5929,N_5128);
xor U6523 (N_6523,N_4543,N_4386);
nand U6524 (N_6524,N_4002,N_4590);
and U6525 (N_6525,N_4342,N_4039);
xor U6526 (N_6526,N_5669,N_4410);
xnor U6527 (N_6527,N_4357,N_4240);
xnor U6528 (N_6528,N_4084,N_5374);
nor U6529 (N_6529,N_5618,N_4698);
nand U6530 (N_6530,N_4851,N_4161);
nand U6531 (N_6531,N_5924,N_5495);
nor U6532 (N_6532,N_5406,N_4733);
nor U6533 (N_6533,N_5200,N_4568);
nand U6534 (N_6534,N_5423,N_5626);
or U6535 (N_6535,N_5691,N_4907);
nand U6536 (N_6536,N_4473,N_4427);
nand U6537 (N_6537,N_4891,N_5443);
xor U6538 (N_6538,N_5310,N_5253);
xor U6539 (N_6539,N_4272,N_5453);
and U6540 (N_6540,N_5845,N_5698);
xnor U6541 (N_6541,N_5605,N_5485);
nand U6542 (N_6542,N_5558,N_5168);
nor U6543 (N_6543,N_4462,N_4253);
nor U6544 (N_6544,N_4091,N_5977);
xor U6545 (N_6545,N_5861,N_4863);
nand U6546 (N_6546,N_5223,N_4025);
nand U6547 (N_6547,N_5178,N_5642);
or U6548 (N_6548,N_5851,N_4641);
xor U6549 (N_6549,N_5695,N_5328);
xnor U6550 (N_6550,N_4061,N_5549);
nor U6551 (N_6551,N_4368,N_5516);
xor U6552 (N_6552,N_5850,N_5435);
or U6553 (N_6553,N_4383,N_4204);
and U6554 (N_6554,N_4968,N_5211);
xnor U6555 (N_6555,N_4296,N_5563);
nor U6556 (N_6556,N_4331,N_4369);
nor U6557 (N_6557,N_5592,N_4391);
or U6558 (N_6558,N_5660,N_5448);
nand U6559 (N_6559,N_4978,N_5819);
nor U6560 (N_6560,N_5524,N_5975);
nand U6561 (N_6561,N_5003,N_4606);
nor U6562 (N_6562,N_4228,N_5297);
xor U6563 (N_6563,N_4601,N_4869);
nand U6564 (N_6564,N_5326,N_5195);
xor U6565 (N_6565,N_4536,N_5976);
or U6566 (N_6566,N_4416,N_4617);
xor U6567 (N_6567,N_5442,N_4660);
nor U6568 (N_6568,N_5868,N_4613);
nand U6569 (N_6569,N_4344,N_5979);
or U6570 (N_6570,N_5433,N_4385);
nand U6571 (N_6571,N_4982,N_4186);
and U6572 (N_6572,N_4397,N_4121);
nor U6573 (N_6573,N_4239,N_5866);
nor U6574 (N_6574,N_4149,N_5027);
and U6575 (N_6575,N_4755,N_5438);
nand U6576 (N_6576,N_5867,N_5768);
and U6577 (N_6577,N_5146,N_5349);
or U6578 (N_6578,N_4694,N_4432);
xnor U6579 (N_6579,N_4831,N_4299);
and U6580 (N_6580,N_4323,N_4495);
nor U6581 (N_6581,N_4835,N_5317);
or U6582 (N_6582,N_4356,N_5992);
nor U6583 (N_6583,N_4564,N_4459);
nand U6584 (N_6584,N_4849,N_5968);
or U6585 (N_6585,N_4073,N_4305);
and U6586 (N_6586,N_4236,N_5910);
nand U6587 (N_6587,N_4890,N_5969);
or U6588 (N_6588,N_4361,N_5500);
or U6589 (N_6589,N_5070,N_5057);
or U6590 (N_6590,N_4783,N_4743);
nand U6591 (N_6591,N_5072,N_5622);
nand U6592 (N_6592,N_5154,N_5713);
xnor U6593 (N_6593,N_5414,N_4188);
nor U6594 (N_6594,N_4311,N_5344);
nor U6595 (N_6595,N_5997,N_5207);
or U6596 (N_6596,N_5990,N_4638);
and U6597 (N_6597,N_5044,N_4340);
xnor U6598 (N_6598,N_5215,N_4892);
nand U6599 (N_6599,N_4238,N_4033);
or U6600 (N_6600,N_4351,N_4059);
xnor U6601 (N_6601,N_5600,N_5896);
nand U6602 (N_6602,N_5984,N_4609);
or U6603 (N_6603,N_4275,N_5012);
nor U6604 (N_6604,N_5390,N_4824);
nor U6605 (N_6605,N_4836,N_4417);
nor U6606 (N_6606,N_4881,N_5298);
nor U6607 (N_6607,N_4819,N_4255);
and U6608 (N_6608,N_5325,N_5737);
or U6609 (N_6609,N_5350,N_4829);
or U6610 (N_6610,N_4879,N_4655);
nand U6611 (N_6611,N_4486,N_5419);
or U6612 (N_6612,N_5884,N_4697);
nor U6613 (N_6613,N_5360,N_5854);
and U6614 (N_6614,N_4811,N_5235);
nand U6615 (N_6615,N_5047,N_4791);
nand U6616 (N_6616,N_5675,N_4502);
nand U6617 (N_6617,N_4266,N_5117);
or U6618 (N_6618,N_4456,N_5887);
xor U6619 (N_6619,N_5258,N_4795);
nand U6620 (N_6620,N_4157,N_4052);
xnor U6621 (N_6621,N_4379,N_4545);
xor U6622 (N_6622,N_5589,N_5426);
nand U6623 (N_6623,N_4205,N_4394);
nor U6624 (N_6624,N_4759,N_5243);
and U6625 (N_6625,N_4950,N_5844);
nand U6626 (N_6626,N_5790,N_5091);
and U6627 (N_6627,N_5620,N_5842);
and U6628 (N_6628,N_5125,N_5722);
nor U6629 (N_6629,N_5921,N_4620);
nor U6630 (N_6630,N_5252,N_4095);
and U6631 (N_6631,N_5554,N_4768);
nor U6632 (N_6632,N_5490,N_5425);
xnor U6633 (N_6633,N_4533,N_4648);
xor U6634 (N_6634,N_4173,N_5339);
or U6635 (N_6635,N_5923,N_4537);
or U6636 (N_6636,N_5061,N_4145);
xor U6637 (N_6637,N_5189,N_4060);
nor U6638 (N_6638,N_5193,N_4782);
nor U6639 (N_6639,N_4700,N_5333);
nor U6640 (N_6640,N_5829,N_5242);
nand U6641 (N_6641,N_4172,N_5305);
nor U6642 (N_6642,N_4681,N_5208);
xnor U6643 (N_6643,N_5408,N_5477);
and U6644 (N_6644,N_4630,N_5631);
nand U6645 (N_6645,N_4956,N_5657);
nor U6646 (N_6646,N_4049,N_4673);
nand U6647 (N_6647,N_5486,N_4962);
xor U6648 (N_6648,N_5043,N_5460);
xor U6649 (N_6649,N_5169,N_4349);
nor U6650 (N_6650,N_5413,N_4983);
nor U6651 (N_6651,N_4012,N_5385);
nor U6652 (N_6652,N_4195,N_5687);
or U6653 (N_6653,N_4880,N_4870);
xnor U6654 (N_6654,N_4019,N_5781);
and U6655 (N_6655,N_4520,N_4951);
or U6656 (N_6656,N_4637,N_5048);
or U6657 (N_6657,N_4169,N_5841);
and U6658 (N_6658,N_4728,N_5183);
or U6659 (N_6659,N_4684,N_5798);
and U6660 (N_6660,N_5102,N_5103);
or U6661 (N_6661,N_5148,N_4201);
and U6662 (N_6662,N_4254,N_5312);
nand U6663 (N_6663,N_5772,N_4906);
nand U6664 (N_6664,N_4429,N_5045);
xnor U6665 (N_6665,N_4208,N_5251);
nand U6666 (N_6666,N_4283,N_5753);
xnor U6667 (N_6667,N_5529,N_4089);
xnor U6668 (N_6668,N_5457,N_5821);
or U6669 (N_6669,N_4026,N_5158);
or U6670 (N_6670,N_5777,N_4388);
xor U6671 (N_6671,N_4494,N_5804);
nand U6672 (N_6672,N_5095,N_4164);
and U6673 (N_6673,N_4527,N_5391);
nand U6674 (N_6674,N_5938,N_4852);
xor U6675 (N_6675,N_5489,N_4136);
xnor U6676 (N_6676,N_4830,N_5367);
xnor U6677 (N_6677,N_4367,N_5693);
and U6678 (N_6678,N_4850,N_4438);
or U6679 (N_6679,N_5302,N_5925);
nand U6680 (N_6680,N_4511,N_5040);
xor U6681 (N_6681,N_4341,N_4695);
nor U6682 (N_6682,N_5233,N_5096);
xnor U6683 (N_6683,N_5136,N_5640);
nor U6684 (N_6684,N_5092,N_5249);
nand U6685 (N_6685,N_4554,N_5634);
or U6686 (N_6686,N_5250,N_4287);
nand U6687 (N_6687,N_5810,N_5807);
nand U6688 (N_6688,N_5282,N_5711);
nand U6689 (N_6689,N_4350,N_4908);
xnor U6690 (N_6690,N_4602,N_5218);
nand U6691 (N_6691,N_4823,N_4940);
or U6692 (N_6692,N_4160,N_5371);
or U6693 (N_6693,N_5831,N_5094);
xor U6694 (N_6694,N_5666,N_4512);
xnor U6695 (N_6695,N_5877,N_5901);
and U6696 (N_6696,N_5272,N_5582);
nand U6697 (N_6697,N_5269,N_5430);
nand U6698 (N_6698,N_4058,N_4967);
xnor U6699 (N_6699,N_4102,N_5519);
or U6700 (N_6700,N_5593,N_4334);
nand U6701 (N_6701,N_5731,N_4659);
nand U6702 (N_6702,N_4326,N_5521);
nand U6703 (N_6703,N_4828,N_5288);
xor U6704 (N_6704,N_5763,N_5985);
and U6705 (N_6705,N_5418,N_5479);
xnor U6706 (N_6706,N_5144,N_4359);
nor U6707 (N_6707,N_5899,N_5372);
nor U6708 (N_6708,N_5551,N_4882);
nor U6709 (N_6709,N_4036,N_5967);
xnor U6710 (N_6710,N_5900,N_5116);
nand U6711 (N_6711,N_5595,N_5743);
or U6712 (N_6712,N_4769,N_4156);
nor U6713 (N_6713,N_5919,N_4038);
or U6714 (N_6714,N_4481,N_5389);
xnor U6715 (N_6715,N_4786,N_4454);
nand U6716 (N_6716,N_5784,N_5482);
or U6717 (N_6717,N_4229,N_4469);
xor U6718 (N_6718,N_5032,N_5894);
xor U6719 (N_6719,N_4947,N_5303);
or U6720 (N_6720,N_5680,N_4267);
nand U6721 (N_6721,N_5155,N_4261);
or U6722 (N_6722,N_5493,N_5717);
and U6723 (N_6723,N_5386,N_4929);
nor U6724 (N_6724,N_4626,N_4897);
nor U6725 (N_6725,N_5869,N_5662);
or U6726 (N_6726,N_4577,N_5561);
nor U6727 (N_6727,N_5616,N_4524);
nor U6728 (N_6728,N_5903,N_4899);
and U6729 (N_6729,N_5780,N_4398);
xor U6730 (N_6730,N_5547,N_4354);
or U6731 (N_6731,N_4460,N_4519);
and U6732 (N_6732,N_5090,N_4718);
nand U6733 (N_6733,N_5080,N_5455);
nand U6734 (N_6734,N_4872,N_5715);
nand U6735 (N_6735,N_5721,N_5499);
and U6736 (N_6736,N_5480,N_4813);
or U6737 (N_6737,N_4594,N_5015);
xor U6738 (N_6738,N_5507,N_5002);
and U6739 (N_6739,N_5260,N_4110);
xnor U6740 (N_6740,N_4288,N_5130);
nand U6741 (N_6741,N_5127,N_4115);
nand U6742 (N_6742,N_4937,N_5611);
nor U6743 (N_6743,N_4315,N_4846);
nand U6744 (N_6744,N_5732,N_4569);
and U6745 (N_6745,N_4806,N_4489);
nand U6746 (N_6746,N_5963,N_5658);
or U6747 (N_6747,N_4193,N_4963);
or U6748 (N_6748,N_4646,N_4373);
nand U6749 (N_6749,N_5533,N_5655);
and U6750 (N_6750,N_4764,N_4374);
or U6751 (N_6751,N_5366,N_4015);
nand U6752 (N_6752,N_5106,N_4574);
and U6753 (N_6753,N_4832,N_5228);
nor U6754 (N_6754,N_5562,N_4612);
nand U6755 (N_6755,N_5627,N_5411);
or U6756 (N_6756,N_5275,N_4274);
or U6757 (N_6757,N_4103,N_4428);
and U6758 (N_6758,N_4809,N_4976);
nand U6759 (N_6759,N_5779,N_5245);
and U6760 (N_6760,N_5427,N_5384);
xnor U6761 (N_6761,N_5783,N_4285);
xnor U6762 (N_6762,N_4316,N_5587);
nor U6763 (N_6763,N_4966,N_5750);
and U6764 (N_6764,N_5462,N_4466);
or U6765 (N_6765,N_5141,N_5556);
xnor U6766 (N_6766,N_5741,N_4037);
nand U6767 (N_6767,N_4960,N_4139);
and U6768 (N_6768,N_5539,N_4444);
nor U6769 (N_6769,N_4970,N_4029);
and U6770 (N_6770,N_5708,N_4717);
nand U6771 (N_6771,N_4713,N_4016);
xor U6772 (N_6772,N_5013,N_5053);
and U6773 (N_6773,N_5165,N_5081);
or U6774 (N_6774,N_5120,N_5818);
nor U6775 (N_6775,N_4547,N_5572);
and U6776 (N_6776,N_4663,N_4446);
or U6777 (N_6777,N_4842,N_5907);
or U6778 (N_6778,N_5705,N_4284);
or U6779 (N_6779,N_5054,N_5809);
nor U6780 (N_6780,N_5294,N_4624);
nor U6781 (N_6781,N_4635,N_5239);
or U6782 (N_6782,N_4734,N_4534);
nand U6783 (N_6783,N_4483,N_4001);
and U6784 (N_6784,N_5670,N_5577);
nand U6785 (N_6785,N_5424,N_5906);
and U6786 (N_6786,N_4306,N_4461);
nor U6787 (N_6787,N_4561,N_4991);
nand U6788 (N_6788,N_4200,N_4948);
nand U6789 (N_6789,N_4833,N_5636);
xnor U6790 (N_6790,N_4150,N_5580);
or U6791 (N_6791,N_5112,N_4250);
xor U6792 (N_6792,N_4639,N_5498);
xor U6793 (N_6793,N_5915,N_5814);
nor U6794 (N_6794,N_5735,N_4244);
nand U6795 (N_6795,N_4556,N_4154);
nor U6796 (N_6796,N_5579,N_5362);
or U6797 (N_6797,N_4333,N_4170);
xor U6798 (N_6798,N_4370,N_4715);
or U6799 (N_6799,N_5016,N_5514);
and U6800 (N_6800,N_4182,N_5761);
xnor U6801 (N_6801,N_4221,N_4687);
nand U6802 (N_6802,N_4625,N_4062);
nand U6803 (N_6803,N_4632,N_4129);
xor U6804 (N_6804,N_4278,N_4196);
nand U6805 (N_6805,N_4152,N_4808);
nand U6806 (N_6806,N_5143,N_4292);
or U6807 (N_6807,N_4030,N_5206);
nor U6808 (N_6808,N_4898,N_5908);
xnor U6809 (N_6809,N_5381,N_5050);
xnor U6810 (N_6810,N_4737,N_5674);
nor U6811 (N_6811,N_4011,N_5871);
and U6812 (N_6812,N_5537,N_5684);
or U6813 (N_6813,N_5342,N_5210);
xor U6814 (N_6814,N_5766,N_5030);
nand U6815 (N_6815,N_4525,N_4692);
nand U6816 (N_6816,N_5060,N_4310);
or U6817 (N_6817,N_4751,N_4901);
nor U6818 (N_6818,N_5287,N_4399);
xnor U6819 (N_6819,N_4888,N_4071);
nor U6820 (N_6820,N_4245,N_4559);
and U6821 (N_6821,N_4678,N_5451);
and U6822 (N_6822,N_5284,N_4973);
or U6823 (N_6823,N_4796,N_5062);
and U6824 (N_6824,N_5621,N_5681);
xor U6825 (N_6825,N_4412,N_4276);
nor U6826 (N_6826,N_4971,N_4219);
xor U6827 (N_6827,N_5849,N_5162);
or U6828 (N_6828,N_5240,N_5281);
or U6829 (N_6829,N_5797,N_4941);
or U6830 (N_6830,N_5009,N_4847);
nand U6831 (N_6831,N_5573,N_4441);
xnor U6832 (N_6832,N_4668,N_4180);
nor U6833 (N_6833,N_5276,N_4056);
and U6834 (N_6834,N_5775,N_5569);
and U6835 (N_6835,N_4194,N_4669);
or U6836 (N_6836,N_4422,N_5199);
and U6837 (N_6837,N_5859,N_5108);
nand U6838 (N_6838,N_4701,N_4451);
and U6839 (N_6839,N_4579,N_5540);
nor U6840 (N_6840,N_4249,N_4259);
nor U6841 (N_6841,N_4517,N_4599);
xor U6842 (N_6842,N_5891,N_5712);
nand U6843 (N_6843,N_5286,N_4787);
xor U6844 (N_6844,N_5656,N_5308);
and U6845 (N_6845,N_4726,N_5560);
xor U6846 (N_6846,N_4176,N_4790);
and U6847 (N_6847,N_5131,N_5217);
xor U6848 (N_6848,N_5022,N_5668);
xor U6849 (N_6849,N_4345,N_5525);
xnor U6850 (N_6850,N_4330,N_4366);
and U6851 (N_6851,N_5974,N_5170);
and U6852 (N_6852,N_4957,N_5506);
nand U6853 (N_6853,N_5447,N_5309);
xor U6854 (N_6854,N_5134,N_5937);
xor U6855 (N_6855,N_5926,N_4818);
and U6856 (N_6856,N_5653,N_4778);
and U6857 (N_6857,N_4837,N_5745);
nor U6858 (N_6858,N_4113,N_4418);
nor U6859 (N_6859,N_5794,N_5369);
nor U6860 (N_6860,N_5789,N_4591);
xor U6861 (N_6861,N_5632,N_4223);
or U6862 (N_6862,N_4433,N_5639);
nor U6863 (N_6863,N_5801,N_4148);
xor U6864 (N_6864,N_5313,N_4319);
and U6865 (N_6865,N_5755,N_5966);
and U6866 (N_6866,N_4471,N_4184);
xor U6867 (N_6867,N_5110,N_5947);
xnor U6868 (N_6868,N_4010,N_5628);
or U6869 (N_6869,N_5278,N_5538);
and U6870 (N_6870,N_4964,N_4689);
nand U6871 (N_6871,N_5129,N_4925);
xor U6872 (N_6872,N_4853,N_4175);
nand U6873 (N_6873,N_5823,N_5161);
nand U6874 (N_6874,N_5380,N_4526);
or U6875 (N_6875,N_4516,N_4450);
or U6876 (N_6876,N_5028,N_4945);
xor U6877 (N_6877,N_5359,N_4953);
xor U6878 (N_6878,N_4623,N_4098);
and U6879 (N_6879,N_4990,N_4270);
nand U6880 (N_6880,N_5986,N_5492);
nand U6881 (N_6881,N_5837,N_5364);
nand U6882 (N_6882,N_4403,N_5119);
or U6883 (N_6883,N_4927,N_4308);
nand U6884 (N_6884,N_5259,N_4522);
xor U6885 (N_6885,N_5725,N_4562);
xor U6886 (N_6886,N_5555,N_4277);
xor U6887 (N_6887,N_4709,N_4248);
nor U6888 (N_6888,N_5000,N_5363);
nand U6889 (N_6889,N_5336,N_5318);
xor U6890 (N_6890,N_4028,N_4472);
and U6891 (N_6891,N_4174,N_4862);
xor U6892 (N_6892,N_4158,N_4260);
xnor U6893 (N_6893,N_4414,N_4291);
and U6894 (N_6894,N_4567,N_5459);
nand U6895 (N_6895,N_5672,N_4910);
nor U6896 (N_6896,N_5707,N_4587);
xor U6897 (N_6897,N_5512,N_4207);
nand U6898 (N_6898,N_4770,N_5058);
nand U6899 (N_6899,N_5751,N_4008);
xor U6900 (N_6900,N_4903,N_5607);
nor U6901 (N_6901,N_5597,N_5671);
or U6902 (N_6902,N_5153,N_4621);
nand U6903 (N_6903,N_4252,N_5470);
xor U6904 (N_6904,N_5151,N_4338);
nor U6905 (N_6905,N_4309,N_4271);
xor U6906 (N_6906,N_5023,N_4732);
and U6907 (N_6907,N_4336,N_4069);
nand U6908 (N_6908,N_4895,N_5332);
nand U6909 (N_6909,N_5330,N_5552);
xnor U6910 (N_6910,N_5728,N_4297);
nand U6911 (N_6911,N_5230,N_5311);
xnor U6912 (N_6912,N_4064,N_5202);
and U6913 (N_6913,N_4224,N_4703);
or U6914 (N_6914,N_5370,N_4400);
and U6915 (N_6915,N_4074,N_5716);
nor U6916 (N_6916,N_4531,N_5953);
xor U6917 (N_6917,N_4738,N_4484);
xnor U6918 (N_6918,N_4736,N_5651);
nand U6919 (N_6919,N_5257,N_4649);
nor U6920 (N_6920,N_5301,N_5071);
xor U6921 (N_6921,N_5033,N_4445);
or U6922 (N_6922,N_4644,N_4263);
nor U6923 (N_6923,N_4871,N_4875);
nand U6924 (N_6924,N_5403,N_4523);
and U6925 (N_6925,N_5960,N_4985);
nor U6926 (N_6926,N_5101,N_5274);
or U6927 (N_6927,N_4328,N_4452);
nand U6928 (N_6928,N_5008,N_4705);
and U6929 (N_6929,N_5484,N_4946);
nor U6930 (N_6930,N_4151,N_5690);
and U6931 (N_6931,N_5166,N_5069);
or U6932 (N_6932,N_5179,N_4141);
and U6933 (N_6933,N_5461,N_5702);
xnor U6934 (N_6934,N_5703,N_4754);
xnor U6935 (N_6935,N_4138,N_4844);
and U6936 (N_6936,N_4108,N_4500);
nor U6937 (N_6937,N_4977,N_5998);
or U6938 (N_6938,N_5429,N_4295);
nor U6939 (N_6939,N_5685,N_4375);
nor U6940 (N_6940,N_4320,N_5699);
xor U6941 (N_6941,N_5476,N_5663);
xnor U6942 (N_6942,N_5739,N_5099);
xor U6943 (N_6943,N_4670,N_5541);
and U6944 (N_6944,N_5785,N_4654);
nor U6945 (N_6945,N_5337,N_4380);
or U6946 (N_6946,N_4080,N_4693);
nand U6947 (N_6947,N_5300,N_4926);
nor U6948 (N_6948,N_5067,N_5398);
xnor U6949 (N_6949,N_4864,N_5928);
nor U6950 (N_6950,N_4805,N_5890);
xor U6951 (N_6951,N_4708,N_4155);
xor U6952 (N_6952,N_5216,N_4608);
xor U6953 (N_6953,N_4035,N_4865);
or U6954 (N_6954,N_5601,N_5001);
nand U6955 (N_6955,N_4749,N_4704);
xnor U6956 (N_6956,N_5834,N_4118);
and U6957 (N_6957,N_5248,N_5471);
xnor U6958 (N_6958,N_4425,N_5192);
nor U6959 (N_6959,N_4044,N_4436);
and U6960 (N_6960,N_5603,N_4756);
nor U6961 (N_6961,N_4918,N_4592);
nor U6962 (N_6962,N_5643,N_5181);
and U6963 (N_6963,N_4099,N_4090);
nand U6964 (N_6964,N_4022,N_5951);
or U6965 (N_6965,N_4740,N_5532);
and U6966 (N_6966,N_5440,N_5039);
and U6967 (N_6967,N_4401,N_4377);
and U6968 (N_6968,N_5864,N_5629);
or U6969 (N_6969,N_4857,N_5686);
xor U6970 (N_6970,N_5522,N_5952);
and U6971 (N_6971,N_5943,N_5689);
and U6972 (N_6972,N_5078,N_5238);
nand U6973 (N_6973,N_5188,N_5964);
and U6974 (N_6974,N_5222,N_5704);
and U6975 (N_6975,N_4465,N_5791);
and U6976 (N_6976,N_5586,N_5756);
xnor U6977 (N_6977,N_4582,N_5083);
nand U6978 (N_6978,N_4247,N_4464);
nand U6979 (N_6979,N_5346,N_4936);
or U6980 (N_6980,N_4699,N_5853);
and U6981 (N_6981,N_5933,N_4411);
and U6982 (N_6982,N_4431,N_4092);
and U6983 (N_6983,N_5449,N_5234);
and U6984 (N_6984,N_4043,N_5186);
xor U6985 (N_6985,N_4557,N_5962);
nand U6986 (N_6986,N_4696,N_5468);
xor U6987 (N_6987,N_5004,N_5895);
nor U6988 (N_6988,N_5688,N_4822);
nand U6989 (N_6989,N_5184,N_4573);
xor U6990 (N_6990,N_4112,N_5730);
nor U6991 (N_6991,N_4449,N_5650);
nand U6992 (N_6992,N_4911,N_5543);
nor U6993 (N_6993,N_5799,N_4147);
or U6994 (N_6994,N_5983,N_4021);
nor U6995 (N_6995,N_5517,N_5862);
nor U6996 (N_6996,N_4777,N_4631);
nor U6997 (N_6997,N_5174,N_4604);
or U6998 (N_6998,N_5954,N_4817);
or U6999 (N_6999,N_5481,N_4213);
xor U7000 (N_7000,N_4740,N_5307);
nor U7001 (N_7001,N_4995,N_5436);
nor U7002 (N_7002,N_5310,N_4706);
nand U7003 (N_7003,N_4380,N_4265);
or U7004 (N_7004,N_4400,N_5333);
or U7005 (N_7005,N_5982,N_5058);
nor U7006 (N_7006,N_5016,N_5702);
nand U7007 (N_7007,N_4183,N_4672);
or U7008 (N_7008,N_5264,N_4287);
and U7009 (N_7009,N_4045,N_5883);
xor U7010 (N_7010,N_5552,N_5804);
xnor U7011 (N_7011,N_4737,N_4924);
and U7012 (N_7012,N_4062,N_4758);
nor U7013 (N_7013,N_4685,N_5020);
xor U7014 (N_7014,N_5040,N_4984);
or U7015 (N_7015,N_5084,N_4074);
nand U7016 (N_7016,N_4234,N_4995);
nor U7017 (N_7017,N_5879,N_4632);
xor U7018 (N_7018,N_5649,N_5405);
and U7019 (N_7019,N_4580,N_5764);
xnor U7020 (N_7020,N_5396,N_4872);
and U7021 (N_7021,N_5317,N_4355);
nand U7022 (N_7022,N_4325,N_5738);
and U7023 (N_7023,N_5586,N_4134);
nor U7024 (N_7024,N_5998,N_5461);
nor U7025 (N_7025,N_4117,N_5627);
nor U7026 (N_7026,N_5810,N_4886);
nor U7027 (N_7027,N_4518,N_4262);
or U7028 (N_7028,N_5509,N_5443);
or U7029 (N_7029,N_4169,N_5377);
xor U7030 (N_7030,N_5980,N_4363);
nor U7031 (N_7031,N_5558,N_4972);
nor U7032 (N_7032,N_4761,N_4750);
nor U7033 (N_7033,N_4161,N_5504);
and U7034 (N_7034,N_4769,N_4757);
nand U7035 (N_7035,N_4220,N_5466);
or U7036 (N_7036,N_4421,N_4466);
nor U7037 (N_7037,N_5074,N_4870);
nor U7038 (N_7038,N_4891,N_5156);
or U7039 (N_7039,N_5889,N_5148);
nor U7040 (N_7040,N_4318,N_5819);
and U7041 (N_7041,N_4641,N_5354);
and U7042 (N_7042,N_5930,N_4941);
and U7043 (N_7043,N_4494,N_4163);
nand U7044 (N_7044,N_5741,N_5459);
xnor U7045 (N_7045,N_4355,N_5624);
nand U7046 (N_7046,N_4523,N_5098);
nor U7047 (N_7047,N_5222,N_4492);
or U7048 (N_7048,N_5210,N_5341);
and U7049 (N_7049,N_5606,N_5764);
or U7050 (N_7050,N_5089,N_5205);
and U7051 (N_7051,N_5680,N_5700);
and U7052 (N_7052,N_5738,N_5251);
nand U7053 (N_7053,N_5092,N_4821);
xnor U7054 (N_7054,N_4497,N_4340);
nand U7055 (N_7055,N_5703,N_4400);
or U7056 (N_7056,N_5106,N_5138);
nand U7057 (N_7057,N_5471,N_5453);
xor U7058 (N_7058,N_5921,N_5161);
xor U7059 (N_7059,N_4534,N_5677);
nand U7060 (N_7060,N_4221,N_5004);
and U7061 (N_7061,N_4129,N_4607);
or U7062 (N_7062,N_5422,N_4324);
nand U7063 (N_7063,N_4644,N_4533);
nor U7064 (N_7064,N_5477,N_4045);
xnor U7065 (N_7065,N_5737,N_5744);
nor U7066 (N_7066,N_4001,N_4856);
and U7067 (N_7067,N_5636,N_5870);
nand U7068 (N_7068,N_5780,N_5514);
nand U7069 (N_7069,N_4470,N_5028);
or U7070 (N_7070,N_4263,N_5207);
nor U7071 (N_7071,N_5013,N_5078);
nor U7072 (N_7072,N_4668,N_4804);
or U7073 (N_7073,N_5598,N_4887);
nor U7074 (N_7074,N_5857,N_5781);
nand U7075 (N_7075,N_5542,N_4661);
nand U7076 (N_7076,N_5090,N_4473);
xnor U7077 (N_7077,N_5885,N_4124);
and U7078 (N_7078,N_5071,N_4586);
xor U7079 (N_7079,N_5767,N_4340);
and U7080 (N_7080,N_4346,N_4893);
xnor U7081 (N_7081,N_5380,N_4862);
nor U7082 (N_7082,N_4060,N_5011);
and U7083 (N_7083,N_4399,N_5096);
xnor U7084 (N_7084,N_5343,N_4510);
nand U7085 (N_7085,N_4700,N_4092);
xor U7086 (N_7086,N_5052,N_5748);
nor U7087 (N_7087,N_5819,N_5576);
and U7088 (N_7088,N_4626,N_4002);
nand U7089 (N_7089,N_4449,N_4406);
or U7090 (N_7090,N_5558,N_4455);
nand U7091 (N_7091,N_5221,N_5404);
or U7092 (N_7092,N_4830,N_5099);
or U7093 (N_7093,N_4171,N_4545);
xnor U7094 (N_7094,N_4583,N_4281);
or U7095 (N_7095,N_4319,N_4732);
or U7096 (N_7096,N_5642,N_4672);
nor U7097 (N_7097,N_4157,N_5000);
and U7098 (N_7098,N_5805,N_5059);
and U7099 (N_7099,N_4054,N_4806);
nor U7100 (N_7100,N_5840,N_4716);
and U7101 (N_7101,N_5537,N_5787);
nor U7102 (N_7102,N_5289,N_4299);
xnor U7103 (N_7103,N_5948,N_4565);
or U7104 (N_7104,N_5099,N_5175);
xnor U7105 (N_7105,N_4079,N_4618);
and U7106 (N_7106,N_4362,N_4520);
or U7107 (N_7107,N_5149,N_5007);
xnor U7108 (N_7108,N_4856,N_4836);
xnor U7109 (N_7109,N_5356,N_5541);
xor U7110 (N_7110,N_5753,N_5581);
and U7111 (N_7111,N_4864,N_5966);
or U7112 (N_7112,N_4902,N_5782);
nand U7113 (N_7113,N_5314,N_5025);
nor U7114 (N_7114,N_5263,N_4782);
and U7115 (N_7115,N_5782,N_5369);
nor U7116 (N_7116,N_5583,N_4773);
or U7117 (N_7117,N_4846,N_4677);
or U7118 (N_7118,N_5186,N_5440);
xnor U7119 (N_7119,N_5069,N_4918);
xor U7120 (N_7120,N_5216,N_5228);
nand U7121 (N_7121,N_4862,N_5886);
nor U7122 (N_7122,N_4974,N_5027);
xor U7123 (N_7123,N_5363,N_5161);
nand U7124 (N_7124,N_4299,N_5529);
xnor U7125 (N_7125,N_4408,N_5549);
nand U7126 (N_7126,N_4982,N_4612);
and U7127 (N_7127,N_4811,N_5728);
nand U7128 (N_7128,N_4341,N_5188);
xnor U7129 (N_7129,N_5540,N_5821);
xnor U7130 (N_7130,N_5426,N_4356);
xor U7131 (N_7131,N_5066,N_5016);
nor U7132 (N_7132,N_5533,N_4507);
xnor U7133 (N_7133,N_4388,N_5054);
nand U7134 (N_7134,N_5831,N_5157);
and U7135 (N_7135,N_5829,N_4459);
nand U7136 (N_7136,N_5900,N_4054);
nand U7137 (N_7137,N_4912,N_4489);
xor U7138 (N_7138,N_5795,N_5828);
nand U7139 (N_7139,N_5084,N_5605);
nor U7140 (N_7140,N_5081,N_4826);
nand U7141 (N_7141,N_5528,N_5320);
or U7142 (N_7142,N_4805,N_4270);
nand U7143 (N_7143,N_5345,N_5798);
or U7144 (N_7144,N_5535,N_4479);
or U7145 (N_7145,N_4259,N_5323);
and U7146 (N_7146,N_5142,N_5943);
xnor U7147 (N_7147,N_4600,N_5957);
nor U7148 (N_7148,N_5086,N_4833);
or U7149 (N_7149,N_4097,N_5269);
nor U7150 (N_7150,N_4508,N_5270);
nor U7151 (N_7151,N_4346,N_4293);
nor U7152 (N_7152,N_4299,N_4906);
xor U7153 (N_7153,N_5209,N_5199);
xnor U7154 (N_7154,N_5245,N_4539);
and U7155 (N_7155,N_5965,N_5047);
and U7156 (N_7156,N_4771,N_4463);
xor U7157 (N_7157,N_5241,N_5205);
nor U7158 (N_7158,N_5623,N_4796);
and U7159 (N_7159,N_4076,N_5376);
or U7160 (N_7160,N_5794,N_5212);
or U7161 (N_7161,N_4783,N_5740);
nand U7162 (N_7162,N_5532,N_4185);
xor U7163 (N_7163,N_4393,N_5830);
xnor U7164 (N_7164,N_5037,N_4930);
xor U7165 (N_7165,N_5298,N_4643);
nor U7166 (N_7166,N_4340,N_5938);
nand U7167 (N_7167,N_5231,N_4973);
or U7168 (N_7168,N_5339,N_5743);
nor U7169 (N_7169,N_5544,N_4777);
and U7170 (N_7170,N_5337,N_5965);
nor U7171 (N_7171,N_4737,N_4970);
nand U7172 (N_7172,N_4905,N_4215);
and U7173 (N_7173,N_5263,N_4241);
nand U7174 (N_7174,N_4862,N_5971);
nor U7175 (N_7175,N_4924,N_5239);
xor U7176 (N_7176,N_4982,N_4853);
and U7177 (N_7177,N_5035,N_4819);
xor U7178 (N_7178,N_4019,N_4794);
and U7179 (N_7179,N_5118,N_4228);
and U7180 (N_7180,N_5703,N_5576);
nor U7181 (N_7181,N_4458,N_5888);
or U7182 (N_7182,N_5326,N_5032);
nand U7183 (N_7183,N_5460,N_5602);
xor U7184 (N_7184,N_4710,N_5323);
and U7185 (N_7185,N_5861,N_4893);
or U7186 (N_7186,N_4986,N_4785);
or U7187 (N_7187,N_5643,N_5317);
and U7188 (N_7188,N_5139,N_5393);
nor U7189 (N_7189,N_5846,N_5621);
xnor U7190 (N_7190,N_5989,N_5096);
nor U7191 (N_7191,N_4324,N_4420);
or U7192 (N_7192,N_5250,N_5326);
xor U7193 (N_7193,N_5624,N_4964);
xor U7194 (N_7194,N_5189,N_4044);
nor U7195 (N_7195,N_5715,N_4991);
xor U7196 (N_7196,N_4305,N_5626);
xor U7197 (N_7197,N_5867,N_4051);
and U7198 (N_7198,N_5268,N_4985);
xnor U7199 (N_7199,N_4800,N_5467);
nor U7200 (N_7200,N_5914,N_5377);
xor U7201 (N_7201,N_4439,N_4432);
and U7202 (N_7202,N_5173,N_5656);
or U7203 (N_7203,N_4869,N_5072);
and U7204 (N_7204,N_4481,N_4579);
nor U7205 (N_7205,N_4660,N_5518);
nand U7206 (N_7206,N_5254,N_4969);
xor U7207 (N_7207,N_4070,N_4453);
nor U7208 (N_7208,N_5009,N_5375);
and U7209 (N_7209,N_4875,N_4822);
xor U7210 (N_7210,N_5604,N_4949);
nor U7211 (N_7211,N_4621,N_4580);
nor U7212 (N_7212,N_4627,N_5880);
or U7213 (N_7213,N_4314,N_4693);
and U7214 (N_7214,N_4067,N_5091);
nor U7215 (N_7215,N_4418,N_5933);
and U7216 (N_7216,N_4771,N_4975);
and U7217 (N_7217,N_4231,N_4945);
and U7218 (N_7218,N_5491,N_5091);
or U7219 (N_7219,N_5093,N_5491);
nor U7220 (N_7220,N_4229,N_5042);
nor U7221 (N_7221,N_4843,N_4331);
nor U7222 (N_7222,N_4312,N_4040);
nand U7223 (N_7223,N_5777,N_5197);
and U7224 (N_7224,N_4445,N_4859);
and U7225 (N_7225,N_4080,N_4167);
and U7226 (N_7226,N_4994,N_4974);
nand U7227 (N_7227,N_4171,N_4054);
or U7228 (N_7228,N_5973,N_5757);
nand U7229 (N_7229,N_4751,N_4608);
nor U7230 (N_7230,N_5042,N_5453);
or U7231 (N_7231,N_4582,N_4055);
and U7232 (N_7232,N_4710,N_4567);
or U7233 (N_7233,N_5151,N_4691);
nand U7234 (N_7234,N_4375,N_4247);
nor U7235 (N_7235,N_4539,N_5482);
or U7236 (N_7236,N_4235,N_5557);
or U7237 (N_7237,N_4299,N_5833);
xor U7238 (N_7238,N_4773,N_5031);
nand U7239 (N_7239,N_4501,N_5382);
xor U7240 (N_7240,N_4917,N_5664);
nor U7241 (N_7241,N_5506,N_4429);
and U7242 (N_7242,N_5958,N_5774);
nor U7243 (N_7243,N_5035,N_5085);
xor U7244 (N_7244,N_5167,N_4370);
nand U7245 (N_7245,N_5611,N_4223);
nor U7246 (N_7246,N_4987,N_4407);
nor U7247 (N_7247,N_4960,N_5596);
or U7248 (N_7248,N_5821,N_5827);
nand U7249 (N_7249,N_5193,N_5811);
and U7250 (N_7250,N_4452,N_4220);
nand U7251 (N_7251,N_4776,N_5994);
nor U7252 (N_7252,N_4587,N_5227);
and U7253 (N_7253,N_4542,N_4232);
and U7254 (N_7254,N_5560,N_5646);
and U7255 (N_7255,N_4084,N_5986);
xnor U7256 (N_7256,N_5503,N_5347);
or U7257 (N_7257,N_5083,N_4062);
nand U7258 (N_7258,N_5476,N_4474);
or U7259 (N_7259,N_5130,N_4902);
or U7260 (N_7260,N_5796,N_4728);
and U7261 (N_7261,N_4444,N_4171);
nor U7262 (N_7262,N_4611,N_5087);
xnor U7263 (N_7263,N_5423,N_5502);
nand U7264 (N_7264,N_5312,N_4332);
and U7265 (N_7265,N_5120,N_4588);
nor U7266 (N_7266,N_5052,N_4623);
and U7267 (N_7267,N_5268,N_5816);
nand U7268 (N_7268,N_5174,N_4223);
xnor U7269 (N_7269,N_5766,N_5599);
nor U7270 (N_7270,N_5711,N_4936);
and U7271 (N_7271,N_5004,N_5821);
nand U7272 (N_7272,N_4626,N_4770);
xnor U7273 (N_7273,N_4880,N_4495);
nor U7274 (N_7274,N_5113,N_4703);
or U7275 (N_7275,N_4834,N_4035);
nand U7276 (N_7276,N_4035,N_4097);
nand U7277 (N_7277,N_5928,N_5972);
nor U7278 (N_7278,N_4313,N_5078);
nor U7279 (N_7279,N_5512,N_4525);
nand U7280 (N_7280,N_4116,N_5938);
or U7281 (N_7281,N_5291,N_4330);
xnor U7282 (N_7282,N_5402,N_5403);
nand U7283 (N_7283,N_4043,N_4242);
nand U7284 (N_7284,N_5785,N_4681);
nor U7285 (N_7285,N_4199,N_4610);
nand U7286 (N_7286,N_5979,N_4554);
and U7287 (N_7287,N_4822,N_5054);
nand U7288 (N_7288,N_4836,N_4226);
nor U7289 (N_7289,N_4385,N_5184);
nand U7290 (N_7290,N_4303,N_4476);
or U7291 (N_7291,N_5372,N_5832);
nor U7292 (N_7292,N_5833,N_5950);
and U7293 (N_7293,N_4765,N_4201);
nor U7294 (N_7294,N_4684,N_5427);
and U7295 (N_7295,N_5061,N_5265);
xor U7296 (N_7296,N_4036,N_5056);
xnor U7297 (N_7297,N_4557,N_5558);
nor U7298 (N_7298,N_4843,N_4391);
nand U7299 (N_7299,N_5226,N_4728);
nor U7300 (N_7300,N_5497,N_4012);
or U7301 (N_7301,N_5061,N_4884);
xor U7302 (N_7302,N_5133,N_5754);
nand U7303 (N_7303,N_5941,N_5284);
xor U7304 (N_7304,N_5503,N_4961);
and U7305 (N_7305,N_4301,N_5339);
xnor U7306 (N_7306,N_4365,N_4325);
nand U7307 (N_7307,N_4608,N_4332);
nor U7308 (N_7308,N_5265,N_5218);
nor U7309 (N_7309,N_4584,N_4590);
or U7310 (N_7310,N_5979,N_4959);
nor U7311 (N_7311,N_4068,N_4243);
nor U7312 (N_7312,N_4159,N_5693);
nor U7313 (N_7313,N_5127,N_5597);
and U7314 (N_7314,N_4928,N_5473);
nor U7315 (N_7315,N_4575,N_4664);
or U7316 (N_7316,N_5326,N_4771);
xor U7317 (N_7317,N_5888,N_5232);
or U7318 (N_7318,N_5178,N_5801);
nand U7319 (N_7319,N_5735,N_4322);
and U7320 (N_7320,N_4122,N_5426);
nor U7321 (N_7321,N_4864,N_5306);
nor U7322 (N_7322,N_5830,N_4865);
nor U7323 (N_7323,N_5090,N_4938);
xnor U7324 (N_7324,N_4284,N_5949);
nor U7325 (N_7325,N_5838,N_5481);
nand U7326 (N_7326,N_4516,N_5579);
nand U7327 (N_7327,N_5275,N_5795);
nand U7328 (N_7328,N_5914,N_5103);
xor U7329 (N_7329,N_4452,N_5339);
or U7330 (N_7330,N_4072,N_5371);
nand U7331 (N_7331,N_4512,N_4526);
nand U7332 (N_7332,N_4714,N_5719);
nor U7333 (N_7333,N_4250,N_5201);
nand U7334 (N_7334,N_4426,N_4786);
and U7335 (N_7335,N_5432,N_4104);
xor U7336 (N_7336,N_5570,N_5949);
and U7337 (N_7337,N_4807,N_5606);
and U7338 (N_7338,N_4784,N_4023);
nand U7339 (N_7339,N_4726,N_5602);
nand U7340 (N_7340,N_5646,N_5605);
nand U7341 (N_7341,N_4026,N_5892);
and U7342 (N_7342,N_5984,N_5346);
nand U7343 (N_7343,N_4202,N_5886);
xor U7344 (N_7344,N_4739,N_5711);
nand U7345 (N_7345,N_4639,N_4927);
nand U7346 (N_7346,N_4288,N_4868);
xor U7347 (N_7347,N_5396,N_5541);
xnor U7348 (N_7348,N_4831,N_5270);
and U7349 (N_7349,N_4140,N_4451);
or U7350 (N_7350,N_5841,N_4731);
and U7351 (N_7351,N_4848,N_4872);
or U7352 (N_7352,N_4611,N_4711);
nand U7353 (N_7353,N_5285,N_5602);
and U7354 (N_7354,N_4415,N_5656);
or U7355 (N_7355,N_4561,N_5910);
and U7356 (N_7356,N_4672,N_5561);
or U7357 (N_7357,N_4707,N_5646);
nor U7358 (N_7358,N_4411,N_5817);
nor U7359 (N_7359,N_5336,N_4447);
nand U7360 (N_7360,N_5399,N_5184);
or U7361 (N_7361,N_5311,N_5022);
xnor U7362 (N_7362,N_5304,N_5068);
or U7363 (N_7363,N_4918,N_4980);
nor U7364 (N_7364,N_5739,N_4035);
and U7365 (N_7365,N_5601,N_5938);
nor U7366 (N_7366,N_4913,N_5596);
nand U7367 (N_7367,N_4865,N_4968);
nand U7368 (N_7368,N_4691,N_5649);
nor U7369 (N_7369,N_4678,N_5488);
nor U7370 (N_7370,N_5710,N_5936);
nor U7371 (N_7371,N_5253,N_5072);
and U7372 (N_7372,N_4362,N_5432);
nor U7373 (N_7373,N_5921,N_4075);
xor U7374 (N_7374,N_4572,N_5905);
and U7375 (N_7375,N_4811,N_5748);
and U7376 (N_7376,N_4624,N_5576);
xor U7377 (N_7377,N_4649,N_5336);
or U7378 (N_7378,N_5983,N_5948);
xnor U7379 (N_7379,N_4393,N_5467);
nand U7380 (N_7380,N_5513,N_5360);
nor U7381 (N_7381,N_4062,N_4675);
xor U7382 (N_7382,N_4964,N_4239);
nor U7383 (N_7383,N_5432,N_4718);
xnor U7384 (N_7384,N_4050,N_4784);
or U7385 (N_7385,N_5054,N_4099);
and U7386 (N_7386,N_5956,N_4390);
nor U7387 (N_7387,N_4406,N_4854);
nand U7388 (N_7388,N_5106,N_5728);
and U7389 (N_7389,N_4266,N_4843);
and U7390 (N_7390,N_5182,N_4603);
xnor U7391 (N_7391,N_4425,N_5646);
xor U7392 (N_7392,N_4553,N_4978);
and U7393 (N_7393,N_4367,N_5020);
and U7394 (N_7394,N_5612,N_4192);
xor U7395 (N_7395,N_5857,N_4280);
xnor U7396 (N_7396,N_5863,N_4569);
xor U7397 (N_7397,N_4421,N_5757);
and U7398 (N_7398,N_5775,N_4495);
and U7399 (N_7399,N_4543,N_5912);
xor U7400 (N_7400,N_4609,N_5854);
nand U7401 (N_7401,N_4898,N_4593);
xor U7402 (N_7402,N_4212,N_5422);
or U7403 (N_7403,N_5658,N_5707);
nor U7404 (N_7404,N_4284,N_4938);
nor U7405 (N_7405,N_5718,N_4849);
xor U7406 (N_7406,N_5580,N_4866);
nor U7407 (N_7407,N_4587,N_5698);
and U7408 (N_7408,N_5103,N_5662);
or U7409 (N_7409,N_5226,N_4044);
and U7410 (N_7410,N_4355,N_5032);
xor U7411 (N_7411,N_5640,N_5324);
and U7412 (N_7412,N_5578,N_4397);
or U7413 (N_7413,N_4046,N_5063);
nand U7414 (N_7414,N_5240,N_4902);
or U7415 (N_7415,N_4809,N_5387);
or U7416 (N_7416,N_4917,N_5827);
and U7417 (N_7417,N_4028,N_5052);
nor U7418 (N_7418,N_5393,N_4096);
nand U7419 (N_7419,N_5910,N_4823);
nor U7420 (N_7420,N_4926,N_4210);
or U7421 (N_7421,N_4916,N_4955);
xor U7422 (N_7422,N_4202,N_5418);
nor U7423 (N_7423,N_5296,N_4847);
and U7424 (N_7424,N_4990,N_4105);
nand U7425 (N_7425,N_4617,N_5996);
nand U7426 (N_7426,N_4258,N_5968);
xor U7427 (N_7427,N_4806,N_5226);
nand U7428 (N_7428,N_5772,N_5846);
nand U7429 (N_7429,N_5022,N_4781);
xnor U7430 (N_7430,N_4072,N_4410);
nor U7431 (N_7431,N_4918,N_4761);
nor U7432 (N_7432,N_4056,N_5360);
and U7433 (N_7433,N_5895,N_4504);
xnor U7434 (N_7434,N_4214,N_4397);
or U7435 (N_7435,N_5085,N_5526);
or U7436 (N_7436,N_5922,N_5234);
nor U7437 (N_7437,N_5521,N_4802);
xor U7438 (N_7438,N_4428,N_4806);
nand U7439 (N_7439,N_4998,N_4867);
nand U7440 (N_7440,N_4907,N_4637);
nor U7441 (N_7441,N_4946,N_4460);
nor U7442 (N_7442,N_4541,N_4901);
xor U7443 (N_7443,N_4138,N_4962);
or U7444 (N_7444,N_5214,N_5369);
nand U7445 (N_7445,N_4777,N_5499);
nor U7446 (N_7446,N_4902,N_5251);
xor U7447 (N_7447,N_4655,N_5708);
nor U7448 (N_7448,N_4690,N_5431);
nand U7449 (N_7449,N_5296,N_4709);
nand U7450 (N_7450,N_4384,N_5256);
or U7451 (N_7451,N_4526,N_5464);
xor U7452 (N_7452,N_4944,N_5976);
nand U7453 (N_7453,N_5169,N_4190);
or U7454 (N_7454,N_5347,N_4989);
or U7455 (N_7455,N_5554,N_4719);
or U7456 (N_7456,N_4813,N_4703);
nand U7457 (N_7457,N_4602,N_4565);
or U7458 (N_7458,N_4648,N_5201);
and U7459 (N_7459,N_5479,N_5294);
xor U7460 (N_7460,N_5740,N_5158);
and U7461 (N_7461,N_4582,N_5439);
nor U7462 (N_7462,N_4335,N_4958);
xnor U7463 (N_7463,N_5442,N_4477);
xnor U7464 (N_7464,N_5782,N_4208);
nand U7465 (N_7465,N_4357,N_5661);
and U7466 (N_7466,N_4750,N_4499);
or U7467 (N_7467,N_5175,N_4220);
nor U7468 (N_7468,N_5570,N_4612);
and U7469 (N_7469,N_4160,N_4514);
xor U7470 (N_7470,N_5872,N_5630);
nand U7471 (N_7471,N_5128,N_5862);
nand U7472 (N_7472,N_4690,N_5907);
or U7473 (N_7473,N_4822,N_5853);
or U7474 (N_7474,N_5411,N_5319);
nand U7475 (N_7475,N_5634,N_4761);
or U7476 (N_7476,N_5035,N_4134);
and U7477 (N_7477,N_4924,N_5119);
nor U7478 (N_7478,N_5104,N_5694);
nand U7479 (N_7479,N_4136,N_4732);
nor U7480 (N_7480,N_4024,N_5497);
nor U7481 (N_7481,N_5790,N_4503);
xnor U7482 (N_7482,N_5430,N_4249);
and U7483 (N_7483,N_5833,N_5569);
xnor U7484 (N_7484,N_4542,N_5485);
or U7485 (N_7485,N_4974,N_4488);
or U7486 (N_7486,N_5275,N_5131);
nand U7487 (N_7487,N_5723,N_4489);
and U7488 (N_7488,N_4089,N_5617);
xor U7489 (N_7489,N_5157,N_4482);
xnor U7490 (N_7490,N_5015,N_5327);
nor U7491 (N_7491,N_5715,N_5377);
or U7492 (N_7492,N_5510,N_4260);
or U7493 (N_7493,N_5353,N_4539);
nor U7494 (N_7494,N_5878,N_5434);
nand U7495 (N_7495,N_5190,N_5698);
nand U7496 (N_7496,N_5624,N_5917);
nand U7497 (N_7497,N_5044,N_4118);
nor U7498 (N_7498,N_4851,N_4149);
nor U7499 (N_7499,N_4687,N_5038);
or U7500 (N_7500,N_4747,N_4053);
nor U7501 (N_7501,N_4237,N_4841);
or U7502 (N_7502,N_5279,N_4949);
or U7503 (N_7503,N_5127,N_5606);
and U7504 (N_7504,N_5236,N_4185);
or U7505 (N_7505,N_4308,N_5311);
and U7506 (N_7506,N_4986,N_4897);
nor U7507 (N_7507,N_5286,N_4516);
and U7508 (N_7508,N_4449,N_5973);
and U7509 (N_7509,N_4741,N_5729);
xnor U7510 (N_7510,N_4062,N_4572);
and U7511 (N_7511,N_5722,N_5661);
xnor U7512 (N_7512,N_4188,N_5626);
xnor U7513 (N_7513,N_4959,N_5485);
nand U7514 (N_7514,N_4096,N_4749);
or U7515 (N_7515,N_5491,N_4199);
nor U7516 (N_7516,N_5885,N_4386);
nand U7517 (N_7517,N_5972,N_4772);
nand U7518 (N_7518,N_5065,N_4893);
xor U7519 (N_7519,N_5132,N_4896);
nor U7520 (N_7520,N_4672,N_4784);
xnor U7521 (N_7521,N_5489,N_5907);
xnor U7522 (N_7522,N_4934,N_5575);
nor U7523 (N_7523,N_5240,N_5241);
or U7524 (N_7524,N_5865,N_5503);
and U7525 (N_7525,N_5512,N_5015);
or U7526 (N_7526,N_5153,N_4339);
nor U7527 (N_7527,N_5066,N_5456);
or U7528 (N_7528,N_4844,N_5541);
nand U7529 (N_7529,N_5916,N_4760);
xnor U7530 (N_7530,N_5684,N_5165);
nor U7531 (N_7531,N_5229,N_5065);
and U7532 (N_7532,N_4114,N_4812);
nand U7533 (N_7533,N_4358,N_4991);
or U7534 (N_7534,N_5820,N_5256);
nand U7535 (N_7535,N_4395,N_4787);
nand U7536 (N_7536,N_5290,N_4132);
xnor U7537 (N_7537,N_5415,N_4288);
or U7538 (N_7538,N_5003,N_5706);
xnor U7539 (N_7539,N_5739,N_5858);
and U7540 (N_7540,N_5888,N_4343);
nand U7541 (N_7541,N_4654,N_5339);
or U7542 (N_7542,N_5842,N_5105);
or U7543 (N_7543,N_4071,N_4656);
nor U7544 (N_7544,N_5256,N_5567);
or U7545 (N_7545,N_5285,N_5104);
xor U7546 (N_7546,N_4030,N_5232);
nor U7547 (N_7547,N_4807,N_4695);
or U7548 (N_7548,N_5238,N_4661);
xor U7549 (N_7549,N_4922,N_4968);
nand U7550 (N_7550,N_5439,N_4013);
or U7551 (N_7551,N_4871,N_5024);
or U7552 (N_7552,N_4627,N_5956);
nor U7553 (N_7553,N_4235,N_4422);
and U7554 (N_7554,N_4328,N_4600);
and U7555 (N_7555,N_5949,N_5696);
nor U7556 (N_7556,N_5914,N_5012);
nor U7557 (N_7557,N_4232,N_5693);
and U7558 (N_7558,N_4846,N_4808);
xnor U7559 (N_7559,N_4663,N_4304);
xnor U7560 (N_7560,N_4213,N_5605);
or U7561 (N_7561,N_5175,N_5503);
nor U7562 (N_7562,N_4094,N_5468);
xor U7563 (N_7563,N_5425,N_5553);
nor U7564 (N_7564,N_5563,N_5867);
xor U7565 (N_7565,N_4344,N_5882);
or U7566 (N_7566,N_4861,N_4319);
xor U7567 (N_7567,N_4039,N_4763);
and U7568 (N_7568,N_4947,N_4908);
and U7569 (N_7569,N_5833,N_4690);
and U7570 (N_7570,N_5348,N_4737);
and U7571 (N_7571,N_4684,N_5675);
nand U7572 (N_7572,N_4857,N_4455);
nand U7573 (N_7573,N_4044,N_5832);
or U7574 (N_7574,N_5161,N_4405);
nand U7575 (N_7575,N_5995,N_4673);
or U7576 (N_7576,N_4187,N_5729);
and U7577 (N_7577,N_4281,N_5279);
and U7578 (N_7578,N_5631,N_5952);
and U7579 (N_7579,N_4709,N_5628);
nor U7580 (N_7580,N_4073,N_4706);
nor U7581 (N_7581,N_5219,N_5870);
and U7582 (N_7582,N_5232,N_4231);
xor U7583 (N_7583,N_4930,N_5116);
or U7584 (N_7584,N_5175,N_5759);
nand U7585 (N_7585,N_5808,N_5902);
nand U7586 (N_7586,N_4930,N_4299);
xnor U7587 (N_7587,N_4181,N_5605);
nand U7588 (N_7588,N_4499,N_5635);
or U7589 (N_7589,N_4085,N_4150);
or U7590 (N_7590,N_4634,N_4410);
or U7591 (N_7591,N_4915,N_5918);
and U7592 (N_7592,N_5520,N_5644);
or U7593 (N_7593,N_4052,N_4337);
nand U7594 (N_7594,N_5248,N_4364);
nand U7595 (N_7595,N_5431,N_4490);
xor U7596 (N_7596,N_5877,N_5418);
xnor U7597 (N_7597,N_4251,N_4822);
and U7598 (N_7598,N_5986,N_4644);
or U7599 (N_7599,N_5223,N_5906);
xor U7600 (N_7600,N_5850,N_4237);
xor U7601 (N_7601,N_4134,N_4845);
xor U7602 (N_7602,N_4186,N_5504);
or U7603 (N_7603,N_4713,N_5119);
and U7604 (N_7604,N_5770,N_5141);
nor U7605 (N_7605,N_4778,N_5874);
nor U7606 (N_7606,N_4438,N_5606);
and U7607 (N_7607,N_5958,N_5269);
xnor U7608 (N_7608,N_5678,N_5281);
nor U7609 (N_7609,N_5963,N_5981);
or U7610 (N_7610,N_4018,N_4360);
or U7611 (N_7611,N_5683,N_4293);
xor U7612 (N_7612,N_5919,N_5647);
and U7613 (N_7613,N_5389,N_5225);
xnor U7614 (N_7614,N_4149,N_4089);
nor U7615 (N_7615,N_5062,N_5886);
nor U7616 (N_7616,N_5153,N_4201);
and U7617 (N_7617,N_5502,N_4283);
or U7618 (N_7618,N_5949,N_4436);
and U7619 (N_7619,N_5538,N_5495);
xnor U7620 (N_7620,N_5373,N_5899);
nor U7621 (N_7621,N_4887,N_4757);
xor U7622 (N_7622,N_5263,N_4894);
nor U7623 (N_7623,N_4362,N_5798);
xor U7624 (N_7624,N_5892,N_4234);
or U7625 (N_7625,N_5088,N_4119);
nor U7626 (N_7626,N_4702,N_4368);
xor U7627 (N_7627,N_5569,N_5425);
or U7628 (N_7628,N_4092,N_5395);
nor U7629 (N_7629,N_5216,N_5920);
xnor U7630 (N_7630,N_5378,N_4883);
and U7631 (N_7631,N_4757,N_4018);
xor U7632 (N_7632,N_4226,N_4269);
xnor U7633 (N_7633,N_4127,N_4599);
nor U7634 (N_7634,N_5937,N_4572);
and U7635 (N_7635,N_4647,N_4323);
nor U7636 (N_7636,N_4675,N_5220);
xor U7637 (N_7637,N_5563,N_5352);
nand U7638 (N_7638,N_5436,N_5901);
or U7639 (N_7639,N_4309,N_4366);
or U7640 (N_7640,N_5849,N_5618);
and U7641 (N_7641,N_5885,N_4072);
and U7642 (N_7642,N_4022,N_5774);
and U7643 (N_7643,N_5813,N_5135);
xnor U7644 (N_7644,N_4440,N_5630);
nand U7645 (N_7645,N_4646,N_4757);
or U7646 (N_7646,N_5446,N_4773);
nor U7647 (N_7647,N_4583,N_5326);
xnor U7648 (N_7648,N_5088,N_4751);
xor U7649 (N_7649,N_5858,N_4335);
nor U7650 (N_7650,N_4575,N_4607);
nand U7651 (N_7651,N_4184,N_5453);
or U7652 (N_7652,N_5068,N_5932);
nand U7653 (N_7653,N_4267,N_4925);
nand U7654 (N_7654,N_4812,N_4579);
nand U7655 (N_7655,N_4358,N_5609);
and U7656 (N_7656,N_5804,N_4952);
xnor U7657 (N_7657,N_5207,N_5576);
xnor U7658 (N_7658,N_5667,N_4050);
or U7659 (N_7659,N_4615,N_5593);
or U7660 (N_7660,N_4322,N_4701);
and U7661 (N_7661,N_4277,N_4397);
xor U7662 (N_7662,N_4035,N_5712);
and U7663 (N_7663,N_4356,N_5784);
xnor U7664 (N_7664,N_4961,N_5005);
nand U7665 (N_7665,N_5522,N_5905);
or U7666 (N_7666,N_5306,N_4043);
and U7667 (N_7667,N_5096,N_5748);
xor U7668 (N_7668,N_5608,N_5627);
or U7669 (N_7669,N_4424,N_4357);
nand U7670 (N_7670,N_4208,N_4620);
nand U7671 (N_7671,N_4541,N_4354);
and U7672 (N_7672,N_5148,N_5717);
nand U7673 (N_7673,N_4386,N_5534);
xor U7674 (N_7674,N_5555,N_5938);
and U7675 (N_7675,N_5625,N_5169);
or U7676 (N_7676,N_4001,N_5123);
xnor U7677 (N_7677,N_4760,N_5765);
nand U7678 (N_7678,N_4428,N_5720);
nand U7679 (N_7679,N_4507,N_4087);
nor U7680 (N_7680,N_4330,N_5288);
nand U7681 (N_7681,N_5266,N_5651);
or U7682 (N_7682,N_5690,N_4191);
nand U7683 (N_7683,N_5320,N_5593);
nor U7684 (N_7684,N_5812,N_4904);
or U7685 (N_7685,N_4294,N_4839);
nor U7686 (N_7686,N_4432,N_5516);
xnor U7687 (N_7687,N_4429,N_5348);
nand U7688 (N_7688,N_5843,N_4606);
nand U7689 (N_7689,N_5791,N_5353);
and U7690 (N_7690,N_5357,N_4330);
or U7691 (N_7691,N_4089,N_5852);
or U7692 (N_7692,N_4973,N_5814);
and U7693 (N_7693,N_5743,N_4234);
nand U7694 (N_7694,N_5645,N_4955);
or U7695 (N_7695,N_4836,N_5618);
xor U7696 (N_7696,N_4359,N_5222);
or U7697 (N_7697,N_4768,N_4160);
or U7698 (N_7698,N_5300,N_4248);
and U7699 (N_7699,N_5579,N_4282);
nand U7700 (N_7700,N_5136,N_5601);
nand U7701 (N_7701,N_5364,N_5988);
or U7702 (N_7702,N_5766,N_4888);
nor U7703 (N_7703,N_4543,N_4302);
nor U7704 (N_7704,N_4612,N_4467);
or U7705 (N_7705,N_5361,N_4019);
or U7706 (N_7706,N_5412,N_5080);
xor U7707 (N_7707,N_4271,N_4872);
or U7708 (N_7708,N_4637,N_5461);
or U7709 (N_7709,N_5190,N_4646);
or U7710 (N_7710,N_4750,N_5029);
nand U7711 (N_7711,N_5232,N_5118);
xor U7712 (N_7712,N_4278,N_4766);
nor U7713 (N_7713,N_4309,N_5221);
and U7714 (N_7714,N_5703,N_4249);
nand U7715 (N_7715,N_5796,N_5578);
and U7716 (N_7716,N_5647,N_4784);
xor U7717 (N_7717,N_4022,N_5070);
xor U7718 (N_7718,N_4585,N_5340);
nor U7719 (N_7719,N_5849,N_5870);
or U7720 (N_7720,N_5507,N_4415);
nand U7721 (N_7721,N_5080,N_4860);
xnor U7722 (N_7722,N_4937,N_5715);
nand U7723 (N_7723,N_5500,N_5950);
and U7724 (N_7724,N_4992,N_5026);
nand U7725 (N_7725,N_5273,N_4587);
nand U7726 (N_7726,N_5121,N_4952);
or U7727 (N_7727,N_4320,N_4728);
or U7728 (N_7728,N_5562,N_5111);
xnor U7729 (N_7729,N_4911,N_5023);
nand U7730 (N_7730,N_5725,N_5013);
or U7731 (N_7731,N_4879,N_4925);
xnor U7732 (N_7732,N_5152,N_4047);
nor U7733 (N_7733,N_5792,N_4461);
and U7734 (N_7734,N_5552,N_5543);
nor U7735 (N_7735,N_4556,N_5102);
nand U7736 (N_7736,N_4584,N_5152);
xor U7737 (N_7737,N_4647,N_5691);
and U7738 (N_7738,N_4720,N_5004);
nand U7739 (N_7739,N_5498,N_5581);
xor U7740 (N_7740,N_4257,N_4785);
or U7741 (N_7741,N_4743,N_4151);
nand U7742 (N_7742,N_4669,N_5141);
xnor U7743 (N_7743,N_5595,N_4470);
or U7744 (N_7744,N_4419,N_5911);
and U7745 (N_7745,N_4853,N_4521);
nand U7746 (N_7746,N_5697,N_5259);
nand U7747 (N_7747,N_4431,N_4159);
nor U7748 (N_7748,N_4146,N_4150);
nand U7749 (N_7749,N_5376,N_4590);
nand U7750 (N_7750,N_5518,N_5666);
nand U7751 (N_7751,N_4021,N_4281);
nor U7752 (N_7752,N_5307,N_4944);
xor U7753 (N_7753,N_4885,N_4210);
and U7754 (N_7754,N_5155,N_5487);
or U7755 (N_7755,N_5318,N_4216);
or U7756 (N_7756,N_5316,N_4700);
xnor U7757 (N_7757,N_4254,N_5691);
and U7758 (N_7758,N_4559,N_4656);
and U7759 (N_7759,N_5395,N_4614);
xnor U7760 (N_7760,N_5006,N_5464);
or U7761 (N_7761,N_4766,N_5820);
and U7762 (N_7762,N_5552,N_4235);
and U7763 (N_7763,N_5004,N_4498);
and U7764 (N_7764,N_4769,N_5487);
xnor U7765 (N_7765,N_5934,N_4930);
nand U7766 (N_7766,N_4462,N_4159);
xnor U7767 (N_7767,N_5710,N_4410);
nor U7768 (N_7768,N_5139,N_5012);
nor U7769 (N_7769,N_5569,N_4206);
and U7770 (N_7770,N_5115,N_5996);
nand U7771 (N_7771,N_4374,N_4600);
or U7772 (N_7772,N_5797,N_5756);
nor U7773 (N_7773,N_4334,N_4717);
nor U7774 (N_7774,N_5235,N_4514);
nand U7775 (N_7775,N_5730,N_5949);
nand U7776 (N_7776,N_5320,N_4226);
and U7777 (N_7777,N_5589,N_4500);
xor U7778 (N_7778,N_5451,N_4736);
nor U7779 (N_7779,N_5533,N_4610);
xor U7780 (N_7780,N_4066,N_4879);
and U7781 (N_7781,N_4961,N_5567);
xor U7782 (N_7782,N_4473,N_4317);
and U7783 (N_7783,N_5459,N_4993);
nor U7784 (N_7784,N_4091,N_5885);
or U7785 (N_7785,N_5518,N_4817);
xor U7786 (N_7786,N_4159,N_4379);
nand U7787 (N_7787,N_5932,N_4933);
or U7788 (N_7788,N_4971,N_4671);
nor U7789 (N_7789,N_5594,N_4105);
nand U7790 (N_7790,N_4955,N_5187);
nand U7791 (N_7791,N_5372,N_5074);
or U7792 (N_7792,N_4123,N_4799);
xor U7793 (N_7793,N_4026,N_5547);
nor U7794 (N_7794,N_4274,N_5233);
xnor U7795 (N_7795,N_5078,N_5207);
and U7796 (N_7796,N_4731,N_5147);
nand U7797 (N_7797,N_5743,N_4762);
nor U7798 (N_7798,N_5734,N_5984);
or U7799 (N_7799,N_4938,N_4570);
xnor U7800 (N_7800,N_4510,N_4832);
nand U7801 (N_7801,N_4515,N_5427);
or U7802 (N_7802,N_4247,N_4520);
nor U7803 (N_7803,N_5133,N_5851);
or U7804 (N_7804,N_5672,N_4851);
and U7805 (N_7805,N_4886,N_4198);
xor U7806 (N_7806,N_5948,N_5898);
xnor U7807 (N_7807,N_4350,N_5430);
or U7808 (N_7808,N_4651,N_5125);
xnor U7809 (N_7809,N_5970,N_5732);
xor U7810 (N_7810,N_4506,N_4309);
and U7811 (N_7811,N_4010,N_4934);
nor U7812 (N_7812,N_4951,N_5652);
nand U7813 (N_7813,N_5346,N_4232);
nand U7814 (N_7814,N_4810,N_4857);
nand U7815 (N_7815,N_5270,N_5333);
nand U7816 (N_7816,N_5266,N_4059);
xnor U7817 (N_7817,N_5595,N_5381);
and U7818 (N_7818,N_4552,N_4514);
nand U7819 (N_7819,N_4096,N_5206);
or U7820 (N_7820,N_4854,N_5711);
nor U7821 (N_7821,N_5455,N_4903);
nor U7822 (N_7822,N_5010,N_5119);
and U7823 (N_7823,N_4333,N_5116);
nor U7824 (N_7824,N_4435,N_4791);
and U7825 (N_7825,N_5476,N_5820);
or U7826 (N_7826,N_4192,N_5572);
nand U7827 (N_7827,N_5223,N_4206);
nand U7828 (N_7828,N_4283,N_5611);
nor U7829 (N_7829,N_5783,N_4914);
nand U7830 (N_7830,N_5277,N_5707);
xnor U7831 (N_7831,N_4356,N_4244);
nor U7832 (N_7832,N_5323,N_5932);
or U7833 (N_7833,N_5533,N_5252);
nand U7834 (N_7834,N_4248,N_5754);
nand U7835 (N_7835,N_5163,N_5029);
nor U7836 (N_7836,N_5067,N_5583);
and U7837 (N_7837,N_4618,N_4533);
nor U7838 (N_7838,N_4274,N_4483);
xor U7839 (N_7839,N_4820,N_5133);
or U7840 (N_7840,N_4231,N_5815);
nor U7841 (N_7841,N_4680,N_4947);
xnor U7842 (N_7842,N_4166,N_5238);
and U7843 (N_7843,N_4312,N_5218);
nand U7844 (N_7844,N_5320,N_4054);
nand U7845 (N_7845,N_4239,N_5983);
nor U7846 (N_7846,N_5151,N_5131);
or U7847 (N_7847,N_5646,N_4849);
nor U7848 (N_7848,N_4169,N_4279);
nor U7849 (N_7849,N_4049,N_4945);
xnor U7850 (N_7850,N_5090,N_4227);
or U7851 (N_7851,N_4980,N_4833);
nand U7852 (N_7852,N_5312,N_4944);
xor U7853 (N_7853,N_5821,N_4948);
xnor U7854 (N_7854,N_5668,N_5547);
nor U7855 (N_7855,N_4862,N_5697);
nor U7856 (N_7856,N_5315,N_4516);
or U7857 (N_7857,N_4220,N_5473);
and U7858 (N_7858,N_5079,N_5775);
nor U7859 (N_7859,N_5380,N_5433);
xor U7860 (N_7860,N_4319,N_4455);
xor U7861 (N_7861,N_4406,N_4668);
nand U7862 (N_7862,N_4295,N_4866);
or U7863 (N_7863,N_5850,N_4966);
nand U7864 (N_7864,N_5707,N_4750);
and U7865 (N_7865,N_4620,N_4303);
or U7866 (N_7866,N_4149,N_5547);
nand U7867 (N_7867,N_4676,N_4190);
xnor U7868 (N_7868,N_5159,N_5639);
and U7869 (N_7869,N_5378,N_4594);
or U7870 (N_7870,N_5291,N_5171);
xnor U7871 (N_7871,N_4636,N_5954);
and U7872 (N_7872,N_5174,N_4574);
nor U7873 (N_7873,N_5073,N_4279);
and U7874 (N_7874,N_4672,N_4394);
or U7875 (N_7875,N_4480,N_4972);
and U7876 (N_7876,N_4707,N_5933);
or U7877 (N_7877,N_4880,N_4606);
nor U7878 (N_7878,N_4867,N_4008);
and U7879 (N_7879,N_5198,N_5039);
nand U7880 (N_7880,N_4347,N_5819);
nand U7881 (N_7881,N_4649,N_5683);
nor U7882 (N_7882,N_4220,N_4687);
nand U7883 (N_7883,N_4494,N_4543);
and U7884 (N_7884,N_5271,N_4420);
xnor U7885 (N_7885,N_4003,N_4545);
nor U7886 (N_7886,N_5983,N_4671);
nand U7887 (N_7887,N_4509,N_5713);
or U7888 (N_7888,N_5813,N_5693);
or U7889 (N_7889,N_4678,N_4826);
or U7890 (N_7890,N_5154,N_4706);
and U7891 (N_7891,N_4650,N_4051);
or U7892 (N_7892,N_4675,N_5818);
nand U7893 (N_7893,N_4622,N_4692);
and U7894 (N_7894,N_5162,N_5260);
nand U7895 (N_7895,N_4355,N_4310);
nor U7896 (N_7896,N_4661,N_4820);
nand U7897 (N_7897,N_4150,N_5723);
and U7898 (N_7898,N_5138,N_4809);
xnor U7899 (N_7899,N_5295,N_4118);
nand U7900 (N_7900,N_5103,N_5654);
nand U7901 (N_7901,N_5260,N_5779);
nand U7902 (N_7902,N_4035,N_4209);
nand U7903 (N_7903,N_4632,N_5468);
xor U7904 (N_7904,N_5434,N_4723);
nand U7905 (N_7905,N_4731,N_5272);
nor U7906 (N_7906,N_4228,N_4199);
nand U7907 (N_7907,N_4770,N_4283);
or U7908 (N_7908,N_4449,N_5236);
nor U7909 (N_7909,N_5251,N_5163);
and U7910 (N_7910,N_5382,N_5268);
or U7911 (N_7911,N_5029,N_4907);
or U7912 (N_7912,N_4070,N_4152);
nand U7913 (N_7913,N_5026,N_5024);
nand U7914 (N_7914,N_4726,N_5870);
and U7915 (N_7915,N_4360,N_5482);
and U7916 (N_7916,N_4214,N_5721);
xor U7917 (N_7917,N_4630,N_5651);
nor U7918 (N_7918,N_5638,N_4385);
and U7919 (N_7919,N_4117,N_5472);
xor U7920 (N_7920,N_5136,N_4986);
nor U7921 (N_7921,N_5060,N_4750);
and U7922 (N_7922,N_5213,N_5492);
or U7923 (N_7923,N_5499,N_5146);
xnor U7924 (N_7924,N_4142,N_5883);
nor U7925 (N_7925,N_5982,N_4400);
nor U7926 (N_7926,N_5382,N_4342);
and U7927 (N_7927,N_4132,N_5330);
and U7928 (N_7928,N_5181,N_5541);
or U7929 (N_7929,N_5802,N_5539);
nand U7930 (N_7930,N_5008,N_4128);
or U7931 (N_7931,N_4574,N_5981);
nor U7932 (N_7932,N_5793,N_5590);
or U7933 (N_7933,N_5638,N_4478);
nor U7934 (N_7934,N_5150,N_5229);
xnor U7935 (N_7935,N_4638,N_5076);
xnor U7936 (N_7936,N_4761,N_4099);
nor U7937 (N_7937,N_5263,N_4415);
and U7938 (N_7938,N_5318,N_5589);
or U7939 (N_7939,N_4622,N_4831);
nand U7940 (N_7940,N_5037,N_5908);
or U7941 (N_7941,N_4438,N_5750);
nand U7942 (N_7942,N_5508,N_5721);
nand U7943 (N_7943,N_4120,N_4076);
and U7944 (N_7944,N_4385,N_5924);
nor U7945 (N_7945,N_4756,N_4202);
or U7946 (N_7946,N_5929,N_4520);
and U7947 (N_7947,N_4287,N_5831);
nand U7948 (N_7948,N_4951,N_4035);
xor U7949 (N_7949,N_4236,N_4324);
xnor U7950 (N_7950,N_5390,N_4928);
and U7951 (N_7951,N_5815,N_5990);
and U7952 (N_7952,N_5108,N_4176);
and U7953 (N_7953,N_5486,N_4341);
nor U7954 (N_7954,N_4215,N_4080);
nand U7955 (N_7955,N_4494,N_4767);
xor U7956 (N_7956,N_4702,N_5896);
nand U7957 (N_7957,N_4826,N_4268);
and U7958 (N_7958,N_4700,N_5784);
nand U7959 (N_7959,N_5079,N_5038);
nor U7960 (N_7960,N_4766,N_4365);
nand U7961 (N_7961,N_5834,N_5638);
nor U7962 (N_7962,N_4300,N_5692);
nor U7963 (N_7963,N_4188,N_4465);
nand U7964 (N_7964,N_4256,N_5598);
xnor U7965 (N_7965,N_5259,N_4321);
nor U7966 (N_7966,N_5591,N_5889);
nand U7967 (N_7967,N_5347,N_4912);
or U7968 (N_7968,N_4381,N_5709);
xnor U7969 (N_7969,N_4114,N_4086);
nor U7970 (N_7970,N_4606,N_4755);
or U7971 (N_7971,N_4262,N_4999);
xor U7972 (N_7972,N_4860,N_4821);
xor U7973 (N_7973,N_4438,N_4114);
and U7974 (N_7974,N_5503,N_5461);
and U7975 (N_7975,N_5662,N_4578);
xnor U7976 (N_7976,N_4514,N_4584);
nor U7977 (N_7977,N_5621,N_5496);
nor U7978 (N_7978,N_4963,N_4334);
xnor U7979 (N_7979,N_4986,N_4722);
xor U7980 (N_7980,N_5678,N_4044);
or U7981 (N_7981,N_5169,N_4249);
and U7982 (N_7982,N_4556,N_4705);
nor U7983 (N_7983,N_4955,N_4430);
or U7984 (N_7984,N_5891,N_4671);
nand U7985 (N_7985,N_5926,N_5465);
or U7986 (N_7986,N_4739,N_4130);
or U7987 (N_7987,N_4034,N_4989);
nor U7988 (N_7988,N_4717,N_5826);
nor U7989 (N_7989,N_4578,N_4210);
and U7990 (N_7990,N_5565,N_5733);
and U7991 (N_7991,N_5166,N_5545);
nand U7992 (N_7992,N_4674,N_4042);
or U7993 (N_7993,N_5928,N_5965);
and U7994 (N_7994,N_5270,N_4398);
nor U7995 (N_7995,N_5878,N_5338);
nand U7996 (N_7996,N_5315,N_5740);
xnor U7997 (N_7997,N_5094,N_4446);
and U7998 (N_7998,N_5706,N_5276);
or U7999 (N_7999,N_5067,N_4734);
and U8000 (N_8000,N_7248,N_6125);
nand U8001 (N_8001,N_6628,N_7242);
nor U8002 (N_8002,N_7118,N_7320);
nor U8003 (N_8003,N_6327,N_6720);
nor U8004 (N_8004,N_6278,N_7909);
and U8005 (N_8005,N_6520,N_7838);
or U8006 (N_8006,N_6467,N_7938);
nor U8007 (N_8007,N_6683,N_7314);
or U8008 (N_8008,N_7109,N_7408);
and U8009 (N_8009,N_6198,N_6359);
and U8010 (N_8010,N_7936,N_7973);
or U8011 (N_8011,N_6139,N_6430);
and U8012 (N_8012,N_6210,N_6355);
and U8013 (N_8013,N_7734,N_6225);
or U8014 (N_8014,N_6867,N_7986);
nand U8015 (N_8015,N_6681,N_6256);
or U8016 (N_8016,N_6161,N_6824);
or U8017 (N_8017,N_6484,N_6252);
and U8018 (N_8018,N_7181,N_7223);
xnor U8019 (N_8019,N_6343,N_6267);
xnor U8020 (N_8020,N_7797,N_6341);
nor U8021 (N_8021,N_6477,N_7985);
and U8022 (N_8022,N_7081,N_7824);
and U8023 (N_8023,N_7769,N_7130);
nor U8024 (N_8024,N_7550,N_7673);
and U8025 (N_8025,N_6096,N_7955);
or U8026 (N_8026,N_6623,N_6969);
or U8027 (N_8027,N_7645,N_7156);
or U8028 (N_8028,N_6007,N_6769);
nor U8029 (N_8029,N_6751,N_7175);
or U8030 (N_8030,N_6967,N_6631);
nor U8031 (N_8031,N_6912,N_7179);
and U8032 (N_8032,N_6910,N_7937);
and U8033 (N_8033,N_7716,N_7856);
nand U8034 (N_8034,N_6478,N_7153);
or U8035 (N_8035,N_6464,N_7335);
xor U8036 (N_8036,N_7245,N_7813);
and U8037 (N_8037,N_6428,N_7215);
xnor U8038 (N_8038,N_7384,N_7726);
and U8039 (N_8039,N_7641,N_6024);
or U8040 (N_8040,N_6978,N_7024);
xnor U8041 (N_8041,N_6568,N_6587);
nand U8042 (N_8042,N_7880,N_6823);
nor U8043 (N_8043,N_6090,N_6586);
nor U8044 (N_8044,N_6600,N_7648);
or U8045 (N_8045,N_6879,N_6009);
nand U8046 (N_8046,N_7939,N_7547);
and U8047 (N_8047,N_6119,N_7117);
or U8048 (N_8048,N_7947,N_6023);
nor U8049 (N_8049,N_7960,N_6851);
or U8050 (N_8050,N_7950,N_6909);
xor U8051 (N_8051,N_7662,N_7089);
nand U8052 (N_8052,N_6483,N_7587);
or U8053 (N_8053,N_7876,N_6271);
xnor U8054 (N_8054,N_7221,N_6987);
nor U8055 (N_8055,N_6329,N_7386);
nand U8056 (N_8056,N_7885,N_7398);
nor U8057 (N_8057,N_7478,N_7329);
and U8058 (N_8058,N_7093,N_6444);
or U8059 (N_8059,N_6764,N_7006);
and U8060 (N_8060,N_6898,N_6196);
nor U8061 (N_8061,N_7189,N_6420);
nor U8062 (N_8062,N_7476,N_6168);
and U8063 (N_8063,N_6490,N_6924);
or U8064 (N_8064,N_6195,N_7954);
nand U8065 (N_8065,N_6092,N_6440);
nand U8066 (N_8066,N_6018,N_7513);
or U8067 (N_8067,N_7490,N_7239);
or U8068 (N_8068,N_7790,N_6050);
and U8069 (N_8069,N_6858,N_7290);
nor U8070 (N_8070,N_7427,N_7139);
or U8071 (N_8071,N_7007,N_7459);
nand U8072 (N_8072,N_6356,N_7514);
nand U8073 (N_8073,N_6560,N_7857);
nor U8074 (N_8074,N_6553,N_7186);
and U8075 (N_8075,N_7890,N_7423);
nand U8076 (N_8076,N_6905,N_6614);
and U8077 (N_8077,N_7581,N_6411);
nor U8078 (N_8078,N_7968,N_6738);
nand U8079 (N_8079,N_6358,N_7562);
nand U8080 (N_8080,N_7259,N_7703);
nor U8081 (N_8081,N_6468,N_6321);
and U8082 (N_8082,N_6543,N_7681);
xnor U8083 (N_8083,N_7898,N_6556);
nand U8084 (N_8084,N_7772,N_6991);
xnor U8085 (N_8085,N_6122,N_7545);
nand U8086 (N_8086,N_6274,N_7049);
nor U8087 (N_8087,N_7128,N_6871);
nand U8088 (N_8088,N_7832,N_7343);
nor U8089 (N_8089,N_6227,N_7251);
nor U8090 (N_8090,N_6181,N_6776);
nor U8091 (N_8091,N_7820,N_6629);
and U8092 (N_8092,N_6432,N_7348);
nand U8093 (N_8093,N_6272,N_7231);
or U8094 (N_8094,N_7722,N_7426);
or U8095 (N_8095,N_7225,N_6521);
or U8096 (N_8096,N_7262,N_6123);
and U8097 (N_8097,N_7725,N_7786);
nand U8098 (N_8098,N_7578,N_6812);
xnor U8099 (N_8099,N_6756,N_7352);
nor U8100 (N_8100,N_6856,N_7387);
and U8101 (N_8101,N_6998,N_7429);
or U8102 (N_8102,N_6584,N_6646);
xor U8103 (N_8103,N_6796,N_7217);
or U8104 (N_8104,N_7601,N_6708);
nand U8105 (N_8105,N_7064,N_7462);
nor U8106 (N_8106,N_7777,N_7041);
and U8107 (N_8107,N_6627,N_6844);
and U8108 (N_8108,N_6697,N_7733);
nand U8109 (N_8109,N_6204,N_6249);
nor U8110 (N_8110,N_6676,N_7299);
xnor U8111 (N_8111,N_7001,N_6514);
and U8112 (N_8112,N_6216,N_6895);
or U8113 (N_8113,N_7380,N_7235);
or U8114 (N_8114,N_6157,N_6340);
and U8115 (N_8115,N_6182,N_7430);
or U8116 (N_8116,N_6784,N_7405);
and U8117 (N_8117,N_6583,N_6962);
nor U8118 (N_8118,N_6183,N_7188);
and U8119 (N_8119,N_6760,N_7162);
and U8120 (N_8120,N_6828,N_6263);
nand U8121 (N_8121,N_7792,N_7543);
nand U8122 (N_8122,N_7759,N_6965);
xnor U8123 (N_8123,N_7600,N_7308);
or U8124 (N_8124,N_7702,N_6400);
or U8125 (N_8125,N_6480,N_7846);
and U8126 (N_8126,N_6840,N_6379);
and U8127 (N_8127,N_6819,N_6863);
nand U8128 (N_8128,N_6067,N_6402);
or U8129 (N_8129,N_7226,N_7551);
and U8130 (N_8130,N_7526,N_6138);
and U8131 (N_8131,N_7931,N_6184);
xnor U8132 (N_8132,N_7812,N_7686);
xor U8133 (N_8133,N_7135,N_7354);
nor U8134 (N_8134,N_7927,N_7032);
and U8135 (N_8135,N_7353,N_7665);
nor U8136 (N_8136,N_6668,N_7101);
xnor U8137 (N_8137,N_6922,N_6956);
nand U8138 (N_8138,N_6606,N_6588);
nor U8139 (N_8139,N_7253,N_7932);
xnor U8140 (N_8140,N_6372,N_7138);
nand U8141 (N_8141,N_6972,N_7187);
nand U8142 (N_8142,N_6816,N_6407);
xor U8143 (N_8143,N_6382,N_7104);
and U8144 (N_8144,N_7701,N_7840);
and U8145 (N_8145,N_7070,N_7014);
xor U8146 (N_8146,N_7373,N_7620);
xnor U8147 (N_8147,N_6744,N_7009);
or U8148 (N_8148,N_7859,N_6339);
nor U8149 (N_8149,N_6911,N_7029);
or U8150 (N_8150,N_6536,N_6305);
or U8151 (N_8151,N_6317,N_7522);
and U8152 (N_8152,N_6386,N_7437);
nand U8153 (N_8153,N_7349,N_7197);
nand U8154 (N_8154,N_7120,N_7424);
or U8155 (N_8155,N_6699,N_6827);
xnor U8156 (N_8156,N_6270,N_6592);
nor U8157 (N_8157,N_6401,N_6617);
xor U8158 (N_8158,N_6916,N_6378);
xor U8159 (N_8159,N_7285,N_6877);
and U8160 (N_8160,N_6745,N_6041);
or U8161 (N_8161,N_7452,N_7180);
or U8162 (N_8162,N_7465,N_6095);
xor U8163 (N_8163,N_6385,N_7787);
xnor U8164 (N_8164,N_7019,N_7244);
nor U8165 (N_8165,N_6893,N_7311);
nor U8166 (N_8166,N_7296,N_6511);
xnor U8167 (N_8167,N_6179,N_7566);
xnor U8168 (N_8168,N_6365,N_6025);
nand U8169 (N_8169,N_7676,N_7413);
or U8170 (N_8170,N_6740,N_7989);
or U8171 (N_8171,N_7229,N_7607);
nand U8172 (N_8172,N_6498,N_7948);
xnor U8173 (N_8173,N_6188,N_7593);
nand U8174 (N_8174,N_7714,N_7473);
and U8175 (N_8175,N_7281,N_7116);
or U8176 (N_8176,N_7778,N_6361);
nand U8177 (N_8177,N_7590,N_6917);
or U8178 (N_8178,N_6647,N_7495);
and U8179 (N_8179,N_6701,N_6752);
nor U8180 (N_8180,N_6381,N_7420);
nor U8181 (N_8181,N_7396,N_6094);
or U8182 (N_8182,N_7737,N_7715);
or U8183 (N_8183,N_7322,N_6940);
and U8184 (N_8184,N_7054,N_6292);
and U8185 (N_8185,N_7502,N_7580);
nand U8186 (N_8186,N_7650,N_6185);
and U8187 (N_8187,N_6442,N_7884);
nand U8188 (N_8188,N_6121,N_7448);
and U8189 (N_8189,N_6667,N_7228);
nand U8190 (N_8190,N_6154,N_7208);
nor U8191 (N_8191,N_7760,N_6416);
nand U8192 (N_8192,N_7306,N_7643);
or U8193 (N_8193,N_6651,N_7933);
or U8194 (N_8194,N_7026,N_7570);
or U8195 (N_8195,N_6475,N_6370);
nand U8196 (N_8196,N_6808,N_6971);
nor U8197 (N_8197,N_6984,N_6896);
or U8198 (N_8198,N_6187,N_7612);
nor U8199 (N_8199,N_6460,N_7119);
xnor U8200 (N_8200,N_7000,N_7941);
nand U8201 (N_8201,N_7864,N_7952);
or U8202 (N_8202,N_7108,N_7970);
and U8203 (N_8203,N_6307,N_6705);
nand U8204 (N_8204,N_6191,N_7381);
xnor U8205 (N_8205,N_7978,N_7125);
xor U8206 (N_8206,N_7624,N_6215);
nor U8207 (N_8207,N_6704,N_7576);
nor U8208 (N_8208,N_6785,N_6749);
xnor U8209 (N_8209,N_6664,N_6211);
and U8210 (N_8210,N_6208,N_7720);
and U8211 (N_8211,N_6450,N_6008);
xor U8212 (N_8212,N_7916,N_7705);
or U8213 (N_8213,N_6481,N_7501);
xnor U8214 (N_8214,N_7359,N_6678);
xnor U8215 (N_8215,N_7503,N_6457);
and U8216 (N_8216,N_6902,N_7444);
and U8217 (N_8217,N_6383,N_6357);
or U8218 (N_8218,N_7222,N_7477);
nor U8219 (N_8219,N_6492,N_7276);
or U8220 (N_8220,N_6354,N_6878);
nand U8221 (N_8221,N_6380,N_7911);
nor U8222 (N_8222,N_7879,N_7757);
nand U8223 (N_8223,N_7067,N_6688);
xor U8224 (N_8224,N_7694,N_6682);
and U8225 (N_8225,N_6253,N_7496);
xnor U8226 (N_8226,N_7484,N_7653);
xor U8227 (N_8227,N_7390,N_6976);
or U8228 (N_8228,N_7270,N_6777);
nor U8229 (N_8229,N_6530,N_6891);
or U8230 (N_8230,N_7061,N_6257);
nor U8231 (N_8231,N_6202,N_6585);
xor U8232 (N_8232,N_6171,N_7919);
and U8233 (N_8233,N_6223,N_6077);
xor U8234 (N_8234,N_7704,N_7140);
nor U8235 (N_8235,N_6063,N_7469);
xor U8236 (N_8236,N_7920,N_6280);
nand U8237 (N_8237,N_6103,N_6805);
and U8238 (N_8238,N_6316,N_6590);
and U8239 (N_8239,N_6616,N_6780);
xor U8240 (N_8240,N_7345,N_6201);
xor U8241 (N_8241,N_6055,N_7666);
nand U8242 (N_8242,N_7371,N_7300);
xnor U8243 (N_8243,N_7058,N_7637);
and U8244 (N_8244,N_7151,N_6194);
or U8245 (N_8245,N_6189,N_6887);
xnor U8246 (N_8246,N_6961,N_6689);
nand U8247 (N_8247,N_6853,N_7869);
nand U8248 (N_8248,N_6608,N_7991);
nand U8249 (N_8249,N_6581,N_7084);
and U8250 (N_8250,N_7539,N_6353);
nand U8251 (N_8251,N_6758,N_7436);
xnor U8252 (N_8252,N_7830,N_6281);
xnor U8253 (N_8253,N_6564,N_6548);
nand U8254 (N_8254,N_7699,N_6410);
nand U8255 (N_8255,N_7871,N_7038);
nand U8256 (N_8256,N_6802,N_7378);
nand U8257 (N_8257,N_7990,N_6883);
nor U8258 (N_8258,N_6698,N_6391);
nor U8259 (N_8259,N_6546,N_6073);
and U8260 (N_8260,N_6562,N_6959);
and U8261 (N_8261,N_7706,N_6578);
and U8262 (N_8262,N_7440,N_7407);
nor U8263 (N_8263,N_7463,N_7540);
nor U8264 (N_8264,N_7795,N_7866);
xnor U8265 (N_8265,N_7282,N_6456);
nor U8266 (N_8266,N_7619,N_6011);
nor U8267 (N_8267,N_7553,N_6632);
xor U8268 (N_8268,N_6645,N_7798);
nor U8269 (N_8269,N_6015,N_7094);
nor U8270 (N_8270,N_6927,N_6065);
nor U8271 (N_8271,N_7975,N_6933);
or U8272 (N_8272,N_7708,N_7525);
nor U8273 (N_8273,N_7988,N_7212);
xor U8274 (N_8274,N_6388,N_6004);
nor U8275 (N_8275,N_6778,N_6044);
nand U8276 (N_8276,N_6944,N_7048);
and U8277 (N_8277,N_7357,N_7040);
and U8278 (N_8278,N_6031,N_7850);
or U8279 (N_8279,N_7297,N_6220);
or U8280 (N_8280,N_6299,N_7512);
nand U8281 (N_8281,N_6241,N_6835);
nand U8282 (N_8282,N_7728,N_7340);
and U8283 (N_8283,N_7843,N_6782);
nor U8284 (N_8284,N_6890,N_6903);
or U8285 (N_8285,N_6958,N_7546);
nand U8286 (N_8286,N_6957,N_7025);
nor U8287 (N_8287,N_7878,N_7154);
nor U8288 (N_8288,N_6126,N_7141);
nand U8289 (N_8289,N_6621,N_7258);
nand U8290 (N_8290,N_6081,N_6322);
and U8291 (N_8291,N_7383,N_6219);
xor U8292 (N_8292,N_7330,N_6247);
nor U8293 (N_8293,N_6135,N_7595);
nor U8294 (N_8294,N_7822,N_7194);
or U8295 (N_8295,N_7174,N_6638);
and U8296 (N_8296,N_6360,N_7983);
and U8297 (N_8297,N_7957,N_6165);
nand U8298 (N_8298,N_6173,N_7516);
nor U8299 (N_8299,N_6527,N_6088);
nor U8300 (N_8300,N_6177,N_7966);
and U8301 (N_8301,N_6557,N_6742);
nand U8302 (N_8302,N_6659,N_7309);
or U8303 (N_8303,N_7500,N_6532);
nor U8304 (N_8304,N_7249,N_6706);
nand U8305 (N_8305,N_7674,N_7984);
and U8306 (N_8306,N_7661,N_7671);
or U8307 (N_8307,N_7124,N_6261);
or U8308 (N_8308,N_6028,N_7214);
nand U8309 (N_8309,N_7523,N_6443);
nor U8310 (N_8310,N_6641,N_7121);
xnor U8311 (N_8311,N_6394,N_6734);
or U8312 (N_8312,N_6397,N_6938);
nor U8313 (N_8313,N_7642,N_7013);
nor U8314 (N_8314,N_6747,N_6038);
or U8315 (N_8315,N_6537,N_6596);
nand U8316 (N_8316,N_6815,N_7099);
xnor U8317 (N_8317,N_6724,N_6414);
or U8318 (N_8318,N_6026,N_7097);
nand U8319 (N_8319,N_6884,N_6016);
nand U8320 (N_8320,N_6045,N_7697);
xor U8321 (N_8321,N_7268,N_6376);
nand U8322 (N_8322,N_7710,N_7542);
or U8323 (N_8323,N_6533,N_7132);
nor U8324 (N_8324,N_6949,N_6674);
or U8325 (N_8325,N_6097,N_7834);
xor U8326 (N_8326,N_6845,N_6213);
or U8327 (N_8327,N_6921,N_6937);
nand U8328 (N_8328,N_6367,N_7889);
nor U8329 (N_8329,N_7867,N_6577);
nor U8330 (N_8330,N_7411,N_7442);
nor U8331 (N_8331,N_7161,N_6612);
and U8332 (N_8332,N_6132,N_7280);
or U8333 (N_8333,N_7206,N_6419);
or U8334 (N_8334,N_7807,N_6797);
nand U8335 (N_8335,N_7216,N_7134);
or U8336 (N_8336,N_6860,N_6363);
nor U8337 (N_8337,N_7964,N_6714);
and U8338 (N_8338,N_6846,N_7126);
nand U8339 (N_8339,N_7485,N_6572);
nor U8340 (N_8340,N_6968,N_6035);
nor U8341 (N_8341,N_7981,N_6159);
and U8342 (N_8342,N_7374,N_6574);
nor U8343 (N_8343,N_7574,N_7611);
and U8344 (N_8344,N_7457,N_6791);
nor U8345 (N_8345,N_6595,N_6848);
and U8346 (N_8346,N_6610,N_6152);
nand U8347 (N_8347,N_7802,N_6350);
nand U8348 (N_8348,N_6839,N_7895);
and U8349 (N_8349,N_6652,N_6634);
or U8350 (N_8350,N_6392,N_6488);
and U8351 (N_8351,N_6136,N_6452);
or U8352 (N_8352,N_6174,N_6781);
or U8353 (N_8353,N_7450,N_6140);
nor U8354 (N_8354,N_7839,N_7821);
and U8355 (N_8355,N_6282,N_6426);
xor U8356 (N_8356,N_7998,N_6294);
or U8357 (N_8357,N_7963,N_6607);
nor U8358 (N_8358,N_7923,N_7604);
nor U8359 (N_8359,N_7096,N_6995);
or U8360 (N_8360,N_7515,N_7488);
or U8361 (N_8361,N_6807,N_6020);
xnor U8362 (N_8362,N_7199,N_6345);
nand U8363 (N_8363,N_6087,N_6966);
nand U8364 (N_8364,N_6002,N_7896);
xor U8365 (N_8365,N_7063,N_6774);
or U8366 (N_8366,N_6197,N_6541);
nor U8367 (N_8367,N_7819,N_7605);
nand U8368 (N_8368,N_7532,N_6462);
or U8369 (N_8369,N_6232,N_7046);
xor U8370 (N_8370,N_6642,N_7805);
and U8371 (N_8371,N_7266,N_6315);
nor U8372 (N_8372,N_7767,N_7967);
or U8373 (N_8373,N_6108,N_7844);
nor U8374 (N_8374,N_7305,N_6438);
nor U8375 (N_8375,N_6377,N_6311);
xnor U8376 (N_8376,N_7914,N_7635);
nand U8377 (N_8377,N_6763,N_7959);
nand U8378 (N_8378,N_6500,N_6874);
nor U8379 (N_8379,N_6233,N_7918);
xnor U8380 (N_8380,N_6806,N_7803);
nor U8381 (N_8381,N_7557,N_6512);
and U8382 (N_8382,N_6830,N_7237);
or U8383 (N_8383,N_7055,N_7184);
or U8384 (N_8384,N_6466,N_7868);
and U8385 (N_8385,N_6799,N_6408);
and U8386 (N_8386,N_7855,N_7971);
or U8387 (N_8387,N_6078,N_6000);
or U8388 (N_8388,N_7569,N_6996);
xor U8389 (N_8389,N_6037,N_6279);
and U8390 (N_8390,N_6214,N_6670);
xor U8391 (N_8391,N_7507,N_6021);
nand U8392 (N_8392,N_6489,N_7443);
or U8393 (N_8393,N_6680,N_6167);
xor U8394 (N_8394,N_7901,N_6145);
or U8395 (N_8395,N_7874,N_6342);
nor U8396 (N_8396,N_6981,N_7446);
nor U8397 (N_8397,N_7649,N_7627);
nor U8398 (N_8398,N_7086,N_6993);
xor U8399 (N_8399,N_6019,N_7316);
and U8400 (N_8400,N_7050,N_7066);
or U8401 (N_8401,N_6602,N_7492);
xor U8402 (N_8402,N_7454,N_7368);
xor U8403 (N_8403,N_7735,N_6399);
nor U8404 (N_8404,N_7409,N_7887);
nand U8405 (N_8405,N_7092,N_6766);
xor U8406 (N_8406,N_6335,N_7730);
nand U8407 (N_8407,N_7888,N_7471);
xnor U8408 (N_8408,N_7265,N_7913);
or U8409 (N_8409,N_7634,N_7756);
or U8410 (N_8410,N_6569,N_7614);
and U8411 (N_8411,N_7136,N_6690);
nor U8412 (N_8412,N_6719,N_7535);
and U8413 (N_8413,N_6047,N_7934);
nand U8414 (N_8414,N_7801,N_7486);
nor U8415 (N_8415,N_6114,N_6926);
xor U8416 (N_8416,N_6731,N_7291);
and U8417 (N_8417,N_6482,N_6287);
or U8418 (N_8418,N_6507,N_7780);
nand U8419 (N_8419,N_7617,N_7205);
nor U8420 (N_8420,N_7897,N_6324);
xnor U8421 (N_8421,N_7034,N_6499);
nor U8422 (N_8422,N_6547,N_6712);
nand U8423 (N_8423,N_7509,N_7418);
or U8424 (N_8424,N_7173,N_7928);
xnor U8425 (N_8425,N_6373,N_6296);
nor U8426 (N_8426,N_6349,N_7852);
nor U8427 (N_8427,N_6695,N_7679);
nor U8428 (N_8428,N_6212,N_7060);
and U8429 (N_8429,N_7115,N_7949);
and U8430 (N_8430,N_6618,N_7908);
or U8431 (N_8431,N_6346,N_7982);
nor U8432 (N_8432,N_6395,N_7749);
nand U8433 (N_8433,N_6900,N_7201);
nor U8434 (N_8434,N_6264,N_7499);
or U8435 (N_8435,N_7062,N_6091);
and U8436 (N_8436,N_6721,N_6609);
xnor U8437 (N_8437,N_7935,N_6277);
nor U8438 (N_8438,N_6469,N_7388);
xor U8439 (N_8439,N_7393,N_6199);
or U8440 (N_8440,N_6371,N_6773);
xor U8441 (N_8441,N_7365,N_6254);
nand U8442 (N_8442,N_7538,N_6566);
and U8443 (N_8443,N_7399,N_6105);
or U8444 (N_8444,N_6406,N_6694);
and U8445 (N_8445,N_7623,N_7994);
nor U8446 (N_8446,N_6348,N_7762);
and U8447 (N_8447,N_7745,N_6338);
nor U8448 (N_8448,N_7747,N_7346);
nor U8449 (N_8449,N_7709,N_6137);
nor U8450 (N_8450,N_7695,N_6528);
and U8451 (N_8451,N_6071,N_6593);
nand U8452 (N_8452,N_6567,N_6571);
and U8453 (N_8453,N_6064,N_7831);
and U8454 (N_8454,N_7858,N_6117);
and U8455 (N_8455,N_7678,N_6258);
nor U8456 (N_8456,N_6043,N_7339);
nor U8457 (N_8457,N_6765,N_6923);
nand U8458 (N_8458,N_6209,N_7961);
or U8459 (N_8459,N_6857,N_6729);
and U8460 (N_8460,N_6175,N_6473);
nor U8461 (N_8461,N_7647,N_7327);
xnor U8462 (N_8462,N_7761,N_6237);
nand U8463 (N_8463,N_7788,N_7669);
and U8464 (N_8464,N_7255,N_7035);
or U8465 (N_8465,N_7401,N_7690);
nor U8466 (N_8466,N_7603,N_6675);
and U8467 (N_8467,N_7338,N_7571);
nor U8468 (N_8468,N_7129,N_6711);
nor U8469 (N_8469,N_7360,N_6915);
xor U8470 (N_8470,N_6876,N_6613);
nand U8471 (N_8471,N_7766,N_7972);
nor U8472 (N_8472,N_6955,N_6034);
nand U8473 (N_8473,N_7247,N_7015);
nand U8474 (N_8474,N_6529,N_6415);
or U8475 (N_8475,N_6084,N_6746);
xor U8476 (N_8476,N_7583,N_7626);
nand U8477 (N_8477,N_7683,N_7075);
and U8478 (N_8478,N_6149,N_6293);
nand U8479 (N_8479,N_7011,N_7246);
and U8480 (N_8480,N_6673,N_7243);
and U8481 (N_8481,N_6238,N_6029);
or U8482 (N_8482,N_6522,N_7375);
nand U8483 (N_8483,N_7230,N_6717);
and U8484 (N_8484,N_6417,N_7692);
xnor U8485 (N_8485,N_7713,N_6207);
nor U8486 (N_8486,N_6800,N_6169);
or U8487 (N_8487,N_6289,N_7377);
and U8488 (N_8488,N_7763,N_6767);
nand U8489 (N_8489,N_7765,N_7404);
nor U8490 (N_8490,N_6771,N_7417);
nand U8491 (N_8491,N_7750,N_6040);
nor U8492 (N_8492,N_6542,N_7775);
or U8493 (N_8493,N_7740,N_7344);
nor U8494 (N_8494,N_7438,N_6153);
or U8495 (N_8495,N_6463,N_7664);
and U8496 (N_8496,N_7412,N_6288);
xnor U8497 (N_8497,N_7057,N_6396);
nor U8498 (N_8498,N_7472,N_7351);
xnor U8499 (N_8499,N_6795,N_7886);
or U8500 (N_8500,N_6575,N_7165);
or U8501 (N_8501,N_6899,N_6474);
nor U8502 (N_8502,N_6932,N_6244);
nor U8503 (N_8503,N_7332,N_6620);
xor U8504 (N_8504,N_7743,N_6573);
nand U8505 (N_8505,N_7524,N_6850);
xnor U8506 (N_8506,N_7150,N_7877);
xor U8507 (N_8507,N_7579,N_6222);
nor U8508 (N_8508,N_6435,N_6418);
and U8509 (N_8509,N_7675,N_7278);
xnor U8510 (N_8510,N_7475,N_6085);
xor U8511 (N_8511,N_7588,N_7123);
xor U8512 (N_8512,N_7688,N_6504);
nor U8513 (N_8513,N_6821,N_7080);
xor U8514 (N_8514,N_6446,N_6326);
and U8515 (N_8515,N_6068,N_7198);
xnor U8516 (N_8516,N_6847,N_6671);
and U8517 (N_8517,N_6741,N_6082);
nand U8518 (N_8518,N_7814,N_7631);
nand U8519 (N_8519,N_6075,N_6558);
nor U8520 (N_8520,N_7313,N_6591);
or U8521 (N_8521,N_7751,N_6471);
nand U8522 (N_8522,N_7144,N_7263);
nor U8523 (N_8523,N_7657,N_7808);
or U8524 (N_8524,N_6089,N_7541);
nand U8525 (N_8525,N_6496,N_6393);
nor U8526 (N_8526,N_6046,N_7828);
nand U8527 (N_8527,N_6424,N_7148);
or U8528 (N_8528,N_6952,N_6759);
nor U8529 (N_8529,N_6885,N_6003);
and U8530 (N_8530,N_7302,N_6868);
nand U8531 (N_8531,N_6404,N_6757);
xor U8532 (N_8532,N_6875,N_6754);
and U8533 (N_8533,N_7053,N_6579);
nor U8534 (N_8534,N_7930,N_6973);
nand U8535 (N_8535,N_7912,N_6323);
nor U8536 (N_8536,N_7382,N_6156);
or U8537 (N_8537,N_6265,N_7155);
or U8538 (N_8538,N_6104,N_6672);
nor U8539 (N_8539,N_6369,N_6255);
nor U8540 (N_8540,N_7112,N_6702);
or U8541 (N_8541,N_6990,N_6389);
xnor U8542 (N_8542,N_6193,N_7273);
or U8543 (N_8543,N_7369,N_6163);
and U8544 (N_8544,N_6989,N_7656);
or U8545 (N_8545,N_7693,N_6459);
xnor U8546 (N_8546,N_7434,N_6820);
nand U8547 (N_8547,N_7953,N_6918);
nand U8548 (N_8548,N_6873,N_6658);
xor U8549 (N_8549,N_7905,N_6516);
nand U8550 (N_8550,N_6559,N_7680);
nand U8551 (N_8551,N_7347,N_7558);
or U8552 (N_8552,N_6787,N_7536);
nand U8553 (N_8553,N_7872,N_7881);
and U8554 (N_8554,N_7143,N_7289);
xnor U8555 (N_8555,N_7892,N_6409);
xor U8556 (N_8556,N_7773,N_6637);
and U8557 (N_8557,N_7875,N_6398);
and U8558 (N_8558,N_6124,N_7091);
and U8559 (N_8559,N_6344,N_7341);
or U8560 (N_8560,N_7870,N_6120);
nand U8561 (N_8561,N_7453,N_7027);
and U8562 (N_8562,N_6841,N_7506);
nand U8563 (N_8563,N_7068,N_6328);
nand U8564 (N_8564,N_6913,N_7083);
nand U8565 (N_8565,N_7331,N_7530);
or U8566 (N_8566,N_6906,N_7836);
and U8567 (N_8567,N_6116,N_6811);
and U8568 (N_8568,N_7696,N_7017);
and U8569 (N_8569,N_7277,N_6930);
nand U8570 (N_8570,N_6657,N_7196);
and U8571 (N_8571,N_6775,N_7482);
xor U8572 (N_8572,N_6226,N_7774);
xor U8573 (N_8573,N_6640,N_7287);
and U8574 (N_8574,N_7944,N_6331);
nor U8575 (N_8575,N_7312,N_7979);
xor U8576 (N_8576,N_7043,N_6999);
xnor U8577 (N_8577,N_7392,N_6524);
or U8578 (N_8578,N_7395,N_6836);
xor U8579 (N_8579,N_6737,N_7433);
or U8580 (N_8580,N_6098,N_6375);
nand U8581 (N_8581,N_6042,N_6718);
and U8582 (N_8582,N_6242,N_7071);
nor U8583 (N_8583,N_7894,N_6325);
or U8584 (N_8584,N_6582,N_7700);
or U8585 (N_8585,N_7494,N_7724);
and U8586 (N_8586,N_7195,N_6881);
nand U8587 (N_8587,N_6615,N_7211);
or U8588 (N_8588,N_7157,N_7862);
xnor U8589 (N_8589,N_6865,N_7644);
nor U8590 (N_8590,N_7079,N_7668);
nor U8591 (N_8591,N_6235,N_7833);
or U8592 (N_8592,N_6997,N_7639);
nand U8593 (N_8593,N_6421,N_7028);
nand U8594 (N_8594,N_6384,N_7193);
xor U8595 (N_8595,N_6837,N_7582);
nand U8596 (N_8596,N_6655,N_7589);
or U8597 (N_8597,N_6988,N_6790);
or U8598 (N_8598,N_6268,N_6832);
nand U8599 (N_8599,N_6260,N_7002);
nor U8600 (N_8600,N_7817,N_7293);
nand U8601 (N_8601,N_7487,N_6243);
nand U8602 (N_8602,N_7996,N_7727);
nor U8603 (N_8603,N_6493,N_7622);
or U8604 (N_8604,N_7133,N_6928);
nor U8605 (N_8605,N_6535,N_7865);
nor U8606 (N_8606,N_7047,N_6313);
nor U8607 (N_8607,N_7234,N_6713);
or U8608 (N_8608,N_6166,N_6352);
nor U8609 (N_8609,N_6603,N_6437);
xnor U8610 (N_8610,N_7873,N_6920);
nand U8611 (N_8611,N_7292,N_7698);
nor U8612 (N_8612,N_6228,N_6240);
and U8613 (N_8613,N_7575,N_6601);
and U8614 (N_8614,N_6423,N_7511);
nand U8615 (N_8615,N_7660,N_7303);
nor U8616 (N_8616,N_7307,N_6519);
and U8617 (N_8617,N_7044,N_6735);
nor U8618 (N_8618,N_7572,N_7158);
nand U8619 (N_8619,N_6190,N_6405);
nor U8620 (N_8620,N_6710,N_7183);
nand U8621 (N_8621,N_6129,N_6058);
nand U8622 (N_8622,N_6945,N_6831);
or U8623 (N_8623,N_6368,N_7585);
or U8624 (N_8624,N_6192,N_7997);
nor U8625 (N_8625,N_7826,N_7010);
and U8626 (N_8626,N_7168,N_7045);
or U8627 (N_8627,N_6643,N_7385);
or U8628 (N_8628,N_6703,N_7284);
and U8629 (N_8629,N_6290,N_6684);
and U8630 (N_8630,N_7483,N_6864);
nand U8631 (N_8631,N_6074,N_6833);
nand U8632 (N_8632,N_7742,N_7753);
nor U8633 (N_8633,N_6661,N_7748);
xnor U8634 (N_8634,N_7883,N_7391);
xnor U8635 (N_8635,N_7602,N_6901);
and U8636 (N_8636,N_6286,N_7519);
nor U8637 (N_8637,N_7269,N_6245);
nand U8638 (N_8638,N_6297,N_7922);
and U8639 (N_8639,N_6630,N_6334);
xnor U8640 (N_8640,N_7712,N_7491);
or U8641 (N_8641,N_6146,N_6218);
nand U8642 (N_8642,N_6691,N_6598);
nand U8643 (N_8643,N_6069,N_6538);
or U8644 (N_8644,N_7793,N_6622);
and U8645 (N_8645,N_6312,N_7310);
nand U8646 (N_8646,N_7779,N_7213);
nand U8647 (N_8647,N_7853,N_6862);
xor U8648 (N_8648,N_7497,N_6309);
xor U8649 (N_8649,N_7560,N_7992);
and U8650 (N_8650,N_7882,N_7451);
nor U8651 (N_8651,N_7456,N_7167);
or U8652 (N_8652,N_7841,N_6448);
xnor U8653 (N_8653,N_7356,N_6010);
xor U8654 (N_8654,N_6838,N_6054);
nor U8655 (N_8655,N_6118,N_7220);
xnor U8656 (N_8656,N_6455,N_7202);
nand U8657 (N_8657,N_6061,N_6470);
nor U8658 (N_8658,N_7899,N_6934);
nand U8659 (N_8659,N_6128,N_6723);
xnor U8660 (N_8660,N_7264,N_7731);
and U8661 (N_8661,N_6515,N_7609);
nor U8662 (N_8662,N_6770,N_6472);
xnor U8663 (N_8663,N_6318,N_6130);
nand U8664 (N_8664,N_6251,N_7466);
xnor U8665 (N_8665,N_6413,N_6142);
xor U8666 (N_8666,N_6950,N_6649);
and U8667 (N_8667,N_6486,N_7283);
nor U8668 (N_8668,N_6291,N_6206);
nand U8669 (N_8669,N_7073,N_7517);
and U8670 (N_8670,N_7238,N_7672);
xnor U8671 (N_8671,N_6155,N_6813);
and U8672 (N_8672,N_7659,N_6205);
nand U8673 (N_8673,N_7677,N_7554);
nor U8674 (N_8674,N_7837,N_7719);
xnor U8675 (N_8675,N_6809,N_6727);
nand U8676 (N_8676,N_6465,N_7379);
and U8677 (N_8677,N_6056,N_7470);
nor U8678 (N_8678,N_6725,N_6872);
xnor U8679 (N_8679,N_7372,N_7510);
and U8680 (N_8680,N_6093,N_6870);
nand U8681 (N_8681,N_6433,N_6259);
xnor U8682 (N_8682,N_7711,N_6929);
nor U8683 (N_8683,N_6677,N_6036);
xor U8684 (N_8684,N_7078,N_7563);
and U8685 (N_8685,N_7192,N_7616);
or U8686 (N_8686,N_7410,N_6692);
nor U8687 (N_8687,N_6427,N_7394);
and U8688 (N_8688,N_7036,N_6611);
xnor U8689 (N_8689,N_7561,N_7361);
or U8690 (N_8690,N_7783,N_6434);
or U8691 (N_8691,N_7037,N_7319);
nor U8692 (N_8692,N_6822,N_7921);
and U8693 (N_8693,N_7304,N_6390);
nand U8694 (N_8694,N_7823,N_7439);
or U8695 (N_8695,N_6508,N_6626);
nand U8696 (N_8696,N_6888,N_7317);
and U8697 (N_8697,N_7529,N_6476);
and U8698 (N_8698,N_6669,N_6302);
nand U8699 (N_8699,N_6964,N_7738);
nor U8700 (N_8700,N_7321,N_7518);
or U8701 (N_8701,N_6453,N_6861);
nand U8702 (N_8702,N_7827,N_6027);
nor U8703 (N_8703,N_6889,N_6604);
nand U8704 (N_8704,N_7236,N_6221);
nor U8705 (N_8705,N_7549,N_7107);
xor U8706 (N_8706,N_7333,N_7358);
nand U8707 (N_8707,N_6495,N_7568);
xor U8708 (N_8708,N_6908,N_6148);
xnor U8709 (N_8709,N_7033,N_7721);
nand U8710 (N_8710,N_7977,N_6180);
and U8711 (N_8711,N_7400,N_7425);
xnor U8712 (N_8712,N_6979,N_7207);
nand U8713 (N_8713,N_7537,N_7829);
and U8714 (N_8714,N_7275,N_6374);
or U8715 (N_8715,N_7818,N_6239);
and U8716 (N_8716,N_7298,N_7785);
and U8717 (N_8717,N_6295,N_7219);
nor U8718 (N_8718,N_6513,N_7638);
xor U8719 (N_8719,N_6366,N_7599);
or U8720 (N_8720,N_6992,N_7271);
or U8721 (N_8721,N_6494,N_7781);
nand U8722 (N_8722,N_7816,N_6447);
and U8723 (N_8723,N_7461,N_7825);
and U8724 (N_8724,N_6314,N_7528);
nand U8725 (N_8725,N_7111,N_7164);
nand U8726 (N_8726,N_7565,N_6186);
xnor U8727 (N_8727,N_6510,N_7663);
and U8728 (N_8728,N_6320,N_7854);
or U8729 (N_8729,N_6052,N_7445);
nand U8730 (N_8730,N_7191,N_6422);
nor U8731 (N_8731,N_6269,N_7629);
and U8732 (N_8732,N_7210,N_7056);
or U8733 (N_8733,N_6479,N_7008);
nand U8734 (N_8734,N_7481,N_7020);
nand U8735 (N_8735,N_7039,N_6429);
xor U8736 (N_8736,N_6762,N_6005);
xnor U8737 (N_8737,N_7946,N_7995);
nor U8738 (N_8738,N_6539,N_6234);
nand U8739 (N_8739,N_7567,N_7159);
xnor U8740 (N_8740,N_7288,N_6852);
nand U8741 (N_8741,N_6246,N_6485);
nand U8742 (N_8742,N_6347,N_7204);
nand U8743 (N_8743,N_7993,N_7640);
or U8744 (N_8744,N_6554,N_7171);
xor U8745 (N_8745,N_7004,N_6788);
nand U8746 (N_8746,N_6109,N_6855);
and U8747 (N_8747,N_6250,N_7106);
and U8748 (N_8748,N_7707,N_6273);
nand U8749 (N_8749,N_7597,N_7910);
and U8750 (N_8750,N_6070,N_7435);
nand U8751 (N_8751,N_7023,N_7342);
and U8752 (N_8752,N_7907,N_7924);
xor U8753 (N_8753,N_7504,N_6013);
nor U8754 (N_8754,N_7687,N_7630);
xnor U8755 (N_8755,N_6663,N_6436);
or U8756 (N_8756,N_7279,N_7615);
nand U8757 (N_8757,N_7799,N_6276);
nor U8758 (N_8758,N_7085,N_7098);
or U8759 (N_8759,N_6057,N_7464);
and U8760 (N_8760,N_6894,N_7958);
and U8761 (N_8761,N_6076,N_7110);
and U8762 (N_8762,N_7428,N_6101);
nor U8763 (N_8763,N_6960,N_6062);
and U8764 (N_8764,N_6006,N_7256);
nand U8765 (N_8765,N_7209,N_6080);
xnor U8766 (N_8766,N_7127,N_6115);
nand U8767 (N_8767,N_7969,N_7052);
nand U8768 (N_8768,N_6589,N_7328);
and U8769 (N_8769,N_6935,N_7744);
or U8770 (N_8770,N_7754,N_7337);
nand U8771 (N_8771,N_6563,N_6113);
and U8772 (N_8772,N_6946,N_6203);
nand U8773 (N_8773,N_7069,N_6387);
xnor U8774 (N_8774,N_6597,N_7416);
xnor U8775 (N_8775,N_7200,N_6750);
nor U8776 (N_8776,N_6985,N_6412);
and U8777 (N_8777,N_7533,N_7636);
nor U8778 (N_8778,N_6941,N_7421);
nor U8779 (N_8779,N_7218,N_7489);
nor U8780 (N_8780,N_7422,N_7042);
nand U8781 (N_8781,N_7012,N_7625);
or U8782 (N_8782,N_7861,N_7527);
nand U8783 (N_8783,N_7460,N_7628);
and U8784 (N_8784,N_7355,N_7739);
xor U8785 (N_8785,N_6625,N_7531);
nand U8786 (N_8786,N_6753,N_7403);
and U8787 (N_8787,N_7021,N_7318);
and U8788 (N_8788,N_7670,N_6033);
nand U8789 (N_8789,N_6817,N_6728);
or U8790 (N_8790,N_6656,N_6977);
xor U8791 (N_8791,N_6818,N_7474);
and U8792 (N_8792,N_7586,N_6685);
nand U8793 (N_8793,N_7552,N_7367);
xnor U8794 (N_8794,N_6914,N_6308);
and U8795 (N_8795,N_6502,N_6943);
nand U8796 (N_8796,N_7521,N_7315);
nor U8797 (N_8797,N_6696,N_7018);
nand U8798 (N_8798,N_7178,N_7286);
and U8799 (N_8799,N_6049,N_6783);
and U8800 (N_8800,N_6150,N_6869);
nor U8801 (N_8801,N_6403,N_6106);
xnor U8802 (N_8802,N_7493,N_6351);
nor U8803 (N_8803,N_6039,N_6079);
nor U8804 (N_8804,N_7224,N_6147);
xnor U8805 (N_8805,N_7847,N_6772);
nor U8806 (N_8806,N_6127,N_7652);
and U8807 (N_8807,N_6266,N_6112);
nand U8808 (N_8808,N_7172,N_7362);
or U8809 (N_8809,N_7016,N_6953);
nand U8810 (N_8810,N_7606,N_6882);
nand U8811 (N_8811,N_7447,N_6285);
xor U8812 (N_8812,N_6229,N_7806);
or U8813 (N_8813,N_7942,N_6102);
or U8814 (N_8814,N_7431,N_6051);
xnor U8815 (N_8815,N_6866,N_6523);
nor U8816 (N_8816,N_7350,N_7689);
xor U8817 (N_8817,N_7682,N_6650);
or U8818 (N_8818,N_7845,N_7102);
nand U8819 (N_8819,N_7684,N_6275);
nor U8820 (N_8820,N_7718,N_7146);
xnor U8821 (N_8821,N_6525,N_6665);
or U8822 (N_8822,N_6635,N_7573);
nor U8823 (N_8823,N_6158,N_7940);
nand U8824 (N_8824,N_6176,N_7945);
nand U8825 (N_8825,N_7272,N_6099);
nand U8826 (N_8826,N_7863,N_6144);
nor U8827 (N_8827,N_6059,N_7632);
nand U8828 (N_8828,N_6501,N_7592);
nor U8829 (N_8829,N_7613,N_7241);
and U8830 (N_8830,N_7943,N_6304);
nand U8831 (N_8831,N_7131,N_6134);
or U8832 (N_8832,N_7090,N_6552);
and U8833 (N_8833,N_6636,N_7893);
nor U8834 (N_8834,N_7903,N_7406);
and U8835 (N_8835,N_7325,N_6505);
nand U8836 (N_8836,N_6743,N_7336);
nand U8837 (N_8837,N_7752,N_6594);
nor U8838 (N_8838,N_6301,N_7182);
nor U8839 (N_8839,N_7082,N_7294);
xnor U8840 (N_8840,N_6733,N_7851);
or U8841 (N_8841,N_6722,N_6540);
nor U8842 (N_8842,N_6970,N_7800);
nand U8843 (N_8843,N_7114,N_6164);
or U8844 (N_8844,N_6693,N_6810);
or U8845 (N_8845,N_6425,N_6826);
nand U8846 (N_8846,N_6798,N_7402);
nand U8847 (N_8847,N_6599,N_7758);
nand U8848 (N_8848,N_6892,N_7770);
nand U8849 (N_8849,N_7902,N_7260);
and U8850 (N_8850,N_6644,N_6441);
and U8851 (N_8851,N_7925,N_7685);
nor U8852 (N_8852,N_7577,N_6732);
nand U8853 (N_8853,N_7441,N_6503);
xor U8854 (N_8854,N_7295,N_6333);
or U8855 (N_8855,N_7776,N_7419);
nand U8856 (N_8856,N_7796,N_6451);
and U8857 (N_8857,N_7559,N_6716);
nor U8858 (N_8858,N_6829,N_7065);
nor U8859 (N_8859,N_6100,N_6761);
xnor U8860 (N_8860,N_6555,N_7505);
and U8861 (N_8861,N_7654,N_7729);
or U8862 (N_8862,N_7176,N_6880);
xor U8863 (N_8863,N_7003,N_7074);
nor U8864 (N_8864,N_7646,N_7584);
and U8865 (N_8865,N_7113,N_7261);
nand U8866 (N_8866,N_6662,N_6200);
or U8867 (N_8867,N_7555,N_6886);
nor U8868 (N_8868,N_6975,N_7432);
xnor U8869 (N_8869,N_6231,N_6686);
and U8870 (N_8870,N_7598,N_6550);
or U8871 (N_8871,N_6794,N_7962);
or U8872 (N_8872,N_6963,N_6904);
xor U8873 (N_8873,N_6679,N_6298);
and U8874 (N_8874,N_7667,N_6730);
nand U8875 (N_8875,N_6700,N_7926);
nor U8876 (N_8876,N_6283,N_6531);
nor U8877 (N_8877,N_6217,N_6300);
nand U8878 (N_8878,N_7480,N_6983);
or U8879 (N_8879,N_6624,N_7250);
and U8880 (N_8880,N_7891,N_6709);
xor U8881 (N_8881,N_7051,N_6947);
and U8882 (N_8882,N_7804,N_7784);
nor U8883 (N_8883,N_7915,N_6224);
nand U8884 (N_8884,N_6925,N_6951);
xor U8885 (N_8885,N_7771,N_7254);
nor U8886 (N_8886,N_6633,N_7232);
xor U8887 (N_8887,N_7951,N_6160);
and U8888 (N_8888,N_7257,N_7621);
or U8889 (N_8889,N_7651,N_6801);
nand U8890 (N_8890,N_7789,N_6110);
or U8891 (N_8891,N_6162,N_7768);
nand U8892 (N_8892,N_6032,N_7147);
nor U8893 (N_8893,N_6534,N_7534);
nor U8894 (N_8894,N_6942,N_7142);
nand U8895 (N_8895,N_7240,N_6248);
nand U8896 (N_8896,N_7556,N_6337);
nor U8897 (N_8897,N_6726,N_7811);
xor U8898 (N_8898,N_7976,N_6549);
xnor U8899 (N_8899,N_6580,N_7965);
and U8900 (N_8900,N_6936,N_7326);
xnor U8901 (N_8901,N_7468,N_7455);
nand U8902 (N_8902,N_7177,N_7149);
and U8903 (N_8903,N_7906,N_7520);
nand U8904 (N_8904,N_6907,N_7397);
nand U8905 (N_8905,N_6178,N_7904);
or U8906 (N_8906,N_7544,N_6060);
and U8907 (N_8907,N_6445,N_7633);
nand U8908 (N_8908,N_7185,N_7324);
nand U8909 (N_8909,N_6362,N_6001);
nor U8910 (N_8910,N_6687,N_7956);
nand U8911 (N_8911,N_7366,N_7810);
and U8912 (N_8912,N_6653,N_6994);
nor U8913 (N_8913,N_7746,N_7364);
nor U8914 (N_8914,N_6141,N_7005);
and U8915 (N_8915,N_7301,N_7618);
or U8916 (N_8916,N_6948,N_6506);
nand U8917 (N_8917,N_6825,N_7999);
nand U8918 (N_8918,N_6517,N_6230);
nor U8919 (N_8919,N_6639,N_7596);
nor U8920 (N_8920,N_6748,N_6814);
or U8921 (N_8921,N_6458,N_7170);
nand U8922 (N_8922,N_6803,N_6561);
and U8923 (N_8923,N_6364,N_7087);
and U8924 (N_8924,N_6793,N_7103);
xor U8925 (N_8925,N_6012,N_7498);
xnor U8926 (N_8926,N_6332,N_7608);
nor U8927 (N_8927,N_6066,N_7145);
nand U8928 (N_8928,N_6319,N_7031);
nand U8929 (N_8929,N_6449,N_6431);
or U8930 (N_8930,N_7610,N_7163);
xnor U8931 (N_8931,N_6048,N_6954);
nor U8932 (N_8932,N_6565,N_6014);
nand U8933 (N_8933,N_7059,N_6786);
nor U8934 (N_8934,N_6974,N_7233);
and U8935 (N_8935,N_7974,N_7137);
xor U8936 (N_8936,N_7691,N_7389);
and U8937 (N_8937,N_7166,N_6619);
and U8938 (N_8938,N_7467,N_6804);
nor U8939 (N_8939,N_7794,N_6654);
xnor U8940 (N_8940,N_7848,N_6854);
or U8941 (N_8941,N_7723,N_7900);
and U8942 (N_8942,N_7203,N_7076);
nand U8943 (N_8943,N_7414,N_7860);
or U8944 (N_8944,N_6660,N_6792);
xor U8945 (N_8945,N_7842,N_6236);
and U8946 (N_8946,N_7980,N_6336);
or U8947 (N_8947,N_6072,N_7169);
nor U8948 (N_8948,N_6570,N_6897);
nor U8949 (N_8949,N_7987,N_7449);
nor U8950 (N_8950,N_7741,N_6170);
and U8951 (N_8951,N_6310,N_7594);
and U8952 (N_8952,N_6306,N_7363);
nor U8953 (N_8953,N_6133,N_6834);
xor U8954 (N_8954,N_6131,N_7849);
nand U8955 (N_8955,N_6518,N_6859);
or U8956 (N_8956,N_7458,N_7508);
nor U8957 (N_8957,N_6017,N_7088);
nor U8958 (N_8958,N_6939,N_6111);
nor U8959 (N_8959,N_7274,N_6053);
nand U8960 (N_8960,N_6768,N_7479);
nand U8961 (N_8961,N_7190,N_7252);
or U8962 (N_8962,N_7030,N_6982);
or U8963 (N_8963,N_6461,N_7415);
xor U8964 (N_8964,N_7755,N_7370);
or U8965 (N_8965,N_6736,N_6980);
and U8966 (N_8966,N_7736,N_6986);
and U8967 (N_8967,N_6605,N_6666);
nor U8968 (N_8968,N_7717,N_7548);
nand U8969 (N_8969,N_6330,N_6739);
xnor U8970 (N_8970,N_7022,N_7591);
xor U8971 (N_8971,N_7564,N_6931);
or U8972 (N_8972,N_6707,N_6030);
or U8973 (N_8973,N_6284,N_7732);
and U8974 (N_8974,N_7334,N_7072);
nand U8975 (N_8975,N_7152,N_6551);
nand U8976 (N_8976,N_6151,N_6487);
and U8977 (N_8977,N_7267,N_7376);
nor U8978 (N_8978,N_6919,N_6143);
nor U8979 (N_8979,N_6755,N_6779);
nor U8980 (N_8980,N_7095,N_6454);
or U8981 (N_8981,N_6172,N_6022);
xnor U8982 (N_8982,N_7815,N_7917);
nor U8983 (N_8983,N_7809,N_7791);
and U8984 (N_8984,N_6648,N_6789);
nor U8985 (N_8985,N_7105,N_6545);
xnor U8986 (N_8986,N_7782,N_7835);
xnor U8987 (N_8987,N_7658,N_6083);
xnor U8988 (N_8988,N_6849,N_7323);
or U8989 (N_8989,N_6086,N_6262);
xor U8990 (N_8990,N_6576,N_6303);
xor U8991 (N_8991,N_6491,N_7655);
xor U8992 (N_8992,N_7160,N_6509);
nand U8993 (N_8993,N_6843,N_7227);
and U8994 (N_8994,N_7077,N_6439);
and U8995 (N_8995,N_6842,N_6526);
xor U8996 (N_8996,N_7122,N_6497);
nand U8997 (N_8997,N_7100,N_6544);
nand U8998 (N_8998,N_6107,N_7764);
nor U8999 (N_8999,N_6715,N_7929);
or U9000 (N_9000,N_6573,N_6620);
and U9001 (N_9001,N_6976,N_7710);
or U9002 (N_9002,N_7708,N_6137);
and U9003 (N_9003,N_7588,N_6035);
and U9004 (N_9004,N_6481,N_6722);
nor U9005 (N_9005,N_6193,N_7507);
nor U9006 (N_9006,N_7121,N_6235);
and U9007 (N_9007,N_6755,N_7811);
or U9008 (N_9008,N_7203,N_6407);
nand U9009 (N_9009,N_7734,N_7853);
xor U9010 (N_9010,N_7722,N_6277);
nand U9011 (N_9011,N_6427,N_6690);
and U9012 (N_9012,N_7764,N_7100);
or U9013 (N_9013,N_7000,N_6504);
or U9014 (N_9014,N_6155,N_7658);
and U9015 (N_9015,N_7046,N_7653);
nor U9016 (N_9016,N_6134,N_7567);
and U9017 (N_9017,N_6408,N_7898);
xor U9018 (N_9018,N_7428,N_7117);
or U9019 (N_9019,N_6740,N_6746);
nand U9020 (N_9020,N_7578,N_6764);
nand U9021 (N_9021,N_7486,N_7547);
or U9022 (N_9022,N_6126,N_6132);
xor U9023 (N_9023,N_7717,N_6063);
and U9024 (N_9024,N_7090,N_7742);
xor U9025 (N_9025,N_7531,N_7069);
nor U9026 (N_9026,N_7358,N_7386);
nand U9027 (N_9027,N_6260,N_6937);
nor U9028 (N_9028,N_6255,N_6909);
nor U9029 (N_9029,N_6891,N_7070);
xnor U9030 (N_9030,N_6136,N_7214);
and U9031 (N_9031,N_7447,N_6551);
xor U9032 (N_9032,N_7088,N_7004);
and U9033 (N_9033,N_7946,N_7594);
or U9034 (N_9034,N_6748,N_7058);
or U9035 (N_9035,N_7685,N_7985);
nor U9036 (N_9036,N_7417,N_7624);
and U9037 (N_9037,N_6072,N_6597);
and U9038 (N_9038,N_6511,N_6759);
or U9039 (N_9039,N_6450,N_7040);
and U9040 (N_9040,N_6631,N_7083);
xnor U9041 (N_9041,N_7474,N_7767);
nor U9042 (N_9042,N_6451,N_7760);
and U9043 (N_9043,N_7710,N_6846);
or U9044 (N_9044,N_7980,N_6706);
nor U9045 (N_9045,N_6700,N_7611);
nor U9046 (N_9046,N_7701,N_6186);
nand U9047 (N_9047,N_7651,N_7827);
nand U9048 (N_9048,N_7632,N_7380);
and U9049 (N_9049,N_7766,N_7842);
xor U9050 (N_9050,N_6618,N_6341);
xor U9051 (N_9051,N_7247,N_6935);
and U9052 (N_9052,N_7589,N_7279);
nor U9053 (N_9053,N_7450,N_6874);
nor U9054 (N_9054,N_6365,N_6320);
xor U9055 (N_9055,N_6389,N_7608);
or U9056 (N_9056,N_6207,N_7349);
or U9057 (N_9057,N_6244,N_6942);
nand U9058 (N_9058,N_7205,N_7515);
xnor U9059 (N_9059,N_6201,N_7634);
and U9060 (N_9060,N_6324,N_7399);
xnor U9061 (N_9061,N_6327,N_6349);
xnor U9062 (N_9062,N_7631,N_6896);
nor U9063 (N_9063,N_6667,N_7314);
nand U9064 (N_9064,N_7890,N_6863);
nand U9065 (N_9065,N_7692,N_7282);
and U9066 (N_9066,N_6431,N_6772);
xnor U9067 (N_9067,N_7983,N_6140);
nor U9068 (N_9068,N_7258,N_7191);
or U9069 (N_9069,N_6682,N_6707);
or U9070 (N_9070,N_7920,N_6708);
or U9071 (N_9071,N_6735,N_7099);
nand U9072 (N_9072,N_6970,N_6173);
or U9073 (N_9073,N_7863,N_6187);
nand U9074 (N_9074,N_6024,N_6007);
and U9075 (N_9075,N_7263,N_6497);
or U9076 (N_9076,N_6087,N_7769);
and U9077 (N_9077,N_6276,N_6041);
nor U9078 (N_9078,N_7376,N_6163);
and U9079 (N_9079,N_6489,N_7019);
nand U9080 (N_9080,N_6477,N_6641);
or U9081 (N_9081,N_7272,N_7784);
or U9082 (N_9082,N_7701,N_6107);
and U9083 (N_9083,N_6470,N_7754);
or U9084 (N_9084,N_7698,N_7288);
nand U9085 (N_9085,N_6185,N_7331);
and U9086 (N_9086,N_6433,N_6059);
and U9087 (N_9087,N_7834,N_7895);
or U9088 (N_9088,N_6676,N_7365);
nor U9089 (N_9089,N_6470,N_7899);
nand U9090 (N_9090,N_6225,N_6938);
nor U9091 (N_9091,N_6492,N_6157);
xor U9092 (N_9092,N_6980,N_6652);
or U9093 (N_9093,N_7136,N_7191);
or U9094 (N_9094,N_6303,N_7165);
and U9095 (N_9095,N_7766,N_6819);
nand U9096 (N_9096,N_6100,N_6623);
or U9097 (N_9097,N_7544,N_6808);
and U9098 (N_9098,N_7632,N_6991);
nor U9099 (N_9099,N_6771,N_7088);
nor U9100 (N_9100,N_6015,N_7664);
nand U9101 (N_9101,N_7404,N_6695);
nand U9102 (N_9102,N_7406,N_7969);
and U9103 (N_9103,N_6315,N_7011);
or U9104 (N_9104,N_6316,N_6195);
nor U9105 (N_9105,N_6072,N_6788);
nand U9106 (N_9106,N_7495,N_7567);
nor U9107 (N_9107,N_6012,N_6061);
and U9108 (N_9108,N_6967,N_7090);
nand U9109 (N_9109,N_7420,N_7319);
nand U9110 (N_9110,N_7055,N_6379);
nand U9111 (N_9111,N_6538,N_6356);
and U9112 (N_9112,N_6442,N_6039);
xnor U9113 (N_9113,N_7444,N_6623);
and U9114 (N_9114,N_6248,N_7660);
nor U9115 (N_9115,N_6561,N_7072);
or U9116 (N_9116,N_7531,N_6681);
nor U9117 (N_9117,N_7968,N_6730);
xnor U9118 (N_9118,N_7123,N_6519);
or U9119 (N_9119,N_6832,N_6673);
xor U9120 (N_9120,N_7977,N_7347);
nand U9121 (N_9121,N_6019,N_7283);
nand U9122 (N_9122,N_7585,N_6698);
nand U9123 (N_9123,N_6774,N_7561);
nand U9124 (N_9124,N_6584,N_6215);
xor U9125 (N_9125,N_6695,N_7689);
and U9126 (N_9126,N_7504,N_6695);
and U9127 (N_9127,N_6296,N_6969);
nand U9128 (N_9128,N_7898,N_7573);
nor U9129 (N_9129,N_6498,N_6992);
nand U9130 (N_9130,N_7818,N_6677);
or U9131 (N_9131,N_6356,N_6264);
or U9132 (N_9132,N_7863,N_7038);
nand U9133 (N_9133,N_7926,N_7364);
or U9134 (N_9134,N_7668,N_7478);
nand U9135 (N_9135,N_7499,N_6151);
or U9136 (N_9136,N_6192,N_7041);
nor U9137 (N_9137,N_7016,N_6790);
nand U9138 (N_9138,N_7333,N_7929);
or U9139 (N_9139,N_6857,N_6465);
nor U9140 (N_9140,N_7600,N_6901);
or U9141 (N_9141,N_7112,N_6355);
or U9142 (N_9142,N_7946,N_6953);
or U9143 (N_9143,N_6402,N_6755);
xnor U9144 (N_9144,N_6281,N_6754);
or U9145 (N_9145,N_6171,N_6122);
or U9146 (N_9146,N_7565,N_7139);
xnor U9147 (N_9147,N_6111,N_6902);
and U9148 (N_9148,N_6563,N_7327);
or U9149 (N_9149,N_7045,N_6993);
xnor U9150 (N_9150,N_6078,N_7978);
and U9151 (N_9151,N_7041,N_7355);
nand U9152 (N_9152,N_7420,N_7871);
and U9153 (N_9153,N_6321,N_7072);
or U9154 (N_9154,N_6701,N_7854);
or U9155 (N_9155,N_7921,N_7234);
or U9156 (N_9156,N_6860,N_7825);
or U9157 (N_9157,N_7706,N_6070);
or U9158 (N_9158,N_6432,N_6813);
nor U9159 (N_9159,N_6685,N_6551);
nand U9160 (N_9160,N_6489,N_7920);
and U9161 (N_9161,N_6042,N_7996);
or U9162 (N_9162,N_7091,N_6812);
nand U9163 (N_9163,N_7626,N_6215);
and U9164 (N_9164,N_6487,N_7015);
xor U9165 (N_9165,N_7500,N_6166);
xor U9166 (N_9166,N_6981,N_7503);
nor U9167 (N_9167,N_6458,N_6220);
and U9168 (N_9168,N_6931,N_6394);
nor U9169 (N_9169,N_6010,N_6863);
and U9170 (N_9170,N_7694,N_6638);
or U9171 (N_9171,N_7552,N_6711);
or U9172 (N_9172,N_6068,N_6210);
nand U9173 (N_9173,N_6938,N_6141);
xor U9174 (N_9174,N_7367,N_6041);
nor U9175 (N_9175,N_7881,N_7364);
xnor U9176 (N_9176,N_7301,N_6697);
nor U9177 (N_9177,N_6669,N_6535);
or U9178 (N_9178,N_7574,N_6954);
and U9179 (N_9179,N_6607,N_6102);
nor U9180 (N_9180,N_6096,N_7429);
nand U9181 (N_9181,N_6708,N_6349);
xnor U9182 (N_9182,N_6420,N_6409);
nand U9183 (N_9183,N_7133,N_6718);
nor U9184 (N_9184,N_7004,N_6529);
or U9185 (N_9185,N_6946,N_6395);
and U9186 (N_9186,N_6183,N_6580);
nor U9187 (N_9187,N_7208,N_7312);
and U9188 (N_9188,N_7345,N_7816);
nor U9189 (N_9189,N_7333,N_6699);
nor U9190 (N_9190,N_7859,N_6881);
xnor U9191 (N_9191,N_6421,N_6351);
nand U9192 (N_9192,N_7014,N_7455);
nand U9193 (N_9193,N_6998,N_7699);
or U9194 (N_9194,N_7596,N_6386);
nor U9195 (N_9195,N_7275,N_7404);
xor U9196 (N_9196,N_7892,N_7221);
nor U9197 (N_9197,N_6142,N_7483);
xnor U9198 (N_9198,N_6148,N_7203);
or U9199 (N_9199,N_7459,N_7613);
nand U9200 (N_9200,N_6021,N_6935);
nand U9201 (N_9201,N_7247,N_6333);
nor U9202 (N_9202,N_6569,N_7795);
or U9203 (N_9203,N_6997,N_7339);
and U9204 (N_9204,N_6721,N_6056);
nand U9205 (N_9205,N_7104,N_7762);
nand U9206 (N_9206,N_6825,N_7978);
and U9207 (N_9207,N_6404,N_7173);
nand U9208 (N_9208,N_6556,N_6822);
nand U9209 (N_9209,N_7907,N_7029);
nor U9210 (N_9210,N_7795,N_7699);
xnor U9211 (N_9211,N_6471,N_7589);
or U9212 (N_9212,N_6022,N_7258);
xor U9213 (N_9213,N_6243,N_7402);
xnor U9214 (N_9214,N_6602,N_7261);
or U9215 (N_9215,N_6210,N_7457);
nand U9216 (N_9216,N_7923,N_6434);
xnor U9217 (N_9217,N_6674,N_7149);
xor U9218 (N_9218,N_7383,N_7587);
nor U9219 (N_9219,N_7145,N_7418);
nor U9220 (N_9220,N_7537,N_7524);
or U9221 (N_9221,N_7610,N_6285);
xnor U9222 (N_9222,N_7846,N_6898);
and U9223 (N_9223,N_7992,N_6086);
nand U9224 (N_9224,N_6230,N_6466);
xnor U9225 (N_9225,N_7115,N_6453);
and U9226 (N_9226,N_6349,N_6566);
xnor U9227 (N_9227,N_7451,N_6646);
xnor U9228 (N_9228,N_7415,N_6635);
nor U9229 (N_9229,N_7623,N_7741);
nand U9230 (N_9230,N_7758,N_7645);
nor U9231 (N_9231,N_6641,N_6867);
nand U9232 (N_9232,N_7970,N_7205);
nor U9233 (N_9233,N_7746,N_6469);
and U9234 (N_9234,N_6574,N_6502);
and U9235 (N_9235,N_7500,N_7813);
nand U9236 (N_9236,N_7283,N_6079);
nand U9237 (N_9237,N_6363,N_7431);
and U9238 (N_9238,N_6975,N_7855);
nor U9239 (N_9239,N_6851,N_7188);
or U9240 (N_9240,N_6229,N_6234);
nor U9241 (N_9241,N_7408,N_6757);
and U9242 (N_9242,N_6999,N_7795);
and U9243 (N_9243,N_7156,N_6964);
or U9244 (N_9244,N_7530,N_6740);
xor U9245 (N_9245,N_7892,N_7270);
nor U9246 (N_9246,N_6316,N_6865);
nand U9247 (N_9247,N_6824,N_7030);
and U9248 (N_9248,N_7722,N_6858);
nor U9249 (N_9249,N_6333,N_6343);
nand U9250 (N_9250,N_7240,N_7327);
nor U9251 (N_9251,N_7293,N_6486);
nor U9252 (N_9252,N_6752,N_7826);
nand U9253 (N_9253,N_7819,N_7248);
nand U9254 (N_9254,N_6507,N_7243);
nor U9255 (N_9255,N_7154,N_7970);
and U9256 (N_9256,N_6446,N_7666);
nor U9257 (N_9257,N_6200,N_6116);
nor U9258 (N_9258,N_7400,N_7200);
nor U9259 (N_9259,N_7239,N_6407);
and U9260 (N_9260,N_7061,N_7740);
or U9261 (N_9261,N_7977,N_7697);
and U9262 (N_9262,N_7992,N_7780);
nand U9263 (N_9263,N_6248,N_7178);
nor U9264 (N_9264,N_6674,N_6289);
nand U9265 (N_9265,N_6717,N_7709);
nor U9266 (N_9266,N_7135,N_6991);
nor U9267 (N_9267,N_6287,N_7579);
xnor U9268 (N_9268,N_7019,N_7913);
and U9269 (N_9269,N_6608,N_7351);
nor U9270 (N_9270,N_6142,N_6914);
nor U9271 (N_9271,N_7411,N_7957);
xnor U9272 (N_9272,N_7079,N_6202);
and U9273 (N_9273,N_6978,N_7878);
nor U9274 (N_9274,N_7863,N_7548);
and U9275 (N_9275,N_6989,N_6176);
nor U9276 (N_9276,N_6237,N_7928);
or U9277 (N_9277,N_6549,N_6161);
nand U9278 (N_9278,N_7342,N_6786);
and U9279 (N_9279,N_6858,N_6618);
or U9280 (N_9280,N_6155,N_7104);
nand U9281 (N_9281,N_6587,N_7756);
xnor U9282 (N_9282,N_7165,N_6953);
and U9283 (N_9283,N_7416,N_6673);
xor U9284 (N_9284,N_6211,N_7586);
nand U9285 (N_9285,N_6018,N_6782);
nor U9286 (N_9286,N_7613,N_7769);
nor U9287 (N_9287,N_6891,N_6069);
and U9288 (N_9288,N_6884,N_7471);
and U9289 (N_9289,N_6558,N_7164);
nand U9290 (N_9290,N_6307,N_7486);
nor U9291 (N_9291,N_6670,N_7657);
and U9292 (N_9292,N_7688,N_7229);
nor U9293 (N_9293,N_7695,N_6433);
or U9294 (N_9294,N_7754,N_6615);
nor U9295 (N_9295,N_6108,N_7485);
nor U9296 (N_9296,N_6963,N_6878);
nand U9297 (N_9297,N_7066,N_7090);
nor U9298 (N_9298,N_6871,N_7854);
nand U9299 (N_9299,N_7631,N_7357);
nor U9300 (N_9300,N_6426,N_7949);
nor U9301 (N_9301,N_7993,N_7820);
nor U9302 (N_9302,N_7695,N_7472);
and U9303 (N_9303,N_7511,N_6076);
and U9304 (N_9304,N_6603,N_7211);
or U9305 (N_9305,N_7729,N_7360);
nor U9306 (N_9306,N_6073,N_7331);
nand U9307 (N_9307,N_7840,N_6852);
nor U9308 (N_9308,N_7496,N_7704);
or U9309 (N_9309,N_7619,N_7266);
nand U9310 (N_9310,N_7592,N_7193);
or U9311 (N_9311,N_6213,N_6625);
and U9312 (N_9312,N_7722,N_6719);
nand U9313 (N_9313,N_6486,N_7576);
xor U9314 (N_9314,N_6804,N_7470);
nand U9315 (N_9315,N_6230,N_7971);
xor U9316 (N_9316,N_7026,N_7574);
or U9317 (N_9317,N_6425,N_6095);
nand U9318 (N_9318,N_6591,N_6962);
nand U9319 (N_9319,N_7565,N_7795);
or U9320 (N_9320,N_7498,N_6868);
nor U9321 (N_9321,N_7609,N_6045);
or U9322 (N_9322,N_7322,N_6949);
xnor U9323 (N_9323,N_6314,N_6414);
and U9324 (N_9324,N_6674,N_7654);
xnor U9325 (N_9325,N_7657,N_7364);
or U9326 (N_9326,N_6503,N_6691);
or U9327 (N_9327,N_6925,N_6426);
nand U9328 (N_9328,N_6843,N_6229);
and U9329 (N_9329,N_6184,N_7065);
nand U9330 (N_9330,N_7299,N_6175);
and U9331 (N_9331,N_6556,N_6792);
and U9332 (N_9332,N_7468,N_7466);
xor U9333 (N_9333,N_6662,N_6778);
nor U9334 (N_9334,N_7973,N_7558);
nand U9335 (N_9335,N_7401,N_6896);
and U9336 (N_9336,N_7782,N_6525);
xnor U9337 (N_9337,N_6573,N_7248);
nand U9338 (N_9338,N_7170,N_7207);
or U9339 (N_9339,N_6541,N_6006);
and U9340 (N_9340,N_7444,N_7233);
nand U9341 (N_9341,N_7123,N_6451);
nor U9342 (N_9342,N_6078,N_7881);
nor U9343 (N_9343,N_6689,N_7932);
xor U9344 (N_9344,N_7896,N_6722);
xor U9345 (N_9345,N_6208,N_7179);
xor U9346 (N_9346,N_6831,N_7781);
and U9347 (N_9347,N_6694,N_6804);
and U9348 (N_9348,N_6535,N_7415);
nor U9349 (N_9349,N_6091,N_6750);
nor U9350 (N_9350,N_7346,N_7554);
or U9351 (N_9351,N_7059,N_7354);
nand U9352 (N_9352,N_7183,N_6125);
or U9353 (N_9353,N_6975,N_6137);
nor U9354 (N_9354,N_7517,N_7392);
nor U9355 (N_9355,N_6664,N_7646);
or U9356 (N_9356,N_7731,N_7162);
nand U9357 (N_9357,N_6613,N_7293);
xor U9358 (N_9358,N_6112,N_6805);
and U9359 (N_9359,N_6839,N_6623);
and U9360 (N_9360,N_7361,N_7384);
and U9361 (N_9361,N_6234,N_7352);
nor U9362 (N_9362,N_7068,N_7548);
xor U9363 (N_9363,N_7693,N_6471);
nand U9364 (N_9364,N_6374,N_6297);
nor U9365 (N_9365,N_7664,N_7333);
and U9366 (N_9366,N_6110,N_6023);
nor U9367 (N_9367,N_6181,N_6991);
xnor U9368 (N_9368,N_6574,N_7624);
xnor U9369 (N_9369,N_7431,N_6353);
nor U9370 (N_9370,N_7914,N_6306);
or U9371 (N_9371,N_6626,N_6788);
nor U9372 (N_9372,N_7950,N_7172);
and U9373 (N_9373,N_7400,N_7030);
xnor U9374 (N_9374,N_6132,N_6551);
nor U9375 (N_9375,N_6327,N_6540);
nor U9376 (N_9376,N_6388,N_6185);
or U9377 (N_9377,N_7157,N_6619);
nor U9378 (N_9378,N_6257,N_6303);
xor U9379 (N_9379,N_7851,N_6603);
or U9380 (N_9380,N_7759,N_7887);
xnor U9381 (N_9381,N_6308,N_7826);
and U9382 (N_9382,N_7546,N_6782);
nor U9383 (N_9383,N_7419,N_7083);
and U9384 (N_9384,N_7221,N_7582);
xnor U9385 (N_9385,N_7243,N_6016);
or U9386 (N_9386,N_7264,N_7916);
and U9387 (N_9387,N_6715,N_6863);
nand U9388 (N_9388,N_7488,N_6814);
xnor U9389 (N_9389,N_6199,N_7324);
nand U9390 (N_9390,N_7210,N_7963);
xnor U9391 (N_9391,N_6302,N_6041);
xnor U9392 (N_9392,N_6091,N_6720);
or U9393 (N_9393,N_6571,N_7719);
xor U9394 (N_9394,N_6616,N_7486);
and U9395 (N_9395,N_6233,N_7095);
and U9396 (N_9396,N_6993,N_7395);
nand U9397 (N_9397,N_6998,N_7989);
xor U9398 (N_9398,N_7725,N_7428);
nand U9399 (N_9399,N_6158,N_6229);
or U9400 (N_9400,N_6562,N_6651);
xnor U9401 (N_9401,N_7948,N_6244);
nand U9402 (N_9402,N_6263,N_7182);
nor U9403 (N_9403,N_7294,N_6585);
and U9404 (N_9404,N_7190,N_6370);
or U9405 (N_9405,N_6530,N_6744);
and U9406 (N_9406,N_7799,N_7540);
and U9407 (N_9407,N_6852,N_6846);
or U9408 (N_9408,N_6705,N_6479);
nand U9409 (N_9409,N_6600,N_7374);
or U9410 (N_9410,N_6037,N_7626);
nand U9411 (N_9411,N_7627,N_6549);
xnor U9412 (N_9412,N_6098,N_6012);
nor U9413 (N_9413,N_7457,N_6839);
and U9414 (N_9414,N_7807,N_7732);
and U9415 (N_9415,N_6400,N_6801);
or U9416 (N_9416,N_7305,N_6878);
or U9417 (N_9417,N_6419,N_7999);
and U9418 (N_9418,N_6418,N_7223);
or U9419 (N_9419,N_7425,N_7095);
nand U9420 (N_9420,N_6581,N_6761);
xor U9421 (N_9421,N_6268,N_7040);
and U9422 (N_9422,N_6420,N_6943);
and U9423 (N_9423,N_6929,N_7022);
and U9424 (N_9424,N_7191,N_6004);
xnor U9425 (N_9425,N_6895,N_7931);
or U9426 (N_9426,N_6910,N_7819);
or U9427 (N_9427,N_6832,N_7942);
nor U9428 (N_9428,N_7998,N_6734);
nand U9429 (N_9429,N_7218,N_7634);
nor U9430 (N_9430,N_6164,N_7516);
or U9431 (N_9431,N_7000,N_7039);
nand U9432 (N_9432,N_6684,N_7629);
or U9433 (N_9433,N_7975,N_6109);
and U9434 (N_9434,N_6065,N_6047);
nand U9435 (N_9435,N_7491,N_7418);
or U9436 (N_9436,N_6819,N_6590);
xor U9437 (N_9437,N_6101,N_7197);
or U9438 (N_9438,N_7500,N_7507);
and U9439 (N_9439,N_6785,N_7760);
nand U9440 (N_9440,N_7762,N_7633);
nand U9441 (N_9441,N_7807,N_6049);
xnor U9442 (N_9442,N_7335,N_7078);
nand U9443 (N_9443,N_6600,N_7012);
and U9444 (N_9444,N_7960,N_7001);
nor U9445 (N_9445,N_6496,N_6409);
nor U9446 (N_9446,N_6832,N_6707);
xor U9447 (N_9447,N_7688,N_7712);
and U9448 (N_9448,N_7118,N_6489);
and U9449 (N_9449,N_7579,N_7451);
nor U9450 (N_9450,N_6249,N_7288);
and U9451 (N_9451,N_7667,N_7379);
nand U9452 (N_9452,N_6753,N_6817);
nor U9453 (N_9453,N_7394,N_6543);
nand U9454 (N_9454,N_7375,N_7811);
or U9455 (N_9455,N_7740,N_7113);
and U9456 (N_9456,N_6583,N_6256);
nand U9457 (N_9457,N_6618,N_7853);
nand U9458 (N_9458,N_7056,N_7756);
and U9459 (N_9459,N_7153,N_7904);
nor U9460 (N_9460,N_7597,N_7537);
nor U9461 (N_9461,N_7058,N_7406);
xnor U9462 (N_9462,N_7204,N_7865);
xnor U9463 (N_9463,N_6578,N_6598);
nor U9464 (N_9464,N_6182,N_7523);
or U9465 (N_9465,N_6542,N_7349);
xnor U9466 (N_9466,N_7689,N_6873);
xor U9467 (N_9467,N_7251,N_7141);
xor U9468 (N_9468,N_7096,N_7827);
or U9469 (N_9469,N_6747,N_7164);
xnor U9470 (N_9470,N_6618,N_6647);
and U9471 (N_9471,N_6332,N_6520);
nand U9472 (N_9472,N_7649,N_6946);
and U9473 (N_9473,N_6176,N_7103);
xor U9474 (N_9474,N_6099,N_6498);
or U9475 (N_9475,N_6988,N_7141);
or U9476 (N_9476,N_6961,N_7776);
and U9477 (N_9477,N_6329,N_6642);
nor U9478 (N_9478,N_7136,N_7486);
or U9479 (N_9479,N_7420,N_7440);
or U9480 (N_9480,N_7550,N_6974);
or U9481 (N_9481,N_6554,N_7016);
nor U9482 (N_9482,N_7390,N_7887);
nor U9483 (N_9483,N_7910,N_6948);
nor U9484 (N_9484,N_6293,N_7977);
xor U9485 (N_9485,N_7483,N_6328);
nand U9486 (N_9486,N_6188,N_7367);
xor U9487 (N_9487,N_7286,N_7514);
nand U9488 (N_9488,N_6603,N_6905);
nand U9489 (N_9489,N_7479,N_6944);
nand U9490 (N_9490,N_6108,N_7325);
xnor U9491 (N_9491,N_6604,N_7926);
nor U9492 (N_9492,N_7328,N_6380);
nor U9493 (N_9493,N_7243,N_6953);
nand U9494 (N_9494,N_7886,N_7492);
and U9495 (N_9495,N_6983,N_7494);
nor U9496 (N_9496,N_7362,N_6283);
or U9497 (N_9497,N_7860,N_6142);
nor U9498 (N_9498,N_7213,N_6283);
and U9499 (N_9499,N_6387,N_7409);
nand U9500 (N_9500,N_6984,N_7902);
nor U9501 (N_9501,N_7341,N_7256);
xnor U9502 (N_9502,N_7745,N_7175);
xor U9503 (N_9503,N_6221,N_7475);
nor U9504 (N_9504,N_7819,N_6465);
and U9505 (N_9505,N_7346,N_7374);
nand U9506 (N_9506,N_6730,N_6331);
or U9507 (N_9507,N_7972,N_6790);
or U9508 (N_9508,N_7327,N_7324);
or U9509 (N_9509,N_6094,N_7956);
and U9510 (N_9510,N_7292,N_7082);
and U9511 (N_9511,N_6443,N_6261);
xor U9512 (N_9512,N_7103,N_6713);
nor U9513 (N_9513,N_7184,N_6915);
nor U9514 (N_9514,N_7770,N_7557);
nand U9515 (N_9515,N_7239,N_7768);
or U9516 (N_9516,N_7662,N_7709);
xor U9517 (N_9517,N_7815,N_7254);
nand U9518 (N_9518,N_6352,N_7118);
nor U9519 (N_9519,N_6791,N_7897);
nor U9520 (N_9520,N_6834,N_6664);
and U9521 (N_9521,N_7611,N_7409);
xnor U9522 (N_9522,N_7013,N_7800);
and U9523 (N_9523,N_7233,N_7471);
nor U9524 (N_9524,N_6997,N_7748);
or U9525 (N_9525,N_7834,N_7465);
nor U9526 (N_9526,N_6960,N_6655);
xnor U9527 (N_9527,N_6113,N_6408);
and U9528 (N_9528,N_6691,N_6939);
nor U9529 (N_9529,N_7499,N_6308);
and U9530 (N_9530,N_7616,N_7573);
nand U9531 (N_9531,N_6235,N_6422);
nand U9532 (N_9532,N_7694,N_6911);
xnor U9533 (N_9533,N_6291,N_7641);
nand U9534 (N_9534,N_7931,N_6186);
or U9535 (N_9535,N_6276,N_7772);
nand U9536 (N_9536,N_7435,N_7695);
xor U9537 (N_9537,N_6157,N_6247);
and U9538 (N_9538,N_6706,N_7593);
nor U9539 (N_9539,N_7504,N_7626);
and U9540 (N_9540,N_7269,N_6740);
or U9541 (N_9541,N_7109,N_6054);
and U9542 (N_9542,N_6957,N_6409);
nor U9543 (N_9543,N_6995,N_7082);
nor U9544 (N_9544,N_6209,N_7565);
or U9545 (N_9545,N_6036,N_6793);
nand U9546 (N_9546,N_6136,N_6470);
and U9547 (N_9547,N_7432,N_6080);
xnor U9548 (N_9548,N_6228,N_6269);
nor U9549 (N_9549,N_6998,N_7355);
nand U9550 (N_9550,N_6765,N_7655);
nor U9551 (N_9551,N_7645,N_7583);
nand U9552 (N_9552,N_7084,N_7746);
and U9553 (N_9553,N_7836,N_7867);
and U9554 (N_9554,N_7729,N_6021);
or U9555 (N_9555,N_6582,N_7044);
and U9556 (N_9556,N_6885,N_7197);
nor U9557 (N_9557,N_6553,N_7882);
nor U9558 (N_9558,N_7926,N_6365);
nor U9559 (N_9559,N_7068,N_6848);
nor U9560 (N_9560,N_6476,N_7453);
nand U9561 (N_9561,N_6609,N_6039);
or U9562 (N_9562,N_7017,N_7186);
xor U9563 (N_9563,N_7309,N_7895);
nand U9564 (N_9564,N_6112,N_6680);
and U9565 (N_9565,N_6694,N_7465);
xnor U9566 (N_9566,N_6778,N_6129);
nand U9567 (N_9567,N_6288,N_7761);
or U9568 (N_9568,N_6029,N_7521);
and U9569 (N_9569,N_7229,N_7922);
or U9570 (N_9570,N_6381,N_7171);
or U9571 (N_9571,N_7029,N_6250);
nor U9572 (N_9572,N_6845,N_7284);
xnor U9573 (N_9573,N_6564,N_7399);
nand U9574 (N_9574,N_7645,N_6275);
xnor U9575 (N_9575,N_6538,N_6566);
or U9576 (N_9576,N_7222,N_7739);
or U9577 (N_9577,N_6949,N_7659);
and U9578 (N_9578,N_6166,N_6122);
and U9579 (N_9579,N_6852,N_7399);
and U9580 (N_9580,N_6020,N_6362);
and U9581 (N_9581,N_7174,N_7953);
nor U9582 (N_9582,N_6827,N_7065);
xor U9583 (N_9583,N_7409,N_6320);
xnor U9584 (N_9584,N_7288,N_7738);
or U9585 (N_9585,N_6067,N_6211);
nand U9586 (N_9586,N_7966,N_6213);
nand U9587 (N_9587,N_6136,N_6322);
or U9588 (N_9588,N_6980,N_7829);
and U9589 (N_9589,N_7010,N_7102);
nand U9590 (N_9590,N_6557,N_7718);
nor U9591 (N_9591,N_7742,N_7232);
or U9592 (N_9592,N_7917,N_7655);
nand U9593 (N_9593,N_7411,N_7753);
or U9594 (N_9594,N_7849,N_6658);
xor U9595 (N_9595,N_7678,N_7623);
xor U9596 (N_9596,N_7821,N_7324);
xor U9597 (N_9597,N_7848,N_6704);
nand U9598 (N_9598,N_6462,N_6872);
xor U9599 (N_9599,N_6078,N_7412);
nand U9600 (N_9600,N_7853,N_6299);
nand U9601 (N_9601,N_7096,N_6878);
or U9602 (N_9602,N_6112,N_6058);
nand U9603 (N_9603,N_7081,N_7491);
nand U9604 (N_9604,N_7762,N_6413);
and U9605 (N_9605,N_6209,N_7450);
and U9606 (N_9606,N_7709,N_6321);
xor U9607 (N_9607,N_7121,N_6901);
nor U9608 (N_9608,N_7286,N_6185);
and U9609 (N_9609,N_7478,N_7447);
nor U9610 (N_9610,N_6585,N_6134);
xor U9611 (N_9611,N_6475,N_7536);
xor U9612 (N_9612,N_7362,N_6949);
nor U9613 (N_9613,N_6295,N_6456);
nand U9614 (N_9614,N_7843,N_6368);
nor U9615 (N_9615,N_6637,N_6809);
or U9616 (N_9616,N_6933,N_7657);
nand U9617 (N_9617,N_7956,N_6846);
xor U9618 (N_9618,N_7145,N_6842);
or U9619 (N_9619,N_6016,N_7812);
and U9620 (N_9620,N_6193,N_6204);
xnor U9621 (N_9621,N_7555,N_7960);
and U9622 (N_9622,N_6966,N_6565);
or U9623 (N_9623,N_6676,N_7260);
or U9624 (N_9624,N_6381,N_6241);
nand U9625 (N_9625,N_6099,N_6888);
xor U9626 (N_9626,N_6203,N_7163);
nor U9627 (N_9627,N_7879,N_7782);
nand U9628 (N_9628,N_6985,N_7277);
or U9629 (N_9629,N_7629,N_7968);
nor U9630 (N_9630,N_7097,N_7372);
nor U9631 (N_9631,N_7094,N_6239);
and U9632 (N_9632,N_6273,N_6177);
nand U9633 (N_9633,N_7921,N_6846);
or U9634 (N_9634,N_6638,N_7332);
and U9635 (N_9635,N_7839,N_6883);
and U9636 (N_9636,N_6160,N_7457);
xor U9637 (N_9637,N_7337,N_7315);
and U9638 (N_9638,N_7385,N_7903);
and U9639 (N_9639,N_6924,N_6103);
xnor U9640 (N_9640,N_7883,N_7636);
nand U9641 (N_9641,N_7446,N_6056);
and U9642 (N_9642,N_6207,N_7291);
nor U9643 (N_9643,N_7676,N_7218);
or U9644 (N_9644,N_6247,N_7468);
or U9645 (N_9645,N_7622,N_7508);
nand U9646 (N_9646,N_7639,N_6600);
nand U9647 (N_9647,N_6675,N_6421);
or U9648 (N_9648,N_6904,N_7499);
or U9649 (N_9649,N_6234,N_7080);
xor U9650 (N_9650,N_7502,N_6159);
or U9651 (N_9651,N_6648,N_7053);
xnor U9652 (N_9652,N_7383,N_6386);
nand U9653 (N_9653,N_7117,N_7855);
and U9654 (N_9654,N_6596,N_6443);
nand U9655 (N_9655,N_6239,N_7003);
nor U9656 (N_9656,N_7532,N_6409);
and U9657 (N_9657,N_6442,N_6101);
or U9658 (N_9658,N_7927,N_6634);
and U9659 (N_9659,N_6023,N_6875);
and U9660 (N_9660,N_6438,N_7003);
or U9661 (N_9661,N_6560,N_7670);
or U9662 (N_9662,N_7345,N_7875);
or U9663 (N_9663,N_6657,N_7772);
or U9664 (N_9664,N_6207,N_6577);
or U9665 (N_9665,N_6953,N_7876);
nor U9666 (N_9666,N_6606,N_6526);
xnor U9667 (N_9667,N_6064,N_7958);
nand U9668 (N_9668,N_7707,N_7545);
nor U9669 (N_9669,N_6797,N_7176);
or U9670 (N_9670,N_6833,N_7722);
xor U9671 (N_9671,N_7988,N_7722);
or U9672 (N_9672,N_7462,N_7303);
nor U9673 (N_9673,N_6958,N_6739);
and U9674 (N_9674,N_7043,N_6623);
xnor U9675 (N_9675,N_6869,N_6808);
nor U9676 (N_9676,N_7876,N_6268);
or U9677 (N_9677,N_7613,N_6198);
xnor U9678 (N_9678,N_7642,N_6133);
and U9679 (N_9679,N_7267,N_7694);
and U9680 (N_9680,N_7210,N_6114);
and U9681 (N_9681,N_6128,N_7825);
xor U9682 (N_9682,N_6533,N_6926);
nor U9683 (N_9683,N_7124,N_6231);
or U9684 (N_9684,N_6563,N_7565);
nand U9685 (N_9685,N_6877,N_7662);
or U9686 (N_9686,N_6429,N_6514);
xnor U9687 (N_9687,N_6165,N_7428);
xor U9688 (N_9688,N_7187,N_7672);
nand U9689 (N_9689,N_6298,N_7253);
and U9690 (N_9690,N_6163,N_6740);
xnor U9691 (N_9691,N_6703,N_6360);
nor U9692 (N_9692,N_6682,N_6470);
and U9693 (N_9693,N_6134,N_6430);
or U9694 (N_9694,N_6965,N_6749);
or U9695 (N_9695,N_6600,N_6213);
and U9696 (N_9696,N_7913,N_7724);
nand U9697 (N_9697,N_7106,N_7921);
and U9698 (N_9698,N_6403,N_7472);
xor U9699 (N_9699,N_6108,N_6391);
nand U9700 (N_9700,N_6430,N_6713);
and U9701 (N_9701,N_7525,N_6782);
nand U9702 (N_9702,N_7999,N_7277);
and U9703 (N_9703,N_6827,N_6058);
xor U9704 (N_9704,N_6584,N_6503);
xnor U9705 (N_9705,N_7459,N_6776);
and U9706 (N_9706,N_7152,N_7825);
and U9707 (N_9707,N_7223,N_7018);
and U9708 (N_9708,N_7842,N_7584);
nor U9709 (N_9709,N_7784,N_6089);
xor U9710 (N_9710,N_6116,N_6797);
or U9711 (N_9711,N_6355,N_7785);
and U9712 (N_9712,N_6331,N_7242);
nand U9713 (N_9713,N_6384,N_6617);
or U9714 (N_9714,N_7085,N_6936);
nor U9715 (N_9715,N_6890,N_7953);
nand U9716 (N_9716,N_6591,N_6785);
xor U9717 (N_9717,N_7687,N_6760);
and U9718 (N_9718,N_6401,N_7115);
and U9719 (N_9719,N_7035,N_7929);
xor U9720 (N_9720,N_6692,N_7513);
and U9721 (N_9721,N_7386,N_6729);
nor U9722 (N_9722,N_7239,N_6863);
nor U9723 (N_9723,N_7331,N_6142);
nand U9724 (N_9724,N_6734,N_7428);
and U9725 (N_9725,N_6010,N_7268);
xor U9726 (N_9726,N_7352,N_7248);
or U9727 (N_9727,N_6046,N_7182);
and U9728 (N_9728,N_6298,N_7543);
or U9729 (N_9729,N_6974,N_6945);
or U9730 (N_9730,N_6999,N_7862);
or U9731 (N_9731,N_7380,N_7152);
nand U9732 (N_9732,N_7986,N_6183);
xnor U9733 (N_9733,N_7025,N_7057);
and U9734 (N_9734,N_6175,N_7327);
and U9735 (N_9735,N_6752,N_6796);
nand U9736 (N_9736,N_6215,N_7711);
xnor U9737 (N_9737,N_6455,N_6139);
and U9738 (N_9738,N_6859,N_7859);
xnor U9739 (N_9739,N_6317,N_6000);
nand U9740 (N_9740,N_6716,N_7027);
nor U9741 (N_9741,N_6881,N_7128);
nor U9742 (N_9742,N_7912,N_6386);
xnor U9743 (N_9743,N_7155,N_7163);
nor U9744 (N_9744,N_7026,N_6153);
nor U9745 (N_9745,N_6960,N_7998);
and U9746 (N_9746,N_6232,N_7762);
nor U9747 (N_9747,N_6411,N_7741);
or U9748 (N_9748,N_6839,N_7942);
and U9749 (N_9749,N_7432,N_7509);
nand U9750 (N_9750,N_6729,N_6632);
or U9751 (N_9751,N_6795,N_6164);
nand U9752 (N_9752,N_7785,N_7815);
xor U9753 (N_9753,N_7487,N_7003);
or U9754 (N_9754,N_6871,N_6511);
xnor U9755 (N_9755,N_7978,N_6813);
xnor U9756 (N_9756,N_7234,N_6028);
nand U9757 (N_9757,N_6768,N_7230);
nand U9758 (N_9758,N_6531,N_7008);
and U9759 (N_9759,N_6618,N_7049);
nor U9760 (N_9760,N_7048,N_6813);
nand U9761 (N_9761,N_7157,N_7757);
nand U9762 (N_9762,N_6341,N_7182);
nor U9763 (N_9763,N_6027,N_6688);
nand U9764 (N_9764,N_7510,N_6982);
nand U9765 (N_9765,N_6141,N_7760);
or U9766 (N_9766,N_7147,N_6941);
and U9767 (N_9767,N_7124,N_6241);
nand U9768 (N_9768,N_7270,N_6663);
and U9769 (N_9769,N_7451,N_7424);
and U9770 (N_9770,N_7734,N_6031);
nand U9771 (N_9771,N_7241,N_6987);
and U9772 (N_9772,N_7905,N_7674);
and U9773 (N_9773,N_7586,N_6227);
and U9774 (N_9774,N_6090,N_7080);
nand U9775 (N_9775,N_7870,N_7205);
nor U9776 (N_9776,N_6287,N_7330);
xor U9777 (N_9777,N_7293,N_6829);
xor U9778 (N_9778,N_7932,N_6948);
and U9779 (N_9779,N_7861,N_6563);
or U9780 (N_9780,N_7404,N_7704);
or U9781 (N_9781,N_7271,N_7533);
xor U9782 (N_9782,N_6372,N_6016);
xor U9783 (N_9783,N_7299,N_7490);
and U9784 (N_9784,N_6844,N_7245);
and U9785 (N_9785,N_7501,N_6205);
nand U9786 (N_9786,N_6768,N_6803);
xnor U9787 (N_9787,N_7574,N_6873);
nand U9788 (N_9788,N_7432,N_7436);
or U9789 (N_9789,N_6842,N_7982);
and U9790 (N_9790,N_7094,N_6073);
and U9791 (N_9791,N_7350,N_7933);
and U9792 (N_9792,N_6685,N_6540);
and U9793 (N_9793,N_6542,N_7225);
or U9794 (N_9794,N_7326,N_7273);
xor U9795 (N_9795,N_7192,N_6342);
nor U9796 (N_9796,N_7708,N_6091);
and U9797 (N_9797,N_7674,N_6109);
nand U9798 (N_9798,N_6440,N_6821);
and U9799 (N_9799,N_7252,N_7957);
and U9800 (N_9800,N_6789,N_7529);
nor U9801 (N_9801,N_6190,N_6451);
nor U9802 (N_9802,N_6461,N_6219);
and U9803 (N_9803,N_7664,N_6968);
nor U9804 (N_9804,N_6941,N_6965);
nor U9805 (N_9805,N_6966,N_6702);
nor U9806 (N_9806,N_6844,N_7500);
nand U9807 (N_9807,N_6567,N_7984);
or U9808 (N_9808,N_7311,N_6165);
or U9809 (N_9809,N_6923,N_6786);
nor U9810 (N_9810,N_6904,N_7745);
nand U9811 (N_9811,N_6485,N_7762);
nand U9812 (N_9812,N_6895,N_7143);
xnor U9813 (N_9813,N_7080,N_6363);
or U9814 (N_9814,N_6432,N_6135);
and U9815 (N_9815,N_6395,N_6724);
nand U9816 (N_9816,N_6548,N_6876);
nor U9817 (N_9817,N_7310,N_6105);
nand U9818 (N_9818,N_7227,N_7390);
xor U9819 (N_9819,N_6993,N_6774);
xnor U9820 (N_9820,N_6708,N_6692);
nand U9821 (N_9821,N_6917,N_7131);
xnor U9822 (N_9822,N_6324,N_6719);
and U9823 (N_9823,N_6014,N_7941);
or U9824 (N_9824,N_6394,N_6954);
and U9825 (N_9825,N_7949,N_6345);
nor U9826 (N_9826,N_6704,N_7047);
or U9827 (N_9827,N_6348,N_6516);
nand U9828 (N_9828,N_7679,N_7189);
and U9829 (N_9829,N_6430,N_6445);
nand U9830 (N_9830,N_7852,N_7060);
xor U9831 (N_9831,N_6903,N_6562);
nand U9832 (N_9832,N_7550,N_7621);
or U9833 (N_9833,N_7294,N_7398);
nand U9834 (N_9834,N_6438,N_7348);
and U9835 (N_9835,N_7068,N_7185);
and U9836 (N_9836,N_6625,N_6273);
nor U9837 (N_9837,N_6070,N_7391);
nor U9838 (N_9838,N_6888,N_6874);
nor U9839 (N_9839,N_7597,N_6857);
nand U9840 (N_9840,N_7941,N_6741);
nand U9841 (N_9841,N_6058,N_6845);
or U9842 (N_9842,N_6137,N_6449);
and U9843 (N_9843,N_7648,N_6460);
or U9844 (N_9844,N_7767,N_7436);
xor U9845 (N_9845,N_7335,N_7336);
nand U9846 (N_9846,N_7368,N_6258);
nor U9847 (N_9847,N_7660,N_6944);
or U9848 (N_9848,N_7767,N_6395);
nand U9849 (N_9849,N_6583,N_6414);
nand U9850 (N_9850,N_6719,N_6472);
xnor U9851 (N_9851,N_7494,N_6112);
or U9852 (N_9852,N_7695,N_7970);
nand U9853 (N_9853,N_6106,N_7349);
xor U9854 (N_9854,N_6082,N_7363);
and U9855 (N_9855,N_6560,N_6343);
nand U9856 (N_9856,N_7634,N_7204);
nor U9857 (N_9857,N_6312,N_6600);
or U9858 (N_9858,N_6429,N_6765);
nor U9859 (N_9859,N_6137,N_6933);
or U9860 (N_9860,N_6130,N_7395);
or U9861 (N_9861,N_6590,N_7785);
and U9862 (N_9862,N_7193,N_7208);
and U9863 (N_9863,N_7570,N_7485);
nor U9864 (N_9864,N_6102,N_7234);
nand U9865 (N_9865,N_6874,N_7364);
xnor U9866 (N_9866,N_7496,N_6912);
and U9867 (N_9867,N_6917,N_6816);
xor U9868 (N_9868,N_7592,N_7845);
and U9869 (N_9869,N_7740,N_7493);
and U9870 (N_9870,N_7446,N_6418);
and U9871 (N_9871,N_7540,N_6863);
or U9872 (N_9872,N_6099,N_6014);
and U9873 (N_9873,N_7993,N_6334);
nand U9874 (N_9874,N_6222,N_6751);
nor U9875 (N_9875,N_6590,N_7756);
nand U9876 (N_9876,N_7977,N_7796);
nor U9877 (N_9877,N_7023,N_6826);
nor U9878 (N_9878,N_6535,N_7189);
xnor U9879 (N_9879,N_6844,N_7655);
nor U9880 (N_9880,N_7131,N_6584);
and U9881 (N_9881,N_7347,N_6745);
or U9882 (N_9882,N_7536,N_7291);
xor U9883 (N_9883,N_6960,N_7188);
or U9884 (N_9884,N_6213,N_7747);
nor U9885 (N_9885,N_7775,N_7373);
xnor U9886 (N_9886,N_6403,N_7097);
nor U9887 (N_9887,N_7784,N_7038);
and U9888 (N_9888,N_7781,N_7683);
nand U9889 (N_9889,N_6640,N_7550);
xnor U9890 (N_9890,N_7072,N_7597);
xnor U9891 (N_9891,N_7914,N_7082);
xor U9892 (N_9892,N_6747,N_6660);
xor U9893 (N_9893,N_7506,N_6832);
nor U9894 (N_9894,N_7839,N_7174);
nor U9895 (N_9895,N_6472,N_6242);
nor U9896 (N_9896,N_7489,N_7663);
xor U9897 (N_9897,N_6234,N_6968);
nand U9898 (N_9898,N_6498,N_6691);
and U9899 (N_9899,N_6022,N_7749);
nor U9900 (N_9900,N_7723,N_6088);
nand U9901 (N_9901,N_7091,N_6689);
xnor U9902 (N_9902,N_7111,N_6895);
and U9903 (N_9903,N_6429,N_6566);
nand U9904 (N_9904,N_6393,N_7310);
and U9905 (N_9905,N_6962,N_7320);
and U9906 (N_9906,N_7923,N_7043);
xor U9907 (N_9907,N_6899,N_6191);
nand U9908 (N_9908,N_7115,N_7886);
xor U9909 (N_9909,N_7804,N_7600);
or U9910 (N_9910,N_7457,N_7221);
xnor U9911 (N_9911,N_6239,N_6309);
nor U9912 (N_9912,N_6501,N_6439);
and U9913 (N_9913,N_7765,N_6442);
nor U9914 (N_9914,N_6830,N_7358);
nor U9915 (N_9915,N_6703,N_6655);
xnor U9916 (N_9916,N_7687,N_6880);
or U9917 (N_9917,N_6616,N_7858);
nor U9918 (N_9918,N_6712,N_7221);
or U9919 (N_9919,N_7557,N_6202);
or U9920 (N_9920,N_7645,N_7717);
and U9921 (N_9921,N_7797,N_6737);
and U9922 (N_9922,N_6451,N_6264);
nor U9923 (N_9923,N_7517,N_6655);
and U9924 (N_9924,N_6406,N_7522);
or U9925 (N_9925,N_7633,N_6397);
and U9926 (N_9926,N_7064,N_6593);
or U9927 (N_9927,N_7261,N_6522);
nand U9928 (N_9928,N_6246,N_7697);
nor U9929 (N_9929,N_6061,N_7528);
or U9930 (N_9930,N_7767,N_6906);
and U9931 (N_9931,N_6533,N_7394);
and U9932 (N_9932,N_6955,N_6472);
or U9933 (N_9933,N_7656,N_7088);
nand U9934 (N_9934,N_6366,N_6086);
xnor U9935 (N_9935,N_6025,N_6977);
nand U9936 (N_9936,N_7107,N_7397);
or U9937 (N_9937,N_6831,N_6024);
or U9938 (N_9938,N_7307,N_6549);
nand U9939 (N_9939,N_7247,N_7258);
xor U9940 (N_9940,N_7246,N_6475);
nor U9941 (N_9941,N_7907,N_6295);
nand U9942 (N_9942,N_7045,N_6584);
or U9943 (N_9943,N_6397,N_6042);
nor U9944 (N_9944,N_6228,N_6372);
nand U9945 (N_9945,N_6490,N_7462);
xor U9946 (N_9946,N_7142,N_6406);
or U9947 (N_9947,N_7047,N_6635);
or U9948 (N_9948,N_6245,N_6548);
and U9949 (N_9949,N_7187,N_6955);
and U9950 (N_9950,N_6653,N_6918);
nand U9951 (N_9951,N_6773,N_7907);
nor U9952 (N_9952,N_6033,N_6752);
or U9953 (N_9953,N_7987,N_6578);
or U9954 (N_9954,N_6796,N_7831);
and U9955 (N_9955,N_6474,N_7942);
nor U9956 (N_9956,N_7321,N_7673);
or U9957 (N_9957,N_7517,N_7814);
or U9958 (N_9958,N_6018,N_7791);
nand U9959 (N_9959,N_7404,N_6198);
xor U9960 (N_9960,N_6407,N_6569);
or U9961 (N_9961,N_7974,N_6395);
xnor U9962 (N_9962,N_7662,N_7968);
and U9963 (N_9963,N_6747,N_6188);
xor U9964 (N_9964,N_7411,N_6972);
xor U9965 (N_9965,N_6404,N_7638);
xor U9966 (N_9966,N_6035,N_7517);
xnor U9967 (N_9967,N_6041,N_7087);
nand U9968 (N_9968,N_7719,N_7847);
nand U9969 (N_9969,N_6988,N_7274);
nor U9970 (N_9970,N_7427,N_7857);
nor U9971 (N_9971,N_7364,N_7348);
nand U9972 (N_9972,N_7003,N_6727);
and U9973 (N_9973,N_7208,N_6525);
or U9974 (N_9974,N_6181,N_6398);
nor U9975 (N_9975,N_6516,N_6373);
and U9976 (N_9976,N_6744,N_7012);
xnor U9977 (N_9977,N_6332,N_7356);
and U9978 (N_9978,N_7542,N_7188);
and U9979 (N_9979,N_6637,N_7929);
nor U9980 (N_9980,N_7106,N_6520);
nor U9981 (N_9981,N_6401,N_6667);
and U9982 (N_9982,N_7354,N_7052);
xor U9983 (N_9983,N_6025,N_6133);
nor U9984 (N_9984,N_6428,N_7987);
and U9985 (N_9985,N_6911,N_7691);
xnor U9986 (N_9986,N_6543,N_7456);
and U9987 (N_9987,N_7572,N_6400);
xor U9988 (N_9988,N_6130,N_7021);
and U9989 (N_9989,N_6921,N_7452);
nor U9990 (N_9990,N_6907,N_6515);
nand U9991 (N_9991,N_6256,N_6160);
nor U9992 (N_9992,N_7157,N_6328);
nor U9993 (N_9993,N_7870,N_6772);
xnor U9994 (N_9994,N_6214,N_6142);
and U9995 (N_9995,N_7327,N_6784);
nand U9996 (N_9996,N_7431,N_7914);
nand U9997 (N_9997,N_6228,N_7775);
xnor U9998 (N_9998,N_6429,N_6945);
xor U9999 (N_9999,N_7918,N_6287);
xor U10000 (N_10000,N_9455,N_8611);
nand U10001 (N_10001,N_9881,N_9832);
nor U10002 (N_10002,N_9748,N_8005);
xor U10003 (N_10003,N_9260,N_9936);
nand U10004 (N_10004,N_9271,N_8038);
nor U10005 (N_10005,N_8167,N_8511);
nand U10006 (N_10006,N_9988,N_8693);
or U10007 (N_10007,N_9266,N_9813);
nand U10008 (N_10008,N_8116,N_9328);
nand U10009 (N_10009,N_9002,N_9851);
nor U10010 (N_10010,N_9032,N_9931);
or U10011 (N_10011,N_9450,N_9010);
xor U10012 (N_10012,N_8315,N_9040);
nand U10013 (N_10013,N_8425,N_9990);
nor U10014 (N_10014,N_9318,N_9131);
xnor U10015 (N_10015,N_8615,N_8781);
xnor U10016 (N_10016,N_9740,N_8719);
and U10017 (N_10017,N_8412,N_9322);
and U10018 (N_10018,N_9289,N_8861);
nand U10019 (N_10019,N_9228,N_8322);
nor U10020 (N_10020,N_8193,N_8572);
nand U10021 (N_10021,N_8902,N_8003);
nor U10022 (N_10022,N_8512,N_8788);
nand U10023 (N_10023,N_9900,N_8605);
xor U10024 (N_10024,N_8879,N_8523);
nor U10025 (N_10025,N_8629,N_9980);
xor U10026 (N_10026,N_9241,N_9841);
xnor U10027 (N_10027,N_8330,N_8585);
or U10028 (N_10028,N_9685,N_8077);
nor U10029 (N_10029,N_9071,N_9247);
xor U10030 (N_10030,N_8667,N_9424);
xor U10031 (N_10031,N_8048,N_8524);
or U10032 (N_10032,N_9155,N_8111);
and U10033 (N_10033,N_8503,N_8892);
nor U10034 (N_10034,N_9970,N_8303);
nor U10035 (N_10035,N_8718,N_8215);
nand U10036 (N_10036,N_8029,N_8906);
nand U10037 (N_10037,N_9300,N_9205);
and U10038 (N_10038,N_8026,N_8784);
or U10039 (N_10039,N_8098,N_8969);
or U10040 (N_10040,N_9188,N_9705);
or U10041 (N_10041,N_8008,N_8117);
and U10042 (N_10042,N_9103,N_8327);
nand U10043 (N_10043,N_9817,N_8817);
or U10044 (N_10044,N_8390,N_9622);
or U10045 (N_10045,N_9839,N_9068);
and U10046 (N_10046,N_9716,N_9430);
nor U10047 (N_10047,N_8610,N_8494);
and U10048 (N_10048,N_9320,N_8772);
nand U10049 (N_10049,N_8378,N_8289);
or U10050 (N_10050,N_8483,N_8741);
nor U10051 (N_10051,N_9976,N_8086);
xor U10052 (N_10052,N_9274,N_8314);
or U10053 (N_10053,N_8006,N_9476);
xnor U10054 (N_10054,N_8721,N_9079);
and U10055 (N_10055,N_8326,N_9466);
nand U10056 (N_10056,N_8195,N_9122);
or U10057 (N_10057,N_9711,N_9303);
and U10058 (N_10058,N_9855,N_8963);
nand U10059 (N_10059,N_8368,N_9761);
xor U10060 (N_10060,N_9550,N_9845);
and U10061 (N_10061,N_8044,N_8183);
or U10062 (N_10062,N_8847,N_9655);
xor U10063 (N_10063,N_8675,N_9077);
nor U10064 (N_10064,N_9235,N_8119);
nor U10065 (N_10065,N_9779,N_9911);
xnor U10066 (N_10066,N_9145,N_9333);
xnor U10067 (N_10067,N_9408,N_9072);
nand U10068 (N_10068,N_9771,N_9517);
nand U10069 (N_10069,N_9882,N_8220);
nor U10070 (N_10070,N_8934,N_9887);
or U10071 (N_10071,N_9059,N_9651);
nor U10072 (N_10072,N_8375,N_9793);
xnor U10073 (N_10073,N_8915,N_9116);
or U10074 (N_10074,N_8544,N_8971);
nand U10075 (N_10075,N_8826,N_8468);
or U10076 (N_10076,N_9947,N_8956);
and U10077 (N_10077,N_9600,N_9258);
or U10078 (N_10078,N_8185,N_8261);
nor U10079 (N_10079,N_9799,N_8932);
or U10080 (N_10080,N_9297,N_9073);
xnor U10081 (N_10081,N_9594,N_8304);
nand U10082 (N_10082,N_8133,N_8809);
nand U10083 (N_10083,N_8489,N_9843);
xnor U10084 (N_10084,N_9050,N_9286);
or U10085 (N_10085,N_9733,N_9764);
nor U10086 (N_10086,N_8241,N_9309);
or U10087 (N_10087,N_9330,N_9807);
nor U10088 (N_10088,N_8866,N_9162);
and U10089 (N_10089,N_9509,N_8361);
nand U10090 (N_10090,N_8992,N_9618);
nor U10091 (N_10091,N_8914,N_9027);
xor U10092 (N_10092,N_9663,N_8701);
xnor U10093 (N_10093,N_8131,N_8991);
nor U10094 (N_10094,N_9080,N_8886);
or U10095 (N_10095,N_9569,N_9730);
xnor U10096 (N_10096,N_9499,N_9680);
or U10097 (N_10097,N_8064,N_9113);
xnor U10098 (N_10098,N_9387,N_8568);
or U10099 (N_10099,N_8001,N_9662);
nand U10100 (N_10100,N_8025,N_9511);
nand U10101 (N_10101,N_9780,N_9454);
nor U10102 (N_10102,N_9969,N_9206);
or U10103 (N_10103,N_9270,N_8296);
nand U10104 (N_10104,N_9405,N_9874);
nor U10105 (N_10105,N_9777,N_9507);
nor U10106 (N_10106,N_8706,N_9323);
nand U10107 (N_10107,N_9042,N_8834);
nand U10108 (N_10108,N_8732,N_8125);
xor U10109 (N_10109,N_8715,N_9446);
and U10110 (N_10110,N_9496,N_9060);
nor U10111 (N_10111,N_9383,N_9488);
nor U10112 (N_10112,N_8587,N_8273);
and U10113 (N_10113,N_9642,N_9821);
or U10114 (N_10114,N_8597,N_9223);
nand U10115 (N_10115,N_8050,N_9391);
and U10116 (N_10116,N_9413,N_9175);
or U10117 (N_10117,N_8299,N_9472);
nand U10118 (N_10118,N_9802,N_9789);
xor U10119 (N_10119,N_8197,N_9182);
and U10120 (N_10120,N_9835,N_8310);
nor U10121 (N_10121,N_8609,N_9142);
or U10122 (N_10122,N_8118,N_8663);
nor U10123 (N_10123,N_8940,N_8030);
and U10124 (N_10124,N_8600,N_8281);
nand U10125 (N_10125,N_8164,N_8759);
or U10126 (N_10126,N_9571,N_9935);
xnor U10127 (N_10127,N_9406,N_9197);
nor U10128 (N_10128,N_8067,N_8104);
nand U10129 (N_10129,N_8716,N_9232);
nor U10130 (N_10130,N_8399,N_9867);
or U10131 (N_10131,N_8175,N_8893);
nor U10132 (N_10132,N_8516,N_9313);
nand U10133 (N_10133,N_9301,N_9461);
nor U10134 (N_10134,N_9443,N_9484);
xor U10135 (N_10135,N_9973,N_9012);
nor U10136 (N_10136,N_9453,N_9778);
nor U10137 (N_10137,N_8520,N_8336);
xor U10138 (N_10138,N_8124,N_8618);
and U10139 (N_10139,N_9132,N_8564);
nand U10140 (N_10140,N_9146,N_8577);
nand U10141 (N_10141,N_8152,N_9880);
and U10142 (N_10142,N_9026,N_9772);
nand U10143 (N_10143,N_9553,N_9918);
or U10144 (N_10144,N_9008,N_9902);
nor U10145 (N_10145,N_8002,N_8205);
nor U10146 (N_10146,N_8224,N_8981);
or U10147 (N_10147,N_8946,N_9372);
or U10148 (N_10148,N_9619,N_9017);
xnor U10149 (N_10149,N_8422,N_9833);
nor U10150 (N_10150,N_8084,N_9883);
and U10151 (N_10151,N_8232,N_9910);
or U10152 (N_10152,N_9563,N_9515);
nor U10153 (N_10153,N_9785,N_9668);
nand U10154 (N_10154,N_9808,N_9554);
xor U10155 (N_10155,N_8376,N_9321);
nand U10156 (N_10156,N_8669,N_9677);
or U10157 (N_10157,N_9204,N_8009);
nand U10158 (N_10158,N_8628,N_9334);
xnor U10159 (N_10159,N_9127,N_8821);
xor U10160 (N_10160,N_8911,N_9312);
nand U10161 (N_10161,N_9107,N_8080);
xor U10162 (N_10162,N_9991,N_8773);
xor U10163 (N_10163,N_9643,N_8710);
nand U10164 (N_10164,N_9720,N_9277);
xnor U10165 (N_10165,N_8441,N_8022);
xor U10166 (N_10166,N_9912,N_9997);
nor U10167 (N_10167,N_9719,N_9064);
nand U10168 (N_10168,N_8952,N_8749);
and U10169 (N_10169,N_9279,N_8907);
or U10170 (N_10170,N_9775,N_9884);
nand U10171 (N_10171,N_8360,N_8181);
xor U10172 (N_10172,N_9056,N_9745);
nor U10173 (N_10173,N_8582,N_8043);
nor U10174 (N_10174,N_8603,N_8862);
xor U10175 (N_10175,N_9921,N_9765);
nor U10176 (N_10176,N_8411,N_8332);
and U10177 (N_10177,N_9061,N_8988);
and U10178 (N_10178,N_8499,N_9036);
and U10179 (N_10179,N_8871,N_9471);
and U10180 (N_10180,N_9653,N_8632);
nand U10181 (N_10181,N_9169,N_8196);
and U10182 (N_10182,N_9513,N_9192);
and U10183 (N_10183,N_8606,N_9539);
xnor U10184 (N_10184,N_8823,N_8836);
or U10185 (N_10185,N_8254,N_8062);
xnor U10186 (N_10186,N_8127,N_8015);
and U10187 (N_10187,N_8987,N_8623);
or U10188 (N_10188,N_9411,N_8756);
nor U10189 (N_10189,N_9996,N_8820);
nand U10190 (N_10190,N_8334,N_8042);
and U10191 (N_10191,N_8534,N_9019);
nor U10192 (N_10192,N_8157,N_8073);
nand U10193 (N_10193,N_8631,N_8135);
and U10194 (N_10194,N_9822,N_9304);
nor U10195 (N_10195,N_8211,N_8941);
nand U10196 (N_10196,N_8153,N_8931);
or U10197 (N_10197,N_8055,N_9806);
xnor U10198 (N_10198,N_8791,N_9093);
nor U10199 (N_10199,N_8769,N_9152);
nand U10200 (N_10200,N_8673,N_8704);
and U10201 (N_10201,N_8621,N_8156);
xor U10202 (N_10202,N_8364,N_8839);
nand U10203 (N_10203,N_8919,N_9216);
or U10204 (N_10204,N_9287,N_9731);
xor U10205 (N_10205,N_9220,N_9331);
xnor U10206 (N_10206,N_9546,N_8770);
xor U10207 (N_10207,N_8350,N_8060);
nand U10208 (N_10208,N_8052,N_8757);
and U10209 (N_10209,N_8689,N_8264);
and U10210 (N_10210,N_9082,N_9034);
xor U10211 (N_10211,N_8213,N_8172);
and U10212 (N_10212,N_8801,N_8226);
or U10213 (N_10213,N_8640,N_8394);
nor U10214 (N_10214,N_9623,N_8855);
nor U10215 (N_10215,N_9370,N_9746);
nor U10216 (N_10216,N_9664,N_9028);
nor U10217 (N_10217,N_8506,N_9696);
nand U10218 (N_10218,N_8695,N_9830);
nor U10219 (N_10219,N_9459,N_8904);
nor U10220 (N_10220,N_9596,N_8380);
xnor U10221 (N_10221,N_8094,N_8272);
nor U10222 (N_10222,N_8276,N_9015);
or U10223 (N_10223,N_8647,N_8451);
nor U10224 (N_10224,N_8546,N_9528);
xnor U10225 (N_10225,N_9246,N_8837);
or U10226 (N_10226,N_9753,N_9092);
or U10227 (N_10227,N_8790,N_8727);
nand U10228 (N_10228,N_8678,N_9578);
and U10229 (N_10229,N_9626,N_9657);
xnor U10230 (N_10230,N_8184,N_8484);
and U10231 (N_10231,N_9041,N_8918);
nor U10232 (N_10232,N_9491,N_8194);
nor U10233 (N_10233,N_9295,N_9979);
xnor U10234 (N_10234,N_9535,N_9909);
nand U10235 (N_10235,N_9347,N_9354);
or U10236 (N_10236,N_8819,N_8320);
nand U10237 (N_10237,N_9603,N_9847);
nand U10238 (N_10238,N_9311,N_8461);
or U10239 (N_10239,N_9441,N_9009);
xnor U10240 (N_10240,N_9003,N_9234);
nor U10241 (N_10241,N_8528,N_8301);
nor U10242 (N_10242,N_9429,N_8537);
nor U10243 (N_10243,N_8027,N_9972);
and U10244 (N_10244,N_8795,N_9757);
and U10245 (N_10245,N_8702,N_8259);
nor U10246 (N_10246,N_8216,N_9704);
or U10247 (N_10247,N_8723,N_9742);
and U10248 (N_10248,N_8517,N_8056);
or U10249 (N_10249,N_9203,N_8341);
nand U10250 (N_10250,N_9613,N_9736);
or U10251 (N_10251,N_8011,N_9726);
xnor U10252 (N_10252,N_9358,N_8711);
and U10253 (N_10253,N_9269,N_9872);
and U10254 (N_10254,N_8308,N_8481);
xor U10255 (N_10255,N_9097,N_8527);
xnor U10256 (N_10256,N_9126,N_9302);
and U10257 (N_10257,N_9683,N_9776);
nor U10258 (N_10258,N_8717,N_8804);
xor U10259 (N_10259,N_8671,N_8171);
and U10260 (N_10260,N_8031,N_9315);
nand U10261 (N_10261,N_8400,N_9708);
nor U10262 (N_10262,N_9434,N_9389);
xor U10263 (N_10263,N_9635,N_8613);
or U10264 (N_10264,N_9467,N_9904);
nand U10265 (N_10265,N_8265,N_8087);
or U10266 (N_10266,N_8140,N_8901);
and U10267 (N_10267,N_8649,N_8426);
or U10268 (N_10268,N_9219,N_8943);
or U10269 (N_10269,N_9282,N_9352);
nand U10270 (N_10270,N_9095,N_8730);
and U10271 (N_10271,N_9656,N_8746);
xor U10272 (N_10272,N_9209,N_8782);
and U10273 (N_10273,N_9157,N_8852);
or U10274 (N_10274,N_8463,N_9862);
xnor U10275 (N_10275,N_9148,N_8446);
xnor U10276 (N_10276,N_8720,N_8707);
and U10277 (N_10277,N_8382,N_8256);
or U10278 (N_10278,N_9575,N_8559);
or U10279 (N_10279,N_9795,N_8436);
nand U10280 (N_10280,N_9572,N_9689);
or U10281 (N_10281,N_9964,N_9725);
and U10282 (N_10282,N_9280,N_9549);
or U10283 (N_10283,N_8251,N_8342);
and U10284 (N_10284,N_9185,N_8173);
or U10285 (N_10285,N_8571,N_8287);
or U10286 (N_10286,N_9150,N_8604);
nor U10287 (N_10287,N_8432,N_8046);
xnor U10288 (N_10288,N_8557,N_9831);
xnor U10289 (N_10289,N_8177,N_8305);
or U10290 (N_10290,N_9426,N_9410);
nand U10291 (N_10291,N_9005,N_9285);
and U10292 (N_10292,N_8561,N_9512);
xor U10293 (N_10293,N_9350,N_8404);
nor U10294 (N_10294,N_8225,N_8986);
or U10295 (N_10295,N_8085,N_9013);
and U10296 (N_10296,N_8555,N_8169);
and U10297 (N_10297,N_8724,N_9161);
nor U10298 (N_10298,N_9500,N_9633);
and U10299 (N_10299,N_9977,N_9458);
or U10300 (N_10300,N_8661,N_9035);
nand U10301 (N_10301,N_8204,N_9382);
nand U10302 (N_10302,N_8200,N_9335);
nor U10303 (N_10303,N_8983,N_8266);
nand U10304 (N_10304,N_8136,N_9200);
and U10305 (N_10305,N_8897,N_8831);
or U10306 (N_10306,N_9937,N_9201);
xor U10307 (N_10307,N_9449,N_8596);
and U10308 (N_10308,N_8574,N_8589);
or U10309 (N_10309,N_9412,N_9589);
and U10310 (N_10310,N_8250,N_9089);
xor U10311 (N_10311,N_8161,N_8535);
nor U10312 (N_10312,N_8480,N_9006);
or U10313 (N_10313,N_8418,N_8004);
xor U10314 (N_10314,N_8779,N_8958);
nor U10315 (N_10315,N_8685,N_8047);
or U10316 (N_10316,N_8850,N_8165);
nor U10317 (N_10317,N_8947,N_8595);
xnor U10318 (N_10318,N_8909,N_8887);
and U10319 (N_10319,N_9374,N_8318);
and U10320 (N_10320,N_8796,N_8584);
or U10321 (N_10321,N_8263,N_9968);
and U10322 (N_10322,N_9118,N_9191);
xnor U10323 (N_10323,N_9403,N_8323);
nor U10324 (N_10324,N_9621,N_8237);
and U10325 (N_10325,N_8634,N_9136);
or U10326 (N_10326,N_8828,N_8592);
xor U10327 (N_10327,N_9063,N_8096);
and U10328 (N_10328,N_8579,N_9542);
and U10329 (N_10329,N_8469,N_9735);
nand U10330 (N_10330,N_9878,N_9377);
nor U10331 (N_10331,N_9172,N_8541);
nor U10332 (N_10332,N_9508,N_8286);
xor U10333 (N_10333,N_9556,N_9431);
or U10334 (N_10334,N_9233,N_8872);
nor U10335 (N_10335,N_8114,N_9164);
or U10336 (N_10336,N_9557,N_9432);
or U10337 (N_10337,N_8550,N_8182);
nor U10338 (N_10338,N_9767,N_9422);
and U10339 (N_10339,N_9956,N_8666);
xnor U10340 (N_10340,N_9692,N_9661);
or U10341 (N_10341,N_9243,N_9697);
xnor U10342 (N_10342,N_8884,N_9686);
or U10343 (N_10343,N_8061,N_8291);
nand U10344 (N_10344,N_9390,N_8646);
and U10345 (N_10345,N_8994,N_8763);
xnor U10346 (N_10346,N_9611,N_8674);
nand U10347 (N_10347,N_8424,N_9986);
or U10348 (N_10348,N_8134,N_9787);
nand U10349 (N_10349,N_9473,N_8057);
nand U10350 (N_10350,N_8275,N_8755);
or U10351 (N_10351,N_9570,N_8648);
nand U10352 (N_10352,N_8176,N_9165);
and U10353 (N_10353,N_9187,N_9420);
nor U10354 (N_10354,N_8921,N_9871);
or U10355 (N_10355,N_8799,N_8542);
or U10356 (N_10356,N_8900,N_9464);
and U10357 (N_10357,N_9916,N_8874);
nor U10358 (N_10358,N_9987,N_9958);
and U10359 (N_10359,N_9421,N_9530);
nand U10360 (N_10360,N_8538,N_8764);
xor U10361 (N_10361,N_9166,N_9824);
or U10362 (N_10362,N_8507,N_9029);
nor U10363 (N_10363,N_9826,N_9951);
nor U10364 (N_10364,N_9102,N_8903);
nand U10365 (N_10365,N_8875,N_9180);
and U10366 (N_10366,N_9877,N_8435);
xor U10367 (N_10367,N_9447,N_8221);
nand U10368 (N_10368,N_9924,N_8454);
or U10369 (N_10369,N_8331,N_9690);
nor U10370 (N_10370,N_9751,N_9717);
and U10371 (N_10371,N_8976,N_9394);
nor U10372 (N_10372,N_9226,N_9151);
nand U10373 (N_10373,N_8032,N_8252);
nand U10374 (N_10374,N_8543,N_9489);
or U10375 (N_10375,N_8533,N_8684);
nor U10376 (N_10376,N_8954,N_8810);
nor U10377 (N_10377,N_9744,N_8898);
and U10378 (N_10378,N_9231,N_9111);
or U10379 (N_10379,N_8464,N_9852);
or U10380 (N_10380,N_9244,N_9186);
nand U10381 (N_10381,N_8825,N_8668);
xor U10382 (N_10382,N_9114,N_9189);
nor U10383 (N_10383,N_8267,N_8680);
xor U10384 (N_10384,N_9124,N_9520);
or U10385 (N_10385,N_8908,N_9982);
and U10386 (N_10386,N_8913,N_9129);
nor U10387 (N_10387,N_9478,N_9229);
nand U10388 (N_10388,N_9953,N_9090);
nor U10389 (N_10389,N_8740,N_8442);
nor U10390 (N_10390,N_8815,N_9094);
and U10391 (N_10391,N_9054,N_8794);
xor U10392 (N_10392,N_9159,N_9339);
nor U10393 (N_10393,N_8137,N_8832);
nand U10394 (N_10394,N_8206,N_9171);
xnor U10395 (N_10395,N_9108,N_9899);
nor U10396 (N_10396,N_8588,N_9263);
xnor U10397 (N_10397,N_9629,N_8475);
nand U10398 (N_10398,N_8294,N_8558);
xnor U10399 (N_10399,N_9120,N_8083);
nor U10400 (N_10400,N_9485,N_9875);
nand U10401 (N_10401,N_8849,N_8985);
nor U10402 (N_10402,N_8515,N_8486);
nor U10403 (N_10403,N_9030,N_8452);
xor U10404 (N_10404,N_9070,N_8800);
nand U10405 (N_10405,N_8466,N_9173);
xor U10406 (N_10406,N_9342,N_8502);
nand U10407 (N_10407,N_8622,N_9290);
nor U10408 (N_10408,N_8998,N_8149);
nor U10409 (N_10409,N_8822,N_9606);
xor U10410 (N_10410,N_9268,N_9588);
and U10411 (N_10411,N_8020,N_8745);
and U10412 (N_10412,N_9396,N_8926);
or U10413 (N_10413,N_9739,N_9253);
xor U10414 (N_10414,N_8536,N_8396);
or U10415 (N_10415,N_8487,N_9052);
and U10416 (N_10416,N_9722,N_9965);
nand U10417 (N_10417,N_8888,N_8729);
and U10418 (N_10418,N_9768,N_8238);
and U10419 (N_10419,N_9409,N_9415);
xnor U10420 (N_10420,N_9984,N_8846);
xnor U10421 (N_10421,N_9153,N_8369);
and U10422 (N_10422,N_8269,N_8090);
xor U10423 (N_10423,N_9259,N_9844);
or U10424 (N_10424,N_8462,N_8290);
or U10425 (N_10425,N_9738,N_8231);
xnor U10426 (N_10426,N_8567,N_8863);
xor U10427 (N_10427,N_8392,N_8655);
xor U10428 (N_10428,N_8692,N_8491);
or U10429 (N_10429,N_8880,N_9544);
or U10430 (N_10430,N_8105,N_9962);
and U10431 (N_10431,N_8362,N_9856);
xor U10432 (N_10432,N_8889,N_9506);
and U10433 (N_10433,N_8359,N_8682);
or U10434 (N_10434,N_8858,N_8662);
and U10435 (N_10435,N_9440,N_8805);
or U10436 (N_10436,N_9305,N_9325);
nor U10437 (N_10437,N_8235,N_9590);
nand U10438 (N_10438,N_8122,N_8955);
nor U10439 (N_10439,N_8973,N_9110);
nor U10440 (N_10440,N_8239,N_9088);
xor U10441 (N_10441,N_9591,N_9062);
nor U10442 (N_10442,N_8722,N_9853);
nand U10443 (N_10443,N_9130,N_8219);
and U10444 (N_10444,N_8753,N_9273);
or U10445 (N_10445,N_8316,N_8285);
nor U10446 (N_10446,N_9562,N_9075);
nand U10447 (N_10447,N_8222,N_8599);
nor U10448 (N_10448,N_8270,N_9811);
nand U10449 (N_10449,N_9823,N_8188);
nand U10450 (N_10450,N_8586,N_9938);
nand U10451 (N_10451,N_8594,N_8728);
and U10452 (N_10452,N_9617,N_8321);
and U10453 (N_10453,N_9149,N_9084);
nand U10454 (N_10454,N_8547,N_9001);
and U10455 (N_10455,N_8700,N_8126);
and U10456 (N_10456,N_8824,N_9537);
nand U10457 (N_10457,N_8258,N_8514);
nor U10458 (N_10458,N_8645,N_9104);
xor U10459 (N_10459,N_9210,N_9154);
nand U10460 (N_10460,N_9178,N_8793);
nor U10461 (N_10461,N_8340,N_9992);
nor U10462 (N_10462,N_9700,N_8509);
nand U10463 (N_10463,N_8708,N_9943);
nor U10464 (N_10464,N_8590,N_8385);
and U10465 (N_10465,N_9820,N_8179);
xnor U10466 (N_10466,N_9645,N_9341);
or U10467 (N_10467,N_9362,N_8797);
nor U10468 (N_10468,N_8970,N_9516);
nor U10469 (N_10469,N_8313,N_9974);
nand U10470 (N_10470,N_8141,N_9654);
or U10471 (N_10471,N_8051,N_8653);
nand U10472 (N_10472,N_9602,N_9814);
or U10473 (N_10473,N_8786,N_9254);
xnor U10474 (N_10474,N_9039,N_9023);
xor U10475 (N_10475,N_8242,N_8665);
nand U10476 (N_10476,N_9766,N_9388);
nand U10477 (N_10477,N_8933,N_9928);
nor U10478 (N_10478,N_8413,N_9067);
nand U10479 (N_10479,N_9545,N_8068);
nor U10480 (N_10480,N_8317,N_8996);
or U10481 (N_10481,N_8964,N_8899);
and U10482 (N_10482,N_8246,N_8065);
nor U10483 (N_10483,N_8761,N_8416);
or U10484 (N_10484,N_9846,N_8762);
xnor U10485 (N_10485,N_8848,N_9801);
or U10486 (N_10486,N_8798,N_8882);
or U10487 (N_10487,N_9284,N_8227);
and U10488 (N_10488,N_8891,N_8208);
or U10489 (N_10489,N_8614,N_9317);
xor U10490 (N_10490,N_8274,N_8860);
and U10491 (N_10491,N_9298,N_8278);
xnor U10492 (N_10492,N_8843,N_9582);
and U10493 (N_10493,N_8551,N_8950);
or U10494 (N_10494,N_8620,N_8642);
nand U10495 (N_10495,N_8488,N_9100);
nor U10496 (N_10496,N_8990,N_9428);
and U10497 (N_10497,N_9773,N_9140);
and U10498 (N_10498,N_9291,N_8935);
and U10499 (N_10499,N_9927,N_9989);
nand U10500 (N_10500,N_9218,N_8333);
or U10501 (N_10501,N_8324,N_8896);
nor U10502 (N_10502,N_9105,N_9763);
nor U10503 (N_10503,N_8792,N_8760);
and U10504 (N_10504,N_9595,N_8808);
nand U10505 (N_10505,N_8737,N_8429);
and U10506 (N_10506,N_9800,N_9861);
nor U10507 (N_10507,N_9137,N_9527);
and U10508 (N_10508,N_9143,N_9385);
xnor U10509 (N_10509,N_8552,N_9345);
nor U10510 (N_10510,N_9208,N_9184);
and U10511 (N_10511,N_8082,N_8785);
nor U10512 (N_10512,N_8071,N_8767);
nand U10513 (N_10513,N_8198,N_9160);
and U10514 (N_10514,N_8110,N_8381);
nor U10515 (N_10515,N_8490,N_8053);
and U10516 (N_10516,N_8041,N_9402);
or U10517 (N_10517,N_9177,N_9293);
nand U10518 (N_10518,N_9275,N_9599);
xnor U10519 (N_10519,N_9194,N_9397);
nand U10520 (N_10520,N_8018,N_8774);
and U10521 (N_10521,N_8100,N_9715);
nor U10522 (N_10522,N_8501,N_9893);
xor U10523 (N_10523,N_8417,N_8076);
xor U10524 (N_10524,N_9905,N_9957);
nor U10525 (N_10525,N_9559,N_8223);
and U10526 (N_10526,N_8878,N_8393);
xor U10527 (N_10527,N_9442,N_9580);
nor U10528 (N_10528,N_8070,N_8271);
xor U10529 (N_10529,N_8151,N_8924);
xor U10530 (N_10530,N_8450,N_9190);
and U10531 (N_10531,N_8873,N_9224);
xor U10532 (N_10532,N_8868,N_9262);
or U10533 (N_10533,N_8431,N_8108);
nand U10534 (N_10534,N_8058,N_9433);
and U10535 (N_10535,N_8163,N_9538);
nand U10536 (N_10536,N_9349,N_8158);
and U10537 (N_10537,N_8207,N_8549);
nand U10538 (N_10538,N_9156,N_8999);
nand U10539 (N_10539,N_8566,N_9360);
nand U10540 (N_10540,N_9344,N_8279);
nor U10541 (N_10541,N_8641,N_9518);
xnor U10542 (N_10542,N_9363,N_9607);
nand U10543 (N_10543,N_9529,N_9400);
nor U10544 (N_10544,N_8420,N_9815);
nand U10545 (N_10545,N_8939,N_8023);
nand U10546 (N_10546,N_8159,N_9324);
nor U10547 (N_10547,N_8748,N_9043);
nand U10548 (N_10548,N_9020,N_8859);
or U10549 (N_10549,N_8074,N_9865);
or U10550 (N_10550,N_9359,N_8017);
and U10551 (N_10551,N_9837,N_8107);
and U10552 (N_10552,N_9487,N_8470);
or U10553 (N_10553,N_8965,N_9584);
xnor U10554 (N_10554,N_8492,N_9797);
or U10555 (N_10555,N_8218,N_9998);
nand U10556 (N_10556,N_8777,N_8853);
nand U10557 (N_10557,N_9435,N_8768);
xnor U10558 (N_10558,N_8099,N_9999);
nand U10559 (N_10559,N_8402,N_9727);
nor U10560 (N_10560,N_8602,N_9490);
or U10561 (N_10561,N_9502,N_9141);
xnor U10562 (N_10562,N_9695,N_8309);
nand U10563 (N_10563,N_9098,N_9198);
or U10564 (N_10564,N_8372,N_9381);
nand U10565 (N_10565,N_8690,N_8510);
nor U10566 (N_10566,N_9714,N_9868);
and U10567 (N_10567,N_8423,N_8019);
nand U10568 (N_10568,N_8691,N_9648);
xnor U10569 (N_10569,N_9828,N_9407);
xnor U10570 (N_10570,N_8395,N_9525);
or U10571 (N_10571,N_8325,N_9678);
nand U10572 (N_10572,N_9051,N_9933);
nand U10573 (N_10573,N_9055,N_9115);
nand U10574 (N_10574,N_8942,N_8917);
xor U10575 (N_10575,N_9630,N_9479);
nor U10576 (N_10576,N_8681,N_9628);
and U10577 (N_10577,N_8563,N_8637);
or U10578 (N_10578,N_8170,N_8654);
xnor U10579 (N_10579,N_8129,N_9762);
xor U10580 (N_10580,N_8953,N_8093);
nor U10581 (N_10581,N_9886,N_9585);
nand U10582 (N_10582,N_9960,N_8443);
nor U10583 (N_10583,N_8138,N_8012);
and U10584 (N_10584,N_8072,N_8957);
nor U10585 (N_10585,N_8598,N_8453);
or U10586 (N_10586,N_9790,N_9625);
xnor U10587 (N_10587,N_8460,N_8840);
nand U10588 (N_10588,N_8639,N_9759);
nand U10589 (N_10589,N_9134,N_8980);
or U10590 (N_10590,N_9605,N_8199);
nor U10591 (N_10591,N_8297,N_9966);
nand U10592 (N_10592,N_8575,N_9047);
or U10593 (N_10593,N_9256,N_9995);
or U10594 (N_10594,N_9950,N_8013);
or U10595 (N_10595,N_8039,N_9698);
xnor U10596 (N_10596,N_9379,N_9214);
nand U10597 (N_10597,N_9650,N_9007);
xor U10598 (N_10598,N_8300,N_8033);
nor U10599 (N_10599,N_9250,N_8066);
nor U10600 (N_10600,N_8989,N_8930);
or U10601 (N_10601,N_9337,N_8356);
and U10602 (N_10602,N_8895,N_8696);
nor U10603 (N_10603,N_9368,N_8750);
xnor U10604 (N_10604,N_8240,N_9873);
nand U10605 (N_10605,N_9249,N_9373);
nand U10606 (N_10606,N_9675,N_8292);
and U10607 (N_10607,N_8201,N_9087);
or U10608 (N_10608,N_9798,N_8659);
nor U10609 (N_10609,N_8439,N_8531);
nand U10610 (N_10610,N_8508,N_8697);
nor U10611 (N_10611,N_9948,N_8203);
or U10612 (N_10612,N_8277,N_9548);
nor U10613 (N_10613,N_8744,N_9652);
xnor U10614 (N_10614,N_9281,N_9737);
and U10615 (N_10615,N_8739,N_8789);
and U10616 (N_10616,N_9294,N_9125);
and U10617 (N_10617,N_9213,N_9632);
or U10618 (N_10618,N_8458,N_8865);
and U10619 (N_10619,N_8168,N_9401);
or U10620 (N_10620,N_8869,N_8670);
and U10621 (N_10621,N_9579,N_8189);
and U10622 (N_10622,N_9215,N_9326);
xnor U10623 (N_10623,N_9804,N_8410);
nand U10624 (N_10624,N_9091,N_9624);
and U10625 (N_10625,N_8521,N_8608);
or U10626 (N_10626,N_8236,N_9492);
and U10627 (N_10627,N_9031,N_8293);
nand U10628 (N_10628,N_9769,N_8705);
nand U10629 (N_10629,N_9573,N_9338);
nand U10630 (N_10630,N_8174,N_9919);
and U10631 (N_10631,N_9850,N_9465);
xnor U10632 (N_10632,N_9794,N_9497);
xor U10633 (N_10633,N_8383,N_8624);
and U10634 (N_10634,N_8374,N_8630);
xor U10635 (N_10635,N_9451,N_9004);
nand U10636 (N_10636,N_8112,N_9897);
and U10637 (N_10637,N_9519,N_8519);
nor U10638 (N_10638,N_9076,N_8190);
nor U10639 (N_10639,N_9671,N_8155);
xnor U10640 (N_10640,N_8186,N_9915);
xnor U10641 (N_10641,N_9532,N_9901);
nor U10642 (N_10642,N_9819,N_8440);
xnor U10643 (N_10643,N_9949,N_9083);
xnor U10644 (N_10644,N_9760,N_9267);
and U10645 (N_10645,N_9702,N_9576);
xnor U10646 (N_10646,N_8262,N_8143);
nor U10647 (N_10647,N_8816,N_8095);
and U10648 (N_10648,N_8081,N_8433);
xor U10649 (N_10649,N_8765,N_9818);
nand U10650 (N_10650,N_8343,N_8348);
xor U10651 (N_10651,N_9750,N_8363);
nand U10652 (N_10652,N_8776,N_8447);
xor U10653 (N_10653,N_8787,N_8802);
xnor U10654 (N_10654,N_8505,N_9106);
or U10655 (N_10655,N_9469,N_9827);
and U10656 (N_10656,N_8714,N_9016);
and U10657 (N_10657,N_9587,N_9963);
nand U10658 (N_10658,N_9477,N_8713);
nor U10659 (N_10659,N_9898,N_8627);
nor U10660 (N_10660,N_9920,N_9217);
xor U10661 (N_10661,N_8280,N_9914);
or U10662 (N_10662,N_8268,N_9955);
nor U10663 (N_10663,N_8709,N_8960);
nand U10664 (N_10664,N_9086,N_8851);
nor U10665 (N_10665,N_8529,N_8725);
and U10666 (N_10666,N_8306,N_8428);
nor U10667 (N_10667,N_8397,N_8498);
nor U10668 (N_10668,N_9230,N_9892);
and U10669 (N_10669,N_9682,N_8247);
or U10670 (N_10670,N_9895,N_9543);
and U10671 (N_10671,N_9439,N_9954);
xnor U10672 (N_10672,N_9255,N_8638);
and U10673 (N_10673,N_8459,N_8525);
nand U10674 (N_10674,N_8482,N_8672);
xor U10675 (N_10675,N_8069,N_8694);
nand U10676 (N_10676,N_8870,N_8995);
nand U10677 (N_10677,N_8405,N_8747);
and U10678 (N_10678,N_9417,N_9211);
nor U10679 (N_10679,N_8966,N_8625);
and U10680 (N_10680,N_9225,N_8636);
nand U10681 (N_10681,N_9181,N_8255);
xnor U10682 (N_10682,N_8075,N_8109);
nand U10683 (N_10683,N_9803,N_8437);
or U10684 (N_10684,N_9926,N_9592);
nor U10685 (N_10685,N_8409,N_9283);
nor U10686 (N_10686,N_8040,N_8379);
and U10687 (N_10687,N_8972,N_9521);
or U10688 (N_10688,N_9299,N_9248);
or U10689 (N_10689,N_9908,N_9859);
xnor U10690 (N_10690,N_8650,N_9288);
xnor U10691 (N_10691,N_8024,N_8028);
xnor U10692 (N_10692,N_8742,N_9631);
nor U10693 (N_10693,N_9179,N_9706);
or U10694 (N_10694,N_8230,N_9838);
nand U10695 (N_10695,N_8283,N_9480);
or U10696 (N_10696,N_9174,N_9482);
nand U10697 (N_10697,N_8427,N_9792);
nor U10698 (N_10698,N_9242,N_8307);
xnor U10699 (N_10699,N_8679,N_8228);
xor U10700 (N_10700,N_8778,N_9566);
and U10701 (N_10701,N_8936,N_8754);
nand U10702 (N_10702,N_9743,N_9365);
xnor U10703 (N_10703,N_9723,N_9869);
nand U10704 (N_10704,N_8389,N_9109);
or U10705 (N_10705,N_9022,N_9749);
or U10706 (N_10706,N_9308,N_9307);
or U10707 (N_10707,N_8191,N_9257);
and U10708 (N_10708,N_9264,N_8803);
and U10709 (N_10709,N_9251,N_8731);
or U10710 (N_10710,N_9456,N_9679);
nor U10711 (N_10711,N_9860,N_9014);
xnor U10712 (N_10712,N_8967,N_8007);
and U10713 (N_10713,N_8091,N_8829);
xor U10714 (N_10714,N_9366,N_8894);
nand U10715 (N_10715,N_8187,N_8856);
nand U10716 (N_10716,N_9448,N_9475);
or U10717 (N_10717,N_8591,N_9975);
xnor U10718 (N_10718,N_9889,N_9646);
nand U10719 (N_10719,N_9033,N_9598);
and U10720 (N_10720,N_8814,N_9567);
and U10721 (N_10721,N_8386,N_9236);
nand U10722 (N_10722,N_8421,N_9786);
nand U10723 (N_10723,N_9687,N_8049);
nor U10724 (N_10724,N_9734,N_8726);
nand U10725 (N_10725,N_9474,N_9340);
nand U10726 (N_10726,N_8734,N_9540);
xnor U10727 (N_10727,N_8975,N_9791);
xor U10728 (N_10728,N_9025,N_8493);
or U10729 (N_10729,N_8997,N_8388);
or U10730 (N_10730,N_8581,N_9701);
or U10731 (N_10731,N_8526,N_8751);
or U10732 (N_10732,N_9614,N_8354);
or U10733 (N_10733,N_8319,N_8813);
or U10734 (N_10734,N_8123,N_9199);
or U10735 (N_10735,N_9386,N_8842);
nor U10736 (N_10736,N_9292,N_9903);
nor U10737 (N_10737,N_8927,N_9934);
nor U10738 (N_10738,N_8733,N_8302);
nand U10739 (N_10739,N_8312,N_9351);
and U10740 (N_10740,N_8154,N_9158);
or U10741 (N_10741,N_9673,N_8532);
or U10742 (N_10742,N_9522,N_8063);
nand U10743 (N_10743,N_8403,N_9728);
nor U10744 (N_10744,N_9332,N_9644);
nand U10745 (N_10745,N_9375,N_9392);
xor U10746 (N_10746,N_8735,N_9674);
nor U10747 (N_10747,N_8827,N_8780);
or U10748 (N_10748,N_8573,N_8664);
and U10749 (N_10749,N_9355,N_8877);
nand U10750 (N_10750,N_9196,N_8479);
and U10751 (N_10751,N_8530,N_8658);
and U10752 (N_10752,N_8035,N_8612);
or U10753 (N_10753,N_9896,N_8101);
and U10754 (N_10754,N_8144,N_9096);
xnor U10755 (N_10755,N_8473,N_8337);
nand U10756 (N_10756,N_9681,N_9812);
and U10757 (N_10757,N_9048,N_8962);
and U10758 (N_10758,N_9276,N_8830);
and U10759 (N_10759,N_8037,N_8401);
or U10760 (N_10760,N_8984,N_8288);
nand U10761 (N_10761,N_8097,N_9774);
or U10762 (N_10762,N_8580,N_8406);
or U10763 (N_10763,N_8890,N_9636);
nand U10764 (N_10764,N_8465,N_8928);
or U10765 (N_10765,N_9597,N_8036);
nand U10766 (N_10766,N_8835,N_8113);
and U10767 (N_10767,N_8556,N_8139);
and U10768 (N_10768,N_8329,N_9504);
or U10769 (N_10769,N_8651,N_9427);
xnor U10770 (N_10770,N_8295,N_9634);
and U10771 (N_10771,N_9058,N_9755);
and U10772 (N_10772,N_9505,N_9069);
xor U10773 (N_10773,N_8993,N_8477);
and U10774 (N_10774,N_9404,N_9081);
xor U10775 (N_10775,N_9782,N_8346);
nor U10776 (N_10776,N_8249,N_8766);
or U10777 (N_10777,N_8883,N_9848);
and U10778 (N_10778,N_9876,N_8545);
nand U10779 (N_10779,N_9581,N_9959);
xor U10780 (N_10780,N_9913,N_8601);
nand U10781 (N_10781,N_8398,N_8366);
or U10782 (N_10782,N_9195,N_8353);
and U10783 (N_10783,N_9721,N_8683);
nand U10784 (N_10784,N_8147,N_8092);
nand U10785 (N_10785,N_8497,N_9222);
or U10786 (N_10786,N_8513,N_8478);
nor U10787 (N_10787,N_8078,N_8518);
xor U10788 (N_10788,N_8539,N_8414);
xnor U10789 (N_10789,N_8660,N_9425);
xnor U10790 (N_10790,N_9560,N_8938);
and U10791 (N_10791,N_9796,N_9045);
or U10792 (N_10792,N_9501,N_8818);
nand U10793 (N_10793,N_9356,N_9825);
and U10794 (N_10794,N_9836,N_8626);
xnor U10795 (N_10795,N_8607,N_8656);
or U10796 (N_10796,N_8845,N_8021);
nor U10797 (N_10797,N_9176,N_9608);
nor U10798 (N_10798,N_9810,N_9265);
xnor U10799 (N_10799,N_9741,N_9864);
or U10800 (N_10800,N_9423,N_9128);
nand U10801 (N_10801,N_8365,N_9946);
xnor U10802 (N_10802,N_8234,N_8961);
and U10803 (N_10803,N_9816,N_8948);
and U10804 (N_10804,N_9565,N_9117);
nand U10805 (N_10805,N_9718,N_9547);
nand U10806 (N_10806,N_8560,N_8145);
xnor U10807 (N_10807,N_9894,N_9486);
xnor U10808 (N_10808,N_8089,N_8178);
nand U10809 (N_10809,N_8373,N_9610);
xnor U10810 (N_10810,N_8010,N_9561);
or U10811 (N_10811,N_8054,N_9952);
nand U10812 (N_10812,N_8743,N_9930);
nand U10813 (N_10813,N_8949,N_9568);
or U10814 (N_10814,N_8347,N_9649);
nand U10815 (N_10815,N_8253,N_9452);
xor U10816 (N_10816,N_9367,N_8146);
nand U10817 (N_10817,N_8160,N_8657);
and U10818 (N_10818,N_9170,N_9944);
and U10819 (N_10819,N_8016,N_9694);
xnor U10820 (N_10820,N_9221,N_9416);
nor U10821 (N_10821,N_9135,N_9238);
nand U10822 (N_10822,N_9627,N_9346);
xnor U10823 (N_10823,N_9000,N_9316);
xnor U10824 (N_10824,N_9053,N_9364);
or U10825 (N_10825,N_9667,N_8202);
nor U10826 (N_10826,N_9239,N_8844);
or U10827 (N_10827,N_8982,N_8457);
and U10828 (N_10828,N_8652,N_8349);
or U10829 (N_10829,N_9857,N_8540);
and U10830 (N_10830,N_8328,N_9639);
and U10831 (N_10831,N_8339,N_8217);
xnor U10832 (N_10832,N_8120,N_9057);
nand U10833 (N_10833,N_9523,N_9393);
xor U10834 (N_10834,N_9376,N_9922);
nor U10835 (N_10835,N_8712,N_8775);
nand U10836 (N_10836,N_8384,N_9809);
and U10837 (N_10837,N_9670,N_9524);
and U10838 (N_10838,N_9227,N_9202);
or U10839 (N_10839,N_8686,N_8593);
and U10840 (N_10840,N_8687,N_9669);
xor U10841 (N_10841,N_9783,N_9510);
nand U10842 (N_10842,N_9252,N_8311);
or U10843 (N_10843,N_9037,N_8644);
xnor U10844 (N_10844,N_8243,N_9336);
and U10845 (N_10845,N_9119,N_9747);
xnor U10846 (N_10846,N_8355,N_8841);
or U10847 (N_10847,N_9620,N_9395);
and U10848 (N_10848,N_9533,N_9536);
nand U10849 (N_10849,N_8944,N_8643);
nand U10850 (N_10850,N_9398,N_9212);
nor U10851 (N_10851,N_8922,N_9245);
xnor U10852 (N_10852,N_8979,N_9468);
and U10853 (N_10853,N_8485,N_9462);
nand U10854 (N_10854,N_8617,N_9784);
nor U10855 (N_10855,N_9353,N_9945);
nand U10856 (N_10856,N_9724,N_9985);
nand U10857 (N_10857,N_9314,N_8929);
nor U10858 (N_10858,N_9460,N_9099);
nor U10859 (N_10859,N_9961,N_8358);
or U10860 (N_10860,N_9018,N_9541);
xnor U10861 (N_10861,N_9327,N_9470);
and U10862 (N_10862,N_9615,N_8244);
nand U10863 (N_10863,N_9531,N_8857);
and U10864 (N_10864,N_9770,N_9138);
nand U10865 (N_10865,N_9641,N_9445);
nor U10866 (N_10866,N_9457,N_9666);
nand U10867 (N_10867,N_8115,N_9361);
xnor U10868 (N_10868,N_8476,N_9240);
nand U10869 (N_10869,N_9319,N_8854);
nand U10870 (N_10870,N_8806,N_9534);
and U10871 (N_10871,N_8419,N_9418);
nor U10872 (N_10872,N_9296,N_8391);
and U10873 (N_10873,N_9752,N_9583);
nor U10874 (N_10874,N_8467,N_8260);
nor U10875 (N_10875,N_9437,N_8838);
nor U10876 (N_10876,N_9967,N_9660);
and U10877 (N_10877,N_8977,N_8209);
nor U10878 (N_10878,N_8752,N_8867);
and U10879 (N_10879,N_9858,N_9123);
or U10880 (N_10880,N_8738,N_9101);
nor U10881 (N_10881,N_8583,N_9699);
and U10882 (N_10882,N_8282,N_9849);
xnor U10883 (N_10883,N_8298,N_8912);
or U10884 (N_10884,N_8616,N_9493);
and U10885 (N_10885,N_9994,N_9971);
or U10886 (N_10886,N_9498,N_9854);
or U10887 (N_10887,N_8522,N_9637);
xnor U10888 (N_10888,N_8434,N_8688);
xor U10889 (N_10889,N_8807,N_8758);
nand U10890 (N_10890,N_8079,N_8703);
or U10891 (N_10891,N_9929,N_9729);
xnor U10892 (N_10892,N_9574,N_8471);
xor U10893 (N_10893,N_9078,N_9709);
and U10894 (N_10894,N_8881,N_9710);
nor U10895 (N_10895,N_8210,N_9676);
or U10896 (N_10896,N_8248,N_8864);
nor U10897 (N_10897,N_9183,N_8554);
nand U10898 (N_10898,N_8142,N_8034);
nor U10899 (N_10899,N_8059,N_9049);
or U10900 (N_10900,N_8925,N_9074);
xnor U10901 (N_10901,N_9640,N_9348);
nand U10902 (N_10902,N_8106,N_8677);
and U10903 (N_10903,N_8920,N_9066);
nor U10904 (N_10904,N_9011,N_9917);
nor U10905 (N_10905,N_9558,N_9713);
and U10906 (N_10906,N_9842,N_8338);
nor U10907 (N_10907,N_9371,N_8132);
nand U10908 (N_10908,N_8548,N_9399);
nand U10909 (N_10909,N_8430,N_9601);
nor U10910 (N_10910,N_9419,N_8284);
and U10911 (N_10911,N_8387,N_8166);
nand U10912 (N_10912,N_9993,N_8130);
xor U10913 (N_10913,N_9380,N_8968);
xor U10914 (N_10914,N_9834,N_9261);
nor U10915 (N_10915,N_8974,N_8014);
and U10916 (N_10916,N_9925,N_9941);
and U10917 (N_10917,N_8951,N_9586);
nor U10918 (N_10918,N_8923,N_9616);
or U10919 (N_10919,N_8345,N_9940);
or U10920 (N_10920,N_8910,N_9983);
nor U10921 (N_10921,N_8905,N_9444);
nand U10922 (N_10922,N_9357,N_8698);
xnor U10923 (N_10923,N_8495,N_9085);
and U10924 (N_10924,N_9665,N_9414);
and U10925 (N_10925,N_8257,N_8496);
or U10926 (N_10926,N_8959,N_9932);
nor U10927 (N_10927,N_8500,N_8578);
nor U10928 (N_10928,N_8212,N_9658);
xor U10929 (N_10929,N_9038,N_9555);
xnor U10930 (N_10930,N_9237,N_8102);
xor U10931 (N_10931,N_9907,N_9612);
nor U10932 (N_10932,N_8504,N_9754);
and U10933 (N_10933,N_9781,N_9890);
xnor U10934 (N_10934,N_8576,N_8876);
nand U10935 (N_10935,N_8455,N_8699);
xnor U10936 (N_10936,N_9306,N_9503);
nor U10937 (N_10937,N_9526,N_9438);
nand U10938 (N_10938,N_9638,N_9436);
or U10939 (N_10939,N_8103,N_8438);
nand U10940 (N_10940,N_8811,N_9888);
xnor U10941 (N_10941,N_9481,N_9044);
nor U10942 (N_10942,N_8344,N_9147);
xor U10943 (N_10943,N_9840,N_8335);
nor U10944 (N_10944,N_8415,N_8121);
and U10945 (N_10945,N_9046,N_8357);
xor U10946 (N_10946,N_8945,N_9310);
nor U10947 (N_10947,N_8445,N_8562);
nand U10948 (N_10948,N_8377,N_8474);
nand U10949 (N_10949,N_9703,N_8407);
nor U10950 (N_10950,N_8162,N_9144);
nand U10951 (N_10951,N_8000,N_9193);
or U10952 (N_10952,N_9978,N_9788);
nor U10953 (N_10953,N_9829,N_9923);
nand U10954 (N_10954,N_8916,N_8448);
and U10955 (N_10955,N_9939,N_9712);
or U10956 (N_10956,N_9278,N_8245);
and U10957 (N_10957,N_8472,N_9167);
nor U10958 (N_10958,N_9942,N_8676);
nand U10959 (N_10959,N_9981,N_9024);
nand U10960 (N_10960,N_9343,N_8565);
or U10961 (N_10961,N_9688,N_9732);
nor U10962 (N_10962,N_9604,N_8150);
nor U10963 (N_10963,N_9577,N_8088);
nor U10964 (N_10964,N_9609,N_9378);
or U10965 (N_10965,N_9659,N_8885);
or U10966 (N_10966,N_9021,N_9065);
nor U10967 (N_10967,N_8456,N_9891);
and U10968 (N_10968,N_8978,N_8444);
and U10969 (N_10969,N_8569,N_9494);
nor U10970 (N_10970,N_9133,N_9870);
nand U10971 (N_10971,N_9707,N_9805);
xor U10972 (N_10972,N_9272,N_8370);
or U10973 (N_10973,N_9879,N_9495);
nor U10974 (N_10974,N_9756,N_8619);
or U10975 (N_10975,N_9121,N_9551);
xor U10976 (N_10976,N_9691,N_9112);
nor U10977 (N_10977,N_9885,N_9906);
nor U10978 (N_10978,N_8449,N_9384);
xor U10979 (N_10979,N_8371,N_8352);
and U10980 (N_10980,N_9866,N_9647);
xor U10981 (N_10981,N_8229,N_8812);
or U10982 (N_10982,N_9483,N_8570);
and U10983 (N_10983,N_8045,N_8736);
or U10984 (N_10984,N_9672,N_8771);
or U10985 (N_10985,N_9463,N_9863);
or U10986 (N_10986,N_9163,N_8367);
xnor U10987 (N_10987,N_9593,N_9369);
or U10988 (N_10988,N_9514,N_9329);
nand U10989 (N_10989,N_8937,N_8633);
and U10990 (N_10990,N_8180,N_8233);
xnor U10991 (N_10991,N_8214,N_8833);
and U10992 (N_10992,N_8783,N_9139);
nor U10993 (N_10993,N_8635,N_9693);
nor U10994 (N_10994,N_9168,N_9758);
xnor U10995 (N_10995,N_8148,N_8192);
nand U10996 (N_10996,N_9207,N_8408);
and U10997 (N_10997,N_9684,N_9552);
or U10998 (N_10998,N_9564,N_8553);
nor U10999 (N_10999,N_8351,N_8128);
nor U11000 (N_11000,N_9715,N_9363);
nand U11001 (N_11001,N_8556,N_8553);
nor U11002 (N_11002,N_8694,N_9982);
nor U11003 (N_11003,N_9432,N_9574);
nand U11004 (N_11004,N_8270,N_8912);
nand U11005 (N_11005,N_8947,N_9911);
and U11006 (N_11006,N_8654,N_9477);
or U11007 (N_11007,N_8233,N_9225);
xor U11008 (N_11008,N_9506,N_9216);
nor U11009 (N_11009,N_8355,N_8566);
xor U11010 (N_11010,N_8171,N_9716);
nor U11011 (N_11011,N_9935,N_9937);
xor U11012 (N_11012,N_9895,N_9771);
or U11013 (N_11013,N_9716,N_9471);
and U11014 (N_11014,N_8061,N_8027);
xor U11015 (N_11015,N_8755,N_9935);
nor U11016 (N_11016,N_9990,N_8935);
nand U11017 (N_11017,N_9451,N_9159);
nor U11018 (N_11018,N_9353,N_8919);
nand U11019 (N_11019,N_8555,N_8420);
xnor U11020 (N_11020,N_9237,N_8182);
and U11021 (N_11021,N_9972,N_8741);
nand U11022 (N_11022,N_9196,N_8005);
nand U11023 (N_11023,N_8116,N_8526);
xnor U11024 (N_11024,N_9745,N_9000);
nand U11025 (N_11025,N_8271,N_8791);
nand U11026 (N_11026,N_8511,N_9428);
xnor U11027 (N_11027,N_8224,N_9254);
nor U11028 (N_11028,N_8807,N_8361);
and U11029 (N_11029,N_9440,N_9151);
and U11030 (N_11030,N_9261,N_8802);
and U11031 (N_11031,N_9293,N_8285);
or U11032 (N_11032,N_8050,N_9947);
and U11033 (N_11033,N_8205,N_9178);
xor U11034 (N_11034,N_8815,N_8035);
and U11035 (N_11035,N_8807,N_9209);
or U11036 (N_11036,N_9967,N_9693);
or U11037 (N_11037,N_8930,N_8362);
and U11038 (N_11038,N_9590,N_8519);
nor U11039 (N_11039,N_9924,N_9500);
xor U11040 (N_11040,N_9710,N_8291);
nor U11041 (N_11041,N_9742,N_8052);
nand U11042 (N_11042,N_8040,N_9752);
xor U11043 (N_11043,N_9267,N_9337);
nand U11044 (N_11044,N_9074,N_8364);
nand U11045 (N_11045,N_9318,N_9465);
and U11046 (N_11046,N_9754,N_9190);
nor U11047 (N_11047,N_8970,N_8700);
xor U11048 (N_11048,N_8384,N_9657);
xnor U11049 (N_11049,N_9364,N_8748);
nor U11050 (N_11050,N_9997,N_8830);
nand U11051 (N_11051,N_8208,N_8640);
and U11052 (N_11052,N_8052,N_8054);
nand U11053 (N_11053,N_9313,N_9911);
xnor U11054 (N_11054,N_9653,N_9210);
nand U11055 (N_11055,N_9086,N_9348);
nor U11056 (N_11056,N_8125,N_8367);
nor U11057 (N_11057,N_9695,N_9295);
and U11058 (N_11058,N_9321,N_8317);
xnor U11059 (N_11059,N_8325,N_9199);
nor U11060 (N_11060,N_9365,N_8060);
and U11061 (N_11061,N_9328,N_9073);
nor U11062 (N_11062,N_8717,N_9886);
nand U11063 (N_11063,N_9730,N_9941);
xor U11064 (N_11064,N_9606,N_9617);
or U11065 (N_11065,N_8604,N_8665);
nand U11066 (N_11066,N_8509,N_9397);
nor U11067 (N_11067,N_9561,N_9515);
or U11068 (N_11068,N_8115,N_9779);
and U11069 (N_11069,N_8022,N_9778);
xor U11070 (N_11070,N_9411,N_8946);
or U11071 (N_11071,N_9666,N_8957);
nor U11072 (N_11072,N_8041,N_9261);
and U11073 (N_11073,N_9389,N_8968);
nand U11074 (N_11074,N_9969,N_9200);
and U11075 (N_11075,N_8837,N_9562);
nor U11076 (N_11076,N_8143,N_8991);
xor U11077 (N_11077,N_9351,N_8955);
nand U11078 (N_11078,N_8316,N_9522);
nor U11079 (N_11079,N_8633,N_8317);
xnor U11080 (N_11080,N_9630,N_9980);
or U11081 (N_11081,N_9992,N_8648);
nor U11082 (N_11082,N_8893,N_9986);
or U11083 (N_11083,N_9065,N_8421);
xor U11084 (N_11084,N_8730,N_9945);
xor U11085 (N_11085,N_8170,N_9808);
or U11086 (N_11086,N_9192,N_8772);
nor U11087 (N_11087,N_9953,N_8430);
xnor U11088 (N_11088,N_8229,N_9933);
or U11089 (N_11089,N_8444,N_9810);
nand U11090 (N_11090,N_8104,N_9009);
nor U11091 (N_11091,N_9431,N_9720);
or U11092 (N_11092,N_8168,N_8699);
nor U11093 (N_11093,N_9021,N_9834);
nor U11094 (N_11094,N_9237,N_9008);
xor U11095 (N_11095,N_9638,N_8278);
or U11096 (N_11096,N_9537,N_9387);
xor U11097 (N_11097,N_8445,N_8813);
xnor U11098 (N_11098,N_9559,N_8369);
xor U11099 (N_11099,N_8307,N_8501);
and U11100 (N_11100,N_9057,N_9697);
xnor U11101 (N_11101,N_9305,N_9250);
xnor U11102 (N_11102,N_8743,N_9295);
or U11103 (N_11103,N_8663,N_9973);
nor U11104 (N_11104,N_9200,N_8942);
or U11105 (N_11105,N_9446,N_8101);
xnor U11106 (N_11106,N_8192,N_8853);
nor U11107 (N_11107,N_9701,N_8510);
and U11108 (N_11108,N_9972,N_9984);
or U11109 (N_11109,N_9177,N_8203);
and U11110 (N_11110,N_8685,N_8563);
or U11111 (N_11111,N_9780,N_8644);
nand U11112 (N_11112,N_8736,N_9203);
or U11113 (N_11113,N_8864,N_8267);
xor U11114 (N_11114,N_8098,N_8477);
xor U11115 (N_11115,N_8208,N_9140);
and U11116 (N_11116,N_8221,N_9752);
and U11117 (N_11117,N_9724,N_9996);
and U11118 (N_11118,N_9292,N_8851);
and U11119 (N_11119,N_9821,N_8437);
and U11120 (N_11120,N_9598,N_8840);
xnor U11121 (N_11121,N_9648,N_9454);
xnor U11122 (N_11122,N_8468,N_9390);
xnor U11123 (N_11123,N_9010,N_8670);
or U11124 (N_11124,N_9646,N_8668);
or U11125 (N_11125,N_8903,N_9873);
and U11126 (N_11126,N_8443,N_9306);
nor U11127 (N_11127,N_8206,N_9086);
nand U11128 (N_11128,N_8753,N_8343);
nand U11129 (N_11129,N_8483,N_8439);
or U11130 (N_11130,N_8841,N_8953);
xnor U11131 (N_11131,N_9602,N_9359);
nor U11132 (N_11132,N_8141,N_8469);
or U11133 (N_11133,N_9581,N_8912);
nand U11134 (N_11134,N_8739,N_9806);
or U11135 (N_11135,N_9272,N_8553);
nand U11136 (N_11136,N_8863,N_9877);
xor U11137 (N_11137,N_8244,N_8491);
or U11138 (N_11138,N_9047,N_9069);
nor U11139 (N_11139,N_8454,N_9570);
or U11140 (N_11140,N_8865,N_8619);
and U11141 (N_11141,N_8761,N_9913);
nor U11142 (N_11142,N_8936,N_9831);
or U11143 (N_11143,N_8502,N_8756);
nor U11144 (N_11144,N_8820,N_9163);
or U11145 (N_11145,N_8821,N_9178);
nand U11146 (N_11146,N_8708,N_8912);
and U11147 (N_11147,N_9112,N_9455);
nand U11148 (N_11148,N_8630,N_9831);
and U11149 (N_11149,N_9363,N_8205);
or U11150 (N_11150,N_9956,N_9985);
xnor U11151 (N_11151,N_8498,N_8629);
nand U11152 (N_11152,N_8196,N_9612);
and U11153 (N_11153,N_9299,N_9664);
and U11154 (N_11154,N_8457,N_9325);
nand U11155 (N_11155,N_8615,N_8330);
or U11156 (N_11156,N_9932,N_8569);
xnor U11157 (N_11157,N_8553,N_9357);
nor U11158 (N_11158,N_9262,N_8443);
and U11159 (N_11159,N_8413,N_9777);
nor U11160 (N_11160,N_9420,N_8514);
nor U11161 (N_11161,N_8961,N_9111);
nor U11162 (N_11162,N_8179,N_8676);
nor U11163 (N_11163,N_9760,N_8891);
or U11164 (N_11164,N_9480,N_8820);
nor U11165 (N_11165,N_8586,N_9372);
nand U11166 (N_11166,N_8456,N_9343);
xnor U11167 (N_11167,N_8370,N_9834);
nor U11168 (N_11168,N_8999,N_9149);
nand U11169 (N_11169,N_8161,N_9671);
or U11170 (N_11170,N_9923,N_8600);
nand U11171 (N_11171,N_9526,N_9289);
nor U11172 (N_11172,N_9730,N_9502);
nor U11173 (N_11173,N_8970,N_8536);
nor U11174 (N_11174,N_9285,N_9516);
nand U11175 (N_11175,N_8276,N_8212);
and U11176 (N_11176,N_9987,N_8592);
nand U11177 (N_11177,N_8025,N_8232);
and U11178 (N_11178,N_9498,N_9071);
nand U11179 (N_11179,N_9858,N_8073);
nor U11180 (N_11180,N_9211,N_8895);
and U11181 (N_11181,N_9593,N_8720);
or U11182 (N_11182,N_8616,N_8800);
and U11183 (N_11183,N_8707,N_9587);
nand U11184 (N_11184,N_9187,N_8848);
and U11185 (N_11185,N_9556,N_8889);
nand U11186 (N_11186,N_9926,N_9471);
and U11187 (N_11187,N_9799,N_8126);
nor U11188 (N_11188,N_9432,N_8359);
or U11189 (N_11189,N_8820,N_8729);
nand U11190 (N_11190,N_8432,N_9694);
xor U11191 (N_11191,N_9403,N_8809);
and U11192 (N_11192,N_9048,N_8505);
xor U11193 (N_11193,N_8367,N_9848);
or U11194 (N_11194,N_9272,N_9744);
or U11195 (N_11195,N_9178,N_8966);
nor U11196 (N_11196,N_9433,N_8001);
or U11197 (N_11197,N_8940,N_8406);
nor U11198 (N_11198,N_9888,N_9403);
nor U11199 (N_11199,N_9643,N_8271);
or U11200 (N_11200,N_9952,N_9804);
xor U11201 (N_11201,N_9524,N_9828);
nand U11202 (N_11202,N_8791,N_8035);
and U11203 (N_11203,N_9013,N_8805);
and U11204 (N_11204,N_9604,N_8506);
nand U11205 (N_11205,N_8934,N_8126);
xnor U11206 (N_11206,N_9945,N_9350);
nand U11207 (N_11207,N_8092,N_8648);
xor U11208 (N_11208,N_9799,N_8383);
or U11209 (N_11209,N_8114,N_9296);
nor U11210 (N_11210,N_8797,N_9364);
and U11211 (N_11211,N_8276,N_8844);
nor U11212 (N_11212,N_9500,N_8255);
nand U11213 (N_11213,N_8245,N_8165);
nor U11214 (N_11214,N_8500,N_8726);
and U11215 (N_11215,N_9292,N_9194);
and U11216 (N_11216,N_9018,N_8454);
and U11217 (N_11217,N_9356,N_8535);
nand U11218 (N_11218,N_9472,N_8694);
xnor U11219 (N_11219,N_8833,N_8808);
nor U11220 (N_11220,N_9650,N_8671);
or U11221 (N_11221,N_8454,N_8031);
or U11222 (N_11222,N_8798,N_8490);
nand U11223 (N_11223,N_9059,N_8090);
and U11224 (N_11224,N_8678,N_9074);
nand U11225 (N_11225,N_9107,N_8123);
nand U11226 (N_11226,N_9631,N_8492);
xor U11227 (N_11227,N_9118,N_9957);
nand U11228 (N_11228,N_9400,N_8074);
and U11229 (N_11229,N_9142,N_9544);
nor U11230 (N_11230,N_9194,N_8019);
xnor U11231 (N_11231,N_9163,N_9817);
nor U11232 (N_11232,N_9624,N_9820);
and U11233 (N_11233,N_8047,N_9487);
nand U11234 (N_11234,N_8885,N_9071);
nor U11235 (N_11235,N_9582,N_8147);
or U11236 (N_11236,N_9855,N_8556);
xor U11237 (N_11237,N_8554,N_8677);
xnor U11238 (N_11238,N_9209,N_8705);
nand U11239 (N_11239,N_9117,N_8533);
xnor U11240 (N_11240,N_9191,N_8446);
nand U11241 (N_11241,N_8278,N_8240);
xor U11242 (N_11242,N_9469,N_8919);
xnor U11243 (N_11243,N_9481,N_9963);
xnor U11244 (N_11244,N_8599,N_9360);
nor U11245 (N_11245,N_9976,N_8505);
and U11246 (N_11246,N_9978,N_8510);
and U11247 (N_11247,N_9834,N_8560);
nand U11248 (N_11248,N_8253,N_8492);
xor U11249 (N_11249,N_9008,N_9569);
xnor U11250 (N_11250,N_9074,N_8547);
xnor U11251 (N_11251,N_9941,N_9065);
nor U11252 (N_11252,N_9337,N_8856);
or U11253 (N_11253,N_9069,N_8569);
nor U11254 (N_11254,N_8611,N_8612);
nand U11255 (N_11255,N_8267,N_8233);
and U11256 (N_11256,N_9032,N_9704);
or U11257 (N_11257,N_9494,N_9529);
and U11258 (N_11258,N_9272,N_8838);
and U11259 (N_11259,N_9264,N_9614);
xor U11260 (N_11260,N_9722,N_8029);
nand U11261 (N_11261,N_9775,N_8199);
nor U11262 (N_11262,N_9691,N_8553);
xnor U11263 (N_11263,N_9316,N_8375);
xnor U11264 (N_11264,N_8381,N_9480);
xor U11265 (N_11265,N_9483,N_8883);
xor U11266 (N_11266,N_8215,N_8060);
nand U11267 (N_11267,N_9781,N_8673);
nor U11268 (N_11268,N_9634,N_8499);
nor U11269 (N_11269,N_8838,N_8794);
xor U11270 (N_11270,N_8204,N_9262);
xnor U11271 (N_11271,N_8289,N_8810);
or U11272 (N_11272,N_8657,N_8074);
and U11273 (N_11273,N_9532,N_9963);
nor U11274 (N_11274,N_9671,N_9533);
and U11275 (N_11275,N_8541,N_8848);
nor U11276 (N_11276,N_8605,N_9554);
and U11277 (N_11277,N_9913,N_8364);
and U11278 (N_11278,N_8066,N_9242);
nor U11279 (N_11279,N_8079,N_9704);
nand U11280 (N_11280,N_9656,N_8346);
nor U11281 (N_11281,N_9255,N_8898);
nor U11282 (N_11282,N_9813,N_8271);
and U11283 (N_11283,N_8974,N_9397);
nand U11284 (N_11284,N_8594,N_8557);
or U11285 (N_11285,N_9545,N_9343);
xnor U11286 (N_11286,N_8192,N_8873);
nor U11287 (N_11287,N_9290,N_8323);
and U11288 (N_11288,N_9407,N_8943);
and U11289 (N_11289,N_8936,N_8011);
or U11290 (N_11290,N_9392,N_8247);
and U11291 (N_11291,N_9850,N_9509);
and U11292 (N_11292,N_9396,N_8231);
nand U11293 (N_11293,N_9027,N_9978);
nor U11294 (N_11294,N_9282,N_8562);
and U11295 (N_11295,N_9871,N_8206);
nor U11296 (N_11296,N_8845,N_8548);
and U11297 (N_11297,N_8491,N_8181);
or U11298 (N_11298,N_9647,N_9255);
xnor U11299 (N_11299,N_9977,N_8253);
nand U11300 (N_11300,N_9831,N_8588);
nor U11301 (N_11301,N_9628,N_9378);
xnor U11302 (N_11302,N_9061,N_8594);
nor U11303 (N_11303,N_8602,N_8049);
xnor U11304 (N_11304,N_8276,N_9098);
and U11305 (N_11305,N_9172,N_8497);
xnor U11306 (N_11306,N_8168,N_8991);
nor U11307 (N_11307,N_8423,N_9848);
or U11308 (N_11308,N_8212,N_9585);
and U11309 (N_11309,N_8594,N_9485);
nand U11310 (N_11310,N_9244,N_9343);
and U11311 (N_11311,N_9486,N_9543);
or U11312 (N_11312,N_8579,N_8972);
xnor U11313 (N_11313,N_9928,N_9201);
or U11314 (N_11314,N_9982,N_8687);
nor U11315 (N_11315,N_8750,N_9407);
or U11316 (N_11316,N_9060,N_9526);
and U11317 (N_11317,N_8059,N_9913);
xor U11318 (N_11318,N_8772,N_9526);
or U11319 (N_11319,N_8000,N_8676);
and U11320 (N_11320,N_9935,N_8561);
nor U11321 (N_11321,N_9632,N_8066);
nor U11322 (N_11322,N_8690,N_9933);
xor U11323 (N_11323,N_9831,N_8185);
or U11324 (N_11324,N_8093,N_8539);
and U11325 (N_11325,N_8903,N_9089);
and U11326 (N_11326,N_8220,N_9361);
or U11327 (N_11327,N_8549,N_9558);
and U11328 (N_11328,N_8856,N_8441);
or U11329 (N_11329,N_8121,N_8729);
or U11330 (N_11330,N_9467,N_9399);
and U11331 (N_11331,N_8412,N_8220);
and U11332 (N_11332,N_8881,N_8541);
and U11333 (N_11333,N_8194,N_9773);
and U11334 (N_11334,N_8521,N_8771);
nor U11335 (N_11335,N_8849,N_8471);
or U11336 (N_11336,N_8667,N_8859);
and U11337 (N_11337,N_9886,N_9274);
xor U11338 (N_11338,N_9878,N_9132);
xor U11339 (N_11339,N_9504,N_9024);
or U11340 (N_11340,N_9795,N_8061);
nand U11341 (N_11341,N_9680,N_9116);
xnor U11342 (N_11342,N_9826,N_8189);
and U11343 (N_11343,N_8046,N_8226);
xnor U11344 (N_11344,N_8083,N_8869);
and U11345 (N_11345,N_8361,N_9557);
and U11346 (N_11346,N_8744,N_9360);
nor U11347 (N_11347,N_9571,N_8696);
and U11348 (N_11348,N_9529,N_8725);
xor U11349 (N_11349,N_8739,N_9292);
nand U11350 (N_11350,N_8314,N_9631);
nor U11351 (N_11351,N_9424,N_9183);
or U11352 (N_11352,N_9259,N_9884);
xnor U11353 (N_11353,N_9537,N_9160);
or U11354 (N_11354,N_9129,N_8920);
and U11355 (N_11355,N_9860,N_9581);
nand U11356 (N_11356,N_8104,N_8837);
xor U11357 (N_11357,N_9363,N_9388);
and U11358 (N_11358,N_9423,N_9630);
or U11359 (N_11359,N_9817,N_9916);
nor U11360 (N_11360,N_9519,N_9593);
nand U11361 (N_11361,N_9542,N_9606);
or U11362 (N_11362,N_8542,N_8455);
and U11363 (N_11363,N_8298,N_9848);
or U11364 (N_11364,N_9884,N_9213);
or U11365 (N_11365,N_8177,N_9634);
and U11366 (N_11366,N_8249,N_9768);
xnor U11367 (N_11367,N_8891,N_9803);
nor U11368 (N_11368,N_8613,N_9760);
xnor U11369 (N_11369,N_9869,N_8967);
xor U11370 (N_11370,N_8256,N_8579);
or U11371 (N_11371,N_8145,N_9926);
and U11372 (N_11372,N_8019,N_9908);
and U11373 (N_11373,N_9851,N_9414);
xnor U11374 (N_11374,N_9229,N_8329);
or U11375 (N_11375,N_8617,N_9643);
nand U11376 (N_11376,N_9031,N_8844);
nor U11377 (N_11377,N_9034,N_8626);
or U11378 (N_11378,N_8292,N_9826);
nand U11379 (N_11379,N_9253,N_9814);
and U11380 (N_11380,N_9495,N_8927);
xor U11381 (N_11381,N_9444,N_9109);
nand U11382 (N_11382,N_9587,N_9841);
nand U11383 (N_11383,N_8038,N_9310);
xnor U11384 (N_11384,N_9478,N_9207);
nand U11385 (N_11385,N_8507,N_9279);
and U11386 (N_11386,N_8514,N_9991);
nor U11387 (N_11387,N_9232,N_9664);
or U11388 (N_11388,N_8848,N_9140);
nor U11389 (N_11389,N_9141,N_8793);
or U11390 (N_11390,N_8244,N_8431);
nand U11391 (N_11391,N_9149,N_9086);
and U11392 (N_11392,N_9703,N_9169);
nor U11393 (N_11393,N_8104,N_8614);
xor U11394 (N_11394,N_9939,N_9016);
nand U11395 (N_11395,N_9371,N_9644);
or U11396 (N_11396,N_9815,N_8983);
nor U11397 (N_11397,N_8351,N_8633);
xnor U11398 (N_11398,N_9105,N_9057);
and U11399 (N_11399,N_9851,N_8247);
and U11400 (N_11400,N_9602,N_9050);
and U11401 (N_11401,N_9428,N_8872);
nand U11402 (N_11402,N_8824,N_9922);
nand U11403 (N_11403,N_9613,N_9305);
nand U11404 (N_11404,N_8330,N_8690);
nand U11405 (N_11405,N_9920,N_9362);
nor U11406 (N_11406,N_9722,N_8938);
nand U11407 (N_11407,N_9509,N_8824);
and U11408 (N_11408,N_9572,N_9579);
xor U11409 (N_11409,N_8723,N_8889);
or U11410 (N_11410,N_9183,N_8808);
or U11411 (N_11411,N_8899,N_8106);
nand U11412 (N_11412,N_9801,N_9253);
or U11413 (N_11413,N_9985,N_8347);
xor U11414 (N_11414,N_8453,N_8309);
nand U11415 (N_11415,N_9513,N_8553);
nor U11416 (N_11416,N_9565,N_9685);
and U11417 (N_11417,N_9208,N_9786);
nand U11418 (N_11418,N_9214,N_9850);
nand U11419 (N_11419,N_8212,N_8878);
nor U11420 (N_11420,N_8417,N_8936);
nor U11421 (N_11421,N_8171,N_9624);
and U11422 (N_11422,N_8387,N_9701);
and U11423 (N_11423,N_9527,N_9390);
or U11424 (N_11424,N_9156,N_9088);
or U11425 (N_11425,N_8643,N_8344);
or U11426 (N_11426,N_9607,N_8977);
nor U11427 (N_11427,N_8427,N_9781);
and U11428 (N_11428,N_9524,N_8620);
nor U11429 (N_11429,N_9069,N_9035);
or U11430 (N_11430,N_8027,N_8780);
and U11431 (N_11431,N_8054,N_9676);
nor U11432 (N_11432,N_8328,N_8614);
nand U11433 (N_11433,N_8859,N_8339);
nand U11434 (N_11434,N_9334,N_9236);
xnor U11435 (N_11435,N_8292,N_8515);
xnor U11436 (N_11436,N_8047,N_8142);
nand U11437 (N_11437,N_8305,N_8956);
or U11438 (N_11438,N_9016,N_8251);
xor U11439 (N_11439,N_8485,N_8726);
nand U11440 (N_11440,N_9768,N_8843);
or U11441 (N_11441,N_8152,N_8759);
xnor U11442 (N_11442,N_8578,N_9535);
nor U11443 (N_11443,N_9112,N_9151);
nor U11444 (N_11444,N_8837,N_9922);
nor U11445 (N_11445,N_9553,N_9232);
xor U11446 (N_11446,N_8393,N_8366);
nand U11447 (N_11447,N_9293,N_9098);
or U11448 (N_11448,N_9451,N_8084);
or U11449 (N_11449,N_9454,N_8642);
xor U11450 (N_11450,N_8145,N_9124);
or U11451 (N_11451,N_8275,N_8632);
nor U11452 (N_11452,N_9289,N_8999);
nor U11453 (N_11453,N_8195,N_8179);
and U11454 (N_11454,N_9928,N_8579);
nand U11455 (N_11455,N_8177,N_8096);
xor U11456 (N_11456,N_9591,N_8667);
nor U11457 (N_11457,N_9734,N_9316);
nor U11458 (N_11458,N_8565,N_9214);
xnor U11459 (N_11459,N_8748,N_8333);
or U11460 (N_11460,N_9977,N_9214);
xor U11461 (N_11461,N_9782,N_8819);
or U11462 (N_11462,N_8706,N_8845);
or U11463 (N_11463,N_8435,N_8325);
and U11464 (N_11464,N_8663,N_9606);
or U11465 (N_11465,N_9116,N_9597);
nand U11466 (N_11466,N_9283,N_9667);
xnor U11467 (N_11467,N_8435,N_8022);
xor U11468 (N_11468,N_9857,N_8728);
nand U11469 (N_11469,N_8849,N_8818);
and U11470 (N_11470,N_9953,N_8466);
and U11471 (N_11471,N_8460,N_9951);
nor U11472 (N_11472,N_9080,N_9714);
or U11473 (N_11473,N_8981,N_8580);
or U11474 (N_11474,N_8176,N_9945);
or U11475 (N_11475,N_8493,N_9778);
or U11476 (N_11476,N_8729,N_8179);
nor U11477 (N_11477,N_8954,N_9896);
nand U11478 (N_11478,N_8301,N_8047);
or U11479 (N_11479,N_8662,N_9377);
or U11480 (N_11480,N_8973,N_8210);
nor U11481 (N_11481,N_8746,N_8435);
or U11482 (N_11482,N_9304,N_9508);
nand U11483 (N_11483,N_9565,N_9638);
and U11484 (N_11484,N_9643,N_8214);
nor U11485 (N_11485,N_8019,N_8536);
nand U11486 (N_11486,N_9404,N_8154);
xor U11487 (N_11487,N_8810,N_9859);
nand U11488 (N_11488,N_8204,N_8111);
and U11489 (N_11489,N_8333,N_8764);
xor U11490 (N_11490,N_8144,N_9558);
nor U11491 (N_11491,N_8566,N_8037);
xor U11492 (N_11492,N_9911,N_8641);
nor U11493 (N_11493,N_8987,N_9764);
or U11494 (N_11494,N_8015,N_8773);
nor U11495 (N_11495,N_9065,N_9950);
xor U11496 (N_11496,N_8495,N_8607);
nor U11497 (N_11497,N_8797,N_9093);
and U11498 (N_11498,N_9001,N_9819);
nand U11499 (N_11499,N_9021,N_9772);
or U11500 (N_11500,N_8445,N_8414);
nor U11501 (N_11501,N_9873,N_9477);
xor U11502 (N_11502,N_8639,N_9334);
nor U11503 (N_11503,N_9371,N_8984);
and U11504 (N_11504,N_8942,N_9094);
nor U11505 (N_11505,N_8620,N_9704);
nand U11506 (N_11506,N_9398,N_9745);
nand U11507 (N_11507,N_8793,N_8799);
and U11508 (N_11508,N_8339,N_8871);
nand U11509 (N_11509,N_8759,N_8964);
nor U11510 (N_11510,N_8603,N_9025);
nor U11511 (N_11511,N_8308,N_8255);
nand U11512 (N_11512,N_9343,N_8709);
nand U11513 (N_11513,N_8971,N_8317);
xnor U11514 (N_11514,N_8983,N_9747);
xnor U11515 (N_11515,N_8029,N_9652);
nor U11516 (N_11516,N_9508,N_9152);
nand U11517 (N_11517,N_8969,N_9600);
nor U11518 (N_11518,N_8350,N_9252);
xnor U11519 (N_11519,N_8105,N_9319);
xnor U11520 (N_11520,N_9473,N_8991);
nand U11521 (N_11521,N_9221,N_8551);
and U11522 (N_11522,N_8366,N_9047);
or U11523 (N_11523,N_9706,N_9574);
or U11524 (N_11524,N_8128,N_8209);
xor U11525 (N_11525,N_8024,N_8813);
xor U11526 (N_11526,N_8506,N_8279);
xor U11527 (N_11527,N_8213,N_8948);
nand U11528 (N_11528,N_9364,N_9386);
xor U11529 (N_11529,N_8111,N_8672);
or U11530 (N_11530,N_8781,N_8959);
xor U11531 (N_11531,N_8886,N_8095);
or U11532 (N_11532,N_9530,N_8999);
nand U11533 (N_11533,N_9726,N_8647);
nand U11534 (N_11534,N_9370,N_9904);
nor U11535 (N_11535,N_8781,N_9638);
nor U11536 (N_11536,N_8642,N_8471);
nand U11537 (N_11537,N_8272,N_8012);
nand U11538 (N_11538,N_9665,N_8849);
nor U11539 (N_11539,N_8475,N_8479);
and U11540 (N_11540,N_9301,N_9719);
nor U11541 (N_11541,N_8261,N_8371);
or U11542 (N_11542,N_8834,N_9145);
and U11543 (N_11543,N_9298,N_9384);
nand U11544 (N_11544,N_9249,N_8732);
nand U11545 (N_11545,N_8785,N_8937);
xnor U11546 (N_11546,N_8816,N_9590);
or U11547 (N_11547,N_9533,N_9221);
or U11548 (N_11548,N_8457,N_8413);
and U11549 (N_11549,N_8515,N_8152);
nand U11550 (N_11550,N_8800,N_9451);
nor U11551 (N_11551,N_8651,N_8664);
or U11552 (N_11552,N_8698,N_9680);
nand U11553 (N_11553,N_9758,N_9684);
nand U11554 (N_11554,N_8472,N_8148);
xor U11555 (N_11555,N_9006,N_8989);
nand U11556 (N_11556,N_9198,N_9890);
xnor U11557 (N_11557,N_9707,N_9000);
nand U11558 (N_11558,N_9721,N_8992);
nand U11559 (N_11559,N_9787,N_8831);
or U11560 (N_11560,N_9930,N_8144);
xor U11561 (N_11561,N_9590,N_9781);
nor U11562 (N_11562,N_8106,N_8662);
nand U11563 (N_11563,N_8882,N_9435);
nor U11564 (N_11564,N_8189,N_8404);
nor U11565 (N_11565,N_9351,N_8911);
nand U11566 (N_11566,N_8760,N_8327);
or U11567 (N_11567,N_8556,N_9515);
and U11568 (N_11568,N_9370,N_8709);
and U11569 (N_11569,N_8513,N_8447);
and U11570 (N_11570,N_8660,N_8555);
or U11571 (N_11571,N_9409,N_8852);
and U11572 (N_11572,N_9525,N_8924);
nor U11573 (N_11573,N_8211,N_8092);
nor U11574 (N_11574,N_9548,N_9192);
nand U11575 (N_11575,N_9566,N_8208);
xnor U11576 (N_11576,N_8760,N_9111);
or U11577 (N_11577,N_8807,N_9428);
nand U11578 (N_11578,N_8594,N_9735);
nand U11579 (N_11579,N_9928,N_8185);
and U11580 (N_11580,N_9166,N_8630);
or U11581 (N_11581,N_8328,N_9345);
nor U11582 (N_11582,N_8836,N_9233);
nor U11583 (N_11583,N_8250,N_8799);
nor U11584 (N_11584,N_9041,N_8253);
and U11585 (N_11585,N_9544,N_9499);
xnor U11586 (N_11586,N_8355,N_8117);
nand U11587 (N_11587,N_9398,N_8167);
or U11588 (N_11588,N_9756,N_9535);
nor U11589 (N_11589,N_9140,N_8622);
nand U11590 (N_11590,N_9913,N_8753);
xor U11591 (N_11591,N_8158,N_8200);
and U11592 (N_11592,N_8094,N_8422);
nor U11593 (N_11593,N_8146,N_8952);
xnor U11594 (N_11594,N_9585,N_9642);
or U11595 (N_11595,N_9179,N_9172);
or U11596 (N_11596,N_9045,N_9841);
and U11597 (N_11597,N_8109,N_9741);
nor U11598 (N_11598,N_8008,N_8687);
xor U11599 (N_11599,N_8801,N_9577);
nor U11600 (N_11600,N_9294,N_9074);
or U11601 (N_11601,N_8027,N_8595);
or U11602 (N_11602,N_9586,N_9097);
and U11603 (N_11603,N_8841,N_8828);
or U11604 (N_11604,N_8664,N_9227);
nor U11605 (N_11605,N_9472,N_9406);
and U11606 (N_11606,N_8460,N_8337);
nand U11607 (N_11607,N_9902,N_8097);
and U11608 (N_11608,N_8176,N_8119);
or U11609 (N_11609,N_9919,N_9272);
nand U11610 (N_11610,N_8855,N_9351);
nand U11611 (N_11611,N_8876,N_8990);
nand U11612 (N_11612,N_9589,N_9857);
nor U11613 (N_11613,N_9282,N_9954);
nor U11614 (N_11614,N_8663,N_9691);
or U11615 (N_11615,N_9460,N_9457);
nor U11616 (N_11616,N_8984,N_9258);
xor U11617 (N_11617,N_8425,N_8917);
nor U11618 (N_11618,N_8090,N_8114);
and U11619 (N_11619,N_8624,N_9798);
or U11620 (N_11620,N_8074,N_8028);
and U11621 (N_11621,N_9251,N_9978);
and U11622 (N_11622,N_8877,N_9508);
or U11623 (N_11623,N_8471,N_8826);
xor U11624 (N_11624,N_8265,N_8025);
nand U11625 (N_11625,N_8799,N_9050);
xnor U11626 (N_11626,N_9463,N_9198);
and U11627 (N_11627,N_9957,N_8920);
or U11628 (N_11628,N_9889,N_9514);
or U11629 (N_11629,N_9490,N_9356);
nor U11630 (N_11630,N_9047,N_9270);
or U11631 (N_11631,N_8355,N_8817);
nor U11632 (N_11632,N_9843,N_9308);
and U11633 (N_11633,N_9231,N_8900);
xor U11634 (N_11634,N_9304,N_9177);
nand U11635 (N_11635,N_9652,N_9103);
xor U11636 (N_11636,N_9342,N_8169);
nand U11637 (N_11637,N_8920,N_9639);
nor U11638 (N_11638,N_9233,N_9554);
or U11639 (N_11639,N_8194,N_9145);
xnor U11640 (N_11640,N_9985,N_9239);
and U11641 (N_11641,N_9416,N_9980);
or U11642 (N_11642,N_8800,N_9566);
xnor U11643 (N_11643,N_8333,N_8550);
nor U11644 (N_11644,N_9983,N_8737);
nand U11645 (N_11645,N_8683,N_8106);
nand U11646 (N_11646,N_8143,N_8481);
nand U11647 (N_11647,N_8953,N_8862);
nor U11648 (N_11648,N_9130,N_9221);
xnor U11649 (N_11649,N_9954,N_8416);
nand U11650 (N_11650,N_9160,N_8008);
or U11651 (N_11651,N_9477,N_8490);
nand U11652 (N_11652,N_8464,N_8143);
or U11653 (N_11653,N_9707,N_8360);
and U11654 (N_11654,N_9875,N_9178);
and U11655 (N_11655,N_9363,N_8401);
xnor U11656 (N_11656,N_9641,N_8446);
nor U11657 (N_11657,N_8849,N_8501);
nand U11658 (N_11658,N_9711,N_9094);
nand U11659 (N_11659,N_8712,N_8985);
and U11660 (N_11660,N_8029,N_9042);
or U11661 (N_11661,N_8739,N_8305);
nor U11662 (N_11662,N_9127,N_9735);
and U11663 (N_11663,N_8840,N_9569);
nand U11664 (N_11664,N_9198,N_9664);
xnor U11665 (N_11665,N_8611,N_9706);
nor U11666 (N_11666,N_8250,N_8581);
nor U11667 (N_11667,N_8490,N_9067);
and U11668 (N_11668,N_8468,N_9607);
or U11669 (N_11669,N_8573,N_8474);
xnor U11670 (N_11670,N_9869,N_8094);
and U11671 (N_11671,N_9629,N_8079);
xnor U11672 (N_11672,N_9813,N_8962);
xor U11673 (N_11673,N_9724,N_8332);
nand U11674 (N_11674,N_8730,N_8611);
or U11675 (N_11675,N_8478,N_8968);
nor U11676 (N_11676,N_8865,N_9804);
nor U11677 (N_11677,N_8810,N_8733);
nand U11678 (N_11678,N_9451,N_9751);
and U11679 (N_11679,N_9074,N_9854);
and U11680 (N_11680,N_8988,N_8497);
and U11681 (N_11681,N_9689,N_9738);
nor U11682 (N_11682,N_9823,N_8403);
nor U11683 (N_11683,N_8261,N_9220);
nand U11684 (N_11684,N_8349,N_9984);
nand U11685 (N_11685,N_9746,N_9254);
nand U11686 (N_11686,N_8975,N_8969);
nor U11687 (N_11687,N_8941,N_9980);
nor U11688 (N_11688,N_9464,N_8490);
nor U11689 (N_11689,N_9499,N_8680);
xor U11690 (N_11690,N_8732,N_9819);
nor U11691 (N_11691,N_9097,N_8871);
or U11692 (N_11692,N_9745,N_9546);
or U11693 (N_11693,N_9333,N_9611);
nand U11694 (N_11694,N_9263,N_8418);
nand U11695 (N_11695,N_8664,N_9111);
and U11696 (N_11696,N_8748,N_9722);
xnor U11697 (N_11697,N_9157,N_8512);
and U11698 (N_11698,N_9777,N_8532);
and U11699 (N_11699,N_8853,N_9961);
and U11700 (N_11700,N_8825,N_8475);
xnor U11701 (N_11701,N_9695,N_9385);
nand U11702 (N_11702,N_9679,N_9853);
nand U11703 (N_11703,N_9631,N_9482);
nand U11704 (N_11704,N_8089,N_9221);
nor U11705 (N_11705,N_9835,N_9111);
xnor U11706 (N_11706,N_9093,N_8645);
and U11707 (N_11707,N_8296,N_9682);
nand U11708 (N_11708,N_9214,N_9297);
nor U11709 (N_11709,N_9099,N_8978);
or U11710 (N_11710,N_9684,N_9066);
or U11711 (N_11711,N_9377,N_8945);
nand U11712 (N_11712,N_9416,N_8384);
nand U11713 (N_11713,N_9493,N_8897);
xor U11714 (N_11714,N_8302,N_9745);
nand U11715 (N_11715,N_8999,N_9099);
xor U11716 (N_11716,N_9420,N_9404);
or U11717 (N_11717,N_9417,N_8860);
nand U11718 (N_11718,N_9293,N_9445);
nor U11719 (N_11719,N_8028,N_8653);
and U11720 (N_11720,N_8537,N_8382);
xnor U11721 (N_11721,N_8455,N_8310);
and U11722 (N_11722,N_9797,N_9497);
or U11723 (N_11723,N_8914,N_8595);
nor U11724 (N_11724,N_8785,N_9070);
xnor U11725 (N_11725,N_8065,N_8313);
and U11726 (N_11726,N_8762,N_8032);
or U11727 (N_11727,N_9184,N_8371);
and U11728 (N_11728,N_8881,N_9878);
or U11729 (N_11729,N_9645,N_9246);
nor U11730 (N_11730,N_9937,N_9037);
and U11731 (N_11731,N_9535,N_9324);
nand U11732 (N_11732,N_9277,N_8596);
and U11733 (N_11733,N_9745,N_8272);
and U11734 (N_11734,N_9650,N_9219);
nor U11735 (N_11735,N_9760,N_9909);
nand U11736 (N_11736,N_8014,N_9493);
or U11737 (N_11737,N_9867,N_9073);
xor U11738 (N_11738,N_9238,N_9608);
xnor U11739 (N_11739,N_9605,N_9325);
nor U11740 (N_11740,N_8790,N_8410);
and U11741 (N_11741,N_9529,N_9621);
nand U11742 (N_11742,N_9647,N_9199);
and U11743 (N_11743,N_8252,N_8144);
xor U11744 (N_11744,N_8247,N_9843);
and U11745 (N_11745,N_9956,N_9912);
or U11746 (N_11746,N_8791,N_8860);
nor U11747 (N_11747,N_8982,N_8334);
and U11748 (N_11748,N_9789,N_8718);
or U11749 (N_11749,N_8633,N_8649);
and U11750 (N_11750,N_9666,N_8572);
or U11751 (N_11751,N_8733,N_9800);
and U11752 (N_11752,N_8998,N_9820);
and U11753 (N_11753,N_8130,N_8355);
or U11754 (N_11754,N_9981,N_8482);
nor U11755 (N_11755,N_8677,N_8799);
xnor U11756 (N_11756,N_8998,N_9281);
nor U11757 (N_11757,N_8353,N_9961);
nand U11758 (N_11758,N_8728,N_8709);
and U11759 (N_11759,N_9556,N_8370);
xnor U11760 (N_11760,N_9377,N_8613);
xnor U11761 (N_11761,N_8629,N_9211);
or U11762 (N_11762,N_9985,N_9476);
or U11763 (N_11763,N_8047,N_9753);
nand U11764 (N_11764,N_9768,N_8873);
and U11765 (N_11765,N_8497,N_9223);
or U11766 (N_11766,N_8474,N_8916);
xor U11767 (N_11767,N_9333,N_9377);
nor U11768 (N_11768,N_8430,N_9043);
nor U11769 (N_11769,N_9735,N_9870);
xor U11770 (N_11770,N_9696,N_8425);
xnor U11771 (N_11771,N_8539,N_8066);
and U11772 (N_11772,N_9306,N_9201);
nand U11773 (N_11773,N_8523,N_8950);
or U11774 (N_11774,N_9586,N_8629);
xor U11775 (N_11775,N_9044,N_9369);
and U11776 (N_11776,N_9899,N_8036);
and U11777 (N_11777,N_9985,N_9853);
nor U11778 (N_11778,N_9789,N_9310);
xnor U11779 (N_11779,N_9149,N_9627);
and U11780 (N_11780,N_9725,N_8533);
nand U11781 (N_11781,N_9264,N_9237);
and U11782 (N_11782,N_9906,N_9624);
or U11783 (N_11783,N_8783,N_8312);
or U11784 (N_11784,N_8608,N_9691);
and U11785 (N_11785,N_9758,N_9992);
nor U11786 (N_11786,N_9393,N_9203);
or U11787 (N_11787,N_8642,N_8222);
or U11788 (N_11788,N_8218,N_8069);
nand U11789 (N_11789,N_9590,N_8415);
or U11790 (N_11790,N_8017,N_9460);
nand U11791 (N_11791,N_9841,N_9748);
nand U11792 (N_11792,N_9558,N_8124);
or U11793 (N_11793,N_9613,N_8925);
nand U11794 (N_11794,N_9423,N_9967);
nand U11795 (N_11795,N_8262,N_9059);
or U11796 (N_11796,N_8119,N_9758);
or U11797 (N_11797,N_8666,N_8990);
nor U11798 (N_11798,N_8000,N_9073);
nand U11799 (N_11799,N_8170,N_8872);
and U11800 (N_11800,N_9797,N_8831);
or U11801 (N_11801,N_9144,N_9434);
and U11802 (N_11802,N_9216,N_8861);
and U11803 (N_11803,N_8660,N_8942);
nor U11804 (N_11804,N_9282,N_8000);
and U11805 (N_11805,N_8837,N_8166);
nand U11806 (N_11806,N_9795,N_8767);
nor U11807 (N_11807,N_9656,N_8218);
nor U11808 (N_11808,N_8707,N_9269);
nor U11809 (N_11809,N_8507,N_9855);
or U11810 (N_11810,N_9657,N_8514);
and U11811 (N_11811,N_8134,N_9784);
nand U11812 (N_11812,N_8353,N_9693);
xor U11813 (N_11813,N_9181,N_8144);
nor U11814 (N_11814,N_8032,N_9067);
or U11815 (N_11815,N_9194,N_8818);
or U11816 (N_11816,N_8626,N_8346);
or U11817 (N_11817,N_9692,N_9384);
and U11818 (N_11818,N_9561,N_9542);
and U11819 (N_11819,N_8380,N_8632);
xor U11820 (N_11820,N_8848,N_9835);
or U11821 (N_11821,N_9035,N_9472);
and U11822 (N_11822,N_8979,N_9659);
xor U11823 (N_11823,N_9192,N_9640);
nand U11824 (N_11824,N_9364,N_8709);
nand U11825 (N_11825,N_8359,N_8497);
or U11826 (N_11826,N_8630,N_9619);
nor U11827 (N_11827,N_8911,N_8917);
nor U11828 (N_11828,N_9643,N_9802);
nand U11829 (N_11829,N_8058,N_9745);
and U11830 (N_11830,N_8972,N_8211);
or U11831 (N_11831,N_9039,N_8115);
xnor U11832 (N_11832,N_9092,N_9929);
and U11833 (N_11833,N_9343,N_9386);
nand U11834 (N_11834,N_8211,N_8043);
nor U11835 (N_11835,N_9738,N_8828);
or U11836 (N_11836,N_8290,N_9437);
or U11837 (N_11837,N_8186,N_9149);
xnor U11838 (N_11838,N_8611,N_8978);
and U11839 (N_11839,N_9328,N_8803);
and U11840 (N_11840,N_9612,N_9046);
xor U11841 (N_11841,N_8252,N_8136);
and U11842 (N_11842,N_8480,N_9463);
nor U11843 (N_11843,N_8977,N_9980);
and U11844 (N_11844,N_8925,N_9323);
and U11845 (N_11845,N_9190,N_8890);
nand U11846 (N_11846,N_8014,N_9104);
and U11847 (N_11847,N_8941,N_8684);
nor U11848 (N_11848,N_9233,N_9053);
and U11849 (N_11849,N_8801,N_8178);
xor U11850 (N_11850,N_9489,N_9221);
nor U11851 (N_11851,N_9852,N_9007);
or U11852 (N_11852,N_8724,N_9712);
or U11853 (N_11853,N_8507,N_8746);
and U11854 (N_11854,N_9904,N_8435);
xnor U11855 (N_11855,N_9962,N_9452);
and U11856 (N_11856,N_8963,N_9009);
or U11857 (N_11857,N_9325,N_8603);
nor U11858 (N_11858,N_8997,N_8916);
and U11859 (N_11859,N_8316,N_8899);
or U11860 (N_11860,N_8258,N_8487);
or U11861 (N_11861,N_8555,N_9217);
nand U11862 (N_11862,N_8983,N_8237);
xnor U11863 (N_11863,N_8294,N_9594);
and U11864 (N_11864,N_8923,N_9199);
and U11865 (N_11865,N_9825,N_8832);
or U11866 (N_11866,N_9664,N_9156);
xnor U11867 (N_11867,N_9788,N_8475);
or U11868 (N_11868,N_9529,N_8263);
and U11869 (N_11869,N_8023,N_8363);
or U11870 (N_11870,N_9697,N_9595);
nor U11871 (N_11871,N_8037,N_8578);
nand U11872 (N_11872,N_8078,N_8893);
and U11873 (N_11873,N_8422,N_8580);
nand U11874 (N_11874,N_8037,N_8996);
xor U11875 (N_11875,N_9872,N_8809);
nor U11876 (N_11876,N_9893,N_9406);
or U11877 (N_11877,N_9646,N_8579);
xor U11878 (N_11878,N_9543,N_8874);
xnor U11879 (N_11879,N_9094,N_9936);
nor U11880 (N_11880,N_9808,N_8407);
xnor U11881 (N_11881,N_9009,N_9938);
or U11882 (N_11882,N_8344,N_8972);
nand U11883 (N_11883,N_8497,N_8734);
xnor U11884 (N_11884,N_9220,N_9247);
nand U11885 (N_11885,N_9554,N_8539);
or U11886 (N_11886,N_9116,N_8894);
nor U11887 (N_11887,N_8870,N_9172);
nor U11888 (N_11888,N_9848,N_9037);
nand U11889 (N_11889,N_8596,N_8407);
or U11890 (N_11890,N_9137,N_9876);
and U11891 (N_11891,N_9621,N_9006);
xor U11892 (N_11892,N_9029,N_8822);
and U11893 (N_11893,N_9927,N_9206);
or U11894 (N_11894,N_9262,N_8775);
or U11895 (N_11895,N_9930,N_9858);
nand U11896 (N_11896,N_8797,N_8097);
and U11897 (N_11897,N_9209,N_9601);
nand U11898 (N_11898,N_9120,N_8858);
nand U11899 (N_11899,N_8527,N_9227);
nand U11900 (N_11900,N_8533,N_8398);
nor U11901 (N_11901,N_9916,N_9411);
nand U11902 (N_11902,N_8976,N_8699);
nand U11903 (N_11903,N_8148,N_8646);
and U11904 (N_11904,N_8202,N_9793);
nand U11905 (N_11905,N_8465,N_9662);
xnor U11906 (N_11906,N_9602,N_9400);
or U11907 (N_11907,N_8106,N_8517);
xor U11908 (N_11908,N_8242,N_8928);
nor U11909 (N_11909,N_8045,N_9617);
and U11910 (N_11910,N_9479,N_9108);
xnor U11911 (N_11911,N_9405,N_8542);
nor U11912 (N_11912,N_9399,N_9577);
nand U11913 (N_11913,N_8916,N_8564);
nor U11914 (N_11914,N_8876,N_9253);
and U11915 (N_11915,N_8811,N_9945);
and U11916 (N_11916,N_9857,N_9591);
or U11917 (N_11917,N_8090,N_9328);
and U11918 (N_11918,N_9790,N_8704);
or U11919 (N_11919,N_9497,N_8610);
nor U11920 (N_11920,N_8727,N_8890);
or U11921 (N_11921,N_8478,N_9098);
xor U11922 (N_11922,N_8903,N_8097);
xnor U11923 (N_11923,N_9504,N_8723);
or U11924 (N_11924,N_8820,N_8506);
and U11925 (N_11925,N_8154,N_9959);
xnor U11926 (N_11926,N_9927,N_9758);
xor U11927 (N_11927,N_9062,N_9824);
xor U11928 (N_11928,N_9506,N_9238);
nor U11929 (N_11929,N_8361,N_9022);
and U11930 (N_11930,N_8422,N_9063);
xor U11931 (N_11931,N_8223,N_9816);
nor U11932 (N_11932,N_9809,N_9000);
or U11933 (N_11933,N_8892,N_8448);
nor U11934 (N_11934,N_9699,N_9567);
nor U11935 (N_11935,N_8408,N_8980);
nand U11936 (N_11936,N_8765,N_8680);
nand U11937 (N_11937,N_9098,N_9373);
and U11938 (N_11938,N_9273,N_9715);
nor U11939 (N_11939,N_8213,N_8368);
nor U11940 (N_11940,N_8742,N_9032);
or U11941 (N_11941,N_8836,N_9623);
or U11942 (N_11942,N_8934,N_8506);
nand U11943 (N_11943,N_9661,N_8114);
xor U11944 (N_11944,N_9460,N_8162);
nand U11945 (N_11945,N_9618,N_9034);
nor U11946 (N_11946,N_8681,N_8564);
xor U11947 (N_11947,N_9046,N_8012);
and U11948 (N_11948,N_8662,N_9807);
nand U11949 (N_11949,N_8004,N_8771);
nor U11950 (N_11950,N_8698,N_8876);
or U11951 (N_11951,N_8014,N_9761);
nor U11952 (N_11952,N_8743,N_9394);
nand U11953 (N_11953,N_8093,N_8678);
and U11954 (N_11954,N_9624,N_8090);
nor U11955 (N_11955,N_8474,N_8519);
nand U11956 (N_11956,N_8118,N_8271);
nand U11957 (N_11957,N_9789,N_8724);
nor U11958 (N_11958,N_8385,N_8334);
xor U11959 (N_11959,N_8844,N_8677);
nor U11960 (N_11960,N_8930,N_9246);
and U11961 (N_11961,N_8603,N_8939);
nand U11962 (N_11962,N_9341,N_9359);
or U11963 (N_11963,N_9292,N_9565);
or U11964 (N_11964,N_9694,N_8391);
xnor U11965 (N_11965,N_9830,N_9200);
xnor U11966 (N_11966,N_8278,N_8073);
nor U11967 (N_11967,N_9994,N_9285);
or U11968 (N_11968,N_8680,N_9372);
or U11969 (N_11969,N_9203,N_9633);
nand U11970 (N_11970,N_8518,N_8734);
nor U11971 (N_11971,N_9125,N_8624);
xnor U11972 (N_11972,N_9085,N_9132);
or U11973 (N_11973,N_8809,N_8080);
nand U11974 (N_11974,N_9878,N_9414);
nand U11975 (N_11975,N_9904,N_9402);
nand U11976 (N_11976,N_9566,N_8643);
xor U11977 (N_11977,N_9138,N_8668);
nor U11978 (N_11978,N_9219,N_9749);
and U11979 (N_11979,N_9857,N_9926);
nand U11980 (N_11980,N_9571,N_8691);
nand U11981 (N_11981,N_9692,N_8420);
nand U11982 (N_11982,N_8079,N_8800);
and U11983 (N_11983,N_8604,N_8313);
and U11984 (N_11984,N_9359,N_8782);
and U11985 (N_11985,N_9129,N_8313);
and U11986 (N_11986,N_8307,N_9574);
nand U11987 (N_11987,N_9186,N_8525);
nand U11988 (N_11988,N_9572,N_9003);
xor U11989 (N_11989,N_8192,N_8287);
nand U11990 (N_11990,N_8258,N_8155);
nor U11991 (N_11991,N_8544,N_9924);
and U11992 (N_11992,N_8469,N_9921);
xnor U11993 (N_11993,N_8309,N_8071);
xnor U11994 (N_11994,N_9658,N_8490);
nand U11995 (N_11995,N_8999,N_9632);
nand U11996 (N_11996,N_9749,N_9740);
nand U11997 (N_11997,N_9616,N_8590);
nor U11998 (N_11998,N_8682,N_9285);
nor U11999 (N_11999,N_9725,N_8188);
xor U12000 (N_12000,N_10750,N_10204);
nor U12001 (N_12001,N_10517,N_10669);
nand U12002 (N_12002,N_10234,N_10846);
and U12003 (N_12003,N_11828,N_11370);
or U12004 (N_12004,N_11315,N_11490);
and U12005 (N_12005,N_11641,N_10504);
or U12006 (N_12006,N_10715,N_11115);
or U12007 (N_12007,N_10957,N_10743);
nand U12008 (N_12008,N_10171,N_10326);
nand U12009 (N_12009,N_11918,N_10036);
xnor U12010 (N_12010,N_11710,N_10488);
or U12011 (N_12011,N_10191,N_10676);
xor U12012 (N_12012,N_10105,N_10694);
nor U12013 (N_12013,N_11708,N_10052);
nand U12014 (N_12014,N_11645,N_10128);
and U12015 (N_12015,N_11650,N_11247);
nand U12016 (N_12016,N_11352,N_11427);
and U12017 (N_12017,N_11254,N_10018);
nor U12018 (N_12018,N_11736,N_11237);
or U12019 (N_12019,N_11627,N_11465);
nand U12020 (N_12020,N_11161,N_11099);
nand U12021 (N_12021,N_10997,N_11761);
and U12022 (N_12022,N_10027,N_11114);
or U12023 (N_12023,N_10183,N_10355);
nor U12024 (N_12024,N_10535,N_10524);
or U12025 (N_12025,N_10042,N_11872);
and U12026 (N_12026,N_10407,N_10713);
nor U12027 (N_12027,N_11207,N_11258);
or U12028 (N_12028,N_11299,N_10554);
and U12029 (N_12029,N_10124,N_11076);
or U12030 (N_12030,N_11686,N_10097);
nor U12031 (N_12031,N_11524,N_10560);
and U12032 (N_12032,N_10531,N_11735);
and U12033 (N_12033,N_11950,N_11006);
and U12034 (N_12034,N_11663,N_10935);
and U12035 (N_12035,N_10207,N_10500);
or U12036 (N_12036,N_10521,N_11599);
nor U12037 (N_12037,N_10405,N_11265);
and U12038 (N_12038,N_11621,N_11907);
and U12039 (N_12039,N_11437,N_11540);
nor U12040 (N_12040,N_11833,N_10712);
nor U12041 (N_12041,N_11978,N_11184);
and U12042 (N_12042,N_10605,N_11267);
xor U12043 (N_12043,N_11008,N_11345);
nand U12044 (N_12044,N_10224,N_10248);
and U12045 (N_12045,N_10762,N_11638);
xnor U12046 (N_12046,N_11797,N_10785);
xor U12047 (N_12047,N_11232,N_11187);
or U12048 (N_12048,N_11609,N_10366);
and U12049 (N_12049,N_10084,N_11654);
nor U12050 (N_12050,N_11239,N_10928);
xnor U12051 (N_12051,N_11457,N_11805);
and U12052 (N_12052,N_10189,N_10037);
or U12053 (N_12053,N_10327,N_11477);
xor U12054 (N_12054,N_10000,N_11405);
or U12055 (N_12055,N_10100,N_10873);
and U12056 (N_12056,N_10122,N_11067);
nor U12057 (N_12057,N_10950,N_11618);
and U12058 (N_12058,N_11100,N_11139);
nand U12059 (N_12059,N_10158,N_11803);
or U12060 (N_12060,N_11070,N_10907);
nand U12061 (N_12061,N_11940,N_11052);
xnor U12062 (N_12062,N_10291,N_11857);
xnor U12063 (N_12063,N_11439,N_10969);
nor U12064 (N_12064,N_11440,N_11055);
and U12065 (N_12065,N_11140,N_10344);
and U12066 (N_12066,N_10684,N_11225);
or U12067 (N_12067,N_10832,N_10468);
xnor U12068 (N_12068,N_10369,N_10575);
nor U12069 (N_12069,N_10316,N_11616);
xnor U12070 (N_12070,N_11913,N_10401);
or U12071 (N_12071,N_10566,N_11269);
or U12072 (N_12072,N_11279,N_11531);
and U12073 (N_12073,N_11914,N_10467);
nor U12074 (N_12074,N_10686,N_11066);
and U12075 (N_12075,N_11051,N_11798);
and U12076 (N_12076,N_11335,N_10840);
nor U12077 (N_12077,N_10745,N_11189);
xor U12078 (N_12078,N_10254,N_10179);
nand U12079 (N_12079,N_10862,N_11271);
nand U12080 (N_12080,N_10809,N_11785);
and U12081 (N_12081,N_10173,N_10511);
xor U12082 (N_12082,N_10379,N_11569);
xor U12083 (N_12083,N_10077,N_10800);
nand U12084 (N_12084,N_11823,N_10081);
xor U12085 (N_12085,N_10239,N_11044);
xnor U12086 (N_12086,N_11580,N_10876);
and U12087 (N_12087,N_11520,N_11392);
or U12088 (N_12088,N_11473,N_11215);
or U12089 (N_12089,N_10583,N_11478);
xnor U12090 (N_12090,N_10614,N_10390);
nor U12091 (N_12091,N_10092,N_11202);
nor U12092 (N_12092,N_10573,N_11112);
xor U12093 (N_12093,N_11351,N_11741);
nand U12094 (N_12094,N_11018,N_11098);
nor U12095 (N_12095,N_11312,N_11211);
xor U12096 (N_12096,N_10044,N_10858);
or U12097 (N_12097,N_10340,N_11962);
or U12098 (N_12098,N_10587,N_10222);
xnor U12099 (N_12099,N_11314,N_10623);
nand U12100 (N_12100,N_11246,N_10424);
or U12101 (N_12101,N_11992,N_10240);
nor U12102 (N_12102,N_10600,N_11860);
nand U12103 (N_12103,N_11414,N_11298);
nand U12104 (N_12104,N_10104,N_10886);
and U12105 (N_12105,N_11159,N_10242);
nand U12106 (N_12106,N_10157,N_11623);
xor U12107 (N_12107,N_10164,N_11772);
and U12108 (N_12108,N_11585,N_10579);
and U12109 (N_12109,N_11373,N_10578);
nand U12110 (N_12110,N_11192,N_10720);
xor U12111 (N_12111,N_10402,N_10045);
or U12112 (N_12112,N_10759,N_11219);
xor U12113 (N_12113,N_11123,N_10910);
or U12114 (N_12114,N_11101,N_10082);
nand U12115 (N_12115,N_11594,N_11197);
xnor U12116 (N_12116,N_10079,N_10703);
nor U12117 (N_12117,N_10269,N_10760);
nand U12118 (N_12118,N_11777,N_10914);
nand U12119 (N_12119,N_10542,N_10046);
nand U12120 (N_12120,N_11989,N_10861);
and U12121 (N_12121,N_11086,N_10755);
nor U12122 (N_12122,N_10272,N_11723);
nor U12123 (N_12123,N_11206,N_10702);
nor U12124 (N_12124,N_10496,N_10048);
and U12125 (N_12125,N_10658,N_10475);
or U12126 (N_12126,N_11394,N_11261);
nor U12127 (N_12127,N_10252,N_10498);
nand U12128 (N_12128,N_11285,N_11304);
nor U12129 (N_12129,N_10491,N_10300);
nand U12130 (N_12130,N_10662,N_11297);
nor U12131 (N_12131,N_11276,N_10385);
or U12132 (N_12132,N_10533,N_11890);
nor U12133 (N_12133,N_11379,N_10106);
nor U12134 (N_12134,N_10210,N_11092);
or U12135 (N_12135,N_11631,N_11303);
and U12136 (N_12136,N_10732,N_10541);
or U12137 (N_12137,N_10228,N_10130);
nand U12138 (N_12138,N_10083,N_10411);
xor U12139 (N_12139,N_11482,N_11689);
nand U12140 (N_12140,N_11732,N_11849);
and U12141 (N_12141,N_10493,N_10434);
nand U12142 (N_12142,N_11886,N_11792);
nor U12143 (N_12143,N_10415,N_11449);
nor U12144 (N_12144,N_10992,N_11658);
xor U12145 (N_12145,N_11445,N_10911);
or U12146 (N_12146,N_11648,N_10453);
xnor U12147 (N_12147,N_10723,N_11718);
or U12148 (N_12148,N_11858,N_10386);
or U12149 (N_12149,N_10973,N_10552);
and U12150 (N_12150,N_11999,N_11391);
nand U12151 (N_12151,N_10038,N_10708);
nand U12152 (N_12152,N_10471,N_11701);
nor U12153 (N_12153,N_11005,N_11712);
nor U12154 (N_12154,N_11652,N_11894);
nand U12155 (N_12155,N_10089,N_11773);
or U12156 (N_12156,N_11775,N_11038);
nand U12157 (N_12157,N_10577,N_10982);
nand U12158 (N_12158,N_11063,N_11542);
xnor U12159 (N_12159,N_10636,N_11725);
nand U12160 (N_12160,N_10315,N_10019);
nand U12161 (N_12161,N_10430,N_11291);
nand U12162 (N_12162,N_11850,N_11330);
nand U12163 (N_12163,N_11558,N_11510);
nor U12164 (N_12164,N_10134,N_11240);
nor U12165 (N_12165,N_10514,N_10963);
and U12166 (N_12166,N_10435,N_11767);
and U12167 (N_12167,N_11488,N_11050);
nand U12168 (N_12168,N_10264,N_10879);
xor U12169 (N_12169,N_11132,N_11548);
or U12170 (N_12170,N_11015,N_11178);
and U12171 (N_12171,N_10867,N_10767);
nor U12172 (N_12172,N_11948,N_10007);
or U12173 (N_12173,N_10944,N_10329);
and U12174 (N_12174,N_11353,N_11912);
nand U12175 (N_12175,N_10241,N_10141);
nor U12176 (N_12176,N_10748,N_10024);
nor U12177 (N_12177,N_11619,N_11466);
and U12178 (N_12178,N_10547,N_11952);
or U12179 (N_12179,N_11447,N_11576);
xnor U12180 (N_12180,N_11892,N_10463);
nand U12181 (N_12181,N_10103,N_11878);
or U12182 (N_12182,N_10393,N_11643);
nor U12183 (N_12183,N_11471,N_10129);
or U12184 (N_12184,N_11980,N_11448);
xor U12185 (N_12185,N_10165,N_10839);
nand U12186 (N_12186,N_11518,N_10472);
nor U12187 (N_12187,N_11917,N_11231);
or U12188 (N_12188,N_10348,N_10659);
xnor U12189 (N_12189,N_11145,N_10529);
xnor U12190 (N_12190,N_10645,N_11400);
or U12191 (N_12191,N_11812,N_10070);
xnor U12192 (N_12192,N_11719,N_11093);
and U12193 (N_12193,N_11410,N_10449);
nor U12194 (N_12194,N_10816,N_10553);
and U12195 (N_12195,N_11456,N_11757);
nand U12196 (N_12196,N_11097,N_10352);
xnor U12197 (N_12197,N_11366,N_11257);
or U12198 (N_12198,N_11674,N_10971);
and U12199 (N_12199,N_10526,N_10318);
nand U12200 (N_12200,N_10328,N_11613);
nor U12201 (N_12201,N_11975,N_11581);
and U12202 (N_12202,N_10633,N_10267);
xor U12203 (N_12203,N_10069,N_10829);
or U12204 (N_12204,N_11561,N_11896);
xor U12205 (N_12205,N_11227,N_10375);
nor U12206 (N_12206,N_11056,N_10559);
nand U12207 (N_12207,N_10395,N_11393);
nor U12208 (N_12208,N_11997,N_10683);
and U12209 (N_12209,N_11588,N_10392);
or U12210 (N_12210,N_11446,N_10638);
and U12211 (N_12211,N_11344,N_11452);
nor U12212 (N_12212,N_11504,N_11855);
or U12213 (N_12213,N_11769,N_10656);
nand U12214 (N_12214,N_11944,N_10934);
and U12215 (N_12215,N_10906,N_10570);
and U12216 (N_12216,N_11799,N_10296);
nand U12217 (N_12217,N_11739,N_10590);
or U12218 (N_12218,N_11001,N_10032);
or U12219 (N_12219,N_10235,N_11497);
nand U12220 (N_12220,N_11234,N_10855);
or U12221 (N_12221,N_11004,N_10075);
nor U12222 (N_12222,N_11626,N_10029);
xor U12223 (N_12223,N_10953,N_11983);
nand U12224 (N_12224,N_11200,N_11483);
xnor U12225 (N_12225,N_10078,N_10895);
nor U12226 (N_12226,N_11970,N_11957);
and U12227 (N_12227,N_11859,N_10637);
xor U12228 (N_12228,N_11696,N_11876);
and U12229 (N_12229,N_11186,N_11527);
nand U12230 (N_12230,N_11821,N_10875);
and U12231 (N_12231,N_11933,N_11172);
nor U12232 (N_12232,N_10331,N_10890);
nor U12233 (N_12233,N_10783,N_11880);
or U12234 (N_12234,N_11310,N_10260);
nand U12235 (N_12235,N_11791,N_11094);
nand U12236 (N_12236,N_10006,N_11426);
or U12237 (N_12237,N_10850,N_10295);
xnor U12238 (N_12238,N_10555,N_11176);
xor U12239 (N_12239,N_11517,N_10887);
or U12240 (N_12240,N_10464,N_10143);
nor U12241 (N_12241,N_11287,N_11195);
xor U12242 (N_12242,N_11943,N_11721);
nand U12243 (N_12243,N_10247,N_10818);
nand U12244 (N_12244,N_10916,N_10279);
and U12245 (N_12245,N_10212,N_11144);
or U12246 (N_12246,N_10305,N_10287);
or U12247 (N_12247,N_11556,N_10571);
and U12248 (N_12248,N_11358,N_10396);
xnor U12249 (N_12249,N_10093,N_10619);
and U12250 (N_12250,N_10400,N_11700);
and U12251 (N_12251,N_10330,N_11143);
xnor U12252 (N_12252,N_10642,N_11407);
nand U12253 (N_12253,N_10597,N_10624);
or U12254 (N_12254,N_10478,N_11945);
xor U12255 (N_12255,N_11503,N_11692);
or U12256 (N_12256,N_10409,N_10803);
xnor U12257 (N_12257,N_11307,N_11031);
xnor U12258 (N_12258,N_11549,N_10815);
nor U12259 (N_12259,N_11953,N_11597);
xor U12260 (N_12260,N_10101,N_10211);
and U12261 (N_12261,N_10231,N_10489);
nand U12262 (N_12262,N_11770,N_11709);
nor U12263 (N_12263,N_11583,N_11949);
or U12264 (N_12264,N_10664,N_10917);
nor U12265 (N_12265,N_10451,N_10088);
nor U12266 (N_12266,N_10268,N_11079);
nor U12267 (N_12267,N_11260,N_10109);
or U12268 (N_12268,N_10959,N_10121);
nand U12269 (N_12269,N_10680,N_10205);
and U12270 (N_12270,N_10925,N_10342);
or U12271 (N_12271,N_10841,N_10062);
xnor U12272 (N_12272,N_10596,N_10051);
nand U12273 (N_12273,N_11898,N_11519);
xor U12274 (N_12274,N_11988,N_10232);
and U12275 (N_12275,N_11993,N_11996);
nor U12276 (N_12276,N_11378,N_10756);
nand U12277 (N_12277,N_10817,N_11946);
and U12278 (N_12278,N_11263,N_10852);
nand U12279 (N_12279,N_10607,N_11835);
xor U12280 (N_12280,N_11047,N_11694);
nor U12281 (N_12281,N_11105,N_10281);
or U12282 (N_12282,N_11302,N_11406);
nand U12283 (N_12283,N_11214,N_10085);
nand U12284 (N_12284,N_11110,N_11045);
and U12285 (N_12285,N_10180,N_10771);
nand U12286 (N_12286,N_11695,N_10398);
or U12287 (N_12287,N_11657,N_11308);
or U12288 (N_12288,N_11827,N_11058);
nand U12289 (N_12289,N_10967,N_11578);
or U12290 (N_12290,N_11409,N_11377);
nor U12291 (N_12291,N_10512,N_10580);
nor U12292 (N_12292,N_11435,N_10350);
xor U12293 (N_12293,N_11586,N_11175);
or U12294 (N_12294,N_10091,N_11321);
xor U12295 (N_12295,N_11673,N_11491);
or U12296 (N_12296,N_11074,N_11774);
nand U12297 (N_12297,N_10482,N_11879);
and U12298 (N_12298,N_11444,N_10813);
nor U12299 (N_12299,N_11591,N_10376);
and U12300 (N_12300,N_11198,N_10990);
or U12301 (N_12301,N_10501,N_10665);
or U12302 (N_12302,N_10788,N_10156);
or U12303 (N_12303,N_10194,N_10486);
and U12304 (N_12304,N_11131,N_10643);
or U12305 (N_12305,N_10111,N_10470);
or U12306 (N_12306,N_11371,N_11493);
nand U12307 (N_12307,N_10761,N_10799);
nor U12308 (N_12308,N_11472,N_11705);
or U12309 (N_12309,N_10615,N_11174);
nor U12310 (N_12310,N_11489,N_10445);
nor U12311 (N_12311,N_10538,N_10657);
and U12312 (N_12312,N_10058,N_10192);
and U12313 (N_12313,N_10516,N_10892);
and U12314 (N_12314,N_10290,N_11750);
and U12315 (N_12315,N_10253,N_11380);
and U12316 (N_12316,N_10126,N_10259);
xnor U12317 (N_12317,N_10135,N_11108);
xor U12318 (N_12318,N_11221,N_10087);
and U12319 (N_12319,N_10292,N_11104);
xor U12320 (N_12320,N_11218,N_10807);
or U12321 (N_12321,N_10576,N_10874);
xnor U12322 (N_12322,N_10943,N_10975);
nand U12323 (N_12323,N_10394,N_11963);
nand U12324 (N_12324,N_10722,N_10080);
nand U12325 (N_12325,N_10276,N_11249);
nor U12326 (N_12326,N_10933,N_11508);
nor U12327 (N_12327,N_10185,N_11758);
nor U12328 (N_12328,N_11523,N_11057);
nand U12329 (N_12329,N_10026,N_11755);
and U12330 (N_12330,N_10688,N_10920);
nand U12331 (N_12331,N_11951,N_10112);
nand U12332 (N_12332,N_11039,N_11317);
or U12333 (N_12333,N_11925,N_11653);
nor U12334 (N_12334,N_10341,N_11162);
nor U12335 (N_12335,N_10528,N_11655);
xor U12336 (N_12336,N_11505,N_11554);
nand U12337 (N_12337,N_11041,N_11820);
nand U12338 (N_12338,N_11550,N_10711);
or U12339 (N_12339,N_11095,N_10682);
or U12340 (N_12340,N_11802,N_11078);
or U12341 (N_12341,N_10842,N_10776);
nor U12342 (N_12342,N_10851,N_11964);
nor U12343 (N_12343,N_10900,N_11844);
or U12344 (N_12344,N_10979,N_10951);
nor U12345 (N_12345,N_10002,N_10978);
nor U12346 (N_12346,N_11242,N_11651);
nand U12347 (N_12347,N_10380,N_10361);
and U12348 (N_12348,N_10221,N_10283);
or U12349 (N_12349,N_10494,N_11486);
xnor U12350 (N_12350,N_11368,N_10181);
nand U12351 (N_12351,N_11752,N_11087);
xnor U12352 (N_12352,N_10996,N_10793);
and U12353 (N_12353,N_10685,N_10197);
or U12354 (N_12354,N_11020,N_11316);
or U12355 (N_12355,N_11711,N_11029);
and U12356 (N_12356,N_10769,N_11134);
nor U12357 (N_12357,N_11359,N_11669);
and U12358 (N_12358,N_10055,N_10994);
and U12359 (N_12359,N_10454,N_11048);
or U12360 (N_12360,N_10698,N_10585);
or U12361 (N_12361,N_10833,N_11248);
xnor U12362 (N_12362,N_10335,N_11411);
xor U12363 (N_12363,N_10277,N_11834);
nand U12364 (N_12364,N_10525,N_11332);
nor U12365 (N_12365,N_10056,N_10926);
xor U12366 (N_12366,N_11969,N_11415);
nor U12367 (N_12367,N_11152,N_11203);
nand U12368 (N_12368,N_11116,N_11915);
nor U12369 (N_12369,N_11156,N_10714);
nor U12370 (N_12370,N_11971,N_11570);
and U12371 (N_12371,N_10459,N_10499);
xnor U12372 (N_12372,N_11387,N_11367);
or U12373 (N_12373,N_11751,N_10823);
nor U12374 (N_12374,N_10719,N_10530);
nand U12375 (N_12375,N_11463,N_10557);
and U12376 (N_12376,N_11481,N_10617);
and U12377 (N_12377,N_10319,N_10918);
or U12378 (N_12378,N_10064,N_11822);
xnor U12379 (N_12379,N_11256,N_11148);
nand U12380 (N_12380,N_11529,N_10594);
or U12381 (N_12381,N_10515,N_10307);
nand U12382 (N_12382,N_11683,N_11611);
nand U12383 (N_12383,N_10695,N_11111);
nor U12384 (N_12384,N_10730,N_11796);
nand U12385 (N_12385,N_10540,N_10948);
nor U12386 (N_12386,N_11264,N_11629);
nand U12387 (N_12387,N_10437,N_11838);
or U12388 (N_12388,N_11984,N_10608);
xnor U12389 (N_12389,N_10215,N_10008);
or U12390 (N_12390,N_10015,N_11272);
nor U12391 (N_12391,N_11080,N_11604);
nand U12392 (N_12392,N_10962,N_11932);
nor U12393 (N_12393,N_10791,N_11054);
and U12394 (N_12394,N_10621,N_11296);
nand U12395 (N_12395,N_10286,N_10707);
xnor U12396 (N_12396,N_11438,N_10902);
xnor U12397 (N_12397,N_10323,N_10821);
or U12398 (N_12398,N_11120,N_11781);
nand U12399 (N_12399,N_10298,N_10622);
xor U12400 (N_12400,N_10336,N_10774);
nand U12401 (N_12401,N_10261,N_10250);
nand U12402 (N_12402,N_11521,N_11672);
xor U12403 (N_12403,N_10020,N_11091);
nand U12404 (N_12404,N_10220,N_11506);
nor U12405 (N_12405,N_11598,N_10837);
nand U12406 (N_12406,N_10946,N_10847);
xor U12407 (N_12407,N_11829,N_10808);
or U12408 (N_12408,N_10419,N_10337);
xnor U12409 (N_12409,N_11343,N_10391);
nand U12410 (N_12410,N_11729,N_10144);
or U12411 (N_12411,N_10280,N_10303);
xnor U12412 (N_12412,N_10147,N_11662);
xor U12413 (N_12413,N_11128,N_11553);
and U12414 (N_12414,N_11348,N_10439);
xnor U12415 (N_12415,N_11153,N_11022);
nand U12416 (N_12416,N_10945,N_10717);
xor U12417 (N_12417,N_10003,N_10017);
nand U12418 (N_12418,N_10773,N_11903);
nor U12419 (N_12419,N_10216,N_11244);
xor U12420 (N_12420,N_11329,N_10740);
xnor U12421 (N_12421,N_10728,N_11560);
or U12422 (N_12422,N_10661,N_10034);
nor U12423 (N_12423,N_11081,N_11530);
nor U12424 (N_12424,N_10765,N_10537);
xor U12425 (N_12425,N_10923,N_10629);
nor U12426 (N_12426,N_11690,N_10519);
nor U12427 (N_12427,N_10060,N_11564);
xor U12428 (N_12428,N_11401,N_10937);
nand U12429 (N_12429,N_11061,N_10116);
nand U12430 (N_12430,N_11408,N_11223);
nor U12431 (N_12431,N_10870,N_10218);
xor U12432 (N_12432,N_11607,N_11010);
or U12433 (N_12433,N_10359,N_11171);
and U12434 (N_12434,N_11698,N_10263);
nand U12435 (N_12435,N_10090,N_11562);
or U12436 (N_12436,N_11906,N_10061);
nor U12437 (N_12437,N_11941,N_11809);
and U12438 (N_12438,N_10028,N_10119);
or U12439 (N_12439,N_10536,N_11337);
xor U12440 (N_12440,N_11138,N_11845);
or U12441 (N_12441,N_10481,N_10174);
or U12442 (N_12442,N_10227,N_11266);
nand U12443 (N_12443,N_11023,N_10324);
nand U12444 (N_12444,N_10522,N_11893);
nand U12445 (N_12445,N_11470,N_10299);
or U12446 (N_12446,N_10729,N_10961);
nor U12447 (N_12447,N_10539,N_10446);
or U12448 (N_12448,N_10160,N_11125);
nand U12449 (N_12449,N_10199,N_10011);
nor U12450 (N_12450,N_11816,N_11868);
or U12451 (N_12451,N_10110,N_10562);
and U12452 (N_12452,N_10041,N_11458);
nand U12453 (N_12453,N_10801,N_11697);
nor U12454 (N_12454,N_10831,N_10966);
and U12455 (N_12455,N_11713,N_11442);
xor U12456 (N_12456,N_10262,N_10927);
nor U12457 (N_12457,N_11973,N_11327);
nand U12458 (N_12458,N_11572,N_11660);
nor U12459 (N_12459,N_10754,N_10746);
or U12460 (N_12460,N_11402,N_10878);
or U12461 (N_12461,N_11986,N_10175);
and U12462 (N_12462,N_10634,N_11222);
xnor U12463 (N_12463,N_10903,N_10751);
and U12464 (N_12464,N_10830,N_10441);
or U12465 (N_12465,N_10880,N_10378);
nor U12466 (N_12466,N_10766,N_11012);
and U12467 (N_12467,N_11069,N_11848);
xor U12468 (N_12468,N_11756,N_10689);
or U12469 (N_12469,N_10931,N_10170);
xor U12470 (N_12470,N_11461,N_10347);
or U12471 (N_12471,N_11824,N_10374);
and U12472 (N_12472,N_11661,N_11547);
nand U12473 (N_12473,N_10010,N_10545);
or U12474 (N_12474,N_11117,N_10304);
and U12475 (N_12475,N_11182,N_11362);
and U12476 (N_12476,N_10915,N_10314);
or U12477 (N_12477,N_11930,N_11533);
and U12478 (N_12478,N_11028,N_10819);
and U12479 (N_12479,N_11679,N_11863);
nor U12480 (N_12480,N_11082,N_11236);
and U12481 (N_12481,N_10737,N_11682);
and U12482 (N_12482,N_11744,N_10289);
nand U12483 (N_12483,N_10700,N_11372);
xor U12484 (N_12484,N_10922,N_10403);
or U12485 (N_12485,N_10193,N_10693);
or U12486 (N_12486,N_11854,N_11688);
nand U12487 (N_12487,N_10094,N_11825);
xnor U12488 (N_12488,N_11567,N_11574);
nor U12489 (N_12489,N_10367,N_11687);
nor U12490 (N_12490,N_10368,N_11453);
nand U12491 (N_12491,N_10995,N_10243);
nor U12492 (N_12492,N_10428,N_10136);
nor U12493 (N_12493,N_10609,N_11188);
or U12494 (N_12494,N_10270,N_11191);
and U12495 (N_12495,N_10462,N_10527);
nor U12496 (N_12496,N_11836,N_10891);
nand U12497 (N_12497,N_10245,N_10673);
or U12498 (N_12498,N_10416,N_10627);
xnor U12499 (N_12499,N_10125,N_10589);
or U12500 (N_12500,N_10477,N_11479);
or U12501 (N_12501,N_11455,N_10679);
or U12502 (N_12502,N_10814,N_10138);
and U12503 (N_12503,N_11590,N_11612);
nand U12504 (N_12504,N_10704,N_11177);
or U12505 (N_12505,N_10692,N_10864);
or U12506 (N_12506,N_11990,N_11764);
xor U12507 (N_12507,N_10167,N_10388);
xor U12508 (N_12508,N_10804,N_11670);
xor U12509 (N_12509,N_11397,N_10616);
and U12510 (N_12510,N_10789,N_11107);
and U12511 (N_12511,N_10490,N_10955);
nand U12512 (N_12512,N_11727,N_11800);
and U12513 (N_12513,N_11085,N_11742);
nor U12514 (N_12514,N_11575,N_10716);
xor U12515 (N_12515,N_10397,N_11753);
and U12516 (N_12516,N_10025,N_10230);
and U12517 (N_12517,N_11905,N_11810);
and U12518 (N_12518,N_10178,N_10865);
nor U12519 (N_12519,N_10567,N_10768);
nand U12520 (N_12520,N_10384,N_11147);
or U12521 (N_12521,N_10273,N_10588);
nor U12522 (N_12522,N_10909,N_11165);
and U12523 (N_12523,N_10671,N_10418);
nor U12524 (N_12524,N_10929,N_11190);
and U12525 (N_12525,N_11013,N_10544);
xnor U12526 (N_12526,N_11924,N_10806);
and U12527 (N_12527,N_11121,N_11938);
nand U12528 (N_12528,N_11077,N_11636);
and U12529 (N_12529,N_11675,N_10255);
nand U12530 (N_12530,N_11538,N_11862);
nand U12531 (N_12531,N_11386,N_10881);
nor U12532 (N_12532,N_11421,N_11419);
or U12533 (N_12533,N_11939,N_11059);
nand U12534 (N_12534,N_10236,N_10137);
and U12535 (N_12535,N_10860,N_11342);
or U12536 (N_12536,N_10321,N_11677);
or U12537 (N_12537,N_10854,N_10675);
xnor U12538 (N_12538,N_11856,N_10882);
and U12539 (N_12539,N_11127,N_10572);
xnor U12540 (N_12540,N_11780,N_10741);
xnor U12541 (N_12541,N_11846,N_10952);
xor U12542 (N_12542,N_11920,N_10857);
xor U12543 (N_12543,N_11644,N_11309);
nor U12544 (N_12544,N_10274,N_11601);
and U12545 (N_12545,N_10140,N_11667);
nand U12546 (N_12546,N_11096,N_11904);
and U12547 (N_12547,N_11776,N_11385);
and U12548 (N_12548,N_11160,N_10991);
or U12549 (N_12549,N_11328,N_11228);
or U12550 (N_12550,N_10523,N_10031);
and U12551 (N_12551,N_11630,N_10942);
or U12552 (N_12552,N_11902,N_11842);
nand U12553 (N_12553,N_10726,N_10980);
or U12554 (N_12554,N_10389,N_11155);
nand U12555 (N_12555,N_11967,N_11639);
nor U12556 (N_12556,N_10947,N_10826);
xor U12557 (N_12557,N_11746,N_10452);
xnor U12558 (N_12558,N_11224,N_10606);
xnor U12559 (N_12559,N_11668,N_10063);
or U12560 (N_12560,N_10266,N_11584);
or U12561 (N_12561,N_10338,N_11484);
nand U12562 (N_12562,N_11295,N_10423);
or U12563 (N_12563,N_10422,N_11532);
and U12564 (N_12564,N_10897,N_10432);
xnor U12565 (N_12565,N_11417,N_11864);
xnor U12566 (N_12566,N_11173,N_10099);
nand U12567 (N_12567,N_10381,N_10047);
nand U12568 (N_12568,N_10310,N_10758);
xnor U12569 (N_12569,N_11889,N_11625);
nand U12570 (N_12570,N_11974,N_10113);
or U12571 (N_12571,N_10738,N_11715);
nor U12572 (N_12572,N_10427,N_10710);
nand U12573 (N_12573,N_11494,N_10625);
nand U12574 (N_12574,N_10131,N_11882);
nand U12575 (N_12575,N_11771,N_11977);
and U12576 (N_12576,N_11288,N_10039);
nor U12577 (N_12577,N_10763,N_11875);
xnor U12578 (N_12578,N_10460,N_10311);
xnor U12579 (N_12579,N_10667,N_11420);
nand U12580 (N_12580,N_11418,N_11795);
or U12581 (N_12581,N_11541,N_10440);
nand U12582 (N_12582,N_10182,N_11360);
nand U12583 (N_12583,N_10561,N_10556);
nand U12584 (N_12584,N_11867,N_11179);
xnor U12585 (N_12585,N_10655,N_11126);
nand U12586 (N_12586,N_11642,N_10014);
nand U12587 (N_12587,N_11496,N_11021);
or U12588 (N_12588,N_11592,N_10697);
nand U12589 (N_12589,N_11281,N_10360);
or U12590 (N_12590,N_10293,N_11436);
xor U12591 (N_12591,N_10200,N_11571);
xnor U12592 (N_12592,N_11350,N_10456);
nor U12593 (N_12593,N_11960,N_10053);
xor U12594 (N_12594,N_11158,N_10598);
nor U12595 (N_12595,N_11253,N_10772);
nand U12596 (N_12596,N_10306,N_11551);
nand U12597 (N_12597,N_10322,N_10214);
xnor U12598 (N_12598,N_11181,N_11535);
nor U12599 (N_12599,N_11596,N_11664);
xnor U12600 (N_12600,N_10644,N_10172);
xor U12601 (N_12601,N_10646,N_11492);
nor U12602 (N_12602,N_11433,N_10320);
nand U12603 (N_12603,N_10154,N_11030);
or U12604 (N_12604,N_11154,N_10889);
or U12605 (N_12605,N_11305,N_11804);
nor U12606 (N_12606,N_10022,N_11589);
or U12607 (N_12607,N_11888,N_11071);
nor U12608 (N_12608,N_10412,N_11961);
nor U12609 (N_12609,N_11404,N_11416);
xnor U12610 (N_12610,N_11916,N_10825);
xnor U12611 (N_12611,N_11300,N_11422);
nor U12612 (N_12612,N_10353,N_10436);
and U12613 (N_12613,N_10004,N_11994);
or U12614 (N_12614,N_11759,N_11640);
or U12615 (N_12615,N_11106,N_11313);
nor U12616 (N_12616,N_11566,N_10848);
xor U12617 (N_12617,N_11003,N_11255);
and U12618 (N_12618,N_10166,N_11251);
xor U12619 (N_12619,N_10649,N_11927);
and U12620 (N_12620,N_11837,N_11793);
xnor U12621 (N_12621,N_10599,N_11122);
and U12622 (N_12622,N_10668,N_10313);
nand U12623 (N_12623,N_11334,N_11220);
nor U12624 (N_12624,N_10884,N_11819);
nor U12625 (N_12625,N_11617,N_11766);
and U12626 (N_12626,N_10753,N_11754);
or U12627 (N_12627,N_11680,N_11928);
xor U12628 (N_12628,N_11037,N_10654);
nor U12629 (N_12629,N_11881,N_11016);
and U12630 (N_12630,N_10581,N_10420);
or U12631 (N_12631,N_10278,N_11090);
and U12632 (N_12632,N_10958,N_10853);
nor U12633 (N_12633,N_11602,N_11998);
xor U12634 (N_12634,N_11163,N_10349);
nor U12635 (N_12635,N_11579,N_10357);
and U12636 (N_12636,N_10551,N_10301);
nand U12637 (N_12637,N_11783,N_11462);
nor U12638 (N_12638,N_10744,N_10071);
xor U12639 (N_12639,N_10223,N_11852);
xor U12640 (N_12640,N_11318,N_10176);
and U12641 (N_12641,N_11374,N_11811);
xor U12642 (N_12642,N_10812,N_10308);
and U12643 (N_12643,N_10153,N_10899);
xnor U12644 (N_12644,N_10198,N_11789);
nor U12645 (N_12645,N_10203,N_11454);
nand U12646 (N_12646,N_10410,N_10339);
or U12647 (N_12647,N_11982,N_10709);
nor U12648 (N_12648,N_11119,N_10114);
nand U12649 (N_12649,N_10696,N_11790);
or U12650 (N_12650,N_10507,N_11637);
nand U12651 (N_12651,N_10001,N_10565);
xnor U12652 (N_12652,N_10663,N_10602);
and U12653 (N_12653,N_10188,N_10213);
nor U12654 (N_12654,N_10059,N_10288);
or U12655 (N_12655,N_11763,N_11363);
nor U12656 (N_12656,N_11024,N_10872);
nor U12657 (N_12657,N_11624,N_11649);
nand U12658 (N_12658,N_11068,N_11025);
nand U12659 (N_12659,N_11209,N_11724);
xor U12660 (N_12660,N_10186,N_11060);
xor U12661 (N_12661,N_10387,N_10246);
and U12662 (N_12662,N_11423,N_10632);
nand U12663 (N_12663,N_11083,N_10219);
xor U12664 (N_12664,N_10976,N_10736);
or U12665 (N_12665,N_11730,N_10780);
nor U12666 (N_12666,N_11931,N_11043);
nor U12667 (N_12667,N_10977,N_10844);
and U12668 (N_12668,N_11921,N_11544);
or U12669 (N_12669,N_11923,N_10706);
nor U12670 (N_12670,N_10510,N_10256);
nand U12671 (N_12671,N_10894,N_11942);
or U12672 (N_12672,N_11376,N_11606);
nor U12673 (N_12673,N_10351,N_11620);
nor U12674 (N_12674,N_11545,N_11046);
xnor U12675 (N_12675,N_10721,N_10601);
nor U12676 (N_12676,N_11784,N_10325);
and U12677 (N_12677,N_10168,N_11684);
and U12678 (N_12678,N_10838,N_10724);
and U12679 (N_12679,N_11522,N_11384);
xnor U12680 (N_12680,N_11947,N_10752);
nor U12681 (N_12681,N_11459,N_11347);
and U12682 (N_12682,N_10066,N_10939);
or U12683 (N_12683,N_10792,N_10905);
nand U12684 (N_12684,N_11167,N_10586);
or U12685 (N_12685,N_11565,N_11259);
and U12686 (N_12686,N_10009,N_10827);
xor U12687 (N_12687,N_10406,N_10797);
or U12688 (N_12688,N_11537,N_10040);
nor U12689 (N_12689,N_10981,N_11897);
and U12690 (N_12690,N_10480,N_10265);
xor U12691 (N_12691,N_10152,N_10784);
nor U12692 (N_12692,N_11443,N_10108);
nand U12693 (N_12693,N_11278,N_11885);
or U12694 (N_12694,N_10508,N_11217);
nor U12695 (N_12695,N_11027,N_11103);
nand U12696 (N_12696,N_10725,N_10201);
nand U12697 (N_12697,N_10563,N_11216);
and U12698 (N_12698,N_10972,N_10364);
nor U12699 (N_12699,N_11765,N_10098);
or U12700 (N_12700,N_10505,N_11388);
nor U12701 (N_12701,N_11487,N_10513);
and U12702 (N_12702,N_11428,N_11146);
and U12703 (N_12703,N_11270,N_10569);
nor U12704 (N_12704,N_10169,N_11113);
xnor U12705 (N_12705,N_10237,N_11934);
xor U12706 (N_12706,N_11600,N_10913);
nor U12707 (N_12707,N_10595,N_11678);
nor U12708 (N_12708,N_11324,N_10983);
and U12709 (N_12709,N_10096,N_10885);
nand U12710 (N_12710,N_11954,N_11170);
nor U12711 (N_12711,N_11891,N_11451);
nand U12712 (N_12712,N_11072,N_11036);
xnor U12713 (N_12713,N_11717,N_11995);
xnor U12714 (N_12714,N_11851,N_11685);
or U12715 (N_12715,N_10546,N_11734);
xor U12716 (N_12716,N_11341,N_10444);
xnor U12717 (N_12717,N_10438,N_10651);
xor U12718 (N_12718,N_10960,N_10824);
nor U12719 (N_12719,N_10485,N_10309);
nor U12720 (N_12720,N_11424,N_11084);
and U12721 (N_12721,N_11608,N_10970);
nor U12722 (N_12722,N_11722,N_11509);
and U12723 (N_12723,N_11681,N_10777);
nand U12724 (N_12724,N_11635,N_10086);
nand U12725 (N_12725,N_11065,N_11647);
nor U12726 (N_12726,N_10564,N_10233);
and U12727 (N_12727,N_10795,N_10998);
nand U12728 (N_12728,N_11511,N_11002);
nor U12729 (N_12729,N_10370,N_11129);
nor U12730 (N_12730,N_11073,N_10620);
and U12731 (N_12731,N_10333,N_10054);
nand U12732 (N_12732,N_11831,N_11011);
xor U12733 (N_12733,N_10612,N_11294);
xor U12734 (N_12734,N_11495,N_11277);
or U12735 (N_12735,N_11830,N_11089);
and U12736 (N_12736,N_10782,N_11760);
nand U12737 (N_12737,N_10989,N_10835);
xnor U12738 (N_12738,N_11749,N_10778);
or U12739 (N_12739,N_11124,N_11513);
or U12740 (N_12740,N_10701,N_11460);
or U12741 (N_12741,N_11981,N_10450);
or U12742 (N_12742,N_10447,N_11728);
xnor U12743 (N_12743,N_11208,N_11853);
nor U12744 (N_12744,N_10150,N_11390);
nand U12745 (N_12745,N_10414,N_11534);
nand U12746 (N_12746,N_10345,N_10805);
or U12747 (N_12747,N_11817,N_11157);
xor U12748 (N_12748,N_10779,N_11238);
xor U12749 (N_12749,N_11413,N_11861);
nand U12750 (N_12750,N_10127,N_10371);
or U12751 (N_12751,N_11895,N_10672);
or U12752 (N_12752,N_10057,N_11137);
xor U12753 (N_12753,N_10095,N_10458);
nand U12754 (N_12754,N_10718,N_10123);
or U12755 (N_12755,N_10734,N_11869);
nand U12756 (N_12756,N_11748,N_11659);
and U12757 (N_12757,N_10487,N_10217);
nand U12758 (N_12758,N_11032,N_11229);
or U12759 (N_12759,N_10343,N_10699);
and U12760 (N_12760,N_11212,N_10016);
or U12761 (N_12761,N_11908,N_11233);
and U12762 (N_12762,N_11737,N_11480);
or U12763 (N_12763,N_10354,N_10764);
nand U12764 (N_12764,N_11432,N_10358);
or U12765 (N_12765,N_11331,N_11704);
xnor U12766 (N_12766,N_10503,N_11322);
nor U12767 (N_12767,N_11919,N_10650);
xor U12768 (N_12768,N_11693,N_11871);
or U12769 (N_12769,N_10811,N_10653);
and U12770 (N_12770,N_11501,N_10834);
and U12771 (N_12771,N_11130,N_11349);
nor U12772 (N_12772,N_11557,N_10877);
xnor U12773 (N_12773,N_10238,N_10988);
and U12774 (N_12774,N_10558,N_11356);
or U12775 (N_12775,N_10102,N_11361);
xnor U12776 (N_12776,N_10334,N_11778);
nor U12777 (N_12777,N_10936,N_11714);
nand U12778 (N_12778,N_11500,N_11369);
and U12779 (N_12779,N_10749,N_11498);
nor U12780 (N_12780,N_10030,N_10727);
xor U12781 (N_12781,N_10940,N_10965);
nand U12782 (N_12782,N_11301,N_10187);
nor U12783 (N_12783,N_10798,N_10687);
xor U12784 (N_12784,N_11656,N_10896);
nand U12785 (N_12785,N_11204,N_10781);
nor U12786 (N_12786,N_11235,N_11840);
xor U12787 (N_12787,N_11166,N_10346);
xnor U12788 (N_12788,N_11292,N_10635);
nand U12789 (N_12789,N_11633,N_11149);
xor U12790 (N_12790,N_11252,N_11909);
nor U12791 (N_12791,N_10072,N_10822);
and U12792 (N_12792,N_11526,N_10641);
nand U12793 (N_12793,N_10448,N_11788);
nor U12794 (N_12794,N_11014,N_11033);
or U12795 (N_12795,N_10628,N_10074);
xnor U12796 (N_12796,N_11847,N_10465);
nand U12797 (N_12797,N_11808,N_10639);
and U12798 (N_12798,N_11826,N_11040);
nand U12799 (N_12799,N_10520,N_11365);
and U12800 (N_12800,N_10365,N_10431);
and U12801 (N_12801,N_11109,N_10495);
xnor U12802 (N_12802,N_11434,N_11716);
nand U12803 (N_12803,N_11064,N_10757);
nor U12804 (N_12804,N_10866,N_10742);
nand U12805 (N_12805,N_11412,N_10161);
nor U12806 (N_12806,N_11676,N_11273);
or U12807 (N_12807,N_10146,N_10257);
nor U12808 (N_12808,N_11603,N_11877);
nand U12809 (N_12809,N_11587,N_10404);
xnor U12810 (N_12810,N_11007,N_10382);
xnor U12811 (N_12811,N_11136,N_11142);
or U12812 (N_12812,N_10229,N_11745);
nor U12813 (N_12813,N_11671,N_10362);
or U12814 (N_12814,N_11552,N_10426);
nor U12815 (N_12815,N_11333,N_11213);
nor U12816 (N_12816,N_11665,N_10985);
nor U12817 (N_12817,N_10574,N_11720);
xor U12818 (N_12818,N_11150,N_10856);
or U12819 (N_12819,N_11017,N_11956);
nand U12820 (N_12820,N_11180,N_10845);
nand U12821 (N_12821,N_11610,N_11118);
nand U12822 (N_12822,N_10202,N_10443);
nand U12823 (N_12823,N_10312,N_10139);
and U12824 (N_12824,N_11818,N_10275);
and U12825 (N_12825,N_11762,N_11987);
xnor U12826 (N_12826,N_10787,N_10294);
and U12827 (N_12827,N_10993,N_11364);
or U12828 (N_12828,N_11241,N_10509);
nand U12829 (N_12829,N_11615,N_11843);
nor U12830 (N_12830,N_11782,N_11666);
or U12831 (N_12831,N_11185,N_11141);
nor U12832 (N_12832,N_10549,N_10548);
or U12833 (N_12833,N_11201,N_10868);
or U12834 (N_12834,N_11283,N_11595);
nor U12835 (N_12835,N_10466,N_10888);
and U12836 (N_12836,N_10859,N_11972);
or U12837 (N_12837,N_11976,N_11210);
nor U12838 (N_12838,N_10532,N_10012);
xor U12839 (N_12839,N_10151,N_11747);
nand U12840 (N_12840,N_10999,N_11926);
nor U12841 (N_12841,N_10155,N_10433);
nand U12842 (N_12842,N_10775,N_10476);
nor U12843 (N_12843,N_11807,N_11965);
nor U12844 (N_12844,N_10429,N_10249);
nor U12845 (N_12845,N_11357,N_11922);
nand U12846 (N_12846,N_10483,N_10497);
and U12847 (N_12847,N_11555,N_11568);
nor U12848 (N_12848,N_10408,N_11102);
or U12849 (N_12849,N_10023,N_11884);
nor U12850 (N_12850,N_11866,N_11474);
or U12851 (N_12851,N_10790,N_10670);
nand U12852 (N_12852,N_11250,N_10674);
xnor U12853 (N_12853,N_11164,N_10731);
or U12854 (N_12854,N_11429,N_10603);
and U12855 (N_12855,N_11382,N_10425);
xnor U12856 (N_12856,N_10148,N_10584);
or U12857 (N_12857,N_10869,N_11968);
and U12858 (N_12858,N_11703,N_11469);
xor U12859 (N_12859,N_11282,N_11403);
and U12860 (N_12860,N_10986,N_10747);
nand U12861 (N_12861,N_11691,N_11991);
nand U12862 (N_12862,N_11306,N_11733);
xnor U12863 (N_12863,N_10770,N_11430);
and U12864 (N_12864,N_11499,N_10372);
nor U12865 (N_12865,N_11936,N_11468);
nand U12866 (N_12866,N_10492,N_10484);
or U12867 (N_12867,N_11290,N_11814);
nor U12868 (N_12868,N_10863,N_10117);
xnor U12869 (N_12869,N_11628,N_11467);
and U12870 (N_12870,N_10473,N_10893);
nand U12871 (N_12871,N_10904,N_11289);
nor U12872 (N_12872,N_11937,N_10912);
nand U12873 (N_12873,N_11326,N_11035);
nor U12874 (N_12874,N_10049,N_11026);
nand U12875 (N_12875,N_10457,N_11275);
nand U12876 (N_12876,N_10518,N_11813);
nor U12877 (N_12877,N_10332,N_11614);
and U12878 (N_12878,N_10363,N_10921);
or U12879 (N_12879,N_11815,N_11009);
or U12880 (N_12880,N_10043,N_10132);
and U12881 (N_12881,N_11707,N_10383);
or U12882 (N_12882,N_10626,N_11582);
nand U12883 (N_12883,N_11516,N_11274);
and U12884 (N_12884,N_11841,N_11262);
nor U12885 (N_12885,N_11911,N_10317);
nor U12886 (N_12886,N_11355,N_10149);
nor U12887 (N_12887,N_11955,N_11806);
or U12888 (N_12888,N_11726,N_10021);
nand U12889 (N_12889,N_11338,N_10284);
nor U12890 (N_12890,N_11389,N_10206);
and U12891 (N_12891,N_10984,N_10195);
xnor U12892 (N_12892,N_10118,N_11502);
and U12893 (N_12893,N_11464,N_11515);
nor U12894 (N_12894,N_11740,N_11062);
and U12895 (N_12895,N_11768,N_10613);
nand U12896 (N_12896,N_11563,N_11396);
nor U12897 (N_12897,N_11336,N_10282);
xor U12898 (N_12898,N_10941,N_10604);
and U12899 (N_12899,N_10442,N_10068);
and U12900 (N_12900,N_10794,N_10209);
or U12901 (N_12901,N_11958,N_11019);
nor U12902 (N_12902,N_11706,N_11199);
nor U12903 (N_12903,N_10133,N_11512);
nand U12904 (N_12904,N_10506,N_10162);
or U12905 (N_12905,N_10681,N_10285);
xor U12906 (N_12906,N_10593,N_10163);
nor U12907 (N_12907,N_10677,N_11985);
nand U12908 (N_12908,N_11485,N_11743);
xor U12909 (N_12909,N_10073,N_10631);
and U12910 (N_12910,N_11395,N_10107);
nand U12911 (N_12911,N_11959,N_10691);
and U12912 (N_12912,N_10647,N_11546);
nor U12913 (N_12913,N_10469,N_10244);
nor U12914 (N_12914,N_11883,N_11398);
nand U12915 (N_12915,N_10502,N_10810);
xor U12916 (N_12916,N_11731,N_10226);
xnor U12917 (N_12917,N_11787,N_11441);
nor U12918 (N_12918,N_11779,N_10297);
nor U12919 (N_12919,N_11320,N_11622);
nor U12920 (N_12920,N_10678,N_10735);
or U12921 (N_12921,N_11593,N_10258);
or U12922 (N_12922,N_10733,N_11738);
and U12923 (N_12923,N_10919,N_10611);
or U12924 (N_12924,N_11979,N_11507);
nand U12925 (N_12925,N_10225,N_11966);
and U12926 (N_12926,N_11194,N_11929);
and U12927 (N_12927,N_10908,N_11801);
or U12928 (N_12928,N_10115,N_11381);
and U12929 (N_12929,N_10968,N_11873);
nand U12930 (N_12930,N_11049,N_10786);
nand U12931 (N_12931,N_11325,N_10159);
nand U12932 (N_12932,N_10050,N_10196);
xor U12933 (N_12933,N_10543,N_11632);
and U12934 (N_12934,N_11293,N_10836);
or U12935 (N_12935,N_11476,N_10871);
or U12936 (N_12936,N_11901,N_10930);
and U12937 (N_12937,N_11899,N_11539);
nand U12938 (N_12938,N_10474,N_10802);
nor U12939 (N_12939,N_11168,N_10550);
nand U12940 (N_12940,N_11431,N_10302);
nand U12941 (N_12941,N_10142,N_10076);
and U12942 (N_12942,N_11786,N_10630);
xor U12943 (N_12943,N_11605,N_10065);
nand U12944 (N_12944,N_11870,N_11354);
and U12945 (N_12945,N_10796,N_10067);
and U12946 (N_12946,N_11346,N_10705);
or U12947 (N_12947,N_10399,N_10177);
nor U12948 (N_12948,N_10901,N_10421);
or U12949 (N_12949,N_10828,N_11311);
or U12950 (N_12950,N_10190,N_11536);
xnor U12951 (N_12951,N_11268,N_10592);
xor U12952 (N_12952,N_10120,N_10251);
nor U12953 (N_12953,N_10356,N_10974);
xnor U12954 (N_12954,N_10479,N_11935);
or U12955 (N_12955,N_11399,N_10949);
nand U12956 (N_12956,N_10640,N_11475);
nor U12957 (N_12957,N_11205,N_11528);
and U12958 (N_12958,N_10954,N_10924);
and U12959 (N_12959,N_11577,N_10739);
and U12960 (N_12960,N_10883,N_11900);
nand U12961 (N_12961,N_11230,N_11196);
and U12962 (N_12962,N_11832,N_11053);
and U12963 (N_12963,N_10373,N_10849);
nand U12964 (N_12964,N_10618,N_10568);
nor U12965 (N_12965,N_11286,N_10648);
nor U12966 (N_12966,N_11284,N_11646);
xor U12967 (N_12967,N_10660,N_11245);
and U12968 (N_12968,N_10652,N_11887);
nor U12969 (N_12969,N_11088,N_11559);
or U12970 (N_12970,N_11339,N_11525);
nor U12971 (N_12971,N_11383,N_10690);
nor U12972 (N_12972,N_11702,N_11169);
and U12973 (N_12973,N_10145,N_11910);
nand U12974 (N_12974,N_10932,N_11280);
nor U12975 (N_12975,N_11042,N_11634);
nand U12976 (N_12976,N_10013,N_11000);
nor U12977 (N_12977,N_10987,N_10377);
or U12978 (N_12978,N_11425,N_11193);
and U12979 (N_12979,N_11226,N_11243);
nor U12980 (N_12980,N_11794,N_11514);
nor U12981 (N_12981,N_10461,N_10582);
xnor U12982 (N_12982,N_11319,N_10938);
nand U12983 (N_12983,N_11135,N_11874);
nor U12984 (N_12984,N_11340,N_10964);
nor U12985 (N_12985,N_10035,N_10843);
nand U12986 (N_12986,N_10956,N_11375);
xor U12987 (N_12987,N_10184,N_11865);
and U12988 (N_12988,N_11450,N_10610);
nand U12989 (N_12989,N_11699,N_10417);
nor U12990 (N_12990,N_11133,N_11151);
xnor U12991 (N_12991,N_11183,N_10005);
nand U12992 (N_12992,N_11034,N_10591);
xnor U12993 (N_12993,N_10208,N_10271);
and U12994 (N_12994,N_11573,N_11323);
xor U12995 (N_12995,N_10666,N_11839);
nor U12996 (N_12996,N_10534,N_10820);
nor U12997 (N_12997,N_10898,N_10455);
or U12998 (N_12998,N_10033,N_11543);
xor U12999 (N_12999,N_10413,N_11075);
and U13000 (N_13000,N_11516,N_10043);
and U13001 (N_13001,N_10746,N_10498);
nand U13002 (N_13002,N_10801,N_10221);
nor U13003 (N_13003,N_10070,N_10821);
nand U13004 (N_13004,N_10083,N_11887);
or U13005 (N_13005,N_10287,N_11004);
nor U13006 (N_13006,N_10911,N_10053);
nand U13007 (N_13007,N_10793,N_11795);
nor U13008 (N_13008,N_11801,N_11862);
nand U13009 (N_13009,N_11330,N_11438);
nor U13010 (N_13010,N_10339,N_10267);
nor U13011 (N_13011,N_10107,N_10706);
xnor U13012 (N_13012,N_11253,N_10657);
nor U13013 (N_13013,N_11937,N_10475);
or U13014 (N_13014,N_10851,N_10340);
or U13015 (N_13015,N_10369,N_11255);
nor U13016 (N_13016,N_10666,N_11319);
nor U13017 (N_13017,N_10105,N_10659);
nand U13018 (N_13018,N_10592,N_10853);
nand U13019 (N_13019,N_10549,N_10952);
or U13020 (N_13020,N_11238,N_10479);
nand U13021 (N_13021,N_11872,N_10833);
nor U13022 (N_13022,N_11436,N_11874);
and U13023 (N_13023,N_11897,N_10698);
nand U13024 (N_13024,N_11603,N_11721);
xnor U13025 (N_13025,N_11594,N_10470);
xor U13026 (N_13026,N_10845,N_11568);
or U13027 (N_13027,N_10917,N_11302);
and U13028 (N_13028,N_11066,N_10668);
and U13029 (N_13029,N_10701,N_10508);
and U13030 (N_13030,N_11598,N_10140);
and U13031 (N_13031,N_11410,N_11344);
or U13032 (N_13032,N_10168,N_10906);
and U13033 (N_13033,N_10477,N_11508);
nand U13034 (N_13034,N_10794,N_10687);
nand U13035 (N_13035,N_10220,N_11372);
or U13036 (N_13036,N_10562,N_10143);
nor U13037 (N_13037,N_11092,N_11399);
or U13038 (N_13038,N_10109,N_11485);
nor U13039 (N_13039,N_10797,N_10756);
or U13040 (N_13040,N_11877,N_10633);
and U13041 (N_13041,N_10590,N_10401);
or U13042 (N_13042,N_10609,N_10940);
nor U13043 (N_13043,N_11966,N_11289);
and U13044 (N_13044,N_11661,N_11399);
and U13045 (N_13045,N_11933,N_11390);
and U13046 (N_13046,N_10091,N_11728);
or U13047 (N_13047,N_10379,N_10342);
xnor U13048 (N_13048,N_11540,N_11659);
nand U13049 (N_13049,N_10072,N_10657);
and U13050 (N_13050,N_11448,N_11166);
or U13051 (N_13051,N_10879,N_10351);
or U13052 (N_13052,N_10365,N_10750);
and U13053 (N_13053,N_10292,N_11221);
and U13054 (N_13054,N_11787,N_10922);
nor U13055 (N_13055,N_10850,N_11800);
and U13056 (N_13056,N_10586,N_11833);
xor U13057 (N_13057,N_11071,N_11494);
and U13058 (N_13058,N_11288,N_10020);
or U13059 (N_13059,N_11989,N_11891);
or U13060 (N_13060,N_10656,N_11248);
xor U13061 (N_13061,N_11125,N_10100);
xor U13062 (N_13062,N_11461,N_10538);
and U13063 (N_13063,N_11811,N_11956);
or U13064 (N_13064,N_10848,N_10750);
nand U13065 (N_13065,N_10481,N_11802);
or U13066 (N_13066,N_10626,N_10684);
or U13067 (N_13067,N_11999,N_11393);
nor U13068 (N_13068,N_10774,N_10334);
xnor U13069 (N_13069,N_11117,N_10887);
nand U13070 (N_13070,N_10926,N_10808);
and U13071 (N_13071,N_11302,N_11672);
nand U13072 (N_13072,N_10296,N_10320);
xnor U13073 (N_13073,N_11061,N_10587);
nor U13074 (N_13074,N_11754,N_10682);
nor U13075 (N_13075,N_11869,N_10493);
and U13076 (N_13076,N_11427,N_10880);
and U13077 (N_13077,N_11846,N_11663);
nand U13078 (N_13078,N_11257,N_10015);
nor U13079 (N_13079,N_10974,N_11670);
xor U13080 (N_13080,N_10979,N_10194);
nor U13081 (N_13081,N_10617,N_10942);
or U13082 (N_13082,N_11017,N_10310);
and U13083 (N_13083,N_11767,N_11097);
or U13084 (N_13084,N_11833,N_11600);
and U13085 (N_13085,N_10634,N_10621);
and U13086 (N_13086,N_11268,N_10203);
nor U13087 (N_13087,N_10745,N_10050);
nand U13088 (N_13088,N_10977,N_10204);
nand U13089 (N_13089,N_11954,N_10530);
or U13090 (N_13090,N_11899,N_10134);
xnor U13091 (N_13091,N_10140,N_11751);
and U13092 (N_13092,N_11644,N_10875);
nor U13093 (N_13093,N_11772,N_11673);
nand U13094 (N_13094,N_11495,N_10963);
nand U13095 (N_13095,N_11019,N_11028);
or U13096 (N_13096,N_10818,N_11349);
and U13097 (N_13097,N_10869,N_10348);
nand U13098 (N_13098,N_10915,N_10361);
xor U13099 (N_13099,N_10088,N_11308);
nand U13100 (N_13100,N_10875,N_10244);
and U13101 (N_13101,N_10502,N_11331);
nand U13102 (N_13102,N_10559,N_11505);
xnor U13103 (N_13103,N_11559,N_11701);
or U13104 (N_13104,N_11055,N_10486);
nand U13105 (N_13105,N_10190,N_11553);
or U13106 (N_13106,N_10820,N_10288);
and U13107 (N_13107,N_10161,N_10750);
and U13108 (N_13108,N_10392,N_11779);
and U13109 (N_13109,N_11429,N_10109);
xor U13110 (N_13110,N_11166,N_10733);
nand U13111 (N_13111,N_11789,N_10959);
xor U13112 (N_13112,N_11217,N_10921);
nor U13113 (N_13113,N_10857,N_11330);
or U13114 (N_13114,N_10448,N_11711);
or U13115 (N_13115,N_11871,N_11882);
nor U13116 (N_13116,N_10623,N_11774);
or U13117 (N_13117,N_10182,N_10639);
or U13118 (N_13118,N_11595,N_11478);
nand U13119 (N_13119,N_10692,N_11799);
nand U13120 (N_13120,N_10053,N_10045);
or U13121 (N_13121,N_11919,N_10798);
or U13122 (N_13122,N_11505,N_11279);
nand U13123 (N_13123,N_11055,N_11962);
nand U13124 (N_13124,N_11131,N_10356);
nand U13125 (N_13125,N_10812,N_11972);
nand U13126 (N_13126,N_11356,N_11191);
nand U13127 (N_13127,N_10385,N_10082);
nand U13128 (N_13128,N_10100,N_10310);
or U13129 (N_13129,N_11774,N_11582);
nor U13130 (N_13130,N_10138,N_10252);
and U13131 (N_13131,N_11214,N_10429);
nand U13132 (N_13132,N_11253,N_10911);
nand U13133 (N_13133,N_10285,N_10192);
nand U13134 (N_13134,N_10661,N_10196);
nand U13135 (N_13135,N_11821,N_10691);
nand U13136 (N_13136,N_11799,N_10644);
nand U13137 (N_13137,N_10993,N_11528);
and U13138 (N_13138,N_10936,N_11676);
or U13139 (N_13139,N_10157,N_11766);
nor U13140 (N_13140,N_10847,N_11169);
nor U13141 (N_13141,N_11980,N_11136);
or U13142 (N_13142,N_10731,N_10141);
nand U13143 (N_13143,N_10102,N_11396);
or U13144 (N_13144,N_10282,N_10645);
nand U13145 (N_13145,N_10673,N_11663);
xnor U13146 (N_13146,N_11702,N_10596);
nand U13147 (N_13147,N_11915,N_10853);
or U13148 (N_13148,N_11631,N_11812);
xor U13149 (N_13149,N_11552,N_10882);
or U13150 (N_13150,N_10846,N_10086);
xnor U13151 (N_13151,N_11288,N_10716);
or U13152 (N_13152,N_11118,N_11657);
nand U13153 (N_13153,N_11945,N_10326);
xnor U13154 (N_13154,N_10848,N_10691);
nand U13155 (N_13155,N_11864,N_10036);
nor U13156 (N_13156,N_10152,N_11224);
xnor U13157 (N_13157,N_10542,N_11540);
xor U13158 (N_13158,N_11908,N_10418);
nand U13159 (N_13159,N_11079,N_11185);
and U13160 (N_13160,N_11190,N_11823);
nor U13161 (N_13161,N_10907,N_11494);
and U13162 (N_13162,N_10606,N_10720);
and U13163 (N_13163,N_11963,N_11479);
nor U13164 (N_13164,N_11782,N_10746);
xor U13165 (N_13165,N_10100,N_11862);
nand U13166 (N_13166,N_11582,N_11016);
and U13167 (N_13167,N_11195,N_11923);
nor U13168 (N_13168,N_11566,N_10672);
xnor U13169 (N_13169,N_11643,N_11347);
or U13170 (N_13170,N_10466,N_10485);
nor U13171 (N_13171,N_10567,N_11261);
xnor U13172 (N_13172,N_10967,N_10557);
or U13173 (N_13173,N_11883,N_11388);
xor U13174 (N_13174,N_10286,N_11457);
or U13175 (N_13175,N_10670,N_11701);
nor U13176 (N_13176,N_11978,N_10928);
nor U13177 (N_13177,N_10409,N_10029);
nand U13178 (N_13178,N_11778,N_11609);
nand U13179 (N_13179,N_10150,N_10088);
and U13180 (N_13180,N_11355,N_11966);
nand U13181 (N_13181,N_11405,N_10864);
and U13182 (N_13182,N_11901,N_11699);
nor U13183 (N_13183,N_10701,N_11234);
nand U13184 (N_13184,N_10695,N_10446);
or U13185 (N_13185,N_11871,N_11346);
or U13186 (N_13186,N_11586,N_11730);
xnor U13187 (N_13187,N_10019,N_10743);
nor U13188 (N_13188,N_11817,N_10276);
and U13189 (N_13189,N_10395,N_11894);
and U13190 (N_13190,N_10805,N_10381);
xor U13191 (N_13191,N_10423,N_10534);
or U13192 (N_13192,N_10585,N_10304);
xnor U13193 (N_13193,N_10299,N_10568);
and U13194 (N_13194,N_10896,N_11634);
nor U13195 (N_13195,N_10133,N_11601);
and U13196 (N_13196,N_10507,N_10108);
xor U13197 (N_13197,N_11821,N_10784);
xor U13198 (N_13198,N_11630,N_11367);
nand U13199 (N_13199,N_10274,N_10682);
and U13200 (N_13200,N_11998,N_11044);
xor U13201 (N_13201,N_11532,N_11568);
nand U13202 (N_13202,N_11529,N_11956);
xor U13203 (N_13203,N_11841,N_10028);
and U13204 (N_13204,N_11137,N_11257);
xnor U13205 (N_13205,N_10519,N_10916);
and U13206 (N_13206,N_10069,N_10050);
nor U13207 (N_13207,N_10521,N_10158);
nor U13208 (N_13208,N_11932,N_10624);
and U13209 (N_13209,N_10872,N_10601);
xnor U13210 (N_13210,N_11495,N_10377);
nand U13211 (N_13211,N_11837,N_11354);
or U13212 (N_13212,N_10280,N_11178);
and U13213 (N_13213,N_10929,N_10621);
or U13214 (N_13214,N_10993,N_10287);
nor U13215 (N_13215,N_10177,N_10247);
nand U13216 (N_13216,N_10274,N_11927);
or U13217 (N_13217,N_10840,N_10253);
nor U13218 (N_13218,N_10944,N_11216);
xor U13219 (N_13219,N_10204,N_10433);
nand U13220 (N_13220,N_11343,N_10808);
nor U13221 (N_13221,N_11828,N_10991);
and U13222 (N_13222,N_11137,N_11314);
or U13223 (N_13223,N_10200,N_10058);
xor U13224 (N_13224,N_11660,N_10246);
xnor U13225 (N_13225,N_11537,N_11000);
nand U13226 (N_13226,N_11781,N_11501);
nor U13227 (N_13227,N_10797,N_10783);
nand U13228 (N_13228,N_10739,N_10548);
and U13229 (N_13229,N_10601,N_10931);
or U13230 (N_13230,N_11141,N_11878);
and U13231 (N_13231,N_11729,N_11568);
xnor U13232 (N_13232,N_10724,N_11310);
and U13233 (N_13233,N_10358,N_10801);
or U13234 (N_13234,N_10499,N_11040);
xor U13235 (N_13235,N_10917,N_11488);
xor U13236 (N_13236,N_11442,N_10520);
and U13237 (N_13237,N_11709,N_11455);
or U13238 (N_13238,N_10549,N_10786);
or U13239 (N_13239,N_11217,N_10946);
xnor U13240 (N_13240,N_11382,N_10435);
nor U13241 (N_13241,N_10335,N_10372);
xnor U13242 (N_13242,N_10313,N_11879);
xnor U13243 (N_13243,N_10249,N_10841);
nor U13244 (N_13244,N_10333,N_10218);
or U13245 (N_13245,N_11224,N_11726);
nor U13246 (N_13246,N_11825,N_11745);
and U13247 (N_13247,N_10367,N_10565);
nor U13248 (N_13248,N_10036,N_10456);
nand U13249 (N_13249,N_10495,N_11365);
nor U13250 (N_13250,N_11257,N_10401);
xnor U13251 (N_13251,N_11249,N_10024);
nand U13252 (N_13252,N_11380,N_11916);
nor U13253 (N_13253,N_10830,N_11467);
nor U13254 (N_13254,N_11790,N_11418);
xor U13255 (N_13255,N_11695,N_10466);
nor U13256 (N_13256,N_10010,N_11659);
or U13257 (N_13257,N_11227,N_11867);
xor U13258 (N_13258,N_10452,N_11341);
nand U13259 (N_13259,N_11330,N_10908);
nor U13260 (N_13260,N_11759,N_10376);
nor U13261 (N_13261,N_11618,N_10637);
nor U13262 (N_13262,N_11610,N_11437);
nor U13263 (N_13263,N_11812,N_11541);
or U13264 (N_13264,N_11486,N_10804);
nand U13265 (N_13265,N_10289,N_11063);
xnor U13266 (N_13266,N_11782,N_11952);
xor U13267 (N_13267,N_11817,N_10448);
or U13268 (N_13268,N_10849,N_11142);
xor U13269 (N_13269,N_10421,N_10663);
nand U13270 (N_13270,N_11620,N_10234);
or U13271 (N_13271,N_11762,N_10815);
or U13272 (N_13272,N_10257,N_10217);
and U13273 (N_13273,N_11177,N_10028);
and U13274 (N_13274,N_10280,N_11452);
nor U13275 (N_13275,N_10699,N_11399);
and U13276 (N_13276,N_10013,N_10706);
nand U13277 (N_13277,N_10328,N_10213);
and U13278 (N_13278,N_10921,N_11733);
nor U13279 (N_13279,N_11678,N_11101);
nand U13280 (N_13280,N_11903,N_10894);
nand U13281 (N_13281,N_10776,N_11462);
nor U13282 (N_13282,N_10209,N_10256);
nand U13283 (N_13283,N_11765,N_11240);
nor U13284 (N_13284,N_11265,N_11649);
nor U13285 (N_13285,N_11962,N_10231);
or U13286 (N_13286,N_11104,N_10806);
xnor U13287 (N_13287,N_11085,N_10520);
and U13288 (N_13288,N_11628,N_11609);
nand U13289 (N_13289,N_11891,N_11276);
or U13290 (N_13290,N_10372,N_11638);
nand U13291 (N_13291,N_10938,N_10032);
and U13292 (N_13292,N_10028,N_10615);
nand U13293 (N_13293,N_11469,N_11530);
nor U13294 (N_13294,N_10491,N_11930);
nand U13295 (N_13295,N_11935,N_10174);
nand U13296 (N_13296,N_10272,N_11351);
xor U13297 (N_13297,N_10788,N_11250);
and U13298 (N_13298,N_11087,N_10494);
nand U13299 (N_13299,N_10894,N_10743);
and U13300 (N_13300,N_10299,N_10326);
nand U13301 (N_13301,N_11815,N_11616);
and U13302 (N_13302,N_11571,N_10505);
xor U13303 (N_13303,N_11451,N_10183);
or U13304 (N_13304,N_11410,N_11436);
nor U13305 (N_13305,N_10098,N_10995);
xor U13306 (N_13306,N_11018,N_11997);
or U13307 (N_13307,N_11896,N_10221);
xnor U13308 (N_13308,N_11677,N_11167);
xnor U13309 (N_13309,N_10710,N_11751);
and U13310 (N_13310,N_11924,N_11284);
or U13311 (N_13311,N_11961,N_11244);
and U13312 (N_13312,N_11962,N_10738);
nor U13313 (N_13313,N_11647,N_11657);
nor U13314 (N_13314,N_10299,N_11744);
nand U13315 (N_13315,N_10226,N_10889);
nor U13316 (N_13316,N_10813,N_11169);
or U13317 (N_13317,N_11131,N_11157);
or U13318 (N_13318,N_11417,N_10451);
nand U13319 (N_13319,N_11250,N_11355);
nor U13320 (N_13320,N_11706,N_11827);
or U13321 (N_13321,N_10450,N_10879);
or U13322 (N_13322,N_10338,N_10180);
and U13323 (N_13323,N_11918,N_10862);
xnor U13324 (N_13324,N_11861,N_10745);
nor U13325 (N_13325,N_10867,N_11938);
xor U13326 (N_13326,N_11274,N_10043);
and U13327 (N_13327,N_10749,N_10118);
and U13328 (N_13328,N_11380,N_10929);
nand U13329 (N_13329,N_11766,N_11889);
or U13330 (N_13330,N_11022,N_11150);
nor U13331 (N_13331,N_11920,N_10291);
nor U13332 (N_13332,N_10490,N_10924);
or U13333 (N_13333,N_10894,N_10416);
and U13334 (N_13334,N_10542,N_11608);
xor U13335 (N_13335,N_11575,N_11926);
nand U13336 (N_13336,N_10049,N_10091);
or U13337 (N_13337,N_10062,N_10906);
and U13338 (N_13338,N_10528,N_11009);
xnor U13339 (N_13339,N_11091,N_10797);
and U13340 (N_13340,N_11868,N_10794);
xor U13341 (N_13341,N_10026,N_11172);
nor U13342 (N_13342,N_10506,N_10293);
and U13343 (N_13343,N_11820,N_11476);
and U13344 (N_13344,N_11044,N_11368);
xnor U13345 (N_13345,N_10388,N_10946);
nor U13346 (N_13346,N_10618,N_10207);
xnor U13347 (N_13347,N_10636,N_11592);
or U13348 (N_13348,N_10754,N_10413);
or U13349 (N_13349,N_10863,N_10321);
xnor U13350 (N_13350,N_10022,N_11016);
nor U13351 (N_13351,N_11864,N_10170);
nor U13352 (N_13352,N_10519,N_11694);
and U13353 (N_13353,N_10603,N_11444);
or U13354 (N_13354,N_10019,N_10939);
and U13355 (N_13355,N_10383,N_10905);
nand U13356 (N_13356,N_11804,N_10688);
xor U13357 (N_13357,N_10320,N_10017);
and U13358 (N_13358,N_10842,N_11043);
xor U13359 (N_13359,N_11154,N_11669);
nand U13360 (N_13360,N_10670,N_10602);
or U13361 (N_13361,N_11360,N_10769);
xnor U13362 (N_13362,N_10118,N_11964);
nor U13363 (N_13363,N_11004,N_11321);
nand U13364 (N_13364,N_10497,N_11656);
nor U13365 (N_13365,N_10764,N_11136);
xor U13366 (N_13366,N_10890,N_11982);
nor U13367 (N_13367,N_10749,N_10160);
and U13368 (N_13368,N_10062,N_11483);
xor U13369 (N_13369,N_10026,N_11425);
and U13370 (N_13370,N_11805,N_11158);
xnor U13371 (N_13371,N_10414,N_11891);
xnor U13372 (N_13372,N_11605,N_10795);
nor U13373 (N_13373,N_11638,N_10534);
and U13374 (N_13374,N_10475,N_11710);
or U13375 (N_13375,N_11900,N_10328);
nand U13376 (N_13376,N_11048,N_10519);
xor U13377 (N_13377,N_11415,N_11983);
or U13378 (N_13378,N_10281,N_11893);
and U13379 (N_13379,N_11892,N_11676);
nand U13380 (N_13380,N_10629,N_11588);
or U13381 (N_13381,N_10679,N_11924);
nor U13382 (N_13382,N_11740,N_11423);
and U13383 (N_13383,N_11542,N_11962);
nand U13384 (N_13384,N_10255,N_11745);
and U13385 (N_13385,N_11186,N_10732);
nand U13386 (N_13386,N_11877,N_10093);
nand U13387 (N_13387,N_10798,N_11204);
and U13388 (N_13388,N_10604,N_11149);
nand U13389 (N_13389,N_10218,N_11661);
xor U13390 (N_13390,N_11168,N_10855);
nand U13391 (N_13391,N_11069,N_11890);
nor U13392 (N_13392,N_10192,N_10639);
xor U13393 (N_13393,N_10854,N_11912);
xnor U13394 (N_13394,N_10505,N_10584);
and U13395 (N_13395,N_11771,N_10800);
xor U13396 (N_13396,N_10237,N_11656);
nor U13397 (N_13397,N_11967,N_11386);
xnor U13398 (N_13398,N_11448,N_11018);
and U13399 (N_13399,N_10894,N_11641);
nor U13400 (N_13400,N_10386,N_11986);
and U13401 (N_13401,N_11995,N_10423);
xor U13402 (N_13402,N_11998,N_11930);
and U13403 (N_13403,N_11460,N_10940);
nor U13404 (N_13404,N_11536,N_10820);
nor U13405 (N_13405,N_11450,N_10196);
xnor U13406 (N_13406,N_11898,N_10590);
nand U13407 (N_13407,N_10324,N_10128);
nor U13408 (N_13408,N_11746,N_10230);
xor U13409 (N_13409,N_10778,N_11582);
nor U13410 (N_13410,N_10469,N_11243);
and U13411 (N_13411,N_11812,N_10993);
xnor U13412 (N_13412,N_10883,N_10985);
or U13413 (N_13413,N_10237,N_10845);
xnor U13414 (N_13414,N_11226,N_10125);
and U13415 (N_13415,N_10038,N_11845);
or U13416 (N_13416,N_11169,N_11023);
or U13417 (N_13417,N_11443,N_11505);
and U13418 (N_13418,N_11306,N_11924);
and U13419 (N_13419,N_10850,N_11853);
nor U13420 (N_13420,N_10333,N_11477);
or U13421 (N_13421,N_11683,N_11293);
xor U13422 (N_13422,N_10367,N_10391);
xnor U13423 (N_13423,N_11873,N_11794);
xor U13424 (N_13424,N_10453,N_11841);
nand U13425 (N_13425,N_11687,N_10384);
xnor U13426 (N_13426,N_11847,N_11098);
nand U13427 (N_13427,N_10776,N_11973);
nor U13428 (N_13428,N_11567,N_10868);
nand U13429 (N_13429,N_11495,N_11595);
nand U13430 (N_13430,N_11208,N_10745);
and U13431 (N_13431,N_10155,N_10291);
nand U13432 (N_13432,N_10160,N_11972);
or U13433 (N_13433,N_10479,N_10005);
and U13434 (N_13434,N_11036,N_11503);
or U13435 (N_13435,N_10856,N_10649);
and U13436 (N_13436,N_11879,N_11973);
and U13437 (N_13437,N_11549,N_10067);
and U13438 (N_13438,N_10971,N_11606);
and U13439 (N_13439,N_10899,N_11378);
nor U13440 (N_13440,N_10619,N_11042);
and U13441 (N_13441,N_10816,N_10840);
and U13442 (N_13442,N_11571,N_11502);
and U13443 (N_13443,N_10536,N_11996);
nor U13444 (N_13444,N_11137,N_10991);
xnor U13445 (N_13445,N_11361,N_10057);
or U13446 (N_13446,N_10498,N_11618);
or U13447 (N_13447,N_11083,N_11433);
and U13448 (N_13448,N_10665,N_11989);
nand U13449 (N_13449,N_11179,N_10951);
xnor U13450 (N_13450,N_10705,N_11704);
xnor U13451 (N_13451,N_11147,N_11194);
or U13452 (N_13452,N_10407,N_11341);
and U13453 (N_13453,N_10831,N_11441);
and U13454 (N_13454,N_11966,N_10058);
nand U13455 (N_13455,N_10344,N_11337);
and U13456 (N_13456,N_10247,N_10994);
and U13457 (N_13457,N_11701,N_11631);
xor U13458 (N_13458,N_11241,N_10150);
nand U13459 (N_13459,N_11756,N_11181);
or U13460 (N_13460,N_11566,N_10216);
or U13461 (N_13461,N_10925,N_10169);
or U13462 (N_13462,N_11601,N_10829);
and U13463 (N_13463,N_11259,N_10246);
or U13464 (N_13464,N_10347,N_10934);
and U13465 (N_13465,N_11907,N_11111);
nor U13466 (N_13466,N_10361,N_11314);
or U13467 (N_13467,N_11566,N_10388);
or U13468 (N_13468,N_11356,N_10467);
nor U13469 (N_13469,N_11255,N_10452);
nor U13470 (N_13470,N_11534,N_11470);
or U13471 (N_13471,N_10599,N_11760);
or U13472 (N_13472,N_10009,N_10175);
or U13473 (N_13473,N_11247,N_11365);
and U13474 (N_13474,N_10533,N_10660);
nand U13475 (N_13475,N_10041,N_10378);
xnor U13476 (N_13476,N_10785,N_10991);
nor U13477 (N_13477,N_11291,N_11152);
or U13478 (N_13478,N_10879,N_11255);
xor U13479 (N_13479,N_10627,N_10955);
or U13480 (N_13480,N_10862,N_10114);
xnor U13481 (N_13481,N_11215,N_10223);
xor U13482 (N_13482,N_10917,N_10796);
nand U13483 (N_13483,N_10952,N_11106);
or U13484 (N_13484,N_10813,N_11736);
xnor U13485 (N_13485,N_10957,N_11764);
xnor U13486 (N_13486,N_11359,N_10803);
nor U13487 (N_13487,N_10275,N_10967);
or U13488 (N_13488,N_11158,N_10778);
xnor U13489 (N_13489,N_10937,N_10285);
or U13490 (N_13490,N_11946,N_10157);
xnor U13491 (N_13491,N_10912,N_10272);
and U13492 (N_13492,N_11623,N_11297);
or U13493 (N_13493,N_10227,N_10797);
nand U13494 (N_13494,N_11804,N_10860);
nand U13495 (N_13495,N_10854,N_11417);
or U13496 (N_13496,N_11861,N_11836);
xnor U13497 (N_13497,N_10247,N_10713);
xnor U13498 (N_13498,N_11666,N_10648);
nor U13499 (N_13499,N_11608,N_10546);
nor U13500 (N_13500,N_10980,N_10845);
or U13501 (N_13501,N_11741,N_10781);
nor U13502 (N_13502,N_11705,N_11897);
nor U13503 (N_13503,N_10488,N_10489);
or U13504 (N_13504,N_11203,N_11439);
or U13505 (N_13505,N_10626,N_10884);
and U13506 (N_13506,N_10744,N_11213);
or U13507 (N_13507,N_10518,N_11284);
or U13508 (N_13508,N_11605,N_10144);
xnor U13509 (N_13509,N_11000,N_11838);
or U13510 (N_13510,N_10290,N_11338);
xor U13511 (N_13511,N_11257,N_11926);
or U13512 (N_13512,N_10186,N_10878);
and U13513 (N_13513,N_10384,N_11681);
or U13514 (N_13514,N_11085,N_11688);
nand U13515 (N_13515,N_10329,N_10343);
nand U13516 (N_13516,N_11498,N_10966);
nor U13517 (N_13517,N_11809,N_11428);
nor U13518 (N_13518,N_11390,N_11599);
nand U13519 (N_13519,N_10581,N_10759);
or U13520 (N_13520,N_11559,N_10347);
xor U13521 (N_13521,N_10425,N_11148);
nand U13522 (N_13522,N_10737,N_10802);
nor U13523 (N_13523,N_10458,N_11198);
or U13524 (N_13524,N_10717,N_10598);
nor U13525 (N_13525,N_11618,N_10924);
nand U13526 (N_13526,N_11625,N_11332);
nor U13527 (N_13527,N_11152,N_10841);
xnor U13528 (N_13528,N_11463,N_10241);
nand U13529 (N_13529,N_10714,N_10971);
and U13530 (N_13530,N_11702,N_11433);
nand U13531 (N_13531,N_11628,N_11910);
nand U13532 (N_13532,N_10982,N_11532);
xor U13533 (N_13533,N_11841,N_11237);
nor U13534 (N_13534,N_11674,N_10512);
and U13535 (N_13535,N_11330,N_11843);
or U13536 (N_13536,N_10429,N_10683);
or U13537 (N_13537,N_10585,N_10715);
nor U13538 (N_13538,N_10380,N_11648);
xnor U13539 (N_13539,N_10088,N_10132);
and U13540 (N_13540,N_11545,N_11131);
or U13541 (N_13541,N_11100,N_11427);
nand U13542 (N_13542,N_11353,N_10126);
nor U13543 (N_13543,N_10918,N_10938);
nand U13544 (N_13544,N_10966,N_11289);
nor U13545 (N_13545,N_11025,N_10350);
nand U13546 (N_13546,N_10974,N_10731);
xor U13547 (N_13547,N_11985,N_11751);
and U13548 (N_13548,N_11876,N_11364);
and U13549 (N_13549,N_11857,N_10975);
and U13550 (N_13550,N_10501,N_10000);
xnor U13551 (N_13551,N_10056,N_10749);
nor U13552 (N_13552,N_11806,N_11072);
nor U13553 (N_13553,N_10079,N_10903);
nand U13554 (N_13554,N_10972,N_11603);
or U13555 (N_13555,N_10177,N_11199);
nand U13556 (N_13556,N_11247,N_10636);
or U13557 (N_13557,N_10190,N_11550);
and U13558 (N_13558,N_11556,N_10484);
nand U13559 (N_13559,N_11922,N_11608);
or U13560 (N_13560,N_11952,N_11634);
xor U13561 (N_13561,N_11803,N_10338);
xnor U13562 (N_13562,N_11338,N_10603);
xnor U13563 (N_13563,N_10749,N_11837);
nor U13564 (N_13564,N_10440,N_10477);
xor U13565 (N_13565,N_10976,N_11486);
nand U13566 (N_13566,N_11384,N_10246);
and U13567 (N_13567,N_11982,N_11390);
and U13568 (N_13568,N_10932,N_11900);
and U13569 (N_13569,N_10163,N_10212);
and U13570 (N_13570,N_11238,N_11832);
nor U13571 (N_13571,N_10525,N_10746);
nand U13572 (N_13572,N_10405,N_11456);
and U13573 (N_13573,N_11535,N_11932);
and U13574 (N_13574,N_10717,N_10649);
nand U13575 (N_13575,N_10703,N_10151);
or U13576 (N_13576,N_11740,N_11204);
xor U13577 (N_13577,N_11574,N_10616);
and U13578 (N_13578,N_10915,N_10577);
or U13579 (N_13579,N_10993,N_11534);
or U13580 (N_13580,N_10998,N_10777);
xnor U13581 (N_13581,N_10925,N_10328);
and U13582 (N_13582,N_10172,N_11732);
xor U13583 (N_13583,N_10509,N_11334);
xnor U13584 (N_13584,N_11346,N_11226);
nor U13585 (N_13585,N_10806,N_10910);
and U13586 (N_13586,N_10653,N_11370);
nor U13587 (N_13587,N_11951,N_10707);
nor U13588 (N_13588,N_11512,N_10644);
nor U13589 (N_13589,N_10262,N_11888);
or U13590 (N_13590,N_10691,N_10804);
xor U13591 (N_13591,N_11733,N_10160);
and U13592 (N_13592,N_11930,N_10060);
nand U13593 (N_13593,N_10656,N_11688);
nor U13594 (N_13594,N_11640,N_11969);
xor U13595 (N_13595,N_11944,N_10171);
nor U13596 (N_13596,N_10630,N_10131);
and U13597 (N_13597,N_10876,N_11790);
nor U13598 (N_13598,N_10382,N_11327);
nand U13599 (N_13599,N_10404,N_10396);
xor U13600 (N_13600,N_11633,N_11043);
or U13601 (N_13601,N_11841,N_11922);
and U13602 (N_13602,N_10015,N_11147);
or U13603 (N_13603,N_11966,N_11928);
and U13604 (N_13604,N_11995,N_11480);
nor U13605 (N_13605,N_10565,N_10704);
xor U13606 (N_13606,N_11916,N_11007);
nand U13607 (N_13607,N_10024,N_11583);
or U13608 (N_13608,N_11201,N_10661);
and U13609 (N_13609,N_11014,N_10173);
xor U13610 (N_13610,N_11578,N_10530);
and U13611 (N_13611,N_11049,N_10928);
xnor U13612 (N_13612,N_11840,N_11052);
nor U13613 (N_13613,N_11967,N_11365);
xor U13614 (N_13614,N_10550,N_10261);
nand U13615 (N_13615,N_11912,N_11531);
and U13616 (N_13616,N_11111,N_11855);
nand U13617 (N_13617,N_11989,N_10472);
nand U13618 (N_13618,N_11943,N_11637);
and U13619 (N_13619,N_10249,N_10088);
and U13620 (N_13620,N_10974,N_10523);
xnor U13621 (N_13621,N_10956,N_11882);
nor U13622 (N_13622,N_10144,N_10178);
nand U13623 (N_13623,N_10821,N_11341);
and U13624 (N_13624,N_11372,N_10598);
nor U13625 (N_13625,N_11939,N_10235);
xor U13626 (N_13626,N_10162,N_10656);
nand U13627 (N_13627,N_11380,N_11267);
xnor U13628 (N_13628,N_11841,N_11687);
nand U13629 (N_13629,N_10342,N_10238);
or U13630 (N_13630,N_10266,N_11556);
nor U13631 (N_13631,N_11142,N_10635);
or U13632 (N_13632,N_11755,N_11056);
or U13633 (N_13633,N_10045,N_10490);
xnor U13634 (N_13634,N_11457,N_10081);
and U13635 (N_13635,N_11172,N_10148);
nand U13636 (N_13636,N_10405,N_10337);
or U13637 (N_13637,N_11689,N_10423);
nand U13638 (N_13638,N_11622,N_10508);
xnor U13639 (N_13639,N_10568,N_10714);
nand U13640 (N_13640,N_10741,N_11887);
nand U13641 (N_13641,N_10757,N_10123);
and U13642 (N_13642,N_10415,N_10720);
or U13643 (N_13643,N_11936,N_10341);
nand U13644 (N_13644,N_11357,N_10511);
and U13645 (N_13645,N_10119,N_11648);
or U13646 (N_13646,N_10566,N_10233);
and U13647 (N_13647,N_11884,N_10543);
nand U13648 (N_13648,N_10538,N_10628);
or U13649 (N_13649,N_10325,N_10842);
nand U13650 (N_13650,N_11838,N_11441);
or U13651 (N_13651,N_11146,N_11303);
or U13652 (N_13652,N_10224,N_11091);
or U13653 (N_13653,N_10094,N_10425);
and U13654 (N_13654,N_11578,N_11493);
nor U13655 (N_13655,N_11817,N_11562);
nand U13656 (N_13656,N_10116,N_11381);
nor U13657 (N_13657,N_11396,N_10442);
and U13658 (N_13658,N_10219,N_11673);
nor U13659 (N_13659,N_11863,N_10004);
nor U13660 (N_13660,N_11037,N_10912);
nor U13661 (N_13661,N_10062,N_11585);
or U13662 (N_13662,N_11104,N_10130);
or U13663 (N_13663,N_10008,N_11833);
nand U13664 (N_13664,N_10518,N_10112);
or U13665 (N_13665,N_11101,N_10983);
nor U13666 (N_13666,N_10352,N_11348);
nand U13667 (N_13667,N_10980,N_11874);
or U13668 (N_13668,N_10766,N_10188);
nand U13669 (N_13669,N_10684,N_11533);
or U13670 (N_13670,N_10007,N_11595);
or U13671 (N_13671,N_10119,N_11283);
or U13672 (N_13672,N_10947,N_10971);
nand U13673 (N_13673,N_10254,N_11430);
xnor U13674 (N_13674,N_10223,N_11912);
nand U13675 (N_13675,N_11762,N_10751);
nor U13676 (N_13676,N_10787,N_11508);
xor U13677 (N_13677,N_11520,N_11350);
nor U13678 (N_13678,N_11103,N_10325);
nand U13679 (N_13679,N_11050,N_11215);
and U13680 (N_13680,N_10898,N_10060);
and U13681 (N_13681,N_11732,N_10100);
nor U13682 (N_13682,N_11339,N_11445);
and U13683 (N_13683,N_10037,N_11184);
xnor U13684 (N_13684,N_11456,N_11892);
xnor U13685 (N_13685,N_10016,N_10372);
and U13686 (N_13686,N_10505,N_10319);
and U13687 (N_13687,N_11646,N_11083);
xor U13688 (N_13688,N_11967,N_11633);
and U13689 (N_13689,N_11682,N_10592);
and U13690 (N_13690,N_10373,N_10692);
nand U13691 (N_13691,N_10867,N_10215);
or U13692 (N_13692,N_11475,N_11953);
and U13693 (N_13693,N_10460,N_10428);
and U13694 (N_13694,N_11521,N_10542);
or U13695 (N_13695,N_11136,N_10932);
nor U13696 (N_13696,N_11623,N_10215);
and U13697 (N_13697,N_10918,N_11261);
nor U13698 (N_13698,N_11873,N_11826);
xor U13699 (N_13699,N_11410,N_11748);
and U13700 (N_13700,N_10174,N_11312);
or U13701 (N_13701,N_10700,N_10715);
or U13702 (N_13702,N_10068,N_10884);
nor U13703 (N_13703,N_10820,N_10900);
nor U13704 (N_13704,N_11763,N_11700);
nor U13705 (N_13705,N_11079,N_10909);
nor U13706 (N_13706,N_11743,N_10302);
xor U13707 (N_13707,N_10193,N_10728);
nand U13708 (N_13708,N_10292,N_10303);
and U13709 (N_13709,N_11364,N_11154);
nor U13710 (N_13710,N_11886,N_10124);
nor U13711 (N_13711,N_11395,N_10551);
nand U13712 (N_13712,N_10934,N_10961);
nor U13713 (N_13713,N_10900,N_11859);
xor U13714 (N_13714,N_10835,N_11649);
or U13715 (N_13715,N_11748,N_10046);
and U13716 (N_13716,N_11132,N_11372);
or U13717 (N_13717,N_10368,N_10945);
nor U13718 (N_13718,N_10944,N_10769);
nand U13719 (N_13719,N_11388,N_11838);
xor U13720 (N_13720,N_10159,N_11608);
nand U13721 (N_13721,N_11436,N_10557);
xnor U13722 (N_13722,N_10576,N_11588);
nor U13723 (N_13723,N_10777,N_10913);
xor U13724 (N_13724,N_10632,N_10376);
nand U13725 (N_13725,N_10178,N_10892);
and U13726 (N_13726,N_11292,N_10203);
xnor U13727 (N_13727,N_10095,N_10028);
xnor U13728 (N_13728,N_11551,N_11146);
xnor U13729 (N_13729,N_11048,N_11993);
and U13730 (N_13730,N_10950,N_11977);
nand U13731 (N_13731,N_10058,N_11807);
xor U13732 (N_13732,N_10304,N_10311);
and U13733 (N_13733,N_11993,N_10922);
nor U13734 (N_13734,N_11313,N_10273);
or U13735 (N_13735,N_10125,N_10333);
and U13736 (N_13736,N_10468,N_10228);
nand U13737 (N_13737,N_10465,N_10493);
nand U13738 (N_13738,N_11643,N_11580);
xnor U13739 (N_13739,N_11936,N_10648);
or U13740 (N_13740,N_10928,N_11693);
nand U13741 (N_13741,N_10584,N_11683);
or U13742 (N_13742,N_11902,N_10426);
nor U13743 (N_13743,N_11683,N_11718);
nand U13744 (N_13744,N_11465,N_10966);
nand U13745 (N_13745,N_11857,N_11768);
xnor U13746 (N_13746,N_11469,N_10666);
and U13747 (N_13747,N_10527,N_11152);
and U13748 (N_13748,N_11462,N_11945);
nand U13749 (N_13749,N_11191,N_10073);
or U13750 (N_13750,N_11714,N_11083);
or U13751 (N_13751,N_11821,N_10531);
and U13752 (N_13752,N_10222,N_11733);
nor U13753 (N_13753,N_10502,N_10205);
nand U13754 (N_13754,N_11043,N_10735);
nand U13755 (N_13755,N_11616,N_11728);
and U13756 (N_13756,N_10680,N_10567);
nor U13757 (N_13757,N_11045,N_10899);
and U13758 (N_13758,N_11788,N_10769);
or U13759 (N_13759,N_11884,N_10618);
xnor U13760 (N_13760,N_10805,N_10306);
or U13761 (N_13761,N_11456,N_11141);
nor U13762 (N_13762,N_10966,N_10719);
or U13763 (N_13763,N_11864,N_11285);
xor U13764 (N_13764,N_11756,N_10094);
xnor U13765 (N_13765,N_10877,N_11914);
nand U13766 (N_13766,N_11523,N_11683);
and U13767 (N_13767,N_10201,N_11383);
nand U13768 (N_13768,N_11703,N_11295);
nor U13769 (N_13769,N_10731,N_11950);
xnor U13770 (N_13770,N_11172,N_11671);
and U13771 (N_13771,N_10678,N_10407);
and U13772 (N_13772,N_10870,N_11328);
nand U13773 (N_13773,N_11803,N_10004);
nor U13774 (N_13774,N_10406,N_10084);
nand U13775 (N_13775,N_11089,N_10611);
and U13776 (N_13776,N_10330,N_10465);
and U13777 (N_13777,N_11937,N_10590);
and U13778 (N_13778,N_10891,N_10414);
nand U13779 (N_13779,N_10512,N_11607);
xnor U13780 (N_13780,N_11498,N_11654);
or U13781 (N_13781,N_11995,N_11629);
or U13782 (N_13782,N_10040,N_11762);
xnor U13783 (N_13783,N_10751,N_10219);
nand U13784 (N_13784,N_11278,N_11785);
xnor U13785 (N_13785,N_10596,N_11671);
xnor U13786 (N_13786,N_11434,N_10305);
nand U13787 (N_13787,N_11615,N_10282);
and U13788 (N_13788,N_11259,N_11552);
or U13789 (N_13789,N_10354,N_11840);
nand U13790 (N_13790,N_10834,N_11631);
xnor U13791 (N_13791,N_10128,N_10341);
nor U13792 (N_13792,N_10718,N_10581);
nor U13793 (N_13793,N_11324,N_11476);
xnor U13794 (N_13794,N_11006,N_10966);
nor U13795 (N_13795,N_10432,N_11971);
xnor U13796 (N_13796,N_10397,N_10288);
xnor U13797 (N_13797,N_10690,N_10091);
and U13798 (N_13798,N_10794,N_11462);
nand U13799 (N_13799,N_10467,N_10670);
or U13800 (N_13800,N_10425,N_11019);
nand U13801 (N_13801,N_10554,N_10616);
nand U13802 (N_13802,N_11553,N_11913);
or U13803 (N_13803,N_10442,N_10110);
nand U13804 (N_13804,N_11605,N_11696);
nand U13805 (N_13805,N_10614,N_11845);
or U13806 (N_13806,N_10689,N_10273);
and U13807 (N_13807,N_11466,N_11598);
nor U13808 (N_13808,N_11128,N_11524);
nand U13809 (N_13809,N_10134,N_11290);
or U13810 (N_13810,N_10346,N_11070);
nand U13811 (N_13811,N_10413,N_10799);
nor U13812 (N_13812,N_11190,N_10712);
and U13813 (N_13813,N_10269,N_11755);
nand U13814 (N_13814,N_10602,N_11609);
and U13815 (N_13815,N_11338,N_11142);
xor U13816 (N_13816,N_11713,N_11220);
and U13817 (N_13817,N_11399,N_10317);
nand U13818 (N_13818,N_10658,N_10361);
xor U13819 (N_13819,N_11689,N_11247);
nor U13820 (N_13820,N_11436,N_11943);
and U13821 (N_13821,N_10790,N_10274);
or U13822 (N_13822,N_11682,N_10316);
xnor U13823 (N_13823,N_11512,N_10298);
nor U13824 (N_13824,N_11070,N_11705);
and U13825 (N_13825,N_10872,N_10164);
xnor U13826 (N_13826,N_11953,N_11879);
xor U13827 (N_13827,N_10754,N_11550);
xnor U13828 (N_13828,N_11300,N_10278);
or U13829 (N_13829,N_10685,N_10543);
and U13830 (N_13830,N_10639,N_10883);
or U13831 (N_13831,N_10629,N_11839);
or U13832 (N_13832,N_11427,N_11215);
or U13833 (N_13833,N_11785,N_11361);
or U13834 (N_13834,N_10034,N_11112);
nor U13835 (N_13835,N_11679,N_10740);
or U13836 (N_13836,N_10142,N_10303);
nand U13837 (N_13837,N_11566,N_11928);
nand U13838 (N_13838,N_11808,N_11076);
nand U13839 (N_13839,N_10901,N_11480);
xor U13840 (N_13840,N_11692,N_11334);
nor U13841 (N_13841,N_10092,N_11882);
xor U13842 (N_13842,N_10601,N_11830);
or U13843 (N_13843,N_11116,N_11547);
or U13844 (N_13844,N_10574,N_11911);
nor U13845 (N_13845,N_11713,N_11777);
xor U13846 (N_13846,N_11090,N_10164);
or U13847 (N_13847,N_10278,N_11863);
nand U13848 (N_13848,N_10002,N_10475);
nand U13849 (N_13849,N_10802,N_10687);
nor U13850 (N_13850,N_10931,N_10259);
nand U13851 (N_13851,N_10042,N_10030);
xnor U13852 (N_13852,N_10295,N_11381);
nor U13853 (N_13853,N_11494,N_11158);
nor U13854 (N_13854,N_11604,N_10381);
and U13855 (N_13855,N_11584,N_10760);
nor U13856 (N_13856,N_10257,N_11002);
nor U13857 (N_13857,N_10947,N_10370);
nor U13858 (N_13858,N_11026,N_11667);
and U13859 (N_13859,N_11449,N_11381);
xor U13860 (N_13860,N_10494,N_11020);
nand U13861 (N_13861,N_10888,N_10827);
xor U13862 (N_13862,N_11525,N_11819);
and U13863 (N_13863,N_11176,N_10143);
nand U13864 (N_13864,N_10031,N_11004);
and U13865 (N_13865,N_11438,N_10526);
or U13866 (N_13866,N_11774,N_10545);
or U13867 (N_13867,N_10741,N_11680);
and U13868 (N_13868,N_11633,N_10619);
xor U13869 (N_13869,N_10172,N_11924);
and U13870 (N_13870,N_11505,N_10545);
xnor U13871 (N_13871,N_10811,N_11300);
nand U13872 (N_13872,N_10813,N_11935);
nand U13873 (N_13873,N_10172,N_11964);
nand U13874 (N_13874,N_11992,N_10993);
nor U13875 (N_13875,N_10392,N_10177);
or U13876 (N_13876,N_10996,N_10370);
nand U13877 (N_13877,N_11425,N_11843);
xor U13878 (N_13878,N_10405,N_11270);
nor U13879 (N_13879,N_10680,N_11053);
and U13880 (N_13880,N_10348,N_11590);
nand U13881 (N_13881,N_10456,N_10562);
and U13882 (N_13882,N_10487,N_10395);
and U13883 (N_13883,N_10057,N_10641);
xnor U13884 (N_13884,N_11265,N_10012);
xor U13885 (N_13885,N_10738,N_11790);
nand U13886 (N_13886,N_11319,N_11643);
xnor U13887 (N_13887,N_11549,N_10581);
xor U13888 (N_13888,N_11368,N_10678);
nor U13889 (N_13889,N_10788,N_11623);
nand U13890 (N_13890,N_10042,N_11297);
or U13891 (N_13891,N_11918,N_11463);
nand U13892 (N_13892,N_11696,N_10863);
nand U13893 (N_13893,N_11913,N_10126);
nor U13894 (N_13894,N_10451,N_11365);
nor U13895 (N_13895,N_11771,N_10703);
nor U13896 (N_13896,N_10934,N_11625);
xnor U13897 (N_13897,N_11989,N_10570);
nor U13898 (N_13898,N_10688,N_10701);
xnor U13899 (N_13899,N_10977,N_11454);
nor U13900 (N_13900,N_11114,N_10570);
xor U13901 (N_13901,N_11360,N_10015);
or U13902 (N_13902,N_10839,N_11051);
nor U13903 (N_13903,N_10189,N_11230);
nand U13904 (N_13904,N_10132,N_10702);
or U13905 (N_13905,N_11527,N_10615);
xnor U13906 (N_13906,N_11769,N_11730);
nand U13907 (N_13907,N_10363,N_11886);
nor U13908 (N_13908,N_10156,N_11136);
nor U13909 (N_13909,N_11780,N_10157);
or U13910 (N_13910,N_10471,N_10173);
and U13911 (N_13911,N_11821,N_11590);
or U13912 (N_13912,N_10943,N_11565);
xor U13913 (N_13913,N_10277,N_10300);
or U13914 (N_13914,N_10997,N_11213);
and U13915 (N_13915,N_10707,N_10836);
and U13916 (N_13916,N_11367,N_11961);
nand U13917 (N_13917,N_11718,N_11844);
and U13918 (N_13918,N_11519,N_11280);
nand U13919 (N_13919,N_11767,N_10081);
nand U13920 (N_13920,N_10892,N_10721);
xor U13921 (N_13921,N_11384,N_11065);
nand U13922 (N_13922,N_11077,N_10902);
xor U13923 (N_13923,N_11353,N_11175);
and U13924 (N_13924,N_11824,N_11948);
nor U13925 (N_13925,N_11074,N_10078);
nor U13926 (N_13926,N_11774,N_10203);
or U13927 (N_13927,N_11997,N_10174);
and U13928 (N_13928,N_10131,N_10974);
and U13929 (N_13929,N_10321,N_11030);
nand U13930 (N_13930,N_11493,N_11281);
xor U13931 (N_13931,N_11971,N_11177);
nand U13932 (N_13932,N_11755,N_10635);
or U13933 (N_13933,N_11380,N_10388);
or U13934 (N_13934,N_10554,N_10633);
xor U13935 (N_13935,N_11209,N_11356);
xor U13936 (N_13936,N_10561,N_11310);
or U13937 (N_13937,N_11209,N_11702);
and U13938 (N_13938,N_10806,N_10174);
nand U13939 (N_13939,N_10936,N_10332);
nor U13940 (N_13940,N_11289,N_10670);
xor U13941 (N_13941,N_11984,N_10454);
xor U13942 (N_13942,N_11628,N_10979);
nor U13943 (N_13943,N_11122,N_11733);
nand U13944 (N_13944,N_11499,N_10840);
or U13945 (N_13945,N_10234,N_10476);
nor U13946 (N_13946,N_10405,N_10774);
and U13947 (N_13947,N_11888,N_11950);
xor U13948 (N_13948,N_11272,N_10809);
or U13949 (N_13949,N_11321,N_11533);
nor U13950 (N_13950,N_10852,N_11374);
xnor U13951 (N_13951,N_11617,N_11912);
xor U13952 (N_13952,N_11996,N_10736);
and U13953 (N_13953,N_10336,N_10049);
or U13954 (N_13954,N_11700,N_10191);
xnor U13955 (N_13955,N_10431,N_10016);
xnor U13956 (N_13956,N_11363,N_10105);
xor U13957 (N_13957,N_10538,N_11791);
xor U13958 (N_13958,N_10125,N_10017);
or U13959 (N_13959,N_11804,N_11880);
or U13960 (N_13960,N_10544,N_11368);
xnor U13961 (N_13961,N_10162,N_11539);
nor U13962 (N_13962,N_11057,N_10058);
nor U13963 (N_13963,N_10454,N_10295);
nor U13964 (N_13964,N_11439,N_11382);
nor U13965 (N_13965,N_10562,N_11770);
or U13966 (N_13966,N_10872,N_11569);
xnor U13967 (N_13967,N_10972,N_11268);
nand U13968 (N_13968,N_10868,N_10540);
and U13969 (N_13969,N_10640,N_10973);
nand U13970 (N_13970,N_11948,N_10985);
nor U13971 (N_13971,N_10662,N_11308);
nand U13972 (N_13972,N_11343,N_11414);
or U13973 (N_13973,N_11537,N_10242);
or U13974 (N_13974,N_11044,N_10073);
or U13975 (N_13975,N_11357,N_11939);
or U13976 (N_13976,N_10487,N_11583);
or U13977 (N_13977,N_11083,N_11079);
and U13978 (N_13978,N_10772,N_11117);
nand U13979 (N_13979,N_10056,N_11519);
nand U13980 (N_13980,N_10872,N_11166);
nor U13981 (N_13981,N_10585,N_11571);
nand U13982 (N_13982,N_11826,N_11513);
or U13983 (N_13983,N_10556,N_10293);
or U13984 (N_13984,N_11731,N_10026);
nand U13985 (N_13985,N_10012,N_10509);
or U13986 (N_13986,N_11030,N_10749);
nand U13987 (N_13987,N_10438,N_10665);
and U13988 (N_13988,N_11661,N_11924);
or U13989 (N_13989,N_10676,N_10217);
xor U13990 (N_13990,N_10751,N_10672);
and U13991 (N_13991,N_10994,N_11848);
and U13992 (N_13992,N_10888,N_11524);
nor U13993 (N_13993,N_10932,N_11760);
nand U13994 (N_13994,N_10268,N_10466);
or U13995 (N_13995,N_10016,N_11107);
or U13996 (N_13996,N_10438,N_10796);
and U13997 (N_13997,N_10439,N_11108);
or U13998 (N_13998,N_10276,N_10976);
xor U13999 (N_13999,N_11557,N_10368);
xnor U14000 (N_14000,N_12352,N_13219);
or U14001 (N_14001,N_13454,N_12406);
nor U14002 (N_14002,N_13433,N_12617);
or U14003 (N_14003,N_13377,N_12277);
nand U14004 (N_14004,N_12905,N_13175);
and U14005 (N_14005,N_13207,N_12467);
nand U14006 (N_14006,N_13167,N_12493);
nand U14007 (N_14007,N_12180,N_13719);
nand U14008 (N_14008,N_12949,N_12935);
or U14009 (N_14009,N_13336,N_12466);
and U14010 (N_14010,N_12407,N_12542);
nand U14011 (N_14011,N_12117,N_13416);
nor U14012 (N_14012,N_12041,N_13914);
or U14013 (N_14013,N_12890,N_13569);
nand U14014 (N_14014,N_13143,N_12438);
xor U14015 (N_14015,N_13678,N_12071);
and U14016 (N_14016,N_13390,N_13032);
xnor U14017 (N_14017,N_12669,N_13652);
nor U14018 (N_14018,N_13113,N_12484);
and U14019 (N_14019,N_12588,N_12834);
and U14020 (N_14020,N_12820,N_13585);
xnor U14021 (N_14021,N_12631,N_12366);
and U14022 (N_14022,N_13685,N_13999);
nor U14023 (N_14023,N_13758,N_12763);
and U14024 (N_14024,N_12769,N_13245);
xnor U14025 (N_14025,N_12274,N_12263);
nand U14026 (N_14026,N_13636,N_12231);
and U14027 (N_14027,N_13275,N_12673);
nand U14028 (N_14028,N_12513,N_12887);
nor U14029 (N_14029,N_12557,N_13949);
and U14030 (N_14030,N_13943,N_12951);
and U14031 (N_14031,N_12559,N_12402);
or U14032 (N_14032,N_13910,N_13957);
nor U14033 (N_14033,N_13936,N_13461);
or U14034 (N_14034,N_12325,N_12239);
or U14035 (N_14035,N_13791,N_12634);
or U14036 (N_14036,N_13996,N_13519);
nand U14037 (N_14037,N_13903,N_12482);
and U14038 (N_14038,N_13503,N_13169);
nor U14039 (N_14039,N_12595,N_13002);
xor U14040 (N_14040,N_13887,N_13812);
nor U14041 (N_14041,N_13820,N_12740);
xor U14042 (N_14042,N_12236,N_12767);
xor U14043 (N_14043,N_13225,N_13331);
and U14044 (N_14044,N_13562,N_12167);
and U14045 (N_14045,N_12056,N_12799);
xor U14046 (N_14046,N_13967,N_13590);
nor U14047 (N_14047,N_12100,N_13201);
and U14048 (N_14048,N_13299,N_13119);
or U14049 (N_14049,N_12479,N_12967);
nand U14050 (N_14050,N_12638,N_12289);
or U14051 (N_14051,N_13620,N_13923);
nor U14052 (N_14052,N_13533,N_12005);
nor U14053 (N_14053,N_13989,N_13828);
or U14054 (N_14054,N_13558,N_13890);
xnor U14055 (N_14055,N_13520,N_13932);
and U14056 (N_14056,N_12627,N_12343);
nor U14057 (N_14057,N_13718,N_13930);
nand U14058 (N_14058,N_12684,N_13467);
nor U14059 (N_14059,N_13861,N_13640);
or U14060 (N_14060,N_13852,N_12516);
or U14061 (N_14061,N_12065,N_12973);
xnor U14062 (N_14062,N_13919,N_13310);
xor U14063 (N_14063,N_12353,N_13628);
and U14064 (N_14064,N_13931,N_12349);
or U14065 (N_14065,N_12911,N_12830);
nand U14066 (N_14066,N_13252,N_12704);
and U14067 (N_14067,N_13388,N_13609);
or U14068 (N_14068,N_12988,N_12835);
nor U14069 (N_14069,N_12428,N_12031);
and U14070 (N_14070,N_12320,N_12321);
and U14071 (N_14071,N_12028,N_12166);
xnor U14072 (N_14072,N_12546,N_12360);
or U14073 (N_14073,N_13907,N_13523);
or U14074 (N_14074,N_12938,N_13899);
xor U14075 (N_14075,N_13320,N_12244);
nor U14076 (N_14076,N_13742,N_12375);
xnor U14077 (N_14077,N_13840,N_12391);
or U14078 (N_14078,N_13356,N_13613);
xor U14079 (N_14079,N_12473,N_12630);
nand U14080 (N_14080,N_13663,N_13309);
nor U14081 (N_14081,N_13551,N_13060);
nor U14082 (N_14082,N_13363,N_12899);
and U14083 (N_14083,N_13220,N_12223);
or U14084 (N_14084,N_13626,N_13093);
nand U14085 (N_14085,N_13816,N_12163);
nand U14086 (N_14086,N_13328,N_13529);
or U14087 (N_14087,N_13394,N_12836);
nor U14088 (N_14088,N_13401,N_12333);
nor U14089 (N_14089,N_13793,N_13925);
or U14090 (N_14090,N_13188,N_13535);
nor U14091 (N_14091,N_13350,N_13653);
nor U14092 (N_14092,N_13397,N_12765);
nor U14093 (N_14093,N_12145,N_13070);
nor U14094 (N_14094,N_13170,N_12910);
and U14095 (N_14095,N_13236,N_12014);
xor U14096 (N_14096,N_12586,N_13778);
nor U14097 (N_14097,N_13030,N_12664);
nor U14098 (N_14098,N_12114,N_12398);
nor U14099 (N_14099,N_13035,N_12152);
nand U14100 (N_14100,N_12011,N_12787);
nor U14101 (N_14101,N_13057,N_13422);
xnor U14102 (N_14102,N_12917,N_12661);
nand U14103 (N_14103,N_12731,N_12535);
nor U14104 (N_14104,N_12556,N_12703);
nor U14105 (N_14105,N_12168,N_13571);
and U14106 (N_14106,N_13696,N_13260);
or U14107 (N_14107,N_12581,N_13807);
or U14108 (N_14108,N_13884,N_13049);
or U14109 (N_14109,N_12544,N_13792);
and U14110 (N_14110,N_12217,N_12069);
and U14111 (N_14111,N_12299,N_13679);
xnor U14112 (N_14112,N_13763,N_13954);
nand U14113 (N_14113,N_12894,N_12040);
nand U14114 (N_14114,N_12316,N_13565);
xor U14115 (N_14115,N_13818,N_12936);
nand U14116 (N_14116,N_13273,N_13315);
xor U14117 (N_14117,N_13728,N_12611);
or U14118 (N_14118,N_12857,N_13532);
xnor U14119 (N_14119,N_12429,N_13318);
and U14120 (N_14120,N_12816,N_12810);
nand U14121 (N_14121,N_13958,N_13959);
or U14122 (N_14122,N_12749,N_12623);
nand U14123 (N_14123,N_13159,N_12301);
nor U14124 (N_14124,N_12790,N_12906);
nand U14125 (N_14125,N_13337,N_13625);
nor U14126 (N_14126,N_12379,N_12999);
xnor U14127 (N_14127,N_13425,N_13817);
xor U14128 (N_14128,N_12587,N_12425);
nor U14129 (N_14129,N_12435,N_13575);
nand U14130 (N_14130,N_13830,N_13133);
xnor U14131 (N_14131,N_13434,N_12753);
or U14132 (N_14132,N_12451,N_12296);
and U14133 (N_14133,N_12311,N_12807);
nand U14134 (N_14134,N_12276,N_12018);
and U14135 (N_14135,N_13115,N_13526);
or U14136 (N_14136,N_13549,N_13302);
xor U14137 (N_14137,N_13511,N_13018);
and U14138 (N_14138,N_12880,N_13716);
nor U14139 (N_14139,N_12463,N_13373);
nand U14140 (N_14140,N_12786,N_12009);
or U14141 (N_14141,N_12013,N_13859);
nand U14142 (N_14142,N_13886,N_13915);
nand U14143 (N_14143,N_13501,N_12101);
xnor U14144 (N_14144,N_13703,N_13432);
and U14145 (N_14145,N_13136,N_12373);
xor U14146 (N_14146,N_12965,N_12446);
xnor U14147 (N_14147,N_13016,N_13655);
nor U14148 (N_14148,N_13598,N_12002);
nor U14149 (N_14149,N_12308,N_12222);
xnor U14150 (N_14150,N_12822,N_12827);
or U14151 (N_14151,N_12869,N_13146);
xor U14152 (N_14152,N_13068,N_12157);
and U14153 (N_14153,N_13005,N_13749);
nor U14154 (N_14154,N_12972,N_12351);
and U14155 (N_14155,N_13942,N_12777);
nand U14156 (N_14156,N_13627,N_13122);
nand U14157 (N_14157,N_13011,N_13721);
xor U14158 (N_14158,N_13646,N_13864);
xnor U14159 (N_14159,N_13662,N_12292);
nand U14160 (N_14160,N_13066,N_12449);
nand U14161 (N_14161,N_13516,N_12498);
nand U14162 (N_14162,N_13781,N_12327);
nor U14163 (N_14163,N_13645,N_13379);
and U14164 (N_14164,N_12707,N_12464);
and U14165 (N_14165,N_12895,N_12250);
nor U14166 (N_14166,N_12750,N_12698);
nor U14167 (N_14167,N_12653,N_13798);
xor U14168 (N_14168,N_13047,N_12247);
nor U14169 (N_14169,N_12568,N_13405);
nor U14170 (N_14170,N_12229,N_13358);
xor U14171 (N_14171,N_12019,N_12893);
xnor U14172 (N_14172,N_13973,N_12651);
xor U14173 (N_14173,N_13223,N_12552);
and U14174 (N_14174,N_13810,N_13280);
nand U14175 (N_14175,N_13051,N_13862);
xor U14176 (N_14176,N_12758,N_12491);
nand U14177 (N_14177,N_13021,N_13517);
xnor U14178 (N_14178,N_13301,N_12717);
nand U14179 (N_14179,N_12187,N_12162);
nor U14180 (N_14180,N_12774,N_12043);
xor U14181 (N_14181,N_12642,N_13063);
and U14182 (N_14182,N_13956,N_13823);
or U14183 (N_14183,N_12113,N_13217);
or U14184 (N_14184,N_12297,N_13192);
or U14185 (N_14185,N_13563,N_13720);
or U14186 (N_14186,N_13960,N_12317);
or U14187 (N_14187,N_12723,N_12334);
or U14188 (N_14188,N_13286,N_12992);
nor U14189 (N_14189,N_13058,N_13776);
or U14190 (N_14190,N_13639,N_13471);
and U14191 (N_14191,N_13493,N_13908);
or U14192 (N_14192,N_12017,N_12415);
or U14193 (N_14193,N_12455,N_12024);
nand U14194 (N_14194,N_13968,N_12298);
or U14195 (N_14195,N_13061,N_12243);
or U14196 (N_14196,N_13661,N_13492);
xnor U14197 (N_14197,N_13607,N_13616);
and U14198 (N_14198,N_13298,N_12878);
or U14199 (N_14199,N_12094,N_13633);
xnor U14200 (N_14200,N_13868,N_13022);
and U14201 (N_14201,N_12813,N_12189);
xor U14202 (N_14202,N_13677,N_12452);
nor U14203 (N_14203,N_13153,N_12424);
xor U14204 (N_14204,N_13155,N_13335);
and U14205 (N_14205,N_12279,N_13597);
and U14206 (N_14206,N_13477,N_13962);
xor U14207 (N_14207,N_13991,N_12626);
xnor U14208 (N_14208,N_13213,N_13615);
or U14209 (N_14209,N_12092,N_12440);
or U14210 (N_14210,N_12097,N_12105);
nand U14211 (N_14211,N_13249,N_13567);
and U14212 (N_14212,N_13650,N_13450);
xor U14213 (N_14213,N_13193,N_12719);
nor U14214 (N_14214,N_13088,N_12460);
nand U14215 (N_14215,N_12676,N_13067);
and U14216 (N_14216,N_12420,N_12959);
or U14217 (N_14217,N_13787,N_13755);
or U14218 (N_14218,N_13888,N_12561);
nand U14219 (N_14219,N_13893,N_13824);
xor U14220 (N_14220,N_12048,N_12583);
and U14221 (N_14221,N_13024,N_13085);
and U14222 (N_14222,N_12049,N_13026);
xnor U14223 (N_14223,N_13997,N_12828);
or U14224 (N_14224,N_12671,N_13630);
or U14225 (N_14225,N_13165,N_13218);
and U14226 (N_14226,N_12132,N_13419);
xnor U14227 (N_14227,N_12487,N_13885);
xnor U14228 (N_14228,N_13483,N_12710);
xnor U14229 (N_14229,N_12730,N_12982);
xnor U14230 (N_14230,N_13059,N_13319);
nor U14231 (N_14231,N_13684,N_12171);
nand U14232 (N_14232,N_13889,N_12129);
and U14233 (N_14233,N_13330,N_13077);
or U14234 (N_14234,N_12332,N_12093);
or U14235 (N_14235,N_12958,N_12668);
nand U14236 (N_14236,N_13579,N_12852);
nand U14237 (N_14237,N_13995,N_12253);
nand U14238 (N_14238,N_13871,N_13029);
or U14239 (N_14239,N_13242,N_13896);
xor U14240 (N_14240,N_13210,N_12971);
and U14241 (N_14241,N_13349,N_12036);
or U14242 (N_14242,N_13322,N_12739);
or U14243 (N_14243,N_13687,N_13025);
or U14244 (N_14244,N_12089,N_12411);
nor U14245 (N_14245,N_12198,N_12732);
and U14246 (N_14246,N_12670,N_12396);
nand U14247 (N_14247,N_12395,N_13012);
nor U14248 (N_14248,N_13521,N_13439);
xor U14249 (N_14249,N_12979,N_12590);
or U14250 (N_14250,N_13736,N_13782);
xor U14251 (N_14251,N_12335,N_13481);
and U14252 (N_14252,N_13353,N_13268);
xor U14253 (N_14253,N_12675,N_13806);
xor U14254 (N_14254,N_13438,N_13668);
or U14255 (N_14255,N_12682,N_13911);
xnor U14256 (N_14256,N_12647,N_12580);
and U14257 (N_14257,N_12563,N_13140);
nor U14258 (N_14258,N_13504,N_13431);
or U14259 (N_14259,N_12752,N_12862);
or U14260 (N_14260,N_13667,N_12800);
or U14261 (N_14261,N_13804,N_12471);
nor U14262 (N_14262,N_12712,N_12439);
nand U14263 (N_14263,N_12448,N_12672);
nand U14264 (N_14264,N_12727,N_12416);
or U14265 (N_14265,N_13324,N_12578);
nor U14266 (N_14266,N_13568,N_13040);
or U14267 (N_14267,N_13104,N_13171);
nand U14268 (N_14268,N_13725,N_12868);
nor U14269 (N_14269,N_12986,N_12576);
nand U14270 (N_14270,N_13819,N_13935);
or U14271 (N_14271,N_13497,N_13612);
nand U14272 (N_14272,N_12771,N_12004);
xnor U14273 (N_14273,N_12294,N_13842);
xnor U14274 (N_14274,N_12068,N_13970);
xor U14275 (N_14275,N_12457,N_12264);
nand U14276 (N_14276,N_12855,N_12135);
xnor U14277 (N_14277,N_12122,N_12278);
nand U14278 (N_14278,N_13775,N_13710);
nand U14279 (N_14279,N_12064,N_12437);
or U14280 (N_14280,N_13922,N_12572);
and U14281 (N_14281,N_13745,N_13065);
nor U14282 (N_14282,N_13897,N_12687);
and U14283 (N_14283,N_13339,N_13586);
xor U14284 (N_14284,N_13230,N_12692);
nor U14285 (N_14285,N_12007,N_12314);
or U14286 (N_14286,N_12430,N_12228);
nand U14287 (N_14287,N_12271,N_12205);
or U14288 (N_14288,N_12729,N_12077);
or U14289 (N_14289,N_12888,N_12536);
nand U14290 (N_14290,N_12981,N_12322);
or U14291 (N_14291,N_12442,N_12522);
and U14292 (N_14292,N_13580,N_12176);
xor U14293 (N_14293,N_13634,N_13785);
xor U14294 (N_14294,N_13611,N_13447);
nand U14295 (N_14295,N_13478,N_12543);
or U14296 (N_14296,N_13163,N_13333);
nand U14297 (N_14297,N_12609,N_12526);
nor U14298 (N_14298,N_13003,N_13705);
nand U14299 (N_14299,N_12112,N_13891);
nand U14300 (N_14300,N_13559,N_12038);
nand U14301 (N_14301,N_13131,N_13451);
and U14302 (N_14302,N_12921,N_12137);
xnor U14303 (N_14303,N_13768,N_13821);
nand U14304 (N_14304,N_13635,N_12738);
and U14305 (N_14305,N_12047,N_13969);
and U14306 (N_14306,N_12261,N_13622);
xor U14307 (N_14307,N_13283,N_12284);
nand U14308 (N_14308,N_13894,N_13524);
xor U14309 (N_14309,N_12474,N_13654);
nor U14310 (N_14310,N_12884,N_13259);
nor U14311 (N_14311,N_12804,N_12185);
and U14312 (N_14312,N_12136,N_12160);
and U14313 (N_14313,N_12833,N_13522);
nor U14314 (N_14314,N_13534,N_12705);
nand U14315 (N_14315,N_12238,N_13518);
nand U14316 (N_14316,N_13396,N_13340);
and U14317 (N_14317,N_12225,N_13424);
and U14318 (N_14318,N_13883,N_13152);
nor U14319 (N_14319,N_12128,N_13378);
and U14320 (N_14320,N_13099,N_12523);
and U14321 (N_14321,N_12532,N_12268);
and U14322 (N_14322,N_13091,N_12197);
nor U14323 (N_14323,N_12216,N_12757);
xnor U14324 (N_14324,N_12748,N_13987);
nand U14325 (N_14325,N_12764,N_12119);
nand U14326 (N_14326,N_13050,N_13946);
nor U14327 (N_14327,N_13010,N_12643);
or U14328 (N_14328,N_13494,N_12377);
or U14329 (N_14329,N_12659,N_12809);
or U14330 (N_14330,N_12579,N_12472);
and U14331 (N_14331,N_13711,N_12209);
or U14332 (N_14332,N_13849,N_12875);
and U14333 (N_14333,N_13649,N_12574);
and U14334 (N_14334,N_13351,N_12713);
and U14335 (N_14335,N_12995,N_13179);
or U14336 (N_14336,N_12423,N_12055);
or U14337 (N_14337,N_13966,N_13542);
and U14338 (N_14338,N_12272,N_13387);
xor U14339 (N_14339,N_13553,N_13458);
and U14340 (N_14340,N_13561,N_12363);
nand U14341 (N_14341,N_13994,N_12368);
and U14342 (N_14342,N_13411,N_12770);
and U14343 (N_14343,N_12920,N_12076);
nand U14344 (N_14344,N_12666,N_12916);
and U14345 (N_14345,N_12255,N_13566);
xor U14346 (N_14346,N_13069,N_13407);
xnor U14347 (N_14347,N_12519,N_12208);
nor U14348 (N_14348,N_13296,N_12215);
xor U14349 (N_14349,N_13028,N_12956);
nand U14350 (N_14350,N_13362,N_13502);
nor U14351 (N_14351,N_12213,N_12636);
or U14352 (N_14352,N_12953,N_12148);
nor U14353 (N_14353,N_13241,N_13777);
and U14354 (N_14354,N_12389,N_13726);
or U14355 (N_14355,N_12369,N_13581);
or U14356 (N_14356,N_12600,N_12560);
or U14357 (N_14357,N_12831,N_12248);
and U14358 (N_14358,N_12848,N_13248);
xnor U14359 (N_14359,N_12364,N_12450);
nor U14360 (N_14360,N_13371,N_12326);
and U14361 (N_14361,N_13641,N_12497);
nand U14362 (N_14362,N_13090,N_12746);
and U14363 (N_14363,N_12633,N_13345);
nor U14364 (N_14364,N_12371,N_13110);
or U14365 (N_14365,N_13314,N_12404);
xor U14366 (N_14366,N_13409,N_13708);
nand U14367 (N_14367,N_13980,N_13554);
nand U14368 (N_14368,N_12020,N_13948);
nand U14369 (N_14369,N_13666,N_12612);
nand U14370 (N_14370,N_13114,N_13863);
nand U14371 (N_14371,N_12825,N_12507);
or U14372 (N_14372,N_13488,N_12681);
and U14373 (N_14373,N_12978,N_13937);
xnor U14374 (N_14374,N_12859,N_13109);
nor U14375 (N_14375,N_13097,N_13197);
nand U14376 (N_14376,N_12747,N_12086);
xnor U14377 (N_14377,N_13186,N_13490);
and U14378 (N_14378,N_12881,N_13274);
or U14379 (N_14379,N_12454,N_13545);
and U14380 (N_14380,N_12251,N_13130);
xnor U14381 (N_14381,N_13499,N_13469);
nand U14382 (N_14382,N_12146,N_12340);
nand U14383 (N_14383,N_12194,N_13338);
nor U14384 (N_14384,N_13799,N_13972);
and U14385 (N_14385,N_13036,N_13770);
or U14386 (N_14386,N_12997,N_13227);
xor U14387 (N_14387,N_13730,N_13961);
or U14388 (N_14388,N_13858,N_12153);
nor U14389 (N_14389,N_12594,N_12742);
or U14390 (N_14390,N_12249,N_12751);
nor U14391 (N_14391,N_12801,N_13250);
and U14392 (N_14392,N_12537,N_13357);
nor U14393 (N_14393,N_12596,N_13199);
or U14394 (N_14394,N_13107,N_12331);
xnor U14395 (N_14395,N_12081,N_13006);
xor U14396 (N_14396,N_12976,N_13881);
nor U14397 (N_14397,N_13564,N_12341);
nor U14398 (N_14398,N_12791,N_13505);
or U14399 (N_14399,N_12540,N_13277);
nand U14400 (N_14400,N_13284,N_13120);
nor U14401 (N_14401,N_13142,N_13007);
or U14402 (N_14402,N_12485,N_13410);
or U14403 (N_14403,N_13160,N_13211);
nor U14404 (N_14404,N_12754,N_12840);
or U14405 (N_14405,N_13095,N_12718);
nand U14406 (N_14406,N_13832,N_12476);
nor U14407 (N_14407,N_13900,N_13232);
nor U14408 (N_14408,N_12665,N_12269);
nor U14409 (N_14409,N_13463,N_13530);
nand U14410 (N_14410,N_13045,N_12489);
and U14411 (N_14411,N_13148,N_12409);
or U14412 (N_14412,N_12195,N_12904);
or U14413 (N_14413,N_13487,N_12691);
and U14414 (N_14414,N_13865,N_13904);
and U14415 (N_14415,N_12287,N_13604);
nand U14416 (N_14416,N_13453,N_12388);
xnor U14417 (N_14417,N_13417,N_13292);
nand U14418 (N_14418,N_13593,N_12726);
nor U14419 (N_14419,N_12280,N_13573);
nor U14420 (N_14420,N_12344,N_12444);
and U14421 (N_14421,N_12610,N_12577);
or U14422 (N_14422,N_13224,N_12826);
and U14423 (N_14423,N_13311,N_13053);
xnor U14424 (N_14424,N_13669,N_12499);
nor U14425 (N_14425,N_13599,N_13389);
xor U14426 (N_14426,N_13608,N_13675);
nand U14427 (N_14427,N_13054,N_13808);
and U14428 (N_14428,N_12201,N_13084);
and U14429 (N_14429,N_13722,N_12121);
xnor U14430 (N_14430,N_12063,N_12181);
nand U14431 (N_14431,N_12057,N_13243);
nor U14432 (N_14432,N_13731,N_12948);
nand U14433 (N_14433,N_13480,N_12309);
and U14434 (N_14434,N_13360,N_13729);
nand U14435 (N_14435,N_13589,N_13951);
xnor U14436 (N_14436,N_13547,N_13676);
and U14437 (N_14437,N_13205,N_13998);
nand U14438 (N_14438,N_13413,N_13427);
xnor U14439 (N_14439,N_12381,N_13510);
xor U14440 (N_14440,N_12177,N_12734);
and U14441 (N_14441,N_13982,N_12674);
xnor U14442 (N_14442,N_12679,N_13690);
or U14443 (N_14443,N_13906,N_12188);
nor U14444 (N_14444,N_12173,N_12689);
xor U14445 (N_14445,N_12358,N_13577);
or U14446 (N_14446,N_12737,N_13103);
xor U14447 (N_14447,N_13697,N_12374);
and U14448 (N_14448,N_13237,N_12902);
or U14449 (N_14449,N_13860,N_12164);
xnor U14450 (N_14450,N_13262,N_13019);
nor U14451 (N_14451,N_13329,N_13587);
nor U14452 (N_14452,N_12073,N_13541);
nand U14453 (N_14453,N_12245,N_12422);
and U14454 (N_14454,N_12761,N_13303);
nor U14455 (N_14455,N_12170,N_12688);
and U14456 (N_14456,N_13126,N_12490);
nand U14457 (N_14457,N_12156,N_13020);
and U14458 (N_14458,N_12990,N_12974);
or U14459 (N_14459,N_13157,N_12211);
and U14460 (N_14460,N_13285,N_13180);
and U14461 (N_14461,N_13187,N_12743);
xnor U14462 (N_14462,N_12963,N_12517);
nor U14463 (N_14463,N_12006,N_12506);
nor U14464 (N_14464,N_13762,N_12903);
nand U14465 (N_14465,N_12230,N_12601);
xnor U14466 (N_14466,N_12593,N_13671);
nand U14467 (N_14467,N_13595,N_12021);
xnor U14468 (N_14468,N_13073,N_12037);
xor U14469 (N_14469,N_13064,N_13539);
nand U14470 (N_14470,N_13290,N_13557);
and U14471 (N_14471,N_13882,N_12605);
or U14472 (N_14472,N_13673,N_13592);
xor U14473 (N_14473,N_12082,N_12346);
xnor U14474 (N_14474,N_12182,N_12035);
and U14475 (N_14475,N_13624,N_12384);
and U14476 (N_14476,N_12059,N_12237);
xnor U14477 (N_14477,N_13304,N_13112);
and U14478 (N_14478,N_13572,N_12126);
nand U14479 (N_14479,N_12716,N_12591);
xnor U14480 (N_14480,N_12102,N_12789);
nor U14481 (N_14481,N_13732,N_12961);
nor U14482 (N_14482,N_13147,N_13276);
or U14483 (N_14483,N_13443,N_12923);
and U14484 (N_14484,N_12350,N_12851);
and U14485 (N_14485,N_13801,N_12257);
nor U14486 (N_14486,N_12867,N_13000);
nor U14487 (N_14487,N_12539,N_13141);
xor U14488 (N_14488,N_13717,N_12566);
and U14489 (N_14489,N_12370,N_12027);
and U14490 (N_14490,N_12735,N_13246);
xnor U14491 (N_14491,N_13263,N_12655);
nand U14492 (N_14492,N_12456,N_12138);
nor U14493 (N_14493,N_12419,N_12418);
xor U14494 (N_14494,N_12662,N_12240);
and U14495 (N_14495,N_12792,N_12599);
xor U14496 (N_14496,N_13365,N_12143);
or U14497 (N_14497,N_12202,N_13042);
or U14498 (N_14498,N_13605,N_12199);
xor U14499 (N_14499,N_12045,N_12051);
xor U14500 (N_14500,N_12829,N_13039);
or U14501 (N_14501,N_12702,N_12179);
and U14502 (N_14502,N_13015,N_12762);
nor U14503 (N_14503,N_13172,N_13149);
nand U14504 (N_14504,N_12678,N_13596);
and U14505 (N_14505,N_13437,N_12246);
nand U14506 (N_14506,N_12015,N_13295);
and U14507 (N_14507,N_12838,N_13933);
nand U14508 (N_14508,N_12426,N_13746);
nand U14509 (N_14509,N_12155,N_13741);
and U14510 (N_14510,N_12336,N_12072);
nand U14511 (N_14511,N_13209,N_13326);
or U14512 (N_14512,N_12562,N_13222);
and U14513 (N_14513,N_13766,N_12950);
xor U14514 (N_14514,N_12219,N_13934);
nand U14515 (N_14515,N_13606,N_12896);
nor U14516 (N_14516,N_12337,N_13857);
or U14517 (N_14517,N_13963,N_12741);
nor U14518 (N_14518,N_13430,N_12412);
nor U14519 (N_14519,N_13965,N_13601);
nor U14520 (N_14520,N_13917,N_13537);
xnor U14521 (N_14521,N_12414,N_13856);
or U14522 (N_14522,N_12026,N_12721);
nor U14523 (N_14523,N_13929,N_12928);
nor U14524 (N_14524,N_13603,N_12818);
or U14525 (N_14525,N_12260,N_12866);
nor U14526 (N_14526,N_12275,N_12533);
or U14527 (N_14527,N_12232,N_13198);
nor U14528 (N_14528,N_13183,N_13367);
xnor U14529 (N_14529,N_13976,N_12078);
and U14530 (N_14530,N_13964,N_12772);
nand U14531 (N_14531,N_13046,N_12150);
nand U14532 (N_14532,N_12977,N_13753);
nand U14533 (N_14533,N_12161,N_13752);
nor U14534 (N_14534,N_12553,N_13033);
nor U14535 (N_14535,N_12405,N_12776);
and U14536 (N_14536,N_12549,N_13783);
nor U14537 (N_14537,N_12806,N_13484);
nand U14538 (N_14538,N_13756,N_12115);
xnor U14539 (N_14539,N_12940,N_12053);
nor U14540 (N_14540,N_13829,N_13052);
xnor U14541 (N_14541,N_13588,N_12470);
xnor U14542 (N_14542,N_12361,N_12952);
xor U14543 (N_14543,N_12192,N_12860);
nand U14544 (N_14544,N_13658,N_13751);
xor U14545 (N_14545,N_12125,N_13709);
nor U14546 (N_14546,N_12106,N_12012);
or U14547 (N_14547,N_12547,N_12622);
nand U14548 (N_14548,N_12443,N_12025);
and U14549 (N_14549,N_13202,N_13027);
nor U14550 (N_14550,N_13121,N_12259);
or U14551 (N_14551,N_13670,N_13546);
xnor U14552 (N_14552,N_12964,N_12955);
and U14553 (N_14553,N_13444,N_13261);
and U14554 (N_14554,N_13918,N_13664);
or U14555 (N_14555,N_12481,N_13706);
nor U14556 (N_14556,N_12962,N_13233);
and U14557 (N_14557,N_12569,N_12632);
nand U14558 (N_14558,N_12032,N_13312);
nor U14559 (N_14559,N_12725,N_12110);
or U14560 (N_14560,N_12795,N_13306);
xor U14561 (N_14561,N_13185,N_12530);
nor U14562 (N_14562,N_12602,N_12385);
and U14563 (N_14563,N_12720,N_12354);
and U14564 (N_14564,N_13062,N_12159);
nor U14565 (N_14565,N_13081,N_13578);
xnor U14566 (N_14566,N_13814,N_13491);
xor U14567 (N_14567,N_12957,N_12355);
xnor U14568 (N_14568,N_12803,N_12736);
nor U14569 (N_14569,N_13347,N_13092);
xnor U14570 (N_14570,N_12483,N_13023);
xor U14571 (N_14571,N_12891,N_12494);
or U14572 (N_14572,N_12103,N_12722);
nand U14573 (N_14573,N_13154,N_12468);
nand U14574 (N_14574,N_12204,N_12987);
and U14575 (N_14575,N_13354,N_13240);
nor U14576 (N_14576,N_12847,N_12254);
xor U14577 (N_14577,N_12436,N_12515);
and U14578 (N_14578,N_13769,N_12313);
and U14579 (N_14579,N_13150,N_13985);
xor U14580 (N_14580,N_12760,N_13089);
nor U14581 (N_14581,N_12628,N_13531);
nand U14582 (N_14582,N_12066,N_13376);
nand U14583 (N_14583,N_13743,N_12323);
or U14584 (N_14584,N_12706,N_13452);
and U14585 (N_14585,N_13525,N_12714);
or U14586 (N_14586,N_12733,N_12500);
nor U14587 (N_14587,N_13257,N_13548);
nor U14588 (N_14588,N_12131,N_12879);
nor U14589 (N_14589,N_13316,N_13744);
xnor U14590 (N_14590,N_13208,N_13657);
nor U14591 (N_14591,N_13323,N_13941);
xnor U14592 (N_14592,N_13123,N_12262);
nand U14593 (N_14593,N_12447,N_12324);
xnor U14594 (N_14594,N_13445,N_13106);
and U14595 (N_14595,N_13370,N_12258);
xor U14596 (N_14596,N_13870,N_13253);
nor U14597 (N_14597,N_12060,N_13833);
xnor U14598 (N_14598,N_13214,N_12067);
xor U14599 (N_14599,N_12648,N_13004);
or U14600 (N_14600,N_13847,N_12808);
xor U14601 (N_14601,N_13009,N_12512);
nand U14602 (N_14602,N_12889,N_12667);
nor U14603 (N_14603,N_12797,N_13239);
nor U14604 (N_14604,N_12584,N_13638);
xnor U14605 (N_14605,N_13307,N_13415);
nand U14606 (N_14606,N_12915,N_12342);
xor U14607 (N_14607,N_13805,N_13825);
nand U14608 (N_14608,N_13361,N_12839);
nor U14609 (N_14609,N_13372,N_13102);
or U14610 (N_14610,N_12782,N_12690);
nand U14611 (N_14611,N_12001,N_13412);
or U14612 (N_14612,N_13181,N_13875);
nor U14613 (N_14613,N_12461,N_13767);
nand U14614 (N_14614,N_13072,N_13228);
and U14615 (N_14615,N_12400,N_13374);
or U14616 (N_14616,N_12635,N_12551);
or U14617 (N_14617,N_12058,N_12193);
and U14618 (N_14618,N_12641,N_12293);
nand U14619 (N_14619,N_13665,N_12039);
nor U14620 (N_14620,N_12780,N_12084);
or U14621 (N_14621,N_13408,N_13289);
nand U14622 (N_14622,N_12759,N_12367);
xor U14623 (N_14623,N_12221,N_13764);
or U14624 (N_14624,N_12850,N_12178);
xnor U14625 (N_14625,N_12942,N_13482);
or U14626 (N_14626,N_12793,N_13912);
or U14627 (N_14627,N_13693,N_12534);
nand U14628 (N_14628,N_12558,N_12550);
and U14629 (N_14629,N_13393,N_13258);
or U14630 (N_14630,N_12802,N_13984);
nor U14631 (N_14631,N_13386,N_13127);
xor U14632 (N_14632,N_13978,N_12983);
nor U14633 (N_14633,N_13462,N_12693);
nand U14634 (N_14634,N_13254,N_13479);
xor U14635 (N_14635,N_13544,N_12434);
nor U14636 (N_14636,N_13294,N_12206);
and U14637 (N_14637,N_13898,N_12925);
or U14638 (N_14638,N_12886,N_13300);
and U14639 (N_14639,N_13464,N_12991);
nand U14640 (N_14640,N_12993,N_13008);
and U14641 (N_14641,N_12527,N_12744);
nand U14642 (N_14642,N_12870,N_12924);
nand U14643 (N_14643,N_12417,N_13576);
nor U14644 (N_14644,N_12842,N_12788);
or U14645 (N_14645,N_13990,N_12510);
xnor U14646 (N_14646,N_13191,N_12885);
and U14647 (N_14647,N_13392,N_12175);
nand U14648 (N_14648,N_12980,N_13688);
xnor U14649 (N_14649,N_12149,N_12922);
nor U14650 (N_14650,N_13086,N_12172);
and U14651 (N_14651,N_13382,N_12382);
nor U14652 (N_14652,N_13927,N_12654);
or U14653 (N_14653,N_12098,N_13125);
and U14654 (N_14654,N_13993,N_12531);
or U14655 (N_14655,N_12318,N_12345);
xnor U14656 (N_14656,N_12918,N_13869);
nand U14657 (N_14657,N_12620,N_13426);
or U14658 (N_14658,N_12427,N_12362);
nand U14659 (N_14659,N_12970,N_12459);
or U14660 (N_14660,N_13905,N_12773);
and U14661 (N_14661,N_12486,N_13031);
nor U14662 (N_14662,N_13822,N_13617);
nor U14663 (N_14663,N_13695,N_13928);
or U14664 (N_14664,N_13118,N_12521);
xor U14665 (N_14665,N_13184,N_13570);
nand U14666 (N_14666,N_12872,N_12016);
nor U14667 (N_14667,N_13853,N_13773);
and U14668 (N_14668,N_13876,N_12235);
and U14669 (N_14669,N_12876,N_12226);
or U14670 (N_14670,N_13508,N_12329);
nand U14671 (N_14671,N_12518,N_13325);
nand U14672 (N_14672,N_13017,N_12203);
nand U14673 (N_14673,N_13293,N_13538);
and U14674 (N_14674,N_12837,N_12091);
and U14675 (N_14675,N_13851,N_12403);
nand U14676 (N_14676,N_13723,N_12637);
nand U14677 (N_14677,N_12652,N_12709);
or U14678 (N_14678,N_13134,N_12541);
or U14679 (N_14679,N_12503,N_12606);
or U14680 (N_14680,N_12554,N_12120);
nor U14681 (N_14681,N_13423,N_13108);
and U14682 (N_14682,N_12658,N_13712);
xnor U14683 (N_14683,N_13880,N_13733);
xor U14684 (N_14684,N_12390,N_13815);
nand U14685 (N_14685,N_13550,N_12573);
nand U14686 (N_14686,N_12812,N_12907);
nand U14687 (N_14687,N_13656,N_12302);
xnor U14688 (N_14688,N_13848,N_12913);
nor U14689 (N_14689,N_13037,N_12919);
or U14690 (N_14690,N_12613,N_13540);
nor U14691 (N_14691,N_13251,N_13867);
nand U14692 (N_14692,N_13648,N_13916);
and U14693 (N_14693,N_13384,N_13145);
and U14694 (N_14694,N_13681,N_13714);
or U14695 (N_14695,N_12234,N_12184);
or U14696 (N_14696,N_13204,N_12393);
and U14697 (N_14697,N_13346,N_12061);
or U14698 (N_14698,N_12989,N_12142);
and U14699 (N_14699,N_13226,N_13271);
or U14700 (N_14700,N_12079,N_13759);
xor U14701 (N_14701,N_13686,N_12282);
nor U14702 (N_14702,N_12858,N_13872);
nand U14703 (N_14703,N_12376,N_13400);
or U14704 (N_14704,N_12968,N_12657);
nand U14705 (N_14705,N_13602,N_13117);
nor U14706 (N_14706,N_13594,N_12941);
nor U14707 (N_14707,N_12107,N_12386);
or U14708 (N_14708,N_13924,N_12421);
xnor U14709 (N_14709,N_12241,N_13178);
nand U14710 (N_14710,N_12985,N_13212);
or U14711 (N_14711,N_13735,N_13485);
or U14712 (N_14712,N_13466,N_12383);
nand U14713 (N_14713,N_12861,N_13836);
xor U14714 (N_14714,N_12931,N_13784);
or U14715 (N_14715,N_12524,N_13348);
or U14716 (N_14716,N_12083,N_13757);
and U14717 (N_14717,N_12085,N_12154);
or U14718 (N_14718,N_12943,N_12697);
nor U14719 (N_14719,N_12629,N_13509);
nor U14720 (N_14720,N_12947,N_12694);
nor U14721 (N_14721,N_12854,N_13790);
and U14722 (N_14722,N_12649,N_13457);
xnor U14723 (N_14723,N_13418,N_13162);
xnor U14724 (N_14724,N_12607,N_12954);
nand U14725 (N_14725,N_13855,N_13238);
xnor U14726 (N_14726,N_13979,N_13327);
nand U14727 (N_14727,N_12224,N_12844);
nand U14728 (N_14728,N_13988,N_12495);
xnor U14729 (N_14729,N_12339,N_12994);
nor U14730 (N_14730,N_13116,N_13297);
nor U14731 (N_14731,N_13895,N_13368);
and U14732 (N_14732,N_12686,N_13156);
and U14733 (N_14733,N_13637,N_13672);
xor U14734 (N_14734,N_12545,N_12212);
or U14735 (N_14735,N_12937,N_13196);
and U14736 (N_14736,N_13168,N_12399);
nor U14737 (N_14737,N_12140,N_13873);
xor U14738 (N_14738,N_12109,N_12305);
and U14739 (N_14739,N_13704,N_13158);
nor U14740 (N_14740,N_12996,N_13385);
or U14741 (N_14741,N_12926,N_13618);
xor U14742 (N_14742,N_13313,N_13473);
and U14743 (N_14743,N_13496,N_12781);
and U14744 (N_14744,N_13078,N_12144);
and U14745 (N_14745,N_12930,N_13449);
or U14746 (N_14746,N_13195,N_12022);
or U14747 (N_14747,N_12295,N_12677);
and U14748 (N_14748,N_12191,N_13429);
nand U14749 (N_14749,N_12571,N_12387);
or U14750 (N_14750,N_12843,N_12514);
and U14751 (N_14751,N_12824,N_12969);
and U14752 (N_14752,N_13802,N_13038);
and U14753 (N_14753,N_13977,N_13441);
xor U14754 (N_14754,N_12075,N_12897);
and U14755 (N_14755,N_12984,N_13839);
xor U14756 (N_14756,N_12564,N_13739);
or U14757 (N_14757,N_13234,N_13920);
nand U14758 (N_14758,N_13421,N_13826);
or U14759 (N_14759,N_13082,N_12619);
and U14760 (N_14760,N_13398,N_13317);
xor U14761 (N_14761,N_12304,N_12283);
nor U14762 (N_14762,N_13265,N_13098);
nand U14763 (N_14763,N_13843,N_12945);
xnor U14764 (N_14764,N_13878,N_13101);
xnor U14765 (N_14765,N_13132,N_12070);
xor U14766 (N_14766,N_13391,N_12307);
and U14767 (N_14767,N_13229,N_13734);
nand U14768 (N_14768,N_13138,N_13001);
and U14769 (N_14769,N_13281,N_13044);
and U14770 (N_14770,N_13137,N_13682);
and U14771 (N_14771,N_13514,N_12042);
nand U14772 (N_14772,N_12646,N_13174);
xnor U14773 (N_14773,N_12501,N_12256);
nor U14774 (N_14774,N_12087,N_12821);
nor U14775 (N_14775,N_13584,N_12823);
and U14776 (N_14776,N_13600,N_13151);
and U14777 (N_14777,N_12575,N_12207);
and U14778 (N_14778,N_13713,N_13794);
nand U14779 (N_14779,N_12528,N_12783);
nor U14780 (N_14780,N_13074,N_12663);
or U14781 (N_14781,N_13139,N_12700);
and U14782 (N_14782,N_12096,N_13111);
or U14783 (N_14783,N_13583,N_13359);
or U14784 (N_14784,N_12784,N_13772);
xor U14785 (N_14785,N_13892,N_13446);
xnor U14786 (N_14786,N_12939,N_13527);
nor U14787 (N_14787,N_12660,N_12873);
nor U14788 (N_14788,N_13194,N_12034);
and U14789 (N_14789,N_13305,N_13144);
nor U14790 (N_14790,N_12794,N_12525);
and U14791 (N_14791,N_13287,N_13692);
or U14792 (N_14792,N_12874,N_12766);
nand U14793 (N_14793,N_12186,N_12357);
nor U14794 (N_14794,N_12372,N_12901);
xnor U14795 (N_14795,N_13560,N_13055);
nand U14796 (N_14796,N_12111,N_12805);
or U14797 (N_14797,N_12745,N_13800);
or U14798 (N_14798,N_13436,N_12008);
and U14799 (N_14799,N_12265,N_13748);
or U14800 (N_14800,N_13623,N_12914);
and U14801 (N_14801,N_13838,N_12401);
nand U14802 (N_14802,N_12715,N_13698);
xnor U14803 (N_14803,N_12779,N_13552);
and U14804 (N_14804,N_12582,N_13267);
nor U14805 (N_14805,N_13789,N_13974);
or U14806 (N_14806,N_13395,N_13342);
nand U14807 (N_14807,N_12849,N_12846);
nor U14808 (N_14808,N_13472,N_12338);
nor U14809 (N_14809,N_12975,N_12252);
or U14810 (N_14810,N_12116,N_12003);
or U14811 (N_14811,N_12378,N_13279);
and U14812 (N_14812,N_12054,N_13375);
nor U14813 (N_14813,N_12465,N_12312);
xor U14814 (N_14814,N_12169,N_13674);
and U14815 (N_14815,N_12865,N_13105);
and U14816 (N_14816,N_13727,N_12392);
xor U14817 (N_14817,N_12010,N_12814);
or U14818 (N_14818,N_12218,N_12397);
nor U14819 (N_14819,N_12927,N_13955);
nand U14820 (N_14820,N_13420,N_13841);
or U14821 (N_14821,N_13164,N_12267);
nor U14822 (N_14822,N_12108,N_12050);
nand U14823 (N_14823,N_12133,N_12477);
nand U14824 (N_14824,N_12529,N_13680);
nand U14825 (N_14825,N_12621,N_13647);
nand U14826 (N_14826,N_12099,N_12330);
nand U14827 (N_14827,N_13428,N_13034);
xor U14828 (N_14828,N_13797,N_12998);
nand U14829 (N_14829,N_13795,N_12196);
nor U14830 (N_14830,N_12410,N_12608);
xor U14831 (N_14831,N_13651,N_13950);
nand U14832 (N_14832,N_13556,N_13435);
nand U14833 (N_14833,N_12062,N_12929);
and U14834 (N_14834,N_13944,N_13272);
or U14835 (N_14835,N_12871,N_13128);
xnor U14836 (N_14836,N_12315,N_12882);
and U14837 (N_14837,N_12639,N_12695);
and U14838 (N_14838,N_13216,N_12614);
nor U14839 (N_14839,N_13707,N_13555);
and U14840 (N_14840,N_13075,N_13383);
or U14841 (N_14841,N_12711,N_13909);
or U14842 (N_14842,N_12408,N_13813);
nor U14843 (N_14843,N_13513,N_13953);
nand U14844 (N_14844,N_13701,N_13381);
xnor U14845 (N_14845,N_13754,N_12139);
nand U14846 (N_14846,N_13921,N_13495);
and U14847 (N_14847,N_13321,N_13811);
or U14848 (N_14848,N_12685,N_13166);
nor U14849 (N_14849,N_13644,N_13135);
or U14850 (N_14850,N_13621,N_13442);
or U14851 (N_14851,N_12347,N_13177);
or U14852 (N_14852,N_13528,N_13738);
xnor U14853 (N_14853,N_13913,N_13689);
xor U14854 (N_14854,N_13014,N_12118);
nand U14855 (N_14855,N_12165,N_12624);
nand U14856 (N_14856,N_13750,N_13334);
and U14857 (N_14857,N_12504,N_13981);
or U14858 (N_14858,N_12598,N_13465);
xnor U14859 (N_14859,N_12227,N_13614);
nand U14860 (N_14860,N_13866,N_12273);
nor U14861 (N_14861,N_12441,N_13879);
nand U14862 (N_14862,N_13715,N_12123);
nand U14863 (N_14863,N_12174,N_12242);
nor U14864 (N_14864,N_12819,N_13013);
or U14865 (N_14865,N_12469,N_13399);
xor U14866 (N_14866,N_13475,N_13737);
nor U14867 (N_14867,N_12863,N_12288);
xnor U14868 (N_14868,N_12492,N_13176);
xor U14869 (N_14869,N_12365,N_13456);
and U14870 (N_14870,N_12616,N_12775);
nor U14871 (N_14871,N_12934,N_13288);
xnor U14872 (N_14872,N_12864,N_12618);
nand U14873 (N_14873,N_13182,N_13844);
nor U14874 (N_14874,N_12946,N_13448);
xnor U14875 (N_14875,N_12900,N_12033);
xnor U14876 (N_14876,N_12755,N_13691);
nor U14877 (N_14877,N_12433,N_13308);
or U14878 (N_14878,N_12088,N_13629);
nand U14879 (N_14879,N_13543,N_13332);
nand U14880 (N_14880,N_12044,N_13945);
xnor U14881 (N_14881,N_12817,N_12431);
xor U14882 (N_14882,N_12845,N_12728);
and U14883 (N_14883,N_13515,N_13854);
nor U14884 (N_14884,N_13780,N_12151);
nor U14885 (N_14885,N_12432,N_12656);
and U14886 (N_14886,N_12565,N_12832);
nor U14887 (N_14887,N_13041,N_12509);
and U14888 (N_14888,N_12090,N_13414);
xor U14889 (N_14889,N_12496,N_13206);
or U14890 (N_14890,N_13076,N_13291);
nor U14891 (N_14891,N_12214,N_13846);
nand U14892 (N_14892,N_13831,N_12286);
and U14893 (N_14893,N_13474,N_13282);
nor U14894 (N_14894,N_13747,N_12696);
xnor U14895 (N_14895,N_13699,N_12683);
xor U14896 (N_14896,N_13278,N_12944);
xor U14897 (N_14897,N_13266,N_13827);
nand U14898 (N_14898,N_12699,N_13235);
and U14899 (N_14899,N_13874,N_12898);
xnor U14900 (N_14900,N_13694,N_12052);
and U14901 (N_14901,N_12220,N_13056);
xnor U14902 (N_14902,N_12290,N_13344);
xor U14903 (N_14903,N_13850,N_12932);
nor U14904 (N_14904,N_12413,N_12328);
nor U14905 (N_14905,N_13809,N_13631);
xor U14906 (N_14906,N_13724,N_13902);
xnor U14907 (N_14907,N_12200,N_12768);
and U14908 (N_14908,N_13244,N_12233);
or U14909 (N_14909,N_13364,N_13403);
and U14910 (N_14910,N_12625,N_13231);
xnor U14911 (N_14911,N_12520,N_13983);
and U14912 (N_14912,N_13079,N_13659);
or U14913 (N_14913,N_13619,N_12548);
xor U14914 (N_14914,N_12359,N_13124);
nor U14915 (N_14915,N_13512,N_13380);
and U14916 (N_14916,N_13269,N_13986);
xor U14917 (N_14917,N_13366,N_12811);
nand U14918 (N_14918,N_13796,N_12134);
nand U14919 (N_14919,N_12841,N_12310);
nor U14920 (N_14920,N_13582,N_12210);
and U14921 (N_14921,N_12306,N_12095);
and U14922 (N_14922,N_13642,N_13643);
nor U14923 (N_14923,N_12597,N_12080);
and U14924 (N_14924,N_12701,N_12270);
nand U14925 (N_14925,N_12615,N_13100);
nor U14926 (N_14926,N_13402,N_13591);
nor U14927 (N_14927,N_13455,N_12570);
nand U14928 (N_14928,N_12892,N_13877);
nand U14929 (N_14929,N_12555,N_13975);
xor U14930 (N_14930,N_12478,N_12592);
xor U14931 (N_14931,N_12266,N_12300);
nand U14932 (N_14932,N_12319,N_13660);
or U14933 (N_14933,N_12458,N_13779);
or U14934 (N_14934,N_13700,N_13161);
or U14935 (N_14935,N_12912,N_13702);
and U14936 (N_14936,N_13940,N_13173);
and U14937 (N_14937,N_12030,N_13460);
or U14938 (N_14938,N_12000,N_13369);
xor U14939 (N_14939,N_12462,N_13489);
and U14940 (N_14940,N_12303,N_12285);
nand U14941 (N_14941,N_13476,N_13837);
and U14942 (N_14942,N_13341,N_12281);
nand U14943 (N_14943,N_12644,N_13264);
nand U14944 (N_14944,N_12029,N_13468);
nand U14945 (N_14945,N_13080,N_12190);
nor U14946 (N_14946,N_12130,N_12511);
xor U14947 (N_14947,N_12567,N_13926);
nand U14948 (N_14948,N_13992,N_12348);
xor U14949 (N_14949,N_13087,N_13406);
nor U14950 (N_14950,N_13574,N_13270);
nand U14951 (N_14951,N_13459,N_12104);
nor U14952 (N_14952,N_13071,N_13939);
nand U14953 (N_14953,N_12488,N_12796);
nor U14954 (N_14954,N_13352,N_12853);
nor U14955 (N_14955,N_13189,N_12966);
or U14956 (N_14956,N_12708,N_12502);
nor U14957 (N_14957,N_13486,N_12445);
nand U14958 (N_14958,N_13835,N_12141);
xnor U14959 (N_14959,N_13083,N_13247);
or U14960 (N_14960,N_12856,N_13094);
nor U14961 (N_14961,N_12147,N_13901);
nor U14962 (N_14962,N_13355,N_13632);
or U14963 (N_14963,N_12909,N_13803);
xor U14964 (N_14964,N_12023,N_13761);
and U14965 (N_14965,N_13788,N_12798);
or U14966 (N_14966,N_13500,N_12394);
nor U14967 (N_14967,N_13043,N_13096);
xor U14968 (N_14968,N_12815,N_12124);
and U14969 (N_14969,N_13498,N_12074);
nand U14970 (N_14970,N_13771,N_12645);
nor U14971 (N_14971,N_13952,N_12908);
nand U14972 (N_14972,N_12756,N_12883);
or U14973 (N_14973,N_12538,N_13834);
xnor U14974 (N_14974,N_12453,N_13404);
or U14975 (N_14975,N_12291,N_13947);
and U14976 (N_14976,N_12778,N_12585);
or U14977 (N_14977,N_13506,N_12640);
or U14978 (N_14978,N_13740,N_13256);
xnor U14979 (N_14979,N_13440,N_13507);
nand U14980 (N_14980,N_13938,N_13536);
and U14981 (N_14981,N_13765,N_13610);
and U14982 (N_14982,N_12158,N_12505);
or U14983 (N_14983,N_12508,N_12127);
or U14984 (N_14984,N_12960,N_12603);
xor U14985 (N_14985,N_13971,N_13221);
and U14986 (N_14986,N_13190,N_13215);
or U14987 (N_14987,N_12356,N_13129);
and U14988 (N_14988,N_13774,N_12650);
or U14989 (N_14989,N_12785,N_13203);
nand U14990 (N_14990,N_13255,N_13343);
nand U14991 (N_14991,N_13048,N_13683);
nor U14992 (N_14992,N_12877,N_12046);
nor U14993 (N_14993,N_12589,N_12480);
nand U14994 (N_14994,N_12724,N_12604);
xnor U14995 (N_14995,N_13470,N_12680);
and U14996 (N_14996,N_13786,N_13845);
xnor U14997 (N_14997,N_13200,N_13760);
xnor U14998 (N_14998,N_12475,N_12183);
nor U14999 (N_14999,N_12380,N_12933);
and U15000 (N_15000,N_12647,N_13800);
or U15001 (N_15001,N_12364,N_12376);
xor U15002 (N_15002,N_13203,N_12660);
or U15003 (N_15003,N_13243,N_12501);
or U15004 (N_15004,N_12286,N_12167);
or U15005 (N_15005,N_12764,N_12223);
nand U15006 (N_15006,N_13457,N_12071);
nand U15007 (N_15007,N_12308,N_13818);
xnor U15008 (N_15008,N_12366,N_12659);
nor U15009 (N_15009,N_13182,N_12171);
xor U15010 (N_15010,N_12572,N_12005);
xor U15011 (N_15011,N_13667,N_12445);
nand U15012 (N_15012,N_13952,N_13128);
nor U15013 (N_15013,N_12816,N_12691);
xnor U15014 (N_15014,N_13555,N_12944);
xnor U15015 (N_15015,N_12660,N_12036);
nand U15016 (N_15016,N_12235,N_12657);
nand U15017 (N_15017,N_13908,N_12024);
and U15018 (N_15018,N_13105,N_13870);
nand U15019 (N_15019,N_13783,N_13206);
nand U15020 (N_15020,N_12570,N_13585);
and U15021 (N_15021,N_12518,N_13709);
nor U15022 (N_15022,N_12047,N_12854);
and U15023 (N_15023,N_12510,N_13288);
nand U15024 (N_15024,N_13530,N_12015);
nor U15025 (N_15025,N_12082,N_13276);
nand U15026 (N_15026,N_12111,N_12469);
or U15027 (N_15027,N_13090,N_12662);
nand U15028 (N_15028,N_13161,N_13280);
xnor U15029 (N_15029,N_12901,N_12792);
xnor U15030 (N_15030,N_13558,N_12146);
xor U15031 (N_15031,N_12230,N_13433);
or U15032 (N_15032,N_13735,N_13767);
or U15033 (N_15033,N_12675,N_13597);
or U15034 (N_15034,N_12681,N_13337);
nor U15035 (N_15035,N_13747,N_13893);
or U15036 (N_15036,N_13053,N_12784);
nand U15037 (N_15037,N_13881,N_12385);
xor U15038 (N_15038,N_13169,N_13378);
xor U15039 (N_15039,N_13064,N_13301);
or U15040 (N_15040,N_13467,N_13287);
or U15041 (N_15041,N_12781,N_13844);
and U15042 (N_15042,N_12126,N_12223);
and U15043 (N_15043,N_12343,N_13907);
or U15044 (N_15044,N_12741,N_12242);
nand U15045 (N_15045,N_13200,N_12945);
xnor U15046 (N_15046,N_13120,N_13179);
or U15047 (N_15047,N_12624,N_13374);
or U15048 (N_15048,N_12419,N_12463);
or U15049 (N_15049,N_13884,N_13253);
and U15050 (N_15050,N_13676,N_12825);
and U15051 (N_15051,N_12099,N_12838);
or U15052 (N_15052,N_13155,N_12200);
or U15053 (N_15053,N_13079,N_13551);
nor U15054 (N_15054,N_12291,N_12162);
xor U15055 (N_15055,N_13378,N_13104);
nand U15056 (N_15056,N_12224,N_13965);
xnor U15057 (N_15057,N_13687,N_13677);
nand U15058 (N_15058,N_12805,N_12786);
nand U15059 (N_15059,N_13195,N_13555);
or U15060 (N_15060,N_12107,N_13233);
and U15061 (N_15061,N_12773,N_12403);
nor U15062 (N_15062,N_13201,N_13737);
nand U15063 (N_15063,N_13790,N_12050);
nor U15064 (N_15064,N_13513,N_12575);
nand U15065 (N_15065,N_12213,N_13653);
or U15066 (N_15066,N_13015,N_12556);
and U15067 (N_15067,N_13517,N_12753);
or U15068 (N_15068,N_13796,N_12509);
or U15069 (N_15069,N_12896,N_13968);
xnor U15070 (N_15070,N_13209,N_12861);
and U15071 (N_15071,N_12239,N_12078);
nor U15072 (N_15072,N_13851,N_13064);
nor U15073 (N_15073,N_12024,N_13741);
and U15074 (N_15074,N_12480,N_12642);
nand U15075 (N_15075,N_13811,N_13249);
or U15076 (N_15076,N_13357,N_12086);
nand U15077 (N_15077,N_12420,N_13859);
xnor U15078 (N_15078,N_13703,N_12863);
nor U15079 (N_15079,N_12037,N_12500);
and U15080 (N_15080,N_13997,N_12437);
or U15081 (N_15081,N_12478,N_12685);
or U15082 (N_15082,N_12829,N_13952);
or U15083 (N_15083,N_13446,N_12448);
and U15084 (N_15084,N_13610,N_13013);
nor U15085 (N_15085,N_12794,N_13052);
and U15086 (N_15086,N_13973,N_12150);
or U15087 (N_15087,N_12579,N_12028);
or U15088 (N_15088,N_13170,N_13861);
nor U15089 (N_15089,N_13241,N_12930);
nor U15090 (N_15090,N_13308,N_12390);
and U15091 (N_15091,N_13724,N_13310);
nand U15092 (N_15092,N_13402,N_13242);
and U15093 (N_15093,N_12686,N_13187);
nor U15094 (N_15094,N_13761,N_13726);
and U15095 (N_15095,N_12742,N_12041);
or U15096 (N_15096,N_13665,N_13413);
nand U15097 (N_15097,N_12573,N_13257);
or U15098 (N_15098,N_13922,N_12754);
or U15099 (N_15099,N_13195,N_12971);
xnor U15100 (N_15100,N_13425,N_12692);
nor U15101 (N_15101,N_13652,N_12157);
or U15102 (N_15102,N_12419,N_13989);
nand U15103 (N_15103,N_13435,N_12284);
and U15104 (N_15104,N_12592,N_12647);
nand U15105 (N_15105,N_13575,N_12943);
nand U15106 (N_15106,N_12852,N_13379);
nand U15107 (N_15107,N_13960,N_12859);
and U15108 (N_15108,N_12053,N_13752);
and U15109 (N_15109,N_13563,N_13843);
xnor U15110 (N_15110,N_13910,N_13879);
nand U15111 (N_15111,N_12411,N_13528);
nand U15112 (N_15112,N_13802,N_12281);
and U15113 (N_15113,N_13759,N_13907);
nand U15114 (N_15114,N_12164,N_12484);
nand U15115 (N_15115,N_13224,N_13984);
or U15116 (N_15116,N_12044,N_13371);
xor U15117 (N_15117,N_13991,N_13976);
xor U15118 (N_15118,N_12892,N_13614);
or U15119 (N_15119,N_12089,N_12496);
or U15120 (N_15120,N_13175,N_12565);
and U15121 (N_15121,N_13738,N_13307);
or U15122 (N_15122,N_12459,N_13860);
nor U15123 (N_15123,N_12196,N_13379);
xor U15124 (N_15124,N_13451,N_13494);
nor U15125 (N_15125,N_13148,N_13364);
or U15126 (N_15126,N_13539,N_13686);
xnor U15127 (N_15127,N_13906,N_13174);
nand U15128 (N_15128,N_12516,N_13318);
xnor U15129 (N_15129,N_12139,N_13280);
or U15130 (N_15130,N_13574,N_13982);
nor U15131 (N_15131,N_12170,N_12348);
and U15132 (N_15132,N_12031,N_12962);
and U15133 (N_15133,N_13202,N_12023);
xor U15134 (N_15134,N_12927,N_13278);
xor U15135 (N_15135,N_12338,N_12309);
nand U15136 (N_15136,N_13138,N_13788);
or U15137 (N_15137,N_13235,N_13773);
xnor U15138 (N_15138,N_13800,N_12088);
or U15139 (N_15139,N_12863,N_12678);
nand U15140 (N_15140,N_13757,N_12528);
and U15141 (N_15141,N_12521,N_12837);
nor U15142 (N_15142,N_13722,N_13274);
nand U15143 (N_15143,N_12927,N_13972);
xor U15144 (N_15144,N_12951,N_13037);
xor U15145 (N_15145,N_13745,N_13585);
and U15146 (N_15146,N_13956,N_12924);
nand U15147 (N_15147,N_13143,N_13111);
or U15148 (N_15148,N_13094,N_12446);
and U15149 (N_15149,N_12221,N_13662);
or U15150 (N_15150,N_12260,N_13474);
nand U15151 (N_15151,N_12021,N_12484);
or U15152 (N_15152,N_13324,N_13691);
and U15153 (N_15153,N_12323,N_13215);
nor U15154 (N_15154,N_13730,N_12966);
and U15155 (N_15155,N_12913,N_12302);
xor U15156 (N_15156,N_12574,N_12214);
nor U15157 (N_15157,N_13552,N_13143);
xor U15158 (N_15158,N_13441,N_13611);
or U15159 (N_15159,N_13594,N_12410);
nand U15160 (N_15160,N_13861,N_12938);
and U15161 (N_15161,N_13523,N_12548);
nor U15162 (N_15162,N_12577,N_12070);
xnor U15163 (N_15163,N_13958,N_13305);
or U15164 (N_15164,N_13815,N_12891);
xor U15165 (N_15165,N_13480,N_12216);
nor U15166 (N_15166,N_12440,N_13363);
nor U15167 (N_15167,N_13815,N_13875);
xor U15168 (N_15168,N_13512,N_12096);
nand U15169 (N_15169,N_13444,N_13560);
xor U15170 (N_15170,N_12373,N_12049);
or U15171 (N_15171,N_13942,N_12295);
or U15172 (N_15172,N_13459,N_13427);
or U15173 (N_15173,N_13849,N_13854);
and U15174 (N_15174,N_13980,N_12146);
nor U15175 (N_15175,N_13182,N_12873);
or U15176 (N_15176,N_13329,N_12152);
and U15177 (N_15177,N_13447,N_13441);
or U15178 (N_15178,N_13173,N_13422);
nor U15179 (N_15179,N_13243,N_12085);
and U15180 (N_15180,N_13129,N_12881);
xor U15181 (N_15181,N_12567,N_12213);
or U15182 (N_15182,N_13847,N_12443);
nor U15183 (N_15183,N_12407,N_13754);
nor U15184 (N_15184,N_12603,N_12228);
or U15185 (N_15185,N_12514,N_12434);
and U15186 (N_15186,N_13390,N_13310);
and U15187 (N_15187,N_12380,N_13734);
xnor U15188 (N_15188,N_12514,N_13785);
or U15189 (N_15189,N_13218,N_12653);
nor U15190 (N_15190,N_13820,N_13913);
or U15191 (N_15191,N_13018,N_12839);
nand U15192 (N_15192,N_12021,N_12472);
nor U15193 (N_15193,N_12854,N_13425);
nor U15194 (N_15194,N_13039,N_12902);
xnor U15195 (N_15195,N_13615,N_12452);
xnor U15196 (N_15196,N_12190,N_13374);
and U15197 (N_15197,N_13902,N_12153);
xor U15198 (N_15198,N_12275,N_12964);
xnor U15199 (N_15199,N_12209,N_12640);
nand U15200 (N_15200,N_13958,N_13451);
xor U15201 (N_15201,N_12820,N_12159);
nand U15202 (N_15202,N_13871,N_12021);
xnor U15203 (N_15203,N_12744,N_12889);
nand U15204 (N_15204,N_12248,N_12236);
xnor U15205 (N_15205,N_12635,N_13603);
nor U15206 (N_15206,N_13472,N_13877);
nor U15207 (N_15207,N_12040,N_13227);
and U15208 (N_15208,N_12113,N_12538);
xor U15209 (N_15209,N_13753,N_12725);
xor U15210 (N_15210,N_13676,N_12920);
nor U15211 (N_15211,N_13666,N_13446);
nand U15212 (N_15212,N_13042,N_12838);
xnor U15213 (N_15213,N_12967,N_12724);
or U15214 (N_15214,N_12474,N_12125);
xnor U15215 (N_15215,N_13570,N_13473);
nor U15216 (N_15216,N_12043,N_12126);
and U15217 (N_15217,N_13904,N_12472);
or U15218 (N_15218,N_13847,N_13079);
xor U15219 (N_15219,N_13721,N_12841);
nor U15220 (N_15220,N_13243,N_12239);
nand U15221 (N_15221,N_12691,N_12175);
nand U15222 (N_15222,N_12749,N_13748);
nor U15223 (N_15223,N_12322,N_13028);
nand U15224 (N_15224,N_12576,N_13760);
or U15225 (N_15225,N_13043,N_13177);
xnor U15226 (N_15226,N_13270,N_13305);
nand U15227 (N_15227,N_13800,N_12830);
xnor U15228 (N_15228,N_13540,N_12488);
nor U15229 (N_15229,N_13755,N_13328);
xnor U15230 (N_15230,N_12456,N_12200);
xnor U15231 (N_15231,N_12813,N_12795);
nand U15232 (N_15232,N_13212,N_12617);
nor U15233 (N_15233,N_12064,N_13162);
nand U15234 (N_15234,N_12350,N_13861);
nand U15235 (N_15235,N_13030,N_12108);
nand U15236 (N_15236,N_12544,N_12533);
nand U15237 (N_15237,N_13140,N_12939);
and U15238 (N_15238,N_12231,N_13750);
nand U15239 (N_15239,N_13016,N_13095);
or U15240 (N_15240,N_12645,N_13492);
nand U15241 (N_15241,N_12539,N_12993);
or U15242 (N_15242,N_12718,N_13679);
xor U15243 (N_15243,N_13100,N_12812);
nand U15244 (N_15244,N_13194,N_12481);
xor U15245 (N_15245,N_12215,N_12717);
or U15246 (N_15246,N_12044,N_13497);
or U15247 (N_15247,N_13244,N_13166);
and U15248 (N_15248,N_13998,N_13393);
nand U15249 (N_15249,N_13257,N_12880);
nor U15250 (N_15250,N_13101,N_13822);
xor U15251 (N_15251,N_13974,N_12192);
xor U15252 (N_15252,N_12023,N_12893);
nor U15253 (N_15253,N_13512,N_13992);
xnor U15254 (N_15254,N_12048,N_13727);
nand U15255 (N_15255,N_13889,N_13017);
nand U15256 (N_15256,N_12451,N_13522);
or U15257 (N_15257,N_12184,N_13130);
nor U15258 (N_15258,N_12305,N_12712);
or U15259 (N_15259,N_13395,N_12112);
or U15260 (N_15260,N_12886,N_13663);
or U15261 (N_15261,N_13460,N_13843);
nand U15262 (N_15262,N_13423,N_12801);
or U15263 (N_15263,N_12612,N_12359);
nor U15264 (N_15264,N_12128,N_13940);
or U15265 (N_15265,N_12613,N_13464);
and U15266 (N_15266,N_13392,N_13544);
nor U15267 (N_15267,N_13045,N_13112);
nor U15268 (N_15268,N_13390,N_13473);
xnor U15269 (N_15269,N_12544,N_13402);
and U15270 (N_15270,N_12734,N_12998);
xnor U15271 (N_15271,N_12985,N_13228);
and U15272 (N_15272,N_13085,N_13762);
xor U15273 (N_15273,N_12928,N_12788);
xor U15274 (N_15274,N_13747,N_12454);
xnor U15275 (N_15275,N_12603,N_12249);
or U15276 (N_15276,N_12232,N_12605);
nand U15277 (N_15277,N_13638,N_13890);
nand U15278 (N_15278,N_13118,N_13505);
nand U15279 (N_15279,N_12675,N_13701);
nand U15280 (N_15280,N_12969,N_13700);
xnor U15281 (N_15281,N_13534,N_12952);
or U15282 (N_15282,N_12116,N_13128);
and U15283 (N_15283,N_12410,N_13700);
nor U15284 (N_15284,N_13636,N_12364);
and U15285 (N_15285,N_13890,N_13221);
nor U15286 (N_15286,N_12334,N_12867);
xor U15287 (N_15287,N_12658,N_12762);
nor U15288 (N_15288,N_13884,N_12635);
nor U15289 (N_15289,N_12589,N_12841);
nor U15290 (N_15290,N_12073,N_12511);
or U15291 (N_15291,N_13680,N_13851);
nand U15292 (N_15292,N_12712,N_13467);
nand U15293 (N_15293,N_13019,N_13423);
and U15294 (N_15294,N_13775,N_13587);
and U15295 (N_15295,N_12413,N_12854);
or U15296 (N_15296,N_13226,N_12279);
xnor U15297 (N_15297,N_13156,N_12452);
or U15298 (N_15298,N_13773,N_12644);
xnor U15299 (N_15299,N_12424,N_12303);
or U15300 (N_15300,N_12679,N_12254);
and U15301 (N_15301,N_12283,N_12882);
xnor U15302 (N_15302,N_13199,N_13303);
nor U15303 (N_15303,N_13406,N_12692);
xor U15304 (N_15304,N_12267,N_12628);
and U15305 (N_15305,N_13235,N_12547);
nor U15306 (N_15306,N_13151,N_12676);
nor U15307 (N_15307,N_13720,N_13011);
xnor U15308 (N_15308,N_12463,N_12641);
and U15309 (N_15309,N_12843,N_12039);
xor U15310 (N_15310,N_12092,N_12469);
nand U15311 (N_15311,N_13628,N_13663);
nor U15312 (N_15312,N_13914,N_13460);
or U15313 (N_15313,N_13530,N_13208);
xnor U15314 (N_15314,N_13666,N_12645);
xor U15315 (N_15315,N_13257,N_12588);
nand U15316 (N_15316,N_13268,N_12997);
nand U15317 (N_15317,N_12209,N_13498);
nand U15318 (N_15318,N_13140,N_13552);
xor U15319 (N_15319,N_12293,N_12407);
and U15320 (N_15320,N_12515,N_13993);
and U15321 (N_15321,N_12232,N_12350);
and U15322 (N_15322,N_12376,N_13450);
and U15323 (N_15323,N_12641,N_13010);
xnor U15324 (N_15324,N_12118,N_12783);
and U15325 (N_15325,N_13418,N_12270);
or U15326 (N_15326,N_12201,N_13605);
and U15327 (N_15327,N_13625,N_13964);
nor U15328 (N_15328,N_13853,N_13983);
or U15329 (N_15329,N_12106,N_13384);
nand U15330 (N_15330,N_12312,N_12142);
nand U15331 (N_15331,N_12107,N_13943);
and U15332 (N_15332,N_13877,N_13241);
nand U15333 (N_15333,N_12032,N_12538);
xnor U15334 (N_15334,N_13226,N_12926);
and U15335 (N_15335,N_12938,N_13539);
nor U15336 (N_15336,N_12697,N_13340);
nor U15337 (N_15337,N_12716,N_12259);
xnor U15338 (N_15338,N_12079,N_12113);
nand U15339 (N_15339,N_12885,N_13587);
nand U15340 (N_15340,N_13462,N_12002);
xor U15341 (N_15341,N_13209,N_13341);
nand U15342 (N_15342,N_13197,N_12378);
nand U15343 (N_15343,N_12688,N_12135);
or U15344 (N_15344,N_13922,N_12799);
and U15345 (N_15345,N_12990,N_13958);
nor U15346 (N_15346,N_13679,N_12543);
or U15347 (N_15347,N_12672,N_13835);
or U15348 (N_15348,N_12660,N_12025);
nand U15349 (N_15349,N_12298,N_13529);
nor U15350 (N_15350,N_12111,N_12317);
xor U15351 (N_15351,N_12956,N_12961);
nor U15352 (N_15352,N_13308,N_13010);
and U15353 (N_15353,N_12309,N_12114);
xor U15354 (N_15354,N_13340,N_12038);
nand U15355 (N_15355,N_13710,N_13963);
or U15356 (N_15356,N_13314,N_12794);
nand U15357 (N_15357,N_12376,N_12403);
nand U15358 (N_15358,N_12775,N_12389);
or U15359 (N_15359,N_13666,N_13431);
xnor U15360 (N_15360,N_12894,N_12244);
and U15361 (N_15361,N_12679,N_12245);
and U15362 (N_15362,N_13146,N_12457);
xor U15363 (N_15363,N_13733,N_13757);
xnor U15364 (N_15364,N_13419,N_12038);
and U15365 (N_15365,N_12503,N_13120);
xor U15366 (N_15366,N_13715,N_12736);
nor U15367 (N_15367,N_13289,N_12907);
nand U15368 (N_15368,N_12139,N_12574);
xor U15369 (N_15369,N_13137,N_13605);
nand U15370 (N_15370,N_13348,N_12316);
nor U15371 (N_15371,N_12232,N_12751);
nor U15372 (N_15372,N_13932,N_13970);
or U15373 (N_15373,N_12262,N_12323);
xor U15374 (N_15374,N_13727,N_13137);
and U15375 (N_15375,N_12311,N_13843);
or U15376 (N_15376,N_12265,N_12628);
xnor U15377 (N_15377,N_12759,N_12001);
nand U15378 (N_15378,N_12225,N_12034);
and U15379 (N_15379,N_12658,N_12157);
xor U15380 (N_15380,N_12704,N_12805);
or U15381 (N_15381,N_13483,N_13253);
nand U15382 (N_15382,N_12564,N_13867);
and U15383 (N_15383,N_12340,N_13573);
nand U15384 (N_15384,N_12279,N_12587);
and U15385 (N_15385,N_13742,N_12925);
and U15386 (N_15386,N_12639,N_13698);
and U15387 (N_15387,N_13390,N_12821);
nand U15388 (N_15388,N_12478,N_13474);
xnor U15389 (N_15389,N_13527,N_12879);
xor U15390 (N_15390,N_13021,N_12397);
or U15391 (N_15391,N_13535,N_13922);
nand U15392 (N_15392,N_12371,N_12194);
nor U15393 (N_15393,N_12164,N_13947);
or U15394 (N_15394,N_12741,N_12726);
or U15395 (N_15395,N_13931,N_12565);
nand U15396 (N_15396,N_12366,N_12073);
nor U15397 (N_15397,N_13191,N_12840);
and U15398 (N_15398,N_12099,N_12334);
nor U15399 (N_15399,N_13637,N_13410);
xnor U15400 (N_15400,N_13934,N_12447);
and U15401 (N_15401,N_13945,N_12878);
and U15402 (N_15402,N_13292,N_13102);
nor U15403 (N_15403,N_13366,N_13875);
and U15404 (N_15404,N_13124,N_12493);
nor U15405 (N_15405,N_12683,N_13649);
or U15406 (N_15406,N_13322,N_12801);
or U15407 (N_15407,N_12656,N_12227);
and U15408 (N_15408,N_13763,N_13253);
xor U15409 (N_15409,N_13669,N_12785);
nand U15410 (N_15410,N_12972,N_12879);
nor U15411 (N_15411,N_13025,N_12694);
or U15412 (N_15412,N_12214,N_12425);
and U15413 (N_15413,N_13633,N_13194);
xnor U15414 (N_15414,N_12893,N_12332);
or U15415 (N_15415,N_13503,N_13027);
and U15416 (N_15416,N_13090,N_13971);
nor U15417 (N_15417,N_13348,N_12144);
nor U15418 (N_15418,N_13004,N_13630);
nor U15419 (N_15419,N_12421,N_12740);
nor U15420 (N_15420,N_13182,N_13034);
xor U15421 (N_15421,N_12288,N_13710);
and U15422 (N_15422,N_13919,N_12894);
nor U15423 (N_15423,N_12556,N_13922);
or U15424 (N_15424,N_13054,N_12013);
or U15425 (N_15425,N_12640,N_13834);
xnor U15426 (N_15426,N_12348,N_12824);
or U15427 (N_15427,N_13167,N_13097);
xor U15428 (N_15428,N_13085,N_12960);
nor U15429 (N_15429,N_13259,N_12354);
xnor U15430 (N_15430,N_13101,N_12524);
nand U15431 (N_15431,N_13051,N_13747);
nand U15432 (N_15432,N_13242,N_13159);
nand U15433 (N_15433,N_13881,N_13708);
nand U15434 (N_15434,N_12652,N_12306);
and U15435 (N_15435,N_13420,N_12557);
xnor U15436 (N_15436,N_13302,N_13113);
and U15437 (N_15437,N_12218,N_13137);
or U15438 (N_15438,N_13990,N_12938);
nor U15439 (N_15439,N_12742,N_13929);
xor U15440 (N_15440,N_12051,N_13965);
nor U15441 (N_15441,N_12571,N_13253);
nor U15442 (N_15442,N_12188,N_13968);
nor U15443 (N_15443,N_13683,N_13208);
xor U15444 (N_15444,N_13514,N_12379);
and U15445 (N_15445,N_12024,N_12580);
nand U15446 (N_15446,N_13149,N_12064);
or U15447 (N_15447,N_12846,N_12266);
nand U15448 (N_15448,N_13245,N_12873);
and U15449 (N_15449,N_12147,N_12830);
xnor U15450 (N_15450,N_12440,N_13197);
and U15451 (N_15451,N_12529,N_13933);
xnor U15452 (N_15452,N_13729,N_13273);
and U15453 (N_15453,N_13695,N_13225);
and U15454 (N_15454,N_13577,N_13335);
xnor U15455 (N_15455,N_12901,N_13559);
and U15456 (N_15456,N_13169,N_13184);
or U15457 (N_15457,N_12199,N_12545);
nor U15458 (N_15458,N_13406,N_13742);
nand U15459 (N_15459,N_12404,N_12820);
nand U15460 (N_15460,N_12984,N_12966);
nor U15461 (N_15461,N_12746,N_13491);
nor U15462 (N_15462,N_12146,N_12710);
nor U15463 (N_15463,N_13975,N_13059);
or U15464 (N_15464,N_12688,N_13653);
xnor U15465 (N_15465,N_13471,N_12387);
and U15466 (N_15466,N_13451,N_13081);
xor U15467 (N_15467,N_12123,N_12611);
nor U15468 (N_15468,N_13202,N_12120);
nand U15469 (N_15469,N_13233,N_12066);
and U15470 (N_15470,N_13761,N_12873);
and U15471 (N_15471,N_13712,N_12823);
and U15472 (N_15472,N_12929,N_13386);
or U15473 (N_15473,N_12678,N_13520);
nor U15474 (N_15474,N_13904,N_12840);
nor U15475 (N_15475,N_13954,N_13623);
and U15476 (N_15476,N_13875,N_13696);
nand U15477 (N_15477,N_13639,N_12620);
or U15478 (N_15478,N_12223,N_13827);
nor U15479 (N_15479,N_12286,N_13088);
nor U15480 (N_15480,N_13909,N_13785);
nor U15481 (N_15481,N_12139,N_12306);
and U15482 (N_15482,N_12805,N_13361);
nand U15483 (N_15483,N_12348,N_12340);
nor U15484 (N_15484,N_12943,N_12091);
and U15485 (N_15485,N_13646,N_13878);
or U15486 (N_15486,N_13869,N_13018);
nor U15487 (N_15487,N_13544,N_12398);
or U15488 (N_15488,N_13911,N_12831);
and U15489 (N_15489,N_12394,N_13905);
nor U15490 (N_15490,N_12384,N_13323);
nand U15491 (N_15491,N_12023,N_13513);
xor U15492 (N_15492,N_13583,N_13488);
nor U15493 (N_15493,N_13274,N_13463);
or U15494 (N_15494,N_12032,N_12808);
xor U15495 (N_15495,N_13304,N_13800);
xnor U15496 (N_15496,N_12225,N_12535);
nand U15497 (N_15497,N_12929,N_12594);
nand U15498 (N_15498,N_13577,N_13206);
or U15499 (N_15499,N_13275,N_13049);
nand U15500 (N_15500,N_13900,N_12054);
nor U15501 (N_15501,N_12643,N_13831);
nand U15502 (N_15502,N_12995,N_12229);
nand U15503 (N_15503,N_13267,N_12706);
nand U15504 (N_15504,N_12048,N_13671);
xor U15505 (N_15505,N_13907,N_12024);
nand U15506 (N_15506,N_12889,N_13382);
or U15507 (N_15507,N_12475,N_13979);
nor U15508 (N_15508,N_12906,N_12330);
and U15509 (N_15509,N_12354,N_13657);
nand U15510 (N_15510,N_12727,N_13487);
nor U15511 (N_15511,N_12211,N_12907);
xor U15512 (N_15512,N_12426,N_13154);
or U15513 (N_15513,N_12557,N_13187);
or U15514 (N_15514,N_13683,N_13773);
nand U15515 (N_15515,N_12428,N_13843);
nand U15516 (N_15516,N_12490,N_12585);
xor U15517 (N_15517,N_12338,N_13715);
nand U15518 (N_15518,N_12722,N_13997);
and U15519 (N_15519,N_12522,N_13015);
and U15520 (N_15520,N_13341,N_13002);
or U15521 (N_15521,N_12306,N_12428);
nand U15522 (N_15522,N_12556,N_12693);
xnor U15523 (N_15523,N_13773,N_12416);
and U15524 (N_15524,N_13901,N_12323);
nand U15525 (N_15525,N_13003,N_13779);
xnor U15526 (N_15526,N_12640,N_12740);
or U15527 (N_15527,N_12906,N_12966);
nand U15528 (N_15528,N_12449,N_12491);
nor U15529 (N_15529,N_12972,N_12232);
or U15530 (N_15530,N_13416,N_13225);
or U15531 (N_15531,N_13147,N_12874);
nor U15532 (N_15532,N_13157,N_12212);
or U15533 (N_15533,N_12830,N_12828);
and U15534 (N_15534,N_13068,N_13934);
or U15535 (N_15535,N_13882,N_13772);
and U15536 (N_15536,N_13229,N_13186);
nand U15537 (N_15537,N_12234,N_13732);
xnor U15538 (N_15538,N_13314,N_13254);
xnor U15539 (N_15539,N_12796,N_12733);
nand U15540 (N_15540,N_13045,N_13380);
nand U15541 (N_15541,N_13991,N_12015);
nor U15542 (N_15542,N_12008,N_12100);
and U15543 (N_15543,N_13046,N_13089);
nand U15544 (N_15544,N_13869,N_12836);
or U15545 (N_15545,N_12783,N_12612);
xnor U15546 (N_15546,N_12570,N_13671);
and U15547 (N_15547,N_12842,N_12200);
nand U15548 (N_15548,N_13765,N_12942);
and U15549 (N_15549,N_12219,N_13568);
nand U15550 (N_15550,N_12472,N_13137);
nor U15551 (N_15551,N_13081,N_12003);
xnor U15552 (N_15552,N_12418,N_13781);
nor U15553 (N_15553,N_12977,N_13151);
and U15554 (N_15554,N_12052,N_13032);
nand U15555 (N_15555,N_12592,N_13768);
nor U15556 (N_15556,N_13513,N_13606);
xor U15557 (N_15557,N_13962,N_12441);
nand U15558 (N_15558,N_13134,N_12205);
nand U15559 (N_15559,N_13780,N_12589);
nand U15560 (N_15560,N_12491,N_13468);
or U15561 (N_15561,N_13298,N_12632);
nand U15562 (N_15562,N_13882,N_13755);
xnor U15563 (N_15563,N_13762,N_13071);
nand U15564 (N_15564,N_12711,N_12297);
nor U15565 (N_15565,N_13926,N_12387);
nand U15566 (N_15566,N_12657,N_13926);
nor U15567 (N_15567,N_13690,N_12149);
nand U15568 (N_15568,N_13318,N_12502);
or U15569 (N_15569,N_12691,N_13796);
nand U15570 (N_15570,N_12982,N_13250);
xor U15571 (N_15571,N_12000,N_13070);
nand U15572 (N_15572,N_13480,N_12639);
nand U15573 (N_15573,N_12520,N_12252);
or U15574 (N_15574,N_13239,N_13029);
or U15575 (N_15575,N_13766,N_13262);
nand U15576 (N_15576,N_12530,N_13143);
nand U15577 (N_15577,N_13893,N_13185);
and U15578 (N_15578,N_13855,N_12420);
nand U15579 (N_15579,N_13557,N_12594);
nor U15580 (N_15580,N_12373,N_12736);
nand U15581 (N_15581,N_13232,N_12224);
nor U15582 (N_15582,N_13190,N_13762);
and U15583 (N_15583,N_12563,N_13760);
nand U15584 (N_15584,N_12592,N_12544);
xnor U15585 (N_15585,N_12939,N_12591);
and U15586 (N_15586,N_13676,N_12017);
xor U15587 (N_15587,N_12056,N_13198);
nor U15588 (N_15588,N_12301,N_12334);
nor U15589 (N_15589,N_12332,N_13359);
xor U15590 (N_15590,N_12259,N_12518);
nand U15591 (N_15591,N_13781,N_12629);
nand U15592 (N_15592,N_12148,N_13433);
xnor U15593 (N_15593,N_13041,N_12858);
or U15594 (N_15594,N_13048,N_12558);
nand U15595 (N_15595,N_13133,N_13508);
xnor U15596 (N_15596,N_13883,N_12899);
nand U15597 (N_15597,N_13871,N_12880);
xnor U15598 (N_15598,N_12426,N_13249);
or U15599 (N_15599,N_13407,N_12668);
and U15600 (N_15600,N_12290,N_12253);
nor U15601 (N_15601,N_12595,N_13746);
or U15602 (N_15602,N_12964,N_13691);
nand U15603 (N_15603,N_13768,N_12879);
or U15604 (N_15604,N_12479,N_12314);
or U15605 (N_15605,N_12587,N_12304);
nand U15606 (N_15606,N_12186,N_13151);
or U15607 (N_15607,N_13742,N_13058);
and U15608 (N_15608,N_12693,N_12316);
or U15609 (N_15609,N_12767,N_13263);
or U15610 (N_15610,N_13077,N_13804);
or U15611 (N_15611,N_13896,N_13360);
nor U15612 (N_15612,N_13387,N_12501);
nor U15613 (N_15613,N_12519,N_13492);
nand U15614 (N_15614,N_13461,N_12900);
xnor U15615 (N_15615,N_12905,N_13658);
and U15616 (N_15616,N_13612,N_12599);
or U15617 (N_15617,N_13710,N_13469);
nor U15618 (N_15618,N_13549,N_13657);
xnor U15619 (N_15619,N_12971,N_13407);
nor U15620 (N_15620,N_12475,N_12493);
and U15621 (N_15621,N_12245,N_12990);
nand U15622 (N_15622,N_13417,N_13850);
or U15623 (N_15623,N_13459,N_12407);
and U15624 (N_15624,N_12630,N_12828);
nand U15625 (N_15625,N_12733,N_12843);
and U15626 (N_15626,N_12982,N_13099);
nor U15627 (N_15627,N_13584,N_12384);
nand U15628 (N_15628,N_12833,N_13857);
nand U15629 (N_15629,N_13167,N_13834);
nand U15630 (N_15630,N_13249,N_13511);
and U15631 (N_15631,N_13007,N_13404);
and U15632 (N_15632,N_12768,N_12165);
xor U15633 (N_15633,N_13026,N_13646);
or U15634 (N_15634,N_13264,N_12072);
or U15635 (N_15635,N_12570,N_12162);
xnor U15636 (N_15636,N_13922,N_13026);
and U15637 (N_15637,N_12433,N_12664);
nor U15638 (N_15638,N_12747,N_12381);
nor U15639 (N_15639,N_13138,N_12331);
and U15640 (N_15640,N_12967,N_12858);
nand U15641 (N_15641,N_12408,N_12309);
nor U15642 (N_15642,N_12002,N_13912);
nor U15643 (N_15643,N_12548,N_12050);
nor U15644 (N_15644,N_12708,N_12419);
xnor U15645 (N_15645,N_12671,N_13833);
nand U15646 (N_15646,N_12706,N_12521);
nor U15647 (N_15647,N_12882,N_13266);
xor U15648 (N_15648,N_12626,N_13304);
nand U15649 (N_15649,N_13752,N_12335);
and U15650 (N_15650,N_12997,N_12399);
nor U15651 (N_15651,N_12247,N_12569);
nor U15652 (N_15652,N_13396,N_13105);
nor U15653 (N_15653,N_12844,N_12816);
or U15654 (N_15654,N_13837,N_13351);
nor U15655 (N_15655,N_12499,N_12894);
or U15656 (N_15656,N_12819,N_12376);
nand U15657 (N_15657,N_13600,N_13606);
and U15658 (N_15658,N_12612,N_12888);
and U15659 (N_15659,N_12942,N_13125);
nor U15660 (N_15660,N_13584,N_12414);
nand U15661 (N_15661,N_13180,N_12185);
nor U15662 (N_15662,N_13741,N_13556);
nor U15663 (N_15663,N_13474,N_12693);
or U15664 (N_15664,N_13714,N_13916);
or U15665 (N_15665,N_12764,N_13496);
nand U15666 (N_15666,N_12840,N_12198);
and U15667 (N_15667,N_13856,N_12676);
xor U15668 (N_15668,N_13284,N_12964);
nand U15669 (N_15669,N_13631,N_13083);
or U15670 (N_15670,N_12036,N_12685);
nand U15671 (N_15671,N_13062,N_12925);
nor U15672 (N_15672,N_13752,N_13026);
xnor U15673 (N_15673,N_13813,N_13218);
xor U15674 (N_15674,N_12622,N_13273);
nor U15675 (N_15675,N_13515,N_13606);
xnor U15676 (N_15676,N_12855,N_13515);
or U15677 (N_15677,N_13388,N_12963);
and U15678 (N_15678,N_13952,N_13906);
and U15679 (N_15679,N_12608,N_13835);
xnor U15680 (N_15680,N_12162,N_12872);
xnor U15681 (N_15681,N_12562,N_12615);
nor U15682 (N_15682,N_12885,N_13546);
and U15683 (N_15683,N_12626,N_12368);
and U15684 (N_15684,N_13391,N_13716);
and U15685 (N_15685,N_13852,N_13269);
nand U15686 (N_15686,N_12855,N_13134);
xnor U15687 (N_15687,N_12564,N_12335);
nand U15688 (N_15688,N_12146,N_12911);
nand U15689 (N_15689,N_12348,N_13017);
and U15690 (N_15690,N_12463,N_12484);
or U15691 (N_15691,N_12677,N_13818);
and U15692 (N_15692,N_13930,N_13264);
and U15693 (N_15693,N_12864,N_13539);
and U15694 (N_15694,N_12009,N_12922);
nor U15695 (N_15695,N_13988,N_12604);
or U15696 (N_15696,N_13312,N_12077);
xnor U15697 (N_15697,N_12654,N_12085);
or U15698 (N_15698,N_13835,N_12110);
and U15699 (N_15699,N_13020,N_13923);
xnor U15700 (N_15700,N_13834,N_12502);
or U15701 (N_15701,N_12566,N_13360);
nor U15702 (N_15702,N_13779,N_13637);
nand U15703 (N_15703,N_13148,N_13080);
xnor U15704 (N_15704,N_12128,N_12611);
nor U15705 (N_15705,N_13712,N_12786);
or U15706 (N_15706,N_12349,N_12469);
and U15707 (N_15707,N_12984,N_12235);
or U15708 (N_15708,N_13766,N_13744);
or U15709 (N_15709,N_12110,N_13622);
or U15710 (N_15710,N_13747,N_12340);
nor U15711 (N_15711,N_13159,N_13130);
or U15712 (N_15712,N_13770,N_13253);
xnor U15713 (N_15713,N_13132,N_13957);
and U15714 (N_15714,N_13509,N_13280);
xnor U15715 (N_15715,N_12379,N_12690);
and U15716 (N_15716,N_12605,N_13114);
xnor U15717 (N_15717,N_12708,N_13636);
nor U15718 (N_15718,N_12835,N_13105);
or U15719 (N_15719,N_12498,N_12743);
nor U15720 (N_15720,N_12836,N_13580);
nor U15721 (N_15721,N_13591,N_12764);
nand U15722 (N_15722,N_12157,N_13895);
nor U15723 (N_15723,N_12050,N_13852);
nand U15724 (N_15724,N_13570,N_12082);
xor U15725 (N_15725,N_12229,N_13782);
nor U15726 (N_15726,N_13713,N_13191);
and U15727 (N_15727,N_13094,N_13648);
nor U15728 (N_15728,N_12306,N_12146);
xnor U15729 (N_15729,N_12015,N_13543);
and U15730 (N_15730,N_13884,N_13001);
nor U15731 (N_15731,N_12987,N_12142);
xnor U15732 (N_15732,N_13130,N_12021);
and U15733 (N_15733,N_13249,N_12427);
nand U15734 (N_15734,N_13840,N_12630);
nand U15735 (N_15735,N_13559,N_13869);
or U15736 (N_15736,N_12852,N_13540);
and U15737 (N_15737,N_12795,N_13408);
or U15738 (N_15738,N_12807,N_12191);
or U15739 (N_15739,N_13579,N_13886);
or U15740 (N_15740,N_13780,N_12026);
nand U15741 (N_15741,N_12442,N_12317);
and U15742 (N_15742,N_12104,N_12207);
or U15743 (N_15743,N_13404,N_13981);
and U15744 (N_15744,N_13425,N_12859);
nand U15745 (N_15745,N_12848,N_13436);
nand U15746 (N_15746,N_13094,N_12718);
xnor U15747 (N_15747,N_13864,N_12596);
nand U15748 (N_15748,N_12973,N_12511);
xor U15749 (N_15749,N_13517,N_13054);
nor U15750 (N_15750,N_12573,N_12437);
nor U15751 (N_15751,N_12331,N_13898);
xor U15752 (N_15752,N_13272,N_13313);
or U15753 (N_15753,N_13439,N_13387);
nand U15754 (N_15754,N_12901,N_13214);
and U15755 (N_15755,N_13186,N_13061);
nor U15756 (N_15756,N_13054,N_12474);
nand U15757 (N_15757,N_13601,N_12302);
nand U15758 (N_15758,N_13463,N_13456);
nand U15759 (N_15759,N_13068,N_12652);
or U15760 (N_15760,N_13115,N_12828);
xor U15761 (N_15761,N_12453,N_12408);
xnor U15762 (N_15762,N_13399,N_13518);
nor U15763 (N_15763,N_13676,N_12821);
nand U15764 (N_15764,N_13909,N_12198);
nor U15765 (N_15765,N_12880,N_12464);
nor U15766 (N_15766,N_12829,N_12132);
xor U15767 (N_15767,N_12020,N_12665);
nand U15768 (N_15768,N_13922,N_13899);
xor U15769 (N_15769,N_13091,N_13716);
nand U15770 (N_15770,N_13405,N_13812);
and U15771 (N_15771,N_13931,N_13050);
nor U15772 (N_15772,N_13299,N_12417);
or U15773 (N_15773,N_12322,N_13544);
xor U15774 (N_15774,N_12544,N_12874);
or U15775 (N_15775,N_13348,N_13833);
or U15776 (N_15776,N_13161,N_12927);
or U15777 (N_15777,N_13864,N_13849);
nor U15778 (N_15778,N_13500,N_13848);
and U15779 (N_15779,N_13371,N_12549);
and U15780 (N_15780,N_13308,N_12869);
and U15781 (N_15781,N_13087,N_13368);
nor U15782 (N_15782,N_12104,N_12186);
nor U15783 (N_15783,N_12381,N_12880);
nor U15784 (N_15784,N_13153,N_12900);
nand U15785 (N_15785,N_12336,N_13880);
nand U15786 (N_15786,N_13126,N_13368);
nor U15787 (N_15787,N_12562,N_12117);
or U15788 (N_15788,N_12991,N_12167);
and U15789 (N_15789,N_12734,N_13100);
or U15790 (N_15790,N_12480,N_12958);
nor U15791 (N_15791,N_12576,N_13865);
and U15792 (N_15792,N_13148,N_12318);
xnor U15793 (N_15793,N_13548,N_13993);
nand U15794 (N_15794,N_13368,N_12824);
nor U15795 (N_15795,N_13201,N_12973);
nor U15796 (N_15796,N_12105,N_12454);
and U15797 (N_15797,N_13561,N_12829);
nand U15798 (N_15798,N_12327,N_12461);
or U15799 (N_15799,N_12419,N_12044);
nand U15800 (N_15800,N_12682,N_13018);
and U15801 (N_15801,N_12677,N_13447);
nand U15802 (N_15802,N_12438,N_12202);
and U15803 (N_15803,N_12945,N_12806);
or U15804 (N_15804,N_13875,N_12840);
and U15805 (N_15805,N_13735,N_12860);
or U15806 (N_15806,N_12009,N_12193);
and U15807 (N_15807,N_12960,N_12972);
xnor U15808 (N_15808,N_12049,N_13534);
or U15809 (N_15809,N_12548,N_13623);
xnor U15810 (N_15810,N_12821,N_12500);
xnor U15811 (N_15811,N_13390,N_12173);
nor U15812 (N_15812,N_12877,N_12015);
nor U15813 (N_15813,N_13581,N_13776);
nand U15814 (N_15814,N_13382,N_12196);
or U15815 (N_15815,N_12793,N_12139);
nor U15816 (N_15816,N_13736,N_12607);
xor U15817 (N_15817,N_13657,N_12102);
or U15818 (N_15818,N_13527,N_12271);
nand U15819 (N_15819,N_13250,N_13298);
and U15820 (N_15820,N_12387,N_12258);
nand U15821 (N_15821,N_13316,N_12887);
and U15822 (N_15822,N_13999,N_12960);
or U15823 (N_15823,N_12358,N_12919);
nor U15824 (N_15824,N_12832,N_13047);
and U15825 (N_15825,N_12449,N_12644);
or U15826 (N_15826,N_13570,N_13265);
xnor U15827 (N_15827,N_13782,N_12114);
or U15828 (N_15828,N_12974,N_12471);
xnor U15829 (N_15829,N_12279,N_12864);
and U15830 (N_15830,N_12062,N_12131);
and U15831 (N_15831,N_12149,N_12981);
or U15832 (N_15832,N_12271,N_12036);
xor U15833 (N_15833,N_12046,N_12834);
and U15834 (N_15834,N_12463,N_12176);
and U15835 (N_15835,N_13855,N_12850);
xor U15836 (N_15836,N_12813,N_13971);
xnor U15837 (N_15837,N_12907,N_13314);
and U15838 (N_15838,N_13029,N_13645);
and U15839 (N_15839,N_13720,N_12521);
nand U15840 (N_15840,N_12698,N_13988);
nand U15841 (N_15841,N_13208,N_13242);
xnor U15842 (N_15842,N_13605,N_12442);
nand U15843 (N_15843,N_13747,N_13540);
and U15844 (N_15844,N_13430,N_12327);
or U15845 (N_15845,N_13484,N_12718);
and U15846 (N_15846,N_12775,N_13413);
or U15847 (N_15847,N_13097,N_13896);
and U15848 (N_15848,N_13003,N_12846);
xnor U15849 (N_15849,N_13480,N_13831);
and U15850 (N_15850,N_12798,N_12536);
nor U15851 (N_15851,N_13552,N_12628);
or U15852 (N_15852,N_12508,N_12667);
and U15853 (N_15853,N_12772,N_13167);
and U15854 (N_15854,N_12528,N_12409);
nand U15855 (N_15855,N_13786,N_13012);
nand U15856 (N_15856,N_12811,N_13595);
nor U15857 (N_15857,N_13846,N_12100);
and U15858 (N_15858,N_13545,N_13539);
xor U15859 (N_15859,N_13102,N_13653);
xor U15860 (N_15860,N_12304,N_13576);
nor U15861 (N_15861,N_13503,N_13395);
nand U15862 (N_15862,N_13768,N_12263);
or U15863 (N_15863,N_12528,N_13370);
nor U15864 (N_15864,N_12705,N_13696);
nand U15865 (N_15865,N_13776,N_12317);
xnor U15866 (N_15866,N_13478,N_12574);
nor U15867 (N_15867,N_12590,N_12858);
xor U15868 (N_15868,N_13060,N_13899);
nand U15869 (N_15869,N_13236,N_12072);
or U15870 (N_15870,N_12068,N_13280);
and U15871 (N_15871,N_13680,N_12299);
nand U15872 (N_15872,N_12924,N_13946);
xor U15873 (N_15873,N_12088,N_12587);
nand U15874 (N_15874,N_13855,N_13718);
xor U15875 (N_15875,N_13681,N_13630);
and U15876 (N_15876,N_13212,N_12436);
nand U15877 (N_15877,N_13330,N_12184);
or U15878 (N_15878,N_12983,N_13382);
nor U15879 (N_15879,N_13904,N_13202);
nor U15880 (N_15880,N_13269,N_12748);
nand U15881 (N_15881,N_13483,N_13029);
xnor U15882 (N_15882,N_12908,N_12140);
or U15883 (N_15883,N_13703,N_13903);
nand U15884 (N_15884,N_12091,N_12929);
nand U15885 (N_15885,N_13600,N_13969);
xnor U15886 (N_15886,N_12581,N_13549);
or U15887 (N_15887,N_12458,N_13852);
nor U15888 (N_15888,N_13115,N_13306);
or U15889 (N_15889,N_12103,N_13167);
nor U15890 (N_15890,N_12964,N_13746);
and U15891 (N_15891,N_13889,N_12398);
xor U15892 (N_15892,N_12757,N_13475);
and U15893 (N_15893,N_12654,N_12041);
nand U15894 (N_15894,N_13934,N_12826);
or U15895 (N_15895,N_12033,N_13796);
or U15896 (N_15896,N_12768,N_13015);
and U15897 (N_15897,N_12895,N_12613);
nor U15898 (N_15898,N_12237,N_12969);
or U15899 (N_15899,N_12674,N_13122);
xnor U15900 (N_15900,N_13876,N_12559);
and U15901 (N_15901,N_13026,N_13023);
or U15902 (N_15902,N_13936,N_13691);
or U15903 (N_15903,N_12730,N_12701);
nand U15904 (N_15904,N_13137,N_13739);
nor U15905 (N_15905,N_12216,N_13953);
nand U15906 (N_15906,N_13566,N_12249);
and U15907 (N_15907,N_12602,N_13748);
or U15908 (N_15908,N_12779,N_13061);
xor U15909 (N_15909,N_12272,N_12017);
nor U15910 (N_15910,N_13303,N_13752);
nor U15911 (N_15911,N_13118,N_12303);
nor U15912 (N_15912,N_13301,N_13050);
nand U15913 (N_15913,N_13243,N_13039);
nor U15914 (N_15914,N_12206,N_13695);
nor U15915 (N_15915,N_13050,N_12840);
nor U15916 (N_15916,N_12233,N_12158);
xor U15917 (N_15917,N_12341,N_13615);
nand U15918 (N_15918,N_12213,N_12966);
nor U15919 (N_15919,N_13621,N_12921);
nor U15920 (N_15920,N_13588,N_13000);
xor U15921 (N_15921,N_13015,N_13977);
xor U15922 (N_15922,N_12476,N_13512);
xor U15923 (N_15923,N_12264,N_12572);
and U15924 (N_15924,N_12935,N_12710);
or U15925 (N_15925,N_13201,N_12307);
nor U15926 (N_15926,N_12748,N_13398);
or U15927 (N_15927,N_13776,N_13595);
nand U15928 (N_15928,N_12759,N_13171);
nand U15929 (N_15929,N_12825,N_12527);
nand U15930 (N_15930,N_13397,N_12639);
and U15931 (N_15931,N_12626,N_13091);
or U15932 (N_15932,N_12143,N_12348);
xor U15933 (N_15933,N_13920,N_13216);
and U15934 (N_15934,N_12466,N_13698);
nor U15935 (N_15935,N_13673,N_13984);
xor U15936 (N_15936,N_12841,N_12210);
xor U15937 (N_15937,N_13561,N_12250);
and U15938 (N_15938,N_13223,N_13091);
and U15939 (N_15939,N_13257,N_12983);
and U15940 (N_15940,N_12971,N_12463);
or U15941 (N_15941,N_13439,N_12016);
nor U15942 (N_15942,N_13412,N_13029);
or U15943 (N_15943,N_12124,N_12608);
xnor U15944 (N_15944,N_12468,N_12872);
nor U15945 (N_15945,N_12641,N_12825);
and U15946 (N_15946,N_12489,N_12692);
nand U15947 (N_15947,N_12934,N_13499);
and U15948 (N_15948,N_12961,N_12489);
xor U15949 (N_15949,N_13840,N_12392);
xor U15950 (N_15950,N_12760,N_12993);
or U15951 (N_15951,N_13427,N_12263);
or U15952 (N_15952,N_12898,N_13739);
nor U15953 (N_15953,N_12512,N_13624);
nand U15954 (N_15954,N_13317,N_12011);
nor U15955 (N_15955,N_12376,N_12106);
nor U15956 (N_15956,N_13797,N_13301);
nand U15957 (N_15957,N_13003,N_13242);
nand U15958 (N_15958,N_12619,N_12898);
or U15959 (N_15959,N_12382,N_12600);
nand U15960 (N_15960,N_12515,N_12021);
or U15961 (N_15961,N_12863,N_13709);
xnor U15962 (N_15962,N_12455,N_13251);
nand U15963 (N_15963,N_12994,N_12862);
xnor U15964 (N_15964,N_12051,N_13503);
and U15965 (N_15965,N_12340,N_12576);
and U15966 (N_15966,N_13647,N_13801);
and U15967 (N_15967,N_13463,N_13245);
nor U15968 (N_15968,N_13814,N_12650);
nor U15969 (N_15969,N_12406,N_12125);
or U15970 (N_15970,N_12014,N_12648);
xor U15971 (N_15971,N_13934,N_12548);
nor U15972 (N_15972,N_12818,N_12187);
and U15973 (N_15973,N_12486,N_12054);
nor U15974 (N_15974,N_13744,N_12101);
nor U15975 (N_15975,N_12571,N_12658);
or U15976 (N_15976,N_13607,N_13925);
xor U15977 (N_15977,N_12094,N_12732);
or U15978 (N_15978,N_13812,N_12307);
nor U15979 (N_15979,N_13600,N_13294);
and U15980 (N_15980,N_12984,N_13005);
nor U15981 (N_15981,N_12219,N_13019);
nor U15982 (N_15982,N_12440,N_13125);
xnor U15983 (N_15983,N_13014,N_12375);
nor U15984 (N_15984,N_12981,N_13406);
nand U15985 (N_15985,N_12639,N_13269);
or U15986 (N_15986,N_13123,N_13670);
and U15987 (N_15987,N_13451,N_13326);
and U15988 (N_15988,N_13073,N_12584);
nor U15989 (N_15989,N_12075,N_13573);
xnor U15990 (N_15990,N_13744,N_13972);
and U15991 (N_15991,N_13072,N_12427);
xnor U15992 (N_15992,N_12535,N_12393);
nand U15993 (N_15993,N_12326,N_12232);
nor U15994 (N_15994,N_12734,N_12317);
xnor U15995 (N_15995,N_12779,N_13393);
nand U15996 (N_15996,N_12245,N_13176);
nand U15997 (N_15997,N_12999,N_13479);
nor U15998 (N_15998,N_12975,N_12210);
and U15999 (N_15999,N_12434,N_13847);
nor U16000 (N_16000,N_14502,N_14997);
nand U16001 (N_16001,N_14040,N_14727);
and U16002 (N_16002,N_15685,N_14057);
xor U16003 (N_16003,N_14840,N_14965);
and U16004 (N_16004,N_14287,N_15654);
or U16005 (N_16005,N_15148,N_14632);
nor U16006 (N_16006,N_15607,N_15163);
nand U16007 (N_16007,N_15938,N_15346);
and U16008 (N_16008,N_14753,N_14741);
and U16009 (N_16009,N_15397,N_14089);
and U16010 (N_16010,N_15307,N_14412);
nor U16011 (N_16011,N_14608,N_15978);
nor U16012 (N_16012,N_14196,N_15395);
nor U16013 (N_16013,N_14655,N_15811);
and U16014 (N_16014,N_15056,N_14529);
and U16015 (N_16015,N_14540,N_15219);
nand U16016 (N_16016,N_15286,N_14691);
nor U16017 (N_16017,N_15314,N_15920);
and U16018 (N_16018,N_14309,N_14630);
or U16019 (N_16019,N_15534,N_14519);
or U16020 (N_16020,N_14807,N_15568);
nand U16021 (N_16021,N_14957,N_15203);
nor U16022 (N_16022,N_14081,N_14269);
and U16023 (N_16023,N_14652,N_14709);
or U16024 (N_16024,N_15466,N_14746);
xnor U16025 (N_16025,N_15726,N_15894);
nand U16026 (N_16026,N_14758,N_15318);
or U16027 (N_16027,N_14112,N_14738);
nor U16028 (N_16028,N_14587,N_14847);
nor U16029 (N_16029,N_14487,N_15470);
nand U16030 (N_16030,N_14201,N_15027);
and U16031 (N_16031,N_15889,N_15038);
nor U16032 (N_16032,N_15487,N_14174);
nor U16033 (N_16033,N_14943,N_15522);
nand U16034 (N_16034,N_14398,N_14233);
and U16035 (N_16035,N_15228,N_15253);
nand U16036 (N_16036,N_14234,N_14853);
xnor U16037 (N_16037,N_15639,N_15009);
and U16038 (N_16038,N_14604,N_15429);
nor U16039 (N_16039,N_14792,N_14590);
nor U16040 (N_16040,N_15097,N_14973);
nor U16041 (N_16041,N_15138,N_14543);
xor U16042 (N_16042,N_14639,N_14078);
xor U16043 (N_16043,N_14416,N_14922);
nand U16044 (N_16044,N_15695,N_14192);
or U16045 (N_16045,N_14161,N_14423);
or U16046 (N_16046,N_15855,N_14938);
nand U16047 (N_16047,N_14051,N_14194);
nand U16048 (N_16048,N_14814,N_14380);
or U16049 (N_16049,N_14681,N_15718);
nor U16050 (N_16050,N_14025,N_15349);
nor U16051 (N_16051,N_14110,N_14743);
or U16052 (N_16052,N_14768,N_15274);
xor U16053 (N_16053,N_15542,N_15198);
or U16054 (N_16054,N_14588,N_15376);
xnor U16055 (N_16055,N_14636,N_14512);
and U16056 (N_16056,N_15705,N_15689);
nor U16057 (N_16057,N_15757,N_15406);
nand U16058 (N_16058,N_15999,N_15847);
and U16059 (N_16059,N_14043,N_15641);
and U16060 (N_16060,N_14185,N_15361);
and U16061 (N_16061,N_14167,N_15371);
xor U16062 (N_16062,N_14933,N_15417);
or U16063 (N_16063,N_15856,N_14061);
xor U16064 (N_16064,N_15142,N_15749);
nor U16065 (N_16065,N_15263,N_15020);
nand U16066 (N_16066,N_15991,N_14300);
nand U16067 (N_16067,N_14831,N_14123);
nand U16068 (N_16068,N_14094,N_14541);
and U16069 (N_16069,N_15881,N_14978);
nand U16070 (N_16070,N_14053,N_14535);
or U16071 (N_16071,N_15330,N_15684);
xnor U16072 (N_16072,N_14224,N_15128);
and U16073 (N_16073,N_15408,N_14808);
or U16074 (N_16074,N_14996,N_15895);
nand U16075 (N_16075,N_14804,N_14118);
nand U16076 (N_16076,N_15779,N_14940);
and U16077 (N_16077,N_14146,N_14248);
or U16078 (N_16078,N_15801,N_14084);
xnor U16079 (N_16079,N_14335,N_15634);
xnor U16080 (N_16080,N_15167,N_15582);
nand U16081 (N_16081,N_14564,N_14376);
or U16082 (N_16082,N_14357,N_14360);
or U16083 (N_16083,N_15019,N_14531);
and U16084 (N_16084,N_15984,N_14657);
nand U16085 (N_16085,N_14607,N_15183);
nand U16086 (N_16086,N_14599,N_14033);
and U16087 (N_16087,N_14782,N_15992);
xnor U16088 (N_16088,N_15182,N_14121);
nor U16089 (N_16089,N_14314,N_15956);
or U16090 (N_16090,N_15465,N_14472);
nand U16091 (N_16091,N_14460,N_14644);
and U16092 (N_16092,N_14346,N_15975);
xnor U16093 (N_16093,N_14769,N_15015);
nand U16094 (N_16094,N_15945,N_15977);
xor U16095 (N_16095,N_14881,N_15277);
xor U16096 (N_16096,N_15325,N_15261);
nand U16097 (N_16097,N_14381,N_14001);
nor U16098 (N_16098,N_14455,N_14092);
xnor U16099 (N_16099,N_14942,N_14833);
nand U16100 (N_16100,N_15815,N_15031);
nand U16101 (N_16101,N_15396,N_15192);
nand U16102 (N_16102,N_15510,N_14260);
nand U16103 (N_16103,N_14690,N_14202);
xor U16104 (N_16104,N_14336,N_14988);
or U16105 (N_16105,N_15890,N_15951);
or U16106 (N_16106,N_15301,N_15653);
xor U16107 (N_16107,N_14851,N_15485);
or U16108 (N_16108,N_15365,N_15401);
nand U16109 (N_16109,N_15870,N_15159);
and U16110 (N_16110,N_14508,N_15717);
nand U16111 (N_16111,N_14748,N_15518);
xor U16112 (N_16112,N_14342,N_15719);
or U16113 (N_16113,N_15958,N_15494);
or U16114 (N_16114,N_15362,N_14030);
nand U16115 (N_16115,N_14023,N_14917);
nor U16116 (N_16116,N_15168,N_14132);
nor U16117 (N_16117,N_14204,N_15593);
and U16118 (N_16118,N_15354,N_15803);
nor U16119 (N_16119,N_14638,N_15981);
or U16120 (N_16120,N_15824,N_14082);
xnor U16121 (N_16121,N_15434,N_15708);
or U16122 (N_16122,N_15216,N_15575);
nand U16123 (N_16123,N_15309,N_15533);
and U16124 (N_16124,N_14715,N_14553);
nand U16125 (N_16125,N_15756,N_15551);
or U16126 (N_16126,N_15094,N_15051);
nor U16127 (N_16127,N_15295,N_14976);
nor U16128 (N_16128,N_14179,N_14819);
nor U16129 (N_16129,N_14296,N_14359);
or U16130 (N_16130,N_15250,N_14492);
nor U16131 (N_16131,N_14718,N_14418);
and U16132 (N_16132,N_14600,N_15730);
nor U16133 (N_16133,N_14151,N_14576);
nor U16134 (N_16134,N_14845,N_15802);
xor U16135 (N_16135,N_15498,N_14232);
and U16136 (N_16136,N_15530,N_15567);
or U16137 (N_16137,N_15058,N_14216);
xor U16138 (N_16138,N_15317,N_15028);
and U16139 (N_16139,N_14706,N_15714);
xor U16140 (N_16140,N_14563,N_14333);
xnor U16141 (N_16141,N_14364,N_14006);
and U16142 (N_16142,N_15449,N_15863);
nor U16143 (N_16143,N_14307,N_15196);
or U16144 (N_16144,N_15191,N_15915);
nand U16145 (N_16145,N_15520,N_14984);
xor U16146 (N_16146,N_15675,N_15215);
nor U16147 (N_16147,N_14742,N_15688);
or U16148 (N_16148,N_15658,N_15060);
nand U16149 (N_16149,N_14325,N_15866);
nand U16150 (N_16150,N_14409,N_15254);
and U16151 (N_16151,N_14760,N_15784);
and U16152 (N_16152,N_15770,N_14169);
xor U16153 (N_16153,N_14949,N_14454);
nor U16154 (N_16154,N_14087,N_15605);
xnor U16155 (N_16155,N_15320,N_15739);
nand U16156 (N_16156,N_14417,N_14008);
nand U16157 (N_16157,N_14446,N_15569);
nand U16158 (N_16158,N_14612,N_15800);
and U16159 (N_16159,N_14953,N_14637);
and U16160 (N_16160,N_14911,N_15900);
nand U16161 (N_16161,N_14343,N_14056);
and U16162 (N_16162,N_15002,N_14730);
nor U16163 (N_16163,N_14824,N_15791);
or U16164 (N_16164,N_14634,N_15189);
nand U16165 (N_16165,N_14207,N_15294);
nor U16166 (N_16166,N_14397,N_14285);
nand U16167 (N_16167,N_15041,N_14931);
xor U16168 (N_16168,N_15130,N_14992);
xnor U16169 (N_16169,N_15502,N_15204);
xnor U16170 (N_16170,N_14827,N_14394);
nor U16171 (N_16171,N_14475,N_14062);
xor U16172 (N_16172,N_14341,N_15422);
and U16173 (N_16173,N_14182,N_15728);
or U16174 (N_16174,N_14131,N_15761);
and U16175 (N_16175,N_15767,N_15143);
and U16176 (N_16176,N_14031,N_14980);
nor U16177 (N_16177,N_14323,N_14313);
and U16178 (N_16178,N_14408,N_15932);
xnor U16179 (N_16179,N_14879,N_15300);
and U16180 (N_16180,N_15202,N_15570);
nand U16181 (N_16181,N_15988,N_15242);
nor U16182 (N_16182,N_14858,N_15360);
and U16183 (N_16183,N_14689,N_15156);
and U16184 (N_16184,N_15591,N_15065);
nand U16185 (N_16185,N_14203,N_15917);
nand U16186 (N_16186,N_15833,N_15876);
and U16187 (N_16187,N_14580,N_14015);
nand U16188 (N_16188,N_15513,N_14361);
nand U16189 (N_16189,N_14319,N_14539);
or U16190 (N_16190,N_15543,N_14405);
or U16191 (N_16191,N_14685,N_15733);
xnor U16192 (N_16192,N_15479,N_15562);
nor U16193 (N_16193,N_14795,N_15854);
nor U16194 (N_16194,N_15971,N_15979);
and U16195 (N_16195,N_14304,N_15586);
or U16196 (N_16196,N_15293,N_14910);
nor U16197 (N_16197,N_14867,N_14733);
nand U16198 (N_16198,N_14303,N_15418);
xor U16199 (N_16199,N_15862,N_14901);
nor U16200 (N_16200,N_15943,N_15305);
xnor U16201 (N_16201,N_15617,N_14291);
nand U16202 (N_16202,N_15554,N_14660);
or U16203 (N_16203,N_15859,N_14666);
nor U16204 (N_16204,N_14515,N_15195);
nand U16205 (N_16205,N_15760,N_15087);
nand U16206 (N_16206,N_15393,N_15967);
nand U16207 (N_16207,N_14068,N_14869);
or U16208 (N_16208,N_15740,N_14915);
xnor U16209 (N_16209,N_14035,N_14072);
nand U16210 (N_16210,N_14048,N_14989);
xor U16211 (N_16211,N_14284,N_14491);
nor U16212 (N_16212,N_15414,N_15768);
nand U16213 (N_16213,N_15339,N_15608);
and U16214 (N_16214,N_14972,N_15332);
nor U16215 (N_16215,N_14547,N_15909);
and U16216 (N_16216,N_15382,N_14778);
and U16217 (N_16217,N_14702,N_14431);
nor U16218 (N_16218,N_14872,N_14424);
nand U16219 (N_16219,N_14740,N_14999);
and U16220 (N_16220,N_14214,N_15882);
xor U16221 (N_16221,N_14560,N_14648);
nand U16222 (N_16222,N_14322,N_14878);
nor U16223 (N_16223,N_15590,N_15524);
and U16224 (N_16224,N_14227,N_14661);
nand U16225 (N_16225,N_15954,N_14402);
and U16226 (N_16226,N_15662,N_15758);
and U16227 (N_16227,N_14631,N_15098);
and U16228 (N_16228,N_15095,N_15257);
or U16229 (N_16229,N_15583,N_15121);
nor U16230 (N_16230,N_14271,N_14886);
nand U16231 (N_16231,N_15231,N_15877);
xor U16232 (N_16232,N_15853,N_14628);
and U16233 (N_16233,N_14974,N_14348);
nor U16234 (N_16234,N_14645,N_15521);
nand U16235 (N_16235,N_14712,N_15721);
xnor U16236 (N_16236,N_14830,N_14926);
or U16237 (N_16237,N_14774,N_14399);
nand U16238 (N_16238,N_15926,N_15319);
nor U16239 (N_16239,N_14002,N_14134);
nor U16240 (N_16240,N_14324,N_14396);
nand U16241 (N_16241,N_14751,N_15334);
xnor U16242 (N_16242,N_14523,N_15503);
nand U16243 (N_16243,N_14622,N_14994);
and U16244 (N_16244,N_15129,N_15244);
nand U16245 (N_16245,N_14102,N_14171);
and U16246 (N_16246,N_14905,N_15112);
nand U16247 (N_16247,N_14286,N_14617);
nor U16248 (N_16248,N_15837,N_14384);
nand U16249 (N_16249,N_14039,N_14744);
xor U16250 (N_16250,N_14267,N_15086);
and U16251 (N_16251,N_14443,N_14242);
or U16252 (N_16252,N_14662,N_14776);
nand U16253 (N_16253,N_14537,N_14559);
nand U16254 (N_16254,N_15676,N_15716);
nand U16255 (N_16255,N_14029,N_14841);
nand U16256 (N_16256,N_14301,N_15432);
nor U16257 (N_16257,N_14725,N_14852);
xor U16258 (N_16258,N_14961,N_14832);
xnor U16259 (N_16259,N_15797,N_15311);
nor U16260 (N_16260,N_14888,N_15029);
or U16261 (N_16261,N_14339,N_15227);
xor U16262 (N_16262,N_15995,N_15378);
nor U16263 (N_16263,N_15117,N_15394);
and U16264 (N_16264,N_14276,N_15172);
and U16265 (N_16265,N_15585,N_15560);
xor U16266 (N_16266,N_14956,N_14249);
or U16267 (N_16267,N_15398,N_15338);
xnor U16268 (N_16268,N_14554,N_14500);
nor U16269 (N_16269,N_15834,N_14592);
xor U16270 (N_16270,N_14433,N_15134);
nor U16271 (N_16271,N_14124,N_14400);
and U16272 (N_16272,N_14370,N_15699);
nor U16273 (N_16273,N_14665,N_14532);
and U16274 (N_16274,N_14119,N_14991);
xnor U16275 (N_16275,N_14135,N_14020);
xor U16276 (N_16276,N_14138,N_14466);
xnor U16277 (N_16277,N_15618,N_14798);
or U16278 (N_16278,N_15913,N_15712);
nor U16279 (N_16279,N_15792,N_15727);
and U16280 (N_16280,N_15576,N_14252);
xor U16281 (N_16281,N_14189,N_14422);
xor U16282 (N_16282,N_15579,N_15315);
xnor U16283 (N_16283,N_14674,N_15679);
xnor U16284 (N_16284,N_14044,N_15645);
nor U16285 (N_16285,N_14012,N_14484);
nor U16286 (N_16286,N_14254,N_15085);
nor U16287 (N_16287,N_14140,N_14385);
nand U16288 (N_16288,N_15668,N_14601);
xor U16289 (N_16289,N_14470,N_14238);
and U16290 (N_16290,N_15114,N_15132);
or U16291 (N_16291,N_15475,N_14904);
and U16292 (N_16292,N_14143,N_15078);
nor U16293 (N_16293,N_14616,N_15423);
or U16294 (N_16294,N_14190,N_15852);
xnor U16295 (N_16295,N_15539,N_15989);
nand U16296 (N_16296,N_14058,N_14425);
and U16297 (N_16297,N_15743,N_15079);
nor U16298 (N_16298,N_14779,N_15828);
nor U16299 (N_16299,N_14211,N_15957);
xor U16300 (N_16300,N_14504,N_15208);
nor U16301 (N_16301,N_15385,N_15843);
nand U16302 (N_16302,N_15033,N_15241);
nor U16303 (N_16303,N_14122,N_15990);
and U16304 (N_16304,N_15302,N_15249);
and U16305 (N_16305,N_14347,N_15947);
and U16306 (N_16306,N_15627,N_15483);
or U16307 (N_16307,N_15729,N_14244);
nor U16308 (N_16308,N_15299,N_15088);
or U16309 (N_16309,N_15936,N_15929);
xnor U16310 (N_16310,N_15342,N_15789);
xor U16311 (N_16311,N_14610,N_15987);
nor U16312 (N_16312,N_15948,N_15883);
nor U16313 (N_16313,N_14401,N_14558);
and U16314 (N_16314,N_14498,N_14593);
or U16315 (N_16315,N_14688,N_14228);
nand U16316 (N_16316,N_15264,N_14351);
nand U16317 (N_16317,N_14337,N_15049);
nand U16318 (N_16318,N_14277,N_14781);
or U16319 (N_16319,N_14461,N_14127);
nand U16320 (N_16320,N_14421,N_14714);
nor U16321 (N_16321,N_14687,N_15872);
nor U16322 (N_16322,N_14683,N_14950);
nand U16323 (N_16323,N_14099,N_14722);
or U16324 (N_16324,N_15152,N_15454);
or U16325 (N_16325,N_15282,N_14280);
nand U16326 (N_16326,N_15912,N_14229);
xnor U16327 (N_16327,N_15446,N_14754);
nand U16328 (N_16328,N_14985,N_15388);
nor U16329 (N_16329,N_14038,N_15357);
nor U16330 (N_16330,N_15648,N_15972);
xor U16331 (N_16331,N_14494,N_14668);
and U16332 (N_16332,N_15275,N_14656);
or U16333 (N_16333,N_15602,N_15303);
nor U16334 (N_16334,N_15723,N_15415);
xor U16335 (N_16335,N_14786,N_15238);
xor U16336 (N_16336,N_14848,N_14268);
or U16337 (N_16337,N_14534,N_15666);
nor U16338 (N_16338,N_15074,N_15290);
or U16339 (N_16339,N_15996,N_14465);
or U16340 (N_16340,N_15817,N_14450);
nor U16341 (N_16341,N_14710,N_15076);
and U16342 (N_16342,N_15443,N_15893);
nand U16343 (N_16343,N_15364,N_15919);
xnor U16344 (N_16344,N_15753,N_14545);
and U16345 (N_16345,N_15306,N_15746);
nand U16346 (N_16346,N_14513,N_14108);
or U16347 (N_16347,N_15775,N_15949);
and U16348 (N_16348,N_15477,N_15983);
or U16349 (N_16349,N_14894,N_14003);
xnor U16350 (N_16350,N_14900,N_14582);
and U16351 (N_16351,N_14226,N_15934);
and U16352 (N_16352,N_14152,N_15867);
or U16353 (N_16353,N_15322,N_15255);
xnor U16354 (N_16354,N_15284,N_14606);
nand U16355 (N_16355,N_15252,N_14505);
and U16356 (N_16356,N_15642,N_14334);
xnor U16357 (N_16357,N_15921,N_14181);
or U16358 (N_16358,N_15935,N_14954);
nor U16359 (N_16359,N_15151,N_14091);
nor U16360 (N_16360,N_15822,N_15829);
nor U16361 (N_16361,N_15384,N_14557);
and U16362 (N_16362,N_14379,N_14705);
nor U16363 (N_16363,N_14614,N_15226);
xor U16364 (N_16364,N_15115,N_15952);
and U16365 (N_16365,N_14664,N_14538);
and U16366 (N_16366,N_14944,N_15043);
xor U16367 (N_16367,N_15964,N_14937);
nand U16368 (N_16368,N_15399,N_15144);
or U16369 (N_16369,N_14154,N_15205);
nand U16370 (N_16370,N_15331,N_15683);
and U16371 (N_16371,N_14389,N_15927);
nor U16372 (N_16372,N_15213,N_14107);
nor U16373 (N_16373,N_15598,N_14749);
nand U16374 (N_16374,N_15835,N_14928);
xnor U16375 (N_16375,N_14948,N_15096);
and U16376 (N_16376,N_14863,N_15161);
nand U16377 (N_16377,N_14589,N_14731);
nor U16378 (N_16378,N_14799,N_14344);
or U16379 (N_16379,N_14549,N_15016);
nor U16380 (N_16380,N_14671,N_15886);
nand U16381 (N_16381,N_15149,N_15545);
or U16382 (N_16382,N_15370,N_15610);
and U16383 (N_16383,N_15544,N_15736);
or U16384 (N_16384,N_15787,N_15891);
and U16385 (N_16385,N_15622,N_14595);
nand U16386 (N_16386,N_15045,N_14097);
nand U16387 (N_16387,N_15109,N_14784);
xnor U16388 (N_16388,N_14736,N_14889);
or U16389 (N_16389,N_14507,N_14857);
or U16390 (N_16390,N_15769,N_14186);
nand U16391 (N_16391,N_14605,N_14159);
nand U16392 (N_16392,N_15044,N_14711);
nor U16393 (N_16393,N_14253,N_15237);
xnor U16394 (N_16394,N_14745,N_15842);
xnor U16395 (N_16395,N_14407,N_14788);
nand U16396 (N_16396,N_15848,N_14987);
nor U16397 (N_16397,N_14468,N_15766);
and U16398 (N_16398,N_15100,N_14149);
and U16399 (N_16399,N_14133,N_15864);
and U16400 (N_16400,N_14104,N_14571);
xnor U16401 (N_16401,N_14675,N_15809);
xnor U16402 (N_16402,N_14704,N_14471);
nor U16403 (N_16403,N_14919,N_15914);
or U16404 (N_16404,N_15786,N_14312);
nor U16405 (N_16405,N_15099,N_15000);
xor U16406 (N_16406,N_14552,N_15555);
or U16407 (N_16407,N_15687,N_15229);
xor U16408 (N_16408,N_15601,N_15230);
or U16409 (N_16409,N_14488,N_14292);
and U16410 (N_16410,N_15785,N_15234);
or U16411 (N_16411,N_15283,N_15421);
or U16412 (N_16412,N_15962,N_15965);
nor U16413 (N_16413,N_14218,N_14449);
and U16414 (N_16414,N_14809,N_15807);
nor U16415 (N_16415,N_15459,N_15865);
xnor U16416 (N_16416,N_15268,N_14198);
nor U16417 (N_16417,N_15006,N_14916);
xnor U16418 (N_16418,N_15133,N_14896);
nor U16419 (N_16419,N_14188,N_15868);
xnor U16420 (N_16420,N_15571,N_14721);
and U16421 (N_16421,N_15968,N_15471);
xnor U16422 (N_16422,N_15742,N_14903);
nand U16423 (N_16423,N_15136,N_14295);
nor U16424 (N_16424,N_14220,N_14923);
nand U16425 (N_16425,N_15774,N_15667);
and U16426 (N_16426,N_14764,N_14236);
nand U16427 (N_16427,N_14843,N_14369);
or U16428 (N_16428,N_15905,N_14970);
or U16429 (N_16429,N_14497,N_14670);
or U16430 (N_16430,N_15146,N_14783);
and U16431 (N_16431,N_15731,N_14028);
xnor U16432 (N_16432,N_15279,N_14761);
and U16433 (N_16433,N_15963,N_15090);
and U16434 (N_16434,N_14642,N_15280);
and U16435 (N_16435,N_15256,N_14945);
and U16436 (N_16436,N_15281,N_14266);
or U16437 (N_16437,N_15720,N_15212);
or U16438 (N_16438,N_15820,N_14305);
or U16439 (N_16439,N_15247,N_15506);
nand U16440 (N_16440,N_14566,N_14105);
xor U16441 (N_16441,N_15516,N_15073);
nor U16442 (N_16442,N_15140,N_15788);
or U16443 (N_16443,N_15336,N_15387);
nand U16444 (N_16444,N_15899,N_15519);
nand U16445 (N_16445,N_15619,N_14701);
nand U16446 (N_16446,N_15181,N_14611);
or U16447 (N_16447,N_14088,N_14215);
nor U16448 (N_16448,N_14850,N_15243);
or U16449 (N_16449,N_15826,N_14747);
nand U16450 (N_16450,N_15973,N_14780);
nand U16451 (N_16451,N_15107,N_14583);
xnor U16452 (N_16452,N_14070,N_14578);
and U16453 (N_16453,N_14835,N_15402);
or U16454 (N_16454,N_15468,N_15851);
nor U16455 (N_16455,N_15537,N_14390);
nor U16456 (N_16456,N_15609,N_14584);
xnor U16457 (N_16457,N_14459,N_14723);
or U16458 (N_16458,N_15898,N_15209);
nand U16459 (N_16459,N_15546,N_15210);
xnor U16460 (N_16460,N_15672,N_14103);
and U16461 (N_16461,N_14136,N_15456);
nand U16462 (N_16462,N_15450,N_15830);
and U16463 (N_16463,N_14909,N_15574);
xor U16464 (N_16464,N_15232,N_14775);
nand U16465 (N_16465,N_14510,N_15939);
nor U16466 (N_16466,N_15072,N_15669);
nand U16467 (N_16467,N_14367,N_15632);
nor U16468 (N_16468,N_15906,N_15052);
or U16469 (N_16469,N_15304,N_15177);
or U16470 (N_16470,N_14150,N_15013);
and U16471 (N_16471,N_14890,N_15188);
xor U16472 (N_16472,N_14713,N_14810);
and U16473 (N_16473,N_15040,N_15258);
and U16474 (N_16474,N_14076,N_14569);
or U16475 (N_16475,N_15748,N_14338);
nand U16476 (N_16476,N_14838,N_14856);
xnor U16477 (N_16477,N_15624,N_14106);
xor U16478 (N_16478,N_14352,N_15347);
nor U16479 (N_16479,N_15677,N_14682);
xnor U16480 (N_16480,N_15904,N_15162);
and U16481 (N_16481,N_15612,N_14598);
nand U16482 (N_16482,N_14871,N_14817);
and U16483 (N_16483,N_14415,N_14283);
nand U16484 (N_16484,N_14789,N_14223);
xnor U16485 (N_16485,N_14330,N_14353);
nor U16486 (N_16486,N_15933,N_15819);
xor U16487 (N_16487,N_15497,N_15273);
and U16488 (N_16488,N_15647,N_14618);
nor U16489 (N_16489,N_14982,N_15923);
nor U16490 (N_16490,N_14290,N_14316);
and U16491 (N_16491,N_14482,N_15224);
or U16492 (N_16492,N_14591,N_14868);
and U16493 (N_16493,N_15505,N_14998);
and U16494 (N_16494,N_15765,N_15158);
xor U16495 (N_16495,N_14109,N_15691);
and U16496 (N_16496,N_14247,N_14279);
nand U16497 (N_16497,N_15550,N_15464);
nor U16498 (N_16498,N_15321,N_15170);
xnor U16499 (N_16499,N_14270,N_14920);
and U16500 (N_16500,N_14597,N_15488);
or U16501 (N_16501,N_15937,N_15104);
and U16502 (N_16502,N_14004,N_15997);
and U16503 (N_16503,N_14126,N_15661);
xor U16504 (N_16504,N_15308,N_15433);
nand U16505 (N_16505,N_15024,N_15441);
or U16506 (N_16506,N_15944,N_14153);
or U16507 (N_16507,N_15630,N_14550);
and U16508 (N_16508,N_15428,N_15467);
nor U16509 (N_16509,N_14172,N_14184);
and U16510 (N_16510,N_14116,N_14083);
and U16511 (N_16511,N_15616,N_14756);
or U16512 (N_16512,N_15804,N_15671);
nand U16513 (N_16513,N_14199,N_14585);
nor U16514 (N_16514,N_15063,N_15069);
or U16515 (N_16515,N_15419,N_14096);
nor U16516 (N_16516,N_14251,N_15702);
and U16517 (N_16517,N_15548,N_14697);
or U16518 (N_16518,N_14680,N_15296);
nor U16519 (N_16519,N_14773,N_14191);
nand U16520 (N_16520,N_15269,N_15246);
and U16521 (N_16521,N_15902,N_14178);
nand U16522 (N_16522,N_14436,N_14093);
nand U16523 (N_16523,N_14791,N_15285);
nand U16524 (N_16524,N_14411,N_15005);
nand U16525 (N_16525,N_14090,N_14877);
or U16526 (N_16526,N_14445,N_14264);
and U16527 (N_16527,N_15629,N_14897);
or U16528 (N_16528,N_15046,N_15011);
or U16529 (N_16529,N_15439,N_15035);
nor U16530 (N_16530,N_15637,N_15751);
and U16531 (N_16531,N_14168,N_14728);
xnor U16532 (N_16532,N_14205,N_15850);
nor U16533 (N_16533,N_15160,N_15493);
nor U16534 (N_16534,N_14986,N_15316);
nand U16535 (N_16535,N_15713,N_14079);
nand U16536 (N_16536,N_15715,N_15931);
or U16537 (N_16537,N_15489,N_14796);
and U16538 (N_16538,N_14241,N_15490);
nor U16539 (N_16539,N_15673,N_15680);
xnor U16540 (N_16540,N_15692,N_14651);
or U16541 (N_16541,N_15794,N_14968);
nand U16542 (N_16542,N_15190,N_14317);
nor U16543 (N_16543,N_15036,N_14113);
or U16544 (N_16544,N_15623,N_15427);
or U16545 (N_16545,N_14511,N_14366);
nand U16546 (N_16546,N_14170,N_15089);
xor U16547 (N_16547,N_15504,N_15444);
or U16548 (N_16548,N_14148,N_15389);
and U16549 (N_16549,N_15119,N_14045);
or U16550 (N_16550,N_15165,N_15141);
nand U16551 (N_16551,N_15001,N_15846);
nor U16552 (N_16552,N_15187,N_15924);
or U16553 (N_16553,N_15123,N_14363);
and U16554 (N_16554,N_14979,N_14427);
nor U16555 (N_16555,N_14646,N_15910);
or U16556 (N_16556,N_15359,N_14293);
xor U16557 (N_16557,N_15875,N_15540);
or U16558 (N_16558,N_15185,N_15452);
nand U16559 (N_16559,N_14086,N_15696);
or U16560 (N_16560,N_14568,N_14054);
or U16561 (N_16561,N_15652,N_15350);
and U16562 (N_16562,N_14927,N_15193);
nand U16563 (N_16563,N_14464,N_15022);
xnor U16564 (N_16564,N_15845,N_14073);
nor U16565 (N_16565,N_14708,N_15959);
and U16566 (N_16566,N_15633,N_15102);
nor U16567 (N_16567,N_15324,N_15960);
xnor U16568 (N_16568,N_14499,N_14556);
nand U16569 (N_16569,N_15486,N_15026);
or U16570 (N_16570,N_15447,N_14692);
nand U16571 (N_16571,N_15549,N_14426);
or U16572 (N_16572,N_15424,N_15626);
xnor U16573 (N_16573,N_15776,N_15874);
xnor U16574 (N_16574,N_15081,N_15062);
nor U16575 (N_16575,N_14255,N_14924);
and U16576 (N_16576,N_14065,N_15225);
xor U16577 (N_16577,N_14759,N_15453);
or U16578 (N_16578,N_15173,N_15741);
nand U16579 (N_16579,N_15631,N_15724);
xnor U16580 (N_16580,N_15903,N_14524);
nor U16581 (N_16581,N_15403,N_15153);
and U16582 (N_16582,N_14913,N_15176);
and U16583 (N_16583,N_14596,N_14142);
nand U16584 (N_16584,N_15781,N_14469);
nand U16585 (N_16585,N_14514,N_14485);
nand U16586 (N_16586,N_15267,N_14624);
and U16587 (N_16587,N_15353,N_14693);
and U16588 (N_16588,N_15816,N_15344);
and U16589 (N_16589,N_14935,N_15372);
nand U16590 (N_16590,N_15596,N_14960);
nand U16591 (N_16591,N_14673,N_15083);
xor U16592 (N_16592,N_14318,N_14320);
and U16593 (N_16593,N_15217,N_14565);
xnor U16594 (N_16594,N_14643,N_14790);
and U16595 (N_16595,N_15014,N_15526);
and U16596 (N_16596,N_14854,N_14849);
nand U16597 (N_16597,N_15496,N_15199);
nor U16598 (N_16598,N_14032,N_14440);
or U16599 (N_16599,N_15759,N_15966);
or U16600 (N_16600,N_14739,N_14555);
or U16601 (N_16601,N_15745,N_14024);
and U16602 (N_16602,N_15067,N_15061);
nor U16603 (N_16603,N_15380,N_14959);
xor U16604 (N_16604,N_15704,N_15106);
and U16605 (N_16605,N_14120,N_14378);
nand U16606 (N_16606,N_14478,N_14572);
nand U16607 (N_16607,N_15523,N_14805);
nor U16608 (N_16608,N_14221,N_15564);
xor U16609 (N_16609,N_15008,N_14581);
or U16610 (N_16610,N_15220,N_15635);
or U16611 (N_16611,N_14212,N_14489);
and U16612 (N_16612,N_14243,N_15145);
and U16613 (N_16613,N_15265,N_14085);
xnor U16614 (N_16614,N_14101,N_14183);
xor U16615 (N_16615,N_15478,N_15461);
nand U16616 (N_16616,N_14162,N_14239);
nand U16617 (N_16617,N_14139,N_14895);
or U16618 (N_16618,N_14518,N_15430);
nand U16619 (N_16619,N_15839,N_14650);
nor U16620 (N_16620,N_14658,N_15722);
and U16621 (N_16621,N_14362,N_14829);
or U16622 (N_16622,N_14430,N_14298);
xnor U16623 (N_16623,N_14479,N_15348);
or U16624 (N_16624,N_15201,N_14542);
or U16625 (N_16625,N_14388,N_15373);
and U16626 (N_16626,N_14823,N_15010);
or U16627 (N_16627,N_14375,N_15869);
nor U16628 (N_16628,N_15122,N_15659);
xnor U16629 (N_16629,N_14561,N_14026);
nor U16630 (N_16630,N_14011,N_14880);
or U16631 (N_16631,N_14975,N_15750);
xor U16632 (N_16632,N_14263,N_15054);
or U16633 (N_16633,N_15536,N_15686);
nor U16634 (N_16634,N_14516,N_15091);
xnor U16635 (N_16635,N_15251,N_14603);
nand U16636 (N_16636,N_15326,N_15458);
nor U16637 (N_16637,N_14129,N_14902);
xnor U16638 (N_16638,N_15640,N_15940);
nand U16639 (N_16639,N_15391,N_14386);
nand U16640 (N_16640,N_14413,N_14551);
or U16641 (N_16641,N_15581,N_14958);
xor U16642 (N_16642,N_14626,N_15657);
and U16643 (N_16643,N_15460,N_14647);
and U16644 (N_16644,N_14165,N_14125);
and U16645 (N_16645,N_14175,N_15532);
or U16646 (N_16646,N_15039,N_15127);
or U16647 (N_16647,N_15514,N_14684);
xor U16648 (N_16648,N_14969,N_14302);
nor U16649 (N_16649,N_15541,N_15599);
xnor U16650 (N_16650,N_15553,N_14594);
nor U16651 (N_16651,N_14256,N_14077);
or U16652 (N_16652,N_15885,N_14354);
nand U16653 (N_16653,N_14050,N_15928);
nor U16654 (N_16654,N_15700,N_14490);
and U16655 (N_16655,N_15682,N_15552);
nor U16656 (N_16656,N_15871,N_14486);
and U16657 (N_16657,N_14635,N_15007);
or U16658 (N_16658,N_14428,N_14602);
or U16659 (N_16659,N_14995,N_15218);
and U16660 (N_16660,N_14641,N_14887);
or U16661 (N_16661,N_15806,N_15171);
xnor U16662 (N_16662,N_15164,N_15594);
and U16663 (N_16663,N_14918,N_15197);
or U16664 (N_16664,N_15313,N_14022);
nand U16665 (N_16665,N_14027,N_14047);
and U16666 (N_16666,N_15764,N_14429);
and U16667 (N_16667,N_15611,N_15796);
or U16668 (N_16668,N_14893,N_15538);
xnor U16669 (N_16669,N_14526,N_14574);
nor U16670 (N_16670,N_14898,N_14870);
nand U16671 (N_16671,N_15790,N_15266);
and U16672 (N_16672,N_14794,N_14177);
nand U16673 (N_16673,N_15946,N_15508);
xnor U16674 (N_16674,N_15101,N_14176);
and U16675 (N_16675,N_14075,N_15352);
nand U16676 (N_16676,N_14404,N_14147);
or U16677 (N_16677,N_14432,N_14437);
or U16678 (N_16678,N_15844,N_14496);
nand U16679 (N_16679,N_15625,N_15420);
nand U16680 (N_16680,N_15077,N_14052);
or U16681 (N_16681,N_15070,N_15911);
or U16682 (N_16682,N_14633,N_14310);
nor U16683 (N_16683,N_14777,N_15287);
nor U16684 (N_16684,N_14623,N_15805);
nor U16685 (N_16685,N_15194,N_14567);
or U16686 (N_16686,N_15017,N_14064);
nand U16687 (N_16687,N_15561,N_14882);
nand U16688 (N_16688,N_14729,N_15278);
nand U16689 (N_16689,N_14137,N_14066);
or U16690 (N_16690,N_15879,N_14629);
nor U16691 (N_16691,N_14517,N_15849);
nand U16692 (N_16692,N_15050,N_14826);
or U16693 (N_16693,N_15773,N_15941);
nand U16694 (N_16694,N_15897,N_15374);
and U16695 (N_16695,N_14005,N_14448);
or U16696 (N_16696,N_15462,N_14820);
nor U16697 (N_16697,N_15474,N_15600);
nor U16698 (N_16698,N_15501,N_14166);
and U16699 (N_16699,N_15413,N_15970);
nand U16700 (N_16700,N_15412,N_15861);
and U16701 (N_16701,N_14230,N_15529);
or U16702 (N_16702,N_14544,N_14420);
xnor U16703 (N_16703,N_14570,N_14921);
or U16704 (N_16704,N_14579,N_15580);
and U16705 (N_16705,N_15025,N_14141);
nand U16706 (N_16706,N_14717,N_14801);
nand U16707 (N_16707,N_14527,N_14816);
nand U16708 (N_16708,N_15950,N_15312);
and U16709 (N_16709,N_14842,N_14281);
nor U16710 (N_16710,N_15492,N_14331);
nor U16711 (N_16711,N_15047,N_15780);
nand U16712 (N_16712,N_14939,N_15711);
nand U16713 (N_16713,N_15832,N_15297);
nand U16714 (N_16714,N_15747,N_14021);
xor U16715 (N_16715,N_15665,N_15131);
or U16716 (N_16716,N_14586,N_14130);
or U16717 (N_16717,N_15725,N_14912);
xnor U16718 (N_16718,N_15615,N_15057);
nor U16719 (N_16719,N_14772,N_14414);
nand U16720 (N_16720,N_15620,N_15463);
xnor U16721 (N_16721,N_15355,N_15732);
nand U16722 (N_16722,N_14520,N_14967);
or U16723 (N_16723,N_14439,N_14536);
xnor U16724 (N_16724,N_14098,N_15823);
xor U16725 (N_16725,N_15873,N_14069);
or U16726 (N_16726,N_14321,N_15698);
xnor U16727 (N_16727,N_15245,N_15435);
or U16728 (N_16728,N_15656,N_14884);
and U16729 (N_16729,N_14195,N_15333);
or U16730 (N_16730,N_14726,N_15528);
nand U16731 (N_16731,N_14262,N_15137);
and U16732 (N_16732,N_14187,N_15603);
nand U16733 (N_16733,N_14231,N_15472);
and U16734 (N_16734,N_14844,N_14158);
or U16735 (N_16735,N_14456,N_14613);
or U16736 (N_16736,N_14180,N_14358);
and U16737 (N_16737,N_15974,N_14846);
nand U16738 (N_16738,N_15507,N_14669);
nand U16739 (N_16739,N_14299,N_15291);
or U16740 (N_16740,N_15451,N_15059);
and U16741 (N_16741,N_14377,N_15329);
xor U16742 (N_16742,N_14699,N_14000);
xor U16743 (N_16743,N_15437,N_14442);
or U16744 (N_16744,N_14625,N_14462);
nor U16745 (N_16745,N_14503,N_14208);
or U16746 (N_16746,N_15240,N_14952);
or U16747 (N_16747,N_15857,N_15709);
and U16748 (N_16748,N_15808,N_15535);
nor U16749 (N_16749,N_15693,N_14382);
nor U16750 (N_16750,N_15587,N_14246);
or U16751 (N_16751,N_14716,N_14501);
or U16752 (N_16752,N_14811,N_15793);
nor U16753 (N_16753,N_14257,N_14493);
nand U16754 (N_16754,N_15955,N_14818);
xor U16755 (N_16755,N_15744,N_15071);
xor U16756 (N_16756,N_15557,N_15386);
nand U16757 (N_16757,N_15664,N_15135);
xnor U16758 (N_16758,N_15222,N_15925);
xor U16759 (N_16759,N_15154,N_15592);
or U16760 (N_16760,N_14573,N_15381);
or U16761 (N_16761,N_15340,N_14451);
nor U16762 (N_16762,N_15207,N_14762);
xnor U16763 (N_16763,N_14947,N_15125);
or U16764 (N_16764,N_15092,N_15084);
nand U16765 (N_16765,N_15239,N_14371);
and U16766 (N_16766,N_15573,N_14365);
xor U16767 (N_16767,N_14946,N_14908);
nand U16768 (N_16768,N_15813,N_15055);
nand U16769 (N_16769,N_14609,N_14441);
nor U16770 (N_16770,N_15755,N_15638);
or U16771 (N_16771,N_15985,N_14990);
and U16772 (N_16772,N_14548,N_15407);
nor U16773 (N_16773,N_15646,N_14821);
or U16774 (N_16774,N_15042,N_15880);
nand U16775 (N_16775,N_14383,N_14672);
or U16776 (N_16776,N_14063,N_15276);
and U16777 (N_16777,N_14080,N_14173);
or U16778 (N_16778,N_14387,N_14458);
xnor U16779 (N_16779,N_15860,N_14328);
and U16780 (N_16780,N_14615,N_14074);
or U16781 (N_16781,N_14013,N_14803);
nand U16782 (N_16782,N_15901,N_14659);
xnor U16783 (N_16783,N_14528,N_15878);
nand U16784 (N_16784,N_14627,N_14533);
or U16785 (N_16785,N_14914,N_14018);
xor U16786 (N_16786,N_15892,N_15559);
nand U16787 (N_16787,N_15918,N_15818);
nor U16788 (N_16788,N_14855,N_14934);
nor U16789 (N_16789,N_14865,N_14345);
xnor U16790 (N_16790,N_15358,N_14834);
or U16791 (N_16791,N_15147,N_15108);
nor U16792 (N_16792,N_14562,N_15175);
and U16793 (N_16793,N_15288,N_14071);
xnor U16794 (N_16794,N_15651,N_15694);
nor U16795 (N_16795,N_15004,N_15425);
or U16796 (N_16796,N_14434,N_14836);
and U16797 (N_16797,N_15838,N_15888);
nor U16798 (N_16798,N_14906,N_15110);
nor U16799 (N_16799,N_14864,N_15066);
or U16800 (N_16800,N_15383,N_15075);
or U16801 (N_16801,N_15233,N_14667);
and U16802 (N_16802,N_14217,N_15584);
nor U16803 (N_16803,N_15821,N_15644);
and U16804 (N_16804,N_15404,N_15426);
or U16805 (N_16805,N_15377,N_14406);
nand U16806 (N_16806,N_14495,N_15476);
nand U16807 (N_16807,N_15980,N_14828);
xor U16808 (N_16808,N_15150,N_15613);
or U16809 (N_16809,N_15998,N_14059);
xor U16810 (N_16810,N_14355,N_14261);
nor U16811 (N_16811,N_15351,N_15908);
and U16812 (N_16812,N_14977,N_15491);
or U16813 (N_16813,N_15595,N_14477);
nand U16814 (N_16814,N_14802,N_14222);
xnor U16815 (N_16815,N_14640,N_15457);
xor U16816 (N_16816,N_15037,N_15179);
xor U16817 (N_16817,N_14907,N_15363);
nor U16818 (N_16818,N_14653,N_15392);
nand U16819 (N_16819,N_15798,N_15678);
and U16820 (N_16820,N_15270,N_15118);
xnor U16821 (N_16821,N_14315,N_14876);
xnor U16822 (N_16822,N_15650,N_15116);
xnor U16823 (N_16823,N_15445,N_14793);
nor U16824 (N_16824,N_14067,N_15120);
xnor U16825 (N_16825,N_14930,N_14200);
or U16826 (N_16826,N_14100,N_14237);
and U16827 (N_16827,N_14210,N_14620);
xnor U16828 (N_16828,N_15649,N_14654);
or U16829 (N_16829,N_15030,N_15221);
xnor U16830 (N_16830,N_15597,N_14546);
and U16831 (N_16831,N_15812,N_15068);
and U16832 (N_16832,N_15368,N_15737);
xnor U16833 (N_16833,N_14311,N_15556);
nor U16834 (N_16834,N_14506,N_15390);
and U16835 (N_16835,N_14395,N_14883);
nand U16836 (N_16836,N_15690,N_14155);
and U16837 (N_16837,N_15831,N_15440);
and U16838 (N_16838,N_15481,N_15021);
nor U16839 (N_16839,N_14825,N_15825);
xnor U16840 (N_16840,N_15588,N_15003);
xor U16841 (N_16841,N_14663,N_14765);
xor U16842 (N_16842,N_14403,N_14332);
nor U16843 (N_16843,N_15922,N_15155);
nor U16844 (N_16844,N_15771,N_15525);
xor U16845 (N_16845,N_15248,N_15994);
nor U16846 (N_16846,N_15763,N_15517);
nor U16847 (N_16847,N_14117,N_15480);
nor U16848 (N_16848,N_14258,N_14463);
or U16849 (N_16849,N_15369,N_14649);
nor U16850 (N_16850,N_14297,N_15734);
nand U16851 (N_16851,N_14235,N_15858);
nor U16852 (N_16852,N_14806,N_14724);
nand U16853 (N_16853,N_14289,N_15993);
xnor U16854 (N_16854,N_15409,N_15986);
nor U16855 (N_16855,N_14755,N_14966);
nor U16856 (N_16856,N_14737,N_14095);
and U16857 (N_16857,N_14014,N_14932);
xnor U16858 (N_16858,N_14964,N_15706);
nor U16859 (N_16859,N_14209,N_14340);
xnor U16860 (N_16860,N_14676,N_14787);
nor U16861 (N_16861,N_14707,N_15080);
xor U16862 (N_16862,N_15126,N_15356);
and U16863 (N_16863,N_15614,N_15674);
and U16864 (N_16864,N_15032,N_15455);
nor U16865 (N_16865,N_15982,N_14481);
xnor U16866 (N_16866,N_14272,N_14875);
or U16867 (N_16867,N_15186,N_14055);
nor U16868 (N_16868,N_15411,N_14797);
nand U16869 (N_16869,N_15200,N_14951);
xnor U16870 (N_16870,N_15499,N_15335);
or U16871 (N_16871,N_14009,N_15660);
xnor U16872 (N_16872,N_14522,N_15442);
or U16873 (N_16873,N_15310,N_14278);
xor U16874 (N_16874,N_15484,N_15018);
or U16875 (N_16875,N_15341,N_15184);
nor U16876 (N_16876,N_14010,N_15367);
and U16877 (N_16877,N_14677,N_14822);
or U16878 (N_16878,N_14509,N_15621);
or U16879 (N_16879,N_14752,N_14925);
or U16880 (N_16880,N_14157,N_15701);
and U16881 (N_16881,N_14483,N_14971);
or U16882 (N_16882,N_15710,N_15782);
and U16883 (N_16883,N_14274,N_14111);
xor U16884 (N_16884,N_15969,N_14837);
nand U16885 (N_16885,N_14873,N_15400);
nor U16886 (N_16886,N_15139,N_14294);
xnor U16887 (N_16887,N_15577,N_14041);
xor U16888 (N_16888,N_14732,N_15515);
nand U16889 (N_16889,N_15558,N_14696);
nand U16890 (N_16890,N_15271,N_15511);
or U16891 (N_16891,N_15942,N_15572);
xor U16892 (N_16892,N_14444,N_15795);
or U16893 (N_16893,N_15178,N_14698);
xor U16894 (N_16894,N_15547,N_14981);
or U16895 (N_16895,N_15841,N_15431);
or U16896 (N_16896,N_15738,N_14273);
nand U16897 (N_16897,N_14525,N_14329);
xnor U16898 (N_16898,N_14929,N_14350);
xor U16899 (N_16899,N_15827,N_15735);
or U16900 (N_16900,N_14373,N_15298);
nor U16901 (N_16901,N_14800,N_14282);
xnor U16902 (N_16902,N_15289,N_14452);
and U16903 (N_16903,N_15328,N_15048);
xor U16904 (N_16904,N_14936,N_15157);
xor U16905 (N_16905,N_14410,N_14750);
nand U16906 (N_16906,N_15214,N_14288);
nor U16907 (N_16907,N_14326,N_14866);
nor U16908 (N_16908,N_15223,N_15482);
nand U16909 (N_16909,N_15469,N_15762);
nand U16910 (N_16910,N_15565,N_14695);
nand U16911 (N_16911,N_14941,N_14530);
xor U16912 (N_16912,N_15814,N_15887);
xnor U16913 (N_16913,N_14476,N_14225);
nand U16914 (N_16914,N_14356,N_14474);
or U16915 (N_16915,N_14453,N_15707);
xnor U16916 (N_16916,N_15500,N_14785);
nor U16917 (N_16917,N_15082,N_14372);
nor U16918 (N_16918,N_15343,N_14619);
nor U16919 (N_16919,N_14193,N_15023);
nand U16920 (N_16920,N_15495,N_14392);
xnor U16921 (N_16921,N_14206,N_14993);
nor U16922 (N_16922,N_14839,N_15643);
or U16923 (N_16923,N_15799,N_14771);
nand U16924 (N_16924,N_14156,N_15976);
or U16925 (N_16925,N_14480,N_15512);
nand U16926 (N_16926,N_15410,N_15907);
and U16927 (N_16927,N_14250,N_14812);
or U16928 (N_16928,N_14016,N_15531);
nor U16929 (N_16929,N_15405,N_15663);
xor U16930 (N_16930,N_14042,N_14678);
and U16931 (N_16931,N_15260,N_14891);
nand U16932 (N_16932,N_15124,N_14621);
and U16933 (N_16933,N_14735,N_14767);
xor U16934 (N_16934,N_15527,N_15448);
and U16935 (N_16935,N_15589,N_14368);
nand U16936 (N_16936,N_15327,N_15375);
nor U16937 (N_16937,N_15752,N_14046);
nor U16938 (N_16938,N_14899,N_14275);
xor U16939 (N_16939,N_14034,N_15053);
xnor U16940 (N_16940,N_14720,N_15236);
nand U16941 (N_16941,N_14435,N_14308);
nand U16942 (N_16942,N_14197,N_14219);
and U16943 (N_16943,N_14265,N_15436);
xor U16944 (N_16944,N_15345,N_15323);
nand U16945 (N_16945,N_15509,N_15566);
nand U16946 (N_16946,N_14962,N_14955);
nand U16947 (N_16947,N_15262,N_15636);
and U16948 (N_16948,N_15166,N_15235);
nand U16949 (N_16949,N_14037,N_14115);
nor U16950 (N_16950,N_14861,N_15655);
xnor U16951 (N_16951,N_15211,N_14144);
and U16952 (N_16952,N_14813,N_15953);
and U16953 (N_16953,N_15272,N_15473);
nor U16954 (N_16954,N_14963,N_14019);
and U16955 (N_16955,N_14885,N_14575);
xnor U16956 (N_16956,N_15169,N_14862);
nor U16957 (N_16957,N_15884,N_15703);
nand U16958 (N_16958,N_14679,N_15416);
and U16959 (N_16959,N_14719,N_14128);
or U16960 (N_16960,N_15111,N_15810);
or U16961 (N_16961,N_14686,N_15777);
nand U16962 (N_16962,N_14763,N_14349);
or U16963 (N_16963,N_14734,N_14145);
xor U16964 (N_16964,N_15292,N_15259);
or U16965 (N_16965,N_15754,N_14017);
xor U16966 (N_16966,N_15366,N_14447);
xnor U16967 (N_16967,N_14766,N_15103);
nand U16968 (N_16968,N_14060,N_14391);
and U16969 (N_16969,N_14694,N_14374);
xor U16970 (N_16970,N_15930,N_14049);
xnor U16971 (N_16971,N_15840,N_15916);
nor U16972 (N_16972,N_14438,N_15093);
nand U16973 (N_16973,N_15896,N_14874);
nand U16974 (N_16974,N_15064,N_14983);
and U16975 (N_16975,N_15606,N_14036);
or U16976 (N_16976,N_14521,N_15180);
xnor U16977 (N_16977,N_15113,N_15034);
nor U16978 (N_16978,N_15206,N_15681);
and U16979 (N_16979,N_14700,N_14815);
or U16980 (N_16980,N_14757,N_15836);
nand U16981 (N_16981,N_14114,N_15961);
or U16982 (N_16982,N_15670,N_14213);
and U16983 (N_16983,N_15337,N_14892);
xor U16984 (N_16984,N_15772,N_14419);
xnor U16985 (N_16985,N_15628,N_14163);
or U16986 (N_16986,N_15012,N_14467);
xnor U16987 (N_16987,N_14007,N_15604);
or U16988 (N_16988,N_14859,N_15778);
or U16989 (N_16989,N_14259,N_15563);
and U16990 (N_16990,N_14770,N_14860);
or U16991 (N_16991,N_15783,N_15174);
nor U16992 (N_16992,N_15105,N_15578);
nor U16993 (N_16993,N_14245,N_14164);
nor U16994 (N_16994,N_15438,N_14457);
xnor U16995 (N_16995,N_14577,N_14327);
nor U16996 (N_16996,N_14703,N_14473);
nand U16997 (N_16997,N_15697,N_14393);
nor U16998 (N_16998,N_15379,N_14306);
nor U16999 (N_16999,N_14160,N_14240);
xnor U17000 (N_17000,N_15447,N_15576);
nor U17001 (N_17001,N_14590,N_15058);
nand U17002 (N_17002,N_15304,N_15114);
nor U17003 (N_17003,N_14848,N_14485);
nand U17004 (N_17004,N_14012,N_14811);
or U17005 (N_17005,N_14943,N_15197);
or U17006 (N_17006,N_14566,N_15381);
xor U17007 (N_17007,N_15731,N_14613);
and U17008 (N_17008,N_15685,N_14508);
nand U17009 (N_17009,N_14544,N_14309);
and U17010 (N_17010,N_15731,N_15702);
and U17011 (N_17011,N_15104,N_15315);
or U17012 (N_17012,N_15850,N_14874);
nor U17013 (N_17013,N_15202,N_14116);
nand U17014 (N_17014,N_14265,N_15688);
nand U17015 (N_17015,N_15097,N_14042);
or U17016 (N_17016,N_14712,N_15827);
nor U17017 (N_17017,N_14956,N_14751);
xor U17018 (N_17018,N_14887,N_15862);
nand U17019 (N_17019,N_14159,N_14375);
and U17020 (N_17020,N_15069,N_14498);
and U17021 (N_17021,N_15036,N_14753);
xnor U17022 (N_17022,N_14623,N_15133);
xnor U17023 (N_17023,N_14594,N_14052);
and U17024 (N_17024,N_14032,N_15392);
nor U17025 (N_17025,N_15666,N_15044);
nand U17026 (N_17026,N_15029,N_15607);
nand U17027 (N_17027,N_15902,N_14675);
xnor U17028 (N_17028,N_14594,N_15780);
and U17029 (N_17029,N_15653,N_14539);
or U17030 (N_17030,N_15975,N_15141);
xnor U17031 (N_17031,N_14456,N_14769);
nor U17032 (N_17032,N_14225,N_14141);
xor U17033 (N_17033,N_14598,N_14049);
and U17034 (N_17034,N_15233,N_15546);
or U17035 (N_17035,N_14040,N_15775);
or U17036 (N_17036,N_15677,N_15649);
or U17037 (N_17037,N_15432,N_15988);
xnor U17038 (N_17038,N_15406,N_14267);
xnor U17039 (N_17039,N_15955,N_14808);
nor U17040 (N_17040,N_14525,N_15737);
xnor U17041 (N_17041,N_14196,N_15780);
nor U17042 (N_17042,N_15839,N_14222);
or U17043 (N_17043,N_14644,N_15634);
or U17044 (N_17044,N_15410,N_14549);
or U17045 (N_17045,N_15842,N_15022);
nand U17046 (N_17046,N_14330,N_14675);
nor U17047 (N_17047,N_14820,N_15220);
or U17048 (N_17048,N_15562,N_14049);
nand U17049 (N_17049,N_14586,N_14335);
nand U17050 (N_17050,N_15648,N_15094);
and U17051 (N_17051,N_14381,N_15305);
nand U17052 (N_17052,N_14061,N_14416);
and U17053 (N_17053,N_15241,N_15016);
nor U17054 (N_17054,N_15580,N_14951);
xnor U17055 (N_17055,N_15898,N_15144);
nand U17056 (N_17056,N_15539,N_15688);
and U17057 (N_17057,N_15673,N_15565);
nor U17058 (N_17058,N_14956,N_15016);
and U17059 (N_17059,N_15969,N_15743);
nand U17060 (N_17060,N_14860,N_15813);
xor U17061 (N_17061,N_14925,N_14349);
nand U17062 (N_17062,N_15971,N_15605);
xor U17063 (N_17063,N_15385,N_15107);
nand U17064 (N_17064,N_15957,N_15746);
or U17065 (N_17065,N_15471,N_15422);
or U17066 (N_17066,N_15106,N_15782);
nand U17067 (N_17067,N_15810,N_14185);
or U17068 (N_17068,N_14230,N_15757);
nand U17069 (N_17069,N_14777,N_14631);
xor U17070 (N_17070,N_15246,N_14838);
nor U17071 (N_17071,N_14854,N_14801);
and U17072 (N_17072,N_15660,N_15141);
nor U17073 (N_17073,N_15428,N_14361);
nand U17074 (N_17074,N_15323,N_15392);
xor U17075 (N_17075,N_14752,N_15838);
and U17076 (N_17076,N_14166,N_14442);
or U17077 (N_17077,N_15028,N_14209);
nor U17078 (N_17078,N_15200,N_15838);
or U17079 (N_17079,N_14915,N_15429);
nor U17080 (N_17080,N_15602,N_15656);
xnor U17081 (N_17081,N_14257,N_15096);
and U17082 (N_17082,N_14803,N_15689);
nand U17083 (N_17083,N_14518,N_15911);
nand U17084 (N_17084,N_15293,N_15640);
xor U17085 (N_17085,N_14114,N_14478);
or U17086 (N_17086,N_15237,N_15886);
xor U17087 (N_17087,N_14821,N_14691);
nand U17088 (N_17088,N_14713,N_14296);
or U17089 (N_17089,N_14621,N_14537);
or U17090 (N_17090,N_15877,N_15156);
xor U17091 (N_17091,N_14626,N_14341);
and U17092 (N_17092,N_15817,N_14559);
xor U17093 (N_17093,N_15580,N_15837);
and U17094 (N_17094,N_14973,N_14410);
nor U17095 (N_17095,N_14148,N_15868);
and U17096 (N_17096,N_14035,N_14857);
xor U17097 (N_17097,N_15089,N_15153);
and U17098 (N_17098,N_14168,N_14143);
and U17099 (N_17099,N_14751,N_14824);
nor U17100 (N_17100,N_14280,N_14133);
and U17101 (N_17101,N_15816,N_14363);
and U17102 (N_17102,N_15057,N_14456);
and U17103 (N_17103,N_15617,N_15405);
and U17104 (N_17104,N_15942,N_14090);
xor U17105 (N_17105,N_15785,N_14778);
and U17106 (N_17106,N_15450,N_14764);
xnor U17107 (N_17107,N_14296,N_14143);
xor U17108 (N_17108,N_15068,N_14379);
nand U17109 (N_17109,N_14220,N_14262);
nor U17110 (N_17110,N_14754,N_14566);
and U17111 (N_17111,N_14703,N_14287);
nand U17112 (N_17112,N_15285,N_14337);
and U17113 (N_17113,N_15812,N_15211);
and U17114 (N_17114,N_15033,N_14624);
nand U17115 (N_17115,N_15604,N_14295);
nand U17116 (N_17116,N_14643,N_14807);
nand U17117 (N_17117,N_15845,N_15448);
nand U17118 (N_17118,N_14589,N_15243);
xor U17119 (N_17119,N_14779,N_15581);
nor U17120 (N_17120,N_15545,N_15357);
nand U17121 (N_17121,N_15701,N_15765);
or U17122 (N_17122,N_14958,N_15314);
nor U17123 (N_17123,N_15937,N_15725);
nor U17124 (N_17124,N_14669,N_14128);
xor U17125 (N_17125,N_14575,N_15131);
nand U17126 (N_17126,N_15193,N_14970);
and U17127 (N_17127,N_15207,N_15096);
nor U17128 (N_17128,N_14222,N_15775);
nand U17129 (N_17129,N_14097,N_14959);
xnor U17130 (N_17130,N_14186,N_14243);
xor U17131 (N_17131,N_15128,N_14808);
xnor U17132 (N_17132,N_14772,N_15567);
xor U17133 (N_17133,N_14083,N_15751);
nand U17134 (N_17134,N_15070,N_15121);
or U17135 (N_17135,N_15416,N_15253);
nor U17136 (N_17136,N_14414,N_14436);
nor U17137 (N_17137,N_14396,N_14423);
nor U17138 (N_17138,N_14713,N_15054);
nand U17139 (N_17139,N_15131,N_14756);
or U17140 (N_17140,N_14755,N_15573);
or U17141 (N_17141,N_15529,N_14402);
or U17142 (N_17142,N_14858,N_15473);
and U17143 (N_17143,N_15109,N_14203);
nand U17144 (N_17144,N_15111,N_14573);
or U17145 (N_17145,N_14090,N_15560);
and U17146 (N_17146,N_15184,N_14518);
nand U17147 (N_17147,N_15158,N_15467);
nand U17148 (N_17148,N_15619,N_14843);
and U17149 (N_17149,N_14046,N_14215);
nor U17150 (N_17150,N_14567,N_15235);
or U17151 (N_17151,N_15993,N_14012);
or U17152 (N_17152,N_14481,N_15127);
or U17153 (N_17153,N_14032,N_15608);
or U17154 (N_17154,N_15643,N_14274);
nor U17155 (N_17155,N_14589,N_14061);
xnor U17156 (N_17156,N_15582,N_14975);
nand U17157 (N_17157,N_14743,N_15294);
nand U17158 (N_17158,N_15387,N_14603);
xor U17159 (N_17159,N_14468,N_14510);
nor U17160 (N_17160,N_14586,N_14860);
nand U17161 (N_17161,N_14143,N_14486);
nand U17162 (N_17162,N_15343,N_15480);
nor U17163 (N_17163,N_15593,N_15386);
xnor U17164 (N_17164,N_14277,N_14942);
or U17165 (N_17165,N_14990,N_15725);
nor U17166 (N_17166,N_14108,N_14674);
and U17167 (N_17167,N_14938,N_14149);
nor U17168 (N_17168,N_14442,N_14981);
and U17169 (N_17169,N_14581,N_15980);
nor U17170 (N_17170,N_14625,N_15170);
or U17171 (N_17171,N_15805,N_15336);
and U17172 (N_17172,N_14915,N_14119);
nand U17173 (N_17173,N_15964,N_14370);
or U17174 (N_17174,N_14573,N_14699);
or U17175 (N_17175,N_15988,N_15213);
xnor U17176 (N_17176,N_14844,N_14381);
xor U17177 (N_17177,N_15335,N_14323);
nand U17178 (N_17178,N_14779,N_14949);
nor U17179 (N_17179,N_15708,N_15863);
nand U17180 (N_17180,N_15602,N_15598);
nor U17181 (N_17181,N_14019,N_15202);
and U17182 (N_17182,N_15776,N_14425);
nand U17183 (N_17183,N_15922,N_15006);
or U17184 (N_17184,N_14726,N_15843);
or U17185 (N_17185,N_14939,N_14864);
xnor U17186 (N_17186,N_14010,N_14899);
and U17187 (N_17187,N_15594,N_14796);
nor U17188 (N_17188,N_15867,N_14781);
nand U17189 (N_17189,N_14175,N_15753);
or U17190 (N_17190,N_14299,N_14499);
and U17191 (N_17191,N_15282,N_15893);
or U17192 (N_17192,N_14589,N_14728);
nor U17193 (N_17193,N_15361,N_14901);
xnor U17194 (N_17194,N_14649,N_15361);
and U17195 (N_17195,N_15920,N_14331);
nand U17196 (N_17196,N_14574,N_15029);
xor U17197 (N_17197,N_15452,N_15896);
nand U17198 (N_17198,N_14267,N_15766);
or U17199 (N_17199,N_15930,N_15826);
nor U17200 (N_17200,N_14129,N_15514);
and U17201 (N_17201,N_14025,N_15152);
or U17202 (N_17202,N_14185,N_15411);
or U17203 (N_17203,N_14487,N_14441);
nor U17204 (N_17204,N_14479,N_14107);
and U17205 (N_17205,N_14977,N_14598);
nand U17206 (N_17206,N_14064,N_14756);
xnor U17207 (N_17207,N_14757,N_14405);
nand U17208 (N_17208,N_15530,N_14555);
and U17209 (N_17209,N_15774,N_14199);
nand U17210 (N_17210,N_14327,N_14403);
xnor U17211 (N_17211,N_14298,N_15061);
nor U17212 (N_17212,N_15240,N_14682);
nand U17213 (N_17213,N_14088,N_15932);
nor U17214 (N_17214,N_14438,N_14119);
and U17215 (N_17215,N_14847,N_14686);
nand U17216 (N_17216,N_15323,N_15962);
nor U17217 (N_17217,N_15933,N_15813);
and U17218 (N_17218,N_15140,N_14653);
nand U17219 (N_17219,N_15074,N_14043);
and U17220 (N_17220,N_15052,N_15740);
xnor U17221 (N_17221,N_15778,N_15717);
nor U17222 (N_17222,N_15208,N_14097);
and U17223 (N_17223,N_14185,N_15429);
nor U17224 (N_17224,N_14490,N_14647);
xnor U17225 (N_17225,N_14501,N_14190);
nand U17226 (N_17226,N_15216,N_15555);
and U17227 (N_17227,N_15062,N_14458);
nand U17228 (N_17228,N_15074,N_14081);
xor U17229 (N_17229,N_15257,N_15924);
nor U17230 (N_17230,N_14335,N_14352);
or U17231 (N_17231,N_14555,N_15326);
nand U17232 (N_17232,N_14381,N_15721);
and U17233 (N_17233,N_14875,N_15094);
xnor U17234 (N_17234,N_15559,N_14037);
and U17235 (N_17235,N_15673,N_15457);
nand U17236 (N_17236,N_14528,N_14666);
or U17237 (N_17237,N_15017,N_15627);
nor U17238 (N_17238,N_14490,N_15694);
nor U17239 (N_17239,N_14882,N_14260);
nor U17240 (N_17240,N_14855,N_15247);
nor U17241 (N_17241,N_15525,N_14470);
and U17242 (N_17242,N_14882,N_14108);
xnor U17243 (N_17243,N_15582,N_15977);
nand U17244 (N_17244,N_14094,N_14372);
or U17245 (N_17245,N_15237,N_15445);
and U17246 (N_17246,N_15446,N_15286);
xnor U17247 (N_17247,N_14438,N_14550);
nand U17248 (N_17248,N_15527,N_15659);
nor U17249 (N_17249,N_15870,N_14114);
and U17250 (N_17250,N_14246,N_14868);
xnor U17251 (N_17251,N_15419,N_14022);
nor U17252 (N_17252,N_14032,N_14104);
nor U17253 (N_17253,N_14372,N_14663);
nand U17254 (N_17254,N_15488,N_14590);
nor U17255 (N_17255,N_15561,N_14071);
xor U17256 (N_17256,N_15251,N_15875);
nor U17257 (N_17257,N_14574,N_15341);
nand U17258 (N_17258,N_15243,N_15296);
or U17259 (N_17259,N_14546,N_15660);
or U17260 (N_17260,N_15726,N_14886);
and U17261 (N_17261,N_14645,N_15294);
and U17262 (N_17262,N_14205,N_15318);
and U17263 (N_17263,N_14044,N_15362);
nor U17264 (N_17264,N_14614,N_14148);
xor U17265 (N_17265,N_14366,N_15754);
and U17266 (N_17266,N_15064,N_14417);
nand U17267 (N_17267,N_15732,N_15477);
or U17268 (N_17268,N_15317,N_14033);
nand U17269 (N_17269,N_15289,N_14553);
and U17270 (N_17270,N_14760,N_14948);
nor U17271 (N_17271,N_15991,N_15881);
xnor U17272 (N_17272,N_14588,N_14532);
or U17273 (N_17273,N_14860,N_15529);
nand U17274 (N_17274,N_15579,N_14900);
or U17275 (N_17275,N_14764,N_15433);
nor U17276 (N_17276,N_15453,N_14766);
nand U17277 (N_17277,N_14948,N_15173);
and U17278 (N_17278,N_15894,N_15564);
and U17279 (N_17279,N_14721,N_15129);
and U17280 (N_17280,N_15082,N_15784);
nand U17281 (N_17281,N_14528,N_14600);
and U17282 (N_17282,N_14061,N_15707);
or U17283 (N_17283,N_14310,N_14470);
and U17284 (N_17284,N_15246,N_14357);
nand U17285 (N_17285,N_15626,N_15904);
xnor U17286 (N_17286,N_15670,N_15188);
nor U17287 (N_17287,N_14997,N_14139);
nand U17288 (N_17288,N_14046,N_14628);
nand U17289 (N_17289,N_15358,N_14145);
nand U17290 (N_17290,N_14142,N_14592);
or U17291 (N_17291,N_15561,N_15422);
xor U17292 (N_17292,N_15431,N_15605);
and U17293 (N_17293,N_14354,N_14414);
nor U17294 (N_17294,N_14780,N_14991);
and U17295 (N_17295,N_15439,N_15644);
or U17296 (N_17296,N_15246,N_15265);
nand U17297 (N_17297,N_14562,N_15418);
nor U17298 (N_17298,N_15148,N_15338);
nand U17299 (N_17299,N_14924,N_14516);
or U17300 (N_17300,N_14199,N_15588);
nand U17301 (N_17301,N_14995,N_15339);
nor U17302 (N_17302,N_15636,N_15682);
xnor U17303 (N_17303,N_14119,N_14444);
and U17304 (N_17304,N_14181,N_15128);
nand U17305 (N_17305,N_14580,N_14125);
or U17306 (N_17306,N_14822,N_14201);
or U17307 (N_17307,N_15597,N_15857);
or U17308 (N_17308,N_14274,N_14748);
nor U17309 (N_17309,N_14804,N_15971);
nor U17310 (N_17310,N_15542,N_14716);
nand U17311 (N_17311,N_15362,N_15126);
xor U17312 (N_17312,N_14643,N_15373);
or U17313 (N_17313,N_14493,N_15010);
and U17314 (N_17314,N_14221,N_15087);
nand U17315 (N_17315,N_14010,N_14041);
and U17316 (N_17316,N_15172,N_14078);
and U17317 (N_17317,N_15515,N_15289);
and U17318 (N_17318,N_15802,N_15060);
nor U17319 (N_17319,N_15742,N_15646);
or U17320 (N_17320,N_14278,N_15766);
or U17321 (N_17321,N_14869,N_15570);
nand U17322 (N_17322,N_15949,N_14133);
nand U17323 (N_17323,N_15002,N_15799);
nor U17324 (N_17324,N_15967,N_15623);
nand U17325 (N_17325,N_15512,N_14632);
or U17326 (N_17326,N_14383,N_15558);
and U17327 (N_17327,N_15355,N_15873);
or U17328 (N_17328,N_14272,N_14334);
xnor U17329 (N_17329,N_14472,N_15876);
xor U17330 (N_17330,N_15456,N_14885);
xnor U17331 (N_17331,N_14641,N_15898);
or U17332 (N_17332,N_15343,N_15556);
and U17333 (N_17333,N_15613,N_15412);
nand U17334 (N_17334,N_15571,N_15835);
xor U17335 (N_17335,N_15964,N_14489);
or U17336 (N_17336,N_15613,N_14432);
xnor U17337 (N_17337,N_15487,N_15990);
or U17338 (N_17338,N_15435,N_14523);
and U17339 (N_17339,N_14651,N_14658);
xnor U17340 (N_17340,N_15575,N_15050);
or U17341 (N_17341,N_14268,N_15926);
nor U17342 (N_17342,N_15781,N_14294);
nor U17343 (N_17343,N_14006,N_15893);
nand U17344 (N_17344,N_14768,N_15227);
and U17345 (N_17345,N_14241,N_15763);
nor U17346 (N_17346,N_15196,N_15675);
or U17347 (N_17347,N_14052,N_15008);
nor U17348 (N_17348,N_15413,N_14660);
nand U17349 (N_17349,N_14096,N_15945);
and U17350 (N_17350,N_15840,N_15027);
or U17351 (N_17351,N_14771,N_15428);
nand U17352 (N_17352,N_14337,N_14713);
and U17353 (N_17353,N_14994,N_15261);
nor U17354 (N_17354,N_15703,N_15623);
xnor U17355 (N_17355,N_15701,N_14193);
or U17356 (N_17356,N_14399,N_15096);
nor U17357 (N_17357,N_15218,N_14206);
or U17358 (N_17358,N_15324,N_14254);
or U17359 (N_17359,N_15233,N_14163);
nand U17360 (N_17360,N_14961,N_15928);
and U17361 (N_17361,N_14620,N_15858);
xnor U17362 (N_17362,N_14561,N_14713);
nand U17363 (N_17363,N_14443,N_15651);
xnor U17364 (N_17364,N_14995,N_15588);
nor U17365 (N_17365,N_14234,N_15403);
xnor U17366 (N_17366,N_15832,N_14351);
nand U17367 (N_17367,N_15848,N_14641);
xnor U17368 (N_17368,N_15981,N_14478);
nand U17369 (N_17369,N_14325,N_14664);
nand U17370 (N_17370,N_14987,N_15752);
nand U17371 (N_17371,N_15358,N_15437);
nand U17372 (N_17372,N_15229,N_14463);
or U17373 (N_17373,N_15491,N_14832);
and U17374 (N_17374,N_14255,N_15770);
nand U17375 (N_17375,N_14432,N_15132);
or U17376 (N_17376,N_15981,N_15866);
nor U17377 (N_17377,N_15376,N_15750);
and U17378 (N_17378,N_14824,N_14450);
nand U17379 (N_17379,N_15656,N_15286);
or U17380 (N_17380,N_15406,N_14107);
and U17381 (N_17381,N_14408,N_15617);
xnor U17382 (N_17382,N_14550,N_14035);
and U17383 (N_17383,N_15461,N_15097);
and U17384 (N_17384,N_14777,N_14244);
and U17385 (N_17385,N_15408,N_15623);
nor U17386 (N_17386,N_14907,N_15831);
nand U17387 (N_17387,N_15666,N_14758);
nor U17388 (N_17388,N_15182,N_15295);
nand U17389 (N_17389,N_15507,N_15343);
nor U17390 (N_17390,N_14438,N_14455);
and U17391 (N_17391,N_15198,N_15599);
or U17392 (N_17392,N_14174,N_14638);
or U17393 (N_17393,N_14645,N_14654);
xnor U17394 (N_17394,N_14541,N_14828);
and U17395 (N_17395,N_14129,N_14816);
or U17396 (N_17396,N_15592,N_14823);
and U17397 (N_17397,N_15897,N_14966);
and U17398 (N_17398,N_14124,N_15342);
nor U17399 (N_17399,N_15723,N_15627);
or U17400 (N_17400,N_14692,N_14484);
xnor U17401 (N_17401,N_15409,N_15059);
or U17402 (N_17402,N_14774,N_15199);
nand U17403 (N_17403,N_14766,N_15555);
nor U17404 (N_17404,N_14065,N_14596);
xor U17405 (N_17405,N_15238,N_15251);
and U17406 (N_17406,N_14843,N_15060);
or U17407 (N_17407,N_15081,N_14464);
xor U17408 (N_17408,N_14971,N_15879);
nor U17409 (N_17409,N_14640,N_15477);
nand U17410 (N_17410,N_14416,N_15054);
nand U17411 (N_17411,N_15122,N_14195);
and U17412 (N_17412,N_14548,N_14526);
nor U17413 (N_17413,N_15627,N_14969);
nor U17414 (N_17414,N_15271,N_14678);
xnor U17415 (N_17415,N_15899,N_15975);
xnor U17416 (N_17416,N_14529,N_14772);
xor U17417 (N_17417,N_15341,N_14023);
or U17418 (N_17418,N_15730,N_15674);
and U17419 (N_17419,N_14127,N_15186);
xor U17420 (N_17420,N_14274,N_14577);
or U17421 (N_17421,N_14182,N_15147);
nand U17422 (N_17422,N_15779,N_14840);
or U17423 (N_17423,N_15182,N_14165);
xnor U17424 (N_17424,N_14648,N_15025);
nand U17425 (N_17425,N_15546,N_14120);
nand U17426 (N_17426,N_15078,N_15727);
xnor U17427 (N_17427,N_15959,N_14201);
nor U17428 (N_17428,N_14622,N_15725);
xor U17429 (N_17429,N_15674,N_15321);
and U17430 (N_17430,N_15793,N_15882);
or U17431 (N_17431,N_15316,N_15357);
and U17432 (N_17432,N_14846,N_15291);
xnor U17433 (N_17433,N_14475,N_14925);
and U17434 (N_17434,N_14971,N_15620);
and U17435 (N_17435,N_14802,N_14877);
and U17436 (N_17436,N_14390,N_15775);
nand U17437 (N_17437,N_15511,N_15516);
nand U17438 (N_17438,N_14832,N_14752);
xor U17439 (N_17439,N_15272,N_15132);
xor U17440 (N_17440,N_15614,N_15804);
or U17441 (N_17441,N_15704,N_14839);
or U17442 (N_17442,N_15863,N_14383);
and U17443 (N_17443,N_15663,N_14062);
xnor U17444 (N_17444,N_14220,N_15757);
nor U17445 (N_17445,N_14792,N_15468);
and U17446 (N_17446,N_15273,N_14030);
or U17447 (N_17447,N_14713,N_14851);
xor U17448 (N_17448,N_14705,N_15107);
nor U17449 (N_17449,N_15022,N_15363);
or U17450 (N_17450,N_15845,N_15651);
and U17451 (N_17451,N_15003,N_15712);
xnor U17452 (N_17452,N_15078,N_15125);
nor U17453 (N_17453,N_15946,N_15228);
nor U17454 (N_17454,N_14709,N_14099);
nand U17455 (N_17455,N_14287,N_15862);
nand U17456 (N_17456,N_14781,N_15321);
nand U17457 (N_17457,N_14276,N_14424);
or U17458 (N_17458,N_15203,N_14704);
nor U17459 (N_17459,N_15514,N_14730);
nor U17460 (N_17460,N_14663,N_14221);
or U17461 (N_17461,N_14196,N_15703);
nand U17462 (N_17462,N_14586,N_15187);
xor U17463 (N_17463,N_15121,N_15035);
nor U17464 (N_17464,N_14879,N_14562);
xnor U17465 (N_17465,N_14482,N_15435);
and U17466 (N_17466,N_15062,N_15105);
nor U17467 (N_17467,N_14823,N_14827);
xnor U17468 (N_17468,N_14476,N_14394);
nor U17469 (N_17469,N_14349,N_15130);
xnor U17470 (N_17470,N_15488,N_14717);
and U17471 (N_17471,N_15549,N_15801);
or U17472 (N_17472,N_15926,N_15308);
or U17473 (N_17473,N_15636,N_15129);
or U17474 (N_17474,N_14008,N_14274);
nor U17475 (N_17475,N_14715,N_14717);
and U17476 (N_17476,N_15173,N_15022);
and U17477 (N_17477,N_15762,N_15391);
and U17478 (N_17478,N_15572,N_15880);
and U17479 (N_17479,N_15612,N_15446);
and U17480 (N_17480,N_14995,N_14268);
or U17481 (N_17481,N_14599,N_14888);
and U17482 (N_17482,N_14873,N_15629);
nand U17483 (N_17483,N_14425,N_14048);
and U17484 (N_17484,N_14340,N_15885);
or U17485 (N_17485,N_15654,N_15633);
and U17486 (N_17486,N_14645,N_14316);
xor U17487 (N_17487,N_14059,N_15571);
nor U17488 (N_17488,N_14788,N_14810);
or U17489 (N_17489,N_14743,N_14095);
nor U17490 (N_17490,N_14199,N_14811);
nor U17491 (N_17491,N_15409,N_14056);
nor U17492 (N_17492,N_15362,N_14269);
and U17493 (N_17493,N_15339,N_14753);
or U17494 (N_17494,N_14879,N_15163);
or U17495 (N_17495,N_15915,N_15254);
or U17496 (N_17496,N_15284,N_15024);
and U17497 (N_17497,N_15531,N_15805);
xnor U17498 (N_17498,N_15857,N_14619);
and U17499 (N_17499,N_15174,N_14605);
xnor U17500 (N_17500,N_15434,N_14051);
nor U17501 (N_17501,N_14386,N_15632);
xor U17502 (N_17502,N_14014,N_15449);
and U17503 (N_17503,N_15879,N_14309);
nand U17504 (N_17504,N_15775,N_15570);
nand U17505 (N_17505,N_14321,N_14192);
and U17506 (N_17506,N_14318,N_15801);
or U17507 (N_17507,N_15011,N_14861);
nor U17508 (N_17508,N_15748,N_15668);
xnor U17509 (N_17509,N_14511,N_15425);
nor U17510 (N_17510,N_15603,N_15445);
and U17511 (N_17511,N_14829,N_15429);
nand U17512 (N_17512,N_14642,N_15363);
or U17513 (N_17513,N_14707,N_15100);
nand U17514 (N_17514,N_15457,N_15715);
and U17515 (N_17515,N_15796,N_15398);
nand U17516 (N_17516,N_14831,N_15302);
nand U17517 (N_17517,N_14591,N_15032);
nor U17518 (N_17518,N_14342,N_15759);
and U17519 (N_17519,N_15480,N_15695);
and U17520 (N_17520,N_15074,N_15634);
nor U17521 (N_17521,N_14946,N_15800);
and U17522 (N_17522,N_15756,N_15791);
and U17523 (N_17523,N_15375,N_15925);
and U17524 (N_17524,N_15251,N_15429);
nand U17525 (N_17525,N_14687,N_15099);
nand U17526 (N_17526,N_14182,N_14710);
and U17527 (N_17527,N_14234,N_15423);
or U17528 (N_17528,N_15785,N_15269);
nor U17529 (N_17529,N_14238,N_15468);
nand U17530 (N_17530,N_14880,N_14896);
nand U17531 (N_17531,N_15096,N_15562);
or U17532 (N_17532,N_14783,N_15466);
or U17533 (N_17533,N_15903,N_15643);
nor U17534 (N_17534,N_15702,N_14592);
nand U17535 (N_17535,N_15031,N_15364);
nand U17536 (N_17536,N_15010,N_15586);
and U17537 (N_17537,N_15111,N_15683);
nand U17538 (N_17538,N_15135,N_15379);
xnor U17539 (N_17539,N_15886,N_15545);
nor U17540 (N_17540,N_14874,N_14590);
xnor U17541 (N_17541,N_14785,N_15596);
xnor U17542 (N_17542,N_14366,N_14520);
and U17543 (N_17543,N_14507,N_14544);
nor U17544 (N_17544,N_14595,N_14961);
or U17545 (N_17545,N_15346,N_14906);
and U17546 (N_17546,N_14628,N_14428);
nor U17547 (N_17547,N_14963,N_15855);
nand U17548 (N_17548,N_14995,N_14844);
nand U17549 (N_17549,N_14484,N_15467);
nor U17550 (N_17550,N_14067,N_14782);
nor U17551 (N_17551,N_14737,N_15085);
nand U17552 (N_17552,N_14138,N_15814);
or U17553 (N_17553,N_14843,N_15332);
and U17554 (N_17554,N_14183,N_15176);
nor U17555 (N_17555,N_15644,N_14794);
xor U17556 (N_17556,N_14497,N_14275);
nand U17557 (N_17557,N_14063,N_15523);
nand U17558 (N_17558,N_14485,N_15503);
nor U17559 (N_17559,N_14909,N_15628);
xnor U17560 (N_17560,N_14426,N_14215);
nor U17561 (N_17561,N_15203,N_14834);
nor U17562 (N_17562,N_14250,N_14350);
nor U17563 (N_17563,N_14450,N_14777);
xor U17564 (N_17564,N_15672,N_14787);
and U17565 (N_17565,N_14596,N_15741);
nand U17566 (N_17566,N_14453,N_15685);
nor U17567 (N_17567,N_15371,N_15599);
nor U17568 (N_17568,N_15093,N_15987);
nor U17569 (N_17569,N_14939,N_14382);
xor U17570 (N_17570,N_14986,N_15197);
and U17571 (N_17571,N_15353,N_15543);
and U17572 (N_17572,N_14991,N_15623);
and U17573 (N_17573,N_15307,N_14149);
nand U17574 (N_17574,N_14021,N_15206);
and U17575 (N_17575,N_15803,N_15708);
or U17576 (N_17576,N_14194,N_15688);
xor U17577 (N_17577,N_14149,N_15958);
and U17578 (N_17578,N_15676,N_15344);
nor U17579 (N_17579,N_14614,N_15734);
xor U17580 (N_17580,N_15488,N_14722);
or U17581 (N_17581,N_14100,N_15569);
nand U17582 (N_17582,N_15233,N_15341);
xnor U17583 (N_17583,N_15324,N_15921);
and U17584 (N_17584,N_15228,N_15029);
nand U17585 (N_17585,N_15963,N_14703);
and U17586 (N_17586,N_14624,N_15900);
nand U17587 (N_17587,N_14607,N_15160);
nand U17588 (N_17588,N_14807,N_15763);
and U17589 (N_17589,N_15250,N_14133);
nand U17590 (N_17590,N_14287,N_15690);
nand U17591 (N_17591,N_15675,N_14093);
and U17592 (N_17592,N_14829,N_14935);
nor U17593 (N_17593,N_14094,N_15364);
xor U17594 (N_17594,N_15916,N_15207);
nor U17595 (N_17595,N_15518,N_14055);
nor U17596 (N_17596,N_14311,N_14576);
nand U17597 (N_17597,N_14927,N_15895);
xor U17598 (N_17598,N_14789,N_15564);
nand U17599 (N_17599,N_14814,N_14177);
nand U17600 (N_17600,N_15685,N_15326);
xnor U17601 (N_17601,N_15053,N_14628);
and U17602 (N_17602,N_14377,N_14311);
xnor U17603 (N_17603,N_14614,N_14541);
xnor U17604 (N_17604,N_14009,N_14204);
xor U17605 (N_17605,N_14851,N_15259);
xor U17606 (N_17606,N_15033,N_15333);
xor U17607 (N_17607,N_14704,N_14453);
and U17608 (N_17608,N_15014,N_14211);
nor U17609 (N_17609,N_14904,N_14460);
xor U17610 (N_17610,N_15374,N_15418);
and U17611 (N_17611,N_14184,N_15548);
or U17612 (N_17612,N_15132,N_14386);
or U17613 (N_17613,N_14842,N_15864);
xor U17614 (N_17614,N_14991,N_15866);
xor U17615 (N_17615,N_15717,N_14213);
and U17616 (N_17616,N_15838,N_14336);
nor U17617 (N_17617,N_14720,N_14293);
nor U17618 (N_17618,N_14543,N_14720);
or U17619 (N_17619,N_15862,N_15978);
and U17620 (N_17620,N_15892,N_14223);
or U17621 (N_17621,N_14051,N_15945);
and U17622 (N_17622,N_14834,N_15530);
or U17623 (N_17623,N_14188,N_14533);
and U17624 (N_17624,N_15797,N_15653);
or U17625 (N_17625,N_15081,N_14485);
and U17626 (N_17626,N_15308,N_15619);
xnor U17627 (N_17627,N_14353,N_14811);
nor U17628 (N_17628,N_15295,N_15602);
or U17629 (N_17629,N_14108,N_15533);
or U17630 (N_17630,N_15076,N_15548);
xor U17631 (N_17631,N_15375,N_15951);
xor U17632 (N_17632,N_15798,N_15589);
xnor U17633 (N_17633,N_15071,N_14673);
or U17634 (N_17634,N_14523,N_14955);
nand U17635 (N_17635,N_15557,N_14414);
xor U17636 (N_17636,N_14184,N_15516);
nand U17637 (N_17637,N_14606,N_15671);
xnor U17638 (N_17638,N_14555,N_15172);
or U17639 (N_17639,N_15249,N_14837);
and U17640 (N_17640,N_15699,N_14019);
or U17641 (N_17641,N_15382,N_15307);
xor U17642 (N_17642,N_15017,N_15492);
nand U17643 (N_17643,N_15167,N_15925);
xnor U17644 (N_17644,N_14438,N_15920);
xnor U17645 (N_17645,N_15312,N_14645);
and U17646 (N_17646,N_14886,N_14077);
xor U17647 (N_17647,N_14942,N_14763);
nor U17648 (N_17648,N_15393,N_14462);
xnor U17649 (N_17649,N_15551,N_15090);
and U17650 (N_17650,N_14011,N_14272);
nand U17651 (N_17651,N_15274,N_15376);
xnor U17652 (N_17652,N_14748,N_15385);
or U17653 (N_17653,N_14451,N_14011);
and U17654 (N_17654,N_15105,N_15581);
or U17655 (N_17655,N_15444,N_14274);
and U17656 (N_17656,N_15994,N_15456);
xor U17657 (N_17657,N_15573,N_14849);
nand U17658 (N_17658,N_14538,N_15861);
nand U17659 (N_17659,N_15021,N_15624);
or U17660 (N_17660,N_15870,N_15355);
xor U17661 (N_17661,N_15780,N_15292);
or U17662 (N_17662,N_15847,N_14204);
and U17663 (N_17663,N_15997,N_15403);
xnor U17664 (N_17664,N_15821,N_15631);
or U17665 (N_17665,N_15868,N_15736);
or U17666 (N_17666,N_15530,N_15206);
nor U17667 (N_17667,N_15743,N_15860);
nand U17668 (N_17668,N_15658,N_15690);
nand U17669 (N_17669,N_14415,N_14584);
nand U17670 (N_17670,N_14433,N_15395);
nand U17671 (N_17671,N_15700,N_14776);
or U17672 (N_17672,N_15704,N_15749);
nand U17673 (N_17673,N_14232,N_15164);
nand U17674 (N_17674,N_14903,N_14610);
and U17675 (N_17675,N_14950,N_14454);
nor U17676 (N_17676,N_14915,N_15687);
nor U17677 (N_17677,N_14855,N_15720);
nor U17678 (N_17678,N_15317,N_14875);
nand U17679 (N_17679,N_15422,N_14338);
nand U17680 (N_17680,N_14443,N_14257);
and U17681 (N_17681,N_14204,N_15112);
or U17682 (N_17682,N_14253,N_15752);
nor U17683 (N_17683,N_15763,N_15738);
or U17684 (N_17684,N_15126,N_14321);
xor U17685 (N_17685,N_15398,N_14048);
nor U17686 (N_17686,N_15657,N_15701);
nor U17687 (N_17687,N_14182,N_15812);
xor U17688 (N_17688,N_15535,N_15039);
and U17689 (N_17689,N_15920,N_14210);
xnor U17690 (N_17690,N_14667,N_14760);
nor U17691 (N_17691,N_15590,N_15471);
xnor U17692 (N_17692,N_15174,N_15715);
xor U17693 (N_17693,N_15781,N_14993);
nor U17694 (N_17694,N_15447,N_14484);
or U17695 (N_17695,N_15021,N_15449);
xnor U17696 (N_17696,N_15103,N_15000);
or U17697 (N_17697,N_15084,N_15558);
and U17698 (N_17698,N_15319,N_15508);
nor U17699 (N_17699,N_14187,N_15891);
xor U17700 (N_17700,N_14468,N_15014);
xnor U17701 (N_17701,N_15195,N_14658);
nand U17702 (N_17702,N_14737,N_14222);
xor U17703 (N_17703,N_15077,N_14190);
nor U17704 (N_17704,N_15851,N_15527);
and U17705 (N_17705,N_14804,N_15949);
and U17706 (N_17706,N_14211,N_14094);
nor U17707 (N_17707,N_14466,N_14928);
xnor U17708 (N_17708,N_15127,N_14878);
nor U17709 (N_17709,N_14612,N_15381);
and U17710 (N_17710,N_14972,N_14262);
nand U17711 (N_17711,N_15359,N_14595);
nor U17712 (N_17712,N_15140,N_15115);
and U17713 (N_17713,N_14830,N_15621);
nor U17714 (N_17714,N_15128,N_14556);
or U17715 (N_17715,N_14133,N_14833);
or U17716 (N_17716,N_14169,N_15514);
and U17717 (N_17717,N_15869,N_14034);
nor U17718 (N_17718,N_14637,N_15709);
xnor U17719 (N_17719,N_14048,N_15418);
nor U17720 (N_17720,N_15458,N_15787);
and U17721 (N_17721,N_14990,N_15576);
nand U17722 (N_17722,N_15111,N_14157);
and U17723 (N_17723,N_15001,N_15349);
and U17724 (N_17724,N_14977,N_15042);
and U17725 (N_17725,N_15127,N_14767);
or U17726 (N_17726,N_15384,N_14924);
xnor U17727 (N_17727,N_14965,N_14301);
nand U17728 (N_17728,N_15361,N_15011);
nand U17729 (N_17729,N_15058,N_15494);
or U17730 (N_17730,N_15092,N_15912);
or U17731 (N_17731,N_14437,N_15189);
xnor U17732 (N_17732,N_14819,N_15183);
xnor U17733 (N_17733,N_15594,N_15251);
or U17734 (N_17734,N_15281,N_14475);
and U17735 (N_17735,N_14946,N_15243);
xnor U17736 (N_17736,N_14463,N_15025);
nor U17737 (N_17737,N_14159,N_14087);
nor U17738 (N_17738,N_15038,N_15256);
nor U17739 (N_17739,N_14693,N_15655);
nand U17740 (N_17740,N_15762,N_15100);
or U17741 (N_17741,N_15640,N_15092);
nor U17742 (N_17742,N_15769,N_14653);
xnor U17743 (N_17743,N_15533,N_14059);
nor U17744 (N_17744,N_14541,N_15464);
nor U17745 (N_17745,N_14318,N_15040);
nor U17746 (N_17746,N_15953,N_14892);
and U17747 (N_17747,N_15075,N_14268);
and U17748 (N_17748,N_14889,N_14953);
and U17749 (N_17749,N_14422,N_14126);
and U17750 (N_17750,N_15759,N_14104);
and U17751 (N_17751,N_14335,N_15714);
xor U17752 (N_17752,N_14947,N_15708);
nor U17753 (N_17753,N_15340,N_15805);
and U17754 (N_17754,N_14015,N_14628);
or U17755 (N_17755,N_14980,N_15696);
nor U17756 (N_17756,N_14712,N_15304);
or U17757 (N_17757,N_14528,N_14028);
nor U17758 (N_17758,N_14198,N_14180);
and U17759 (N_17759,N_14180,N_15693);
and U17760 (N_17760,N_15471,N_14176);
nor U17761 (N_17761,N_15198,N_15107);
and U17762 (N_17762,N_15398,N_15905);
nor U17763 (N_17763,N_14771,N_14544);
nand U17764 (N_17764,N_14182,N_14823);
xor U17765 (N_17765,N_15621,N_14709);
and U17766 (N_17766,N_14970,N_15247);
xnor U17767 (N_17767,N_15563,N_14430);
or U17768 (N_17768,N_15677,N_15943);
xor U17769 (N_17769,N_14860,N_15230);
nand U17770 (N_17770,N_15943,N_14928);
nor U17771 (N_17771,N_14177,N_14497);
nand U17772 (N_17772,N_14303,N_14131);
nor U17773 (N_17773,N_14454,N_15757);
xor U17774 (N_17774,N_14337,N_15979);
xnor U17775 (N_17775,N_15170,N_14595);
and U17776 (N_17776,N_15934,N_15520);
nand U17777 (N_17777,N_14472,N_15556);
and U17778 (N_17778,N_15072,N_15195);
xor U17779 (N_17779,N_14683,N_15793);
nand U17780 (N_17780,N_15612,N_15723);
nand U17781 (N_17781,N_14677,N_15112);
nor U17782 (N_17782,N_14690,N_14893);
nand U17783 (N_17783,N_15843,N_15793);
xor U17784 (N_17784,N_14821,N_15807);
nand U17785 (N_17785,N_15469,N_15893);
nand U17786 (N_17786,N_15319,N_15315);
and U17787 (N_17787,N_15114,N_14214);
xnor U17788 (N_17788,N_14732,N_14794);
nand U17789 (N_17789,N_15333,N_14540);
or U17790 (N_17790,N_14753,N_14869);
nor U17791 (N_17791,N_14117,N_15948);
nand U17792 (N_17792,N_14044,N_14923);
nand U17793 (N_17793,N_15180,N_14971);
nand U17794 (N_17794,N_15839,N_14084);
or U17795 (N_17795,N_14432,N_14291);
or U17796 (N_17796,N_14501,N_15835);
xor U17797 (N_17797,N_14481,N_15426);
nor U17798 (N_17798,N_14228,N_14457);
or U17799 (N_17799,N_15601,N_15244);
and U17800 (N_17800,N_14772,N_14730);
or U17801 (N_17801,N_14247,N_15946);
nor U17802 (N_17802,N_14698,N_14264);
and U17803 (N_17803,N_15186,N_15837);
or U17804 (N_17804,N_15006,N_14915);
nor U17805 (N_17805,N_14253,N_15750);
and U17806 (N_17806,N_14542,N_14691);
xor U17807 (N_17807,N_14143,N_15377);
and U17808 (N_17808,N_15299,N_15291);
and U17809 (N_17809,N_15912,N_14029);
or U17810 (N_17810,N_15674,N_15396);
nand U17811 (N_17811,N_14784,N_15377);
nor U17812 (N_17812,N_15837,N_15869);
nand U17813 (N_17813,N_15949,N_14319);
or U17814 (N_17814,N_15991,N_15295);
xor U17815 (N_17815,N_15056,N_14806);
nor U17816 (N_17816,N_14489,N_14901);
or U17817 (N_17817,N_14536,N_15106);
and U17818 (N_17818,N_15102,N_14172);
xor U17819 (N_17819,N_15591,N_15597);
nor U17820 (N_17820,N_14466,N_14164);
nand U17821 (N_17821,N_14591,N_14434);
nor U17822 (N_17822,N_14659,N_14893);
and U17823 (N_17823,N_14317,N_15346);
nor U17824 (N_17824,N_15038,N_15273);
or U17825 (N_17825,N_14152,N_15374);
nor U17826 (N_17826,N_15561,N_15175);
or U17827 (N_17827,N_15497,N_14481);
xnor U17828 (N_17828,N_14332,N_15721);
or U17829 (N_17829,N_14623,N_14513);
or U17830 (N_17830,N_15824,N_14871);
xor U17831 (N_17831,N_15401,N_15840);
or U17832 (N_17832,N_14799,N_14629);
xnor U17833 (N_17833,N_14676,N_14516);
or U17834 (N_17834,N_14415,N_14661);
nand U17835 (N_17835,N_14182,N_14591);
and U17836 (N_17836,N_15063,N_14332);
xor U17837 (N_17837,N_15737,N_15957);
and U17838 (N_17838,N_14131,N_15061);
xnor U17839 (N_17839,N_15295,N_15950);
and U17840 (N_17840,N_15784,N_14382);
or U17841 (N_17841,N_14084,N_14807);
nor U17842 (N_17842,N_15685,N_14600);
nand U17843 (N_17843,N_14770,N_15751);
xnor U17844 (N_17844,N_14808,N_15430);
xor U17845 (N_17845,N_14225,N_14508);
or U17846 (N_17846,N_14095,N_15694);
xor U17847 (N_17847,N_15873,N_15136);
nor U17848 (N_17848,N_14005,N_15249);
nor U17849 (N_17849,N_15469,N_14602);
and U17850 (N_17850,N_14446,N_15291);
and U17851 (N_17851,N_15796,N_14797);
xor U17852 (N_17852,N_14842,N_14604);
xor U17853 (N_17853,N_14088,N_15446);
nand U17854 (N_17854,N_15273,N_14781);
xor U17855 (N_17855,N_14857,N_14480);
nand U17856 (N_17856,N_15470,N_15098);
nand U17857 (N_17857,N_14881,N_14135);
xnor U17858 (N_17858,N_15829,N_15647);
nand U17859 (N_17859,N_15972,N_14051);
xor U17860 (N_17860,N_15119,N_14633);
and U17861 (N_17861,N_15231,N_14868);
nor U17862 (N_17862,N_15200,N_15726);
or U17863 (N_17863,N_14380,N_14351);
or U17864 (N_17864,N_15195,N_15642);
xnor U17865 (N_17865,N_15991,N_15731);
nand U17866 (N_17866,N_15167,N_14079);
and U17867 (N_17867,N_15046,N_14241);
nand U17868 (N_17868,N_15566,N_15388);
and U17869 (N_17869,N_15965,N_14043);
and U17870 (N_17870,N_15343,N_14884);
xnor U17871 (N_17871,N_14031,N_14124);
or U17872 (N_17872,N_15503,N_14650);
nand U17873 (N_17873,N_15668,N_15137);
or U17874 (N_17874,N_15485,N_15871);
or U17875 (N_17875,N_14937,N_15765);
nand U17876 (N_17876,N_15673,N_14530);
or U17877 (N_17877,N_15610,N_14719);
xnor U17878 (N_17878,N_15024,N_14700);
nand U17879 (N_17879,N_15340,N_14984);
nand U17880 (N_17880,N_15473,N_14046);
nor U17881 (N_17881,N_14995,N_15099);
nor U17882 (N_17882,N_14367,N_14058);
nand U17883 (N_17883,N_15411,N_15439);
nand U17884 (N_17884,N_15445,N_15046);
nor U17885 (N_17885,N_14863,N_15238);
or U17886 (N_17886,N_14747,N_14662);
and U17887 (N_17887,N_14968,N_14717);
and U17888 (N_17888,N_15271,N_15678);
and U17889 (N_17889,N_15610,N_15082);
or U17890 (N_17890,N_14533,N_14914);
and U17891 (N_17891,N_14401,N_15091);
or U17892 (N_17892,N_14764,N_14711);
or U17893 (N_17893,N_15717,N_15949);
nand U17894 (N_17894,N_15865,N_14494);
xor U17895 (N_17895,N_15569,N_14789);
and U17896 (N_17896,N_14312,N_15115);
nand U17897 (N_17897,N_15856,N_14839);
nor U17898 (N_17898,N_15756,N_14467);
xnor U17899 (N_17899,N_14264,N_15208);
xor U17900 (N_17900,N_14426,N_15556);
xnor U17901 (N_17901,N_14021,N_15844);
and U17902 (N_17902,N_14642,N_14509);
xor U17903 (N_17903,N_14994,N_15085);
and U17904 (N_17904,N_15249,N_14949);
or U17905 (N_17905,N_14389,N_14007);
nor U17906 (N_17906,N_14233,N_14295);
or U17907 (N_17907,N_15878,N_15594);
xnor U17908 (N_17908,N_14681,N_14378);
or U17909 (N_17909,N_14895,N_14811);
or U17910 (N_17910,N_15404,N_15784);
xor U17911 (N_17911,N_14826,N_14933);
or U17912 (N_17912,N_15867,N_15747);
nand U17913 (N_17913,N_15447,N_15405);
nand U17914 (N_17914,N_15552,N_14129);
and U17915 (N_17915,N_14249,N_15911);
or U17916 (N_17916,N_15602,N_15002);
nor U17917 (N_17917,N_15450,N_15344);
nand U17918 (N_17918,N_15821,N_14244);
and U17919 (N_17919,N_15877,N_14304);
and U17920 (N_17920,N_14950,N_15728);
nor U17921 (N_17921,N_15918,N_15056);
and U17922 (N_17922,N_14503,N_14983);
and U17923 (N_17923,N_14882,N_14645);
xnor U17924 (N_17924,N_14006,N_15839);
nand U17925 (N_17925,N_15802,N_15116);
xnor U17926 (N_17926,N_14727,N_14321);
nor U17927 (N_17927,N_14831,N_14283);
nand U17928 (N_17928,N_14472,N_14148);
nor U17929 (N_17929,N_14307,N_14840);
nand U17930 (N_17930,N_15853,N_14414);
nor U17931 (N_17931,N_14154,N_14720);
nand U17932 (N_17932,N_14096,N_15483);
or U17933 (N_17933,N_15947,N_15279);
or U17934 (N_17934,N_14124,N_15308);
nor U17935 (N_17935,N_15861,N_14640);
xnor U17936 (N_17936,N_14815,N_15511);
nor U17937 (N_17937,N_15664,N_14513);
nand U17938 (N_17938,N_14116,N_14602);
nand U17939 (N_17939,N_15995,N_15408);
xnor U17940 (N_17940,N_14489,N_14960);
nand U17941 (N_17941,N_14163,N_15641);
nor U17942 (N_17942,N_15540,N_15038);
nor U17943 (N_17943,N_15050,N_14066);
nor U17944 (N_17944,N_15099,N_15890);
and U17945 (N_17945,N_14534,N_15380);
and U17946 (N_17946,N_14982,N_15500);
nand U17947 (N_17947,N_15676,N_15158);
xnor U17948 (N_17948,N_14457,N_15626);
or U17949 (N_17949,N_15600,N_14290);
or U17950 (N_17950,N_14550,N_14577);
nand U17951 (N_17951,N_15806,N_14035);
xnor U17952 (N_17952,N_15699,N_14886);
nor U17953 (N_17953,N_14734,N_14102);
xnor U17954 (N_17954,N_14023,N_15084);
nand U17955 (N_17955,N_14991,N_15021);
and U17956 (N_17956,N_15959,N_15736);
xor U17957 (N_17957,N_15850,N_14125);
and U17958 (N_17958,N_14781,N_14662);
and U17959 (N_17959,N_15089,N_15699);
xor U17960 (N_17960,N_15449,N_15892);
and U17961 (N_17961,N_14659,N_15372);
xnor U17962 (N_17962,N_15881,N_15876);
xnor U17963 (N_17963,N_14403,N_14939);
xnor U17964 (N_17964,N_14139,N_14494);
nand U17965 (N_17965,N_15906,N_14857);
or U17966 (N_17966,N_14474,N_14835);
xnor U17967 (N_17967,N_15201,N_14414);
nand U17968 (N_17968,N_14176,N_14674);
nor U17969 (N_17969,N_15464,N_15283);
xnor U17970 (N_17970,N_14541,N_15907);
nand U17971 (N_17971,N_15929,N_15352);
xnor U17972 (N_17972,N_15764,N_15765);
or U17973 (N_17973,N_15678,N_15926);
or U17974 (N_17974,N_14776,N_15624);
and U17975 (N_17975,N_15231,N_15088);
and U17976 (N_17976,N_15753,N_14492);
and U17977 (N_17977,N_15745,N_15630);
nor U17978 (N_17978,N_15063,N_15331);
nand U17979 (N_17979,N_14231,N_14199);
nor U17980 (N_17980,N_14693,N_15327);
nand U17981 (N_17981,N_14394,N_15723);
xnor U17982 (N_17982,N_15739,N_14166);
or U17983 (N_17983,N_15523,N_14073);
or U17984 (N_17984,N_14487,N_14479);
and U17985 (N_17985,N_14415,N_14195);
xor U17986 (N_17986,N_14376,N_15740);
xnor U17987 (N_17987,N_15152,N_15424);
nand U17988 (N_17988,N_14534,N_14763);
or U17989 (N_17989,N_15235,N_14842);
nor U17990 (N_17990,N_14731,N_14078);
nand U17991 (N_17991,N_15785,N_15263);
and U17992 (N_17992,N_14798,N_15843);
and U17993 (N_17993,N_14441,N_15643);
and U17994 (N_17994,N_15300,N_15698);
and U17995 (N_17995,N_14031,N_14397);
nor U17996 (N_17996,N_15679,N_14910);
and U17997 (N_17997,N_15583,N_14908);
or U17998 (N_17998,N_14217,N_15000);
xor U17999 (N_17999,N_14129,N_15259);
nand U18000 (N_18000,N_17002,N_16443);
and U18001 (N_18001,N_16357,N_16985);
or U18002 (N_18002,N_17775,N_16156);
or U18003 (N_18003,N_17708,N_16368);
nand U18004 (N_18004,N_17857,N_17163);
nand U18005 (N_18005,N_16235,N_17950);
nand U18006 (N_18006,N_17821,N_17494);
and U18007 (N_18007,N_16223,N_17661);
nor U18008 (N_18008,N_16463,N_17651);
nor U18009 (N_18009,N_16339,N_17370);
or U18010 (N_18010,N_16602,N_16640);
nor U18011 (N_18011,N_16575,N_17735);
nor U18012 (N_18012,N_17138,N_17445);
nor U18013 (N_18013,N_17953,N_17529);
and U18014 (N_18014,N_16597,N_17783);
or U18015 (N_18015,N_17923,N_16404);
and U18016 (N_18016,N_17510,N_17200);
and U18017 (N_18017,N_16120,N_16215);
and U18018 (N_18018,N_16583,N_16727);
and U18019 (N_18019,N_17516,N_17013);
and U18020 (N_18020,N_17337,N_17047);
xnor U18021 (N_18021,N_17052,N_17738);
nor U18022 (N_18022,N_16899,N_16166);
xnor U18023 (N_18023,N_16058,N_16721);
nor U18024 (N_18024,N_17543,N_17723);
or U18025 (N_18025,N_16196,N_16941);
and U18026 (N_18026,N_17157,N_17976);
xor U18027 (N_18027,N_17416,N_17823);
nor U18028 (N_18028,N_16651,N_17176);
nor U18029 (N_18029,N_17064,N_17961);
or U18030 (N_18030,N_16806,N_17643);
and U18031 (N_18031,N_17024,N_17262);
nand U18032 (N_18032,N_16359,N_16658);
nand U18033 (N_18033,N_17095,N_17122);
or U18034 (N_18034,N_17703,N_17790);
and U18035 (N_18035,N_17376,N_16674);
and U18036 (N_18036,N_17264,N_16712);
or U18037 (N_18037,N_17880,N_16242);
or U18038 (N_18038,N_16672,N_16479);
nor U18039 (N_18039,N_17518,N_16654);
or U18040 (N_18040,N_16416,N_16092);
or U18041 (N_18041,N_16016,N_17142);
nand U18042 (N_18042,N_16229,N_16613);
and U18043 (N_18043,N_16686,N_16197);
xor U18044 (N_18044,N_17909,N_17758);
nand U18045 (N_18045,N_17873,N_17183);
and U18046 (N_18046,N_16446,N_17637);
nor U18047 (N_18047,N_17087,N_16764);
and U18048 (N_18048,N_16255,N_16670);
or U18049 (N_18049,N_17288,N_16722);
nand U18050 (N_18050,N_17436,N_17496);
or U18051 (N_18051,N_17926,N_16961);
or U18052 (N_18052,N_16834,N_16490);
and U18053 (N_18053,N_17074,N_16250);
or U18054 (N_18054,N_17110,N_17018);
and U18055 (N_18055,N_17294,N_16375);
nor U18056 (N_18056,N_17185,N_16118);
or U18057 (N_18057,N_16800,N_16152);
nand U18058 (N_18058,N_17143,N_17053);
nand U18059 (N_18059,N_17509,N_16681);
or U18060 (N_18060,N_16205,N_17784);
nand U18061 (N_18061,N_17573,N_17903);
xor U18062 (N_18062,N_17302,N_16224);
nor U18063 (N_18063,N_17860,N_16559);
nor U18064 (N_18064,N_16260,N_17048);
or U18065 (N_18065,N_16638,N_17270);
nor U18066 (N_18066,N_16932,N_17676);
nor U18067 (N_18067,N_16923,N_16586);
xnor U18068 (N_18068,N_17710,N_16207);
and U18069 (N_18069,N_17041,N_17554);
xor U18070 (N_18070,N_17888,N_16587);
and U18071 (N_18071,N_16744,N_16927);
nor U18072 (N_18072,N_17447,N_16705);
and U18073 (N_18073,N_16264,N_17653);
nor U18074 (N_18074,N_17442,N_17464);
nand U18075 (N_18075,N_16763,N_16171);
nor U18076 (N_18076,N_16488,N_16667);
and U18077 (N_18077,N_16856,N_16096);
xnor U18078 (N_18078,N_17113,N_16618);
or U18079 (N_18079,N_17646,N_16371);
xnor U18080 (N_18080,N_17353,N_16859);
nand U18081 (N_18081,N_17021,N_17117);
nand U18082 (N_18082,N_17306,N_17852);
xnor U18083 (N_18083,N_16256,N_16194);
and U18084 (N_18084,N_17596,N_17722);
or U18085 (N_18085,N_16087,N_16019);
xnor U18086 (N_18086,N_16792,N_17339);
nand U18087 (N_18087,N_16656,N_16566);
xor U18088 (N_18088,N_16478,N_16348);
or U18089 (N_18089,N_17345,N_16794);
and U18090 (N_18090,N_16939,N_16698);
nand U18091 (N_18091,N_17740,N_17235);
or U18092 (N_18092,N_16541,N_16607);
and U18093 (N_18093,N_16228,N_17806);
or U18094 (N_18094,N_17569,N_16452);
and U18095 (N_18095,N_16950,N_17299);
nor U18096 (N_18096,N_17937,N_16826);
and U18097 (N_18097,N_16955,N_16252);
nand U18098 (N_18098,N_16690,N_17607);
nor U18099 (N_18099,N_17839,N_16027);
and U18100 (N_18100,N_17473,N_17606);
and U18101 (N_18101,N_17290,N_16975);
and U18102 (N_18102,N_17215,N_16270);
nand U18103 (N_18103,N_17156,N_16468);
or U18104 (N_18104,N_17212,N_17896);
xnor U18105 (N_18105,N_17136,N_16759);
xnor U18106 (N_18106,N_17469,N_17556);
and U18107 (N_18107,N_17182,N_17150);
and U18108 (N_18108,N_16983,N_16288);
and U18109 (N_18109,N_17441,N_16878);
nor U18110 (N_18110,N_16053,N_16879);
or U18111 (N_18111,N_17450,N_16007);
nor U18112 (N_18112,N_16810,N_16400);
nand U18113 (N_18113,N_16377,N_16106);
nand U18114 (N_18114,N_17311,N_16465);
nor U18115 (N_18115,N_17466,N_16818);
and U18116 (N_18116,N_17550,N_17906);
nor U18117 (N_18117,N_17387,N_16100);
or U18118 (N_18118,N_16994,N_17181);
and U18119 (N_18119,N_17360,N_17797);
xor U18120 (N_18120,N_16929,N_16451);
nor U18121 (N_18121,N_16259,N_16432);
nand U18122 (N_18122,N_17962,N_16620);
nand U18123 (N_18123,N_17045,N_17497);
and U18124 (N_18124,N_16382,N_16904);
or U18125 (N_18125,N_17378,N_17816);
or U18126 (N_18126,N_16139,N_17978);
nand U18127 (N_18127,N_16931,N_16440);
nand U18128 (N_18128,N_16274,N_16769);
nor U18129 (N_18129,N_17046,N_17170);
and U18130 (N_18130,N_16454,N_17944);
or U18131 (N_18131,N_17366,N_16609);
or U18132 (N_18132,N_16525,N_16655);
nor U18133 (N_18133,N_16268,N_17227);
and U18134 (N_18134,N_16233,N_16206);
nand U18135 (N_18135,N_16009,N_17373);
and U18136 (N_18136,N_17265,N_17603);
xor U18137 (N_18137,N_17928,N_16311);
or U18138 (N_18138,N_17406,N_17620);
nor U18139 (N_18139,N_16063,N_16519);
nand U18140 (N_18140,N_16325,N_16456);
or U18141 (N_18141,N_17462,N_16112);
or U18142 (N_18142,N_17598,N_17491);
xnor U18143 (N_18143,N_16379,N_16304);
xnor U18144 (N_18144,N_16881,N_17774);
nor U18145 (N_18145,N_16491,N_17233);
and U18146 (N_18146,N_17546,N_17530);
and U18147 (N_18147,N_16815,N_16303);
and U18148 (N_18148,N_16489,N_16987);
and U18149 (N_18149,N_16369,N_17963);
xnor U18150 (N_18150,N_17936,N_16949);
xnor U18151 (N_18151,N_17901,N_17879);
xnor U18152 (N_18152,N_16807,N_17418);
and U18153 (N_18153,N_16439,N_17849);
nor U18154 (N_18154,N_16542,N_16854);
or U18155 (N_18155,N_17161,N_16165);
xor U18156 (N_18156,N_17955,N_16410);
or U18157 (N_18157,N_17040,N_17508);
nor U18158 (N_18158,N_16025,N_16663);
and U18159 (N_18159,N_16665,N_16277);
and U18160 (N_18160,N_16765,N_17599);
nand U18161 (N_18161,N_16631,N_16610);
xor U18162 (N_18162,N_17419,N_17446);
and U18163 (N_18163,N_17482,N_16403);
nand U18164 (N_18164,N_16459,N_17335);
nor U18165 (N_18165,N_16175,N_17089);
nor U18166 (N_18166,N_17433,N_16845);
or U18167 (N_18167,N_16911,N_17555);
nand U18168 (N_18168,N_16756,N_17384);
nor U18169 (N_18169,N_16883,N_17776);
nand U18170 (N_18170,N_16389,N_16653);
nand U18171 (N_18171,N_17644,N_16760);
nor U18172 (N_18172,N_17773,N_16540);
or U18173 (N_18173,N_17582,N_16601);
and U18174 (N_18174,N_17078,N_16438);
or U18175 (N_18175,N_17662,N_17241);
and U18176 (N_18176,N_16292,N_17875);
or U18177 (N_18177,N_17781,N_16280);
or U18178 (N_18178,N_16098,N_16392);
nor U18179 (N_18179,N_16507,N_16033);
and U18180 (N_18180,N_17884,N_17291);
nand U18181 (N_18181,N_17260,N_16900);
or U18182 (N_18182,N_17818,N_16317);
xor U18183 (N_18183,N_17871,N_16714);
nand U18184 (N_18184,N_16340,N_16921);
and U18185 (N_18185,N_16185,N_16145);
xor U18186 (N_18186,N_16622,N_17721);
xor U18187 (N_18187,N_16868,N_16189);
xnor U18188 (N_18188,N_16700,N_16436);
and U18189 (N_18189,N_17507,N_17540);
or U18190 (N_18190,N_16405,N_17756);
xnor U18191 (N_18191,N_17899,N_17847);
and U18192 (N_18192,N_16467,N_16547);
nor U18193 (N_18193,N_16528,N_16829);
and U18194 (N_18194,N_16821,N_16361);
or U18195 (N_18195,N_17855,N_16411);
xnor U18196 (N_18196,N_17224,N_16360);
and U18197 (N_18197,N_16257,N_17779);
xnor U18198 (N_18198,N_16676,N_16214);
or U18199 (N_18199,N_16462,N_16203);
xor U18200 (N_18200,N_16937,N_17650);
xor U18201 (N_18201,N_16153,N_17751);
and U18202 (N_18202,N_16430,N_17704);
nand U18203 (N_18203,N_17747,N_16871);
or U18204 (N_18204,N_17254,N_17539);
xor U18205 (N_18205,N_16297,N_16890);
and U18206 (N_18206,N_16835,N_16928);
or U18207 (N_18207,N_16989,N_17440);
and U18208 (N_18208,N_16933,N_17330);
nand U18209 (N_18209,N_17983,N_16604);
nand U18210 (N_18210,N_17697,N_16549);
nand U18211 (N_18211,N_16942,N_16254);
nor U18212 (N_18212,N_16673,N_16837);
nor U18213 (N_18213,N_16953,N_17403);
nand U18214 (N_18214,N_17296,N_17175);
or U18215 (N_18215,N_17870,N_17493);
and U18216 (N_18216,N_16273,N_17451);
or U18217 (N_18217,N_16367,N_17336);
nor U18218 (N_18218,N_17851,N_16159);
nand U18219 (N_18219,N_17481,N_17467);
xnor U18220 (N_18220,N_17794,N_16234);
and U18221 (N_18221,N_17557,N_17067);
xor U18222 (N_18222,N_17568,N_16148);
xor U18223 (N_18223,N_16683,N_17734);
nand U18224 (N_18224,N_16295,N_16778);
and U18225 (N_18225,N_16321,N_17898);
nand U18226 (N_18226,N_17334,N_16570);
or U18227 (N_18227,N_16925,N_17997);
xnor U18228 (N_18228,N_16788,N_17397);
nor U18229 (N_18229,N_17576,N_16567);
nor U18230 (N_18230,N_17027,N_16426);
nor U18231 (N_18231,N_17239,N_16814);
and U18232 (N_18232,N_17631,N_17717);
xnor U18233 (N_18233,N_16823,N_17358);
nand U18234 (N_18234,N_17101,N_17700);
nor U18235 (N_18235,N_17295,N_17489);
or U18236 (N_18236,N_17253,N_17686);
nor U18237 (N_18237,N_17885,N_16743);
xnor U18238 (N_18238,N_16450,N_16523);
nand U18239 (N_18239,N_16804,N_16381);
or U18240 (N_18240,N_17549,N_17275);
xnor U18241 (N_18241,N_17198,N_16038);
or U18242 (N_18242,N_16675,N_16047);
nor U18243 (N_18243,N_16888,N_16715);
xnor U18244 (N_18244,N_16353,N_17544);
xnor U18245 (N_18245,N_17413,N_17084);
xor U18246 (N_18246,N_16230,N_17541);
nand U18247 (N_18247,N_16493,N_16444);
nand U18248 (N_18248,N_17038,N_16569);
and U18249 (N_18249,N_16544,N_17992);
and U18250 (N_18250,N_17395,N_17191);
xor U18251 (N_18251,N_17782,N_17558);
nor U18252 (N_18252,N_17245,N_17553);
nand U18253 (N_18253,N_16202,N_16103);
nand U18254 (N_18254,N_17780,N_17483);
xor U18255 (N_18255,N_16819,N_16924);
or U18256 (N_18256,N_17471,N_17164);
nand U18257 (N_18257,N_17051,N_17169);
nor U18258 (N_18258,N_17513,N_16331);
or U18259 (N_18259,N_16135,N_16090);
xnor U18260 (N_18260,N_17465,N_17144);
and U18261 (N_18261,N_17984,N_17097);
or U18262 (N_18262,N_17055,N_17349);
and U18263 (N_18263,N_17590,N_17907);
and U18264 (N_18264,N_17987,N_17999);
nand U18265 (N_18265,N_16412,N_16515);
nand U18266 (N_18266,N_16825,N_17114);
and U18267 (N_18267,N_16934,N_16212);
nor U18268 (N_18268,N_16780,N_16336);
nand U18269 (N_18269,N_16809,N_17242);
or U18270 (N_18270,N_16969,N_16457);
nand U18271 (N_18271,N_16435,N_17035);
or U18272 (N_18272,N_16115,N_17934);
nand U18273 (N_18273,N_16157,N_17730);
xor U18274 (N_18274,N_16013,N_16434);
or U18275 (N_18275,N_17908,N_17656);
nand U18276 (N_18276,N_16930,N_16948);
nand U18277 (N_18277,N_16827,N_16945);
or U18278 (N_18278,N_17574,N_16739);
or U18279 (N_18279,N_17031,N_16729);
nand U18280 (N_18280,N_17537,N_16101);
or U18281 (N_18281,N_16086,N_16966);
and U18282 (N_18282,N_17970,N_17868);
nor U18283 (N_18283,N_16864,N_16067);
nor U18284 (N_18284,N_16015,N_17993);
or U18285 (N_18285,N_17189,N_17190);
and U18286 (N_18286,N_17272,N_16088);
and U18287 (N_18287,N_17259,N_16838);
nor U18288 (N_18288,N_17461,N_17742);
nor U18289 (N_18289,N_16299,N_17841);
or U18290 (N_18290,N_16487,N_17203);
nor U18291 (N_18291,N_17586,N_17792);
nand U18292 (N_18292,N_17332,N_16737);
xnor U18293 (N_18293,N_17329,N_17531);
or U18294 (N_18294,N_17500,N_17679);
xor U18295 (N_18295,N_17754,N_16483);
xor U18296 (N_18296,N_16352,N_17228);
nor U18297 (N_18297,N_17216,N_17989);
or U18298 (N_18298,N_16240,N_16146);
nor U18299 (N_18299,N_17659,N_16751);
nor U18300 (N_18300,N_16577,N_17398);
and U18301 (N_18301,N_17524,N_17155);
nand U18302 (N_18302,N_16977,N_17913);
nor U18303 (N_18303,N_17402,N_17960);
and U18304 (N_18304,N_17098,N_17042);
xor U18305 (N_18305,N_17344,N_17837);
and U18306 (N_18306,N_17956,N_16776);
nor U18307 (N_18307,N_16247,N_16946);
nand U18308 (N_18308,N_16637,N_17325);
or U18309 (N_18309,N_17567,N_17386);
nand U18310 (N_18310,N_17830,N_16351);
nand U18311 (N_18311,N_17522,N_17129);
nor U18312 (N_18312,N_17526,N_17608);
nor U18313 (N_18313,N_17577,N_17005);
or U18314 (N_18314,N_16574,N_16576);
nor U18315 (N_18315,N_16874,N_17995);
nand U18316 (N_18316,N_16006,N_16679);
nor U18317 (N_18317,N_17111,N_16972);
nor U18318 (N_18318,N_17785,N_16789);
xnor U18319 (N_18319,N_16364,N_16076);
xor U18320 (N_18320,N_16844,N_16530);
nand U18321 (N_18321,N_17059,N_17417);
and U18322 (N_18322,N_16248,N_17625);
nand U18323 (N_18323,N_16278,N_16272);
and U18324 (N_18324,N_16316,N_17848);
nand U18325 (N_18325,N_16652,N_16269);
xor U18326 (N_18326,N_17994,N_16726);
or U18327 (N_18327,N_16867,N_17057);
nor U18328 (N_18328,N_16306,N_16568);
nor U18329 (N_18329,N_17719,N_16554);
nand U18330 (N_18330,N_17204,N_17720);
nor U18331 (N_18331,N_16704,N_17286);
and U18332 (N_18332,N_16901,N_17008);
and U18333 (N_18333,N_16048,N_17752);
xnor U18334 (N_18334,N_16603,N_16908);
nor U18335 (N_18335,N_17617,N_17621);
nor U18336 (N_18336,N_16198,N_16070);
or U18337 (N_18337,N_17869,N_16345);
or U18338 (N_18338,N_17015,N_17105);
nand U18339 (N_18339,N_17083,N_16448);
or U18340 (N_18340,N_16464,N_16407);
and U18341 (N_18341,N_17388,N_17072);
or U18342 (N_18342,N_17864,N_17813);
and U18343 (N_18343,N_17162,N_17106);
and U18344 (N_18344,N_16266,N_17192);
xnor U18345 (N_18345,N_16029,N_17692);
and U18346 (N_18346,N_17385,N_16920);
nand U18347 (N_18347,N_17404,N_16265);
or U18348 (N_18348,N_17412,N_17743);
or U18349 (N_18349,N_17948,N_16851);
nor U18350 (N_18350,N_17560,N_17627);
nand U18351 (N_18351,N_16805,N_17633);
and U18352 (N_18352,N_17248,N_16388);
or U18353 (N_18353,N_17075,N_17043);
nor U18354 (N_18354,N_17152,N_17639);
and U18355 (N_18355,N_17109,N_16329);
and U18356 (N_18356,N_17941,N_17749);
nand U18357 (N_18357,N_17535,N_16719);
and U18358 (N_18358,N_16841,N_17528);
nand U18359 (N_18359,N_17796,N_17480);
or U18360 (N_18360,N_16561,N_17120);
and U18361 (N_18361,N_16619,N_17077);
and U18362 (N_18362,N_16896,N_16614);
or U18363 (N_18363,N_16012,N_17635);
nor U18364 (N_18364,N_16976,N_16645);
nand U18365 (N_18365,N_17564,N_16319);
xnor U18366 (N_18366,N_16536,N_16884);
or U18367 (N_18367,N_16232,N_16555);
or U18368 (N_18368,N_16124,N_16671);
nand U18369 (N_18369,N_16091,N_16177);
nand U18370 (N_18370,N_17660,N_17279);
nand U18371 (N_18371,N_16641,N_17118);
xnor U18372 (N_18372,N_16730,N_17802);
or U18373 (N_18373,N_16831,N_17044);
nor U18374 (N_18374,N_17092,N_16149);
and U18375 (N_18375,N_17019,N_16628);
or U18376 (N_18376,N_16696,N_17408);
or U18377 (N_18377,N_16738,N_16075);
nand U18378 (N_18378,N_17527,N_16307);
nand U18379 (N_18379,N_17793,N_16691);
or U18380 (N_18380,N_17915,N_17093);
or U18381 (N_18381,N_16011,N_16636);
nand U18382 (N_18382,N_16122,N_17640);
xnor U18383 (N_18383,N_17297,N_17060);
nor U18384 (N_18384,N_17929,N_17243);
or U18385 (N_18385,N_16190,N_17916);
nand U18386 (N_18386,N_17671,N_17410);
nor U18387 (N_18387,N_16216,N_17867);
and U18388 (N_18388,N_17379,N_17677);
and U18389 (N_18389,N_16161,N_16060);
or U18390 (N_18390,N_16590,N_16813);
nor U18391 (N_18391,N_16855,N_17593);
and U18392 (N_18392,N_17981,N_17917);
and U18393 (N_18393,N_16220,N_17218);
or U18394 (N_18394,N_17892,N_16922);
and U18395 (N_18395,N_17935,N_17623);
nor U18396 (N_18396,N_16745,N_17430);
xor U18397 (N_18397,N_17769,N_16421);
nand U18398 (N_18398,N_16347,N_16521);
or U18399 (N_18399,N_17277,N_16593);
and U18400 (N_18400,N_17246,N_17853);
nand U18401 (N_18401,N_17237,N_16134);
and U18402 (N_18402,N_16581,N_17112);
and U18403 (N_18403,N_16499,N_16055);
or U18404 (N_18404,N_17287,N_17595);
nand U18405 (N_18405,N_17977,N_17274);
and U18406 (N_18406,N_17392,N_16849);
and U18407 (N_18407,N_17826,N_16936);
xnor U18408 (N_18408,N_17707,N_17069);
nor U18409 (N_18409,N_17611,N_17149);
nand U18410 (N_18410,N_17602,N_16693);
and U18411 (N_18411,N_17820,N_16947);
or U18412 (N_18412,N_16167,N_16370);
or U18413 (N_18413,N_16057,N_17548);
nor U18414 (N_18414,N_17694,N_17396);
or U18415 (N_18415,N_16768,N_17912);
xnor U18416 (N_18416,N_16023,N_16179);
xor U18417 (N_18417,N_17894,N_16282);
and U18418 (N_18418,N_17389,N_17804);
and U18419 (N_18419,N_16423,N_17423);
or U18420 (N_18420,N_17727,N_16591);
nor U18421 (N_18421,N_17099,N_16072);
and U18422 (N_18422,N_16752,N_16938);
or U18423 (N_18423,N_17029,N_16736);
nor U18424 (N_18424,N_16066,N_16384);
xnor U18425 (N_18425,N_17145,N_16850);
or U18426 (N_18426,N_16799,N_17943);
nand U18427 (N_18427,N_16533,N_16968);
nor U18428 (N_18428,N_16287,N_16535);
nor U18429 (N_18429,N_16828,N_17405);
xor U18430 (N_18430,N_17887,N_16082);
and U18431 (N_18431,N_16173,N_17391);
and U18432 (N_18432,N_17657,N_17054);
or U18433 (N_18433,N_16720,N_17897);
xor U18434 (N_18434,N_17814,N_17940);
or U18435 (N_18435,N_17791,N_16741);
nor U18436 (N_18436,N_16915,N_16445);
or U18437 (N_18437,N_16372,N_17835);
xnor U18438 (N_18438,N_17230,N_16300);
xnor U18439 (N_18439,N_17188,N_17016);
or U18440 (N_18440,N_17448,N_16777);
or U18441 (N_18441,N_16427,N_17681);
nor U18442 (N_18442,N_17363,N_16119);
xnor U18443 (N_18443,N_17589,N_16695);
and U18444 (N_18444,N_16046,N_17572);
xor U18445 (N_18445,N_16095,N_16740);
nor U18446 (N_18446,N_16358,N_16885);
nor U18447 (N_18447,N_16332,N_17647);
nor U18448 (N_18448,N_16643,N_16863);
nor U18449 (N_18449,N_16470,N_17303);
nor U18450 (N_18450,N_16772,N_16644);
xnor U18451 (N_18451,N_16703,N_16366);
nand U18452 (N_18452,N_16355,N_16201);
xnor U18453 (N_18453,N_17534,N_17377);
xnor U18454 (N_18454,N_17695,N_16163);
nor U18455 (N_18455,N_16154,N_16391);
nor U18456 (N_18456,N_16138,N_16276);
nand U18457 (N_18457,N_16552,N_17991);
nor U18458 (N_18458,N_16617,N_17371);
and U18459 (N_18459,N_16666,N_16689);
nand U18460 (N_18460,N_16286,N_16164);
nand U18461 (N_18461,N_17369,N_17982);
and U18462 (N_18462,N_17479,N_16694);
nor U18463 (N_18463,N_17859,N_16898);
or U18464 (N_18464,N_17438,N_16495);
nand U18465 (N_18465,N_17478,N_16753);
nor U18466 (N_18466,N_16097,N_17139);
and U18467 (N_18467,N_16279,N_17846);
nand U18468 (N_18468,N_16461,N_16285);
xnor U18469 (N_18469,N_17601,N_16657);
nor U18470 (N_18470,N_16474,N_16022);
or U18471 (N_18471,N_17641,N_16668);
xor U18472 (N_18472,N_16001,N_17998);
and U18473 (N_18473,N_16108,N_17240);
and U18474 (N_18474,N_17836,N_16132);
or U18475 (N_18475,N_16301,N_16526);
xor U18476 (N_18476,N_17352,N_17457);
xnor U18477 (N_18477,N_17990,N_16401);
nor U18478 (N_18478,N_17803,N_17127);
nand U18479 (N_18479,N_17206,N_17975);
nand U18480 (N_18480,N_16244,N_16310);
and U18481 (N_18481,N_17346,N_17737);
nand U18482 (N_18482,N_16349,N_16553);
xor U18483 (N_18483,N_16362,N_17492);
xnor U18484 (N_18484,N_16824,N_16600);
and U18485 (N_18485,N_16709,N_16971);
xnor U18486 (N_18486,N_17037,N_17174);
and U18487 (N_18487,N_17327,N_16639);
or U18488 (N_18488,N_16887,N_16504);
or U18489 (N_18489,N_16383,N_16042);
and U18490 (N_18490,N_17381,N_16188);
and U18491 (N_18491,N_16965,N_16147);
nor U18492 (N_18492,N_17949,N_16169);
nor U18493 (N_18493,N_17362,N_17307);
nand U18494 (N_18494,N_16192,N_16008);
nand U18495 (N_18495,N_17298,N_17931);
or U18496 (N_18496,N_16509,N_17328);
nor U18497 (N_18497,N_16183,N_16718);
xnor U18498 (N_18498,N_17025,N_17160);
xor U18499 (N_18499,N_17914,N_17354);
nor U18500 (N_18500,N_17670,N_16870);
nand U18501 (N_18501,N_17765,N_16830);
xnor U18502 (N_18502,N_17919,N_16724);
nor U18503 (N_18503,N_16988,N_17126);
nand U18504 (N_18504,N_17798,N_16428);
xor U18505 (N_18505,N_16414,N_16612);
or U18506 (N_18506,N_16056,N_17400);
xnor U18507 (N_18507,N_17393,N_16036);
nor U18508 (N_18508,N_17088,N_17439);
and U18509 (N_18509,N_17429,N_17102);
nor U18510 (N_18510,N_17728,N_17748);
xnor U18511 (N_18511,N_16418,N_17865);
nor U18512 (N_18512,N_16333,N_17630);
nor U18513 (N_18513,N_17858,N_17629);
nand U18514 (N_18514,N_17523,N_16518);
and U18515 (N_18515,N_16876,N_17165);
and U18516 (N_18516,N_17255,N_17532);
nor U18517 (N_18517,N_16018,N_17604);
or U18518 (N_18518,N_17273,N_16865);
and U18519 (N_18519,N_17618,N_17636);
nor U18520 (N_18520,N_16589,N_16496);
nand U18521 (N_18521,N_17757,N_17229);
xnor U18522 (N_18522,N_17770,N_17285);
nor U18523 (N_18523,N_17372,N_17761);
nor U18524 (N_18524,N_16466,N_16997);
and U18525 (N_18525,N_17456,N_16781);
xor U18526 (N_18526,N_17407,N_16114);
nor U18527 (N_18527,N_16990,N_17091);
and U18528 (N_18528,N_17714,N_17263);
xnor U18529 (N_18529,N_16127,N_16970);
or U18530 (N_18530,N_17437,N_17173);
or U18531 (N_18531,N_17845,N_16035);
nor U18532 (N_18532,N_16104,N_17746);
or U18533 (N_18533,N_16109,N_16363);
and U18534 (N_18534,N_17614,N_16041);
nand U18535 (N_18535,N_17443,N_16393);
and U18536 (N_18536,N_17073,N_16537);
xor U18537 (N_18537,N_17426,N_17624);
nand U18538 (N_18538,N_17444,N_16130);
or U18539 (N_18539,N_17070,N_16993);
xor U18540 (N_18540,N_17739,N_16294);
nor U18541 (N_18541,N_16062,N_17562);
xor U18542 (N_18542,N_16026,N_16795);
or U18543 (N_18543,N_17147,N_16762);
and U18544 (N_18544,N_17359,N_16543);
or U18545 (N_18545,N_16580,N_16585);
nor U18546 (N_18546,N_17104,N_17186);
nor U18547 (N_18547,N_17881,N_17119);
nand U18548 (N_18548,N_16816,N_17764);
nor U18549 (N_18549,N_16573,N_16774);
and U18550 (N_18550,N_16477,N_16847);
nand U18551 (N_18551,N_17501,N_16356);
or U18552 (N_18552,N_16343,N_17361);
nand U18553 (N_18553,N_17267,N_16548);
xnor U18554 (N_18554,N_17974,N_17221);
nor U18555 (N_18555,N_17502,N_17154);
nand U18556 (N_18556,N_17759,N_17724);
and U18557 (N_18557,N_16895,N_16963);
xnor U18558 (N_18558,N_16064,N_16271);
nand U18559 (N_18559,N_16981,N_16390);
xnor U18560 (N_18560,N_17733,N_16263);
and U18561 (N_18561,N_17414,N_16350);
nor U18562 (N_18562,N_17146,N_17003);
nand U18563 (N_18563,N_16373,N_17503);
or U18564 (N_18564,N_16967,N_16337);
xor U18565 (N_18565,N_17394,N_16852);
and U18566 (N_18566,N_17468,N_17205);
nand U18567 (N_18567,N_16218,N_16320);
xnor U18568 (N_18568,N_16625,N_16860);
and U18569 (N_18569,N_16061,N_17148);
nor U18570 (N_18570,N_16077,N_17570);
nand U18571 (N_18571,N_16960,N_17566);
nor U18572 (N_18572,N_17058,N_17800);
or U18573 (N_18573,N_17932,N_17463);
and U18574 (N_18574,N_16051,N_17725);
and U18575 (N_18575,N_16588,N_16801);
and U18576 (N_18576,N_16754,N_16563);
xnor U18577 (N_18577,N_16406,N_16905);
and U18578 (N_18578,N_16608,N_17023);
xor U18579 (N_18579,N_17945,N_16578);
or U18580 (N_18580,N_17815,N_16733);
or U18581 (N_18581,N_16999,N_17065);
and U18582 (N_18582,N_16980,N_17713);
and U18583 (N_18583,N_17664,N_16913);
nor U18584 (N_18584,N_17202,N_16797);
nor U18585 (N_18585,N_17645,N_17034);
nand U18586 (N_18586,N_17834,N_17036);
nor U18587 (N_18587,N_17827,N_17838);
nor U18588 (N_18588,N_16557,N_17900);
and U18589 (N_18589,N_16723,N_16892);
xnor U18590 (N_18590,N_17390,N_16094);
and U18591 (N_18591,N_16281,N_16974);
nor U18592 (N_18592,N_16502,N_17080);
nand U18593 (N_18593,N_17316,N_16262);
or U18594 (N_18594,N_17684,N_17011);
nor U18595 (N_18595,N_17128,N_16133);
and U18596 (N_18596,N_17768,N_16155);
and U18597 (N_18597,N_16688,N_16142);
xor U18598 (N_18598,N_17196,N_17211);
or U18599 (N_18599,N_17490,N_17214);
nor U18600 (N_18600,N_16918,N_16742);
xor U18601 (N_18601,N_17422,N_16917);
nor U18602 (N_18602,N_17805,N_17284);
or U18603 (N_18603,N_16117,N_16598);
nand U18604 (N_18604,N_17123,N_17715);
nand U18605 (N_18605,N_16111,N_17477);
or U18606 (N_18606,N_17061,N_17166);
and U18607 (N_18607,N_16893,N_16182);
and U18608 (N_18608,N_17323,N_17458);
and U18609 (N_18609,N_17685,N_17996);
xnor U18610 (N_18610,N_17172,N_17665);
or U18611 (N_18611,N_16791,N_17939);
nor U18612 (N_18612,N_17726,N_16661);
and U18613 (N_18613,N_16511,N_16746);
xor U18614 (N_18614,N_17076,N_17004);
nor U18615 (N_18615,N_16749,N_16787);
or U18616 (N_18616,N_17238,N_17232);
and U18617 (N_18617,N_17877,N_17258);
xor U18618 (N_18618,N_17649,N_16584);
xor U18619 (N_18619,N_17605,N_17968);
and U18620 (N_18620,N_17702,N_17952);
nand U18621 (N_18621,N_16014,N_17249);
xnor U18622 (N_18622,N_16028,N_17844);
nand U18623 (N_18623,N_17062,N_16962);
nand U18624 (N_18624,N_17343,N_16912);
and U18625 (N_18625,N_16596,N_17938);
and U18626 (N_18626,N_16894,N_16409);
nor U18627 (N_18627,N_17380,N_17452);
or U18628 (N_18628,N_16484,N_17068);
nand U18629 (N_18629,N_16069,N_17505);
xnor U18630 (N_18630,N_16562,N_16040);
and U18631 (N_18631,N_17799,N_16926);
and U18632 (N_18632,N_17475,N_17760);
nand U18633 (N_18633,N_16181,N_17655);
nor U18634 (N_18634,N_16334,N_16378);
and U18635 (N_18635,N_17459,N_16102);
xnor U18636 (N_18636,N_16677,N_17158);
xnor U18637 (N_18637,N_16328,N_17317);
xnor U18638 (N_18638,N_16200,N_16460);
xnor U18639 (N_18639,N_17890,N_17571);
and U18640 (N_18640,N_16998,N_16275);
and U18641 (N_18641,N_16909,N_17107);
xor U18642 (N_18642,N_17893,N_16080);
nand U18643 (N_18643,N_17786,N_17712);
and U18644 (N_18644,N_16811,N_16506);
nor U18645 (N_18645,N_17079,N_16039);
xnor U18646 (N_18646,N_16706,N_16068);
and U18647 (N_18647,N_17187,N_16785);
or U18648 (N_18648,N_17696,N_17131);
xnor U18649 (N_18649,N_17271,N_17375);
xor U18650 (N_18650,N_16558,N_17292);
nand U18651 (N_18651,N_17231,N_17424);
nand U18652 (N_18652,N_16943,N_17178);
nand U18653 (N_18653,N_17552,N_17470);
nand U18654 (N_18654,N_17269,N_17455);
or U18655 (N_18655,N_17668,N_17547);
or U18656 (N_18656,N_17309,N_16944);
and U18657 (N_18657,N_16128,N_16857);
and U18658 (N_18658,N_17563,N_17988);
nor U18659 (N_18659,N_17753,N_16024);
nand U18660 (N_18660,N_16497,N_16199);
xnor U18661 (N_18661,N_17197,N_16750);
xor U18662 (N_18662,N_17460,N_16872);
xnor U18663 (N_18663,N_17449,N_17066);
xor U18664 (N_18664,N_16386,N_17663);
nand U18665 (N_18665,N_16508,N_16833);
nor U18666 (N_18666,N_16678,N_17687);
or U18667 (N_18667,N_16327,N_17498);
or U18668 (N_18668,N_16178,N_16398);
or U18669 (N_18669,N_16660,N_17979);
xnor U18670 (N_18670,N_17905,N_17201);
nand U18671 (N_18671,N_17351,N_16621);
nand U18672 (N_18672,N_17474,N_16050);
or U18673 (N_18673,N_17276,N_16419);
nand U18674 (N_18674,N_16442,N_17808);
nand U18675 (N_18675,N_16848,N_16168);
nor U18676 (N_18676,N_17026,N_17690);
or U18677 (N_18677,N_17409,N_17542);
and U18678 (N_18678,N_17193,N_17648);
nand U18679 (N_18679,N_16283,N_16241);
xnor U18680 (N_18680,N_16267,N_17310);
nand U18681 (N_18681,N_16458,N_16702);
xnor U18682 (N_18682,N_17810,N_17428);
nor U18683 (N_18683,N_16634,N_16858);
or U18684 (N_18684,N_16662,N_17342);
nor U18685 (N_18685,N_16376,N_16043);
or U18686 (N_18686,N_17718,N_17028);
nand U18687 (N_18687,N_17772,N_16594);
xor U18688 (N_18688,N_17581,N_17545);
or U18689 (N_18689,N_16131,N_16534);
nor U18690 (N_18690,N_17600,N_16326);
nand U18691 (N_18691,N_16059,N_17301);
or U18692 (N_18692,N_17225,N_17415);
or U18693 (N_18693,N_17432,N_16956);
and U18694 (N_18694,N_16437,N_17778);
nor U18695 (N_18695,N_16582,N_16211);
and U18696 (N_18696,N_17100,N_16485);
or U18697 (N_18697,N_17891,N_17071);
xor U18698 (N_18698,N_17850,N_16710);
or U18699 (N_18699,N_16089,N_17304);
and U18700 (N_18700,N_16402,N_17612);
nor U18701 (N_18701,N_16249,N_16044);
and U18702 (N_18702,N_16236,N_17809);
and U18703 (N_18703,N_17367,N_17485);
or U18704 (N_18704,N_16796,N_17251);
nand U18705 (N_18705,N_16227,N_16882);
xor U18706 (N_18706,N_17199,N_16284);
nor U18707 (N_18707,N_16664,N_17506);
or U18708 (N_18708,N_17256,N_16239);
or U18709 (N_18709,N_17082,N_16424);
nor U18710 (N_18710,N_17017,N_17634);
or U18711 (N_18711,N_16812,N_17854);
xnor U18712 (N_18712,N_17876,N_16802);
xnor U18713 (N_18713,N_17427,N_17843);
xnor U18714 (N_18714,N_16298,N_17969);
nor U18715 (N_18715,N_17699,N_16313);
xnor U18716 (N_18716,N_17486,N_16293);
and U18717 (N_18717,N_17210,N_17959);
xor U18718 (N_18718,N_16150,N_16880);
and U18719 (N_18719,N_16991,N_16342);
xor U18720 (N_18720,N_17116,N_17313);
and U18721 (N_18721,N_17504,N_16734);
nand U18722 (N_18722,N_16137,N_17320);
nor U18723 (N_18723,N_16291,N_17933);
nand U18724 (N_18724,N_16659,N_16979);
nor U18725 (N_18725,N_16380,N_17957);
and U18726 (N_18726,N_16503,N_17226);
or U18727 (N_18727,N_17308,N_16251);
xnor U18728 (N_18728,N_17946,N_16222);
and U18729 (N_18729,N_16210,N_16453);
or U18730 (N_18730,N_16571,N_16853);
xnor U18731 (N_18731,N_16482,N_17565);
and U18732 (N_18732,N_16308,N_17840);
nand U18733 (N_18733,N_17039,N_17217);
and U18734 (N_18734,N_16692,N_16606);
or U18735 (N_18735,N_17234,N_16957);
nor U18736 (N_18736,N_17250,N_17137);
nand U18737 (N_18737,N_17745,N_16447);
nand U18738 (N_18738,N_16761,N_17331);
and U18739 (N_18739,N_16984,N_17222);
or U18740 (N_18740,N_17930,N_17476);
nand U18741 (N_18741,N_16842,N_16701);
or U18742 (N_18742,N_16616,N_17856);
or U18743 (N_18743,N_16951,N_17693);
and U18744 (N_18744,N_17878,N_17355);
nand U18745 (N_18745,N_16246,N_16093);
or U18746 (N_18746,N_17584,N_17766);
nand U18747 (N_18747,N_16417,N_17130);
or U18748 (N_18748,N_17682,N_16037);
or U18749 (N_18749,N_16717,N_16045);
nor U18750 (N_18750,N_17401,N_17965);
and U18751 (N_18751,N_17108,N_17266);
nand U18752 (N_18752,N_16650,N_17971);
and U18753 (N_18753,N_16480,N_16318);
xnor U18754 (N_18754,N_16413,N_16599);
or U18755 (N_18755,N_17305,N_16682);
nor U18756 (N_18756,N_17675,N_16790);
xor U18757 (N_18757,N_16116,N_16226);
nor U18758 (N_18758,N_17364,N_16758);
nand U18759 (N_18759,N_17828,N_16422);
and U18760 (N_18760,N_16085,N_16757);
nor U18761 (N_18761,N_16766,N_16209);
xnor U18762 (N_18762,N_17511,N_17863);
nor U18763 (N_18763,N_16314,N_16986);
nor U18764 (N_18764,N_17610,N_17824);
nand U18765 (N_18765,N_16494,N_17587);
nand U18766 (N_18766,N_17125,N_16516);
nand U18767 (N_18767,N_16225,N_16113);
or U18768 (N_18768,N_17895,N_16615);
and U18769 (N_18769,N_16144,N_16204);
xor U18770 (N_18770,N_16958,N_16420);
nor U18771 (N_18771,N_17688,N_17632);
or U18772 (N_18772,N_16649,N_17609);
and U18773 (N_18773,N_16861,N_17338);
xnor U18774 (N_18774,N_17454,N_17030);
nor U18775 (N_18775,N_17348,N_16779);
and U18776 (N_18776,N_17257,N_16500);
or U18777 (N_18777,N_17085,N_16387);
xor U18778 (N_18778,N_16623,N_16897);
xor U18779 (N_18779,N_17911,N_17001);
nand U18780 (N_18780,N_16083,N_17434);
nand U18781 (N_18781,N_16309,N_16498);
and U18782 (N_18782,N_16510,N_17220);
or U18783 (N_18783,N_17678,N_17925);
nor U18784 (N_18784,N_16687,N_16592);
nand U18785 (N_18785,N_17115,N_16513);
or U18786 (N_18786,N_17575,N_16492);
xor U18787 (N_18787,N_16486,N_16020);
and U18788 (N_18788,N_16140,N_17825);
or U18789 (N_18789,N_17788,N_17597);
or U18790 (N_18790,N_16684,N_17951);
nand U18791 (N_18791,N_17318,N_17495);
or U18792 (N_18792,N_17642,N_16034);
nor U18793 (N_18793,N_16839,N_17638);
nor U18794 (N_18794,N_17382,N_17000);
nor U18795 (N_18795,N_16125,N_17014);
xor U18796 (N_18796,N_16550,N_16289);
nand U18797 (N_18797,N_16021,N_17561);
and U18798 (N_18798,N_16074,N_16217);
nor U18799 (N_18799,N_17514,N_16748);
or U18800 (N_18800,N_17219,N_17673);
xor U18801 (N_18801,N_17883,N_16629);
nand U18802 (N_18802,N_17435,N_17588);
nor U18803 (N_18803,N_16646,N_17622);
xor U18804 (N_18804,N_17365,N_16556);
nand U18805 (N_18805,N_17592,N_17559);
or U18806 (N_18806,N_17874,N_16907);
xnor U18807 (N_18807,N_17374,N_16782);
xor U18808 (N_18808,N_16632,N_16529);
or U18809 (N_18809,N_16431,N_17244);
or U18810 (N_18810,N_16449,N_17350);
xnor U18811 (N_18811,N_17683,N_17252);
xor U18812 (N_18812,N_16296,N_17691);
or U18813 (N_18813,N_16875,N_16176);
nor U18814 (N_18814,N_16455,N_17515);
nand U18815 (N_18815,N_16891,N_17616);
xnor U18816 (N_18816,N_16524,N_17972);
or U18817 (N_18817,N_17628,N_16531);
nor U18818 (N_18818,N_17767,N_16121);
nor U18819 (N_18819,N_16725,N_16195);
xor U18820 (N_18820,N_16385,N_17213);
or U18821 (N_18821,N_16512,N_17658);
xnor U18822 (N_18822,N_17777,N_17056);
nand U18823 (N_18823,N_17020,N_16959);
nor U18824 (N_18824,N_17672,N_16635);
and U18825 (N_18825,N_16476,N_17698);
or U18826 (N_18826,N_16397,N_17293);
xnor U18827 (N_18827,N_16073,N_17954);
or U18828 (N_18828,N_16143,N_17420);
or U18829 (N_18829,N_16522,N_16475);
or U18830 (N_18830,N_16180,N_17009);
nand U18831 (N_18831,N_16914,N_17904);
nor U18832 (N_18832,N_16174,N_16982);
and U18833 (N_18833,N_16187,N_17280);
nand U18834 (N_18834,N_16919,N_17533);
nand U18835 (N_18835,N_17519,N_17484);
nor U18836 (N_18836,N_16429,N_17985);
xnor U18837 (N_18837,N_17711,N_16846);
or U18838 (N_18838,N_16213,N_16219);
xor U18839 (N_18839,N_16685,N_17411);
xor U18840 (N_18840,N_17184,N_17247);
nand U18841 (N_18841,N_16595,N_16538);
nor U18842 (N_18842,N_16238,N_17716);
nand U18843 (N_18843,N_17615,N_16151);
xor U18844 (N_18844,N_16123,N_16633);
and U18845 (N_18845,N_17705,N_16886);
xnor U18846 (N_18846,N_16551,N_16071);
or U18847 (N_18847,N_16186,N_16916);
nand U18848 (N_18848,N_16208,N_16395);
xor U18849 (N_18849,N_16099,N_17453);
nor U18850 (N_18850,N_17729,N_17861);
nand U18851 (N_18851,N_17626,N_16669);
nand U18852 (N_18852,N_16258,N_16843);
nor U18853 (N_18853,N_17194,N_17322);
and U18854 (N_18854,N_17973,N_16803);
or U18855 (N_18855,N_16716,N_16747);
or U18856 (N_18856,N_16840,N_17399);
nor U18857 (N_18857,N_17153,N_16049);
nand U18858 (N_18858,N_16707,N_17842);
and U18859 (N_18859,N_17208,N_16611);
and U18860 (N_18860,N_17594,N_16873);
nand U18861 (N_18861,N_16237,N_17171);
nand U18862 (N_18862,N_17578,N_17964);
nand U18863 (N_18863,N_17010,N_17689);
xnor U18864 (N_18864,N_17817,N_16245);
and U18865 (N_18865,N_16877,N_16322);
nor U18866 (N_18866,N_16784,N_17357);
and U18867 (N_18867,N_17583,N_16290);
xor U18868 (N_18868,N_17356,N_17829);
or U18869 (N_18869,N_16532,N_16767);
nand U18870 (N_18870,N_17282,N_16627);
or U18871 (N_18871,N_17179,N_17141);
nand U18872 (N_18872,N_17579,N_16903);
xnor U18873 (N_18873,N_16820,N_16162);
nor U18874 (N_18874,N_16469,N_16084);
nand U18875 (N_18875,N_16869,N_16514);
or U18876 (N_18876,N_16344,N_17732);
or U18877 (N_18877,N_16699,N_16642);
or U18878 (N_18878,N_16732,N_17652);
nand U18879 (N_18879,N_16394,N_16630);
nor U18880 (N_18880,N_16832,N_16808);
nor U18881 (N_18881,N_17763,N_17341);
xor U18882 (N_18882,N_17538,N_17488);
nand U18883 (N_18883,N_16425,N_17525);
nor U18884 (N_18884,N_16231,N_16396);
nor U18885 (N_18885,N_16005,N_16184);
xnor U18886 (N_18886,N_16441,N_17822);
nand U18887 (N_18887,N_16793,N_17585);
nor U18888 (N_18888,N_17086,N_17771);
nand U18889 (N_18889,N_17300,N_17151);
nand U18890 (N_18890,N_16191,N_16910);
and U18891 (N_18891,N_17654,N_16415);
xnor U18892 (N_18892,N_17081,N_17902);
nor U18893 (N_18893,N_17319,N_17709);
xor U18894 (N_18894,N_17315,N_17762);
xnor U18895 (N_18895,N_17882,N_17124);
or U18896 (N_18896,N_17819,N_16564);
and U18897 (N_18897,N_16605,N_16472);
and U18898 (N_18898,N_16032,N_16773);
xor U18899 (N_18899,N_16107,N_16078);
nor U18900 (N_18900,N_17012,N_17674);
and U18901 (N_18901,N_16978,N_17261);
nor U18902 (N_18902,N_17706,N_17324);
or U18903 (N_18903,N_16338,N_16771);
nand U18904 (N_18904,N_17921,N_16110);
nor U18905 (N_18905,N_16302,N_16996);
nand U18906 (N_18906,N_16030,N_17236);
and U18907 (N_18907,N_16624,N_16735);
nor U18908 (N_18908,N_16003,N_17383);
or U18909 (N_18909,N_16579,N_16940);
nor U18910 (N_18910,N_17789,N_16399);
nand U18911 (N_18911,N_17177,N_16973);
or U18912 (N_18912,N_16822,N_16010);
nor U18913 (N_18913,N_16126,N_17967);
xnor U18914 (N_18914,N_16243,N_16365);
xor U18915 (N_18915,N_17787,N_16713);
nand U18916 (N_18916,N_17551,N_17195);
or U18917 (N_18917,N_16798,N_17133);
or U18918 (N_18918,N_16324,N_16786);
and U18919 (N_18919,N_17140,N_17022);
or U18920 (N_18920,N_16374,N_17431);
nor U18921 (N_18921,N_17927,N_16505);
or U18922 (N_18922,N_17103,N_16539);
xnor U18923 (N_18923,N_16065,N_17942);
nand U18924 (N_18924,N_16560,N_17801);
nor U18925 (N_18925,N_16866,N_17812);
nor U18926 (N_18926,N_17918,N_17283);
nor U18927 (N_18927,N_17741,N_17425);
nor U18928 (N_18928,N_17755,N_17520);
or U18929 (N_18929,N_16992,N_17033);
xor U18930 (N_18930,N_17731,N_16565);
or U18931 (N_18931,N_16520,N_16889);
or U18932 (N_18932,N_16648,N_17499);
nand U18933 (N_18933,N_16647,N_16711);
nor U18934 (N_18934,N_16862,N_16952);
or U18935 (N_18935,N_16221,N_17223);
nor U18936 (N_18936,N_17090,N_17872);
xnor U18937 (N_18937,N_16323,N_17159);
or U18938 (N_18938,N_17321,N_16193);
nor U18939 (N_18939,N_16964,N_17886);
or U18940 (N_18940,N_16136,N_16708);
and U18941 (N_18941,N_16906,N_17512);
nand U18942 (N_18942,N_17006,N_17472);
xor U18943 (N_18943,N_16731,N_17866);
nand U18944 (N_18944,N_16545,N_16471);
xnor U18945 (N_18945,N_17667,N_16481);
xor U18946 (N_18946,N_16158,N_16995);
xnor U18947 (N_18947,N_16501,N_16341);
nand U18948 (N_18948,N_17736,N_16354);
xor U18949 (N_18949,N_17278,N_16253);
nand U18950 (N_18950,N_17368,N_17517);
and U18951 (N_18951,N_16755,N_17314);
or U18952 (N_18952,N_16902,N_17831);
or U18953 (N_18953,N_17132,N_16572);
nand U18954 (N_18954,N_17032,N_17920);
or U18955 (N_18955,N_16129,N_17281);
xnor U18956 (N_18956,N_16546,N_16079);
xor U18957 (N_18957,N_17096,N_16775);
nand U18958 (N_18958,N_17121,N_17289);
nand U18959 (N_18959,N_17701,N_17669);
and U18960 (N_18960,N_16017,N_17833);
nand U18961 (N_18961,N_16954,N_17910);
and U18962 (N_18962,N_16160,N_17580);
and U18963 (N_18963,N_17521,N_16004);
nor U18964 (N_18964,N_17666,N_16312);
nand U18965 (N_18965,N_17889,N_16330);
nand U18966 (N_18966,N_17958,N_16172);
and U18967 (N_18967,N_17167,N_16170);
xnor U18968 (N_18968,N_17312,N_17591);
or U18969 (N_18969,N_16141,N_17744);
xnor U18970 (N_18970,N_16680,N_16335);
and U18971 (N_18971,N_17421,N_17207);
and U18972 (N_18972,N_16000,N_16697);
or U18973 (N_18973,N_17613,N_17922);
nand U18974 (N_18974,N_17807,N_17209);
xnor U18975 (N_18975,N_17134,N_17268);
or U18976 (N_18976,N_17832,N_16836);
or U18977 (N_18977,N_16626,N_16770);
xnor U18978 (N_18978,N_17966,N_16315);
nand U18979 (N_18979,N_16346,N_16817);
xnor U18980 (N_18980,N_17347,N_16408);
and U18981 (N_18981,N_17862,N_16527);
nand U18982 (N_18982,N_17619,N_17947);
nor U18983 (N_18983,N_17811,N_16433);
or U18984 (N_18984,N_16002,N_17924);
xor U18985 (N_18985,N_17094,N_17980);
or U18986 (N_18986,N_17135,N_17007);
xnor U18987 (N_18987,N_17487,N_17536);
xor U18988 (N_18988,N_16031,N_17049);
or U18989 (N_18989,N_17168,N_16081);
nor U18990 (N_18990,N_17180,N_17795);
nor U18991 (N_18991,N_17050,N_17750);
and U18992 (N_18992,N_17340,N_17680);
nor U18993 (N_18993,N_16517,N_16473);
nand U18994 (N_18994,N_17333,N_17063);
nor U18995 (N_18995,N_16728,N_16105);
or U18996 (N_18996,N_16305,N_16783);
and U18997 (N_18997,N_16261,N_16054);
xnor U18998 (N_18998,N_17986,N_16935);
and U18999 (N_18999,N_17326,N_16052);
nand U19000 (N_19000,N_16414,N_17511);
nand U19001 (N_19001,N_17520,N_17803);
xor U19002 (N_19002,N_16644,N_16914);
nand U19003 (N_19003,N_17115,N_17222);
and U19004 (N_19004,N_16908,N_16309);
xor U19005 (N_19005,N_17168,N_16449);
nand U19006 (N_19006,N_16792,N_17988);
xor U19007 (N_19007,N_16128,N_16461);
and U19008 (N_19008,N_17274,N_16354);
xor U19009 (N_19009,N_17218,N_16375);
nand U19010 (N_19010,N_17197,N_16867);
xnor U19011 (N_19011,N_17664,N_16483);
and U19012 (N_19012,N_16245,N_17376);
nand U19013 (N_19013,N_17131,N_17577);
xor U19014 (N_19014,N_16864,N_17750);
xnor U19015 (N_19015,N_16099,N_17331);
nand U19016 (N_19016,N_16446,N_17059);
and U19017 (N_19017,N_16621,N_17250);
and U19018 (N_19018,N_17781,N_16663);
nand U19019 (N_19019,N_17517,N_17604);
nor U19020 (N_19020,N_16678,N_17442);
nor U19021 (N_19021,N_17959,N_16595);
nand U19022 (N_19022,N_17217,N_16361);
xor U19023 (N_19023,N_16384,N_17409);
or U19024 (N_19024,N_17472,N_16246);
and U19025 (N_19025,N_16607,N_17310);
nand U19026 (N_19026,N_16324,N_16929);
or U19027 (N_19027,N_17403,N_16369);
nor U19028 (N_19028,N_17661,N_17811);
and U19029 (N_19029,N_17156,N_17077);
and U19030 (N_19030,N_17966,N_17881);
nand U19031 (N_19031,N_16261,N_16080);
nor U19032 (N_19032,N_16584,N_16360);
and U19033 (N_19033,N_16178,N_17707);
or U19034 (N_19034,N_17934,N_17969);
nor U19035 (N_19035,N_17028,N_16713);
or U19036 (N_19036,N_16763,N_17489);
nand U19037 (N_19037,N_16619,N_16453);
or U19038 (N_19038,N_16249,N_16795);
and U19039 (N_19039,N_17539,N_17205);
xnor U19040 (N_19040,N_16879,N_17400);
or U19041 (N_19041,N_17507,N_17708);
xor U19042 (N_19042,N_16033,N_17837);
nand U19043 (N_19043,N_17392,N_16753);
or U19044 (N_19044,N_17216,N_17505);
xor U19045 (N_19045,N_16744,N_17406);
nand U19046 (N_19046,N_16448,N_17373);
and U19047 (N_19047,N_16818,N_17260);
and U19048 (N_19048,N_16845,N_17266);
or U19049 (N_19049,N_16702,N_17155);
xnor U19050 (N_19050,N_17416,N_16192);
or U19051 (N_19051,N_17276,N_16086);
nand U19052 (N_19052,N_16333,N_17415);
or U19053 (N_19053,N_16268,N_16620);
xnor U19054 (N_19054,N_17900,N_17065);
or U19055 (N_19055,N_16240,N_16373);
and U19056 (N_19056,N_16067,N_17457);
nand U19057 (N_19057,N_17560,N_16674);
or U19058 (N_19058,N_17312,N_17465);
xnor U19059 (N_19059,N_17867,N_17668);
and U19060 (N_19060,N_17590,N_17910);
nor U19061 (N_19061,N_16412,N_16452);
and U19062 (N_19062,N_16171,N_17233);
or U19063 (N_19063,N_16563,N_17962);
or U19064 (N_19064,N_16990,N_16840);
or U19065 (N_19065,N_16937,N_17952);
and U19066 (N_19066,N_17711,N_16078);
or U19067 (N_19067,N_17769,N_16893);
or U19068 (N_19068,N_16455,N_16324);
or U19069 (N_19069,N_17711,N_17125);
nand U19070 (N_19070,N_16640,N_17594);
nand U19071 (N_19071,N_17705,N_17145);
xnor U19072 (N_19072,N_16635,N_16164);
nand U19073 (N_19073,N_17590,N_16377);
xor U19074 (N_19074,N_17202,N_17568);
nor U19075 (N_19075,N_17787,N_16036);
nor U19076 (N_19076,N_16661,N_17579);
or U19077 (N_19077,N_17356,N_17497);
and U19078 (N_19078,N_16171,N_17338);
nand U19079 (N_19079,N_16398,N_16597);
or U19080 (N_19080,N_17792,N_17045);
xor U19081 (N_19081,N_16853,N_17818);
nor U19082 (N_19082,N_16046,N_17522);
or U19083 (N_19083,N_16131,N_16376);
and U19084 (N_19084,N_17333,N_16790);
xnor U19085 (N_19085,N_16823,N_16799);
nor U19086 (N_19086,N_16982,N_17955);
or U19087 (N_19087,N_16873,N_17993);
xnor U19088 (N_19088,N_17809,N_16145);
nor U19089 (N_19089,N_17901,N_17611);
and U19090 (N_19090,N_16663,N_17704);
or U19091 (N_19091,N_16238,N_16788);
nor U19092 (N_19092,N_16371,N_16930);
nor U19093 (N_19093,N_17049,N_16781);
and U19094 (N_19094,N_16973,N_17618);
xnor U19095 (N_19095,N_16482,N_16750);
nor U19096 (N_19096,N_16939,N_16371);
and U19097 (N_19097,N_17996,N_16595);
xnor U19098 (N_19098,N_17175,N_17854);
nand U19099 (N_19099,N_16590,N_17965);
or U19100 (N_19100,N_16546,N_17357);
nand U19101 (N_19101,N_16991,N_16382);
nand U19102 (N_19102,N_16934,N_17715);
or U19103 (N_19103,N_16854,N_16063);
xnor U19104 (N_19104,N_16368,N_17029);
nor U19105 (N_19105,N_16550,N_17648);
and U19106 (N_19106,N_17789,N_16929);
and U19107 (N_19107,N_17937,N_17843);
xor U19108 (N_19108,N_16260,N_17849);
xor U19109 (N_19109,N_16025,N_16114);
nand U19110 (N_19110,N_17511,N_16914);
or U19111 (N_19111,N_16281,N_16314);
nand U19112 (N_19112,N_17675,N_16903);
xor U19113 (N_19113,N_16821,N_17848);
or U19114 (N_19114,N_17415,N_16647);
xor U19115 (N_19115,N_17444,N_16772);
nor U19116 (N_19116,N_17096,N_16015);
or U19117 (N_19117,N_17668,N_16746);
or U19118 (N_19118,N_17983,N_17433);
nand U19119 (N_19119,N_16646,N_17777);
nand U19120 (N_19120,N_17639,N_16449);
nor U19121 (N_19121,N_16200,N_17630);
nand U19122 (N_19122,N_17743,N_16297);
or U19123 (N_19123,N_17886,N_17645);
and U19124 (N_19124,N_16219,N_17408);
and U19125 (N_19125,N_16093,N_17931);
nand U19126 (N_19126,N_17090,N_16295);
or U19127 (N_19127,N_16264,N_16950);
nand U19128 (N_19128,N_17506,N_16338);
xor U19129 (N_19129,N_17816,N_16368);
xnor U19130 (N_19130,N_17112,N_16589);
and U19131 (N_19131,N_17155,N_16062);
nor U19132 (N_19132,N_16873,N_17812);
nand U19133 (N_19133,N_17431,N_16836);
nor U19134 (N_19134,N_17307,N_17405);
or U19135 (N_19135,N_16178,N_17946);
nor U19136 (N_19136,N_17564,N_17635);
nand U19137 (N_19137,N_17901,N_17706);
nand U19138 (N_19138,N_17711,N_17136);
nand U19139 (N_19139,N_17936,N_16827);
nor U19140 (N_19140,N_17614,N_16443);
nand U19141 (N_19141,N_17906,N_17160);
nand U19142 (N_19142,N_16511,N_17891);
nand U19143 (N_19143,N_16786,N_17113);
nand U19144 (N_19144,N_17952,N_17814);
or U19145 (N_19145,N_17942,N_16599);
nand U19146 (N_19146,N_16178,N_16176);
nor U19147 (N_19147,N_16976,N_16558);
xor U19148 (N_19148,N_17540,N_16170);
nand U19149 (N_19149,N_17004,N_16256);
nor U19150 (N_19150,N_16082,N_17485);
or U19151 (N_19151,N_17257,N_16002);
and U19152 (N_19152,N_17195,N_16875);
or U19153 (N_19153,N_17434,N_17925);
xnor U19154 (N_19154,N_16753,N_16445);
and U19155 (N_19155,N_16133,N_16482);
or U19156 (N_19156,N_17663,N_17937);
nor U19157 (N_19157,N_16638,N_17522);
nor U19158 (N_19158,N_16025,N_16031);
nand U19159 (N_19159,N_16865,N_17798);
nor U19160 (N_19160,N_17278,N_16357);
nor U19161 (N_19161,N_16363,N_16074);
nor U19162 (N_19162,N_16208,N_17105);
and U19163 (N_19163,N_16088,N_16606);
and U19164 (N_19164,N_17776,N_16435);
nor U19165 (N_19165,N_17895,N_17883);
xnor U19166 (N_19166,N_16728,N_17120);
and U19167 (N_19167,N_16653,N_16779);
nand U19168 (N_19168,N_16972,N_17670);
nor U19169 (N_19169,N_16965,N_16761);
and U19170 (N_19170,N_17615,N_16932);
nor U19171 (N_19171,N_16390,N_17007);
or U19172 (N_19172,N_17793,N_17166);
nand U19173 (N_19173,N_16060,N_16669);
nor U19174 (N_19174,N_16198,N_17223);
nand U19175 (N_19175,N_17251,N_16689);
and U19176 (N_19176,N_17041,N_17953);
nor U19177 (N_19177,N_17096,N_17583);
or U19178 (N_19178,N_16666,N_16809);
nor U19179 (N_19179,N_16454,N_17235);
nand U19180 (N_19180,N_17202,N_16688);
and U19181 (N_19181,N_17333,N_17092);
nand U19182 (N_19182,N_16303,N_16813);
xnor U19183 (N_19183,N_17183,N_16061);
xnor U19184 (N_19184,N_17833,N_16943);
nor U19185 (N_19185,N_16597,N_16698);
or U19186 (N_19186,N_16939,N_16735);
or U19187 (N_19187,N_16165,N_17270);
nand U19188 (N_19188,N_17225,N_17056);
or U19189 (N_19189,N_17546,N_16630);
or U19190 (N_19190,N_16334,N_16451);
nand U19191 (N_19191,N_16885,N_17049);
or U19192 (N_19192,N_16296,N_16498);
and U19193 (N_19193,N_17821,N_16797);
and U19194 (N_19194,N_17995,N_16109);
xor U19195 (N_19195,N_17727,N_16423);
nand U19196 (N_19196,N_16168,N_17125);
xnor U19197 (N_19197,N_16628,N_16119);
xnor U19198 (N_19198,N_17915,N_16180);
and U19199 (N_19199,N_17531,N_16988);
nand U19200 (N_19200,N_17800,N_17391);
and U19201 (N_19201,N_17911,N_17198);
xor U19202 (N_19202,N_17340,N_16981);
nand U19203 (N_19203,N_16136,N_16390);
nor U19204 (N_19204,N_16377,N_17505);
nand U19205 (N_19205,N_16359,N_17368);
xnor U19206 (N_19206,N_17296,N_17210);
and U19207 (N_19207,N_16302,N_17746);
nor U19208 (N_19208,N_17501,N_16670);
xnor U19209 (N_19209,N_17568,N_16640);
or U19210 (N_19210,N_16059,N_16434);
nor U19211 (N_19211,N_17562,N_16064);
nor U19212 (N_19212,N_16784,N_17905);
or U19213 (N_19213,N_16368,N_16302);
nand U19214 (N_19214,N_16193,N_17891);
nor U19215 (N_19215,N_17244,N_17279);
nor U19216 (N_19216,N_17169,N_16500);
nor U19217 (N_19217,N_16359,N_16155);
nor U19218 (N_19218,N_16256,N_17851);
nand U19219 (N_19219,N_16653,N_17084);
and U19220 (N_19220,N_17752,N_16317);
nand U19221 (N_19221,N_16180,N_17928);
nor U19222 (N_19222,N_17838,N_17072);
nand U19223 (N_19223,N_17504,N_16456);
or U19224 (N_19224,N_17095,N_16870);
nor U19225 (N_19225,N_16150,N_17717);
or U19226 (N_19226,N_16353,N_16922);
nand U19227 (N_19227,N_16279,N_17876);
and U19228 (N_19228,N_16171,N_17939);
and U19229 (N_19229,N_16739,N_17269);
xor U19230 (N_19230,N_16774,N_16771);
xor U19231 (N_19231,N_17577,N_16004);
and U19232 (N_19232,N_17455,N_17704);
xor U19233 (N_19233,N_16626,N_16239);
and U19234 (N_19234,N_16078,N_17884);
nor U19235 (N_19235,N_17692,N_17420);
nor U19236 (N_19236,N_17165,N_17935);
and U19237 (N_19237,N_16076,N_17317);
and U19238 (N_19238,N_17743,N_17546);
nand U19239 (N_19239,N_17308,N_17547);
nand U19240 (N_19240,N_17508,N_16275);
xnor U19241 (N_19241,N_17334,N_17596);
and U19242 (N_19242,N_17379,N_16971);
xor U19243 (N_19243,N_16921,N_17834);
or U19244 (N_19244,N_17255,N_16110);
nor U19245 (N_19245,N_16160,N_16576);
nand U19246 (N_19246,N_17186,N_16384);
xnor U19247 (N_19247,N_17489,N_17992);
xor U19248 (N_19248,N_16182,N_17232);
nand U19249 (N_19249,N_16417,N_16584);
and U19250 (N_19250,N_16895,N_17849);
nand U19251 (N_19251,N_16335,N_17481);
nand U19252 (N_19252,N_16057,N_17777);
xor U19253 (N_19253,N_17522,N_16271);
nor U19254 (N_19254,N_16636,N_17832);
xor U19255 (N_19255,N_17157,N_16498);
and U19256 (N_19256,N_17436,N_16657);
and U19257 (N_19257,N_16975,N_16121);
xnor U19258 (N_19258,N_16176,N_17198);
or U19259 (N_19259,N_17302,N_16941);
or U19260 (N_19260,N_17967,N_17438);
nor U19261 (N_19261,N_16961,N_16548);
or U19262 (N_19262,N_17045,N_16674);
or U19263 (N_19263,N_16013,N_16160);
nand U19264 (N_19264,N_16641,N_16912);
or U19265 (N_19265,N_16871,N_17468);
nand U19266 (N_19266,N_17136,N_17771);
nor U19267 (N_19267,N_17587,N_16045);
nand U19268 (N_19268,N_17234,N_17470);
nand U19269 (N_19269,N_17236,N_16662);
and U19270 (N_19270,N_16631,N_16925);
or U19271 (N_19271,N_17384,N_16517);
xnor U19272 (N_19272,N_17545,N_17613);
xor U19273 (N_19273,N_16659,N_16178);
or U19274 (N_19274,N_16233,N_16416);
xor U19275 (N_19275,N_16881,N_16191);
and U19276 (N_19276,N_17943,N_17975);
and U19277 (N_19277,N_17827,N_16238);
xnor U19278 (N_19278,N_17355,N_16472);
nor U19279 (N_19279,N_16518,N_16805);
nand U19280 (N_19280,N_16139,N_16074);
xnor U19281 (N_19281,N_16437,N_17670);
xnor U19282 (N_19282,N_17974,N_16914);
xor U19283 (N_19283,N_17651,N_17435);
xnor U19284 (N_19284,N_17211,N_16766);
and U19285 (N_19285,N_17563,N_17396);
or U19286 (N_19286,N_17902,N_16291);
xor U19287 (N_19287,N_16112,N_17078);
nor U19288 (N_19288,N_16303,N_16079);
or U19289 (N_19289,N_16697,N_16596);
nand U19290 (N_19290,N_16360,N_16374);
and U19291 (N_19291,N_17146,N_17894);
nor U19292 (N_19292,N_17050,N_16216);
or U19293 (N_19293,N_17385,N_17169);
xnor U19294 (N_19294,N_16546,N_17579);
or U19295 (N_19295,N_16002,N_17476);
nor U19296 (N_19296,N_16718,N_16477);
nor U19297 (N_19297,N_16841,N_17336);
xor U19298 (N_19298,N_16398,N_16332);
nand U19299 (N_19299,N_17696,N_16229);
xor U19300 (N_19300,N_17909,N_17325);
nand U19301 (N_19301,N_17471,N_17461);
and U19302 (N_19302,N_16201,N_16871);
and U19303 (N_19303,N_17383,N_16258);
nor U19304 (N_19304,N_16950,N_17800);
xor U19305 (N_19305,N_17776,N_17758);
nand U19306 (N_19306,N_16304,N_16110);
xnor U19307 (N_19307,N_16883,N_16696);
and U19308 (N_19308,N_17639,N_16539);
or U19309 (N_19309,N_17514,N_16236);
nor U19310 (N_19310,N_16996,N_17208);
nand U19311 (N_19311,N_17445,N_16995);
xnor U19312 (N_19312,N_16404,N_16314);
and U19313 (N_19313,N_16663,N_16994);
nor U19314 (N_19314,N_17665,N_16464);
nor U19315 (N_19315,N_16183,N_17103);
or U19316 (N_19316,N_17106,N_16918);
or U19317 (N_19317,N_17215,N_16394);
xnor U19318 (N_19318,N_17216,N_16327);
nand U19319 (N_19319,N_17434,N_16811);
nand U19320 (N_19320,N_17692,N_16763);
xor U19321 (N_19321,N_16181,N_16133);
xor U19322 (N_19322,N_17182,N_16983);
and U19323 (N_19323,N_17135,N_16176);
nand U19324 (N_19324,N_16953,N_17776);
nor U19325 (N_19325,N_16656,N_16922);
or U19326 (N_19326,N_17712,N_16452);
and U19327 (N_19327,N_17355,N_17059);
and U19328 (N_19328,N_16441,N_17452);
nor U19329 (N_19329,N_17689,N_16673);
nor U19330 (N_19330,N_17661,N_17212);
nand U19331 (N_19331,N_17429,N_16794);
or U19332 (N_19332,N_17339,N_16262);
xor U19333 (N_19333,N_16010,N_17921);
nand U19334 (N_19334,N_16464,N_17689);
nand U19335 (N_19335,N_16155,N_17131);
or U19336 (N_19336,N_16192,N_17059);
xor U19337 (N_19337,N_17147,N_17962);
or U19338 (N_19338,N_16659,N_17669);
xor U19339 (N_19339,N_17449,N_17688);
or U19340 (N_19340,N_17904,N_17204);
and U19341 (N_19341,N_17543,N_17572);
nor U19342 (N_19342,N_17296,N_17878);
or U19343 (N_19343,N_17558,N_16318);
nor U19344 (N_19344,N_16394,N_17491);
nor U19345 (N_19345,N_17922,N_17781);
xor U19346 (N_19346,N_17059,N_16856);
xor U19347 (N_19347,N_16118,N_16890);
xor U19348 (N_19348,N_17769,N_16814);
or U19349 (N_19349,N_17136,N_17882);
xnor U19350 (N_19350,N_16140,N_16173);
nand U19351 (N_19351,N_16268,N_16527);
nor U19352 (N_19352,N_17451,N_16160);
nand U19353 (N_19353,N_17965,N_16688);
xnor U19354 (N_19354,N_17095,N_17926);
or U19355 (N_19355,N_16281,N_17481);
and U19356 (N_19356,N_17683,N_17886);
nor U19357 (N_19357,N_16096,N_17665);
xnor U19358 (N_19358,N_16775,N_16595);
and U19359 (N_19359,N_16838,N_17641);
xnor U19360 (N_19360,N_16596,N_16906);
or U19361 (N_19361,N_17569,N_16980);
nand U19362 (N_19362,N_16332,N_17757);
nor U19363 (N_19363,N_16035,N_16176);
and U19364 (N_19364,N_17232,N_16599);
or U19365 (N_19365,N_17022,N_17815);
xor U19366 (N_19366,N_17188,N_16816);
xnor U19367 (N_19367,N_16068,N_16584);
nor U19368 (N_19368,N_16977,N_16901);
nand U19369 (N_19369,N_16754,N_16466);
or U19370 (N_19370,N_17548,N_16535);
nand U19371 (N_19371,N_17852,N_16508);
nand U19372 (N_19372,N_17663,N_16562);
nand U19373 (N_19373,N_17486,N_17864);
xnor U19374 (N_19374,N_16026,N_16626);
xor U19375 (N_19375,N_17624,N_16049);
and U19376 (N_19376,N_16690,N_16485);
nand U19377 (N_19377,N_16800,N_16445);
xnor U19378 (N_19378,N_16589,N_17848);
nand U19379 (N_19379,N_16523,N_16923);
nand U19380 (N_19380,N_17844,N_16075);
xnor U19381 (N_19381,N_16836,N_17293);
nand U19382 (N_19382,N_16894,N_17982);
xor U19383 (N_19383,N_17301,N_17771);
xnor U19384 (N_19384,N_17882,N_16979);
or U19385 (N_19385,N_16052,N_17669);
nor U19386 (N_19386,N_16998,N_17285);
nand U19387 (N_19387,N_16234,N_17765);
nand U19388 (N_19388,N_17077,N_16921);
xnor U19389 (N_19389,N_16122,N_17915);
xnor U19390 (N_19390,N_16972,N_17323);
nand U19391 (N_19391,N_17077,N_17011);
nand U19392 (N_19392,N_16321,N_17314);
xor U19393 (N_19393,N_16714,N_16460);
xor U19394 (N_19394,N_16053,N_16123);
and U19395 (N_19395,N_17471,N_17549);
nor U19396 (N_19396,N_17053,N_16770);
and U19397 (N_19397,N_16069,N_17686);
and U19398 (N_19398,N_16286,N_17495);
nand U19399 (N_19399,N_16845,N_17486);
nor U19400 (N_19400,N_17784,N_17009);
nor U19401 (N_19401,N_17613,N_16394);
and U19402 (N_19402,N_17078,N_17312);
xnor U19403 (N_19403,N_17566,N_17880);
nand U19404 (N_19404,N_17096,N_17623);
and U19405 (N_19405,N_17892,N_17093);
xnor U19406 (N_19406,N_16717,N_16027);
or U19407 (N_19407,N_16985,N_16878);
nand U19408 (N_19408,N_17538,N_16593);
or U19409 (N_19409,N_16545,N_16048);
and U19410 (N_19410,N_16860,N_17642);
nor U19411 (N_19411,N_17275,N_17278);
and U19412 (N_19412,N_17760,N_17337);
nor U19413 (N_19413,N_17453,N_16691);
xnor U19414 (N_19414,N_16631,N_16963);
nor U19415 (N_19415,N_17300,N_16315);
nand U19416 (N_19416,N_17654,N_17443);
nand U19417 (N_19417,N_16885,N_16829);
xor U19418 (N_19418,N_16462,N_17380);
nand U19419 (N_19419,N_17628,N_16546);
and U19420 (N_19420,N_16108,N_16863);
nand U19421 (N_19421,N_16949,N_17199);
xnor U19422 (N_19422,N_17392,N_17968);
nor U19423 (N_19423,N_17552,N_16674);
or U19424 (N_19424,N_16116,N_16180);
or U19425 (N_19425,N_17785,N_17780);
xnor U19426 (N_19426,N_17953,N_17940);
and U19427 (N_19427,N_17214,N_17272);
nor U19428 (N_19428,N_17149,N_16321);
and U19429 (N_19429,N_17195,N_16049);
and U19430 (N_19430,N_17273,N_17379);
xor U19431 (N_19431,N_17958,N_17716);
nand U19432 (N_19432,N_17407,N_16047);
and U19433 (N_19433,N_17704,N_16628);
nand U19434 (N_19434,N_17815,N_16415);
or U19435 (N_19435,N_16360,N_16037);
nor U19436 (N_19436,N_17136,N_16578);
and U19437 (N_19437,N_17099,N_17026);
and U19438 (N_19438,N_16038,N_16431);
or U19439 (N_19439,N_17221,N_16542);
xor U19440 (N_19440,N_16273,N_16114);
and U19441 (N_19441,N_16649,N_17969);
and U19442 (N_19442,N_16977,N_17452);
nor U19443 (N_19443,N_16137,N_16550);
nand U19444 (N_19444,N_16939,N_17462);
nor U19445 (N_19445,N_17704,N_17239);
nand U19446 (N_19446,N_17744,N_17305);
xor U19447 (N_19447,N_17296,N_16930);
or U19448 (N_19448,N_16316,N_16474);
or U19449 (N_19449,N_16306,N_17802);
and U19450 (N_19450,N_17734,N_17671);
xnor U19451 (N_19451,N_16274,N_17763);
nor U19452 (N_19452,N_16162,N_16960);
nor U19453 (N_19453,N_16213,N_16664);
nand U19454 (N_19454,N_16443,N_17375);
nand U19455 (N_19455,N_17702,N_16035);
nand U19456 (N_19456,N_17254,N_16944);
nand U19457 (N_19457,N_17399,N_17422);
xnor U19458 (N_19458,N_16917,N_17563);
or U19459 (N_19459,N_16049,N_16105);
xnor U19460 (N_19460,N_17890,N_17820);
and U19461 (N_19461,N_17624,N_16285);
or U19462 (N_19462,N_16451,N_17617);
xor U19463 (N_19463,N_17008,N_17559);
and U19464 (N_19464,N_17990,N_16083);
nand U19465 (N_19465,N_17425,N_16140);
nor U19466 (N_19466,N_17264,N_16796);
or U19467 (N_19467,N_17559,N_16538);
nor U19468 (N_19468,N_17417,N_17291);
and U19469 (N_19469,N_16986,N_16240);
nor U19470 (N_19470,N_17566,N_16821);
nor U19471 (N_19471,N_17317,N_17087);
or U19472 (N_19472,N_16872,N_17785);
nor U19473 (N_19473,N_16401,N_16398);
and U19474 (N_19474,N_16203,N_17650);
and U19475 (N_19475,N_16751,N_17452);
nor U19476 (N_19476,N_16793,N_17005);
and U19477 (N_19477,N_17898,N_16982);
nand U19478 (N_19478,N_17526,N_16468);
or U19479 (N_19479,N_17994,N_16506);
and U19480 (N_19480,N_17544,N_16110);
nand U19481 (N_19481,N_16162,N_16531);
nand U19482 (N_19482,N_16358,N_17386);
nor U19483 (N_19483,N_16146,N_17204);
and U19484 (N_19484,N_17284,N_17614);
xnor U19485 (N_19485,N_17614,N_17871);
nor U19486 (N_19486,N_17509,N_17213);
and U19487 (N_19487,N_17939,N_16278);
or U19488 (N_19488,N_17241,N_16875);
or U19489 (N_19489,N_16275,N_17047);
or U19490 (N_19490,N_16188,N_17819);
and U19491 (N_19491,N_16370,N_17223);
and U19492 (N_19492,N_16546,N_16578);
and U19493 (N_19493,N_17188,N_16356);
xnor U19494 (N_19494,N_17193,N_17023);
nor U19495 (N_19495,N_16920,N_17743);
nand U19496 (N_19496,N_16296,N_16337);
nor U19497 (N_19497,N_16106,N_16974);
xor U19498 (N_19498,N_17855,N_16508);
nand U19499 (N_19499,N_16094,N_17021);
nand U19500 (N_19500,N_17597,N_17668);
xnor U19501 (N_19501,N_16438,N_17662);
nand U19502 (N_19502,N_17609,N_16845);
or U19503 (N_19503,N_16555,N_17150);
or U19504 (N_19504,N_16686,N_17638);
and U19505 (N_19505,N_17441,N_17727);
or U19506 (N_19506,N_17407,N_17169);
or U19507 (N_19507,N_17745,N_17553);
or U19508 (N_19508,N_16374,N_16587);
or U19509 (N_19509,N_17427,N_17094);
and U19510 (N_19510,N_17408,N_16997);
and U19511 (N_19511,N_16760,N_17211);
or U19512 (N_19512,N_17794,N_16942);
or U19513 (N_19513,N_17252,N_16046);
xnor U19514 (N_19514,N_16705,N_16365);
xnor U19515 (N_19515,N_17007,N_17842);
nor U19516 (N_19516,N_16057,N_17002);
nor U19517 (N_19517,N_16011,N_16905);
and U19518 (N_19518,N_16405,N_17194);
nor U19519 (N_19519,N_16676,N_17380);
and U19520 (N_19520,N_16325,N_16604);
or U19521 (N_19521,N_17337,N_16012);
xnor U19522 (N_19522,N_17593,N_17113);
nor U19523 (N_19523,N_17559,N_17776);
nand U19524 (N_19524,N_17652,N_16225);
or U19525 (N_19525,N_16033,N_17037);
and U19526 (N_19526,N_16142,N_17952);
nor U19527 (N_19527,N_16566,N_16018);
and U19528 (N_19528,N_17003,N_16884);
xnor U19529 (N_19529,N_16843,N_16654);
or U19530 (N_19530,N_16740,N_17516);
nor U19531 (N_19531,N_17146,N_17887);
and U19532 (N_19532,N_16319,N_17254);
and U19533 (N_19533,N_16901,N_17445);
xor U19534 (N_19534,N_16693,N_17083);
nand U19535 (N_19535,N_16642,N_17409);
nor U19536 (N_19536,N_17805,N_16486);
nor U19537 (N_19537,N_17281,N_17378);
nand U19538 (N_19538,N_17613,N_16105);
or U19539 (N_19539,N_17562,N_16954);
or U19540 (N_19540,N_17014,N_17538);
nand U19541 (N_19541,N_17437,N_17545);
and U19542 (N_19542,N_16345,N_16728);
nand U19543 (N_19543,N_17613,N_16883);
xnor U19544 (N_19544,N_17031,N_16230);
or U19545 (N_19545,N_16719,N_17486);
and U19546 (N_19546,N_17658,N_17905);
or U19547 (N_19547,N_16774,N_17162);
and U19548 (N_19548,N_17707,N_17563);
xnor U19549 (N_19549,N_17975,N_16564);
or U19550 (N_19550,N_16835,N_16255);
and U19551 (N_19551,N_16291,N_17699);
xor U19552 (N_19552,N_17904,N_16357);
xor U19553 (N_19553,N_17800,N_17730);
nand U19554 (N_19554,N_17408,N_16503);
xnor U19555 (N_19555,N_16043,N_16976);
and U19556 (N_19556,N_17437,N_16975);
xnor U19557 (N_19557,N_16121,N_16236);
xnor U19558 (N_19558,N_16450,N_16561);
nand U19559 (N_19559,N_16401,N_16052);
xnor U19560 (N_19560,N_16199,N_16272);
nor U19561 (N_19561,N_16348,N_17633);
or U19562 (N_19562,N_17988,N_16742);
and U19563 (N_19563,N_16341,N_17831);
xnor U19564 (N_19564,N_16668,N_17229);
and U19565 (N_19565,N_17951,N_17733);
or U19566 (N_19566,N_16836,N_16480);
xnor U19567 (N_19567,N_16515,N_16675);
nor U19568 (N_19568,N_17240,N_17347);
or U19569 (N_19569,N_17680,N_16502);
nand U19570 (N_19570,N_16260,N_16134);
nand U19571 (N_19571,N_16944,N_16140);
nor U19572 (N_19572,N_16425,N_16885);
and U19573 (N_19573,N_17048,N_17538);
nor U19574 (N_19574,N_17273,N_17658);
xor U19575 (N_19575,N_16324,N_16083);
nor U19576 (N_19576,N_17865,N_17764);
and U19577 (N_19577,N_17112,N_16414);
nor U19578 (N_19578,N_16898,N_16299);
nor U19579 (N_19579,N_17484,N_17175);
nand U19580 (N_19580,N_16256,N_16617);
nand U19581 (N_19581,N_16509,N_17532);
nand U19582 (N_19582,N_16428,N_17255);
and U19583 (N_19583,N_16936,N_17975);
and U19584 (N_19584,N_17215,N_17872);
nand U19585 (N_19585,N_17002,N_17457);
xnor U19586 (N_19586,N_17248,N_16792);
and U19587 (N_19587,N_17767,N_17500);
and U19588 (N_19588,N_17519,N_16632);
and U19589 (N_19589,N_16762,N_17799);
xnor U19590 (N_19590,N_16014,N_16688);
nand U19591 (N_19591,N_16888,N_17483);
xnor U19592 (N_19592,N_17079,N_16590);
nor U19593 (N_19593,N_17288,N_16729);
or U19594 (N_19594,N_17782,N_17695);
or U19595 (N_19595,N_16950,N_17420);
or U19596 (N_19596,N_17501,N_17859);
nor U19597 (N_19597,N_16426,N_16807);
or U19598 (N_19598,N_16124,N_16458);
nor U19599 (N_19599,N_17251,N_17687);
and U19600 (N_19600,N_17455,N_16066);
nand U19601 (N_19601,N_16210,N_16499);
xnor U19602 (N_19602,N_17104,N_16510);
nand U19603 (N_19603,N_17936,N_16963);
nand U19604 (N_19604,N_17090,N_17212);
or U19605 (N_19605,N_16516,N_16563);
or U19606 (N_19606,N_16062,N_16548);
or U19607 (N_19607,N_16158,N_17651);
or U19608 (N_19608,N_17973,N_16955);
nor U19609 (N_19609,N_17724,N_16964);
xnor U19610 (N_19610,N_17481,N_16802);
xor U19611 (N_19611,N_16413,N_17865);
nor U19612 (N_19612,N_17351,N_16259);
xnor U19613 (N_19613,N_17381,N_17034);
nand U19614 (N_19614,N_17006,N_16975);
nor U19615 (N_19615,N_16113,N_17638);
nor U19616 (N_19616,N_17192,N_16104);
nand U19617 (N_19617,N_17989,N_17680);
xnor U19618 (N_19618,N_17964,N_16681);
nand U19619 (N_19619,N_17886,N_17127);
or U19620 (N_19620,N_17593,N_17719);
xnor U19621 (N_19621,N_16816,N_17084);
nor U19622 (N_19622,N_16383,N_17053);
nor U19623 (N_19623,N_17760,N_17016);
nor U19624 (N_19624,N_17186,N_16072);
or U19625 (N_19625,N_16019,N_16858);
nand U19626 (N_19626,N_17052,N_16279);
xor U19627 (N_19627,N_16256,N_16692);
nand U19628 (N_19628,N_16392,N_16795);
xnor U19629 (N_19629,N_17835,N_16226);
xor U19630 (N_19630,N_16128,N_17598);
xor U19631 (N_19631,N_17482,N_16029);
or U19632 (N_19632,N_16476,N_17539);
and U19633 (N_19633,N_16618,N_17370);
or U19634 (N_19634,N_17858,N_17135);
xor U19635 (N_19635,N_17992,N_16908);
nand U19636 (N_19636,N_17156,N_17849);
or U19637 (N_19637,N_16057,N_17887);
nor U19638 (N_19638,N_16001,N_17867);
and U19639 (N_19639,N_17762,N_17693);
nor U19640 (N_19640,N_17804,N_16875);
nand U19641 (N_19641,N_16278,N_16843);
nand U19642 (N_19642,N_16549,N_16068);
xor U19643 (N_19643,N_17199,N_17391);
and U19644 (N_19644,N_16253,N_16459);
or U19645 (N_19645,N_17574,N_16171);
nand U19646 (N_19646,N_17124,N_16011);
nor U19647 (N_19647,N_16841,N_16050);
and U19648 (N_19648,N_17348,N_16251);
nand U19649 (N_19649,N_16872,N_17029);
nand U19650 (N_19650,N_17214,N_16472);
nor U19651 (N_19651,N_17871,N_16364);
xor U19652 (N_19652,N_16637,N_17659);
xor U19653 (N_19653,N_17240,N_16270);
nand U19654 (N_19654,N_17456,N_16858);
nor U19655 (N_19655,N_16739,N_16720);
or U19656 (N_19656,N_16756,N_17775);
and U19657 (N_19657,N_16360,N_16500);
or U19658 (N_19658,N_17631,N_16776);
nor U19659 (N_19659,N_16913,N_16209);
and U19660 (N_19660,N_16761,N_16794);
or U19661 (N_19661,N_17708,N_17682);
and U19662 (N_19662,N_16944,N_16736);
xor U19663 (N_19663,N_17271,N_16415);
nand U19664 (N_19664,N_16394,N_16952);
or U19665 (N_19665,N_16613,N_17869);
or U19666 (N_19666,N_16953,N_16193);
xor U19667 (N_19667,N_17168,N_17042);
xnor U19668 (N_19668,N_16211,N_16956);
and U19669 (N_19669,N_16115,N_17895);
and U19670 (N_19670,N_17819,N_17496);
and U19671 (N_19671,N_17686,N_17129);
nand U19672 (N_19672,N_17540,N_17175);
or U19673 (N_19673,N_16210,N_17710);
nor U19674 (N_19674,N_17815,N_16684);
nor U19675 (N_19675,N_16686,N_17624);
nand U19676 (N_19676,N_16836,N_16865);
xnor U19677 (N_19677,N_16462,N_16527);
xor U19678 (N_19678,N_16857,N_16934);
nand U19679 (N_19679,N_17608,N_16495);
nand U19680 (N_19680,N_16769,N_16792);
nand U19681 (N_19681,N_17523,N_17632);
xor U19682 (N_19682,N_16960,N_17106);
or U19683 (N_19683,N_16311,N_17214);
nand U19684 (N_19684,N_17147,N_16969);
nor U19685 (N_19685,N_17332,N_16385);
and U19686 (N_19686,N_17582,N_17752);
and U19687 (N_19687,N_16949,N_16187);
xnor U19688 (N_19688,N_16245,N_16421);
xnor U19689 (N_19689,N_17932,N_17805);
and U19690 (N_19690,N_17949,N_16667);
or U19691 (N_19691,N_16559,N_16257);
and U19692 (N_19692,N_16976,N_16851);
nand U19693 (N_19693,N_16225,N_17383);
nand U19694 (N_19694,N_17711,N_17733);
nand U19695 (N_19695,N_16149,N_16813);
and U19696 (N_19696,N_16047,N_16296);
nor U19697 (N_19697,N_16672,N_16009);
xor U19698 (N_19698,N_16653,N_17588);
and U19699 (N_19699,N_17113,N_17426);
xnor U19700 (N_19700,N_16597,N_16897);
nand U19701 (N_19701,N_16936,N_17040);
nand U19702 (N_19702,N_16499,N_16215);
nor U19703 (N_19703,N_16704,N_17676);
and U19704 (N_19704,N_17446,N_16286);
and U19705 (N_19705,N_17633,N_16556);
nand U19706 (N_19706,N_17052,N_16368);
nand U19707 (N_19707,N_16764,N_17987);
xor U19708 (N_19708,N_17046,N_16966);
nand U19709 (N_19709,N_17934,N_17271);
or U19710 (N_19710,N_17243,N_16176);
nand U19711 (N_19711,N_16676,N_16175);
nor U19712 (N_19712,N_17033,N_16549);
or U19713 (N_19713,N_16214,N_16997);
nand U19714 (N_19714,N_17912,N_17235);
xor U19715 (N_19715,N_17260,N_17319);
nand U19716 (N_19716,N_17973,N_17088);
or U19717 (N_19717,N_16481,N_16196);
or U19718 (N_19718,N_17959,N_16697);
nand U19719 (N_19719,N_17865,N_16684);
xnor U19720 (N_19720,N_17965,N_17836);
xnor U19721 (N_19721,N_16781,N_17021);
and U19722 (N_19722,N_17824,N_17008);
nand U19723 (N_19723,N_17902,N_16359);
nand U19724 (N_19724,N_17075,N_16573);
and U19725 (N_19725,N_16307,N_16884);
and U19726 (N_19726,N_17136,N_17180);
nand U19727 (N_19727,N_17799,N_16413);
and U19728 (N_19728,N_16574,N_16756);
or U19729 (N_19729,N_17779,N_16158);
nor U19730 (N_19730,N_16567,N_16932);
nor U19731 (N_19731,N_17536,N_17023);
or U19732 (N_19732,N_17266,N_16695);
xnor U19733 (N_19733,N_17235,N_16976);
xor U19734 (N_19734,N_17944,N_16901);
nor U19735 (N_19735,N_17023,N_16047);
xor U19736 (N_19736,N_17352,N_17546);
xnor U19737 (N_19737,N_17069,N_17148);
nand U19738 (N_19738,N_17655,N_16247);
nor U19739 (N_19739,N_17562,N_16348);
and U19740 (N_19740,N_16095,N_16480);
nor U19741 (N_19741,N_16173,N_16981);
nor U19742 (N_19742,N_17950,N_16339);
xnor U19743 (N_19743,N_17713,N_17575);
xor U19744 (N_19744,N_16735,N_17651);
nand U19745 (N_19745,N_17496,N_17934);
or U19746 (N_19746,N_17645,N_16873);
or U19747 (N_19747,N_17090,N_16081);
xor U19748 (N_19748,N_17279,N_16051);
nor U19749 (N_19749,N_16926,N_17855);
xor U19750 (N_19750,N_16428,N_16888);
nand U19751 (N_19751,N_16992,N_17679);
nor U19752 (N_19752,N_16913,N_17710);
and U19753 (N_19753,N_17378,N_16919);
and U19754 (N_19754,N_16157,N_16678);
xnor U19755 (N_19755,N_16673,N_16214);
and U19756 (N_19756,N_16519,N_17845);
and U19757 (N_19757,N_16955,N_17026);
and U19758 (N_19758,N_16654,N_16437);
nor U19759 (N_19759,N_16899,N_17332);
nand U19760 (N_19760,N_17623,N_16354);
nand U19761 (N_19761,N_16205,N_17861);
xnor U19762 (N_19762,N_16321,N_17218);
xor U19763 (N_19763,N_17751,N_16663);
and U19764 (N_19764,N_17022,N_16898);
xnor U19765 (N_19765,N_16189,N_16074);
xnor U19766 (N_19766,N_17947,N_17096);
or U19767 (N_19767,N_16914,N_17683);
nor U19768 (N_19768,N_17568,N_16421);
and U19769 (N_19769,N_16300,N_17756);
xor U19770 (N_19770,N_17127,N_17456);
and U19771 (N_19771,N_17876,N_16124);
or U19772 (N_19772,N_17653,N_17834);
and U19773 (N_19773,N_17122,N_16446);
and U19774 (N_19774,N_16269,N_16942);
nand U19775 (N_19775,N_16482,N_16648);
nand U19776 (N_19776,N_17349,N_16000);
and U19777 (N_19777,N_17074,N_17435);
xnor U19778 (N_19778,N_17034,N_17316);
or U19779 (N_19779,N_16613,N_16737);
xor U19780 (N_19780,N_17046,N_17181);
xor U19781 (N_19781,N_17140,N_17666);
nand U19782 (N_19782,N_16530,N_17046);
nor U19783 (N_19783,N_16386,N_16533);
and U19784 (N_19784,N_16048,N_17985);
and U19785 (N_19785,N_17400,N_16558);
and U19786 (N_19786,N_16878,N_16125);
and U19787 (N_19787,N_17223,N_16202);
or U19788 (N_19788,N_17257,N_16786);
xnor U19789 (N_19789,N_16160,N_16268);
xor U19790 (N_19790,N_17205,N_17701);
xor U19791 (N_19791,N_17418,N_17613);
or U19792 (N_19792,N_17315,N_17247);
or U19793 (N_19793,N_17907,N_17496);
and U19794 (N_19794,N_16881,N_16516);
nand U19795 (N_19795,N_17101,N_17528);
nor U19796 (N_19796,N_17353,N_16529);
xnor U19797 (N_19797,N_17335,N_17404);
nand U19798 (N_19798,N_16939,N_16709);
nor U19799 (N_19799,N_17557,N_16611);
xor U19800 (N_19800,N_16814,N_17751);
and U19801 (N_19801,N_16638,N_17289);
nor U19802 (N_19802,N_16890,N_16069);
and U19803 (N_19803,N_17139,N_16293);
nor U19804 (N_19804,N_17787,N_16647);
or U19805 (N_19805,N_17576,N_17660);
and U19806 (N_19806,N_16471,N_16188);
or U19807 (N_19807,N_17373,N_17424);
nand U19808 (N_19808,N_17130,N_16367);
nor U19809 (N_19809,N_16727,N_17579);
nor U19810 (N_19810,N_17109,N_17655);
xor U19811 (N_19811,N_16345,N_16313);
and U19812 (N_19812,N_16760,N_16064);
xnor U19813 (N_19813,N_16174,N_16808);
nand U19814 (N_19814,N_17841,N_17566);
nand U19815 (N_19815,N_17602,N_17523);
nand U19816 (N_19816,N_16499,N_16343);
and U19817 (N_19817,N_17927,N_16324);
xor U19818 (N_19818,N_17170,N_17343);
xnor U19819 (N_19819,N_17573,N_16591);
and U19820 (N_19820,N_17771,N_16625);
nor U19821 (N_19821,N_17431,N_17506);
xor U19822 (N_19822,N_16506,N_17141);
or U19823 (N_19823,N_16382,N_17869);
xor U19824 (N_19824,N_16680,N_17349);
or U19825 (N_19825,N_17988,N_17319);
xor U19826 (N_19826,N_17745,N_17455);
nand U19827 (N_19827,N_17151,N_16671);
and U19828 (N_19828,N_17788,N_16179);
and U19829 (N_19829,N_17421,N_16887);
nor U19830 (N_19830,N_17904,N_17020);
nand U19831 (N_19831,N_17870,N_16581);
nor U19832 (N_19832,N_16053,N_17768);
nand U19833 (N_19833,N_17618,N_16916);
nand U19834 (N_19834,N_17395,N_16946);
nand U19835 (N_19835,N_17601,N_16049);
nand U19836 (N_19836,N_16947,N_17194);
nand U19837 (N_19837,N_16426,N_17608);
xor U19838 (N_19838,N_17036,N_16521);
nor U19839 (N_19839,N_17213,N_16748);
nand U19840 (N_19840,N_16328,N_17998);
xor U19841 (N_19841,N_17228,N_17125);
nor U19842 (N_19842,N_16693,N_17574);
xor U19843 (N_19843,N_17137,N_17249);
or U19844 (N_19844,N_16623,N_17457);
xnor U19845 (N_19845,N_17092,N_17807);
nor U19846 (N_19846,N_17898,N_16412);
and U19847 (N_19847,N_17118,N_17008);
nand U19848 (N_19848,N_16910,N_17695);
nor U19849 (N_19849,N_17535,N_16691);
or U19850 (N_19850,N_17089,N_16138);
or U19851 (N_19851,N_16436,N_16140);
or U19852 (N_19852,N_16483,N_16409);
and U19853 (N_19853,N_17649,N_16159);
nor U19854 (N_19854,N_17408,N_17115);
nor U19855 (N_19855,N_17771,N_16448);
nand U19856 (N_19856,N_17986,N_16711);
xor U19857 (N_19857,N_17531,N_16328);
and U19858 (N_19858,N_17686,N_17110);
and U19859 (N_19859,N_16039,N_17284);
nor U19860 (N_19860,N_16573,N_16207);
xor U19861 (N_19861,N_16033,N_17031);
or U19862 (N_19862,N_16360,N_17776);
nor U19863 (N_19863,N_17483,N_16287);
nand U19864 (N_19864,N_17532,N_16918);
nand U19865 (N_19865,N_16906,N_17105);
nor U19866 (N_19866,N_16334,N_17089);
and U19867 (N_19867,N_16785,N_16338);
and U19868 (N_19868,N_16481,N_17452);
or U19869 (N_19869,N_17926,N_17434);
or U19870 (N_19870,N_16703,N_16420);
or U19871 (N_19871,N_16015,N_17264);
nor U19872 (N_19872,N_17470,N_16195);
nand U19873 (N_19873,N_17662,N_16952);
and U19874 (N_19874,N_17726,N_17503);
nand U19875 (N_19875,N_16135,N_17854);
and U19876 (N_19876,N_16221,N_17498);
xor U19877 (N_19877,N_16311,N_16417);
and U19878 (N_19878,N_16175,N_16526);
and U19879 (N_19879,N_17036,N_16987);
xor U19880 (N_19880,N_17435,N_17126);
or U19881 (N_19881,N_17764,N_17128);
nor U19882 (N_19882,N_16188,N_17020);
or U19883 (N_19883,N_17026,N_16850);
or U19884 (N_19884,N_16079,N_16277);
or U19885 (N_19885,N_16132,N_16149);
and U19886 (N_19886,N_17295,N_16179);
or U19887 (N_19887,N_16855,N_17204);
nand U19888 (N_19888,N_16641,N_16848);
nor U19889 (N_19889,N_17608,N_16153);
nor U19890 (N_19890,N_17824,N_17538);
and U19891 (N_19891,N_16736,N_16838);
xor U19892 (N_19892,N_16762,N_16447);
and U19893 (N_19893,N_16365,N_16959);
nand U19894 (N_19894,N_17468,N_17767);
and U19895 (N_19895,N_17111,N_17872);
and U19896 (N_19896,N_17075,N_17743);
nand U19897 (N_19897,N_16966,N_16764);
xor U19898 (N_19898,N_16685,N_16857);
and U19899 (N_19899,N_16091,N_16241);
xnor U19900 (N_19900,N_17831,N_17952);
or U19901 (N_19901,N_16365,N_17529);
nand U19902 (N_19902,N_17581,N_17809);
and U19903 (N_19903,N_17679,N_17538);
xnor U19904 (N_19904,N_16555,N_17338);
and U19905 (N_19905,N_17371,N_16177);
nand U19906 (N_19906,N_16781,N_16590);
nand U19907 (N_19907,N_16667,N_16374);
nor U19908 (N_19908,N_16380,N_16045);
and U19909 (N_19909,N_17502,N_17226);
or U19910 (N_19910,N_16382,N_17445);
nor U19911 (N_19911,N_17619,N_16417);
and U19912 (N_19912,N_16719,N_16321);
nand U19913 (N_19913,N_16464,N_16390);
and U19914 (N_19914,N_16606,N_17642);
and U19915 (N_19915,N_16672,N_17352);
or U19916 (N_19916,N_16959,N_16323);
xor U19917 (N_19917,N_17141,N_17412);
nor U19918 (N_19918,N_16814,N_16870);
xnor U19919 (N_19919,N_17821,N_16979);
or U19920 (N_19920,N_16750,N_17629);
xnor U19921 (N_19921,N_16916,N_17025);
xnor U19922 (N_19922,N_17201,N_17806);
and U19923 (N_19923,N_16531,N_16544);
nand U19924 (N_19924,N_16704,N_16490);
nand U19925 (N_19925,N_16812,N_17345);
or U19926 (N_19926,N_17616,N_17567);
and U19927 (N_19927,N_16563,N_16682);
nor U19928 (N_19928,N_17850,N_16530);
nor U19929 (N_19929,N_17808,N_16477);
nor U19930 (N_19930,N_16777,N_17513);
nand U19931 (N_19931,N_17439,N_17243);
nand U19932 (N_19932,N_17295,N_16489);
nand U19933 (N_19933,N_17063,N_16629);
or U19934 (N_19934,N_16105,N_16976);
nor U19935 (N_19935,N_17849,N_17640);
nor U19936 (N_19936,N_17056,N_17441);
xnor U19937 (N_19937,N_16277,N_17454);
and U19938 (N_19938,N_16111,N_17935);
xor U19939 (N_19939,N_17969,N_16987);
nand U19940 (N_19940,N_17341,N_16721);
nor U19941 (N_19941,N_16950,N_16893);
nand U19942 (N_19942,N_17322,N_16939);
or U19943 (N_19943,N_16399,N_17553);
or U19944 (N_19944,N_17266,N_16631);
or U19945 (N_19945,N_16055,N_17255);
or U19946 (N_19946,N_17055,N_17574);
or U19947 (N_19947,N_17570,N_16760);
nor U19948 (N_19948,N_17702,N_16011);
nand U19949 (N_19949,N_17518,N_16499);
nand U19950 (N_19950,N_16079,N_17780);
or U19951 (N_19951,N_17841,N_17130);
nand U19952 (N_19952,N_17458,N_16618);
nor U19953 (N_19953,N_16243,N_16460);
or U19954 (N_19954,N_17613,N_16866);
and U19955 (N_19955,N_17808,N_17301);
and U19956 (N_19956,N_16088,N_17359);
nor U19957 (N_19957,N_16996,N_17618);
or U19958 (N_19958,N_16661,N_16009);
nand U19959 (N_19959,N_16472,N_17609);
nor U19960 (N_19960,N_17691,N_16384);
or U19961 (N_19961,N_17684,N_17919);
nand U19962 (N_19962,N_16484,N_16042);
or U19963 (N_19963,N_17747,N_16202);
xor U19964 (N_19964,N_16661,N_16461);
nor U19965 (N_19965,N_16316,N_17584);
nor U19966 (N_19966,N_16785,N_17539);
xnor U19967 (N_19967,N_16675,N_17356);
and U19968 (N_19968,N_17895,N_16947);
or U19969 (N_19969,N_16017,N_16783);
nor U19970 (N_19970,N_16451,N_16771);
nand U19971 (N_19971,N_16644,N_17039);
or U19972 (N_19972,N_16111,N_17585);
and U19973 (N_19973,N_17187,N_17435);
and U19974 (N_19974,N_16967,N_17841);
xnor U19975 (N_19975,N_16293,N_17832);
or U19976 (N_19976,N_16927,N_16622);
nor U19977 (N_19977,N_17098,N_16763);
nor U19978 (N_19978,N_16751,N_16265);
and U19979 (N_19979,N_17961,N_17681);
or U19980 (N_19980,N_16481,N_17290);
and U19981 (N_19981,N_17967,N_17717);
nor U19982 (N_19982,N_17193,N_16621);
xnor U19983 (N_19983,N_16521,N_17753);
xnor U19984 (N_19984,N_17581,N_17102);
nor U19985 (N_19985,N_16064,N_17269);
and U19986 (N_19986,N_17636,N_16675);
or U19987 (N_19987,N_17582,N_16115);
nor U19988 (N_19988,N_16560,N_16923);
xnor U19989 (N_19989,N_17147,N_16012);
or U19990 (N_19990,N_16834,N_16473);
and U19991 (N_19991,N_17775,N_16070);
xor U19992 (N_19992,N_17023,N_17587);
nor U19993 (N_19993,N_16766,N_17387);
or U19994 (N_19994,N_16512,N_16875);
nor U19995 (N_19995,N_17573,N_16994);
xnor U19996 (N_19996,N_16158,N_16577);
nand U19997 (N_19997,N_16952,N_17919);
nand U19998 (N_19998,N_17270,N_16573);
nor U19999 (N_19999,N_17475,N_17266);
and U20000 (N_20000,N_18000,N_19825);
nor U20001 (N_20001,N_19473,N_19816);
nand U20002 (N_20002,N_18113,N_19516);
xor U20003 (N_20003,N_19806,N_19480);
nor U20004 (N_20004,N_19501,N_19441);
and U20005 (N_20005,N_18177,N_19222);
and U20006 (N_20006,N_18183,N_18696);
xor U20007 (N_20007,N_18964,N_19803);
or U20008 (N_20008,N_18044,N_18294);
or U20009 (N_20009,N_18943,N_19013);
xnor U20010 (N_20010,N_19419,N_18078);
xor U20011 (N_20011,N_18868,N_19517);
xor U20012 (N_20012,N_18881,N_19583);
xor U20013 (N_20013,N_18494,N_19664);
nor U20014 (N_20014,N_19867,N_18380);
nor U20015 (N_20015,N_18255,N_18398);
nor U20016 (N_20016,N_18709,N_19336);
xnor U20017 (N_20017,N_18598,N_18094);
nand U20018 (N_20018,N_19903,N_19839);
xnor U20019 (N_20019,N_18188,N_18762);
or U20020 (N_20020,N_19621,N_18351);
or U20021 (N_20021,N_19955,N_19525);
or U20022 (N_20022,N_18182,N_19012);
xnor U20023 (N_20023,N_18370,N_19627);
xnor U20024 (N_20024,N_18835,N_18534);
xnor U20025 (N_20025,N_19310,N_19167);
and U20026 (N_20026,N_19145,N_19019);
and U20027 (N_20027,N_18458,N_19003);
nor U20028 (N_20028,N_19482,N_19027);
nor U20029 (N_20029,N_18514,N_19283);
and U20030 (N_20030,N_18116,N_19998);
nand U20031 (N_20031,N_19017,N_19103);
and U20032 (N_20032,N_19511,N_18129);
nand U20033 (N_20033,N_18437,N_18739);
or U20034 (N_20034,N_18864,N_19932);
or U20035 (N_20035,N_18218,N_19974);
xor U20036 (N_20036,N_18701,N_18633);
nand U20037 (N_20037,N_18411,N_19792);
or U20038 (N_20038,N_19580,N_18510);
and U20039 (N_20039,N_19552,N_19261);
or U20040 (N_20040,N_19328,N_18834);
nor U20041 (N_20041,N_19919,N_19457);
or U20042 (N_20042,N_19978,N_18635);
or U20043 (N_20043,N_18776,N_19692);
xnor U20044 (N_20044,N_19423,N_18065);
xnor U20045 (N_20045,N_18928,N_18756);
xor U20046 (N_20046,N_18721,N_19130);
or U20047 (N_20047,N_19929,N_19312);
nand U20048 (N_20048,N_18276,N_19892);
nand U20049 (N_20049,N_18793,N_19086);
nand U20050 (N_20050,N_19508,N_19970);
nor U20051 (N_20051,N_19590,N_19684);
nand U20052 (N_20052,N_19291,N_18006);
or U20053 (N_20053,N_19064,N_19185);
or U20054 (N_20054,N_18664,N_19871);
and U20055 (N_20055,N_18902,N_18335);
or U20056 (N_20056,N_19172,N_18528);
or U20057 (N_20057,N_19949,N_18125);
and U20058 (N_20058,N_19574,N_19556);
and U20059 (N_20059,N_19622,N_18053);
or U20060 (N_20060,N_18095,N_19895);
nor U20061 (N_20061,N_18471,N_18252);
nand U20062 (N_20062,N_18106,N_19139);
nor U20063 (N_20063,N_19957,N_18666);
and U20064 (N_20064,N_18700,N_19776);
nor U20065 (N_20065,N_18271,N_19496);
xor U20066 (N_20066,N_19104,N_18744);
and U20067 (N_20067,N_19408,N_19240);
or U20068 (N_20068,N_18777,N_18190);
nand U20069 (N_20069,N_19040,N_18518);
nor U20070 (N_20070,N_19376,N_19958);
nand U20071 (N_20071,N_18475,N_19676);
or U20072 (N_20072,N_19371,N_19306);
or U20073 (N_20073,N_18714,N_18054);
and U20074 (N_20074,N_19000,N_18509);
nor U20075 (N_20075,N_18445,N_19568);
nor U20076 (N_20076,N_18041,N_18191);
nand U20077 (N_20077,N_19221,N_19996);
or U20078 (N_20078,N_19450,N_18275);
and U20079 (N_20079,N_19727,N_19788);
or U20080 (N_20080,N_18782,N_19415);
nor U20081 (N_20081,N_19075,N_18951);
or U20082 (N_20082,N_18815,N_18526);
and U20083 (N_20083,N_19366,N_18886);
nor U20084 (N_20084,N_18122,N_18601);
and U20085 (N_20085,N_19883,N_19601);
nand U20086 (N_20086,N_19911,N_18512);
nor U20087 (N_20087,N_18331,N_19407);
or U20088 (N_20088,N_19180,N_18894);
or U20089 (N_20089,N_19295,N_19287);
and U20090 (N_20090,N_19330,N_19435);
xnor U20091 (N_20091,N_19131,N_19625);
nand U20092 (N_20092,N_18356,N_19960);
nand U20093 (N_20093,N_18677,N_18090);
nor U20094 (N_20094,N_18016,N_19355);
or U20095 (N_20095,N_19404,N_19173);
nand U20096 (N_20096,N_18806,N_19512);
xnor U20097 (N_20097,N_18640,N_18719);
nor U20098 (N_20098,N_19581,N_18871);
nand U20099 (N_20099,N_18628,N_19560);
nor U20100 (N_20100,N_19779,N_19117);
nor U20101 (N_20101,N_19785,N_18525);
xnor U20102 (N_20102,N_18329,N_18186);
and U20103 (N_20103,N_18641,N_18736);
or U20104 (N_20104,N_18308,N_18436);
nor U20105 (N_20105,N_18891,N_19662);
nor U20106 (N_20106,N_18315,N_19353);
xor U20107 (N_20107,N_19773,N_18836);
nor U20108 (N_20108,N_18724,N_18660);
nand U20109 (N_20109,N_19398,N_19445);
nand U20110 (N_20110,N_19963,N_18840);
nor U20111 (N_20111,N_19906,N_18029);
xor U20112 (N_20112,N_19712,N_18562);
and U20113 (N_20113,N_19186,N_18631);
nor U20114 (N_20114,N_18690,N_18564);
nand U20115 (N_20115,N_18126,N_19262);
xor U20116 (N_20116,N_18610,N_19354);
nand U20117 (N_20117,N_18219,N_18676);
nand U20118 (N_20118,N_19529,N_19832);
and U20119 (N_20119,N_18524,N_18193);
or U20120 (N_20120,N_19498,N_19746);
xor U20121 (N_20121,N_18319,N_18424);
nand U20122 (N_20122,N_19392,N_19577);
nor U20123 (N_20123,N_18361,N_18763);
and U20124 (N_20124,N_18180,N_19118);
or U20125 (N_20125,N_18703,N_18849);
xor U20126 (N_20126,N_18101,N_19576);
or U20127 (N_20127,N_18487,N_18797);
nor U20128 (N_20128,N_18832,N_18826);
nor U20129 (N_20129,N_19292,N_18649);
xor U20130 (N_20130,N_19536,N_19274);
nand U20131 (N_20131,N_18627,N_19096);
nand U20132 (N_20132,N_18327,N_18028);
or U20133 (N_20133,N_18164,N_18228);
xor U20134 (N_20134,N_19991,N_18673);
or U20135 (N_20135,N_19397,N_18301);
xnor U20136 (N_20136,N_18038,N_19005);
nor U20137 (N_20137,N_19087,N_19632);
xor U20138 (N_20138,N_18481,N_19053);
nor U20139 (N_20139,N_19715,N_19542);
nand U20140 (N_20140,N_18414,N_19899);
and U20141 (N_20141,N_18932,N_19977);
and U20142 (N_20142,N_18148,N_19205);
nand U20143 (N_20143,N_19546,N_19961);
nor U20144 (N_20144,N_18819,N_18742);
or U20145 (N_20145,N_18204,N_19432);
xor U20146 (N_20146,N_19777,N_18372);
xor U20147 (N_20147,N_18937,N_18992);
nor U20148 (N_20148,N_18754,N_18895);
or U20149 (N_20149,N_18682,N_19230);
and U20150 (N_20150,N_18866,N_19414);
xnor U20151 (N_20151,N_19456,N_19597);
nor U20152 (N_20152,N_18305,N_18792);
nand U20153 (N_20153,N_18155,N_18321);
nand U20154 (N_20154,N_19084,N_18720);
or U20155 (N_20155,N_19887,N_19774);
nand U20156 (N_20156,N_18973,N_18553);
or U20157 (N_20157,N_19035,N_18117);
and U20158 (N_20158,N_19361,N_19418);
nor U20159 (N_20159,N_18364,N_18083);
and U20160 (N_20160,N_19898,N_18726);
nor U20161 (N_20161,N_19078,N_19677);
nor U20162 (N_20162,N_18421,N_19613);
nand U20163 (N_20163,N_19935,N_18387);
or U20164 (N_20164,N_18366,N_18069);
xnor U20165 (N_20165,N_19391,N_18771);
nand U20166 (N_20166,N_18059,N_18358);
xnor U20167 (N_20167,N_19528,N_18908);
or U20168 (N_20168,N_18474,N_18824);
and U20169 (N_20169,N_19718,N_18194);
and U20170 (N_20170,N_19151,N_19672);
and U20171 (N_20171,N_18828,N_18657);
nand U20172 (N_20172,N_19997,N_18332);
and U20173 (N_20173,N_19413,N_19810);
nand U20174 (N_20174,N_18718,N_18310);
xor U20175 (N_20175,N_18379,N_19195);
xor U20176 (N_20176,N_18151,N_19559);
nor U20177 (N_20177,N_18061,N_19728);
nand U20178 (N_20178,N_19006,N_18163);
or U20179 (N_20179,N_19447,N_18844);
and U20180 (N_20180,N_19294,N_19537);
nor U20181 (N_20181,N_19438,N_18770);
and U20182 (N_20182,N_19604,N_19535);
nor U20183 (N_20183,N_18527,N_18442);
nor U20184 (N_20184,N_19679,N_19569);
nor U20185 (N_20185,N_18221,N_19610);
nor U20186 (N_20186,N_19538,N_19455);
and U20187 (N_20187,N_18179,N_19217);
xnor U20188 (N_20188,N_18533,N_18587);
nor U20189 (N_20189,N_19124,N_19818);
nor U20190 (N_20190,N_18324,N_19074);
or U20191 (N_20191,N_19479,N_18843);
nor U20192 (N_20192,N_18360,N_18449);
and U20193 (N_20193,N_19156,N_18854);
and U20194 (N_20194,N_19814,N_19859);
or U20195 (N_20195,N_19249,N_18723);
nand U20196 (N_20196,N_18795,N_19179);
nand U20197 (N_20197,N_18713,N_18946);
nand U20198 (N_20198,N_19634,N_18963);
or U20199 (N_20199,N_18671,N_18428);
nor U20200 (N_20200,N_19245,N_19638);
nor U20201 (N_20201,N_18076,N_18341);
nor U20202 (N_20202,N_18769,N_18224);
nand U20203 (N_20203,N_19506,N_19259);
xnor U20204 (N_20204,N_18202,N_18295);
and U20205 (N_20205,N_18270,N_18519);
xor U20206 (N_20206,N_19382,N_19646);
nand U20207 (N_20207,N_19409,N_18561);
xnor U20208 (N_20208,N_19979,N_18551);
and U20209 (N_20209,N_19572,N_18417);
and U20210 (N_20210,N_18800,N_18593);
and U20211 (N_20211,N_18130,N_18277);
nor U20212 (N_20212,N_19439,N_18779);
nand U20213 (N_20213,N_18263,N_18362);
xnor U20214 (N_20214,N_19640,N_19010);
nor U20215 (N_20215,N_18919,N_19891);
nor U20216 (N_20216,N_18269,N_18385);
or U20217 (N_20217,N_19140,N_19459);
xnor U20218 (N_20218,N_19550,N_19851);
nand U20219 (N_20219,N_19736,N_19263);
nand U20220 (N_20220,N_18609,N_19708);
xnor U20221 (N_20221,N_18565,N_19982);
xor U20222 (N_20222,N_18320,N_18419);
nand U20223 (N_20223,N_19034,N_19234);
nor U20224 (N_20224,N_19617,N_18037);
or U20225 (N_20225,N_19828,N_18950);
and U20226 (N_20226,N_18921,N_19789);
nor U20227 (N_20227,N_19349,N_19965);
and U20228 (N_20228,N_18234,N_18406);
xor U20229 (N_20229,N_18001,N_18773);
or U20230 (N_20230,N_18423,N_18585);
xnor U20231 (N_20231,N_18953,N_18761);
xnor U20232 (N_20232,N_19942,N_19214);
nor U20233 (N_20233,N_19723,N_19348);
xnor U20234 (N_20234,N_19062,N_18620);
xor U20235 (N_20235,N_18689,N_18418);
or U20236 (N_20236,N_19948,N_19691);
or U20237 (N_20237,N_19886,N_19155);
nor U20238 (N_20238,N_18281,N_19798);
nor U20239 (N_20239,N_18336,N_18260);
nor U20240 (N_20240,N_19322,N_18634);
nand U20241 (N_20241,N_19200,N_19813);
nand U20242 (N_20242,N_19316,N_19921);
or U20243 (N_20243,N_18933,N_19661);
nand U20244 (N_20244,N_18484,N_19068);
nand U20245 (N_20245,N_18317,N_18354);
or U20246 (N_20246,N_18903,N_19158);
or U20247 (N_20247,N_18994,N_19555);
xor U20248 (N_20248,N_18489,N_19393);
xor U20249 (N_20249,N_19260,N_19476);
nor U20250 (N_20250,N_18692,N_18887);
xnor U20251 (N_20251,N_18209,N_19870);
nor U20252 (N_20252,N_18486,N_19527);
nand U20253 (N_20253,N_18532,N_19338);
or U20254 (N_20254,N_19305,N_18780);
nand U20255 (N_20255,N_18019,N_19620);
nand U20256 (N_20256,N_19319,N_19428);
xor U20257 (N_20257,N_18743,N_19277);
xor U20258 (N_20258,N_19069,N_19317);
xnor U20259 (N_20259,N_18367,N_19043);
and U20260 (N_20260,N_18796,N_19218);
and U20261 (N_20261,N_19499,N_18496);
nor U20262 (N_20262,N_19734,N_19253);
or U20263 (N_20263,N_19163,N_19153);
nor U20264 (N_20264,N_19300,N_18592);
nand U20265 (N_20265,N_18904,N_19220);
or U20266 (N_20266,N_19890,N_19085);
or U20267 (N_20267,N_19372,N_19593);
xnor U20268 (N_20268,N_18923,N_19654);
and U20269 (N_20269,N_18373,N_18146);
xor U20270 (N_20270,N_18922,N_19280);
nand U20271 (N_20271,N_19227,N_19964);
xor U20272 (N_20272,N_19804,N_18389);
and U20273 (N_20273,N_19737,N_19036);
or U20274 (N_20274,N_19095,N_19369);
nand U20275 (N_20275,N_18307,N_18622);
nor U20276 (N_20276,N_19380,N_19464);
nor U20277 (N_20277,N_18216,N_18996);
nand U20278 (N_20278,N_18064,N_19207);
nand U20279 (N_20279,N_19713,N_18642);
xnor U20280 (N_20280,N_19544,N_19115);
nor U20281 (N_20281,N_19193,N_18013);
and U20282 (N_20282,N_18867,N_19709);
xnor U20283 (N_20283,N_18768,N_18759);
xnor U20284 (N_20284,N_19191,N_18972);
or U20285 (N_20285,N_18615,N_18297);
nand U20286 (N_20286,N_18827,N_18876);
nand U20287 (N_20287,N_19648,N_19545);
nor U20288 (N_20288,N_18842,N_19368);
nor U20289 (N_20289,N_18852,N_18060);
and U20290 (N_20290,N_19849,N_19797);
nor U20291 (N_20291,N_19704,N_18390);
xor U20292 (N_20292,N_18258,N_19224);
xnor U20293 (N_20293,N_18326,N_19491);
or U20294 (N_20294,N_18055,N_19643);
and U20295 (N_20295,N_19331,N_19877);
and U20296 (N_20296,N_19563,N_19744);
or U20297 (N_20297,N_18217,N_19543);
or U20298 (N_20298,N_19943,N_19284);
or U20299 (N_20299,N_19817,N_19721);
xor U20300 (N_20300,N_18758,N_19893);
nand U20301 (N_20301,N_18340,N_19566);
nor U20302 (N_20302,N_18222,N_19854);
xnor U20303 (N_20303,N_19902,N_18765);
nand U20304 (N_20304,N_18588,N_18574);
or U20305 (N_20305,N_19930,N_19370);
nand U20306 (N_20306,N_19228,N_19922);
and U20307 (N_20307,N_18926,N_19611);
and U20308 (N_20308,N_18368,N_18621);
nand U20309 (N_20309,N_19440,N_18196);
xor U20310 (N_20310,N_19940,N_18462);
xor U20311 (N_20311,N_19885,N_19141);
nor U20312 (N_20312,N_19874,N_18911);
nor U20313 (N_20313,N_19403,N_19276);
xnor U20314 (N_20314,N_18966,N_18256);
nor U20315 (N_20315,N_19080,N_18002);
nand U20316 (N_20316,N_19226,N_18347);
nor U20317 (N_20317,N_19289,N_18167);
nand U20318 (N_20318,N_19757,N_19099);
xor U20319 (N_20319,N_19833,N_18104);
xor U20320 (N_20320,N_18540,N_19682);
and U20321 (N_20321,N_19796,N_19878);
xor U20322 (N_20322,N_19918,N_18253);
or U20323 (N_20323,N_19908,N_18082);
and U20324 (N_20324,N_18464,N_19838);
nor U20325 (N_20325,N_18755,N_18607);
or U20326 (N_20326,N_18349,N_18650);
xnor U20327 (N_20327,N_18119,N_18654);
and U20328 (N_20328,N_18236,N_18134);
nand U20329 (N_20329,N_19417,N_18045);
nand U20330 (N_20330,N_19855,N_18775);
nor U20331 (N_20331,N_19653,N_18392);
or U20332 (N_20332,N_19425,N_18704);
or U20333 (N_20333,N_18816,N_18403);
nand U20334 (N_20334,N_19586,N_19298);
nand U20335 (N_20335,N_18586,N_19809);
and U20336 (N_20336,N_18446,N_18909);
xnor U20337 (N_20337,N_18995,N_19270);
and U20338 (N_20338,N_18490,N_19791);
and U20339 (N_20339,N_18685,N_18313);
nand U20340 (N_20340,N_18046,N_18400);
and U20341 (N_20341,N_19343,N_19340);
or U20342 (N_20342,N_18751,N_19431);
nor U20343 (N_20343,N_19799,N_18990);
xor U20344 (N_20344,N_18448,N_19714);
or U20345 (N_20345,N_18728,N_19631);
nand U20346 (N_20346,N_18140,N_18791);
xnor U20347 (N_20347,N_18427,N_19802);
xor U20348 (N_20348,N_18873,N_19161);
nand U20349 (N_20349,N_19166,N_19137);
or U20350 (N_20350,N_19599,N_18841);
nand U20351 (N_20351,N_19290,N_18936);
nand U20352 (N_20352,N_19989,N_19889);
nor U20353 (N_20353,N_19110,N_18907);
and U20354 (N_20354,N_19815,N_18479);
nor U20355 (N_20355,N_18342,N_18808);
nand U20356 (N_20356,N_19458,N_18617);
and U20357 (N_20357,N_19533,N_18655);
or U20358 (N_20358,N_18491,N_19988);
xnor U20359 (N_20359,N_18977,N_18910);
or U20360 (N_20360,N_18416,N_18022);
or U20361 (N_20361,N_19696,N_19384);
nand U20362 (N_20362,N_18451,N_19079);
and U20363 (N_20363,N_19987,N_18087);
nand U20364 (N_20364,N_19472,N_19551);
nand U20365 (N_20365,N_19881,N_18401);
or U20366 (N_20366,N_18158,N_19931);
xnor U20367 (N_20367,N_19208,N_19350);
or U20368 (N_20368,N_19042,N_18918);
or U20369 (N_20369,N_18942,N_19745);
xnor U20370 (N_20370,N_18578,N_19897);
nor U20371 (N_20371,N_19624,N_18176);
and U20372 (N_20372,N_18888,N_18093);
nand U20373 (N_20373,N_19507,N_18292);
nand U20374 (N_20374,N_19946,N_19026);
xor U20375 (N_20375,N_18080,N_18750);
nor U20376 (N_20376,N_19474,N_19314);
and U20377 (N_20377,N_18141,N_18377);
or U20378 (N_20378,N_19595,N_18949);
and U20379 (N_20379,N_18860,N_18884);
and U20380 (N_20380,N_18859,N_19377);
nand U20381 (N_20381,N_19285,N_18645);
nand U20382 (N_20382,N_18722,N_18135);
nand U20383 (N_20383,N_18213,N_18955);
nor U20384 (N_20384,N_19044,N_18947);
nor U20385 (N_20385,N_18467,N_19520);
and U20386 (N_20386,N_18012,N_19587);
or U20387 (N_20387,N_19100,N_19334);
nor U20388 (N_20388,N_19198,N_19072);
nand U20389 (N_20389,N_19771,N_19863);
xnor U20390 (N_20390,N_19687,N_19973);
xnor U20391 (N_20391,N_18201,N_19702);
nand U20392 (N_20392,N_19160,N_19526);
or U20393 (N_20393,N_19247,N_18133);
nand U20394 (N_20394,N_18730,N_19357);
nor U20395 (N_20395,N_19652,N_19038);
nand U20396 (N_20396,N_18100,N_18375);
or U20397 (N_20397,N_19282,N_18245);
and U20398 (N_20398,N_19763,N_19420);
or U20399 (N_20399,N_19243,N_18823);
nand U20400 (N_20400,N_19255,N_18981);
and U20401 (N_20401,N_19594,N_19541);
and U20402 (N_20402,N_19557,N_19660);
and U20403 (N_20403,N_19729,N_19783);
or U20404 (N_20404,N_19077,N_19880);
xnor U20405 (N_20405,N_19452,N_19549);
nor U20406 (N_20406,N_19923,N_18070);
or U20407 (N_20407,N_18040,N_18549);
nor U20408 (N_20408,N_18280,N_18466);
and U20409 (N_20409,N_19002,N_19210);
nor U20410 (N_20410,N_18684,N_19697);
xor U20411 (N_20411,N_19882,N_19481);
xnor U20412 (N_20412,N_19351,N_18030);
nand U20413 (N_20413,N_19564,N_18906);
xnor U20414 (N_20414,N_18760,N_19494);
xnor U20415 (N_20415,N_19281,N_18382);
nor U20416 (N_20416,N_18517,N_18143);
nor U20417 (N_20417,N_18036,N_18286);
nor U20418 (N_20418,N_18159,N_19216);
nand U20419 (N_20419,N_18212,N_19266);
nand U20420 (N_20420,N_18644,N_19824);
and U20421 (N_20421,N_18629,N_18591);
xor U20422 (N_20422,N_19659,N_19904);
nor U20423 (N_20423,N_18274,N_18801);
or U20424 (N_20424,N_19681,N_18238);
or U20425 (N_20425,N_19983,N_18626);
nand U20426 (N_20426,N_19784,N_18289);
or U20427 (N_20427,N_19782,N_19781);
xnor U20428 (N_20428,N_19386,N_18439);
nand U20429 (N_20429,N_19618,N_18108);
or U20430 (N_20430,N_19256,N_18021);
or U20431 (N_20431,N_18249,N_18830);
or U20432 (N_20432,N_19311,N_19725);
nor U20433 (N_20433,N_19612,N_18530);
and U20434 (N_20434,N_19947,N_19405);
or U20435 (N_20435,N_19915,N_19048);
nor U20436 (N_20436,N_19845,N_19132);
or U20437 (N_20437,N_18814,N_18144);
xor U20438 (N_20438,N_18537,N_18757);
and U20439 (N_20439,N_19683,N_19993);
and U20440 (N_20440,N_19239,N_18987);
xnor U20441 (N_20441,N_18531,N_19204);
nor U20442 (N_20442,N_18251,N_18625);
xor U20443 (N_20443,N_18312,N_18304);
nand U20444 (N_20444,N_19793,N_19296);
xor U20445 (N_20445,N_18848,N_18091);
nor U20446 (N_20446,N_19856,N_19669);
and U20447 (N_20447,N_18374,N_19412);
nand U20448 (N_20448,N_19136,N_18599);
nand U20449 (N_20449,N_19049,N_18659);
nor U20450 (N_20450,N_18042,N_18952);
nor U20451 (N_20451,N_19171,N_18772);
xnor U20452 (N_20452,N_19811,N_18350);
xor U20453 (N_20453,N_18978,N_19668);
xor U20454 (N_20454,N_18968,N_18229);
xor U20455 (N_20455,N_18378,N_19954);
nor U20456 (N_20456,N_19381,N_19258);
nor U20457 (N_20457,N_19717,N_19237);
nor U20458 (N_20458,N_18152,N_18802);
nor U20459 (N_20459,N_19731,N_19790);
nand U20460 (N_20460,N_18915,N_19578);
nor U20461 (N_20461,N_18068,N_19045);
or U20462 (N_20462,N_19812,N_18161);
nand U20463 (N_20463,N_19033,N_18543);
xnor U20464 (N_20464,N_19724,N_19956);
xor U20465 (N_20465,N_18088,N_19250);
nor U20466 (N_20466,N_19926,N_18450);
or U20467 (N_20467,N_18357,N_19209);
and U20468 (N_20468,N_18369,N_18145);
and U20469 (N_20469,N_18242,N_18147);
nand U20470 (N_20470,N_18136,N_19754);
xnor U20471 (N_20471,N_18948,N_18173);
or U20472 (N_20472,N_19972,N_18120);
and U20473 (N_20473,N_18472,N_18982);
nand U20474 (N_20474,N_19823,N_18960);
nand U20475 (N_20475,N_18004,N_19411);
nand U20476 (N_20476,N_18433,N_19076);
or U20477 (N_20477,N_18355,N_19521);
or U20478 (N_20478,N_18536,N_18917);
and U20479 (N_20479,N_18614,N_19772);
xor U20480 (N_20480,N_19711,N_19766);
nand U20481 (N_20481,N_19111,N_18541);
nor U20482 (N_20482,N_19039,N_19359);
or U20483 (N_20483,N_18348,N_19778);
nand U20484 (N_20484,N_18672,N_18480);
xnor U20485 (N_20485,N_18605,N_18399);
nor U20486 (N_20486,N_18371,N_18066);
or U20487 (N_20487,N_19471,N_18516);
nand U20488 (N_20488,N_19320,N_18473);
xnor U20489 (N_20489,N_19037,N_19364);
nor U20490 (N_20490,N_19060,N_19584);
and U20491 (N_20491,N_18170,N_18492);
and U20492 (N_20492,N_19605,N_19344);
or U20493 (N_20493,N_19335,N_19219);
and U20494 (N_20494,N_19341,N_19901);
xor U20495 (N_20495,N_19842,N_18602);
nor U20496 (N_20496,N_19436,N_19827);
nor U20497 (N_20497,N_18817,N_19197);
xnor U20498 (N_20498,N_19875,N_18809);
and U20499 (N_20499,N_19780,N_18014);
xor U20500 (N_20500,N_18097,N_18774);
nand U20501 (N_20501,N_19489,N_18865);
or U20502 (N_20502,N_19705,N_18967);
xnor U20503 (N_20503,N_19109,N_19129);
nand U20504 (N_20504,N_18985,N_19135);
xor U20505 (N_20505,N_19698,N_18272);
and U20506 (N_20506,N_19389,N_19969);
nor U20507 (N_20507,N_19951,N_18482);
nand U20508 (N_20508,N_19673,N_19463);
and U20509 (N_20509,N_18105,N_19945);
xnor U20510 (N_20510,N_19387,N_19189);
or U20511 (N_20511,N_19061,N_19843);
and U20512 (N_20512,N_18314,N_18608);
nor U20513 (N_20513,N_18231,N_18813);
or U20514 (N_20514,N_18745,N_18885);
xor U20515 (N_20515,N_18556,N_18807);
and U20516 (N_20516,N_19154,N_19645);
nand U20517 (N_20517,N_18988,N_18637);
nor U20518 (N_20518,N_19092,N_19514);
or U20519 (N_20519,N_18681,N_18396);
or U20520 (N_20520,N_19461,N_18753);
nor U20521 (N_20521,N_19223,N_18893);
or U20522 (N_20522,N_19764,N_18613);
nor U20523 (N_20523,N_18638,N_18927);
nand U20524 (N_20524,N_19082,N_19735);
nand U20525 (N_20525,N_18052,N_19468);
nor U20526 (N_20526,N_18944,N_19888);
and U20527 (N_20527,N_18440,N_19505);
xor U20528 (N_20528,N_19488,N_18160);
nand U20529 (N_20529,N_18573,N_18507);
nand U20530 (N_20530,N_18504,N_18711);
nor U20531 (N_20531,N_18208,N_19795);
nand U20532 (N_20532,N_19275,N_18595);
nand U20533 (N_20533,N_19860,N_18282);
nor U20534 (N_20534,N_18568,N_18077);
xor U20535 (N_20535,N_19607,N_18693);
nor U20536 (N_20536,N_18092,N_19623);
and U20537 (N_20537,N_19573,N_19626);
or U20538 (N_20538,N_18624,N_18497);
and U20539 (N_20539,N_19912,N_18020);
or U20540 (N_20540,N_18215,N_18579);
and U20541 (N_20541,N_18109,N_18612);
and U20542 (N_20542,N_18557,N_18862);
nor U20543 (N_20543,N_19531,N_19628);
or U20544 (N_20544,N_18548,N_18461);
and U20545 (N_20545,N_19199,N_19365);
nand U20546 (N_20546,N_18334,N_19424);
nor U20547 (N_20547,N_18432,N_18288);
nand U20548 (N_20548,N_18422,N_19119);
nor U20549 (N_20549,N_19671,N_19030);
nor U20550 (N_20550,N_19190,N_19530);
xnor U20551 (N_20551,N_19858,N_19966);
xnor U20552 (N_20552,N_19378,N_19808);
or U20553 (N_20553,N_19278,N_18575);
nor U20554 (N_20554,N_18511,N_19504);
nor U20555 (N_20555,N_19460,N_18858);
nor U20556 (N_20556,N_18485,N_18837);
nor U20557 (N_20557,N_18426,N_18137);
or U20558 (N_20558,N_19232,N_18778);
nand U20559 (N_20559,N_18583,N_19656);
xor U20560 (N_20560,N_18407,N_19004);
and U20561 (N_20561,N_18971,N_18408);
xor U20562 (N_20562,N_19127,N_18596);
and U20563 (N_20563,N_18050,N_19760);
and U20564 (N_20564,N_18630,N_18788);
and U20565 (N_20565,N_18618,N_18184);
xor U20566 (N_20566,N_18391,N_18425);
xnor U20567 (N_20567,N_18740,N_18405);
nor U20568 (N_20568,N_19024,N_19992);
or U20569 (N_20569,N_19990,N_18805);
or U20570 (N_20570,N_18710,N_18452);
nor U20571 (N_20571,N_18296,N_19133);
xnor U20572 (N_20572,N_18047,N_18804);
or U20573 (N_20573,N_18443,N_19934);
or U20574 (N_20574,N_18063,N_19647);
or U20575 (N_20575,N_18455,N_18247);
and U20576 (N_20576,N_18538,N_18725);
nand U20577 (N_20577,N_18822,N_19689);
or U20578 (N_20578,N_19694,N_19719);
nor U20579 (N_20579,N_19165,N_18192);
nand U20580 (N_20580,N_19920,N_18956);
and U20581 (N_20581,N_18096,N_19269);
or U20582 (N_20582,N_18913,N_18225);
and U20583 (N_20583,N_19388,N_19787);
or U20584 (N_20584,N_19644,N_19655);
nand U20585 (N_20585,N_18268,N_19775);
and U20586 (N_20586,N_18024,N_19325);
nor U20587 (N_20587,N_18431,N_18393);
nand U20588 (N_20588,N_18243,N_18847);
xor U20589 (N_20589,N_18043,N_19478);
nor U20590 (N_20590,N_18246,N_18941);
xnor U20591 (N_20591,N_18781,N_18554);
or U20592 (N_20592,N_19649,N_19342);
nand U20593 (N_20593,N_18178,N_19326);
or U20594 (N_20594,N_18007,N_19279);
nand U20595 (N_20595,N_19770,N_19688);
or U20596 (N_20596,N_19502,N_19009);
xor U20597 (N_20597,N_18899,N_19434);
nand U20598 (N_20598,N_19571,N_18890);
nand U20599 (N_20599,N_18169,N_19288);
nand U20600 (N_20600,N_18594,N_18318);
or U20601 (N_20601,N_19937,N_19018);
and U20602 (N_20602,N_18600,N_19635);
or U20603 (N_20603,N_19121,N_18211);
nand U20604 (N_20604,N_18732,N_19339);
xor U20605 (N_20605,N_19807,N_19448);
or U20606 (N_20606,N_19105,N_19609);
nor U20607 (N_20607,N_19707,N_18969);
and U20608 (N_20608,N_19503,N_19188);
xnor U20609 (N_20609,N_18878,N_19443);
and U20610 (N_20610,N_18027,N_19307);
and U20611 (N_20611,N_19134,N_18185);
nand U20612 (N_20612,N_19924,N_19606);
or U20613 (N_20613,N_18883,N_18309);
and U20614 (N_20614,N_19466,N_19927);
or U20615 (N_20615,N_19701,N_18611);
or U20616 (N_20616,N_18924,N_19841);
nor U20617 (N_20617,N_18997,N_18468);
nand U20618 (N_20618,N_19410,N_19272);
or U20619 (N_20619,N_18581,N_19985);
and U20620 (N_20620,N_18085,N_19089);
and U20621 (N_20621,N_18717,N_18572);
or U20622 (N_20622,N_19169,N_19008);
nand U20623 (N_20623,N_18283,N_19251);
or U20624 (N_20624,N_19716,N_18189);
nor U20625 (N_20625,N_18560,N_19203);
or U20626 (N_20626,N_18026,N_18785);
nor U20627 (N_20627,N_18619,N_19323);
nor U20628 (N_20628,N_19112,N_19057);
xor U20629 (N_20629,N_18197,N_19025);
nor U20630 (N_20630,N_18799,N_19446);
xor U20631 (N_20631,N_19710,N_19582);
nor U20632 (N_20632,N_18821,N_18741);
or U20633 (N_20633,N_18935,N_19952);
nand U20634 (N_20634,N_18975,N_19540);
nand U20635 (N_20635,N_19767,N_19152);
nor U20636 (N_20636,N_19083,N_18670);
nor U20637 (N_20637,N_18647,N_19029);
nand U20638 (N_20638,N_18940,N_19318);
xor U20639 (N_20639,N_19358,N_19670);
nand U20640 (N_20640,N_19286,N_19144);
nand U20641 (N_20641,N_19603,N_18171);
and U20642 (N_20642,N_19485,N_19925);
xor U20643 (N_20643,N_18623,N_18175);
xnor U20644 (N_20644,N_18686,N_19202);
or U20645 (N_20645,N_19031,N_19123);
xor U20646 (N_20646,N_18863,N_18976);
nor U20647 (N_20647,N_19588,N_19248);
and U20648 (N_20648,N_19675,N_19229);
or U20649 (N_20649,N_19686,N_18291);
nand U20650 (N_20650,N_19641,N_18220);
nor U20651 (N_20651,N_19265,N_19056);
and U20652 (N_20652,N_19884,N_19562);
and U20653 (N_20653,N_19532,N_18338);
xnor U20654 (N_20654,N_19495,N_19829);
nand U20655 (N_20655,N_18123,N_18099);
or U20656 (N_20656,N_18790,N_19475);
nand U20657 (N_20657,N_19196,N_18846);
xor U20658 (N_20658,N_19437,N_19106);
xor U20659 (N_20659,N_18306,N_19449);
nand U20660 (N_20660,N_19055,N_19861);
or U20661 (N_20661,N_18727,N_19907);
xor U20662 (N_20662,N_19914,N_18035);
nor U20663 (N_20663,N_18789,N_19786);
nand U20664 (N_20664,N_18833,N_18845);
nor U20665 (N_20665,N_19835,N_19433);
and U20666 (N_20666,N_18339,N_18715);
xor U20667 (N_20667,N_18547,N_19722);
or U20668 (N_20668,N_18302,N_19558);
or U20669 (N_20669,N_18707,N_18748);
xor U20670 (N_20670,N_19637,N_18850);
nand U20671 (N_20671,N_18034,N_19373);
or U20672 (N_20672,N_19741,N_18244);
and U20673 (N_20673,N_18111,N_18265);
xor U20674 (N_20674,N_19743,N_18386);
nor U20675 (N_20675,N_18005,N_18829);
or U20676 (N_20676,N_19876,N_18746);
xor U20677 (N_20677,N_18737,N_19794);
nand U20678 (N_20678,N_19490,N_19215);
nor U20679 (N_20679,N_19332,N_19213);
and U20680 (N_20680,N_19699,N_18930);
and U20681 (N_20681,N_18203,N_18838);
or U20682 (N_20682,N_19194,N_18454);
nand U20683 (N_20683,N_18230,N_18311);
nand U20684 (N_20684,N_19362,N_19852);
or U20685 (N_20685,N_19302,N_18632);
nand U20686 (N_20686,N_19091,N_18345);
xor U20687 (N_20687,N_18142,N_19650);
nor U20688 (N_20688,N_18920,N_18457);
xor U20689 (N_20689,N_18818,N_19020);
nor U20690 (N_20690,N_18009,N_19749);
xnor U20691 (N_20691,N_18662,N_19703);
and U20692 (N_20692,N_19162,N_19515);
xor U20693 (N_20693,N_18520,N_19642);
nor U20694 (N_20694,N_19848,N_19327);
and U20695 (N_20695,N_19873,N_19826);
nor U20696 (N_20696,N_19984,N_18278);
nand U20697 (N_20697,N_19356,N_18665);
and U20698 (N_20698,N_19548,N_18279);
or U20699 (N_20699,N_18266,N_18102);
and U20700 (N_20700,N_18984,N_18465);
and U20701 (N_20701,N_19928,N_18870);
xnor U20702 (N_20702,N_19001,N_18051);
and U20703 (N_20703,N_19422,N_18498);
xor U20704 (N_20704,N_18898,N_18181);
or U20705 (N_20705,N_19896,N_18460);
or U20706 (N_20706,N_18438,N_18831);
nand U20707 (N_20707,N_18115,N_18934);
nand U20708 (N_20708,N_18254,N_18323);
and U20709 (N_20709,N_19981,N_19201);
nand U20710 (N_20710,N_18057,N_19971);
and U20711 (N_20711,N_19830,N_19667);
xnor U20712 (N_20712,N_18545,N_18646);
or U20713 (N_20713,N_18786,N_19534);
and U20714 (N_20714,N_19379,N_19938);
xor U20715 (N_20715,N_18232,N_19321);
xnor U20716 (N_20716,N_18901,N_19021);
or U20717 (N_20717,N_19192,N_18025);
nor U20718 (N_20718,N_19941,N_18882);
or U20719 (N_20719,N_18039,N_19451);
xnor U20720 (N_20720,N_18128,N_19147);
and U20721 (N_20721,N_18453,N_19244);
nor U20722 (N_20722,N_19759,N_18259);
xnor U20723 (N_20723,N_19374,N_19995);
xor U20724 (N_20724,N_18316,N_19519);
or U20725 (N_20725,N_18515,N_18154);
nor U20726 (N_20726,N_18110,N_19090);
nand U20727 (N_20727,N_19071,N_18648);
and U20728 (N_20728,N_19383,N_19944);
or U20729 (N_20729,N_18787,N_19591);
nor U20730 (N_20730,N_18003,N_19128);
and U20731 (N_20731,N_18322,N_19615);
or U20732 (N_20732,N_19674,N_19453);
or U20733 (N_20733,N_18521,N_19264);
and U20734 (N_20734,N_19868,N_18430);
or U20735 (N_20735,N_19146,N_19968);
xnor U20736 (N_20736,N_18875,N_19333);
and U20737 (N_20737,N_19846,N_19765);
and U20738 (N_20738,N_18300,N_19665);
and U20739 (N_20739,N_18149,N_19257);
or U20740 (N_20740,N_18678,N_19235);
nand U20741 (N_20741,N_18731,N_18674);
nand U20742 (N_20742,N_19396,N_18384);
nor U20743 (N_20743,N_18290,N_19097);
nand U20744 (N_20744,N_18199,N_19769);
nand U20745 (N_20745,N_18571,N_19657);
nand U20746 (N_20746,N_19421,N_18668);
and U20747 (N_20747,N_18879,N_19567);
or U20748 (N_20748,N_18079,N_18980);
nor U20749 (N_20749,N_19297,N_18925);
xor U20750 (N_20750,N_19916,N_18851);
or U20751 (N_20751,N_18825,N_18764);
or U20752 (N_20752,N_19487,N_19268);
and U20753 (N_20753,N_18359,N_18839);
or U20754 (N_20754,N_18444,N_18706);
nand U20755 (N_20755,N_18098,N_18330);
nand U20756 (N_20756,N_18957,N_18086);
or U20757 (N_20757,N_19206,N_18394);
and U20758 (N_20758,N_18880,N_18476);
or U20759 (N_20759,N_18112,N_18694);
and U20760 (N_20760,N_18395,N_18415);
or U20761 (N_20761,N_19953,N_19212);
xor U20762 (N_20762,N_18337,N_19732);
nand U20763 (N_20763,N_19894,N_19962);
xor U20764 (N_20764,N_18505,N_18567);
and U20765 (N_20765,N_18705,N_18993);
nand U20766 (N_20766,N_19821,N_18139);
or U20767 (N_20767,N_18699,N_18033);
nand U20768 (N_20768,N_18223,N_19477);
and U20769 (N_20769,N_18958,N_19975);
or U20770 (N_20770,N_19363,N_18855);
or U20771 (N_20771,N_18166,N_19986);
nor U20772 (N_20772,N_18409,N_19303);
nand U20773 (N_20773,N_19367,N_19678);
nor U20774 (N_20774,N_18734,N_18580);
or U20775 (N_20775,N_18877,N_18661);
and U20776 (N_20776,N_19236,N_19761);
nand U20777 (N_20777,N_18397,N_18979);
nor U20778 (N_20778,N_18938,N_19385);
xnor U20779 (N_20779,N_19840,N_18157);
xnor U20780 (N_20780,N_19999,N_18240);
nand U20781 (N_20781,N_19753,N_18501);
or U20782 (N_20782,N_18071,N_18008);
or U20783 (N_20783,N_19050,N_18089);
nor U20784 (N_20784,N_19107,N_19748);
and U20785 (N_20785,N_18766,N_19596);
or U20786 (N_20786,N_19047,N_18695);
nand U20787 (N_20787,N_19028,N_19122);
or U20788 (N_20788,N_18861,N_19909);
nor U20789 (N_20789,N_19299,N_18535);
or U20790 (N_20790,N_18555,N_19304);
or U20791 (N_20791,N_19345,N_18303);
nor U20792 (N_20792,N_18074,N_18413);
nor U20793 (N_20793,N_19430,N_18798);
nor U20794 (N_20794,N_19058,N_18441);
xnor U20795 (N_20795,N_19170,N_19598);
xnor U20796 (N_20796,N_18293,N_18702);
and U20797 (N_20797,N_19685,N_18939);
and U20798 (N_20798,N_19347,N_18931);
nor U20799 (N_20799,N_19465,N_19523);
xor U20800 (N_20800,N_19094,N_19469);
or U20801 (N_20801,N_18912,N_19865);
xnor U20802 (N_20802,N_18118,N_18636);
or U20803 (N_20803,N_19950,N_18559);
xnor U20804 (N_20804,N_18162,N_19492);
or U20805 (N_20805,N_19510,N_18767);
or U20806 (N_20806,N_18563,N_19706);
xnor U20807 (N_20807,N_18570,N_19395);
xnor U20808 (N_20808,N_19066,N_19666);
nor U20809 (N_20809,N_19565,N_18900);
or U20810 (N_20810,N_19522,N_18299);
nand U20811 (N_20811,N_19337,N_19175);
and U20812 (N_20812,N_18914,N_18698);
and U20813 (N_20813,N_19267,N_18285);
and U20814 (N_20814,N_18729,N_18072);
or U20815 (N_20815,N_18214,N_18523);
and U20816 (N_20816,N_19313,N_18542);
xor U20817 (N_20817,N_18172,N_18153);
or U20818 (N_20818,N_18897,N_18062);
and U20819 (N_20819,N_19168,N_18522);
nor U20820 (N_20820,N_18206,N_18352);
xor U20821 (N_20821,N_19241,N_19579);
nor U20822 (N_20822,N_19739,N_19273);
and U20823 (N_20823,N_18168,N_18127);
xor U20824 (N_20824,N_18048,N_19114);
or U20825 (N_20825,N_19619,N_19755);
nor U20826 (N_20826,N_19231,N_18138);
and U20827 (N_20827,N_19143,N_18667);
and U20828 (N_20828,N_19108,N_18584);
nor U20829 (N_20829,N_18388,N_18284);
and U20830 (N_20830,N_18539,N_19416);
or U20831 (N_20831,N_18658,N_18150);
or U20832 (N_20832,N_18683,N_18056);
xor U20833 (N_20833,N_18896,N_19088);
xnor U20834 (N_20834,N_19400,N_19148);
or U20835 (N_20835,N_19116,N_19150);
or U20836 (N_20836,N_19750,N_18566);
nand U20837 (N_20837,N_18346,N_19073);
nor U20838 (N_20838,N_19633,N_18546);
xor U20839 (N_20839,N_19102,N_18961);
nor U20840 (N_20840,N_19254,N_19561);
or U20841 (N_20841,N_18032,N_18257);
or U20842 (N_20842,N_18353,N_19837);
and U20843 (N_20843,N_18656,N_19801);
nor U20844 (N_20844,N_19011,N_18500);
or U20845 (N_20845,N_19513,N_18018);
or U20846 (N_20846,N_18735,N_18435);
or U20847 (N_20847,N_19589,N_19182);
nor U20848 (N_20848,N_18716,N_18343);
nand U20849 (N_20849,N_18929,N_19401);
and U20850 (N_20850,N_19742,N_19138);
nor U20851 (N_20851,N_19933,N_18132);
or U20852 (N_20852,N_19980,N_18402);
or U20853 (N_20853,N_19177,N_18084);
nand U20854 (N_20854,N_19959,N_19157);
nor U20855 (N_20855,N_19467,N_18198);
or U20856 (N_20856,N_18207,N_18011);
xor U20857 (N_20857,N_19046,N_19426);
nand U20858 (N_20858,N_18049,N_18738);
xor U20859 (N_20859,N_18675,N_18639);
and U20860 (N_20860,N_18241,N_19752);
nor U20861 (N_20861,N_18502,N_19518);
or U20862 (N_20862,N_18820,N_18067);
nor U20863 (N_20863,N_18983,N_19149);
or U20864 (N_20864,N_19315,N_18488);
or U20865 (N_20865,N_18747,N_18250);
and U20866 (N_20866,N_19429,N_19857);
or U20867 (N_20867,N_18783,N_19442);
or U20868 (N_20868,N_18794,N_19233);
nand U20869 (N_20869,N_19271,N_18603);
nor U20870 (N_20870,N_18872,N_18954);
nand U20871 (N_20871,N_19023,N_19629);
xor U20872 (N_20872,N_19484,N_18998);
xor U20873 (N_20873,N_18333,N_18606);
nor U20874 (N_20874,N_19836,N_18187);
or U20875 (N_20875,N_19126,N_19098);
nor U20876 (N_20876,N_18965,N_18200);
and U20877 (N_20877,N_18708,N_19720);
xor U20878 (N_20878,N_18463,N_19740);
and U20879 (N_20879,N_19636,N_19639);
and U20880 (N_20880,N_18652,N_18365);
nor U20881 (N_20881,N_18569,N_19905);
and U20882 (N_20882,N_18195,N_19850);
or U20883 (N_20883,N_18237,N_19994);
xnor U20884 (N_20884,N_18687,N_19913);
xor U20885 (N_20885,N_18651,N_18114);
nor U20886 (N_20886,N_18239,N_19015);
nor U20887 (N_20887,N_19246,N_18383);
or U20888 (N_20888,N_19462,N_18325);
nor U20889 (N_20889,N_19600,N_19575);
and U20890 (N_20890,N_18962,N_19178);
nand U20891 (N_20891,N_18493,N_19065);
or U20892 (N_20892,N_18749,N_18529);
xnor U20893 (N_20893,N_19159,N_19493);
nor U20894 (N_20894,N_19070,N_19444);
or U20895 (N_20895,N_19308,N_18227);
nand U20896 (N_20896,N_18031,N_18404);
or U20897 (N_20897,N_19486,N_18697);
and U20898 (N_20898,N_19051,N_18174);
xnor U20899 (N_20899,N_19900,N_19360);
or U20900 (N_20900,N_19032,N_19756);
nor U20901 (N_20901,N_19939,N_18691);
nand U20902 (N_20902,N_19805,N_18889);
xor U20903 (N_20903,N_18597,N_19470);
nand U20904 (N_20904,N_18503,N_19872);
or U20905 (N_20905,N_19142,N_19834);
or U20906 (N_20906,N_18058,N_18680);
nand U20907 (N_20907,N_18905,N_18477);
xnor U20908 (N_20908,N_19093,N_19125);
and U20909 (N_20909,N_19614,N_19866);
xor U20910 (N_20910,N_19483,N_19554);
and U20911 (N_20911,N_18073,N_18248);
or U20912 (N_20912,N_19054,N_19352);
and U20913 (N_20913,N_19427,N_19524);
nand U20914 (N_20914,N_18226,N_18328);
nor U20915 (N_20915,N_19976,N_19663);
nor U20916 (N_20916,N_19176,N_19187);
nand U20917 (N_20917,N_19819,N_18544);
and U20918 (N_20918,N_18121,N_19346);
and U20919 (N_20919,N_18075,N_18945);
xor U20920 (N_20920,N_18210,N_19570);
or U20921 (N_20921,N_19910,N_18023);
xnor U20922 (N_20922,N_18959,N_19181);
nand U20923 (N_20923,N_18856,N_19751);
nand U20924 (N_20924,N_19651,N_18550);
nand U20925 (N_20925,N_19014,N_18381);
nor U20926 (N_20926,N_18679,N_19917);
xor U20927 (N_20927,N_19879,N_19497);
nand U20928 (N_20928,N_18991,N_19238);
xor U20929 (N_20929,N_19164,N_19936);
xor U20930 (N_20930,N_18376,N_18970);
xor U20931 (N_20931,N_18233,N_18429);
and U20932 (N_20932,N_18298,N_19738);
nor U20933 (N_20933,N_19041,N_18582);
or U20934 (N_20934,N_19184,N_18558);
nor U20935 (N_20935,N_19831,N_18459);
nor U20936 (N_20936,N_18590,N_18495);
and U20937 (N_20937,N_18410,N_19768);
and U20938 (N_20938,N_18469,N_19183);
xnor U20939 (N_20939,N_19007,N_18420);
xor U20940 (N_20940,N_18478,N_18103);
and U20941 (N_20941,N_18124,N_18508);
nand U20942 (N_20942,N_19869,N_19067);
and U20943 (N_20943,N_19113,N_18669);
nor U20944 (N_20944,N_18287,N_19242);
or U20945 (N_20945,N_18506,N_19800);
nor U20946 (N_20946,N_19101,N_18363);
and U20947 (N_20947,N_19690,N_18974);
or U20948 (N_20948,N_18456,N_19822);
and U20949 (N_20949,N_18989,N_19120);
or U20950 (N_20950,N_19630,N_19390);
nor U20951 (N_20951,N_18552,N_19547);
nor U20952 (N_20952,N_19329,N_18010);
xnor U20953 (N_20953,N_18604,N_19693);
nand U20954 (N_20954,N_18688,N_19726);
nor U20955 (N_20955,N_19844,N_19616);
xor U20956 (N_20956,N_19225,N_19309);
or U20957 (N_20957,N_18663,N_19293);
and U20958 (N_20958,N_18643,N_18470);
or U20959 (N_20959,N_19862,N_19700);
nor U20960 (N_20960,N_19592,N_18081);
xnor U20961 (N_20961,N_18810,N_19730);
or U20962 (N_20962,N_18344,N_18156);
and U20963 (N_20963,N_19500,N_19324);
xor U20964 (N_20964,N_18916,N_19758);
nand U20965 (N_20965,N_19375,N_19394);
or U20966 (N_20966,N_18892,N_18264);
and U20967 (N_20967,N_19585,N_19695);
nand U20968 (N_20968,N_19608,N_18513);
nand U20969 (N_20969,N_19658,N_18412);
or U20970 (N_20970,N_18589,N_18576);
xor U20971 (N_20971,N_18235,N_19174);
or U20972 (N_20972,N_18986,N_19820);
and U20973 (N_20973,N_18577,N_18811);
or U20974 (N_20974,N_18853,N_19864);
and U20975 (N_20975,N_18483,N_19211);
xnor U20976 (N_20976,N_18999,N_18712);
nand U20977 (N_20977,N_19539,N_18812);
xor U20978 (N_20978,N_19602,N_18434);
and U20979 (N_20979,N_19252,N_19022);
xor U20980 (N_20980,N_19847,N_18267);
or U20981 (N_20981,N_18784,N_19059);
and U20982 (N_20982,N_19016,N_19063);
and U20983 (N_20983,N_18874,N_19402);
nand U20984 (N_20984,N_19553,N_19406);
xnor U20985 (N_20985,N_18857,N_18499);
nor U20986 (N_20986,N_19680,N_18653);
nor U20987 (N_20987,N_18273,N_18261);
nand U20988 (N_20988,N_19509,N_18165);
or U20989 (N_20989,N_19762,N_19052);
nand U20990 (N_20990,N_19454,N_18752);
or U20991 (N_20991,N_18107,N_19301);
or U20992 (N_20992,N_18733,N_18205);
nor U20993 (N_20993,N_18131,N_18447);
nand U20994 (N_20994,N_18262,N_19733);
xor U20995 (N_20995,N_19399,N_19853);
nand U20996 (N_20996,N_18869,N_19081);
and U20997 (N_20997,N_19967,N_18803);
and U20998 (N_20998,N_18015,N_18017);
nor U20999 (N_20999,N_18616,N_19747);
or U21000 (N_21000,N_18329,N_18368);
nand U21001 (N_21001,N_19032,N_18089);
and U21002 (N_21002,N_18164,N_18981);
nand U21003 (N_21003,N_19449,N_19919);
nor U21004 (N_21004,N_18856,N_18298);
or U21005 (N_21005,N_19226,N_18832);
xnor U21006 (N_21006,N_19927,N_18157);
nand U21007 (N_21007,N_18486,N_18722);
or U21008 (N_21008,N_18566,N_19063);
and U21009 (N_21009,N_18243,N_19999);
xor U21010 (N_21010,N_18186,N_19760);
or U21011 (N_21011,N_18072,N_18994);
xnor U21012 (N_21012,N_18306,N_19628);
nand U21013 (N_21013,N_18541,N_18512);
or U21014 (N_21014,N_19244,N_19013);
xor U21015 (N_21015,N_18082,N_18249);
and U21016 (N_21016,N_19959,N_18111);
xor U21017 (N_21017,N_18750,N_18722);
xnor U21018 (N_21018,N_18781,N_19626);
xor U21019 (N_21019,N_19185,N_19271);
nor U21020 (N_21020,N_19540,N_18037);
xnor U21021 (N_21021,N_19658,N_19082);
or U21022 (N_21022,N_19365,N_18014);
nor U21023 (N_21023,N_18472,N_19360);
or U21024 (N_21024,N_18246,N_19600);
and U21025 (N_21025,N_18156,N_18704);
xor U21026 (N_21026,N_19458,N_19561);
or U21027 (N_21027,N_19632,N_19954);
and U21028 (N_21028,N_19764,N_19308);
and U21029 (N_21029,N_18336,N_19514);
or U21030 (N_21030,N_19164,N_19235);
and U21031 (N_21031,N_18657,N_18337);
nand U21032 (N_21032,N_19097,N_19235);
nand U21033 (N_21033,N_18489,N_18889);
nand U21034 (N_21034,N_19514,N_19747);
or U21035 (N_21035,N_18729,N_19777);
or U21036 (N_21036,N_18376,N_18875);
nor U21037 (N_21037,N_18476,N_18235);
or U21038 (N_21038,N_19901,N_18981);
xnor U21039 (N_21039,N_18839,N_18999);
xnor U21040 (N_21040,N_18435,N_18975);
xnor U21041 (N_21041,N_18674,N_18764);
nand U21042 (N_21042,N_19904,N_19245);
and U21043 (N_21043,N_18726,N_19260);
nand U21044 (N_21044,N_19473,N_19401);
xnor U21045 (N_21045,N_19514,N_18417);
nor U21046 (N_21046,N_18042,N_18443);
nand U21047 (N_21047,N_19390,N_19722);
xor U21048 (N_21048,N_18425,N_19188);
xnor U21049 (N_21049,N_18687,N_18189);
or U21050 (N_21050,N_19437,N_19580);
and U21051 (N_21051,N_19060,N_18849);
nor U21052 (N_21052,N_18515,N_18367);
and U21053 (N_21053,N_19499,N_19588);
xnor U21054 (N_21054,N_18625,N_19884);
xor U21055 (N_21055,N_19984,N_18065);
and U21056 (N_21056,N_18666,N_19149);
nor U21057 (N_21057,N_19639,N_18539);
nor U21058 (N_21058,N_19744,N_19203);
or U21059 (N_21059,N_18043,N_18157);
and U21060 (N_21060,N_19638,N_18381);
xnor U21061 (N_21061,N_18005,N_18689);
and U21062 (N_21062,N_19438,N_19301);
and U21063 (N_21063,N_19134,N_19229);
nand U21064 (N_21064,N_19411,N_19241);
and U21065 (N_21065,N_19917,N_18017);
nor U21066 (N_21066,N_19102,N_19004);
or U21067 (N_21067,N_18417,N_19934);
xor U21068 (N_21068,N_19089,N_19742);
or U21069 (N_21069,N_19815,N_19804);
xor U21070 (N_21070,N_19026,N_18673);
nand U21071 (N_21071,N_18037,N_18604);
nor U21072 (N_21072,N_19764,N_19969);
or U21073 (N_21073,N_19569,N_19540);
and U21074 (N_21074,N_19407,N_19051);
xor U21075 (N_21075,N_18426,N_18516);
xor U21076 (N_21076,N_18204,N_18714);
and U21077 (N_21077,N_18642,N_19547);
or U21078 (N_21078,N_18245,N_18339);
nor U21079 (N_21079,N_19371,N_18818);
or U21080 (N_21080,N_18841,N_19785);
or U21081 (N_21081,N_18589,N_18431);
and U21082 (N_21082,N_19207,N_19926);
nand U21083 (N_21083,N_19851,N_18236);
xnor U21084 (N_21084,N_19141,N_18029);
and U21085 (N_21085,N_18416,N_19100);
or U21086 (N_21086,N_18167,N_19860);
nand U21087 (N_21087,N_18088,N_19147);
and U21088 (N_21088,N_19918,N_18356);
nand U21089 (N_21089,N_19154,N_18875);
xor U21090 (N_21090,N_19378,N_18528);
and U21091 (N_21091,N_18048,N_19768);
xnor U21092 (N_21092,N_18887,N_18239);
nor U21093 (N_21093,N_19046,N_18938);
xor U21094 (N_21094,N_19761,N_19872);
nand U21095 (N_21095,N_18443,N_19120);
nand U21096 (N_21096,N_19168,N_19739);
and U21097 (N_21097,N_18124,N_18856);
nand U21098 (N_21098,N_18152,N_19961);
or U21099 (N_21099,N_18520,N_19867);
nor U21100 (N_21100,N_18426,N_19431);
nand U21101 (N_21101,N_19305,N_19966);
nor U21102 (N_21102,N_18064,N_18877);
nor U21103 (N_21103,N_18344,N_18055);
xor U21104 (N_21104,N_19557,N_19369);
or U21105 (N_21105,N_19562,N_19936);
nor U21106 (N_21106,N_19383,N_18537);
nand U21107 (N_21107,N_19856,N_19768);
or U21108 (N_21108,N_19699,N_19965);
xor U21109 (N_21109,N_18553,N_19192);
or U21110 (N_21110,N_18332,N_19295);
xnor U21111 (N_21111,N_19831,N_18210);
or U21112 (N_21112,N_19078,N_18507);
nor U21113 (N_21113,N_18399,N_18700);
and U21114 (N_21114,N_18334,N_18359);
or U21115 (N_21115,N_18124,N_19315);
nor U21116 (N_21116,N_19964,N_18884);
and U21117 (N_21117,N_19389,N_19584);
and U21118 (N_21118,N_18300,N_19755);
nor U21119 (N_21119,N_19304,N_19859);
or U21120 (N_21120,N_19801,N_18422);
or U21121 (N_21121,N_19713,N_18185);
or U21122 (N_21122,N_19428,N_18802);
or U21123 (N_21123,N_18030,N_18522);
or U21124 (N_21124,N_18493,N_19512);
and U21125 (N_21125,N_18752,N_19558);
nand U21126 (N_21126,N_19949,N_19887);
or U21127 (N_21127,N_18278,N_19216);
nor U21128 (N_21128,N_19198,N_19860);
or U21129 (N_21129,N_18060,N_19649);
nand U21130 (N_21130,N_19612,N_18041);
or U21131 (N_21131,N_19518,N_19889);
or U21132 (N_21132,N_18522,N_19800);
and U21133 (N_21133,N_18118,N_19023);
or U21134 (N_21134,N_19710,N_19389);
or U21135 (N_21135,N_18119,N_18484);
and U21136 (N_21136,N_19190,N_19418);
and U21137 (N_21137,N_19051,N_18763);
and U21138 (N_21138,N_18070,N_18156);
nor U21139 (N_21139,N_19635,N_18546);
or U21140 (N_21140,N_18504,N_18951);
nor U21141 (N_21141,N_19729,N_19184);
xnor U21142 (N_21142,N_18896,N_18522);
nand U21143 (N_21143,N_18619,N_18201);
nor U21144 (N_21144,N_18039,N_19111);
nor U21145 (N_21145,N_18973,N_19661);
nor U21146 (N_21146,N_18597,N_18451);
nor U21147 (N_21147,N_19525,N_19203);
nor U21148 (N_21148,N_18803,N_18419);
or U21149 (N_21149,N_18728,N_18457);
or U21150 (N_21150,N_18128,N_19274);
xor U21151 (N_21151,N_18120,N_18802);
nand U21152 (N_21152,N_18977,N_19712);
nand U21153 (N_21153,N_19595,N_19299);
nor U21154 (N_21154,N_19876,N_18498);
nand U21155 (N_21155,N_18666,N_19105);
xor U21156 (N_21156,N_19117,N_19084);
and U21157 (N_21157,N_19574,N_18364);
or U21158 (N_21158,N_19567,N_18430);
nand U21159 (N_21159,N_18140,N_18621);
xor U21160 (N_21160,N_18657,N_18791);
nand U21161 (N_21161,N_19838,N_19484);
and U21162 (N_21162,N_18799,N_19918);
nor U21163 (N_21163,N_19772,N_18952);
nand U21164 (N_21164,N_18223,N_19641);
nand U21165 (N_21165,N_19436,N_19495);
nor U21166 (N_21166,N_18251,N_18314);
nor U21167 (N_21167,N_19171,N_19469);
nor U21168 (N_21168,N_19779,N_19251);
or U21169 (N_21169,N_19922,N_19609);
nor U21170 (N_21170,N_18042,N_18212);
nand U21171 (N_21171,N_18476,N_19439);
nand U21172 (N_21172,N_19851,N_19421);
nand U21173 (N_21173,N_19257,N_18088);
xnor U21174 (N_21174,N_18788,N_18910);
xor U21175 (N_21175,N_18741,N_18790);
xnor U21176 (N_21176,N_18096,N_19432);
xnor U21177 (N_21177,N_18541,N_19121);
nand U21178 (N_21178,N_18762,N_19031);
nor U21179 (N_21179,N_19566,N_18400);
nor U21180 (N_21180,N_19103,N_19086);
xor U21181 (N_21181,N_19685,N_19915);
xnor U21182 (N_21182,N_19292,N_18639);
nor U21183 (N_21183,N_18038,N_19967);
xor U21184 (N_21184,N_18352,N_19873);
and U21185 (N_21185,N_19530,N_19577);
xnor U21186 (N_21186,N_18927,N_19268);
nand U21187 (N_21187,N_19904,N_18475);
and U21188 (N_21188,N_18316,N_19538);
nand U21189 (N_21189,N_19777,N_18406);
xor U21190 (N_21190,N_18143,N_18479);
or U21191 (N_21191,N_18009,N_19848);
or U21192 (N_21192,N_19097,N_19679);
nor U21193 (N_21193,N_18566,N_18113);
nand U21194 (N_21194,N_19044,N_18211);
nor U21195 (N_21195,N_18958,N_18813);
and U21196 (N_21196,N_19146,N_19601);
nor U21197 (N_21197,N_19271,N_18852);
nor U21198 (N_21198,N_18658,N_19276);
and U21199 (N_21199,N_19614,N_19062);
xnor U21200 (N_21200,N_18589,N_18924);
nor U21201 (N_21201,N_18642,N_19096);
and U21202 (N_21202,N_18033,N_19827);
nor U21203 (N_21203,N_18160,N_18873);
xor U21204 (N_21204,N_18906,N_18706);
nand U21205 (N_21205,N_18761,N_18127);
nand U21206 (N_21206,N_18183,N_18077);
and U21207 (N_21207,N_19812,N_18100);
nand U21208 (N_21208,N_19344,N_18892);
xnor U21209 (N_21209,N_18328,N_19428);
nor U21210 (N_21210,N_18607,N_18270);
xnor U21211 (N_21211,N_19706,N_18149);
nand U21212 (N_21212,N_19074,N_18807);
xor U21213 (N_21213,N_18880,N_19737);
and U21214 (N_21214,N_19933,N_19720);
nor U21215 (N_21215,N_19549,N_19129);
and U21216 (N_21216,N_18440,N_19810);
xnor U21217 (N_21217,N_19178,N_19692);
nand U21218 (N_21218,N_18068,N_18526);
nand U21219 (N_21219,N_18036,N_19861);
or U21220 (N_21220,N_19552,N_19700);
or U21221 (N_21221,N_19048,N_19262);
and U21222 (N_21222,N_19172,N_19400);
and U21223 (N_21223,N_18191,N_19327);
xor U21224 (N_21224,N_19100,N_18018);
nor U21225 (N_21225,N_19594,N_18526);
xor U21226 (N_21226,N_19286,N_18505);
and U21227 (N_21227,N_19807,N_18849);
xnor U21228 (N_21228,N_19339,N_18716);
or U21229 (N_21229,N_19447,N_19740);
or U21230 (N_21230,N_19120,N_19493);
nand U21231 (N_21231,N_18610,N_19203);
nor U21232 (N_21232,N_19907,N_19326);
or U21233 (N_21233,N_19040,N_18375);
or U21234 (N_21234,N_19896,N_18644);
and U21235 (N_21235,N_19709,N_18830);
xor U21236 (N_21236,N_18423,N_18812);
xnor U21237 (N_21237,N_18101,N_18179);
and U21238 (N_21238,N_19915,N_18909);
and U21239 (N_21239,N_19074,N_19908);
nand U21240 (N_21240,N_19978,N_18702);
and U21241 (N_21241,N_18933,N_18803);
nand U21242 (N_21242,N_19178,N_18101);
nand U21243 (N_21243,N_18371,N_18058);
nand U21244 (N_21244,N_18484,N_19050);
or U21245 (N_21245,N_19471,N_18569);
xor U21246 (N_21246,N_19271,N_19289);
or U21247 (N_21247,N_19193,N_19496);
nor U21248 (N_21248,N_18393,N_19022);
nor U21249 (N_21249,N_19589,N_19373);
and U21250 (N_21250,N_19695,N_18019);
and U21251 (N_21251,N_19363,N_19020);
nor U21252 (N_21252,N_18293,N_19372);
nor U21253 (N_21253,N_18603,N_19939);
nand U21254 (N_21254,N_18885,N_19421);
nand U21255 (N_21255,N_19822,N_19989);
nand U21256 (N_21256,N_19213,N_19526);
nand U21257 (N_21257,N_18140,N_18138);
xor U21258 (N_21258,N_19806,N_18256);
and U21259 (N_21259,N_18146,N_18678);
nand U21260 (N_21260,N_18003,N_18454);
or U21261 (N_21261,N_18691,N_19414);
nor U21262 (N_21262,N_18323,N_18706);
xnor U21263 (N_21263,N_19087,N_19922);
xor U21264 (N_21264,N_18078,N_19787);
nor U21265 (N_21265,N_19671,N_19374);
and U21266 (N_21266,N_18022,N_19704);
nor U21267 (N_21267,N_18168,N_19299);
nand U21268 (N_21268,N_18178,N_18873);
nor U21269 (N_21269,N_18880,N_19806);
nand U21270 (N_21270,N_19031,N_18857);
xor U21271 (N_21271,N_19749,N_18334);
nor U21272 (N_21272,N_18551,N_18894);
nor U21273 (N_21273,N_19775,N_19332);
xor U21274 (N_21274,N_19372,N_19464);
xnor U21275 (N_21275,N_18424,N_19440);
nand U21276 (N_21276,N_18368,N_19414);
and U21277 (N_21277,N_18077,N_19955);
xor U21278 (N_21278,N_18528,N_18446);
nor U21279 (N_21279,N_18393,N_18161);
and U21280 (N_21280,N_19051,N_18582);
nor U21281 (N_21281,N_19347,N_19267);
and U21282 (N_21282,N_18967,N_18839);
nand U21283 (N_21283,N_18058,N_18423);
and U21284 (N_21284,N_18006,N_19206);
or U21285 (N_21285,N_19802,N_19933);
and U21286 (N_21286,N_18014,N_18621);
or U21287 (N_21287,N_19534,N_19223);
nand U21288 (N_21288,N_19898,N_18878);
and U21289 (N_21289,N_19384,N_19964);
xor U21290 (N_21290,N_19262,N_18637);
and U21291 (N_21291,N_19250,N_19950);
xor U21292 (N_21292,N_19791,N_19885);
xor U21293 (N_21293,N_18606,N_18344);
nor U21294 (N_21294,N_18791,N_18720);
xor U21295 (N_21295,N_19779,N_19296);
xor U21296 (N_21296,N_19395,N_18107);
nor U21297 (N_21297,N_19767,N_18431);
nor U21298 (N_21298,N_18026,N_19656);
nor U21299 (N_21299,N_19201,N_19863);
xor U21300 (N_21300,N_19664,N_18517);
and U21301 (N_21301,N_19023,N_19448);
or U21302 (N_21302,N_19583,N_19212);
and U21303 (N_21303,N_19357,N_18404);
nand U21304 (N_21304,N_19824,N_18262);
and U21305 (N_21305,N_18563,N_18717);
nor U21306 (N_21306,N_18552,N_18537);
nor U21307 (N_21307,N_18305,N_18865);
nand U21308 (N_21308,N_18461,N_19049);
or U21309 (N_21309,N_19952,N_18133);
and U21310 (N_21310,N_18181,N_19975);
or U21311 (N_21311,N_18572,N_19181);
nand U21312 (N_21312,N_18098,N_18034);
nor U21313 (N_21313,N_19228,N_18010);
nand U21314 (N_21314,N_19356,N_19822);
nand U21315 (N_21315,N_18913,N_18482);
nor U21316 (N_21316,N_18266,N_19193);
nand U21317 (N_21317,N_19157,N_19167);
or U21318 (N_21318,N_19228,N_19070);
nand U21319 (N_21319,N_18600,N_18068);
nor U21320 (N_21320,N_18836,N_19785);
xor U21321 (N_21321,N_18821,N_18612);
nand U21322 (N_21322,N_19271,N_19843);
or U21323 (N_21323,N_19723,N_18308);
or U21324 (N_21324,N_19336,N_18854);
and U21325 (N_21325,N_18945,N_18942);
nand U21326 (N_21326,N_18056,N_18073);
or U21327 (N_21327,N_18880,N_18673);
nor U21328 (N_21328,N_19329,N_18814);
or U21329 (N_21329,N_19488,N_19445);
and U21330 (N_21330,N_19669,N_19277);
xor U21331 (N_21331,N_18941,N_18501);
or U21332 (N_21332,N_19973,N_19142);
and U21333 (N_21333,N_19847,N_19923);
nand U21334 (N_21334,N_18881,N_18340);
or U21335 (N_21335,N_19116,N_18543);
and U21336 (N_21336,N_18928,N_18419);
nand U21337 (N_21337,N_18318,N_19395);
and U21338 (N_21338,N_18612,N_18490);
and U21339 (N_21339,N_18102,N_18137);
nand U21340 (N_21340,N_18128,N_18573);
or U21341 (N_21341,N_19167,N_19276);
and U21342 (N_21342,N_18146,N_18229);
nor U21343 (N_21343,N_18477,N_19432);
nand U21344 (N_21344,N_19903,N_18883);
xor U21345 (N_21345,N_18032,N_19525);
nand U21346 (N_21346,N_19841,N_19270);
nor U21347 (N_21347,N_19124,N_18519);
xor U21348 (N_21348,N_18750,N_19221);
nor U21349 (N_21349,N_18984,N_19231);
or U21350 (N_21350,N_18160,N_18312);
and U21351 (N_21351,N_19634,N_19920);
or U21352 (N_21352,N_18772,N_19396);
xnor U21353 (N_21353,N_18899,N_19297);
nand U21354 (N_21354,N_18891,N_19035);
nand U21355 (N_21355,N_18586,N_18595);
nor U21356 (N_21356,N_19580,N_18796);
nand U21357 (N_21357,N_19115,N_18930);
xnor U21358 (N_21358,N_19107,N_19968);
or U21359 (N_21359,N_18571,N_19406);
and U21360 (N_21360,N_18367,N_18195);
or U21361 (N_21361,N_19729,N_19810);
nand U21362 (N_21362,N_19891,N_18438);
nor U21363 (N_21363,N_19657,N_18859);
nand U21364 (N_21364,N_18060,N_19773);
and U21365 (N_21365,N_19272,N_18619);
nand U21366 (N_21366,N_18663,N_19031);
nor U21367 (N_21367,N_18913,N_19172);
or U21368 (N_21368,N_19240,N_19719);
nand U21369 (N_21369,N_18918,N_18792);
nor U21370 (N_21370,N_19048,N_18139);
nor U21371 (N_21371,N_19656,N_19213);
or U21372 (N_21372,N_19967,N_19226);
xnor U21373 (N_21373,N_19881,N_18728);
nand U21374 (N_21374,N_18095,N_18032);
nand U21375 (N_21375,N_19368,N_18262);
and U21376 (N_21376,N_19897,N_19087);
and U21377 (N_21377,N_18873,N_19174);
nand U21378 (N_21378,N_18214,N_19450);
nor U21379 (N_21379,N_19187,N_19473);
nor U21380 (N_21380,N_19280,N_18506);
nand U21381 (N_21381,N_18258,N_18030);
or U21382 (N_21382,N_19624,N_18067);
nand U21383 (N_21383,N_18397,N_19682);
and U21384 (N_21384,N_18974,N_19499);
nand U21385 (N_21385,N_18596,N_19545);
nand U21386 (N_21386,N_19967,N_19668);
and U21387 (N_21387,N_18731,N_18000);
nor U21388 (N_21388,N_19179,N_19822);
nor U21389 (N_21389,N_19323,N_18356);
nor U21390 (N_21390,N_18508,N_19497);
nor U21391 (N_21391,N_19440,N_19188);
and U21392 (N_21392,N_18908,N_18370);
xor U21393 (N_21393,N_19381,N_18051);
or U21394 (N_21394,N_18109,N_19115);
or U21395 (N_21395,N_18065,N_19771);
and U21396 (N_21396,N_19922,N_18040);
nand U21397 (N_21397,N_19657,N_19953);
nor U21398 (N_21398,N_18525,N_19715);
xor U21399 (N_21399,N_19007,N_19124);
and U21400 (N_21400,N_19657,N_19644);
nor U21401 (N_21401,N_19787,N_19709);
xor U21402 (N_21402,N_19207,N_18380);
or U21403 (N_21403,N_18008,N_19076);
nor U21404 (N_21404,N_18520,N_19383);
xnor U21405 (N_21405,N_18676,N_19971);
and U21406 (N_21406,N_19638,N_18159);
nor U21407 (N_21407,N_19394,N_19112);
nand U21408 (N_21408,N_19980,N_18372);
and U21409 (N_21409,N_19909,N_19770);
nand U21410 (N_21410,N_19548,N_18836);
nor U21411 (N_21411,N_19877,N_19375);
and U21412 (N_21412,N_18622,N_18249);
nand U21413 (N_21413,N_18340,N_18573);
xor U21414 (N_21414,N_18866,N_19051);
xnor U21415 (N_21415,N_18389,N_19435);
xor U21416 (N_21416,N_18963,N_18340);
nand U21417 (N_21417,N_19769,N_19272);
or U21418 (N_21418,N_18420,N_19656);
and U21419 (N_21419,N_18042,N_19491);
nand U21420 (N_21420,N_18651,N_18351);
nor U21421 (N_21421,N_18704,N_18000);
nor U21422 (N_21422,N_19972,N_18649);
and U21423 (N_21423,N_18961,N_19333);
and U21424 (N_21424,N_19259,N_18917);
nor U21425 (N_21425,N_19493,N_19342);
and U21426 (N_21426,N_18337,N_19047);
xor U21427 (N_21427,N_19329,N_19038);
or U21428 (N_21428,N_19689,N_18406);
or U21429 (N_21429,N_19501,N_19124);
xor U21430 (N_21430,N_19352,N_19013);
or U21431 (N_21431,N_18212,N_18325);
nor U21432 (N_21432,N_18424,N_19674);
nand U21433 (N_21433,N_19006,N_19353);
nor U21434 (N_21434,N_19653,N_19384);
and U21435 (N_21435,N_19755,N_18031);
xnor U21436 (N_21436,N_18666,N_18033);
xnor U21437 (N_21437,N_19797,N_19763);
and U21438 (N_21438,N_18321,N_18484);
or U21439 (N_21439,N_18114,N_18211);
or U21440 (N_21440,N_18824,N_19655);
xor U21441 (N_21441,N_19771,N_18555);
nor U21442 (N_21442,N_18538,N_18745);
or U21443 (N_21443,N_18211,N_18909);
and U21444 (N_21444,N_19583,N_19747);
and U21445 (N_21445,N_18221,N_18176);
nor U21446 (N_21446,N_18931,N_18755);
nor U21447 (N_21447,N_19245,N_19546);
and U21448 (N_21448,N_18231,N_19575);
xor U21449 (N_21449,N_19610,N_19102);
or U21450 (N_21450,N_18719,N_18286);
and U21451 (N_21451,N_19593,N_18374);
and U21452 (N_21452,N_18199,N_19948);
and U21453 (N_21453,N_19021,N_19354);
xnor U21454 (N_21454,N_19952,N_18371);
xor U21455 (N_21455,N_19696,N_18517);
and U21456 (N_21456,N_19771,N_19592);
nand U21457 (N_21457,N_19648,N_18799);
or U21458 (N_21458,N_18894,N_18603);
xnor U21459 (N_21459,N_18766,N_19650);
xor U21460 (N_21460,N_19073,N_18597);
or U21461 (N_21461,N_19831,N_18440);
xnor U21462 (N_21462,N_19185,N_19517);
nand U21463 (N_21463,N_19807,N_18250);
and U21464 (N_21464,N_19841,N_18674);
nand U21465 (N_21465,N_18558,N_19778);
nor U21466 (N_21466,N_18196,N_19198);
nand U21467 (N_21467,N_18874,N_18408);
or U21468 (N_21468,N_18886,N_18803);
nand U21469 (N_21469,N_18746,N_18726);
xor U21470 (N_21470,N_19540,N_19296);
nor U21471 (N_21471,N_18593,N_18162);
or U21472 (N_21472,N_19813,N_18602);
and U21473 (N_21473,N_18679,N_18887);
nor U21474 (N_21474,N_18579,N_18953);
and U21475 (N_21475,N_18660,N_18953);
nand U21476 (N_21476,N_19758,N_18478);
nor U21477 (N_21477,N_19529,N_19494);
nor U21478 (N_21478,N_18412,N_19832);
or U21479 (N_21479,N_18788,N_18308);
xor U21480 (N_21480,N_19659,N_19297);
nand U21481 (N_21481,N_18990,N_18740);
and U21482 (N_21482,N_18928,N_19467);
and U21483 (N_21483,N_18896,N_18716);
or U21484 (N_21484,N_19777,N_18374);
or U21485 (N_21485,N_18199,N_19853);
nand U21486 (N_21486,N_19428,N_19307);
and U21487 (N_21487,N_18758,N_19467);
and U21488 (N_21488,N_18645,N_19867);
xor U21489 (N_21489,N_19932,N_18536);
xnor U21490 (N_21490,N_19378,N_19041);
nand U21491 (N_21491,N_18044,N_18238);
xor U21492 (N_21492,N_19389,N_19287);
or U21493 (N_21493,N_19733,N_18317);
xnor U21494 (N_21494,N_18444,N_18810);
nand U21495 (N_21495,N_19551,N_19579);
and U21496 (N_21496,N_18566,N_19286);
and U21497 (N_21497,N_19496,N_19798);
nand U21498 (N_21498,N_18774,N_19170);
nor U21499 (N_21499,N_18303,N_18020);
and U21500 (N_21500,N_19167,N_19388);
nand U21501 (N_21501,N_18561,N_18339);
or U21502 (N_21502,N_19454,N_18104);
or U21503 (N_21503,N_19987,N_18363);
and U21504 (N_21504,N_19430,N_18426);
xor U21505 (N_21505,N_18148,N_19601);
xor U21506 (N_21506,N_19752,N_18441);
and U21507 (N_21507,N_19854,N_18145);
xnor U21508 (N_21508,N_19052,N_19798);
xor U21509 (N_21509,N_18057,N_19054);
xnor U21510 (N_21510,N_19824,N_19701);
or U21511 (N_21511,N_19723,N_19102);
or U21512 (N_21512,N_18164,N_18369);
nand U21513 (N_21513,N_19924,N_18053);
xnor U21514 (N_21514,N_19428,N_19368);
nor U21515 (N_21515,N_18068,N_18039);
nor U21516 (N_21516,N_19668,N_18022);
xnor U21517 (N_21517,N_19234,N_18029);
nor U21518 (N_21518,N_18677,N_19937);
xor U21519 (N_21519,N_18037,N_18531);
or U21520 (N_21520,N_19210,N_19871);
or U21521 (N_21521,N_19340,N_18528);
or U21522 (N_21522,N_18656,N_19145);
nand U21523 (N_21523,N_18309,N_19852);
or U21524 (N_21524,N_19937,N_18923);
nor U21525 (N_21525,N_19184,N_19422);
nand U21526 (N_21526,N_19293,N_18543);
nand U21527 (N_21527,N_18278,N_18288);
xor U21528 (N_21528,N_19894,N_18956);
xor U21529 (N_21529,N_18225,N_18468);
nand U21530 (N_21530,N_18176,N_18534);
nand U21531 (N_21531,N_18588,N_19592);
xnor U21532 (N_21532,N_18705,N_19012);
nand U21533 (N_21533,N_19220,N_18805);
or U21534 (N_21534,N_19399,N_19913);
nand U21535 (N_21535,N_18411,N_19011);
and U21536 (N_21536,N_19722,N_19658);
xor U21537 (N_21537,N_18631,N_19689);
nor U21538 (N_21538,N_19263,N_19808);
nor U21539 (N_21539,N_19114,N_18781);
and U21540 (N_21540,N_19781,N_19445);
nor U21541 (N_21541,N_18462,N_18273);
nand U21542 (N_21542,N_18873,N_19095);
or U21543 (N_21543,N_18961,N_18905);
xor U21544 (N_21544,N_19348,N_19850);
nand U21545 (N_21545,N_19646,N_19285);
nor U21546 (N_21546,N_19177,N_18512);
nor U21547 (N_21547,N_18253,N_19127);
and U21548 (N_21548,N_19758,N_18897);
nand U21549 (N_21549,N_18843,N_19198);
nor U21550 (N_21550,N_18851,N_19877);
and U21551 (N_21551,N_19202,N_18030);
nor U21552 (N_21552,N_19149,N_19723);
and U21553 (N_21553,N_19634,N_19242);
or U21554 (N_21554,N_19516,N_19818);
and U21555 (N_21555,N_19528,N_19095);
nand U21556 (N_21556,N_18825,N_19785);
nor U21557 (N_21557,N_19874,N_19310);
nand U21558 (N_21558,N_19580,N_18137);
xnor U21559 (N_21559,N_19462,N_19876);
nor U21560 (N_21560,N_19539,N_18965);
nand U21561 (N_21561,N_19836,N_19006);
or U21562 (N_21562,N_19963,N_19832);
nor U21563 (N_21563,N_19553,N_19611);
or U21564 (N_21564,N_18948,N_18899);
nor U21565 (N_21565,N_18098,N_18955);
nor U21566 (N_21566,N_18659,N_18775);
xnor U21567 (N_21567,N_18390,N_19124);
and U21568 (N_21568,N_19802,N_18969);
or U21569 (N_21569,N_19985,N_19867);
and U21570 (N_21570,N_19474,N_19938);
xnor U21571 (N_21571,N_18212,N_18973);
and U21572 (N_21572,N_19257,N_18310);
xor U21573 (N_21573,N_19559,N_18657);
or U21574 (N_21574,N_18579,N_19193);
nor U21575 (N_21575,N_19133,N_19046);
nor U21576 (N_21576,N_19256,N_19973);
or U21577 (N_21577,N_19368,N_18733);
and U21578 (N_21578,N_18711,N_18470);
and U21579 (N_21579,N_18192,N_19109);
or U21580 (N_21580,N_19262,N_19041);
and U21581 (N_21581,N_19325,N_18209);
nand U21582 (N_21582,N_18110,N_18835);
nor U21583 (N_21583,N_19993,N_18463);
nand U21584 (N_21584,N_18987,N_19145);
and U21585 (N_21585,N_18657,N_18686);
or U21586 (N_21586,N_19748,N_19908);
and U21587 (N_21587,N_18182,N_19162);
xnor U21588 (N_21588,N_19516,N_19465);
and U21589 (N_21589,N_18383,N_19270);
xnor U21590 (N_21590,N_19581,N_19683);
or U21591 (N_21591,N_18569,N_19891);
and U21592 (N_21592,N_18568,N_18884);
and U21593 (N_21593,N_19035,N_18316);
nand U21594 (N_21594,N_18858,N_19368);
xor U21595 (N_21595,N_19757,N_19137);
xnor U21596 (N_21596,N_18853,N_19597);
xnor U21597 (N_21597,N_18413,N_19141);
and U21598 (N_21598,N_18255,N_19797);
or U21599 (N_21599,N_18095,N_18989);
xor U21600 (N_21600,N_19896,N_19571);
nor U21601 (N_21601,N_19393,N_19425);
nand U21602 (N_21602,N_19550,N_18490);
and U21603 (N_21603,N_19051,N_19717);
or U21604 (N_21604,N_18663,N_18265);
or U21605 (N_21605,N_19244,N_19526);
or U21606 (N_21606,N_19764,N_19762);
xnor U21607 (N_21607,N_18608,N_18347);
and U21608 (N_21608,N_19272,N_19839);
nand U21609 (N_21609,N_18290,N_18632);
nor U21610 (N_21610,N_19637,N_19915);
and U21611 (N_21611,N_19899,N_18130);
nor U21612 (N_21612,N_18438,N_18546);
or U21613 (N_21613,N_19382,N_19021);
nand U21614 (N_21614,N_18348,N_18684);
and U21615 (N_21615,N_18944,N_19654);
nor U21616 (N_21616,N_19472,N_19498);
and U21617 (N_21617,N_19777,N_19861);
and U21618 (N_21618,N_19446,N_19310);
or U21619 (N_21619,N_19398,N_19093);
nand U21620 (N_21620,N_19374,N_19560);
xor U21621 (N_21621,N_18119,N_19313);
and U21622 (N_21622,N_19947,N_19689);
nor U21623 (N_21623,N_18423,N_18612);
and U21624 (N_21624,N_18045,N_18358);
nor U21625 (N_21625,N_18544,N_18297);
nand U21626 (N_21626,N_19592,N_19689);
xnor U21627 (N_21627,N_18108,N_18579);
xnor U21628 (N_21628,N_19196,N_19945);
nand U21629 (N_21629,N_19039,N_18240);
or U21630 (N_21630,N_19223,N_19025);
or U21631 (N_21631,N_18992,N_19255);
xnor U21632 (N_21632,N_19359,N_18580);
xor U21633 (N_21633,N_18445,N_19080);
xor U21634 (N_21634,N_19133,N_18719);
and U21635 (N_21635,N_18176,N_19473);
and U21636 (N_21636,N_18625,N_19071);
and U21637 (N_21637,N_19637,N_19615);
xor U21638 (N_21638,N_19720,N_19889);
nor U21639 (N_21639,N_18922,N_18843);
and U21640 (N_21640,N_18410,N_18096);
and U21641 (N_21641,N_18974,N_18961);
xor U21642 (N_21642,N_19929,N_18096);
nor U21643 (N_21643,N_19159,N_19681);
or U21644 (N_21644,N_18647,N_18821);
nor U21645 (N_21645,N_18980,N_19055);
xnor U21646 (N_21646,N_18739,N_19716);
xnor U21647 (N_21647,N_19625,N_18913);
nor U21648 (N_21648,N_18458,N_19222);
or U21649 (N_21649,N_18552,N_19222);
nor U21650 (N_21650,N_19863,N_18904);
or U21651 (N_21651,N_18911,N_18536);
or U21652 (N_21652,N_19554,N_19822);
and U21653 (N_21653,N_18522,N_19194);
and U21654 (N_21654,N_19694,N_19936);
xnor U21655 (N_21655,N_18948,N_19735);
nor U21656 (N_21656,N_18627,N_18355);
or U21657 (N_21657,N_19393,N_19787);
nor U21658 (N_21658,N_19924,N_18963);
or U21659 (N_21659,N_19054,N_19103);
or U21660 (N_21660,N_18206,N_19441);
nand U21661 (N_21661,N_18792,N_19705);
xor U21662 (N_21662,N_19767,N_18649);
nor U21663 (N_21663,N_19364,N_19524);
xnor U21664 (N_21664,N_19160,N_19773);
nand U21665 (N_21665,N_19324,N_18062);
or U21666 (N_21666,N_19477,N_19717);
nand U21667 (N_21667,N_18786,N_18340);
or U21668 (N_21668,N_19340,N_19935);
nand U21669 (N_21669,N_19234,N_18148);
nand U21670 (N_21670,N_18840,N_18619);
nor U21671 (N_21671,N_18109,N_19474);
and U21672 (N_21672,N_18154,N_18380);
nor U21673 (N_21673,N_19509,N_18118);
and U21674 (N_21674,N_19828,N_18726);
or U21675 (N_21675,N_19783,N_19727);
nor U21676 (N_21676,N_18198,N_18133);
and U21677 (N_21677,N_18389,N_18228);
and U21678 (N_21678,N_19443,N_19181);
nand U21679 (N_21679,N_19375,N_18195);
or U21680 (N_21680,N_19530,N_19368);
or U21681 (N_21681,N_18103,N_18241);
or U21682 (N_21682,N_18078,N_18526);
and U21683 (N_21683,N_18815,N_19199);
nand U21684 (N_21684,N_18546,N_19294);
and U21685 (N_21685,N_18095,N_18446);
and U21686 (N_21686,N_19859,N_18474);
nand U21687 (N_21687,N_18097,N_18898);
and U21688 (N_21688,N_18578,N_19236);
nand U21689 (N_21689,N_19590,N_19206);
or U21690 (N_21690,N_18526,N_19391);
and U21691 (N_21691,N_18411,N_18698);
or U21692 (N_21692,N_18396,N_18345);
nand U21693 (N_21693,N_18796,N_19976);
or U21694 (N_21694,N_19669,N_19413);
or U21695 (N_21695,N_18613,N_19153);
and U21696 (N_21696,N_19073,N_19764);
nand U21697 (N_21697,N_18875,N_19794);
nor U21698 (N_21698,N_19459,N_19580);
and U21699 (N_21699,N_18073,N_19536);
nor U21700 (N_21700,N_19302,N_18395);
and U21701 (N_21701,N_18836,N_18949);
and U21702 (N_21702,N_19009,N_19844);
nand U21703 (N_21703,N_19324,N_19017);
nor U21704 (N_21704,N_18094,N_19353);
nor U21705 (N_21705,N_18292,N_18764);
xor U21706 (N_21706,N_18319,N_18617);
nor U21707 (N_21707,N_18371,N_18213);
or U21708 (N_21708,N_19120,N_19993);
xor U21709 (N_21709,N_19611,N_18293);
nand U21710 (N_21710,N_18098,N_18870);
nand U21711 (N_21711,N_19201,N_18619);
and U21712 (N_21712,N_19971,N_18113);
nand U21713 (N_21713,N_18664,N_18029);
or U21714 (N_21714,N_18215,N_18736);
nand U21715 (N_21715,N_18574,N_18357);
nand U21716 (N_21716,N_19940,N_19964);
nand U21717 (N_21717,N_18511,N_18836);
nor U21718 (N_21718,N_19173,N_18711);
nand U21719 (N_21719,N_18098,N_18656);
and U21720 (N_21720,N_18836,N_19858);
and U21721 (N_21721,N_18068,N_18843);
or U21722 (N_21722,N_19359,N_18000);
and U21723 (N_21723,N_18038,N_18865);
nor U21724 (N_21724,N_19925,N_19896);
nor U21725 (N_21725,N_18775,N_19593);
xor U21726 (N_21726,N_19183,N_18120);
xor U21727 (N_21727,N_18860,N_19789);
nand U21728 (N_21728,N_19262,N_19074);
nor U21729 (N_21729,N_18406,N_19158);
nor U21730 (N_21730,N_19517,N_19927);
nand U21731 (N_21731,N_19679,N_18830);
xor U21732 (N_21732,N_18664,N_19407);
and U21733 (N_21733,N_18505,N_18660);
and U21734 (N_21734,N_19311,N_19975);
xnor U21735 (N_21735,N_19058,N_18468);
nor U21736 (N_21736,N_18978,N_19107);
nand U21737 (N_21737,N_18227,N_19004);
xor U21738 (N_21738,N_19826,N_18366);
nand U21739 (N_21739,N_19983,N_18125);
nor U21740 (N_21740,N_18407,N_18007);
or U21741 (N_21741,N_18048,N_19343);
and U21742 (N_21742,N_19388,N_19826);
nand U21743 (N_21743,N_19918,N_19459);
xor U21744 (N_21744,N_18100,N_19328);
xor U21745 (N_21745,N_18956,N_18029);
or U21746 (N_21746,N_18948,N_18481);
xor U21747 (N_21747,N_19036,N_18247);
or U21748 (N_21748,N_19172,N_18322);
nand U21749 (N_21749,N_18928,N_19773);
and U21750 (N_21750,N_18397,N_18553);
nor U21751 (N_21751,N_19789,N_19044);
nor U21752 (N_21752,N_19139,N_18012);
nand U21753 (N_21753,N_19065,N_19194);
xnor U21754 (N_21754,N_18245,N_19933);
xnor U21755 (N_21755,N_19829,N_19962);
xnor U21756 (N_21756,N_18476,N_18640);
nor U21757 (N_21757,N_19966,N_19502);
xor U21758 (N_21758,N_19603,N_18026);
xnor U21759 (N_21759,N_18687,N_18092);
xnor U21760 (N_21760,N_18761,N_18499);
and U21761 (N_21761,N_18527,N_18735);
and U21762 (N_21762,N_19413,N_19150);
nor U21763 (N_21763,N_19985,N_18782);
and U21764 (N_21764,N_19391,N_18226);
nand U21765 (N_21765,N_19517,N_18925);
xnor U21766 (N_21766,N_19408,N_18906);
nor U21767 (N_21767,N_18294,N_18950);
nor U21768 (N_21768,N_18943,N_18126);
xor U21769 (N_21769,N_18640,N_18357);
and U21770 (N_21770,N_19398,N_18040);
and U21771 (N_21771,N_18951,N_18224);
nand U21772 (N_21772,N_19074,N_18784);
xnor U21773 (N_21773,N_18693,N_18198);
xnor U21774 (N_21774,N_18959,N_18400);
xnor U21775 (N_21775,N_19092,N_19669);
or U21776 (N_21776,N_19994,N_19670);
xor U21777 (N_21777,N_19064,N_19525);
nor U21778 (N_21778,N_19770,N_18141);
or U21779 (N_21779,N_18623,N_18294);
and U21780 (N_21780,N_18222,N_18071);
nor U21781 (N_21781,N_18109,N_18570);
or U21782 (N_21782,N_18262,N_18109);
nand U21783 (N_21783,N_19904,N_18986);
nand U21784 (N_21784,N_18817,N_19357);
or U21785 (N_21785,N_18009,N_18761);
xnor U21786 (N_21786,N_19298,N_18222);
and U21787 (N_21787,N_19837,N_19865);
nor U21788 (N_21788,N_19446,N_19991);
or U21789 (N_21789,N_18424,N_18280);
xor U21790 (N_21790,N_18883,N_19866);
xnor U21791 (N_21791,N_19372,N_18241);
nor U21792 (N_21792,N_18178,N_18008);
nor U21793 (N_21793,N_18902,N_18372);
xnor U21794 (N_21794,N_18195,N_18293);
xor U21795 (N_21795,N_18262,N_18157);
or U21796 (N_21796,N_19736,N_19744);
xnor U21797 (N_21797,N_19166,N_19748);
xor U21798 (N_21798,N_19967,N_18983);
and U21799 (N_21799,N_18018,N_18205);
xor U21800 (N_21800,N_18291,N_18749);
or U21801 (N_21801,N_18577,N_19845);
nor U21802 (N_21802,N_19744,N_19968);
and U21803 (N_21803,N_18307,N_19728);
and U21804 (N_21804,N_19458,N_19304);
nor U21805 (N_21805,N_18651,N_19178);
nand U21806 (N_21806,N_19459,N_19922);
nand U21807 (N_21807,N_19507,N_19443);
nor U21808 (N_21808,N_18009,N_18427);
nand U21809 (N_21809,N_19541,N_19087);
and U21810 (N_21810,N_18900,N_19415);
nor U21811 (N_21811,N_19313,N_18277);
and U21812 (N_21812,N_19195,N_19833);
or U21813 (N_21813,N_19531,N_18324);
nand U21814 (N_21814,N_18205,N_19449);
nand U21815 (N_21815,N_19156,N_19866);
nand U21816 (N_21816,N_19021,N_19074);
nand U21817 (N_21817,N_19226,N_19314);
xnor U21818 (N_21818,N_19262,N_19058);
nor U21819 (N_21819,N_18261,N_19856);
nor U21820 (N_21820,N_19787,N_19916);
nand U21821 (N_21821,N_18838,N_18542);
nand U21822 (N_21822,N_18203,N_18202);
nor U21823 (N_21823,N_18456,N_18604);
or U21824 (N_21824,N_19088,N_19045);
xor U21825 (N_21825,N_19398,N_18011);
or U21826 (N_21826,N_18782,N_19241);
and U21827 (N_21827,N_18200,N_19343);
xnor U21828 (N_21828,N_18245,N_18184);
nor U21829 (N_21829,N_18430,N_19508);
xor U21830 (N_21830,N_18406,N_19191);
or U21831 (N_21831,N_19735,N_19884);
xnor U21832 (N_21832,N_19455,N_19313);
xnor U21833 (N_21833,N_18319,N_19895);
and U21834 (N_21834,N_18045,N_18927);
or U21835 (N_21835,N_18691,N_18659);
and U21836 (N_21836,N_19127,N_19121);
nor U21837 (N_21837,N_18039,N_18022);
or U21838 (N_21838,N_18962,N_19209);
xnor U21839 (N_21839,N_18514,N_18607);
nand U21840 (N_21840,N_18176,N_18557);
xor U21841 (N_21841,N_18307,N_19666);
or U21842 (N_21842,N_19032,N_19283);
or U21843 (N_21843,N_19982,N_18570);
nand U21844 (N_21844,N_19551,N_18062);
nand U21845 (N_21845,N_19624,N_19326);
xor U21846 (N_21846,N_19104,N_19619);
and U21847 (N_21847,N_18499,N_18831);
xor U21848 (N_21848,N_18684,N_19450);
or U21849 (N_21849,N_19489,N_19606);
and U21850 (N_21850,N_19310,N_18728);
nor U21851 (N_21851,N_19976,N_18139);
or U21852 (N_21852,N_18322,N_18602);
nor U21853 (N_21853,N_18575,N_19522);
or U21854 (N_21854,N_19367,N_18559);
and U21855 (N_21855,N_18973,N_18396);
nand U21856 (N_21856,N_19536,N_19253);
or U21857 (N_21857,N_19557,N_19504);
nand U21858 (N_21858,N_18331,N_19686);
and U21859 (N_21859,N_18013,N_18072);
nor U21860 (N_21860,N_18511,N_19268);
xnor U21861 (N_21861,N_18747,N_18269);
or U21862 (N_21862,N_19541,N_18803);
or U21863 (N_21863,N_18423,N_18888);
or U21864 (N_21864,N_19723,N_19764);
nand U21865 (N_21865,N_18058,N_19212);
xnor U21866 (N_21866,N_19746,N_19779);
xor U21867 (N_21867,N_19414,N_18060);
nand U21868 (N_21868,N_18078,N_19208);
nand U21869 (N_21869,N_18784,N_19211);
nand U21870 (N_21870,N_19514,N_18807);
xor U21871 (N_21871,N_19995,N_19009);
nor U21872 (N_21872,N_18207,N_18483);
or U21873 (N_21873,N_18681,N_19926);
and U21874 (N_21874,N_18479,N_18710);
or U21875 (N_21875,N_18638,N_18837);
xnor U21876 (N_21876,N_18321,N_19057);
nor U21877 (N_21877,N_18453,N_18761);
nand U21878 (N_21878,N_19474,N_18951);
nor U21879 (N_21879,N_18874,N_19592);
or U21880 (N_21880,N_18898,N_18418);
or U21881 (N_21881,N_19124,N_18253);
or U21882 (N_21882,N_19763,N_18944);
and U21883 (N_21883,N_18782,N_19725);
and U21884 (N_21884,N_19016,N_18028);
and U21885 (N_21885,N_18985,N_18950);
nand U21886 (N_21886,N_19037,N_18339);
nor U21887 (N_21887,N_18754,N_19456);
and U21888 (N_21888,N_19180,N_18814);
or U21889 (N_21889,N_19004,N_19904);
and U21890 (N_21890,N_18747,N_18590);
nand U21891 (N_21891,N_18328,N_18195);
and U21892 (N_21892,N_19954,N_18408);
and U21893 (N_21893,N_18405,N_18134);
nand U21894 (N_21894,N_19885,N_18660);
or U21895 (N_21895,N_18490,N_18739);
or U21896 (N_21896,N_19689,N_19067);
or U21897 (N_21897,N_19263,N_18741);
nand U21898 (N_21898,N_19932,N_18882);
nand U21899 (N_21899,N_18824,N_18888);
nor U21900 (N_21900,N_19719,N_19921);
xor U21901 (N_21901,N_18355,N_18580);
and U21902 (N_21902,N_18907,N_19165);
nor U21903 (N_21903,N_18400,N_19646);
nand U21904 (N_21904,N_18744,N_19638);
or U21905 (N_21905,N_18053,N_19431);
or U21906 (N_21906,N_18648,N_19676);
or U21907 (N_21907,N_18217,N_19960);
nor U21908 (N_21908,N_18054,N_19673);
xor U21909 (N_21909,N_18684,N_18772);
nor U21910 (N_21910,N_18169,N_18868);
nor U21911 (N_21911,N_19501,N_18490);
and U21912 (N_21912,N_19305,N_18153);
nor U21913 (N_21913,N_18825,N_19847);
nand U21914 (N_21914,N_19578,N_18302);
or U21915 (N_21915,N_19145,N_18078);
nand U21916 (N_21916,N_18072,N_19045);
or U21917 (N_21917,N_19252,N_18271);
and U21918 (N_21918,N_18376,N_19474);
xnor U21919 (N_21919,N_18823,N_18035);
nor U21920 (N_21920,N_19101,N_18621);
nor U21921 (N_21921,N_18005,N_19448);
and U21922 (N_21922,N_18488,N_18985);
nand U21923 (N_21923,N_18838,N_19709);
nand U21924 (N_21924,N_18163,N_18506);
nand U21925 (N_21925,N_19592,N_18065);
xnor U21926 (N_21926,N_18261,N_19115);
xor U21927 (N_21927,N_18912,N_18471);
xor U21928 (N_21928,N_18821,N_18257);
or U21929 (N_21929,N_18408,N_19195);
or U21930 (N_21930,N_19478,N_19538);
nand U21931 (N_21931,N_19567,N_18387);
nand U21932 (N_21932,N_18413,N_19688);
xor U21933 (N_21933,N_18236,N_19330);
and U21934 (N_21934,N_18314,N_19783);
nand U21935 (N_21935,N_19720,N_18592);
or U21936 (N_21936,N_18372,N_19844);
nand U21937 (N_21937,N_19953,N_18794);
or U21938 (N_21938,N_19396,N_18587);
nor U21939 (N_21939,N_19248,N_18618);
xnor U21940 (N_21940,N_19711,N_19295);
xnor U21941 (N_21941,N_19981,N_18570);
or U21942 (N_21942,N_18066,N_19697);
nor U21943 (N_21943,N_18046,N_19765);
and U21944 (N_21944,N_19127,N_18819);
or U21945 (N_21945,N_19648,N_18396);
or U21946 (N_21946,N_18168,N_19237);
xor U21947 (N_21947,N_18321,N_19782);
nand U21948 (N_21948,N_18498,N_19578);
xor U21949 (N_21949,N_18256,N_18290);
xnor U21950 (N_21950,N_18018,N_19406);
nand U21951 (N_21951,N_18654,N_18599);
xnor U21952 (N_21952,N_19449,N_18181);
nand U21953 (N_21953,N_19239,N_18358);
or U21954 (N_21954,N_19031,N_18650);
and U21955 (N_21955,N_19493,N_18317);
and U21956 (N_21956,N_18370,N_19537);
nor U21957 (N_21957,N_18602,N_19733);
xnor U21958 (N_21958,N_19987,N_19849);
and U21959 (N_21959,N_19887,N_18012);
and U21960 (N_21960,N_18249,N_19149);
nor U21961 (N_21961,N_19092,N_18516);
and U21962 (N_21962,N_18053,N_18086);
nand U21963 (N_21963,N_19310,N_19423);
nand U21964 (N_21964,N_19384,N_19164);
or U21965 (N_21965,N_18662,N_18089);
and U21966 (N_21966,N_19753,N_18682);
xnor U21967 (N_21967,N_19370,N_18065);
or U21968 (N_21968,N_19742,N_18244);
nor U21969 (N_21969,N_19576,N_19543);
nor U21970 (N_21970,N_18182,N_18478);
or U21971 (N_21971,N_19620,N_18201);
and U21972 (N_21972,N_19136,N_19432);
nor U21973 (N_21973,N_18264,N_19855);
nand U21974 (N_21974,N_19166,N_19495);
nand U21975 (N_21975,N_18972,N_18908);
nand U21976 (N_21976,N_18400,N_19023);
or U21977 (N_21977,N_18131,N_19932);
nor U21978 (N_21978,N_18167,N_18051);
nor U21979 (N_21979,N_19057,N_18777);
nor U21980 (N_21980,N_19151,N_18486);
or U21981 (N_21981,N_18316,N_18149);
nor U21982 (N_21982,N_19437,N_19056);
and U21983 (N_21983,N_18418,N_18338);
nand U21984 (N_21984,N_19684,N_19029);
nor U21985 (N_21985,N_19534,N_18551);
nor U21986 (N_21986,N_18158,N_18890);
nor U21987 (N_21987,N_19395,N_18776);
or U21988 (N_21988,N_18818,N_18098);
nor U21989 (N_21989,N_19673,N_18681);
nand U21990 (N_21990,N_19782,N_18364);
and U21991 (N_21991,N_19857,N_18482);
nor U21992 (N_21992,N_18085,N_19071);
or U21993 (N_21993,N_19049,N_19951);
or U21994 (N_21994,N_18054,N_19304);
nand U21995 (N_21995,N_18002,N_19960);
xnor U21996 (N_21996,N_18638,N_19919);
or U21997 (N_21997,N_19538,N_19868);
nand U21998 (N_21998,N_18050,N_19580);
and U21999 (N_21999,N_19421,N_19285);
nor U22000 (N_22000,N_20348,N_21724);
or U22001 (N_22001,N_21068,N_21164);
xnor U22002 (N_22002,N_21761,N_20685);
nor U22003 (N_22003,N_20535,N_21389);
nand U22004 (N_22004,N_20566,N_20222);
xnor U22005 (N_22005,N_21790,N_21643);
nand U22006 (N_22006,N_21634,N_21515);
or U22007 (N_22007,N_21813,N_21689);
and U22008 (N_22008,N_21929,N_20882);
or U22009 (N_22009,N_20610,N_21808);
and U22010 (N_22010,N_21949,N_21685);
and U22011 (N_22011,N_21045,N_21655);
xor U22012 (N_22012,N_20463,N_20925);
nand U22013 (N_22013,N_20819,N_21607);
xor U22014 (N_22014,N_20241,N_21955);
xor U22015 (N_22015,N_20868,N_21281);
or U22016 (N_22016,N_20103,N_21134);
nor U22017 (N_22017,N_20788,N_20702);
and U22018 (N_22018,N_20741,N_21639);
and U22019 (N_22019,N_20804,N_21222);
and U22020 (N_22020,N_20444,N_20753);
nand U22021 (N_22021,N_21087,N_20714);
or U22022 (N_22022,N_20299,N_20924);
nand U22023 (N_22023,N_20305,N_20791);
or U22024 (N_22024,N_21044,N_20235);
or U22025 (N_22025,N_21997,N_21844);
xor U22026 (N_22026,N_21492,N_20242);
nor U22027 (N_22027,N_21864,N_20149);
nor U22028 (N_22028,N_20856,N_20887);
nor U22029 (N_22029,N_20273,N_20757);
or U22030 (N_22030,N_21065,N_21106);
and U22031 (N_22031,N_20328,N_21230);
nand U22032 (N_22032,N_20018,N_21172);
nor U22033 (N_22033,N_21443,N_21446);
or U22034 (N_22034,N_20154,N_20064);
or U22035 (N_22035,N_21345,N_21952);
and U22036 (N_22036,N_20072,N_21484);
or U22037 (N_22037,N_20891,N_21425);
and U22038 (N_22038,N_21283,N_20632);
xor U22039 (N_22039,N_20198,N_21616);
nand U22040 (N_22040,N_20717,N_20726);
and U22041 (N_22041,N_21200,N_21647);
and U22042 (N_22042,N_21941,N_21290);
nor U22043 (N_22043,N_21921,N_20545);
and U22044 (N_22044,N_20326,N_20023);
or U22045 (N_22045,N_21462,N_21510);
and U22046 (N_22046,N_20906,N_21973);
nor U22047 (N_22047,N_20031,N_21171);
xor U22048 (N_22048,N_21173,N_21573);
and U22049 (N_22049,N_21898,N_20596);
xnor U22050 (N_22050,N_21037,N_20503);
xnor U22051 (N_22051,N_20544,N_20042);
nor U22052 (N_22052,N_21207,N_21104);
and U22053 (N_22053,N_21827,N_20773);
nand U22054 (N_22054,N_21320,N_20622);
or U22055 (N_22055,N_21879,N_20693);
nand U22056 (N_22056,N_21257,N_21801);
xnor U22057 (N_22057,N_21971,N_21012);
xnor U22058 (N_22058,N_21220,N_20938);
and U22059 (N_22059,N_21474,N_21985);
nor U22060 (N_22060,N_21742,N_20079);
nor U22061 (N_22061,N_20357,N_21174);
or U22062 (N_22062,N_20621,N_21215);
nand U22063 (N_22063,N_21025,N_20703);
xnor U22064 (N_22064,N_20441,N_20514);
nor U22065 (N_22065,N_21185,N_20112);
or U22066 (N_22066,N_21007,N_20433);
or U22067 (N_22067,N_20897,N_20419);
and U22068 (N_22068,N_21533,N_21935);
xnor U22069 (N_22069,N_20795,N_21888);
nor U22070 (N_22070,N_20571,N_20518);
and U22071 (N_22071,N_21271,N_20803);
xor U22072 (N_22072,N_20495,N_21505);
and U22073 (N_22073,N_20155,N_21361);
or U22074 (N_22074,N_21706,N_20105);
or U22075 (N_22075,N_21204,N_20866);
and U22076 (N_22076,N_21386,N_21117);
xnor U22077 (N_22077,N_20949,N_20705);
nand U22078 (N_22078,N_20044,N_20336);
nor U22079 (N_22079,N_20618,N_20003);
nor U22080 (N_22080,N_20076,N_21370);
xnor U22081 (N_22081,N_21487,N_20979);
xor U22082 (N_22082,N_21429,N_21521);
nand U22083 (N_22083,N_20740,N_21556);
or U22084 (N_22084,N_21940,N_21748);
nand U22085 (N_22085,N_21181,N_20434);
nor U22086 (N_22086,N_20821,N_20500);
nor U22087 (N_22087,N_21870,N_20229);
xnor U22088 (N_22088,N_21658,N_21800);
nor U22089 (N_22089,N_21455,N_21795);
nor U22090 (N_22090,N_21463,N_20701);
and U22091 (N_22091,N_20339,N_21555);
nor U22092 (N_22092,N_21031,N_21956);
xnor U22093 (N_22093,N_20369,N_20333);
xor U22094 (N_22094,N_21387,N_21757);
and U22095 (N_22095,N_20853,N_21596);
xor U22096 (N_22096,N_21401,N_21278);
nand U22097 (N_22097,N_20613,N_21632);
and U22098 (N_22098,N_20445,N_21415);
or U22099 (N_22099,N_21873,N_21541);
nor U22100 (N_22100,N_21201,N_21237);
or U22101 (N_22101,N_21288,N_21002);
nand U22102 (N_22102,N_21552,N_20320);
or U22103 (N_22103,N_20562,N_21231);
nand U22104 (N_22104,N_21308,N_20841);
or U22105 (N_22105,N_21779,N_20450);
nor U22106 (N_22106,N_21226,N_21840);
nand U22107 (N_22107,N_21858,N_21261);
and U22108 (N_22108,N_20776,N_21512);
nand U22109 (N_22109,N_21152,N_20125);
xor U22110 (N_22110,N_20893,N_21525);
xor U22111 (N_22111,N_20310,N_20270);
nand U22112 (N_22112,N_21520,N_21777);
xor U22113 (N_22113,N_21335,N_21809);
and U22114 (N_22114,N_20580,N_21196);
and U22115 (N_22115,N_21625,N_21029);
nand U22116 (N_22116,N_21030,N_20135);
nand U22117 (N_22117,N_21942,N_20986);
and U22118 (N_22118,N_21987,N_20231);
xor U22119 (N_22119,N_21434,N_20142);
nor U22120 (N_22120,N_21179,N_21285);
xnor U22121 (N_22121,N_20658,N_20565);
nor U22122 (N_22122,N_21798,N_20211);
or U22123 (N_22123,N_20722,N_21447);
or U22124 (N_22124,N_21702,N_21250);
or U22125 (N_22125,N_20494,N_21427);
nor U22126 (N_22126,N_20352,N_21523);
or U22127 (N_22127,N_20547,N_20234);
nor U22128 (N_22128,N_21576,N_20291);
nor U22129 (N_22129,N_21460,N_20601);
nand U22130 (N_22130,N_21234,N_20930);
or U22131 (N_22131,N_20199,N_20394);
and U22132 (N_22132,N_20249,N_20708);
or U22133 (N_22133,N_20642,N_20810);
or U22134 (N_22134,N_20523,N_21700);
or U22135 (N_22135,N_20846,N_21327);
or U22136 (N_22136,N_21982,N_20498);
and U22137 (N_22137,N_20051,N_21291);
or U22138 (N_22138,N_21617,N_21468);
nor U22139 (N_22139,N_20030,N_21160);
and U22140 (N_22140,N_21953,N_20360);
xnor U22141 (N_22141,N_21376,N_21225);
xor U22142 (N_22142,N_21395,N_20456);
nand U22143 (N_22143,N_21066,N_21750);
nand U22144 (N_22144,N_20325,N_20627);
xnor U22145 (N_22145,N_21964,N_20491);
and U22146 (N_22146,N_21932,N_21571);
and U22147 (N_22147,N_20090,N_21814);
nand U22148 (N_22148,N_20022,N_21076);
nor U22149 (N_22149,N_20667,N_20109);
or U22150 (N_22150,N_20619,N_20947);
nor U22151 (N_22151,N_21072,N_21875);
and U22152 (N_22152,N_20961,N_20236);
nor U22153 (N_22153,N_21615,N_21522);
and U22154 (N_22154,N_21464,N_20016);
nor U22155 (N_22155,N_20208,N_20455);
nor U22156 (N_22156,N_20747,N_20525);
nor U22157 (N_22157,N_20107,N_20361);
or U22158 (N_22158,N_21493,N_21033);
xnor U22159 (N_22159,N_20269,N_21318);
xnor U22160 (N_22160,N_20818,N_21279);
xor U22161 (N_22161,N_20050,N_20398);
or U22162 (N_22162,N_20307,N_20446);
nor U22163 (N_22163,N_20951,N_21946);
nand U22164 (N_22164,N_20315,N_20383);
xor U22165 (N_22165,N_20426,N_21816);
nor U22166 (N_22166,N_21562,N_20872);
or U22167 (N_22167,N_20624,N_21682);
xnor U22168 (N_22168,N_20247,N_21855);
and U22169 (N_22169,N_21469,N_20449);
and U22170 (N_22170,N_21332,N_21268);
xnor U22171 (N_22171,N_21892,N_21392);
xnor U22172 (N_22172,N_20921,N_20332);
or U22173 (N_22173,N_21040,N_21810);
or U22174 (N_22174,N_21382,N_20528);
or U22175 (N_22175,N_20346,N_21769);
nand U22176 (N_22176,N_20807,N_20008);
or U22177 (N_22177,N_21079,N_21006);
xor U22178 (N_22178,N_21771,N_20935);
nand U22179 (N_22179,N_20848,N_21872);
nand U22180 (N_22180,N_21938,N_21565);
and U22181 (N_22181,N_20423,N_20216);
nor U22182 (N_22182,N_21749,N_20302);
nand U22183 (N_22183,N_21310,N_20709);
nand U22184 (N_22184,N_20255,N_21812);
nor U22185 (N_22185,N_20736,N_21882);
xnor U22186 (N_22186,N_21519,N_21402);
nor U22187 (N_22187,N_21252,N_21055);
or U22188 (N_22188,N_20623,N_20678);
or U22189 (N_22189,N_21101,N_20595);
xnor U22190 (N_22190,N_20052,N_21686);
or U22191 (N_22191,N_21433,N_20611);
or U22192 (N_22192,N_21391,N_20119);
nand U22193 (N_22193,N_21483,N_20330);
nand U22194 (N_22194,N_20928,N_20855);
and U22195 (N_22195,N_20116,N_20732);
xnor U22196 (N_22196,N_21986,N_20400);
xor U22197 (N_22197,N_20864,N_20379);
or U22198 (N_22198,N_21452,N_21516);
or U22199 (N_22199,N_21605,N_20207);
nand U22200 (N_22200,N_20100,N_20675);
xnor U22201 (N_22201,N_20071,N_21111);
or U22202 (N_22202,N_20014,N_21081);
or U22203 (N_22203,N_21128,N_21546);
xnor U22204 (N_22204,N_21497,N_21755);
and U22205 (N_22205,N_20288,N_21550);
xnor U22206 (N_22206,N_21889,N_21450);
nand U22207 (N_22207,N_20243,N_21994);
xor U22208 (N_22208,N_20393,N_20194);
nor U22209 (N_22209,N_21537,N_21919);
or U22210 (N_22210,N_21567,N_20232);
and U22211 (N_22211,N_20965,N_21910);
or U22212 (N_22212,N_21019,N_21539);
or U22213 (N_22213,N_21765,N_21224);
and U22214 (N_22214,N_21059,N_21549);
xnor U22215 (N_22215,N_20962,N_20831);
or U22216 (N_22216,N_20271,N_20727);
nor U22217 (N_22217,N_20614,N_21821);
nand U22218 (N_22218,N_20591,N_20204);
nor U22219 (N_22219,N_20218,N_20173);
xor U22220 (N_22220,N_20783,N_20099);
or U22221 (N_22221,N_20007,N_20911);
xor U22222 (N_22222,N_20964,N_20036);
xnor U22223 (N_22223,N_20480,N_21599);
nand U22224 (N_22224,N_21670,N_21176);
xor U22225 (N_22225,N_20407,N_20088);
nand U22226 (N_22226,N_21815,N_20718);
xnor U22227 (N_22227,N_20942,N_21359);
and U22228 (N_22228,N_20543,N_20669);
or U22229 (N_22229,N_20354,N_21480);
and U22230 (N_22230,N_20275,N_21193);
xnor U22231 (N_22231,N_20188,N_20884);
xnor U22232 (N_22232,N_20552,N_20230);
and U22233 (N_22233,N_21613,N_20899);
nor U22234 (N_22234,N_21362,N_21965);
nand U22235 (N_22235,N_20334,N_20101);
or U22236 (N_22236,N_21566,N_21722);
nor U22237 (N_22237,N_21309,N_20967);
and U22238 (N_22238,N_20822,N_21736);
or U22239 (N_22239,N_21663,N_20277);
nand U22240 (N_22240,N_21314,N_20461);
nand U22241 (N_22241,N_21242,N_20408);
and U22242 (N_22242,N_21557,N_21166);
and U22243 (N_22243,N_20246,N_21822);
nand U22244 (N_22244,N_20129,N_20540);
nor U22245 (N_22245,N_20089,N_21028);
xor U22246 (N_22246,N_20633,N_20548);
xor U22247 (N_22247,N_20663,N_21927);
nand U22248 (N_22248,N_20558,N_20493);
and U22249 (N_22249,N_21577,N_21014);
xnor U22250 (N_22250,N_20802,N_21925);
or U22251 (N_22251,N_20706,N_21851);
xnor U22252 (N_22252,N_21860,N_21159);
xnor U22253 (N_22253,N_20212,N_21021);
nand U22254 (N_22254,N_21284,N_21013);
or U22255 (N_22255,N_20956,N_21619);
or U22256 (N_22256,N_21092,N_20006);
nand U22257 (N_22257,N_21005,N_21529);
or U22258 (N_22258,N_20903,N_21233);
or U22259 (N_22259,N_20733,N_21739);
nand U22260 (N_22260,N_20527,N_21212);
nor U22261 (N_22261,N_20331,N_20752);
and U22262 (N_22262,N_20224,N_20356);
nor U22263 (N_22263,N_20698,N_20327);
or U22264 (N_22264,N_20412,N_21189);
nor U22265 (N_22265,N_21729,N_21060);
xor U22266 (N_22266,N_20021,N_20464);
and U22267 (N_22267,N_21730,N_20377);
nor U22268 (N_22268,N_20995,N_20895);
and U22269 (N_22269,N_21928,N_21770);
nor U22270 (N_22270,N_21175,N_20966);
or U22271 (N_22271,N_21558,N_20359);
nand U22272 (N_22272,N_20997,N_21039);
nor U22273 (N_22273,N_21407,N_21137);
xor U22274 (N_22274,N_20737,N_21954);
xor U22275 (N_22275,N_21177,N_20362);
and U22276 (N_22276,N_21188,N_20998);
nor U22277 (N_22277,N_20832,N_21416);
nand U22278 (N_22278,N_21228,N_21764);
xnor U22279 (N_22279,N_20524,N_20322);
and U22280 (N_22280,N_21967,N_21826);
and U22281 (N_22281,N_21758,N_21397);
and U22282 (N_22282,N_21342,N_21262);
and U22283 (N_22283,N_20617,N_21149);
nand U22284 (N_22284,N_21247,N_20285);
nor U22285 (N_22285,N_21052,N_20556);
and U22286 (N_22286,N_20780,N_21908);
nor U22287 (N_22287,N_20665,N_21939);
or U22288 (N_22288,N_21269,N_21996);
nor U22289 (N_22289,N_20978,N_21687);
or U22290 (N_22290,N_21514,N_21479);
nand U22291 (N_22291,N_20813,N_21618);
nor U22292 (N_22292,N_20634,N_20908);
and U22293 (N_22293,N_21120,N_21951);
xnor U22294 (N_22294,N_21344,N_21354);
xor U22295 (N_22295,N_20108,N_20469);
nor U22296 (N_22296,N_21740,N_20905);
nand U22297 (N_22297,N_21587,N_21854);
or U22298 (N_22298,N_21667,N_21944);
or U22299 (N_22299,N_21375,N_20144);
nand U22300 (N_22300,N_20084,N_21315);
and U22301 (N_22301,N_20343,N_20742);
and U22302 (N_22302,N_21063,N_21714);
xnor U22303 (N_22303,N_21424,N_21334);
and U22304 (N_22304,N_20280,N_20987);
xor U22305 (N_22305,N_20629,N_21961);
nor U22306 (N_22306,N_20782,N_21378);
and U22307 (N_22307,N_21357,N_20662);
nor U22308 (N_22308,N_21136,N_21785);
nand U22309 (N_22309,N_21743,N_20048);
and U22310 (N_22310,N_20228,N_21924);
and U22311 (N_22311,N_21298,N_21646);
or U22312 (N_22312,N_20415,N_21559);
xnor U22313 (N_22313,N_21890,N_20474);
or U22314 (N_22314,N_21979,N_21548);
nand U22315 (N_22315,N_20712,N_21163);
and U22316 (N_22316,N_20594,N_20413);
nand U22317 (N_22317,N_20166,N_21461);
xor U22318 (N_22318,N_21595,N_21883);
and U22319 (N_22319,N_21453,N_20424);
nand U22320 (N_22320,N_20342,N_20248);
xor U22321 (N_22321,N_20133,N_21787);
and U22322 (N_22322,N_21139,N_20857);
xnor U22323 (N_22323,N_20992,N_20862);
and U22324 (N_22324,N_21866,N_21845);
and U22325 (N_22325,N_20176,N_20260);
or U22326 (N_22326,N_20719,N_21995);
or U22327 (N_22327,N_20150,N_21110);
or U22328 (N_22328,N_20656,N_21975);
xor U22329 (N_22329,N_21150,N_21472);
nand U22330 (N_22330,N_21051,N_20881);
nand U22331 (N_22331,N_21992,N_21142);
nand U22332 (N_22332,N_21676,N_21330);
or U22333 (N_22333,N_21394,N_20489);
nor U22334 (N_22334,N_20652,N_21368);
and U22335 (N_22335,N_21209,N_20097);
nor U22336 (N_22336,N_21780,N_21620);
nor U22337 (N_22337,N_21828,N_21095);
or U22338 (N_22338,N_20374,N_20447);
or U22339 (N_22339,N_20182,N_20631);
nor U22340 (N_22340,N_21251,N_21943);
or U22341 (N_22341,N_20878,N_21585);
and U22342 (N_22342,N_20106,N_21151);
nor U22343 (N_22343,N_21598,N_21672);
nand U22344 (N_22344,N_21665,N_20258);
nor U22345 (N_22345,N_20683,N_20314);
nand U22346 (N_22346,N_20438,N_21610);
and U22347 (N_22347,N_21915,N_20420);
or U22348 (N_22348,N_21506,N_21374);
nor U22349 (N_22349,N_21968,N_21448);
or U22350 (N_22350,N_21664,N_20797);
xor U22351 (N_22351,N_20516,N_21048);
and U22352 (N_22352,N_21074,N_20061);
or U22353 (N_22353,N_21263,N_20605);
and U22354 (N_22354,N_21421,N_21373);
xor U22355 (N_22355,N_21756,N_21347);
nand U22356 (N_22356,N_20730,N_20115);
or U22357 (N_22357,N_20297,N_20766);
or U22358 (N_22358,N_21836,N_21738);
nor U22359 (N_22359,N_21984,N_20778);
or U22360 (N_22360,N_21396,N_20227);
nor U22361 (N_22361,N_20148,N_20004);
or U22362 (N_22362,N_21477,N_20684);
and U22363 (N_22363,N_20122,N_21999);
nand U22364 (N_22364,N_21099,N_20127);
and U22365 (N_22365,N_21216,N_20724);
nand U22366 (N_22366,N_20784,N_20179);
nand U22367 (N_22367,N_21069,N_21435);
nor U22368 (N_22368,N_20808,N_20944);
and U22369 (N_22369,N_21123,N_21294);
nor U22370 (N_22370,N_21496,N_21365);
nor U22371 (N_22371,N_20859,N_21265);
xor U22372 (N_22372,N_20606,N_20278);
or U22373 (N_22373,N_20839,N_21426);
or U22374 (N_22374,N_21235,N_21017);
and U22375 (N_22375,N_21126,N_20184);
and U22376 (N_22376,N_20679,N_20536);
nor U22377 (N_22377,N_20825,N_21199);
nand U22378 (N_22378,N_20936,N_21835);
or U22379 (N_22379,N_20830,N_21936);
xnor U22380 (N_22380,N_20993,N_20056);
nand U22381 (N_22381,N_21119,N_21210);
or U22382 (N_22382,N_20147,N_21141);
nor U22383 (N_22383,N_21930,N_20460);
nor U22384 (N_22384,N_20254,N_21922);
nor U22385 (N_22385,N_20777,N_21590);
nor U22386 (N_22386,N_20472,N_21476);
or U22387 (N_22387,N_20588,N_21379);
or U22388 (N_22388,N_21276,N_20095);
nor U22389 (N_22389,N_21097,N_20820);
nand U22390 (N_22390,N_20957,N_21602);
nand U22391 (N_22391,N_20968,N_20032);
nor U22392 (N_22392,N_20468,N_21551);
nor U22393 (N_22393,N_20785,N_21582);
and U22394 (N_22394,N_21720,N_20418);
nand U22395 (N_22395,N_21306,N_20894);
or U22396 (N_22396,N_20687,N_21118);
or U22397 (N_22397,N_20265,N_21513);
nand U22398 (N_22398,N_21471,N_20209);
or U22399 (N_22399,N_21773,N_20110);
and U22400 (N_22400,N_21906,N_21848);
or U22401 (N_22401,N_20599,N_21180);
or U22402 (N_22402,N_21358,N_20217);
nor U22403 (N_22403,N_21923,N_21547);
or U22404 (N_22404,N_21600,N_20927);
and U22405 (N_22405,N_20436,N_21114);
nand U22406 (N_22406,N_20312,N_20983);
nor U22407 (N_22407,N_21403,N_21409);
xor U22408 (N_22408,N_20738,N_20452);
and U22409 (N_22409,N_20244,N_21026);
xor U22410 (N_22410,N_21047,N_20075);
or U22411 (N_22411,N_21653,N_21721);
or U22412 (N_22412,N_20293,N_20430);
and U22413 (N_22413,N_21579,N_20156);
and U22414 (N_22414,N_21684,N_21135);
and U22415 (N_22415,N_21312,N_20542);
nand U22416 (N_22416,N_21793,N_20816);
or U22417 (N_22417,N_20649,N_20324);
xor U22418 (N_22418,N_21331,N_20091);
and U22419 (N_22419,N_21217,N_21989);
nand U22420 (N_22420,N_21274,N_20009);
xnor U22421 (N_22421,N_21132,N_21753);
nor U22422 (N_22422,N_20870,N_21695);
nand U22423 (N_22423,N_21626,N_21668);
nor U22424 (N_22424,N_20584,N_21232);
nor U22425 (N_22425,N_20086,N_21473);
or U22426 (N_22426,N_20837,N_21190);
xnor U22427 (N_22427,N_21837,N_20775);
nor U22428 (N_22428,N_21824,N_20800);
and U22429 (N_22429,N_20237,N_21657);
nand U22430 (N_22430,N_21321,N_20721);
and U22431 (N_22431,N_20402,N_20901);
or U22432 (N_22432,N_21857,N_20187);
or U22433 (N_22433,N_20759,N_20010);
or U22434 (N_22434,N_21666,N_21597);
or U22435 (N_22435,N_20817,N_20466);
and U22436 (N_22436,N_21578,N_21732);
nor U22437 (N_22437,N_21909,N_20760);
xnor U22438 (N_22438,N_20058,N_20892);
xnor U22439 (N_22439,N_21877,N_20405);
nor U22440 (N_22440,N_21023,N_20575);
xor U22441 (N_22441,N_20039,N_21536);
or U22442 (N_22442,N_21897,N_20787);
nor U22443 (N_22443,N_20579,N_20335);
or U22444 (N_22444,N_20401,N_21959);
nand U22445 (N_22445,N_21143,N_20000);
and U22446 (N_22446,N_21355,N_20363);
nor U22447 (N_22447,N_20080,N_20751);
xnor U22448 (N_22448,N_20268,N_20259);
nand U22449 (N_22449,N_20497,N_21441);
nor U22450 (N_22450,N_21680,N_21737);
xnor U22451 (N_22451,N_20852,N_20477);
nor U22452 (N_22452,N_20958,N_20192);
nand U22453 (N_22453,N_21246,N_20786);
xnor U22454 (N_22454,N_20996,N_21299);
or U22455 (N_22455,N_20843,N_21366);
xnor U22456 (N_22456,N_20913,N_21042);
and U22457 (N_22457,N_20272,N_21891);
or U22458 (N_22458,N_20750,N_21887);
nand U22459 (N_22459,N_21349,N_20459);
nor U22460 (N_22460,N_20338,N_20365);
nor U22461 (N_22461,N_20796,N_21213);
nand U22462 (N_22462,N_20409,N_20251);
and U22463 (N_22463,N_21148,N_21078);
and U22464 (N_22464,N_20301,N_21162);
xnor U22465 (N_22465,N_20755,N_20561);
xnor U22466 (N_22466,N_20814,N_20926);
and U22467 (N_22467,N_21904,N_20351);
nor U22468 (N_22468,N_21916,N_20168);
or U22469 (N_22469,N_21363,N_21735);
xnor U22470 (N_22470,N_20533,N_21316);
xnor U22471 (N_22471,N_20537,N_20674);
nand U22472 (N_22472,N_21408,N_21036);
nand U22473 (N_22473,N_20308,N_20482);
xnor U22474 (N_22474,N_21914,N_21811);
xnor U22475 (N_22475,N_20203,N_20758);
nor U22476 (N_22476,N_21445,N_21161);
nor U22477 (N_22477,N_21649,N_20059);
nor U22478 (N_22478,N_20898,N_21621);
and U22479 (N_22479,N_21832,N_21733);
nor U22480 (N_22480,N_20568,N_20851);
nand U22481 (N_22481,N_21699,N_21825);
or U22482 (N_22482,N_20417,N_21988);
nand U22483 (N_22483,N_21459,N_20451);
or U22484 (N_22484,N_21712,N_20661);
and U22485 (N_22485,N_20355,N_20768);
nand U22486 (N_22486,N_21351,N_21384);
or U22487 (N_22487,N_21542,N_21874);
and U22488 (N_22488,N_21829,N_21289);
xnor U22489 (N_22489,N_20651,N_21528);
and U22490 (N_22490,N_20704,N_20849);
nand U22491 (N_22491,N_20429,N_21719);
or U22492 (N_22492,N_20647,N_20769);
nand U22493 (N_22493,N_20347,N_21009);
and U22494 (N_22494,N_20850,N_21301);
and U22495 (N_22495,N_21018,N_21650);
nor U22496 (N_22496,N_21239,N_20492);
or U22497 (N_22497,N_21035,N_20574);
or U22498 (N_22498,N_21432,N_20162);
or U22499 (N_22499,N_21926,N_20519);
or U22500 (N_22500,N_20842,N_21797);
and U22501 (N_22501,N_20102,N_20639);
nor U22502 (N_22502,N_20309,N_21716);
or U22503 (N_22503,N_21096,N_20811);
or U22504 (N_22504,N_20969,N_20070);
nor U22505 (N_22505,N_20515,N_20972);
nor U22506 (N_22506,N_20073,N_20049);
xnor U22507 (N_22507,N_20686,N_20971);
and U22508 (N_22508,N_21871,N_20779);
nand U22509 (N_22509,N_21041,N_21352);
nand U22510 (N_22510,N_21266,N_20794);
and U22511 (N_22511,N_20411,N_21498);
and U22512 (N_22512,N_20483,N_20512);
xor U22513 (N_22513,N_21016,N_20860);
and U22514 (N_22514,N_21186,N_20284);
or U22515 (N_22515,N_20353,N_21962);
xnor U22516 (N_22516,N_21846,N_21774);
nand U22517 (N_22517,N_20549,N_20345);
and U22518 (N_22518,N_20012,N_20991);
nor U22519 (N_22519,N_20520,N_20945);
nor U22520 (N_22520,N_20261,N_21348);
or U22521 (N_22521,N_20457,N_21913);
and U22522 (N_22522,N_20373,N_21146);
nand U22523 (N_22523,N_20300,N_20196);
or U22524 (N_22524,N_20553,N_20676);
nor U22525 (N_22525,N_20932,N_20950);
xnor U22526 (N_22526,N_21184,N_21591);
nand U22527 (N_22527,N_21273,N_20286);
and U22528 (N_22528,N_20055,N_20670);
nand U22529 (N_22529,N_21286,N_21086);
and U22530 (N_22530,N_21131,N_20638);
xor U22531 (N_22531,N_21713,N_20295);
and U22532 (N_22532,N_21776,N_20488);
nand U22533 (N_22533,N_21534,N_21823);
and U22534 (N_22534,N_20238,N_20130);
and U22535 (N_22535,N_21580,N_20691);
or U22536 (N_22536,N_21834,N_20929);
and U22537 (N_22537,N_21561,N_21238);
nor U22538 (N_22538,N_20403,N_20880);
xor U22539 (N_22539,N_20399,N_20541);
nor U22540 (N_22540,N_20387,N_20746);
xor U22541 (N_22541,N_20636,N_21974);
and U22542 (N_22542,N_20762,N_21420);
nor U22543 (N_22543,N_20479,N_21103);
and U22544 (N_22544,N_20875,N_21631);
and U22545 (N_22545,N_20716,N_20970);
nor U22546 (N_22546,N_21532,N_21317);
xor U22547 (N_22547,N_20281,N_21708);
nand U22548 (N_22548,N_21297,N_20038);
xnor U22549 (N_22549,N_20074,N_21588);
or U22550 (N_22550,N_20427,N_21544);
xnor U22551 (N_22551,N_20490,N_21438);
nor U22552 (N_22552,N_20311,N_20121);
xnor U22553 (N_22553,N_21197,N_20630);
nand U22554 (N_22554,N_20161,N_20767);
nor U22555 (N_22555,N_21004,N_21043);
nor U22556 (N_22556,N_21011,N_21381);
nand U22557 (N_22557,N_21698,N_20078);
nor U22558 (N_22558,N_20583,N_21302);
nand U22559 (N_22559,N_20919,N_21731);
nor U22560 (N_22560,N_21454,N_20282);
nor U22561 (N_22561,N_20462,N_21428);
nor U22562 (N_22562,N_21287,N_20191);
nand U22563 (N_22563,N_20729,N_20508);
and U22564 (N_22564,N_21489,N_20664);
nor U22565 (N_22565,N_21198,N_20486);
xnor U22566 (N_22566,N_21990,N_21681);
nor U22567 (N_22567,N_20406,N_21885);
nor U22568 (N_22568,N_21221,N_20013);
and U22569 (N_22569,N_20749,N_21661);
or U22570 (N_22570,N_20589,N_20764);
xor U22571 (N_22571,N_21338,N_21050);
nand U22572 (N_22572,N_20026,N_21648);
and U22573 (N_22573,N_21642,N_21640);
or U22574 (N_22574,N_20564,N_20471);
nand U22575 (N_22575,N_21675,N_21842);
or U22576 (N_22576,N_21191,N_21751);
and U22577 (N_22577,N_21328,N_20174);
xor U22578 (N_22578,N_20046,N_20854);
or U22579 (N_22579,N_20696,N_20313);
nor U22580 (N_22580,N_20694,N_20827);
nor U22581 (N_22581,N_20481,N_21223);
nand U22582 (N_22582,N_21208,N_21282);
nor U22583 (N_22583,N_20973,N_21501);
and U22584 (N_22584,N_21876,N_20643);
nor U22585 (N_22585,N_21745,N_21105);
and U22586 (N_22586,N_20376,N_21538);
nand U22587 (N_22587,N_20578,N_20205);
or U22588 (N_22588,N_21109,N_20989);
and U22589 (N_22589,N_20041,N_20391);
and U22590 (N_22590,N_21027,N_21304);
and U22591 (N_22591,N_20287,N_20392);
or U22592 (N_22592,N_21122,N_21767);
or U22593 (N_22593,N_21073,N_21905);
and U22594 (N_22594,N_20602,N_21659);
nor U22595 (N_22595,N_21490,N_21255);
and U22596 (N_22596,N_20981,N_20124);
or U22597 (N_22597,N_20453,N_20963);
nor U22598 (N_22598,N_21296,N_20226);
nor U22599 (N_22599,N_21966,N_20499);
and U22600 (N_22600,N_21254,N_20098);
and U22601 (N_22601,N_20378,N_20165);
and U22602 (N_22602,N_21917,N_20573);
or U22603 (N_22603,N_21182,N_20990);
nand U22604 (N_22604,N_20180,N_20502);
and U22605 (N_22605,N_21367,N_20020);
and U22606 (N_22606,N_20487,N_21586);
nand U22607 (N_22607,N_21662,N_21195);
xnor U22608 (N_22608,N_20024,N_21145);
nand U22609 (N_22609,N_20195,N_20641);
and U22610 (N_22610,N_20214,N_20114);
xor U22611 (N_22611,N_20735,N_21794);
and U22612 (N_22612,N_20120,N_20890);
or U22613 (N_22613,N_21267,N_21085);
and U22614 (N_22614,N_20319,N_21140);
xnor U22615 (N_22615,N_21937,N_21820);
and U22616 (N_22616,N_20511,N_20739);
xnor U22617 (N_22617,N_21307,N_21084);
or U22618 (N_22618,N_21046,N_21692);
nor U22619 (N_22619,N_20985,N_21504);
nand U22620 (N_22620,N_21157,N_21592);
or U22621 (N_22621,N_20458,N_20298);
or U22622 (N_22622,N_21116,N_20845);
nor U22623 (N_22623,N_20648,N_21518);
and U22624 (N_22624,N_20177,N_20840);
xor U22625 (N_22625,N_20607,N_20337);
xnor U22626 (N_22626,N_21696,N_21673);
or U22627 (N_22627,N_21022,N_20060);
nand U22628 (N_22628,N_21654,N_21067);
nand U22629 (N_22629,N_21248,N_20941);
xnor U22630 (N_22630,N_20657,N_21818);
nand U22631 (N_22631,N_20141,N_20943);
nand U22632 (N_22632,N_21121,N_21495);
and U22633 (N_22633,N_21277,N_20801);
and U22634 (N_22634,N_21108,N_21485);
nor U22635 (N_22635,N_21817,N_20132);
nor U22636 (N_22636,N_20954,N_21313);
and U22637 (N_22637,N_20933,N_20646);
xor U22638 (N_22638,N_20707,N_20526);
nand U22639 (N_22639,N_20546,N_20654);
or U22640 (N_22640,N_20644,N_21934);
nand U22641 (N_22641,N_21693,N_21704);
and U22642 (N_22642,N_20598,N_21847);
xnor U22643 (N_22643,N_21138,N_20946);
or U22644 (N_22644,N_20838,N_20715);
nor U22645 (N_22645,N_20158,N_20096);
nand U22646 (N_22646,N_20485,N_20475);
or U22647 (N_22647,N_20616,N_21978);
nor U22648 (N_22648,N_20539,N_20410);
nand U22649 (N_22649,N_20358,N_20220);
or U22650 (N_22650,N_20428,N_20975);
nor U22651 (N_22651,N_20914,N_20172);
nor U22652 (N_22652,N_20292,N_21957);
nand U22653 (N_22653,N_20874,N_21458);
and U22654 (N_22654,N_20029,N_21604);
nand U22655 (N_22655,N_20823,N_21775);
nand U22656 (N_22656,N_20221,N_20576);
nor U22657 (N_22657,N_20867,N_21154);
nor U22658 (N_22658,N_21669,N_20414);
nand U22659 (N_22659,N_20303,N_20960);
nor U22660 (N_22660,N_20774,N_20323);
nand U22661 (N_22661,N_20183,N_21660);
xor U22662 (N_22662,N_21449,N_21861);
or U22663 (N_22663,N_20812,N_20517);
xnor U22664 (N_22664,N_20390,N_20912);
or U22665 (N_22665,N_21507,N_21214);
nor U22666 (N_22666,N_21205,N_21372);
nand U22667 (N_22667,N_21744,N_21444);
nand U22668 (N_22668,N_21414,N_20530);
and U22669 (N_22669,N_21584,N_21488);
nor U22670 (N_22670,N_21690,N_21614);
nand U22671 (N_22671,N_20045,N_20886);
xor U22672 (N_22672,N_20805,N_21194);
nor U22673 (N_22673,N_21867,N_21895);
nand U22674 (N_22674,N_21423,N_21630);
or U22675 (N_22675,N_20570,N_21833);
xnor U22676 (N_22676,N_20146,N_20210);
nor U22677 (N_22677,N_21056,N_20093);
and U22678 (N_22678,N_20745,N_21945);
and U22679 (N_22679,N_21089,N_21678);
xor U22680 (N_22680,N_21863,N_21113);
nor U22681 (N_22681,N_21003,N_21624);
and U22682 (N_22682,N_21156,N_20999);
nand U22683 (N_22683,N_20223,N_20885);
nand U22684 (N_22684,N_20344,N_20185);
and U22685 (N_22685,N_20085,N_21893);
nor U22686 (N_22686,N_21958,N_21064);
nand U22687 (N_22687,N_21020,N_20910);
xor U22688 (N_22688,N_20743,N_20861);
nor U22689 (N_22689,N_21419,N_21088);
and U22690 (N_22690,N_21998,N_21503);
nor U22691 (N_22691,N_20416,N_21360);
or U22692 (N_22692,N_21881,N_20470);
nor U22693 (N_22693,N_21907,N_20443);
or U22694 (N_22694,N_21170,N_20015);
xor U22695 (N_22695,N_21763,N_21638);
or U22696 (N_22696,N_20835,N_20612);
nor U22697 (N_22697,N_20668,N_20186);
nor U22698 (N_22698,N_21383,N_20824);
and U22699 (N_22699,N_21486,N_21456);
or U22700 (N_22700,N_21575,N_20131);
nor U22701 (N_22701,N_21850,N_21508);
nor U22702 (N_22702,N_21609,N_20635);
nor U22703 (N_22703,N_20994,N_21442);
or U22704 (N_22704,N_21628,N_20290);
nor U22705 (N_22705,N_21969,N_21353);
nor U22706 (N_22706,N_20266,N_20902);
and U22707 (N_22707,N_21805,N_21062);
or U22708 (N_22708,N_20637,N_21760);
nor U22709 (N_22709,N_20609,N_20349);
xnor U22710 (N_22710,N_21192,N_21746);
nor U22711 (N_22711,N_21983,N_20608);
or U22712 (N_22712,N_21491,N_20160);
nand U22713 (N_22713,N_21500,N_20397);
and U22714 (N_22714,N_20035,N_20279);
nand U22715 (N_22715,N_20128,N_21098);
nand U22716 (N_22716,N_20597,N_20711);
xor U22717 (N_22717,N_21762,N_20189);
nand U22718 (N_22718,N_21371,N_20233);
and U22719 (N_22719,N_20871,N_21385);
or U22720 (N_22720,N_21115,N_20863);
nand U22721 (N_22721,N_21244,N_20092);
and U22722 (N_22722,N_21024,N_20368);
or U22723 (N_22723,N_20478,N_21950);
xnor U22724 (N_22724,N_21303,N_20844);
nand U22725 (N_22725,N_21153,N_20876);
nand U22726 (N_22726,N_21710,N_21694);
nor U22727 (N_22727,N_20826,N_21015);
nand U22728 (N_22728,N_20350,N_20171);
xor U22729 (N_22729,N_21405,N_21725);
or U22730 (N_22730,N_21869,N_21784);
or U22731 (N_22731,N_21124,N_21203);
nor U22732 (N_22732,N_21838,N_21804);
and U22733 (N_22733,N_20037,N_21264);
xor U22734 (N_22734,N_20381,N_21008);
xnor U22735 (N_22735,N_20699,N_20916);
and U22736 (N_22736,N_20140,N_20364);
or U22737 (N_22737,N_20620,N_20713);
and U22738 (N_22738,N_21054,N_21517);
nand U22739 (N_22739,N_20467,N_20695);
or U22740 (N_22740,N_20219,N_21900);
nor U22741 (N_22741,N_20940,N_20798);
and U22742 (N_22742,N_21350,N_20959);
or U22743 (N_22743,N_21947,N_20792);
xnor U22744 (N_22744,N_21572,N_20550);
nor U22745 (N_22745,N_20053,N_21717);
or U22746 (N_22746,N_21635,N_20465);
nor U22747 (N_22747,N_21896,N_20673);
nor U22748 (N_22748,N_21807,N_20170);
or U22749 (N_22749,N_21727,N_20370);
and U22750 (N_22750,N_21759,N_20375);
xor U22751 (N_22751,N_21723,N_21241);
or U22752 (N_22752,N_20915,N_20422);
xnor U22753 (N_22753,N_20388,N_21612);
or U22754 (N_22754,N_21791,N_21465);
and U22755 (N_22755,N_20431,N_20593);
and U22756 (N_22756,N_20976,N_21399);
xor U22757 (N_22757,N_21311,N_20501);
and U22758 (N_22758,N_21734,N_21127);
and U22759 (N_22759,N_21683,N_20437);
xor U22760 (N_22760,N_20421,N_21075);
or U22761 (N_22761,N_20628,N_20340);
and U22762 (N_22762,N_21752,N_20239);
and U22763 (N_22763,N_20264,N_21256);
or U22764 (N_22764,N_20560,N_21229);
or U22765 (N_22765,N_21671,N_21754);
xor U22766 (N_22766,N_20920,N_20688);
nor U22767 (N_22767,N_21437,N_21061);
or U22768 (N_22768,N_21183,N_20510);
nand U22769 (N_22769,N_21093,N_21880);
nor U22770 (N_22770,N_20672,N_21583);
nand U22771 (N_22771,N_20939,N_20555);
nand U22772 (N_22772,N_20865,N_21343);
nand U22773 (N_22773,N_20931,N_20666);
nand U22774 (N_22774,N_21918,N_21560);
nand U22775 (N_22775,N_20250,N_21819);
nand U22776 (N_22776,N_20531,N_21865);
and U22777 (N_22777,N_20252,N_20028);
xor U22778 (N_22778,N_20504,N_20934);
xor U22779 (N_22779,N_20081,N_20522);
nand U22780 (N_22780,N_20952,N_20137);
nor U22781 (N_22781,N_20567,N_20581);
xnor U22782 (N_22782,N_20680,N_21475);
or U22783 (N_22783,N_20988,N_20883);
and U22784 (N_22784,N_20681,N_20372);
nand U22785 (N_22785,N_20367,N_20366);
nand U22786 (N_22786,N_21651,N_21707);
xor U22787 (N_22787,N_21130,N_20980);
and U22788 (N_22788,N_20917,N_21786);
xnor U22789 (N_22789,N_21070,N_21623);
xor U22790 (N_22790,N_20771,N_20761);
xor U22791 (N_22791,N_20435,N_20262);
nand U22792 (N_22792,N_21206,N_21057);
xnor U22793 (N_22793,N_21972,N_20329);
and U22794 (N_22794,N_21413,N_21553);
xnor U22795 (N_22795,N_20193,N_20790);
nand U22796 (N_22796,N_20341,N_21406);
or U22797 (N_22797,N_21611,N_21570);
nor U22798 (N_22798,N_21253,N_20159);
or U22799 (N_22799,N_20534,N_21715);
xnor U22800 (N_22800,N_21524,N_21167);
nand U22801 (N_22801,N_20879,N_21728);
nand U22802 (N_22802,N_21129,N_20877);
nor U22803 (N_22803,N_20257,N_21494);
xor U22804 (N_22804,N_20382,N_20833);
and U22805 (N_22805,N_21911,N_20138);
or U22806 (N_22806,N_21531,N_20615);
xnor U22807 (N_22807,N_20948,N_20521);
and U22808 (N_22808,N_20263,N_20118);
xor U22809 (N_22809,N_20017,N_20748);
nand U22810 (N_22810,N_21884,N_20572);
nand U22811 (N_22811,N_20380,N_21789);
or U22812 (N_22812,N_20145,N_21674);
xnor U22813 (N_22813,N_20304,N_21341);
or U22814 (N_22814,N_20505,N_20770);
nand U22815 (N_22815,N_21482,N_20063);
or U22816 (N_22816,N_21411,N_21499);
xnor U22817 (N_22817,N_20799,N_20253);
and U22818 (N_22818,N_20551,N_21899);
or U22819 (N_22819,N_21077,N_21323);
and U22820 (N_22820,N_20834,N_20134);
and U22821 (N_22821,N_20201,N_21364);
xor U22822 (N_22822,N_21100,N_20604);
nor U22823 (N_22823,N_21637,N_20001);
xor U22824 (N_22824,N_21912,N_20386);
or U22825 (N_22825,N_20847,N_20496);
nor U22826 (N_22826,N_20710,N_21568);
xor U22827 (N_22827,N_20563,N_20034);
nor U22828 (N_22828,N_20763,N_21970);
nor U22829 (N_22829,N_21211,N_20240);
or U22830 (N_22830,N_21903,N_20659);
nand U22831 (N_22831,N_20585,N_21202);
and U22832 (N_22832,N_20043,N_21158);
nand U22833 (N_22833,N_21554,N_21859);
xor U22834 (N_22834,N_20754,N_21766);
or U22835 (N_22835,N_20276,N_20215);
and U22836 (N_22836,N_21398,N_21053);
and U22837 (N_22837,N_21102,N_20274);
xnor U22838 (N_22838,N_20117,N_21831);
nand U22839 (N_22839,N_20019,N_21080);
and U22840 (N_22840,N_21878,N_20532);
or U22841 (N_22841,N_21240,N_20723);
or U22842 (N_22842,N_20650,N_20190);
xor U22843 (N_22843,N_21325,N_20828);
and U22844 (N_22844,N_21336,N_21168);
nor U22845 (N_22845,N_21581,N_20725);
or U22846 (N_22846,N_20731,N_20175);
nor U22847 (N_22847,N_21272,N_21430);
and U22848 (N_22848,N_20318,N_21440);
and U22849 (N_22849,N_21701,N_20283);
or U22850 (N_22850,N_21886,N_20087);
nor U22851 (N_22851,N_20645,N_20181);
nand U22852 (N_22852,N_21218,N_21511);
or U22853 (N_22853,N_20289,N_21691);
nand U22854 (N_22854,N_21369,N_21417);
or U22855 (N_22855,N_21305,N_20554);
nor U22856 (N_22856,N_20781,N_21768);
and U22857 (N_22857,N_21718,N_21629);
nand U22858 (N_22858,N_20306,N_20756);
nand U22859 (N_22859,N_20202,N_20371);
nor U22860 (N_22860,N_21622,N_20440);
and U22861 (N_22861,N_21644,N_20033);
xnor U22862 (N_22862,N_21236,N_21976);
and U22863 (N_22863,N_20432,N_21778);
nor U22864 (N_22864,N_21589,N_20067);
nor U22865 (N_22865,N_20586,N_20389);
and U22866 (N_22866,N_21259,N_20626);
nor U22867 (N_22867,N_21219,N_20888);
nand U22868 (N_22868,N_20625,N_20682);
and U22869 (N_22869,N_20169,N_21388);
and U22870 (N_22870,N_20923,N_20152);
and U22871 (N_22871,N_21960,N_21032);
nor U22872 (N_22872,N_20065,N_20937);
nor U22873 (N_22873,N_20027,N_20094);
nor U22874 (N_22874,N_20984,N_21470);
xor U22875 (N_22875,N_21144,N_20557);
and U22876 (N_22876,N_20907,N_20068);
nor U22877 (N_22877,N_21783,N_21377);
xor U22878 (N_22878,N_21090,N_21227);
nor U22879 (N_22879,N_20697,N_20425);
or U22880 (N_22880,N_21133,N_21981);
nor U22881 (N_22881,N_21083,N_20267);
nor U22882 (N_22882,N_20005,N_20772);
nand U22883 (N_22883,N_21481,N_21802);
xnor U22884 (N_22884,N_21841,N_20062);
and U22885 (N_22885,N_20720,N_21393);
xor U22886 (N_22886,N_21569,N_21843);
xor U22887 (N_22887,N_21564,N_20151);
xor U22888 (N_22888,N_20977,N_20384);
nor U22889 (N_22889,N_21980,N_21703);
and U22890 (N_22890,N_20918,N_21527);
or U22891 (N_22891,N_21346,N_21806);
nand U22892 (N_22892,N_21788,N_20590);
nor U22893 (N_22893,N_20002,N_21466);
xor U22894 (N_22894,N_20164,N_21322);
nand U22895 (N_22895,N_21830,N_21410);
nand U22896 (N_22896,N_21530,N_21677);
and U22897 (N_22897,N_21509,N_20765);
xor U22898 (N_22898,N_21478,N_20507);
nor U22899 (N_22899,N_21058,N_20734);
nand U22900 (N_22900,N_20677,N_20197);
nor U22901 (N_22901,N_20439,N_20904);
xor U22902 (N_22902,N_20294,N_20653);
nand U22903 (N_22903,N_21457,N_20922);
or U22904 (N_22904,N_20139,N_21633);
nor U22905 (N_22905,N_21901,N_21792);
xnor U22906 (N_22906,N_21697,N_20054);
nor U22907 (N_22907,N_21094,N_21636);
nor U22908 (N_22908,N_21741,N_21772);
or U22909 (N_22909,N_20484,N_21641);
and U22910 (N_22910,N_21603,N_20025);
or U22911 (N_22911,N_20077,N_21439);
xor U22912 (N_22912,N_20603,N_21404);
nor U22913 (N_22913,N_21799,N_21545);
nor U22914 (N_22914,N_20660,N_21270);
nor U22915 (N_22915,N_20178,N_20083);
and U22916 (N_22916,N_21933,N_21902);
nand U22917 (N_22917,N_21726,N_21178);
and U22918 (N_22918,N_20509,N_21656);
and U22919 (N_22919,N_20111,N_21606);
or U22920 (N_22920,N_21380,N_20974);
or U22921 (N_22921,N_20163,N_21563);
or U22922 (N_22922,N_20900,N_20143);
or U22923 (N_22923,N_20011,N_21243);
nor U22924 (N_22924,N_21329,N_21849);
and U22925 (N_22925,N_20448,N_20316);
nor U22926 (N_22926,N_21991,N_20690);
nand U22927 (N_22927,N_20587,N_21169);
xor U22928 (N_22928,N_20671,N_20225);
and U22929 (N_22929,N_21155,N_20600);
xor U22930 (N_22930,N_20896,N_21862);
xnor U22931 (N_22931,N_20040,N_21535);
xor U22932 (N_22932,N_20806,N_21688);
nand U22933 (N_22933,N_20104,N_20815);
nor U22934 (N_22934,N_21803,N_20057);
nor U22935 (N_22935,N_20396,N_21324);
and U22936 (N_22936,N_21260,N_21010);
and U22937 (N_22937,N_21091,N_20700);
and U22938 (N_22938,N_21977,N_21931);
or U22939 (N_22939,N_21948,N_20317);
and U22940 (N_22940,N_21000,N_21326);
xor U22941 (N_22941,N_21645,N_20442);
and U22942 (N_22942,N_20836,N_21747);
nor U22943 (N_22943,N_20538,N_21337);
and U22944 (N_22944,N_21920,N_21467);
or U22945 (N_22945,N_20385,N_20256);
or U22946 (N_22946,N_20789,N_21082);
nand U22947 (N_22947,N_20123,N_21422);
xor U22948 (N_22948,N_20069,N_20529);
or U22949 (N_22949,N_21333,N_21147);
nor U22950 (N_22950,N_20577,N_21796);
and U22951 (N_22951,N_20793,N_21412);
or U22952 (N_22952,N_20953,N_20955);
or U22953 (N_22953,N_20082,N_21418);
and U22954 (N_22954,N_21339,N_20873);
nand U22955 (N_22955,N_21249,N_20909);
or U22956 (N_22956,N_21868,N_20692);
and U22957 (N_22957,N_20829,N_21574);
xor U22958 (N_22958,N_21601,N_21782);
or U22959 (N_22959,N_20513,N_21853);
xor U22960 (N_22960,N_21608,N_21071);
nand U22961 (N_22961,N_20506,N_21431);
or U22962 (N_22962,N_21390,N_21165);
and U22963 (N_22963,N_20728,N_20296);
nand U22964 (N_22964,N_20476,N_20395);
and U22965 (N_22965,N_20200,N_21340);
and U22966 (N_22966,N_21400,N_21293);
nand U22967 (N_22967,N_20206,N_20569);
xnor U22968 (N_22968,N_21839,N_20066);
xnor U22969 (N_22969,N_20153,N_21245);
or U22970 (N_22970,N_21436,N_20582);
and U22971 (N_22971,N_20245,N_20592);
nor U22972 (N_22972,N_21502,N_21034);
xor U22973 (N_22973,N_21856,N_21258);
nand U22974 (N_22974,N_20126,N_20858);
xor U22975 (N_22975,N_21001,N_20454);
nor U22976 (N_22976,N_20689,N_21187);
xor U22977 (N_22977,N_20167,N_20809);
or U22978 (N_22978,N_21038,N_21852);
nand U22979 (N_22979,N_20113,N_21125);
nor U22980 (N_22980,N_21107,N_20889);
and U22981 (N_22981,N_20744,N_21451);
and U22982 (N_22982,N_21894,N_20655);
nand U22983 (N_22983,N_21280,N_20213);
nand U22984 (N_22984,N_21627,N_21705);
xnor U22985 (N_22985,N_21652,N_20982);
or U22986 (N_22986,N_20404,N_21543);
and U22987 (N_22987,N_21295,N_20869);
and U22988 (N_22988,N_21300,N_20640);
xor U22989 (N_22989,N_21540,N_21709);
or U22990 (N_22990,N_21594,N_21963);
or U22991 (N_22991,N_21049,N_21292);
or U22992 (N_22992,N_21112,N_21275);
xor U22993 (N_22993,N_20136,N_20047);
nand U22994 (N_22994,N_20559,N_21356);
and U22995 (N_22995,N_21711,N_20473);
nand U22996 (N_22996,N_21993,N_21319);
nor U22997 (N_22997,N_21781,N_20321);
xnor U22998 (N_22998,N_20157,N_21593);
nand U22999 (N_22999,N_21526,N_21679);
and U23000 (N_23000,N_20999,N_20269);
nor U23001 (N_23001,N_20713,N_21713);
xor U23002 (N_23002,N_21973,N_20897);
nor U23003 (N_23003,N_20374,N_20957);
nand U23004 (N_23004,N_21273,N_21689);
nand U23005 (N_23005,N_20156,N_20918);
and U23006 (N_23006,N_20374,N_21684);
and U23007 (N_23007,N_21034,N_20094);
nand U23008 (N_23008,N_20242,N_20556);
and U23009 (N_23009,N_20198,N_21549);
nor U23010 (N_23010,N_20828,N_20303);
and U23011 (N_23011,N_20056,N_21613);
nand U23012 (N_23012,N_20917,N_21434);
nand U23013 (N_23013,N_20053,N_21832);
and U23014 (N_23014,N_20884,N_21821);
or U23015 (N_23015,N_21583,N_21362);
xnor U23016 (N_23016,N_20809,N_20030);
xnor U23017 (N_23017,N_20840,N_20019);
nor U23018 (N_23018,N_20689,N_21447);
nand U23019 (N_23019,N_21580,N_20922);
nand U23020 (N_23020,N_21505,N_20880);
or U23021 (N_23021,N_21985,N_21753);
nor U23022 (N_23022,N_21918,N_20140);
or U23023 (N_23023,N_21119,N_21986);
nor U23024 (N_23024,N_21732,N_20512);
and U23025 (N_23025,N_21954,N_21354);
nor U23026 (N_23026,N_21083,N_21838);
xnor U23027 (N_23027,N_21654,N_21772);
nand U23028 (N_23028,N_21177,N_21456);
xor U23029 (N_23029,N_20525,N_20801);
nand U23030 (N_23030,N_20023,N_20131);
nor U23031 (N_23031,N_21879,N_20925);
or U23032 (N_23032,N_21749,N_21591);
or U23033 (N_23033,N_20021,N_21292);
xor U23034 (N_23034,N_21457,N_21570);
and U23035 (N_23035,N_21881,N_21777);
xnor U23036 (N_23036,N_20413,N_21833);
xor U23037 (N_23037,N_21538,N_20743);
nor U23038 (N_23038,N_21447,N_20112);
or U23039 (N_23039,N_21214,N_20865);
xor U23040 (N_23040,N_21635,N_20780);
and U23041 (N_23041,N_21925,N_20204);
and U23042 (N_23042,N_21758,N_21292);
or U23043 (N_23043,N_20275,N_20654);
nand U23044 (N_23044,N_21038,N_20171);
nand U23045 (N_23045,N_21999,N_21199);
xnor U23046 (N_23046,N_20082,N_20213);
or U23047 (N_23047,N_20325,N_20117);
nor U23048 (N_23048,N_20517,N_20535);
xnor U23049 (N_23049,N_20343,N_20092);
nand U23050 (N_23050,N_20710,N_20692);
xor U23051 (N_23051,N_20687,N_20323);
xnor U23052 (N_23052,N_21362,N_20190);
nand U23053 (N_23053,N_21440,N_21066);
xor U23054 (N_23054,N_20147,N_21408);
and U23055 (N_23055,N_20593,N_21220);
nand U23056 (N_23056,N_21355,N_21048);
xnor U23057 (N_23057,N_20465,N_20674);
and U23058 (N_23058,N_20712,N_20877);
nand U23059 (N_23059,N_20165,N_20469);
xnor U23060 (N_23060,N_21579,N_21013);
nor U23061 (N_23061,N_21546,N_21146);
or U23062 (N_23062,N_20885,N_20451);
nand U23063 (N_23063,N_21811,N_21526);
nand U23064 (N_23064,N_20585,N_21666);
nor U23065 (N_23065,N_20205,N_20038);
or U23066 (N_23066,N_20977,N_20522);
nor U23067 (N_23067,N_20166,N_21527);
and U23068 (N_23068,N_20770,N_21182);
xnor U23069 (N_23069,N_20526,N_21902);
and U23070 (N_23070,N_21981,N_20133);
nor U23071 (N_23071,N_20753,N_21007);
xnor U23072 (N_23072,N_21772,N_20523);
nand U23073 (N_23073,N_20189,N_21060);
nor U23074 (N_23074,N_20440,N_20154);
nand U23075 (N_23075,N_21007,N_20389);
xor U23076 (N_23076,N_20570,N_21114);
nand U23077 (N_23077,N_21808,N_21983);
or U23078 (N_23078,N_21981,N_21736);
or U23079 (N_23079,N_20918,N_20043);
and U23080 (N_23080,N_20233,N_21649);
nand U23081 (N_23081,N_20160,N_21630);
nand U23082 (N_23082,N_20763,N_21656);
nor U23083 (N_23083,N_20425,N_21666);
nor U23084 (N_23084,N_20594,N_21986);
xor U23085 (N_23085,N_20769,N_21043);
nor U23086 (N_23086,N_21700,N_20088);
or U23087 (N_23087,N_21748,N_21688);
and U23088 (N_23088,N_20920,N_20738);
nand U23089 (N_23089,N_21387,N_21297);
xnor U23090 (N_23090,N_20612,N_21101);
and U23091 (N_23091,N_21301,N_20377);
and U23092 (N_23092,N_20646,N_20334);
nand U23093 (N_23093,N_21892,N_20023);
and U23094 (N_23094,N_20071,N_20973);
xnor U23095 (N_23095,N_20622,N_20086);
or U23096 (N_23096,N_20960,N_20328);
and U23097 (N_23097,N_20696,N_20674);
nand U23098 (N_23098,N_20429,N_21057);
nor U23099 (N_23099,N_20178,N_21234);
nor U23100 (N_23100,N_20949,N_21601);
nor U23101 (N_23101,N_20882,N_20649);
nand U23102 (N_23102,N_20075,N_20434);
nor U23103 (N_23103,N_20603,N_21209);
nor U23104 (N_23104,N_21365,N_20812);
nand U23105 (N_23105,N_21951,N_20558);
or U23106 (N_23106,N_21163,N_20100);
nand U23107 (N_23107,N_20597,N_21093);
xnor U23108 (N_23108,N_20951,N_20053);
nand U23109 (N_23109,N_20126,N_20613);
nand U23110 (N_23110,N_20785,N_20913);
nand U23111 (N_23111,N_21656,N_20061);
or U23112 (N_23112,N_20918,N_21005);
nand U23113 (N_23113,N_21578,N_21192);
and U23114 (N_23114,N_21549,N_20517);
and U23115 (N_23115,N_21427,N_21053);
nand U23116 (N_23116,N_20259,N_20414);
xnor U23117 (N_23117,N_20125,N_21395);
or U23118 (N_23118,N_21809,N_20667);
xor U23119 (N_23119,N_21003,N_21515);
nand U23120 (N_23120,N_21996,N_20589);
nor U23121 (N_23121,N_21736,N_21392);
nand U23122 (N_23122,N_20055,N_20791);
xnor U23123 (N_23123,N_20681,N_20307);
nor U23124 (N_23124,N_21116,N_20134);
and U23125 (N_23125,N_20122,N_21791);
and U23126 (N_23126,N_20999,N_20851);
and U23127 (N_23127,N_21058,N_20202);
xnor U23128 (N_23128,N_21539,N_20234);
and U23129 (N_23129,N_20768,N_21708);
xor U23130 (N_23130,N_21609,N_21844);
or U23131 (N_23131,N_21559,N_21264);
xor U23132 (N_23132,N_20625,N_20047);
or U23133 (N_23133,N_21771,N_20190);
xor U23134 (N_23134,N_20509,N_21703);
nand U23135 (N_23135,N_20373,N_20919);
xnor U23136 (N_23136,N_21089,N_21122);
nand U23137 (N_23137,N_21756,N_20833);
xor U23138 (N_23138,N_21027,N_21508);
nand U23139 (N_23139,N_20201,N_20003);
nand U23140 (N_23140,N_21351,N_20136);
nand U23141 (N_23141,N_20018,N_20453);
and U23142 (N_23142,N_21960,N_21513);
xor U23143 (N_23143,N_20156,N_21099);
nand U23144 (N_23144,N_21063,N_21702);
nor U23145 (N_23145,N_21111,N_21726);
or U23146 (N_23146,N_20144,N_21966);
nand U23147 (N_23147,N_20978,N_21688);
nor U23148 (N_23148,N_20687,N_20902);
nand U23149 (N_23149,N_20539,N_20144);
or U23150 (N_23150,N_21111,N_20275);
xor U23151 (N_23151,N_21980,N_21847);
nor U23152 (N_23152,N_21530,N_20738);
or U23153 (N_23153,N_21928,N_21911);
or U23154 (N_23154,N_20152,N_20516);
xor U23155 (N_23155,N_21893,N_20664);
nor U23156 (N_23156,N_20935,N_20424);
nand U23157 (N_23157,N_21685,N_21069);
nand U23158 (N_23158,N_20703,N_21357);
or U23159 (N_23159,N_20082,N_20851);
or U23160 (N_23160,N_21561,N_21692);
and U23161 (N_23161,N_21618,N_20112);
xnor U23162 (N_23162,N_21389,N_21094);
nand U23163 (N_23163,N_20358,N_20703);
xnor U23164 (N_23164,N_21267,N_20888);
and U23165 (N_23165,N_21221,N_21628);
xor U23166 (N_23166,N_20067,N_20496);
nor U23167 (N_23167,N_20719,N_20654);
and U23168 (N_23168,N_21924,N_21688);
nand U23169 (N_23169,N_20643,N_21995);
nand U23170 (N_23170,N_20123,N_20933);
or U23171 (N_23171,N_20547,N_20573);
nor U23172 (N_23172,N_20927,N_21287);
and U23173 (N_23173,N_21953,N_20041);
or U23174 (N_23174,N_21654,N_21927);
and U23175 (N_23175,N_20434,N_21848);
nand U23176 (N_23176,N_21217,N_21154);
nand U23177 (N_23177,N_20817,N_21400);
or U23178 (N_23178,N_20074,N_20315);
xor U23179 (N_23179,N_21514,N_20288);
and U23180 (N_23180,N_20926,N_20006);
and U23181 (N_23181,N_21408,N_21555);
nand U23182 (N_23182,N_21055,N_20269);
or U23183 (N_23183,N_20833,N_21388);
or U23184 (N_23184,N_21322,N_21564);
xnor U23185 (N_23185,N_20308,N_21681);
and U23186 (N_23186,N_20320,N_21988);
or U23187 (N_23187,N_20649,N_20044);
nand U23188 (N_23188,N_21176,N_20726);
nor U23189 (N_23189,N_21767,N_21944);
nor U23190 (N_23190,N_21249,N_21166);
nand U23191 (N_23191,N_20785,N_20012);
nand U23192 (N_23192,N_20487,N_21709);
xor U23193 (N_23193,N_20192,N_20220);
nand U23194 (N_23194,N_21653,N_21361);
nand U23195 (N_23195,N_21705,N_20180);
or U23196 (N_23196,N_20481,N_21438);
or U23197 (N_23197,N_21631,N_20486);
or U23198 (N_23198,N_20419,N_21596);
xor U23199 (N_23199,N_20483,N_21653);
xnor U23200 (N_23200,N_20183,N_20531);
nand U23201 (N_23201,N_21433,N_21797);
and U23202 (N_23202,N_20321,N_21815);
and U23203 (N_23203,N_20911,N_21245);
nor U23204 (N_23204,N_20571,N_21306);
xor U23205 (N_23205,N_21615,N_21627);
nand U23206 (N_23206,N_21806,N_20555);
nor U23207 (N_23207,N_21261,N_21201);
or U23208 (N_23208,N_20462,N_21782);
nand U23209 (N_23209,N_20801,N_21572);
xor U23210 (N_23210,N_20457,N_20546);
and U23211 (N_23211,N_20270,N_21742);
and U23212 (N_23212,N_20290,N_20112);
xor U23213 (N_23213,N_21863,N_21137);
and U23214 (N_23214,N_20093,N_20166);
nor U23215 (N_23215,N_20550,N_20108);
nor U23216 (N_23216,N_21188,N_21882);
nand U23217 (N_23217,N_20478,N_20866);
or U23218 (N_23218,N_20689,N_20574);
and U23219 (N_23219,N_20002,N_20559);
xnor U23220 (N_23220,N_21865,N_21068);
and U23221 (N_23221,N_20229,N_21306);
and U23222 (N_23222,N_21679,N_20676);
xor U23223 (N_23223,N_20749,N_20897);
xor U23224 (N_23224,N_20047,N_20697);
and U23225 (N_23225,N_21132,N_20005);
nand U23226 (N_23226,N_21132,N_20120);
nand U23227 (N_23227,N_20630,N_21015);
and U23228 (N_23228,N_20018,N_21814);
and U23229 (N_23229,N_20061,N_20290);
nand U23230 (N_23230,N_21596,N_21300);
xnor U23231 (N_23231,N_20038,N_21519);
xnor U23232 (N_23232,N_20568,N_21046);
xor U23233 (N_23233,N_20356,N_21963);
xor U23234 (N_23234,N_21728,N_21149);
nand U23235 (N_23235,N_21140,N_20798);
xnor U23236 (N_23236,N_20434,N_21415);
or U23237 (N_23237,N_21300,N_21998);
nand U23238 (N_23238,N_21969,N_21457);
and U23239 (N_23239,N_20979,N_20975);
xnor U23240 (N_23240,N_20059,N_21881);
or U23241 (N_23241,N_21263,N_20658);
nand U23242 (N_23242,N_20802,N_21345);
xnor U23243 (N_23243,N_20067,N_20531);
or U23244 (N_23244,N_20906,N_20026);
and U23245 (N_23245,N_21153,N_21963);
xnor U23246 (N_23246,N_20737,N_21677);
xor U23247 (N_23247,N_20973,N_20400);
xor U23248 (N_23248,N_20496,N_20227);
and U23249 (N_23249,N_20635,N_21510);
xor U23250 (N_23250,N_21890,N_20192);
nor U23251 (N_23251,N_20193,N_21250);
or U23252 (N_23252,N_21778,N_20760);
or U23253 (N_23253,N_20476,N_21081);
nand U23254 (N_23254,N_21647,N_20245);
and U23255 (N_23255,N_20721,N_20500);
and U23256 (N_23256,N_20871,N_20910);
and U23257 (N_23257,N_21685,N_20438);
or U23258 (N_23258,N_21461,N_21295);
nor U23259 (N_23259,N_20291,N_20929);
or U23260 (N_23260,N_21044,N_21424);
nor U23261 (N_23261,N_21387,N_20148);
xnor U23262 (N_23262,N_21003,N_20665);
xor U23263 (N_23263,N_20800,N_20358);
nand U23264 (N_23264,N_20383,N_21966);
nor U23265 (N_23265,N_20800,N_21490);
nor U23266 (N_23266,N_21828,N_20656);
nor U23267 (N_23267,N_21698,N_21918);
nand U23268 (N_23268,N_21942,N_21543);
nor U23269 (N_23269,N_21614,N_21353);
and U23270 (N_23270,N_21487,N_20510);
or U23271 (N_23271,N_20097,N_20282);
and U23272 (N_23272,N_21061,N_21685);
nor U23273 (N_23273,N_20348,N_20263);
or U23274 (N_23274,N_20348,N_21475);
and U23275 (N_23275,N_21525,N_21002);
xor U23276 (N_23276,N_20814,N_21313);
or U23277 (N_23277,N_20422,N_21524);
xnor U23278 (N_23278,N_20534,N_21544);
and U23279 (N_23279,N_20074,N_21140);
nor U23280 (N_23280,N_21016,N_21317);
or U23281 (N_23281,N_21382,N_20743);
nor U23282 (N_23282,N_20292,N_20001);
and U23283 (N_23283,N_21662,N_21668);
and U23284 (N_23284,N_21245,N_20559);
and U23285 (N_23285,N_21576,N_21464);
and U23286 (N_23286,N_21248,N_21288);
or U23287 (N_23287,N_21761,N_21583);
nor U23288 (N_23288,N_21895,N_21942);
nor U23289 (N_23289,N_20846,N_20083);
or U23290 (N_23290,N_21745,N_20602);
and U23291 (N_23291,N_21585,N_21622);
and U23292 (N_23292,N_21043,N_21514);
nand U23293 (N_23293,N_20200,N_21020);
nand U23294 (N_23294,N_20551,N_20961);
xor U23295 (N_23295,N_21922,N_20591);
xnor U23296 (N_23296,N_21091,N_20097);
xor U23297 (N_23297,N_20302,N_21965);
nand U23298 (N_23298,N_21613,N_20018);
xor U23299 (N_23299,N_21667,N_21558);
or U23300 (N_23300,N_20870,N_21293);
nand U23301 (N_23301,N_20769,N_21407);
nand U23302 (N_23302,N_21385,N_20951);
nor U23303 (N_23303,N_21388,N_21510);
nand U23304 (N_23304,N_20425,N_20581);
nor U23305 (N_23305,N_20603,N_20450);
and U23306 (N_23306,N_20846,N_20575);
and U23307 (N_23307,N_20984,N_20758);
or U23308 (N_23308,N_20998,N_21214);
nor U23309 (N_23309,N_20675,N_20162);
nand U23310 (N_23310,N_21576,N_20995);
and U23311 (N_23311,N_20464,N_21029);
xor U23312 (N_23312,N_20350,N_20065);
and U23313 (N_23313,N_20638,N_21742);
and U23314 (N_23314,N_20690,N_20567);
xor U23315 (N_23315,N_21088,N_20461);
nor U23316 (N_23316,N_20582,N_20267);
and U23317 (N_23317,N_20826,N_21698);
nand U23318 (N_23318,N_20735,N_21886);
nor U23319 (N_23319,N_21788,N_20071);
nand U23320 (N_23320,N_20422,N_21519);
nor U23321 (N_23321,N_20016,N_21399);
and U23322 (N_23322,N_20105,N_21876);
or U23323 (N_23323,N_20099,N_21771);
nor U23324 (N_23324,N_20992,N_21129);
xor U23325 (N_23325,N_20627,N_20093);
nand U23326 (N_23326,N_20111,N_20861);
nand U23327 (N_23327,N_21487,N_21375);
nor U23328 (N_23328,N_20194,N_21803);
and U23329 (N_23329,N_20612,N_20154);
nand U23330 (N_23330,N_21826,N_21957);
nand U23331 (N_23331,N_20998,N_20359);
xnor U23332 (N_23332,N_21568,N_20233);
xor U23333 (N_23333,N_21767,N_21641);
xor U23334 (N_23334,N_20997,N_20413);
nand U23335 (N_23335,N_21086,N_21175);
or U23336 (N_23336,N_20726,N_20217);
nand U23337 (N_23337,N_21835,N_20464);
and U23338 (N_23338,N_20162,N_21295);
nand U23339 (N_23339,N_21093,N_20567);
xnor U23340 (N_23340,N_20761,N_21237);
xor U23341 (N_23341,N_21647,N_20169);
and U23342 (N_23342,N_21303,N_21957);
and U23343 (N_23343,N_20580,N_21036);
and U23344 (N_23344,N_20405,N_20648);
nor U23345 (N_23345,N_21802,N_20093);
nor U23346 (N_23346,N_21179,N_20264);
and U23347 (N_23347,N_20754,N_21659);
nand U23348 (N_23348,N_20716,N_20434);
nand U23349 (N_23349,N_20559,N_21661);
and U23350 (N_23350,N_20383,N_20656);
or U23351 (N_23351,N_21657,N_21264);
nand U23352 (N_23352,N_20277,N_21459);
xor U23353 (N_23353,N_20196,N_21270);
nand U23354 (N_23354,N_21430,N_21101);
xnor U23355 (N_23355,N_20704,N_20497);
or U23356 (N_23356,N_21999,N_20051);
or U23357 (N_23357,N_20548,N_20045);
nand U23358 (N_23358,N_20155,N_20712);
xnor U23359 (N_23359,N_21565,N_21296);
xor U23360 (N_23360,N_20997,N_20781);
xor U23361 (N_23361,N_21707,N_21033);
or U23362 (N_23362,N_21425,N_20634);
nor U23363 (N_23363,N_20275,N_20044);
xnor U23364 (N_23364,N_21794,N_20337);
or U23365 (N_23365,N_20240,N_21263);
nand U23366 (N_23366,N_21527,N_20162);
xor U23367 (N_23367,N_20091,N_20702);
xor U23368 (N_23368,N_20590,N_21431);
xnor U23369 (N_23369,N_20454,N_20467);
or U23370 (N_23370,N_20737,N_21490);
xor U23371 (N_23371,N_20688,N_21925);
nor U23372 (N_23372,N_21705,N_20328);
xnor U23373 (N_23373,N_21441,N_21465);
nor U23374 (N_23374,N_21179,N_20127);
or U23375 (N_23375,N_20379,N_20054);
xor U23376 (N_23376,N_21878,N_21796);
or U23377 (N_23377,N_20045,N_20066);
and U23378 (N_23378,N_20490,N_21722);
nor U23379 (N_23379,N_21163,N_20829);
xnor U23380 (N_23380,N_21519,N_20230);
nor U23381 (N_23381,N_21816,N_21427);
nand U23382 (N_23382,N_21453,N_21351);
nor U23383 (N_23383,N_21790,N_20720);
and U23384 (N_23384,N_20950,N_21778);
nor U23385 (N_23385,N_20741,N_20204);
and U23386 (N_23386,N_21832,N_21923);
nor U23387 (N_23387,N_20676,N_20006);
xor U23388 (N_23388,N_21620,N_21525);
and U23389 (N_23389,N_20082,N_20221);
xor U23390 (N_23390,N_20540,N_20631);
xor U23391 (N_23391,N_20902,N_21858);
nand U23392 (N_23392,N_20117,N_21359);
xor U23393 (N_23393,N_21680,N_21401);
and U23394 (N_23394,N_21490,N_21781);
xor U23395 (N_23395,N_21866,N_20202);
xnor U23396 (N_23396,N_21109,N_20222);
or U23397 (N_23397,N_20459,N_21972);
or U23398 (N_23398,N_21915,N_21844);
xnor U23399 (N_23399,N_20202,N_21780);
nand U23400 (N_23400,N_20210,N_21378);
or U23401 (N_23401,N_20695,N_21439);
nand U23402 (N_23402,N_21593,N_21672);
nand U23403 (N_23403,N_21582,N_21847);
xor U23404 (N_23404,N_21630,N_21474);
and U23405 (N_23405,N_20292,N_21526);
nor U23406 (N_23406,N_21040,N_21425);
and U23407 (N_23407,N_20698,N_20721);
xor U23408 (N_23408,N_20889,N_21739);
or U23409 (N_23409,N_21261,N_20552);
nor U23410 (N_23410,N_21807,N_20871);
xnor U23411 (N_23411,N_20996,N_20770);
nor U23412 (N_23412,N_20013,N_21219);
nor U23413 (N_23413,N_21517,N_21132);
or U23414 (N_23414,N_21358,N_20302);
or U23415 (N_23415,N_20716,N_20832);
nand U23416 (N_23416,N_20736,N_21237);
nor U23417 (N_23417,N_21885,N_20965);
or U23418 (N_23418,N_20572,N_20056);
and U23419 (N_23419,N_21329,N_21759);
nand U23420 (N_23420,N_20924,N_21431);
nor U23421 (N_23421,N_20312,N_20618);
xnor U23422 (N_23422,N_20573,N_20178);
nor U23423 (N_23423,N_20271,N_20622);
or U23424 (N_23424,N_20143,N_21135);
and U23425 (N_23425,N_20556,N_20847);
and U23426 (N_23426,N_21909,N_21091);
or U23427 (N_23427,N_21429,N_21083);
xnor U23428 (N_23428,N_20418,N_21996);
nand U23429 (N_23429,N_20434,N_20948);
and U23430 (N_23430,N_21724,N_21665);
xnor U23431 (N_23431,N_20732,N_20220);
nor U23432 (N_23432,N_21713,N_20179);
nand U23433 (N_23433,N_20971,N_21899);
nand U23434 (N_23434,N_20311,N_20458);
nor U23435 (N_23435,N_21932,N_20493);
and U23436 (N_23436,N_21630,N_21293);
xor U23437 (N_23437,N_20854,N_20614);
xnor U23438 (N_23438,N_20170,N_21178);
and U23439 (N_23439,N_21890,N_21650);
nor U23440 (N_23440,N_21878,N_20006);
nor U23441 (N_23441,N_21965,N_21923);
xor U23442 (N_23442,N_21250,N_21426);
or U23443 (N_23443,N_21317,N_21123);
and U23444 (N_23444,N_21034,N_20751);
or U23445 (N_23445,N_21008,N_21507);
nand U23446 (N_23446,N_20207,N_20851);
xnor U23447 (N_23447,N_20185,N_20791);
and U23448 (N_23448,N_21494,N_20963);
and U23449 (N_23449,N_21170,N_20632);
nor U23450 (N_23450,N_20177,N_21869);
or U23451 (N_23451,N_20862,N_21133);
or U23452 (N_23452,N_21626,N_21385);
and U23453 (N_23453,N_20010,N_21577);
nor U23454 (N_23454,N_21430,N_20107);
and U23455 (N_23455,N_21998,N_20892);
and U23456 (N_23456,N_20282,N_21060);
xnor U23457 (N_23457,N_20560,N_20677);
and U23458 (N_23458,N_21027,N_20322);
nand U23459 (N_23459,N_21925,N_20270);
xor U23460 (N_23460,N_20668,N_20489);
and U23461 (N_23461,N_21967,N_21389);
or U23462 (N_23462,N_21634,N_20918);
and U23463 (N_23463,N_21968,N_21337);
nand U23464 (N_23464,N_21675,N_20306);
xnor U23465 (N_23465,N_20681,N_21423);
nor U23466 (N_23466,N_20824,N_21159);
nor U23467 (N_23467,N_21259,N_21901);
and U23468 (N_23468,N_21115,N_21930);
xor U23469 (N_23469,N_21292,N_21506);
nor U23470 (N_23470,N_20021,N_21560);
or U23471 (N_23471,N_20326,N_21102);
nor U23472 (N_23472,N_20089,N_20620);
and U23473 (N_23473,N_20896,N_21723);
nand U23474 (N_23474,N_21728,N_21118);
nor U23475 (N_23475,N_20895,N_20517);
xnor U23476 (N_23476,N_20199,N_20335);
or U23477 (N_23477,N_20449,N_20611);
or U23478 (N_23478,N_20927,N_21870);
or U23479 (N_23479,N_20763,N_21024);
and U23480 (N_23480,N_21741,N_20130);
nor U23481 (N_23481,N_20484,N_21935);
xnor U23482 (N_23482,N_21715,N_20445);
nand U23483 (N_23483,N_20322,N_21531);
and U23484 (N_23484,N_21675,N_20908);
nor U23485 (N_23485,N_21148,N_20245);
and U23486 (N_23486,N_20802,N_20012);
nor U23487 (N_23487,N_21021,N_20788);
xnor U23488 (N_23488,N_20052,N_21734);
xnor U23489 (N_23489,N_20586,N_20105);
and U23490 (N_23490,N_20949,N_20562);
nand U23491 (N_23491,N_20238,N_20224);
nor U23492 (N_23492,N_20476,N_21920);
and U23493 (N_23493,N_20807,N_20751);
or U23494 (N_23494,N_21720,N_20262);
or U23495 (N_23495,N_21035,N_21779);
nor U23496 (N_23496,N_20356,N_21065);
or U23497 (N_23497,N_21510,N_20831);
xor U23498 (N_23498,N_21642,N_21628);
and U23499 (N_23499,N_21589,N_20228);
and U23500 (N_23500,N_20793,N_20939);
and U23501 (N_23501,N_21446,N_20295);
nand U23502 (N_23502,N_20486,N_20728);
or U23503 (N_23503,N_20732,N_21267);
or U23504 (N_23504,N_20284,N_21702);
xor U23505 (N_23505,N_20670,N_21646);
and U23506 (N_23506,N_20054,N_21943);
nor U23507 (N_23507,N_20187,N_20915);
or U23508 (N_23508,N_21362,N_21899);
nand U23509 (N_23509,N_20125,N_20300);
nor U23510 (N_23510,N_21222,N_21712);
xnor U23511 (N_23511,N_21611,N_20692);
or U23512 (N_23512,N_20740,N_21701);
nand U23513 (N_23513,N_20943,N_21320);
or U23514 (N_23514,N_20753,N_20528);
xor U23515 (N_23515,N_20282,N_20486);
xor U23516 (N_23516,N_20444,N_21291);
or U23517 (N_23517,N_20874,N_20068);
nor U23518 (N_23518,N_21731,N_21175);
nor U23519 (N_23519,N_20248,N_20466);
and U23520 (N_23520,N_21905,N_21796);
nor U23521 (N_23521,N_21613,N_20137);
and U23522 (N_23522,N_21947,N_20798);
and U23523 (N_23523,N_21943,N_21297);
nand U23524 (N_23524,N_20757,N_20956);
nand U23525 (N_23525,N_20633,N_21166);
nor U23526 (N_23526,N_20755,N_21480);
xor U23527 (N_23527,N_20819,N_20466);
or U23528 (N_23528,N_21862,N_21029);
nand U23529 (N_23529,N_21671,N_20842);
nand U23530 (N_23530,N_20215,N_21412);
and U23531 (N_23531,N_21845,N_21993);
or U23532 (N_23532,N_20756,N_20096);
nor U23533 (N_23533,N_21691,N_21555);
nor U23534 (N_23534,N_21930,N_21951);
or U23535 (N_23535,N_21610,N_20558);
xnor U23536 (N_23536,N_20639,N_21894);
xor U23537 (N_23537,N_20763,N_20247);
xnor U23538 (N_23538,N_20554,N_20205);
and U23539 (N_23539,N_20155,N_21777);
nor U23540 (N_23540,N_21259,N_21162);
and U23541 (N_23541,N_20741,N_21972);
nand U23542 (N_23542,N_20814,N_21551);
nand U23543 (N_23543,N_21904,N_21357);
or U23544 (N_23544,N_21847,N_21130);
xnor U23545 (N_23545,N_21984,N_20693);
nand U23546 (N_23546,N_21043,N_21408);
nor U23547 (N_23547,N_20250,N_20935);
nand U23548 (N_23548,N_21131,N_21759);
xnor U23549 (N_23549,N_20186,N_21385);
nor U23550 (N_23550,N_21648,N_21261);
nor U23551 (N_23551,N_20652,N_20194);
and U23552 (N_23552,N_20634,N_21392);
nand U23553 (N_23553,N_20717,N_21246);
xor U23554 (N_23554,N_20835,N_20246);
xor U23555 (N_23555,N_21386,N_20253);
and U23556 (N_23556,N_21168,N_20043);
nor U23557 (N_23557,N_20097,N_20270);
or U23558 (N_23558,N_21381,N_21974);
xor U23559 (N_23559,N_21551,N_20295);
or U23560 (N_23560,N_21721,N_21054);
xnor U23561 (N_23561,N_21985,N_20906);
nand U23562 (N_23562,N_21437,N_21940);
nor U23563 (N_23563,N_21602,N_21737);
and U23564 (N_23564,N_20067,N_20150);
and U23565 (N_23565,N_20597,N_21067);
or U23566 (N_23566,N_21426,N_21527);
nand U23567 (N_23567,N_20904,N_21888);
nor U23568 (N_23568,N_21222,N_20685);
nor U23569 (N_23569,N_21549,N_20261);
xnor U23570 (N_23570,N_20844,N_21209);
or U23571 (N_23571,N_21069,N_21782);
nand U23572 (N_23572,N_20174,N_20238);
nor U23573 (N_23573,N_20680,N_20172);
nand U23574 (N_23574,N_21842,N_21249);
nor U23575 (N_23575,N_21898,N_20293);
nor U23576 (N_23576,N_21790,N_20462);
and U23577 (N_23577,N_20011,N_20313);
nand U23578 (N_23578,N_21117,N_20466);
xor U23579 (N_23579,N_20882,N_21619);
nor U23580 (N_23580,N_21645,N_21669);
nand U23581 (N_23581,N_20567,N_20450);
or U23582 (N_23582,N_20094,N_21657);
or U23583 (N_23583,N_21275,N_20087);
nand U23584 (N_23584,N_20652,N_20241);
and U23585 (N_23585,N_21679,N_21574);
nand U23586 (N_23586,N_21541,N_20702);
nand U23587 (N_23587,N_20366,N_21952);
nor U23588 (N_23588,N_21936,N_20660);
xor U23589 (N_23589,N_21740,N_20592);
or U23590 (N_23590,N_21441,N_20695);
nor U23591 (N_23591,N_21725,N_21463);
nor U23592 (N_23592,N_20604,N_20765);
nand U23593 (N_23593,N_21778,N_21933);
nand U23594 (N_23594,N_21305,N_21694);
and U23595 (N_23595,N_21331,N_21009);
and U23596 (N_23596,N_20302,N_20257);
nand U23597 (N_23597,N_20447,N_21939);
or U23598 (N_23598,N_21685,N_21145);
xor U23599 (N_23599,N_20612,N_20214);
xnor U23600 (N_23600,N_21540,N_21755);
or U23601 (N_23601,N_21063,N_21733);
nand U23602 (N_23602,N_20063,N_21620);
or U23603 (N_23603,N_21139,N_20672);
and U23604 (N_23604,N_21816,N_21123);
nand U23605 (N_23605,N_20850,N_20001);
and U23606 (N_23606,N_21094,N_20700);
nor U23607 (N_23607,N_21115,N_21080);
nand U23608 (N_23608,N_20241,N_20556);
or U23609 (N_23609,N_20652,N_21638);
or U23610 (N_23610,N_20565,N_20488);
or U23611 (N_23611,N_21961,N_21009);
xnor U23612 (N_23612,N_21232,N_20537);
nand U23613 (N_23613,N_20851,N_20357);
nor U23614 (N_23614,N_20555,N_21849);
xnor U23615 (N_23615,N_21766,N_20587);
xnor U23616 (N_23616,N_20841,N_20517);
or U23617 (N_23617,N_20447,N_21547);
xnor U23618 (N_23618,N_21722,N_21136);
and U23619 (N_23619,N_21357,N_20822);
nand U23620 (N_23620,N_20918,N_21693);
nand U23621 (N_23621,N_20206,N_21516);
and U23622 (N_23622,N_20650,N_20901);
nand U23623 (N_23623,N_21718,N_21885);
or U23624 (N_23624,N_20566,N_20976);
xor U23625 (N_23625,N_20949,N_21678);
nor U23626 (N_23626,N_21132,N_21927);
nor U23627 (N_23627,N_20317,N_20147);
xor U23628 (N_23628,N_20685,N_21491);
nand U23629 (N_23629,N_20931,N_20929);
nand U23630 (N_23630,N_20897,N_21966);
nand U23631 (N_23631,N_21067,N_21035);
or U23632 (N_23632,N_21301,N_21296);
and U23633 (N_23633,N_20159,N_20627);
nand U23634 (N_23634,N_21146,N_20277);
and U23635 (N_23635,N_20564,N_21923);
nand U23636 (N_23636,N_21010,N_20398);
or U23637 (N_23637,N_21427,N_21923);
and U23638 (N_23638,N_20004,N_21019);
nand U23639 (N_23639,N_20499,N_20763);
or U23640 (N_23640,N_21996,N_21484);
xor U23641 (N_23641,N_21022,N_21256);
and U23642 (N_23642,N_21959,N_20821);
or U23643 (N_23643,N_20171,N_21916);
xor U23644 (N_23644,N_20028,N_20057);
xnor U23645 (N_23645,N_20613,N_21430);
nand U23646 (N_23646,N_21674,N_20386);
nor U23647 (N_23647,N_20493,N_20687);
and U23648 (N_23648,N_20438,N_20026);
xnor U23649 (N_23649,N_20150,N_21071);
or U23650 (N_23650,N_20058,N_20555);
and U23651 (N_23651,N_20356,N_20780);
or U23652 (N_23652,N_20229,N_21740);
nand U23653 (N_23653,N_21228,N_20956);
nand U23654 (N_23654,N_20187,N_20467);
or U23655 (N_23655,N_20368,N_20086);
or U23656 (N_23656,N_21486,N_21471);
and U23657 (N_23657,N_21646,N_21260);
nand U23658 (N_23658,N_20456,N_20615);
and U23659 (N_23659,N_21852,N_20151);
xor U23660 (N_23660,N_21099,N_21045);
and U23661 (N_23661,N_21078,N_20338);
nor U23662 (N_23662,N_21731,N_21003);
nand U23663 (N_23663,N_20817,N_20671);
or U23664 (N_23664,N_20827,N_20716);
nor U23665 (N_23665,N_20838,N_20045);
or U23666 (N_23666,N_20391,N_21255);
xnor U23667 (N_23667,N_20137,N_20493);
or U23668 (N_23668,N_20965,N_21303);
xor U23669 (N_23669,N_21132,N_21416);
or U23670 (N_23670,N_21085,N_21727);
nand U23671 (N_23671,N_21228,N_20243);
nand U23672 (N_23672,N_20597,N_20760);
nor U23673 (N_23673,N_21729,N_21460);
nand U23674 (N_23674,N_20671,N_20288);
nor U23675 (N_23675,N_20766,N_21667);
nand U23676 (N_23676,N_21181,N_21066);
and U23677 (N_23677,N_20001,N_20587);
and U23678 (N_23678,N_21349,N_20515);
and U23679 (N_23679,N_20345,N_21784);
nand U23680 (N_23680,N_20989,N_20237);
nand U23681 (N_23681,N_20166,N_21043);
xor U23682 (N_23682,N_21190,N_20853);
nand U23683 (N_23683,N_20103,N_21461);
nor U23684 (N_23684,N_21573,N_20727);
xor U23685 (N_23685,N_20680,N_21551);
and U23686 (N_23686,N_20689,N_21457);
nor U23687 (N_23687,N_21910,N_21633);
and U23688 (N_23688,N_20515,N_21107);
or U23689 (N_23689,N_20873,N_20847);
xor U23690 (N_23690,N_21261,N_21374);
and U23691 (N_23691,N_20917,N_20316);
nor U23692 (N_23692,N_20401,N_21314);
and U23693 (N_23693,N_21656,N_20993);
and U23694 (N_23694,N_21056,N_20170);
or U23695 (N_23695,N_21410,N_21448);
nor U23696 (N_23696,N_21528,N_21853);
nor U23697 (N_23697,N_20089,N_21972);
nor U23698 (N_23698,N_21716,N_21841);
or U23699 (N_23699,N_20766,N_20936);
or U23700 (N_23700,N_21380,N_20521);
nand U23701 (N_23701,N_20277,N_20816);
nor U23702 (N_23702,N_20656,N_21671);
nor U23703 (N_23703,N_20978,N_20256);
nor U23704 (N_23704,N_20029,N_20384);
or U23705 (N_23705,N_21417,N_20029);
nand U23706 (N_23706,N_21860,N_21081);
nor U23707 (N_23707,N_21147,N_21042);
or U23708 (N_23708,N_21813,N_20008);
nand U23709 (N_23709,N_21191,N_20920);
or U23710 (N_23710,N_21988,N_21566);
or U23711 (N_23711,N_20436,N_21636);
nor U23712 (N_23712,N_21444,N_20678);
nor U23713 (N_23713,N_21507,N_21136);
nand U23714 (N_23714,N_21847,N_21299);
nor U23715 (N_23715,N_21276,N_21805);
nor U23716 (N_23716,N_20077,N_21823);
nand U23717 (N_23717,N_20793,N_21709);
nand U23718 (N_23718,N_21350,N_20675);
nor U23719 (N_23719,N_21261,N_20230);
and U23720 (N_23720,N_21354,N_21025);
nor U23721 (N_23721,N_20755,N_20099);
or U23722 (N_23722,N_20302,N_21806);
or U23723 (N_23723,N_21857,N_21581);
or U23724 (N_23724,N_21448,N_20370);
nor U23725 (N_23725,N_20676,N_20090);
nor U23726 (N_23726,N_20596,N_20219);
xnor U23727 (N_23727,N_21669,N_21633);
xnor U23728 (N_23728,N_21872,N_21669);
or U23729 (N_23729,N_20363,N_21052);
nand U23730 (N_23730,N_20034,N_20915);
and U23731 (N_23731,N_20156,N_21491);
nor U23732 (N_23732,N_20963,N_20815);
xor U23733 (N_23733,N_20026,N_20282);
and U23734 (N_23734,N_20792,N_20929);
or U23735 (N_23735,N_21198,N_20129);
or U23736 (N_23736,N_20245,N_21459);
nor U23737 (N_23737,N_20124,N_20411);
and U23738 (N_23738,N_21735,N_20876);
and U23739 (N_23739,N_20459,N_20579);
nand U23740 (N_23740,N_20422,N_21019);
or U23741 (N_23741,N_20559,N_20042);
or U23742 (N_23742,N_20292,N_21436);
or U23743 (N_23743,N_21665,N_21401);
nand U23744 (N_23744,N_21555,N_21675);
or U23745 (N_23745,N_20906,N_21003);
nor U23746 (N_23746,N_21389,N_20797);
or U23747 (N_23747,N_21752,N_21086);
xnor U23748 (N_23748,N_20948,N_21489);
nand U23749 (N_23749,N_21487,N_20529);
and U23750 (N_23750,N_20164,N_21825);
nor U23751 (N_23751,N_21122,N_21188);
or U23752 (N_23752,N_21196,N_21351);
nand U23753 (N_23753,N_20897,N_21240);
nand U23754 (N_23754,N_20431,N_21106);
or U23755 (N_23755,N_20215,N_20305);
xor U23756 (N_23756,N_20445,N_21392);
xnor U23757 (N_23757,N_21139,N_20205);
and U23758 (N_23758,N_21103,N_20785);
nand U23759 (N_23759,N_21043,N_21172);
or U23760 (N_23760,N_20570,N_21594);
nand U23761 (N_23761,N_20247,N_21260);
xor U23762 (N_23762,N_20494,N_20980);
or U23763 (N_23763,N_21066,N_21546);
nand U23764 (N_23764,N_21729,N_20986);
xnor U23765 (N_23765,N_20790,N_21410);
xnor U23766 (N_23766,N_21259,N_21262);
or U23767 (N_23767,N_21795,N_20653);
or U23768 (N_23768,N_20947,N_21232);
xor U23769 (N_23769,N_20276,N_20274);
nor U23770 (N_23770,N_21074,N_20935);
nand U23771 (N_23771,N_20904,N_20974);
or U23772 (N_23772,N_21184,N_20411);
or U23773 (N_23773,N_21532,N_20294);
nor U23774 (N_23774,N_20845,N_20575);
or U23775 (N_23775,N_21313,N_21141);
nor U23776 (N_23776,N_20745,N_21297);
nor U23777 (N_23777,N_20586,N_20175);
and U23778 (N_23778,N_20855,N_20614);
and U23779 (N_23779,N_20408,N_20570);
nor U23780 (N_23780,N_21638,N_21926);
and U23781 (N_23781,N_21762,N_20167);
nand U23782 (N_23782,N_20066,N_20844);
and U23783 (N_23783,N_20634,N_20656);
or U23784 (N_23784,N_21645,N_21563);
xor U23785 (N_23785,N_21272,N_21830);
nand U23786 (N_23786,N_20683,N_20365);
and U23787 (N_23787,N_20059,N_20836);
and U23788 (N_23788,N_21270,N_21329);
xor U23789 (N_23789,N_20719,N_20160);
or U23790 (N_23790,N_21948,N_21112);
nor U23791 (N_23791,N_20708,N_21925);
nand U23792 (N_23792,N_20159,N_21334);
nand U23793 (N_23793,N_20396,N_21973);
nor U23794 (N_23794,N_20982,N_21439);
or U23795 (N_23795,N_21038,N_21514);
or U23796 (N_23796,N_21593,N_20747);
or U23797 (N_23797,N_20124,N_20645);
xnor U23798 (N_23798,N_21442,N_20818);
nor U23799 (N_23799,N_21788,N_20397);
nor U23800 (N_23800,N_20761,N_20229);
or U23801 (N_23801,N_20383,N_21543);
nor U23802 (N_23802,N_20533,N_20834);
nor U23803 (N_23803,N_21115,N_20869);
and U23804 (N_23804,N_20366,N_21157);
xor U23805 (N_23805,N_20515,N_20824);
xor U23806 (N_23806,N_21033,N_20232);
or U23807 (N_23807,N_21263,N_20106);
and U23808 (N_23808,N_20135,N_20214);
or U23809 (N_23809,N_21056,N_21244);
and U23810 (N_23810,N_21655,N_21956);
nor U23811 (N_23811,N_20552,N_20195);
nor U23812 (N_23812,N_21044,N_21687);
or U23813 (N_23813,N_21777,N_20876);
nor U23814 (N_23814,N_21182,N_20447);
nand U23815 (N_23815,N_20348,N_21206);
nand U23816 (N_23816,N_21913,N_21728);
or U23817 (N_23817,N_21217,N_20619);
xor U23818 (N_23818,N_21414,N_20137);
nand U23819 (N_23819,N_20950,N_20804);
nor U23820 (N_23820,N_20517,N_21410);
nor U23821 (N_23821,N_21296,N_20079);
xor U23822 (N_23822,N_20842,N_21504);
or U23823 (N_23823,N_21066,N_21052);
xor U23824 (N_23824,N_21910,N_20982);
and U23825 (N_23825,N_20491,N_21034);
and U23826 (N_23826,N_21768,N_21376);
nand U23827 (N_23827,N_20847,N_21308);
or U23828 (N_23828,N_21819,N_20233);
nand U23829 (N_23829,N_21600,N_20785);
or U23830 (N_23830,N_20686,N_20754);
or U23831 (N_23831,N_20423,N_20752);
and U23832 (N_23832,N_20551,N_20199);
or U23833 (N_23833,N_21501,N_20896);
xnor U23834 (N_23834,N_20238,N_20503);
nor U23835 (N_23835,N_20072,N_21611);
xnor U23836 (N_23836,N_20351,N_21642);
nor U23837 (N_23837,N_21451,N_20189);
and U23838 (N_23838,N_20203,N_21145);
or U23839 (N_23839,N_20440,N_20132);
nand U23840 (N_23840,N_20880,N_21215);
or U23841 (N_23841,N_21148,N_21285);
xor U23842 (N_23842,N_20329,N_21852);
xor U23843 (N_23843,N_20964,N_20682);
or U23844 (N_23844,N_20921,N_20485);
and U23845 (N_23845,N_20174,N_20858);
or U23846 (N_23846,N_20346,N_21970);
nor U23847 (N_23847,N_21486,N_20975);
and U23848 (N_23848,N_20583,N_20216);
and U23849 (N_23849,N_20083,N_20410);
and U23850 (N_23850,N_20124,N_21408);
nand U23851 (N_23851,N_20000,N_20318);
xnor U23852 (N_23852,N_20372,N_20857);
or U23853 (N_23853,N_21890,N_21824);
nor U23854 (N_23854,N_20612,N_21421);
nor U23855 (N_23855,N_21210,N_21989);
nor U23856 (N_23856,N_21974,N_20448);
and U23857 (N_23857,N_21430,N_21428);
nor U23858 (N_23858,N_20732,N_20051);
xor U23859 (N_23859,N_21913,N_20782);
xor U23860 (N_23860,N_20776,N_20222);
or U23861 (N_23861,N_21785,N_21837);
or U23862 (N_23862,N_21747,N_20617);
and U23863 (N_23863,N_20591,N_21086);
or U23864 (N_23864,N_20369,N_20569);
nor U23865 (N_23865,N_20210,N_20488);
or U23866 (N_23866,N_21396,N_21036);
xnor U23867 (N_23867,N_20517,N_20163);
or U23868 (N_23868,N_20725,N_20206);
and U23869 (N_23869,N_20982,N_20547);
and U23870 (N_23870,N_20838,N_20839);
and U23871 (N_23871,N_21565,N_21127);
nand U23872 (N_23872,N_20735,N_21351);
nand U23873 (N_23873,N_20371,N_21209);
and U23874 (N_23874,N_20067,N_21615);
and U23875 (N_23875,N_21680,N_20748);
and U23876 (N_23876,N_20990,N_21789);
nor U23877 (N_23877,N_21979,N_21605);
xnor U23878 (N_23878,N_20288,N_21593);
xor U23879 (N_23879,N_21087,N_20064);
or U23880 (N_23880,N_21139,N_21414);
nand U23881 (N_23881,N_21648,N_21150);
and U23882 (N_23882,N_20849,N_20420);
nor U23883 (N_23883,N_21084,N_20813);
xnor U23884 (N_23884,N_21828,N_21886);
nor U23885 (N_23885,N_21235,N_20473);
and U23886 (N_23886,N_21010,N_20851);
nor U23887 (N_23887,N_20420,N_21245);
or U23888 (N_23888,N_20476,N_21123);
or U23889 (N_23889,N_21518,N_20717);
and U23890 (N_23890,N_21393,N_21564);
and U23891 (N_23891,N_21309,N_21077);
xnor U23892 (N_23892,N_20520,N_21764);
nand U23893 (N_23893,N_21967,N_20395);
xor U23894 (N_23894,N_21628,N_20916);
xor U23895 (N_23895,N_20766,N_21547);
nand U23896 (N_23896,N_21390,N_21687);
nor U23897 (N_23897,N_20756,N_20405);
and U23898 (N_23898,N_21231,N_21053);
or U23899 (N_23899,N_21739,N_21473);
nor U23900 (N_23900,N_21227,N_20915);
nor U23901 (N_23901,N_20120,N_20450);
or U23902 (N_23902,N_21671,N_20645);
nor U23903 (N_23903,N_20093,N_21555);
or U23904 (N_23904,N_21677,N_20319);
xor U23905 (N_23905,N_20061,N_21045);
nor U23906 (N_23906,N_21292,N_21704);
nand U23907 (N_23907,N_20225,N_21503);
nor U23908 (N_23908,N_21419,N_20576);
and U23909 (N_23909,N_21388,N_21707);
and U23910 (N_23910,N_21378,N_21401);
or U23911 (N_23911,N_20067,N_20246);
or U23912 (N_23912,N_20595,N_21210);
or U23913 (N_23913,N_20356,N_21073);
nand U23914 (N_23914,N_20562,N_21136);
xnor U23915 (N_23915,N_21503,N_20670);
or U23916 (N_23916,N_21087,N_20156);
nor U23917 (N_23917,N_20103,N_20362);
nand U23918 (N_23918,N_21740,N_21278);
and U23919 (N_23919,N_20453,N_21344);
nand U23920 (N_23920,N_20983,N_21069);
nand U23921 (N_23921,N_21947,N_21060);
nor U23922 (N_23922,N_20391,N_21138);
nor U23923 (N_23923,N_21609,N_21163);
nand U23924 (N_23924,N_21870,N_21027);
xor U23925 (N_23925,N_20960,N_21945);
xnor U23926 (N_23926,N_20395,N_20388);
nor U23927 (N_23927,N_21033,N_21898);
xnor U23928 (N_23928,N_20500,N_21686);
nor U23929 (N_23929,N_21461,N_21014);
nand U23930 (N_23930,N_21958,N_20761);
and U23931 (N_23931,N_21780,N_21688);
nand U23932 (N_23932,N_21123,N_21799);
nand U23933 (N_23933,N_20989,N_20614);
or U23934 (N_23934,N_20432,N_20268);
nor U23935 (N_23935,N_20707,N_21348);
xor U23936 (N_23936,N_20638,N_21330);
xnor U23937 (N_23937,N_21481,N_21970);
nor U23938 (N_23938,N_20113,N_21271);
nand U23939 (N_23939,N_21989,N_21351);
xor U23940 (N_23940,N_20593,N_20949);
or U23941 (N_23941,N_20512,N_21828);
xnor U23942 (N_23942,N_20023,N_21005);
nand U23943 (N_23943,N_20939,N_21036);
xor U23944 (N_23944,N_20089,N_20913);
or U23945 (N_23945,N_20178,N_21932);
and U23946 (N_23946,N_21807,N_21981);
or U23947 (N_23947,N_21073,N_21188);
or U23948 (N_23948,N_20453,N_20548);
nor U23949 (N_23949,N_20481,N_21389);
xor U23950 (N_23950,N_20547,N_20758);
nand U23951 (N_23951,N_21797,N_21827);
nor U23952 (N_23952,N_20545,N_21285);
xnor U23953 (N_23953,N_20038,N_21417);
nand U23954 (N_23954,N_21165,N_21206);
and U23955 (N_23955,N_20772,N_20759);
nor U23956 (N_23956,N_21778,N_21796);
nand U23957 (N_23957,N_20114,N_20321);
or U23958 (N_23958,N_21860,N_21493);
or U23959 (N_23959,N_20886,N_21711);
and U23960 (N_23960,N_20598,N_20150);
xnor U23961 (N_23961,N_20948,N_21361);
or U23962 (N_23962,N_21573,N_20904);
or U23963 (N_23963,N_20272,N_21026);
xor U23964 (N_23964,N_20698,N_21852);
or U23965 (N_23965,N_21389,N_21874);
xnor U23966 (N_23966,N_20479,N_20169);
nor U23967 (N_23967,N_21238,N_21614);
and U23968 (N_23968,N_20720,N_21175);
or U23969 (N_23969,N_20751,N_20031);
nor U23970 (N_23970,N_21367,N_21460);
nor U23971 (N_23971,N_21040,N_20320);
and U23972 (N_23972,N_21692,N_20298);
and U23973 (N_23973,N_21874,N_20936);
nor U23974 (N_23974,N_21838,N_21567);
and U23975 (N_23975,N_21801,N_21884);
nor U23976 (N_23976,N_20017,N_21977);
or U23977 (N_23977,N_21192,N_21330);
nand U23978 (N_23978,N_21380,N_20109);
and U23979 (N_23979,N_20004,N_20387);
nand U23980 (N_23980,N_20973,N_20521);
or U23981 (N_23981,N_20913,N_20600);
and U23982 (N_23982,N_20579,N_21071);
nand U23983 (N_23983,N_21983,N_20369);
and U23984 (N_23984,N_21501,N_20829);
xnor U23985 (N_23985,N_20137,N_20716);
or U23986 (N_23986,N_21751,N_20792);
and U23987 (N_23987,N_21226,N_21930);
or U23988 (N_23988,N_20296,N_20967);
xor U23989 (N_23989,N_20451,N_20889);
nor U23990 (N_23990,N_20710,N_21529);
nor U23991 (N_23991,N_20514,N_20590);
xnor U23992 (N_23992,N_21258,N_20394);
and U23993 (N_23993,N_21142,N_21081);
xor U23994 (N_23994,N_20037,N_21128);
nor U23995 (N_23995,N_20963,N_21786);
nor U23996 (N_23996,N_20092,N_21793);
nor U23997 (N_23997,N_21090,N_20666);
and U23998 (N_23998,N_21556,N_20332);
and U23999 (N_23999,N_20920,N_20681);
or U24000 (N_24000,N_23154,N_23980);
nand U24001 (N_24001,N_22251,N_23620);
xor U24002 (N_24002,N_23741,N_23318);
xnor U24003 (N_24003,N_22322,N_23405);
nand U24004 (N_24004,N_22441,N_22350);
xor U24005 (N_24005,N_22389,N_22652);
nand U24006 (N_24006,N_22950,N_22498);
or U24007 (N_24007,N_23041,N_23277);
or U24008 (N_24008,N_22957,N_23109);
nor U24009 (N_24009,N_22917,N_22418);
xnor U24010 (N_24010,N_22122,N_22561);
or U24011 (N_24011,N_23909,N_23144);
or U24012 (N_24012,N_22085,N_22696);
nor U24013 (N_24013,N_22523,N_22885);
nand U24014 (N_24014,N_22240,N_23801);
nand U24015 (N_24015,N_23990,N_22203);
xor U24016 (N_24016,N_22244,N_22765);
xor U24017 (N_24017,N_22267,N_23316);
and U24018 (N_24018,N_23789,N_22358);
xnor U24019 (N_24019,N_22433,N_23906);
nand U24020 (N_24020,N_23017,N_23013);
xnor U24021 (N_24021,N_23705,N_22737);
or U24022 (N_24022,N_23214,N_22010);
nor U24023 (N_24023,N_22020,N_23454);
or U24024 (N_24024,N_23252,N_22769);
and U24025 (N_24025,N_22780,N_23900);
nor U24026 (N_24026,N_23201,N_23241);
nand U24027 (N_24027,N_22697,N_22351);
nor U24028 (N_24028,N_23363,N_22406);
nand U24029 (N_24029,N_23351,N_23242);
and U24030 (N_24030,N_23938,N_23519);
xor U24031 (N_24031,N_22083,N_23075);
or U24032 (N_24032,N_22371,N_22397);
nand U24033 (N_24033,N_22205,N_23108);
nand U24034 (N_24034,N_23035,N_22384);
nand U24035 (N_24035,N_23934,N_23279);
or U24036 (N_24036,N_22145,N_22373);
and U24037 (N_24037,N_22223,N_22123);
and U24038 (N_24038,N_23096,N_22431);
nand U24039 (N_24039,N_22931,N_23633);
and U24040 (N_24040,N_23606,N_22781);
nand U24041 (N_24041,N_22288,N_23926);
nor U24042 (N_24042,N_23433,N_23976);
nand U24043 (N_24043,N_23100,N_22269);
nor U24044 (N_24044,N_22374,N_22098);
nand U24045 (N_24045,N_22930,N_22058);
nor U24046 (N_24046,N_22965,N_23314);
xnor U24047 (N_24047,N_23963,N_22045);
xnor U24048 (N_24048,N_23728,N_22790);
nand U24049 (N_24049,N_23731,N_23730);
and U24050 (N_24050,N_23130,N_22743);
xor U24051 (N_24051,N_22339,N_22392);
or U24052 (N_24052,N_22432,N_23739);
nor U24053 (N_24053,N_22257,N_23119);
nand U24054 (N_24054,N_22485,N_22290);
and U24055 (N_24055,N_23682,N_22225);
nor U24056 (N_24056,N_22210,N_23434);
and U24057 (N_24057,N_23590,N_23381);
nor U24058 (N_24058,N_23299,N_22978);
and U24059 (N_24059,N_22693,N_22239);
nor U24060 (N_24060,N_23063,N_22953);
nor U24061 (N_24061,N_23824,N_22943);
nor U24062 (N_24062,N_23210,N_23547);
nor U24063 (N_24063,N_22347,N_22448);
or U24064 (N_24064,N_23868,N_22197);
and U24065 (N_24065,N_23180,N_22548);
nand U24066 (N_24066,N_23892,N_22068);
nand U24067 (N_24067,N_23049,N_23298);
xor U24068 (N_24068,N_22655,N_22609);
or U24069 (N_24069,N_23920,N_23423);
and U24070 (N_24070,N_22755,N_22752);
and U24071 (N_24071,N_22886,N_22846);
nor U24072 (N_24072,N_22720,N_23006);
xor U24073 (N_24073,N_22914,N_23811);
and U24074 (N_24074,N_22165,N_23160);
nand U24075 (N_24075,N_23530,N_22894);
nand U24076 (N_24076,N_22393,N_23585);
and U24077 (N_24077,N_23465,N_23402);
or U24078 (N_24078,N_22834,N_22907);
or U24079 (N_24079,N_22346,N_23643);
xor U24080 (N_24080,N_23168,N_22802);
and U24081 (N_24081,N_23184,N_22836);
nor U24082 (N_24082,N_23131,N_22133);
xor U24083 (N_24083,N_23177,N_22593);
or U24084 (N_24084,N_23630,N_23354);
xor U24085 (N_24085,N_23641,N_23345);
or U24086 (N_24086,N_23735,N_22219);
or U24087 (N_24087,N_23880,N_22578);
nand U24088 (N_24088,N_23818,N_22153);
nor U24089 (N_24089,N_22273,N_23404);
or U24090 (N_24090,N_23974,N_23947);
and U24091 (N_24091,N_22382,N_22237);
nand U24092 (N_24092,N_22956,N_23967);
or U24093 (N_24093,N_23887,N_23674);
xor U24094 (N_24094,N_23376,N_23268);
or U24095 (N_24095,N_22070,N_22478);
nor U24096 (N_24096,N_22893,N_23128);
and U24097 (N_24097,N_22889,N_23280);
and U24098 (N_24098,N_23699,N_22614);
nor U24099 (N_24099,N_22610,N_23807);
xnor U24100 (N_24100,N_23879,N_23635);
xor U24101 (N_24101,N_22899,N_22403);
nand U24102 (N_24102,N_22360,N_23170);
and U24103 (N_24103,N_22856,N_23883);
nand U24104 (N_24104,N_22545,N_23720);
nor U24105 (N_24105,N_22276,N_23118);
or U24106 (N_24106,N_23307,N_22236);
xnor U24107 (N_24107,N_23955,N_22563);
nand U24108 (N_24108,N_22554,N_23271);
and U24109 (N_24109,N_22716,N_23386);
or U24110 (N_24110,N_23684,N_22048);
nand U24111 (N_24111,N_23761,N_23619);
nand U24112 (N_24112,N_23207,N_22014);
nor U24113 (N_24113,N_22046,N_22466);
nand U24114 (N_24114,N_23228,N_23132);
xor U24115 (N_24115,N_22798,N_23962);
xnor U24116 (N_24116,N_22446,N_23841);
nand U24117 (N_24117,N_22952,N_22558);
nand U24118 (N_24118,N_22300,N_23979);
and U24119 (N_24119,N_23670,N_22552);
nand U24120 (N_24120,N_22616,N_22234);
xnor U24121 (N_24121,N_23029,N_22738);
nor U24122 (N_24122,N_22060,N_22143);
or U24123 (N_24123,N_22302,N_23793);
nor U24124 (N_24124,N_22665,N_23021);
xnor U24125 (N_24125,N_23200,N_23320);
or U24126 (N_24126,N_23098,N_23509);
nor U24127 (N_24127,N_22991,N_22401);
and U24128 (N_24128,N_22007,N_22277);
xor U24129 (N_24129,N_22296,N_22844);
or U24130 (N_24130,N_23421,N_22670);
or U24131 (N_24131,N_23165,N_23217);
xor U24132 (N_24132,N_23999,N_23065);
nor U24133 (N_24133,N_23432,N_22641);
nand U24134 (N_24134,N_22581,N_22238);
nand U24135 (N_24135,N_23448,N_22447);
and U24136 (N_24136,N_23708,N_23663);
nor U24137 (N_24137,N_22196,N_22570);
and U24138 (N_24138,N_23992,N_22378);
nor U24139 (N_24139,N_22793,N_23368);
nor U24140 (N_24140,N_22774,N_22119);
and U24141 (N_24141,N_22125,N_22771);
xor U24142 (N_24142,N_23628,N_23863);
xnor U24143 (N_24143,N_23366,N_22586);
xor U24144 (N_24144,N_22486,N_23026);
nand U24145 (N_24145,N_22206,N_22905);
xnor U24146 (N_24146,N_22514,N_23501);
xor U24147 (N_24147,N_23971,N_23870);
nand U24148 (N_24148,N_23559,N_23987);
nand U24149 (N_24149,N_23477,N_23493);
nor U24150 (N_24150,N_23548,N_23072);
nand U24151 (N_24151,N_23073,N_22129);
and U24152 (N_24152,N_22567,N_22672);
or U24153 (N_24153,N_22702,N_22032);
and U24154 (N_24154,N_22161,N_22541);
nand U24155 (N_24155,N_23722,N_23607);
nand U24156 (N_24156,N_22089,N_22929);
nor U24157 (N_24157,N_23498,N_23040);
xor U24158 (N_24158,N_22015,N_22078);
and U24159 (N_24159,N_23986,N_23134);
nor U24160 (N_24160,N_23608,N_23101);
xnor U24161 (N_24161,N_23192,N_23341);
xor U24162 (N_24162,N_22249,N_22369);
nor U24163 (N_24163,N_23324,N_23918);
or U24164 (N_24164,N_22577,N_22660);
xnor U24165 (N_24165,N_23998,N_22380);
nor U24166 (N_24166,N_22892,N_23199);
or U24167 (N_24167,N_23899,N_23092);
or U24168 (N_24168,N_23253,N_23601);
xnor U24169 (N_24169,N_23171,N_23895);
nor U24170 (N_24170,N_23556,N_22183);
nand U24171 (N_24171,N_22517,N_23382);
or U24172 (N_24172,N_23611,N_23779);
and U24173 (N_24173,N_23055,N_22438);
or U24174 (N_24174,N_22345,N_23403);
and U24175 (N_24175,N_22465,N_23531);
or U24176 (N_24176,N_23666,N_23564);
xor U24177 (N_24177,N_22063,N_23413);
nand U24178 (N_24178,N_22867,N_23475);
xnor U24179 (N_24179,N_22612,N_23491);
or U24180 (N_24180,N_22625,N_22149);
or U24181 (N_24181,N_23825,N_23575);
and U24182 (N_24182,N_22022,N_22185);
nor U24183 (N_24183,N_23579,N_22128);
xor U24184 (N_24184,N_23757,N_22118);
xnor U24185 (N_24185,N_23037,N_23336);
nor U24186 (N_24186,N_23284,N_23993);
or U24187 (N_24187,N_22751,N_22450);
xnor U24188 (N_24188,N_23520,N_22766);
xor U24189 (N_24189,N_23169,N_23246);
and U24190 (N_24190,N_23497,N_23675);
and U24191 (N_24191,N_22319,N_22722);
nor U24192 (N_24192,N_23446,N_23983);
xnor U24193 (N_24193,N_23923,N_23410);
and U24194 (N_24194,N_23009,N_23285);
nor U24195 (N_24195,N_22396,N_22939);
xor U24196 (N_24196,N_23309,N_23959);
and U24197 (N_24197,N_22835,N_23780);
nor U24198 (N_24198,N_23267,N_23102);
nand U24199 (N_24199,N_23227,N_22211);
and U24200 (N_24200,N_23347,N_23356);
nand U24201 (N_24201,N_22800,N_22940);
nor U24202 (N_24202,N_22535,N_23353);
xor U24203 (N_24203,N_23183,N_22160);
nor U24204 (N_24204,N_23950,N_23143);
xor U24205 (N_24205,N_23809,N_22687);
xnor U24206 (N_24206,N_22031,N_23945);
and U24207 (N_24207,N_22003,N_22233);
xnor U24208 (N_24208,N_23204,N_23566);
nand U24209 (N_24209,N_23237,N_22194);
or U24210 (N_24210,N_23397,N_23790);
nand U24211 (N_24211,N_23921,N_23594);
xnor U24212 (N_24212,N_22248,N_22445);
or U24213 (N_24213,N_22162,N_23563);
xnor U24214 (N_24214,N_22811,N_22169);
and U24215 (N_24215,N_22908,N_23012);
xnor U24216 (N_24216,N_23944,N_22657);
nand U24217 (N_24217,N_23272,N_23617);
xnor U24218 (N_24218,N_23558,N_23953);
nand U24219 (N_24219,N_22390,N_22011);
and U24220 (N_24220,N_23625,N_22782);
and U24221 (N_24221,N_23034,N_22134);
or U24222 (N_24222,N_23539,N_22414);
nor U24223 (N_24223,N_22324,N_22884);
nand U24224 (N_24224,N_23588,N_23414);
nand U24225 (N_24225,N_22583,N_22503);
xnor U24226 (N_24226,N_23317,N_23360);
nand U24227 (N_24227,N_23703,N_22521);
xnor U24228 (N_24228,N_23834,N_23823);
xor U24229 (N_24229,N_23771,N_23802);
nor U24230 (N_24230,N_23885,N_22824);
or U24231 (N_24231,N_23660,N_22344);
nand U24232 (N_24232,N_22757,N_23435);
nor U24233 (N_24233,N_22792,N_23212);
or U24234 (N_24234,N_22648,N_23653);
xnor U24235 (N_24235,N_22611,N_22964);
xor U24236 (N_24236,N_22840,N_23349);
or U24237 (N_24237,N_23221,N_23615);
nand U24238 (N_24238,N_22180,N_23278);
nor U24239 (N_24239,N_22749,N_23464);
or U24240 (N_24240,N_23849,N_22500);
nand U24241 (N_24241,N_22540,N_23139);
or U24242 (N_24242,N_22565,N_23047);
nand U24243 (N_24243,N_22767,N_23521);
nand U24244 (N_24244,N_22857,N_22411);
or U24245 (N_24245,N_23273,N_22218);
and U24246 (N_24246,N_22712,N_23492);
and U24247 (N_24247,N_22265,N_23600);
xnor U24248 (N_24248,N_22922,N_23513);
xor U24249 (N_24249,N_23562,N_22315);
and U24250 (N_24250,N_23969,N_22264);
or U24251 (N_24251,N_22076,N_23915);
nor U24252 (N_24252,N_22379,N_22684);
nand U24253 (N_24253,N_23460,N_22082);
or U24254 (N_24254,N_22870,N_23455);
nor U24255 (N_24255,N_23773,N_23912);
nand U24256 (N_24256,N_23791,N_22317);
xnor U24257 (N_24257,N_23829,N_23127);
nand U24258 (N_24258,N_23275,N_23541);
nor U24259 (N_24259,N_22963,N_22739);
nand U24260 (N_24260,N_23984,N_23991);
or U24261 (N_24261,N_23438,N_22470);
and U24262 (N_24262,N_22971,N_22801);
or U24263 (N_24263,N_23724,N_22404);
nor U24264 (N_24264,N_23325,N_23815);
or U24265 (N_24265,N_22289,N_22969);
and U24266 (N_24266,N_22226,N_23977);
nand U24267 (N_24267,N_23924,N_22255);
or U24268 (N_24268,N_23255,N_22148);
xnor U24269 (N_24269,N_22510,N_23916);
nor U24270 (N_24270,N_22222,N_22997);
nor U24271 (N_24271,N_23452,N_22762);
nand U24272 (N_24272,N_23147,N_23702);
and U24273 (N_24273,N_23604,N_23262);
xor U24274 (N_24274,N_23798,N_23685);
xor U24275 (N_24275,N_23804,N_22182);
nor U24276 (N_24276,N_23764,N_22826);
xor U24277 (N_24277,N_22776,N_23269);
or U24278 (N_24278,N_23538,N_22910);
and U24279 (N_24279,N_22603,N_22778);
xnor U24280 (N_24280,N_23954,N_22830);
or U24281 (N_24281,N_23932,N_22368);
xor U24282 (N_24282,N_23456,N_23860);
xnor U24283 (N_24283,N_22674,N_23678);
nor U24284 (N_24284,N_23522,N_22278);
and U24285 (N_24285,N_23093,N_22336);
nand U24286 (N_24286,N_22761,N_23067);
nor U24287 (N_24287,N_23332,N_22029);
nor U24288 (N_24288,N_23828,N_22139);
xor U24289 (N_24289,N_22658,N_23573);
nand U24290 (N_24290,N_23297,N_22543);
nand U24291 (N_24291,N_23867,N_23443);
xor U24292 (N_24292,N_23261,N_23442);
and U24293 (N_24293,N_23126,N_23612);
nor U24294 (N_24294,N_23514,N_22443);
xor U24295 (N_24295,N_23239,N_23551);
nand U24296 (N_24296,N_22496,N_22320);
xnor U24297 (N_24297,N_23645,N_22097);
nor U24298 (N_24298,N_23507,N_22945);
nand U24299 (N_24299,N_23406,N_23107);
or U24300 (N_24300,N_23213,N_22906);
and U24301 (N_24301,N_22873,N_23706);
nor U24302 (N_24302,N_23225,N_23140);
nand U24303 (N_24303,N_23133,N_23206);
xor U24304 (N_24304,N_22602,N_22947);
nor U24305 (N_24305,N_23468,N_22629);
nand U24306 (N_24306,N_22462,N_23300);
and U24307 (N_24307,N_22297,N_23240);
and U24308 (N_24308,N_23750,N_23570);
or U24309 (N_24309,N_22456,N_22067);
nor U24310 (N_24310,N_22187,N_23994);
or U24311 (N_24311,N_23597,N_23027);
or U24312 (N_24312,N_23981,N_22310);
and U24313 (N_24313,N_23142,N_23523);
nor U24314 (N_24314,N_22457,N_22656);
and U24315 (N_24315,N_23458,N_23698);
and U24316 (N_24316,N_22301,N_22564);
xnor U24317 (N_24317,N_22831,N_22399);
and U24318 (N_24318,N_22016,N_22281);
nand U24319 (N_24319,N_22174,N_23679);
or U24320 (N_24320,N_23305,N_23677);
xnor U24321 (N_24321,N_22027,N_23748);
nand U24322 (N_24322,N_23024,N_23803);
and U24323 (N_24323,N_22419,N_23765);
nand U24324 (N_24324,N_23135,N_23424);
and U24325 (N_24325,N_22140,N_23669);
nand U24326 (N_24326,N_23744,N_22512);
nor U24327 (N_24327,N_23762,N_22794);
or U24328 (N_24328,N_23484,N_22505);
nor U24329 (N_24329,N_23056,N_23265);
or U24330 (N_24330,N_23772,N_22137);
nand U24331 (N_24331,N_23937,N_23529);
or U24332 (N_24332,N_23589,N_22608);
nand U24333 (N_24333,N_23420,N_22595);
or U24334 (N_24334,N_22176,N_22537);
or U24335 (N_24335,N_22136,N_22591);
xor U24336 (N_24336,N_22633,N_22250);
xnor U24337 (N_24337,N_23767,N_22370);
xnor U24338 (N_24338,N_22103,N_22557);
xnor U24339 (N_24339,N_23110,N_23089);
or U24340 (N_24340,N_23036,N_22460);
xnor U24341 (N_24341,N_23166,N_23871);
or U24342 (N_24342,N_23939,N_22551);
xor U24343 (N_24343,N_22622,N_22903);
or U24344 (N_24344,N_22348,N_23822);
or U24345 (N_24345,N_23572,N_22542);
or U24346 (N_24346,N_23489,N_22051);
nor U24347 (N_24347,N_22335,N_22803);
nand U24348 (N_24348,N_22480,N_23008);
xor U24349 (N_24349,N_22667,N_23494);
nand U24350 (N_24350,N_23161,N_23205);
xnor U24351 (N_24351,N_22705,N_23683);
nand U24352 (N_24352,N_23629,N_22038);
and U24353 (N_24353,N_23931,N_22700);
xor U24354 (N_24354,N_23553,N_22057);
and U24355 (N_24355,N_22475,N_23904);
nor U24356 (N_24356,N_23820,N_23304);
xor U24357 (N_24357,N_22502,N_22261);
and U24358 (N_24358,N_22709,N_22146);
nand U24359 (N_24359,N_23812,N_23658);
and U24360 (N_24360,N_23693,N_22481);
xnor U24361 (N_24361,N_22808,N_22030);
and U24362 (N_24362,N_22483,N_23203);
and U24363 (N_24363,N_22984,N_23232);
nor U24364 (N_24364,N_23786,N_23393);
nor U24365 (N_24365,N_23334,N_22632);
nand U24366 (N_24366,N_23343,N_23624);
xnor U24367 (N_24367,N_23592,N_22094);
nor U24368 (N_24368,N_23408,N_22275);
nand U24369 (N_24369,N_22054,N_22155);
and U24370 (N_24370,N_23196,N_23587);
xor U24371 (N_24371,N_22050,N_22822);
nand U24372 (N_24372,N_22469,N_22796);
and U24373 (N_24373,N_22410,N_23444);
xor U24374 (N_24374,N_22408,N_22472);
xnor U24375 (N_24375,N_22976,N_22574);
nand U24376 (N_24376,N_22627,N_23881);
nand U24377 (N_24377,N_22109,N_22065);
nand U24378 (N_24378,N_23321,N_23734);
or U24379 (N_24379,N_22449,N_22299);
nor U24380 (N_24380,N_23743,N_22074);
nor U24381 (N_24381,N_22178,N_22746);
or U24382 (N_24382,N_23282,N_23542);
or U24383 (N_24383,N_23972,N_23441);
and U24384 (N_24384,N_22960,N_23023);
or U24385 (N_24385,N_22748,N_23537);
nand U24386 (N_24386,N_23188,N_23015);
and U24387 (N_24387,N_22513,N_22004);
and U24388 (N_24388,N_23864,N_23634);
and U24389 (N_24389,N_22691,N_22938);
nor U24390 (N_24390,N_22915,N_23209);
nand U24391 (N_24391,N_22506,N_22066);
nor U24392 (N_24392,N_23701,N_22309);
nand U24393 (N_24393,N_23346,N_22387);
nor U24394 (N_24394,N_23869,N_22572);
and U24395 (N_24395,N_22529,N_23797);
and U24396 (N_24396,N_23535,N_22477);
or U24397 (N_24397,N_22896,N_23051);
nand U24398 (N_24398,N_23568,N_23806);
nor U24399 (N_24399,N_22579,N_22987);
nor U24400 (N_24400,N_22852,N_22839);
nand U24401 (N_24401,N_23555,N_22208);
or U24402 (N_24402,N_22402,N_23311);
xnor U24403 (N_24403,N_23636,N_22644);
nand U24404 (N_24404,N_23123,N_22550);
or U24405 (N_24405,N_23940,N_22817);
nor U24406 (N_24406,N_23358,N_23627);
and U24407 (N_24407,N_23099,N_22809);
nor U24408 (N_24408,N_22902,N_23533);
and U24409 (N_24409,N_22042,N_22772);
or U24410 (N_24410,N_22921,N_22895);
xor U24411 (N_24411,N_22788,N_23893);
nor U24412 (N_24412,N_22400,N_22422);
or U24413 (N_24413,N_23340,N_23988);
nand U24414 (N_24414,N_22292,N_23038);
xnor U24415 (N_24415,N_23374,N_23303);
xnor U24416 (N_24416,N_22663,N_22785);
xor U24417 (N_24417,N_23220,N_22759);
or U24418 (N_24418,N_22192,N_23518);
and U24419 (N_24419,N_22993,N_23956);
nor U24420 (N_24420,N_23230,N_23081);
nor U24421 (N_24421,N_23264,N_22973);
nor U24422 (N_24422,N_22434,N_22594);
xnor U24423 (N_24423,N_22912,N_23391);
or U24424 (N_24424,N_23090,N_22628);
or U24425 (N_24425,N_23859,N_22723);
nand U24426 (N_24426,N_22252,N_23796);
nand U24427 (N_24427,N_22784,N_22685);
and U24428 (N_24428,N_23831,N_23190);
and U24429 (N_24429,N_23447,N_22495);
or U24430 (N_24430,N_22459,N_22688);
and U24431 (N_24431,N_23782,N_22084);
xor U24432 (N_24432,N_23626,N_22911);
nand U24433 (N_24433,N_23163,N_22850);
xor U24434 (N_24434,N_22686,N_22127);
or U24435 (N_24435,N_23256,N_22768);
and U24436 (N_24436,N_22312,N_22209);
or U24437 (N_24437,N_22639,N_23218);
or U24438 (N_24438,N_22282,N_23652);
nor U24439 (N_24439,N_22636,N_22484);
xnor U24440 (N_24440,N_22928,N_23052);
xnor U24441 (N_24441,N_22055,N_22440);
or U24442 (N_24442,N_23364,N_22756);
xor U24443 (N_24443,N_22059,N_23651);
and U24444 (N_24444,N_23655,N_23578);
nand U24445 (N_24445,N_23377,N_22659);
or U24446 (N_24446,N_22843,N_22592);
xnor U24447 (N_24447,N_23357,N_22823);
and U24448 (N_24448,N_23266,N_22235);
nor U24449 (N_24449,N_23445,N_22977);
xnor U24450 (N_24450,N_23153,N_23044);
or U24451 (N_24451,N_23472,N_22888);
and U24452 (N_24452,N_23361,N_23799);
or U24453 (N_24453,N_23754,N_22544);
nor U24454 (N_24454,N_22872,N_23150);
or U24455 (N_24455,N_23544,N_23759);
nor U24456 (N_24456,N_22201,N_23580);
or U24457 (N_24457,N_23479,N_23059);
nor U24458 (N_24458,N_22386,N_22284);
and U24459 (N_24459,N_23223,N_22253);
and U24460 (N_24460,N_23198,N_22955);
nor U24461 (N_24461,N_22718,N_23014);
xor U24462 (N_24462,N_23949,N_22881);
or U24463 (N_24463,N_23736,N_22919);
nor U24464 (N_24464,N_23111,N_22081);
or U24465 (N_24465,N_23574,N_23076);
or U24466 (N_24466,N_23466,N_23640);
xnor U24467 (N_24467,N_23287,N_22428);
or U24468 (N_24468,N_23245,N_23086);
nor U24469 (N_24469,N_22242,N_22154);
xnor U24470 (N_24470,N_22323,N_23890);
and U24471 (N_24471,N_23018,N_22532);
nand U24472 (N_24472,N_23581,N_22337);
or U24473 (N_24473,N_22706,N_23858);
nand U24474 (N_24474,N_23853,N_22962);
and U24475 (N_24475,N_23785,N_22556);
or U24476 (N_24476,N_22651,N_23647);
or U24477 (N_24477,N_23727,N_23610);
nor U24478 (N_24478,N_22522,N_22287);
xnor U24479 (N_24479,N_23191,N_23552);
nand U24480 (N_24480,N_23503,N_23031);
xnor U24481 (N_24481,N_22879,N_22075);
nand U24482 (N_24482,N_22096,N_23756);
xor U24483 (N_24483,N_23776,N_22515);
and U24484 (N_24484,N_23697,N_22062);
nor U24485 (N_24485,N_22329,N_23751);
xnor U24486 (N_24486,N_22647,N_23066);
xnor U24487 (N_24487,N_22304,N_23726);
xnor U24488 (N_24488,N_23914,N_23861);
nor U24489 (N_24489,N_22326,N_22394);
and U24490 (N_24490,N_22135,N_22607);
xor U24491 (N_24491,N_23692,N_23263);
nor U24492 (N_24492,N_22653,N_23339);
nor U24493 (N_24493,N_23409,N_22274);
or U24494 (N_24494,N_23257,N_22927);
nand U24495 (N_24495,N_22724,N_22314);
nand U24496 (N_24496,N_22575,N_23331);
xnor U24497 (N_24497,N_23387,N_22043);
or U24498 (N_24498,N_23810,N_22841);
and U24499 (N_24499,N_23175,N_22388);
and U24500 (N_24500,N_23412,N_23373);
xnor U24501 (N_24501,N_23083,N_23022);
or U24502 (N_24502,N_23695,N_22429);
nor U24503 (N_24503,N_23676,N_22730);
and U24504 (N_24504,N_23483,N_23482);
or U24505 (N_24505,N_22463,N_22241);
nand U24506 (N_24506,N_22626,N_22509);
or U24507 (N_24507,N_22590,N_23827);
nor U24508 (N_24508,N_22604,N_23352);
nand U24509 (N_24509,N_23337,N_22416);
or U24510 (N_24510,N_22559,N_22818);
and U24511 (N_24511,N_23898,N_22151);
xnor U24512 (N_24512,N_22280,N_23054);
and U24513 (N_24513,N_22033,N_22254);
and U24514 (N_24514,N_22362,N_23593);
nand U24515 (N_24515,N_22980,N_23687);
nor U24516 (N_24516,N_22618,N_23462);
nand U24517 (N_24517,N_23486,N_23045);
nor U24518 (N_24518,N_23187,N_22476);
nand U24519 (N_24519,N_23930,N_22126);
or U24520 (N_24520,N_23646,N_23439);
nand U24521 (N_24521,N_22828,N_22854);
nand U24522 (N_24522,N_23019,N_23826);
nor U24523 (N_24523,N_23621,N_22701);
and U24524 (N_24524,N_22167,N_22471);
or U24525 (N_24525,N_23136,N_23896);
nor U24526 (N_24526,N_23536,N_23978);
xor U24527 (N_24527,N_23717,N_23157);
nor U24528 (N_24528,N_23814,N_22147);
and U24529 (N_24529,N_23840,N_22637);
or U24530 (N_24530,N_22833,N_22357);
and U24531 (N_24531,N_23057,N_23661);
nor U24532 (N_24532,N_22023,N_22853);
and U24533 (N_24533,N_23659,N_22571);
nor U24534 (N_24534,N_23689,N_22131);
nand U24535 (N_24535,N_22138,N_23046);
or U24536 (N_24536,N_23813,N_23231);
or U24537 (N_24537,N_22661,N_22061);
nand U24538 (N_24538,N_22729,N_22009);
or U24539 (N_24539,N_23436,N_22095);
and U24540 (N_24540,N_22937,N_23208);
nand U24541 (N_24541,N_23302,N_23768);
and U24542 (N_24542,N_23821,N_23292);
and U24543 (N_24543,N_23583,N_22019);
nand U24544 (N_24544,N_23838,N_22887);
xnor U24545 (N_24545,N_22941,N_22584);
and U24546 (N_24546,N_23080,N_22650);
xnor U24547 (N_24547,N_22420,N_23943);
nand U24548 (N_24548,N_23557,N_22582);
xnor U24549 (N_24549,N_22479,N_23910);
nor U24550 (N_24550,N_22711,N_23700);
or U24551 (N_24551,N_23688,N_22491);
xnor U24552 (N_24552,N_23369,N_22159);
nand U24553 (N_24553,N_22646,N_22717);
and U24554 (N_24554,N_23618,N_22926);
nand U24555 (N_24555,N_23129,N_23159);
and U24556 (N_24556,N_23654,N_22436);
nand U24557 (N_24557,N_23470,N_22795);
and U24558 (N_24558,N_22677,N_22385);
and U24559 (N_24559,N_23857,N_23020);
nor U24560 (N_24560,N_22526,N_23560);
nand U24561 (N_24561,N_23313,N_22130);
and U24562 (N_24562,N_23295,N_23362);
xor U24563 (N_24563,N_22961,N_23389);
and U24564 (N_24564,N_23028,N_23884);
or U24565 (N_24565,N_23179,N_22455);
nor U24566 (N_24566,N_22286,N_23516);
or U24567 (N_24567,N_23459,N_22942);
nor U24568 (N_24568,N_22259,N_22156);
or U24569 (N_24569,N_22698,N_23306);
xnor U24570 (N_24570,N_22263,N_23480);
xor U24571 (N_24571,N_22461,N_23338);
nor U24572 (N_24572,N_22181,N_23524);
nand U24573 (N_24573,N_23960,N_22566);
nand U24574 (N_24574,N_23997,N_23367);
nand U24575 (N_24575,N_23189,N_23105);
or U24576 (N_24576,N_23506,N_22334);
and U24577 (N_24577,N_22707,N_23030);
nor U24578 (N_24578,N_22170,N_22990);
nor U24579 (N_24579,N_22124,N_22008);
nor U24580 (N_24580,N_23379,N_22900);
and U24581 (N_24581,N_22115,N_23996);
or U24582 (N_24582,N_23631,N_22069);
xor U24583 (N_24583,N_23270,N_22342);
or U24584 (N_24584,N_22549,N_23819);
and U24585 (N_24585,N_22635,N_22925);
and U24586 (N_24586,N_23048,N_22682);
and U24587 (N_24587,N_22807,N_23286);
xnor U24588 (N_24588,N_23862,N_23856);
xnor U24589 (N_24589,N_22328,N_22959);
nor U24590 (N_24590,N_22508,N_23005);
nor U24591 (N_24591,N_22972,N_23836);
and U24592 (N_24592,N_22295,N_23847);
or U24593 (N_24593,N_22860,N_22053);
nand U24594 (N_24594,N_23586,N_23673);
xor U24595 (N_24595,N_22601,N_23872);
nor U24596 (N_24596,N_22989,N_23490);
xor U24597 (N_24597,N_22882,N_22524);
nand U24598 (N_24598,N_22375,N_23233);
nor U24599 (N_24599,N_23342,N_23848);
and U24600 (N_24600,N_23243,N_22327);
or U24601 (N_24601,N_22664,N_22909);
nor U24602 (N_24602,N_23752,N_22710);
xor U24603 (N_24603,N_23725,N_23238);
nand U24604 (N_24604,N_22333,N_23886);
or U24605 (N_24605,N_23390,N_23903);
xnor U24606 (N_24606,N_23467,N_23182);
nor U24607 (N_24607,N_23079,N_23158);
nand U24608 (N_24608,N_23528,N_23719);
and U24609 (N_24609,N_22100,N_22804);
xor U24610 (N_24610,N_23417,N_23650);
or U24611 (N_24611,N_23301,N_23584);
nor U24612 (N_24612,N_22731,N_23504);
or U24613 (N_24613,N_23348,N_23576);
xor U24614 (N_24614,N_23396,N_22298);
xor U24615 (N_24615,N_22423,N_23733);
nor U24616 (N_24616,N_22725,N_23155);
nand U24617 (N_24617,N_22190,N_23602);
and U24618 (N_24618,N_22613,N_23260);
or U24619 (N_24619,N_23696,N_22132);
xor U24620 (N_24620,N_22285,N_22488);
xnor U24621 (N_24621,N_23164,N_22858);
nand U24622 (N_24622,N_22740,N_22935);
nor U24623 (N_24623,N_22770,N_23970);
xnor U24624 (N_24624,N_22024,N_22227);
nand U24625 (N_24625,N_22736,N_22837);
nor U24626 (N_24626,N_22934,N_23681);
or U24627 (N_24627,N_22983,N_22158);
nor U24628 (N_24628,N_23973,N_22041);
xor U24629 (N_24629,N_23565,N_23478);
and U24630 (N_24630,N_22539,N_22871);
or U24631 (N_24631,N_22246,N_23355);
nand U24632 (N_24632,N_22534,N_22489);
nor U24633 (N_24633,N_22340,N_23319);
nand U24634 (N_24634,N_22519,N_22415);
and U24635 (N_24635,N_22754,N_22228);
nand U24636 (N_24636,N_22426,N_23487);
nor U24637 (N_24637,N_23437,N_22113);
or U24638 (N_24638,N_22245,N_23113);
and U24639 (N_24639,N_22028,N_23668);
xor U24640 (N_24640,N_22721,N_23917);
and U24641 (N_24641,N_23808,N_22247);
nor U24642 (N_24642,N_23975,N_22681);
nor U24643 (N_24643,N_23738,N_23958);
nor U24644 (N_24644,N_22842,N_22680);
nand U24645 (N_24645,N_23071,N_23665);
xor U24646 (N_24646,N_22487,N_23569);
nand U24647 (N_24647,N_22838,N_23671);
or U24648 (N_24648,N_22948,N_22520);
xor U24649 (N_24649,N_22052,N_22855);
xor U24650 (N_24650,N_22819,N_23137);
nand U24651 (N_24651,N_22553,N_22880);
xnor U24652 (N_24652,N_23656,N_23440);
nor U24653 (N_24653,N_22079,N_22692);
xor U24654 (N_24654,N_22341,N_22606);
xor U24655 (N_24655,N_23913,N_22676);
xor U24656 (N_24656,N_22035,N_22102);
xnor U24657 (N_24657,N_23219,N_22995);
and U24658 (N_24658,N_22600,N_22376);
nand U24659 (N_24659,N_22525,N_22630);
nand U24660 (N_24660,N_22704,N_22427);
and U24661 (N_24661,N_23876,N_22435);
and U24662 (N_24662,N_23657,N_22874);
xor U24663 (N_24663,N_22719,N_23236);
and U24664 (N_24664,N_23429,N_23680);
nand U24665 (N_24665,N_23082,N_23289);
nor U24666 (N_24666,N_23419,N_23901);
or U24667 (N_24667,N_22453,N_22560);
nand U24668 (N_24668,N_22821,N_22256);
nor U24669 (N_24669,N_22979,N_22308);
xor U24670 (N_24670,N_23399,N_22417);
xor U24671 (N_24671,N_22111,N_22642);
or U24672 (N_24672,N_22649,N_23598);
xnor U24673 (N_24673,N_23561,N_23854);
and U24674 (N_24674,N_22332,N_23042);
or U24675 (N_24675,N_22482,N_23525);
nand U24676 (N_24676,N_22865,N_23614);
xor U24677 (N_24677,N_23016,N_23936);
and U24678 (N_24678,N_22034,N_23835);
xnor U24679 (N_24679,N_23070,N_23816);
nand U24680 (N_24680,N_23922,N_23721);
or U24681 (N_24681,N_23222,N_23194);
and U24682 (N_24682,N_22958,N_22527);
or U24683 (N_24683,N_22474,N_22207);
xnor U24684 (N_24684,N_23450,N_23845);
or U24685 (N_24685,N_23897,N_23690);
and U24686 (N_24686,N_22851,N_22012);
nor U24687 (N_24687,N_22923,N_23495);
xnor U24688 (N_24688,N_23426,N_23145);
nand U24689 (N_24689,N_22039,N_22585);
xnor U24690 (N_24690,N_23120,N_23929);
and U24691 (N_24691,N_22671,N_22064);
xor U24692 (N_24692,N_22077,N_23167);
nor U24693 (N_24693,N_23952,N_22377);
nand U24694 (N_24694,N_22813,N_23211);
nor U24695 (N_24695,N_23258,N_23637);
nor U24696 (N_24696,N_22002,N_22981);
nand U24697 (N_24697,N_23254,N_23534);
nor U24698 (N_24698,N_23648,N_23370);
nor U24699 (N_24699,N_22175,N_23686);
and U24700 (N_24700,N_22913,N_23644);
or U24701 (N_24701,N_22425,N_22229);
or U24702 (N_24702,N_23453,N_22631);
nand U24703 (N_24703,N_23502,N_23077);
nand U24704 (N_24704,N_23550,N_23948);
xor U24705 (N_24705,N_22949,N_22005);
nand U24706 (N_24706,N_23982,N_23329);
nand U24707 (N_24707,N_22538,N_22464);
nand U24708 (N_24708,N_23616,N_23599);
nor U24709 (N_24709,N_22862,N_22714);
or U24710 (N_24710,N_22092,N_22338);
nor U24711 (N_24711,N_22025,N_22086);
xor U24712 (N_24712,N_22982,N_23554);
or U24713 (N_24713,N_22679,N_23770);
and U24714 (N_24714,N_23985,N_23380);
and U24715 (N_24715,N_22662,N_23115);
nor U24716 (N_24716,N_23084,N_23778);
nor U24717 (N_24717,N_22198,N_22473);
xnor U24718 (N_24718,N_22305,N_22619);
nand U24719 (N_24719,N_22918,N_23907);
xnor U24720 (N_24720,N_23852,N_22307);
nor U24721 (N_24721,N_23244,N_22444);
xnor U24722 (N_24722,N_22791,N_22499);
and U24723 (N_24723,N_22430,N_23425);
nor U24724 (N_24724,N_22954,N_23638);
and U24725 (N_24725,N_22383,N_22114);
and U24726 (N_24726,N_22279,N_23753);
nand U24727 (N_24727,N_22268,N_22797);
nand U24728 (N_24728,N_23649,N_23463);
nor U24729 (N_24729,N_22547,N_22293);
nor U24730 (N_24730,N_22763,N_22080);
or U24731 (N_24731,N_23335,N_23251);
nand U24732 (N_24732,N_23844,N_23087);
nor U24733 (N_24733,N_23050,N_23125);
or U24734 (N_24734,N_23186,N_23007);
xor U24735 (N_24735,N_22331,N_22088);
and U24736 (N_24736,N_23526,N_23310);
xor U24737 (N_24737,N_23817,N_22573);
or U24738 (N_24738,N_22202,N_22643);
nand U24739 (N_24739,N_22742,N_23508);
nand U24740 (N_24740,N_22232,N_22988);
or U24741 (N_24741,N_23116,N_22398);
xor U24742 (N_24742,N_22589,N_23747);
nor U24743 (N_24743,N_22107,N_22968);
and U24744 (N_24744,N_22177,N_22220);
or U24745 (N_24745,N_22645,N_23176);
xor U24746 (N_24746,N_23234,N_23274);
or U24747 (N_24747,N_22294,N_22087);
nor U24748 (N_24748,N_23141,N_23546);
and U24749 (N_24749,N_23062,N_22090);
nand U24750 (N_24750,N_23935,N_22845);
or U24751 (N_24751,N_22270,N_22617);
nand U24752 (N_24752,N_23249,N_22221);
and U24753 (N_24753,N_22193,N_23742);
xor U24754 (N_24754,N_22204,N_22179);
xor U24755 (N_24755,N_22999,N_22897);
or U24756 (N_24756,N_23001,N_22861);
or U24757 (N_24757,N_23758,N_22623);
or U24758 (N_24758,N_23795,N_22946);
nand U24759 (N_24759,N_23595,N_23333);
nand U24760 (N_24760,N_22878,N_23322);
and U24761 (N_24761,N_23053,N_23609);
nor U24762 (N_24762,N_22599,N_23315);
and U24763 (N_24763,N_22216,N_22173);
nand U24764 (N_24764,N_22355,N_23877);
or U24765 (N_24765,N_23596,N_22006);
and U24766 (N_24766,N_22624,N_22303);
nand U24767 (N_24767,N_22951,N_23216);
xor U24768 (N_24768,N_23185,N_22775);
nor U24769 (N_24769,N_22395,N_22587);
and U24770 (N_24770,N_22727,N_22266);
nand U24771 (N_24771,N_22970,N_22829);
nand U24772 (N_24772,N_23995,N_23148);
and U24773 (N_24773,N_23965,N_23365);
nand U24774 (N_24774,N_22412,N_23103);
xor U24775 (N_24775,N_23485,N_22037);
nor U24776 (N_24776,N_22690,N_22306);
and U24777 (N_24777,N_23121,N_22944);
or U24778 (N_24778,N_22621,N_22356);
and U24779 (N_24779,N_23010,N_22117);
or U24780 (N_24780,N_23830,N_22744);
xnor U24781 (N_24781,N_23989,N_22501);
nor U24782 (N_24782,N_23312,N_23117);
xnor U24783 (N_24783,N_23837,N_22381);
and U24784 (N_24784,N_22104,N_22110);
nand U24785 (N_24785,N_22932,N_22694);
nand U24786 (N_24786,N_23843,N_22354);
nor U24787 (N_24787,N_22451,N_23427);
and U24788 (N_24788,N_22904,N_22974);
xnor U24789 (N_24789,N_23672,N_23451);
nand U24790 (N_24790,N_22848,N_22467);
xor U24791 (N_24791,N_22753,N_22708);
xor U24792 (N_24792,N_23296,N_23415);
nor U24793 (N_24793,N_22184,N_23889);
or U24794 (N_24794,N_22421,N_22750);
or U24795 (N_24795,N_22863,N_22998);
xnor U24796 (N_24796,N_22001,N_23422);
nand U24797 (N_24797,N_22986,N_22875);
xnor U24798 (N_24798,N_23527,N_23713);
nand U24799 (N_24799,N_23933,N_22442);
xnor U24800 (N_24800,N_22966,N_23328);
xor U24801 (N_24801,N_23512,N_22726);
xnor U24802 (N_24802,N_23865,N_23919);
and U24803 (N_24803,N_23088,N_22546);
xnor U24804 (N_24804,N_23715,N_23894);
xor U24805 (N_24805,N_23375,N_23060);
nor U24806 (N_24806,N_23151,N_22214);
or U24807 (N_24807,N_23517,N_22108);
nand U24808 (N_24808,N_22260,N_22689);
or U24809 (N_24809,N_22116,N_23430);
and U24810 (N_24810,N_22898,N_22359);
or U24811 (N_24811,N_23746,N_22364);
xor U24812 (N_24812,N_22195,N_23032);
xor U24813 (N_24813,N_23428,N_23085);
nand U24814 (N_24814,N_23737,N_23411);
and U24815 (N_24815,N_22144,N_23124);
nor U24816 (N_24816,N_23582,N_22013);
xor U24817 (N_24817,N_23833,N_22568);
nor U24818 (N_24818,N_23775,N_23788);
and U24819 (N_24819,N_22231,N_22452);
or U24820 (N_24820,N_23891,N_22199);
xnor U24821 (N_24821,N_22168,N_23064);
nand U24822 (N_24822,N_23878,N_23664);
or U24823 (N_24823,N_22157,N_22112);
and U24824 (N_24824,N_23866,N_22815);
and U24825 (N_24825,N_22779,N_23874);
nor U24826 (N_24826,N_22814,N_23846);
nand U24827 (N_24827,N_22735,N_23248);
nand U24828 (N_24828,N_22200,N_23957);
and U24829 (N_24829,N_23294,N_23662);
xnor U24830 (N_24830,N_23694,N_23718);
nand U24831 (N_24831,N_23774,N_23908);
or U24832 (N_24832,N_22832,N_22353);
nand U24833 (N_24833,N_23290,N_22555);
and U24834 (N_24834,N_23229,N_22877);
and U24835 (N_24835,N_23571,N_22311);
xor U24836 (N_24836,N_23281,N_22047);
nor U24837 (N_24837,N_23716,N_23642);
nand U24838 (N_24838,N_23911,N_22468);
and U24839 (N_24839,N_22106,N_22018);
xor U24840 (N_24840,N_23235,N_23745);
and U24841 (N_24841,N_22760,N_22409);
and U24842 (N_24842,N_22243,N_23925);
nor U24843 (N_24843,N_22536,N_22747);
or U24844 (N_24844,N_23511,N_22597);
or U24845 (N_24845,N_23385,N_22713);
and U24846 (N_24846,N_22580,N_23951);
nor U24847 (N_24847,N_23794,N_22620);
nor U24848 (N_24848,N_22569,N_23384);
xor U24849 (N_24849,N_22864,N_23106);
xor U24850 (N_24850,N_22141,N_22533);
and U24851 (N_24851,N_22741,N_22191);
nor U24852 (N_24852,N_22121,N_22437);
nor U24853 (N_24853,N_23755,N_22890);
nor U24854 (N_24854,N_22000,N_22634);
nand U24855 (N_24855,N_22825,N_22699);
xor U24856 (N_24856,N_23293,N_23882);
nor U24857 (N_24857,N_22217,N_23605);
xor U24858 (N_24858,N_23173,N_23174);
and U24859 (N_24859,N_22424,N_23112);
and U24860 (N_24860,N_23622,N_23283);
nand U24861 (N_24861,N_23691,N_22728);
or U24862 (N_24862,N_22413,N_23777);
nor U24863 (N_24863,N_23549,N_23149);
and U24864 (N_24864,N_22849,N_22789);
xor U24865 (N_24865,N_22812,N_22073);
or U24866 (N_24866,N_23172,N_22330);
xnor U24867 (N_24867,N_22816,N_22827);
and U24868 (N_24868,N_22262,N_23481);
nand U24869 (N_24869,N_22352,N_22695);
nand U24870 (N_24870,N_23011,N_22640);
and U24871 (N_24871,N_23603,N_23567);
and U24872 (N_24872,N_22142,N_22361);
and U24873 (N_24873,N_22212,N_22040);
nor U24874 (N_24874,N_23025,N_22017);
or U24875 (N_24875,N_23074,N_22150);
xnor U24876 (N_24876,N_22044,N_23276);
or U24877 (N_24877,N_22787,N_22596);
nor U24878 (N_24878,N_23156,N_23039);
and U24879 (N_24879,N_23961,N_23888);
nand U24880 (N_24880,N_23288,N_23000);
and U24881 (N_24881,N_22562,N_22847);
nand U24882 (N_24882,N_22876,N_23202);
and U24883 (N_24883,N_23851,N_23395);
xnor U24884 (N_24884,N_22678,N_22891);
or U24885 (N_24885,N_22758,N_22072);
xor U24886 (N_24886,N_23224,N_23033);
or U24887 (N_24887,N_23003,N_22936);
or U24888 (N_24888,N_23146,N_22325);
nand U24889 (N_24889,N_22869,N_23783);
nand U24890 (N_24890,N_23359,N_22933);
xnor U24891 (N_24891,N_22531,N_22091);
nor U24892 (N_24892,N_23418,N_23591);
nor U24893 (N_24893,N_22366,N_22673);
and U24894 (N_24894,N_23577,N_22164);
xor U24895 (N_24895,N_23760,N_23308);
or U24896 (N_24896,N_23097,N_23729);
or U24897 (N_24897,N_22668,N_23850);
nand U24898 (N_24898,N_23613,N_23639);
xor U24899 (N_24899,N_23927,N_23388);
nand U24900 (N_24900,N_22271,N_23043);
nand U24901 (N_24901,N_23732,N_22868);
and U24902 (N_24902,N_22189,N_22093);
or U24903 (N_24903,N_22576,N_22530);
or U24904 (N_24904,N_23138,N_23091);
nor U24905 (N_24905,N_22258,N_22703);
nor U24906 (N_24906,N_22518,N_23545);
xor U24907 (N_24907,N_23247,N_22996);
nor U24908 (N_24908,N_22120,N_22036);
xor U24909 (N_24909,N_23323,N_23500);
xnor U24910 (N_24910,N_23667,N_23723);
xor U24911 (N_24911,N_22654,N_22967);
xor U24912 (N_24912,N_22773,N_22405);
or U24913 (N_24913,N_23152,N_23941);
xnor U24914 (N_24914,N_23061,N_22343);
nor U24915 (N_24915,N_22454,N_22188);
nand U24916 (N_24916,N_22056,N_22407);
and U24917 (N_24917,N_23781,N_23966);
or U24918 (N_24918,N_23496,N_23122);
and U24919 (N_24919,N_22504,N_22171);
and U24920 (N_24920,N_23805,N_23461);
xnor U24921 (N_24921,N_23457,N_23928);
and U24922 (N_24922,N_23942,N_22099);
nand U24923 (N_24923,N_22494,N_23905);
xor U24924 (N_24924,N_23178,N_22230);
nand U24925 (N_24925,N_23499,N_23540);
nor U24926 (N_24926,N_22493,N_23740);
and U24927 (N_24927,N_23712,N_23471);
xnor U24928 (N_24928,N_22186,N_22349);
xor U24929 (N_24929,N_22715,N_23371);
and U24930 (N_24930,N_22916,N_22777);
nor U24931 (N_24931,N_23350,N_23104);
xor U24932 (N_24932,N_23763,N_23855);
and U24933 (N_24933,N_23407,N_22638);
and U24934 (N_24934,N_23505,N_23068);
or U24935 (N_24935,N_22528,N_23095);
nand U24936 (N_24936,N_23709,N_22783);
nand U24937 (N_24937,N_22975,N_22021);
xor U24938 (N_24938,N_23623,N_22985);
nand U24939 (N_24939,N_22321,N_22734);
or U24940 (N_24940,N_22224,N_22490);
and U24941 (N_24941,N_22732,N_23394);
xnor U24942 (N_24942,N_23902,N_22439);
and U24943 (N_24943,N_22666,N_22163);
or U24944 (N_24944,N_22363,N_23398);
and U24945 (N_24945,N_22026,N_23769);
nor U24946 (N_24946,N_23488,N_23532);
xnor U24947 (N_24947,N_22588,N_23832);
xor U24948 (N_24948,N_22213,N_23473);
or U24949 (N_24949,N_23839,N_22598);
xnor U24950 (N_24950,N_22283,N_22272);
or U24951 (N_24951,N_23711,N_22920);
and U24952 (N_24952,N_22806,N_23800);
nand U24953 (N_24953,N_22152,N_22924);
xor U24954 (N_24954,N_22318,N_23476);
or U24955 (N_24955,N_23197,N_23372);
nand U24956 (N_24956,N_22883,N_22901);
and U24957 (N_24957,N_23078,N_23543);
and U24958 (N_24958,N_22166,N_23114);
and U24959 (N_24959,N_22105,N_23707);
and U24960 (N_24960,N_23784,N_22866);
nand U24961 (N_24961,N_23378,N_23792);
nor U24962 (N_24962,N_23327,N_22605);
xnor U24963 (N_24963,N_22764,N_22215);
nor U24964 (N_24964,N_23392,N_22820);
xor U24965 (N_24965,N_23968,N_23004);
xor U24966 (N_24966,N_23449,N_23416);
xor U24967 (N_24967,N_23195,N_23326);
xnor U24968 (N_24968,N_23632,N_23400);
nor U24969 (N_24969,N_23510,N_23162);
and U24970 (N_24970,N_22511,N_22992);
and U24971 (N_24971,N_23215,N_23069);
nor U24972 (N_24972,N_23710,N_23383);
and U24973 (N_24973,N_22365,N_22071);
and U24974 (N_24974,N_23193,N_22516);
nor U24975 (N_24975,N_22615,N_22372);
nor U24976 (N_24976,N_23749,N_22799);
xnor U24977 (N_24977,N_23787,N_22172);
nor U24978 (N_24978,N_22733,N_22810);
xor U24979 (N_24979,N_23291,N_22492);
nand U24980 (N_24980,N_23842,N_23330);
nand U24981 (N_24981,N_22507,N_23469);
and U24982 (N_24982,N_22391,N_23964);
and U24983 (N_24983,N_22291,N_22786);
or U24984 (N_24984,N_23474,N_22313);
nor U24985 (N_24985,N_23181,N_22049);
nor U24986 (N_24986,N_22458,N_23002);
xnor U24987 (N_24987,N_23250,N_22367);
nor U24988 (N_24988,N_23401,N_22805);
nand U24989 (N_24989,N_23344,N_23873);
xnor U24990 (N_24990,N_22316,N_22675);
or U24991 (N_24991,N_23226,N_23946);
nor U24992 (N_24992,N_22101,N_22497);
nor U24993 (N_24993,N_23515,N_22994);
nor U24994 (N_24994,N_22745,N_23094);
nor U24995 (N_24995,N_22683,N_22859);
or U24996 (N_24996,N_23259,N_23058);
or U24997 (N_24997,N_23875,N_22669);
nand U24998 (N_24998,N_23431,N_23714);
nor U24999 (N_24999,N_23766,N_23704);
xnor U25000 (N_25000,N_23759,N_22878);
nor U25001 (N_25001,N_22139,N_23321);
nor U25002 (N_25002,N_22016,N_22620);
or U25003 (N_25003,N_22718,N_23069);
xnor U25004 (N_25004,N_22676,N_22844);
xor U25005 (N_25005,N_22540,N_22766);
nor U25006 (N_25006,N_23085,N_22094);
or U25007 (N_25007,N_22414,N_22130);
or U25008 (N_25008,N_22089,N_22684);
nor U25009 (N_25009,N_22766,N_22402);
xnor U25010 (N_25010,N_22571,N_22867);
and U25011 (N_25011,N_23661,N_23068);
nand U25012 (N_25012,N_23638,N_23691);
xnor U25013 (N_25013,N_23614,N_22268);
or U25014 (N_25014,N_22687,N_23472);
and U25015 (N_25015,N_22881,N_23615);
xnor U25016 (N_25016,N_22794,N_22784);
and U25017 (N_25017,N_23117,N_23418);
xnor U25018 (N_25018,N_22761,N_23727);
nor U25019 (N_25019,N_23085,N_22630);
or U25020 (N_25020,N_23169,N_23938);
and U25021 (N_25021,N_22675,N_22656);
nor U25022 (N_25022,N_22662,N_22405);
xor U25023 (N_25023,N_23817,N_23413);
or U25024 (N_25024,N_23824,N_22687);
and U25025 (N_25025,N_22099,N_22647);
or U25026 (N_25026,N_23252,N_22938);
nor U25027 (N_25027,N_22255,N_23454);
and U25028 (N_25028,N_22089,N_23635);
nor U25029 (N_25029,N_23088,N_22050);
and U25030 (N_25030,N_22215,N_23927);
nor U25031 (N_25031,N_22911,N_22582);
xor U25032 (N_25032,N_22662,N_22001);
nor U25033 (N_25033,N_22233,N_23102);
xor U25034 (N_25034,N_23265,N_23291);
and U25035 (N_25035,N_23947,N_23681);
nor U25036 (N_25036,N_23414,N_23329);
xor U25037 (N_25037,N_22964,N_23354);
or U25038 (N_25038,N_23013,N_23079);
xor U25039 (N_25039,N_23638,N_22754);
or U25040 (N_25040,N_23924,N_23476);
xnor U25041 (N_25041,N_23653,N_23911);
and U25042 (N_25042,N_22886,N_22066);
nor U25043 (N_25043,N_22676,N_22615);
and U25044 (N_25044,N_22375,N_23335);
and U25045 (N_25045,N_22994,N_23512);
and U25046 (N_25046,N_22454,N_22408);
and U25047 (N_25047,N_22473,N_23019);
and U25048 (N_25048,N_23648,N_23078);
nor U25049 (N_25049,N_23439,N_22455);
nand U25050 (N_25050,N_23581,N_22824);
or U25051 (N_25051,N_23518,N_23125);
or U25052 (N_25052,N_23230,N_23456);
nor U25053 (N_25053,N_23813,N_23877);
and U25054 (N_25054,N_22056,N_23918);
nor U25055 (N_25055,N_23997,N_22494);
or U25056 (N_25056,N_23662,N_22894);
or U25057 (N_25057,N_22896,N_23387);
nor U25058 (N_25058,N_22935,N_22036);
or U25059 (N_25059,N_22924,N_23810);
or U25060 (N_25060,N_22044,N_22497);
xnor U25061 (N_25061,N_23778,N_22607);
nor U25062 (N_25062,N_22625,N_23235);
nand U25063 (N_25063,N_23067,N_23341);
or U25064 (N_25064,N_22307,N_22634);
and U25065 (N_25065,N_22387,N_23659);
and U25066 (N_25066,N_22989,N_23426);
nor U25067 (N_25067,N_23229,N_23900);
and U25068 (N_25068,N_23585,N_23710);
or U25069 (N_25069,N_23097,N_22080);
or U25070 (N_25070,N_23378,N_23835);
nand U25071 (N_25071,N_23535,N_22272);
or U25072 (N_25072,N_22978,N_23222);
and U25073 (N_25073,N_22395,N_22065);
xnor U25074 (N_25074,N_22306,N_22219);
and U25075 (N_25075,N_22400,N_23317);
xor U25076 (N_25076,N_23354,N_23583);
and U25077 (N_25077,N_22510,N_22456);
and U25078 (N_25078,N_23711,N_22086);
nand U25079 (N_25079,N_23939,N_23747);
xnor U25080 (N_25080,N_23096,N_22350);
and U25081 (N_25081,N_22306,N_23154);
or U25082 (N_25082,N_22040,N_23103);
xor U25083 (N_25083,N_22572,N_23210);
nor U25084 (N_25084,N_23437,N_22399);
xnor U25085 (N_25085,N_23623,N_22816);
and U25086 (N_25086,N_23593,N_23705);
and U25087 (N_25087,N_23006,N_22759);
xor U25088 (N_25088,N_22019,N_23661);
nor U25089 (N_25089,N_23452,N_23706);
xor U25090 (N_25090,N_22695,N_22721);
nand U25091 (N_25091,N_22558,N_22778);
xor U25092 (N_25092,N_22039,N_22364);
nand U25093 (N_25093,N_23443,N_23119);
nand U25094 (N_25094,N_22525,N_23228);
and U25095 (N_25095,N_23188,N_22496);
or U25096 (N_25096,N_23448,N_22348);
nor U25097 (N_25097,N_22475,N_23685);
nor U25098 (N_25098,N_23246,N_22425);
and U25099 (N_25099,N_22576,N_23609);
and U25100 (N_25100,N_22395,N_23191);
and U25101 (N_25101,N_23542,N_22256);
xnor U25102 (N_25102,N_22532,N_22463);
or U25103 (N_25103,N_22616,N_22739);
or U25104 (N_25104,N_22990,N_22793);
nand U25105 (N_25105,N_22598,N_23913);
and U25106 (N_25106,N_22389,N_22458);
nor U25107 (N_25107,N_23563,N_22407);
xor U25108 (N_25108,N_22104,N_23408);
nor U25109 (N_25109,N_23187,N_23108);
or U25110 (N_25110,N_22003,N_23148);
nand U25111 (N_25111,N_23246,N_22444);
and U25112 (N_25112,N_22401,N_22903);
and U25113 (N_25113,N_22122,N_23822);
and U25114 (N_25114,N_22561,N_23693);
xnor U25115 (N_25115,N_23162,N_23580);
nand U25116 (N_25116,N_23809,N_22692);
nor U25117 (N_25117,N_23391,N_22935);
nor U25118 (N_25118,N_23573,N_23781);
xor U25119 (N_25119,N_22061,N_23774);
and U25120 (N_25120,N_23349,N_23362);
or U25121 (N_25121,N_22484,N_23324);
xor U25122 (N_25122,N_23605,N_23879);
nand U25123 (N_25123,N_22113,N_22855);
and U25124 (N_25124,N_23398,N_22723);
nand U25125 (N_25125,N_22479,N_22250);
xor U25126 (N_25126,N_23253,N_23487);
xor U25127 (N_25127,N_23159,N_22963);
and U25128 (N_25128,N_22240,N_22871);
nor U25129 (N_25129,N_23633,N_23186);
and U25130 (N_25130,N_22734,N_22139);
and U25131 (N_25131,N_22349,N_23942);
or U25132 (N_25132,N_22059,N_23708);
nand U25133 (N_25133,N_22730,N_23164);
nand U25134 (N_25134,N_22617,N_23812);
xnor U25135 (N_25135,N_22497,N_23796);
and U25136 (N_25136,N_23485,N_22650);
nand U25137 (N_25137,N_23717,N_23368);
and U25138 (N_25138,N_22988,N_23628);
xor U25139 (N_25139,N_22422,N_23412);
nor U25140 (N_25140,N_23034,N_22842);
nor U25141 (N_25141,N_22676,N_22910);
nand U25142 (N_25142,N_23015,N_23506);
or U25143 (N_25143,N_23476,N_22128);
xor U25144 (N_25144,N_23674,N_23082);
nand U25145 (N_25145,N_23749,N_22034);
nor U25146 (N_25146,N_23521,N_23524);
nand U25147 (N_25147,N_23245,N_23930);
nor U25148 (N_25148,N_22602,N_22597);
and U25149 (N_25149,N_22186,N_22486);
and U25150 (N_25150,N_22647,N_23951);
and U25151 (N_25151,N_23319,N_22287);
or U25152 (N_25152,N_22389,N_22323);
nor U25153 (N_25153,N_23266,N_23656);
nor U25154 (N_25154,N_23659,N_22562);
or U25155 (N_25155,N_23178,N_23473);
and U25156 (N_25156,N_22396,N_22731);
nand U25157 (N_25157,N_23721,N_23263);
and U25158 (N_25158,N_22812,N_22159);
nand U25159 (N_25159,N_22848,N_22581);
nor U25160 (N_25160,N_23845,N_23790);
nor U25161 (N_25161,N_23093,N_22650);
nand U25162 (N_25162,N_22388,N_23548);
nor U25163 (N_25163,N_23392,N_23681);
and U25164 (N_25164,N_23998,N_23599);
nor U25165 (N_25165,N_22009,N_23829);
or U25166 (N_25166,N_22151,N_22132);
xor U25167 (N_25167,N_22857,N_22243);
and U25168 (N_25168,N_23865,N_22501);
nand U25169 (N_25169,N_22521,N_22569);
or U25170 (N_25170,N_23653,N_22917);
or U25171 (N_25171,N_23758,N_23417);
xnor U25172 (N_25172,N_22467,N_23321);
xnor U25173 (N_25173,N_22941,N_23601);
xnor U25174 (N_25174,N_23874,N_23166);
xnor U25175 (N_25175,N_23197,N_23677);
nand U25176 (N_25176,N_23841,N_22387);
xor U25177 (N_25177,N_23290,N_23480);
nand U25178 (N_25178,N_22154,N_22409);
xnor U25179 (N_25179,N_22331,N_23089);
xor U25180 (N_25180,N_22656,N_23055);
nor U25181 (N_25181,N_22466,N_22022);
xnor U25182 (N_25182,N_22640,N_23264);
nor U25183 (N_25183,N_22669,N_23285);
nor U25184 (N_25184,N_23728,N_23245);
or U25185 (N_25185,N_22392,N_22474);
nand U25186 (N_25186,N_22534,N_23181);
nand U25187 (N_25187,N_22341,N_23955);
xnor U25188 (N_25188,N_22167,N_23963);
nor U25189 (N_25189,N_22300,N_23926);
xor U25190 (N_25190,N_22434,N_22221);
nand U25191 (N_25191,N_23263,N_22349);
and U25192 (N_25192,N_23074,N_22054);
xor U25193 (N_25193,N_22925,N_23200);
or U25194 (N_25194,N_23809,N_22720);
or U25195 (N_25195,N_23381,N_23410);
and U25196 (N_25196,N_23169,N_23848);
nor U25197 (N_25197,N_23100,N_22045);
or U25198 (N_25198,N_23503,N_23959);
and U25199 (N_25199,N_22926,N_23030);
nand U25200 (N_25200,N_22847,N_23835);
or U25201 (N_25201,N_23453,N_23069);
nor U25202 (N_25202,N_23742,N_22024);
xnor U25203 (N_25203,N_22340,N_22156);
nor U25204 (N_25204,N_23283,N_22080);
xnor U25205 (N_25205,N_23869,N_22455);
nor U25206 (N_25206,N_23169,N_23721);
xnor U25207 (N_25207,N_23751,N_23292);
or U25208 (N_25208,N_22984,N_22424);
or U25209 (N_25209,N_23841,N_23493);
and U25210 (N_25210,N_23287,N_22342);
or U25211 (N_25211,N_23191,N_23808);
xnor U25212 (N_25212,N_23235,N_22523);
or U25213 (N_25213,N_23312,N_22034);
nand U25214 (N_25214,N_23397,N_22968);
and U25215 (N_25215,N_22215,N_22958);
and U25216 (N_25216,N_23021,N_22836);
nand U25217 (N_25217,N_23910,N_22978);
nor U25218 (N_25218,N_23519,N_22549);
nor U25219 (N_25219,N_23168,N_23145);
or U25220 (N_25220,N_22527,N_23631);
or U25221 (N_25221,N_23058,N_23299);
xor U25222 (N_25222,N_23470,N_23186);
xor U25223 (N_25223,N_23146,N_22198);
and U25224 (N_25224,N_23426,N_22084);
xnor U25225 (N_25225,N_22054,N_23707);
nand U25226 (N_25226,N_22782,N_22705);
nand U25227 (N_25227,N_22374,N_23462);
nand U25228 (N_25228,N_22292,N_22597);
xor U25229 (N_25229,N_23338,N_23331);
or U25230 (N_25230,N_22960,N_23223);
nor U25231 (N_25231,N_23678,N_23028);
nand U25232 (N_25232,N_22520,N_22879);
nor U25233 (N_25233,N_23833,N_23539);
nand U25234 (N_25234,N_22196,N_23789);
xnor U25235 (N_25235,N_23490,N_23744);
xnor U25236 (N_25236,N_22789,N_22142);
or U25237 (N_25237,N_22329,N_23464);
nor U25238 (N_25238,N_22980,N_23283);
and U25239 (N_25239,N_23154,N_23280);
nand U25240 (N_25240,N_22867,N_22445);
nand U25241 (N_25241,N_23733,N_22225);
xor U25242 (N_25242,N_22516,N_22256);
nor U25243 (N_25243,N_23934,N_22107);
nand U25244 (N_25244,N_23249,N_23152);
nor U25245 (N_25245,N_23390,N_22156);
nand U25246 (N_25246,N_23669,N_22488);
and U25247 (N_25247,N_23971,N_23231);
or U25248 (N_25248,N_22019,N_23936);
and U25249 (N_25249,N_22808,N_23306);
or U25250 (N_25250,N_22436,N_22889);
nor U25251 (N_25251,N_23319,N_22718);
nand U25252 (N_25252,N_22899,N_23515);
xnor U25253 (N_25253,N_23454,N_23534);
nor U25254 (N_25254,N_23596,N_22582);
or U25255 (N_25255,N_22836,N_22426);
and U25256 (N_25256,N_23392,N_22272);
xnor U25257 (N_25257,N_23484,N_23862);
and U25258 (N_25258,N_22707,N_22006);
nor U25259 (N_25259,N_23313,N_23304);
nor U25260 (N_25260,N_22929,N_22596);
nor U25261 (N_25261,N_23517,N_22204);
nor U25262 (N_25262,N_22458,N_22374);
xor U25263 (N_25263,N_22017,N_22792);
and U25264 (N_25264,N_23037,N_23556);
or U25265 (N_25265,N_22002,N_23918);
nand U25266 (N_25266,N_22916,N_22719);
xor U25267 (N_25267,N_22234,N_23149);
and U25268 (N_25268,N_23164,N_23143);
nor U25269 (N_25269,N_23218,N_23924);
nand U25270 (N_25270,N_23957,N_23259);
nor U25271 (N_25271,N_22604,N_23945);
nand U25272 (N_25272,N_22091,N_23642);
and U25273 (N_25273,N_23854,N_23200);
and U25274 (N_25274,N_23765,N_22152);
nor U25275 (N_25275,N_23548,N_22772);
xor U25276 (N_25276,N_23844,N_23472);
xor U25277 (N_25277,N_23504,N_23405);
nor U25278 (N_25278,N_22026,N_23476);
nor U25279 (N_25279,N_22398,N_23260);
or U25280 (N_25280,N_23755,N_23513);
nand U25281 (N_25281,N_23444,N_23723);
xor U25282 (N_25282,N_22411,N_22238);
xnor U25283 (N_25283,N_23524,N_23219);
nand U25284 (N_25284,N_22331,N_22785);
or U25285 (N_25285,N_22128,N_22962);
nor U25286 (N_25286,N_22456,N_23686);
nand U25287 (N_25287,N_23383,N_22162);
or U25288 (N_25288,N_23738,N_23141);
or U25289 (N_25289,N_22627,N_22710);
and U25290 (N_25290,N_23917,N_23193);
nand U25291 (N_25291,N_23503,N_22619);
and U25292 (N_25292,N_22597,N_23502);
nor U25293 (N_25293,N_23337,N_22756);
nand U25294 (N_25294,N_22354,N_22376);
xor U25295 (N_25295,N_22519,N_22910);
and U25296 (N_25296,N_23720,N_22761);
xor U25297 (N_25297,N_23570,N_23643);
xor U25298 (N_25298,N_23738,N_22400);
nor U25299 (N_25299,N_22364,N_23463);
xor U25300 (N_25300,N_23778,N_22425);
xnor U25301 (N_25301,N_23943,N_22121);
xor U25302 (N_25302,N_23593,N_23576);
nor U25303 (N_25303,N_23305,N_23952);
nor U25304 (N_25304,N_23697,N_22810);
xnor U25305 (N_25305,N_22107,N_23064);
or U25306 (N_25306,N_22199,N_23947);
and U25307 (N_25307,N_22149,N_22398);
nor U25308 (N_25308,N_23673,N_22289);
xor U25309 (N_25309,N_23494,N_23061);
nor U25310 (N_25310,N_22063,N_23271);
nand U25311 (N_25311,N_23714,N_23112);
or U25312 (N_25312,N_23670,N_23432);
and U25313 (N_25313,N_23965,N_23240);
nand U25314 (N_25314,N_22340,N_22242);
nand U25315 (N_25315,N_23901,N_23761);
nand U25316 (N_25316,N_22440,N_23369);
xor U25317 (N_25317,N_22479,N_23708);
and U25318 (N_25318,N_22331,N_23828);
nor U25319 (N_25319,N_23544,N_22900);
or U25320 (N_25320,N_23137,N_22707);
nand U25321 (N_25321,N_22432,N_23859);
nand U25322 (N_25322,N_22922,N_22440);
or U25323 (N_25323,N_22840,N_22102);
nor U25324 (N_25324,N_23527,N_22732);
or U25325 (N_25325,N_22029,N_23440);
xor U25326 (N_25326,N_23310,N_22973);
nor U25327 (N_25327,N_23934,N_22329);
nand U25328 (N_25328,N_23490,N_22333);
xor U25329 (N_25329,N_23543,N_23200);
nor U25330 (N_25330,N_22048,N_22832);
or U25331 (N_25331,N_22230,N_22578);
nor U25332 (N_25332,N_22782,N_22387);
and U25333 (N_25333,N_22251,N_22793);
and U25334 (N_25334,N_22931,N_23121);
xnor U25335 (N_25335,N_23453,N_22752);
xnor U25336 (N_25336,N_22758,N_23284);
or U25337 (N_25337,N_23812,N_22475);
or U25338 (N_25338,N_22858,N_22720);
and U25339 (N_25339,N_23411,N_22015);
and U25340 (N_25340,N_23282,N_22011);
nand U25341 (N_25341,N_22570,N_23652);
nor U25342 (N_25342,N_22289,N_22930);
xnor U25343 (N_25343,N_22596,N_23135);
nor U25344 (N_25344,N_22701,N_22278);
or U25345 (N_25345,N_23566,N_22426);
xnor U25346 (N_25346,N_23187,N_23519);
nand U25347 (N_25347,N_22334,N_23154);
nor U25348 (N_25348,N_23484,N_23805);
xor U25349 (N_25349,N_23873,N_23475);
or U25350 (N_25350,N_22164,N_22358);
or U25351 (N_25351,N_23105,N_23619);
and U25352 (N_25352,N_23992,N_23477);
and U25353 (N_25353,N_23528,N_23365);
or U25354 (N_25354,N_23560,N_22957);
nand U25355 (N_25355,N_22980,N_22879);
nand U25356 (N_25356,N_22165,N_23373);
and U25357 (N_25357,N_23850,N_22901);
nor U25358 (N_25358,N_22579,N_23009);
or U25359 (N_25359,N_23471,N_22736);
and U25360 (N_25360,N_22178,N_22869);
or U25361 (N_25361,N_23410,N_22871);
xnor U25362 (N_25362,N_23939,N_23290);
xnor U25363 (N_25363,N_23351,N_22811);
or U25364 (N_25364,N_23328,N_23097);
nor U25365 (N_25365,N_23476,N_22357);
or U25366 (N_25366,N_23881,N_23281);
nand U25367 (N_25367,N_22604,N_23446);
xor U25368 (N_25368,N_23276,N_23460);
nor U25369 (N_25369,N_22033,N_22629);
and U25370 (N_25370,N_23745,N_22961);
and U25371 (N_25371,N_23162,N_22417);
and U25372 (N_25372,N_22407,N_23450);
xnor U25373 (N_25373,N_23067,N_22076);
or U25374 (N_25374,N_22082,N_22461);
or U25375 (N_25375,N_23953,N_22328);
and U25376 (N_25376,N_23935,N_23524);
nor U25377 (N_25377,N_22859,N_23798);
or U25378 (N_25378,N_22146,N_22752);
nor U25379 (N_25379,N_22819,N_22127);
nand U25380 (N_25380,N_23859,N_22047);
nand U25381 (N_25381,N_22123,N_23316);
and U25382 (N_25382,N_22901,N_22922);
xnor U25383 (N_25383,N_23683,N_23839);
nand U25384 (N_25384,N_22052,N_23797);
or U25385 (N_25385,N_22987,N_23942);
xnor U25386 (N_25386,N_22309,N_23800);
nor U25387 (N_25387,N_22976,N_23667);
nand U25388 (N_25388,N_22113,N_22492);
nor U25389 (N_25389,N_23859,N_23977);
and U25390 (N_25390,N_23094,N_22053);
xnor U25391 (N_25391,N_22670,N_23742);
or U25392 (N_25392,N_22544,N_23184);
or U25393 (N_25393,N_23796,N_23500);
or U25394 (N_25394,N_22554,N_23971);
nand U25395 (N_25395,N_22065,N_23226);
nor U25396 (N_25396,N_22343,N_22662);
and U25397 (N_25397,N_22358,N_23843);
or U25398 (N_25398,N_22834,N_22942);
or U25399 (N_25399,N_23356,N_23916);
xor U25400 (N_25400,N_23640,N_22187);
nor U25401 (N_25401,N_23089,N_22440);
and U25402 (N_25402,N_23551,N_22271);
and U25403 (N_25403,N_23813,N_22299);
or U25404 (N_25404,N_23582,N_23971);
or U25405 (N_25405,N_22632,N_23367);
xor U25406 (N_25406,N_22720,N_22860);
xor U25407 (N_25407,N_23957,N_22765);
nor U25408 (N_25408,N_22963,N_23498);
and U25409 (N_25409,N_23656,N_23139);
nor U25410 (N_25410,N_22756,N_22758);
nor U25411 (N_25411,N_23859,N_23866);
and U25412 (N_25412,N_22380,N_22813);
nand U25413 (N_25413,N_23012,N_23563);
or U25414 (N_25414,N_22401,N_23769);
or U25415 (N_25415,N_23879,N_23249);
nand U25416 (N_25416,N_23202,N_23857);
xor U25417 (N_25417,N_23405,N_22830);
and U25418 (N_25418,N_22684,N_22658);
or U25419 (N_25419,N_23339,N_23478);
and U25420 (N_25420,N_23986,N_22164);
or U25421 (N_25421,N_23060,N_22192);
xor U25422 (N_25422,N_23519,N_22265);
nand U25423 (N_25423,N_22020,N_22593);
nor U25424 (N_25424,N_23438,N_23312);
and U25425 (N_25425,N_22193,N_22471);
nor U25426 (N_25426,N_23442,N_23431);
or U25427 (N_25427,N_23335,N_23034);
xor U25428 (N_25428,N_23496,N_23594);
or U25429 (N_25429,N_23173,N_22097);
nor U25430 (N_25430,N_23509,N_23541);
or U25431 (N_25431,N_22450,N_23829);
and U25432 (N_25432,N_22875,N_22402);
or U25433 (N_25433,N_22845,N_22776);
or U25434 (N_25434,N_23239,N_22790);
and U25435 (N_25435,N_23153,N_23834);
or U25436 (N_25436,N_23237,N_23656);
and U25437 (N_25437,N_23542,N_23855);
nor U25438 (N_25438,N_23292,N_22881);
nor U25439 (N_25439,N_22619,N_23273);
xnor U25440 (N_25440,N_22500,N_23528);
xnor U25441 (N_25441,N_22356,N_23615);
and U25442 (N_25442,N_22503,N_23714);
nand U25443 (N_25443,N_23779,N_22235);
nor U25444 (N_25444,N_23856,N_23068);
nand U25445 (N_25445,N_23990,N_22978);
nor U25446 (N_25446,N_22535,N_23918);
nand U25447 (N_25447,N_23143,N_22699);
nor U25448 (N_25448,N_22245,N_22445);
nor U25449 (N_25449,N_23166,N_22842);
or U25450 (N_25450,N_22592,N_22991);
or U25451 (N_25451,N_22178,N_23394);
xor U25452 (N_25452,N_23006,N_22755);
xor U25453 (N_25453,N_23802,N_22478);
or U25454 (N_25454,N_23679,N_22532);
nor U25455 (N_25455,N_22765,N_22939);
nor U25456 (N_25456,N_23052,N_23075);
nand U25457 (N_25457,N_23140,N_23019);
and U25458 (N_25458,N_22280,N_22553);
nor U25459 (N_25459,N_23088,N_23167);
or U25460 (N_25460,N_23566,N_23080);
nand U25461 (N_25461,N_23276,N_22647);
nand U25462 (N_25462,N_23997,N_22659);
and U25463 (N_25463,N_23937,N_22809);
nand U25464 (N_25464,N_22456,N_23313);
nand U25465 (N_25465,N_23884,N_23899);
or U25466 (N_25466,N_23245,N_23206);
nand U25467 (N_25467,N_23923,N_22397);
nand U25468 (N_25468,N_22754,N_22478);
nand U25469 (N_25469,N_23818,N_22809);
xnor U25470 (N_25470,N_23799,N_22334);
xnor U25471 (N_25471,N_23427,N_23318);
or U25472 (N_25472,N_23135,N_22226);
nand U25473 (N_25473,N_22908,N_23550);
and U25474 (N_25474,N_22602,N_23576);
or U25475 (N_25475,N_22908,N_22965);
or U25476 (N_25476,N_23898,N_22201);
and U25477 (N_25477,N_23722,N_22731);
xnor U25478 (N_25478,N_23035,N_22448);
nor U25479 (N_25479,N_22661,N_22215);
nand U25480 (N_25480,N_23658,N_22971);
nor U25481 (N_25481,N_23855,N_23634);
nand U25482 (N_25482,N_23656,N_22314);
nand U25483 (N_25483,N_22756,N_22107);
xnor U25484 (N_25484,N_22646,N_23111);
xnor U25485 (N_25485,N_23167,N_22367);
or U25486 (N_25486,N_22500,N_22030);
or U25487 (N_25487,N_22386,N_23826);
or U25488 (N_25488,N_23268,N_22520);
and U25489 (N_25489,N_23918,N_22417);
and U25490 (N_25490,N_22950,N_23839);
xor U25491 (N_25491,N_23976,N_22708);
nand U25492 (N_25492,N_22758,N_22410);
and U25493 (N_25493,N_22529,N_23538);
nor U25494 (N_25494,N_23614,N_23171);
xor U25495 (N_25495,N_22743,N_23661);
or U25496 (N_25496,N_22019,N_23542);
or U25497 (N_25497,N_22923,N_23283);
xor U25498 (N_25498,N_22536,N_22665);
and U25499 (N_25499,N_23914,N_23257);
nand U25500 (N_25500,N_23791,N_23927);
or U25501 (N_25501,N_23774,N_23880);
nor U25502 (N_25502,N_22326,N_23279);
nand U25503 (N_25503,N_22115,N_23436);
xnor U25504 (N_25504,N_22024,N_22541);
nor U25505 (N_25505,N_22064,N_23650);
nand U25506 (N_25506,N_22319,N_23890);
and U25507 (N_25507,N_23467,N_22524);
xnor U25508 (N_25508,N_22506,N_22407);
or U25509 (N_25509,N_22835,N_23553);
and U25510 (N_25510,N_22678,N_23050);
xor U25511 (N_25511,N_23888,N_23503);
nand U25512 (N_25512,N_22263,N_23128);
xnor U25513 (N_25513,N_23414,N_22941);
nor U25514 (N_25514,N_22177,N_23910);
nand U25515 (N_25515,N_22243,N_22050);
nor U25516 (N_25516,N_23292,N_22447);
nor U25517 (N_25517,N_22478,N_22550);
xnor U25518 (N_25518,N_23935,N_22827);
or U25519 (N_25519,N_23127,N_23787);
nor U25520 (N_25520,N_22841,N_22602);
nand U25521 (N_25521,N_22351,N_23744);
nand U25522 (N_25522,N_22322,N_22686);
or U25523 (N_25523,N_22099,N_23765);
nand U25524 (N_25524,N_23504,N_23541);
nand U25525 (N_25525,N_23022,N_22566);
nand U25526 (N_25526,N_23727,N_22927);
or U25527 (N_25527,N_23608,N_23000);
nand U25528 (N_25528,N_23106,N_22448);
xnor U25529 (N_25529,N_23155,N_23756);
or U25530 (N_25530,N_23787,N_23470);
xor U25531 (N_25531,N_22022,N_23502);
nor U25532 (N_25532,N_22693,N_23929);
xnor U25533 (N_25533,N_23411,N_22809);
and U25534 (N_25534,N_23333,N_23999);
nor U25535 (N_25535,N_22178,N_22701);
or U25536 (N_25536,N_22520,N_22509);
xor U25537 (N_25537,N_22201,N_22446);
nor U25538 (N_25538,N_23119,N_22127);
nand U25539 (N_25539,N_22919,N_23087);
nor U25540 (N_25540,N_22721,N_23004);
xor U25541 (N_25541,N_22265,N_22255);
nor U25542 (N_25542,N_22726,N_23472);
xnor U25543 (N_25543,N_22606,N_22511);
xnor U25544 (N_25544,N_22909,N_22465);
nor U25545 (N_25545,N_23527,N_22914);
nor U25546 (N_25546,N_23226,N_22601);
nand U25547 (N_25547,N_23346,N_23419);
and U25548 (N_25548,N_23340,N_22596);
and U25549 (N_25549,N_22979,N_23313);
or U25550 (N_25550,N_22065,N_23998);
xnor U25551 (N_25551,N_22958,N_22699);
nand U25552 (N_25552,N_22260,N_23475);
or U25553 (N_25553,N_22371,N_23156);
xor U25554 (N_25554,N_22892,N_22496);
or U25555 (N_25555,N_23749,N_22248);
and U25556 (N_25556,N_23886,N_22949);
or U25557 (N_25557,N_22505,N_22164);
xnor U25558 (N_25558,N_23478,N_23042);
nand U25559 (N_25559,N_22288,N_22119);
and U25560 (N_25560,N_22643,N_23084);
nand U25561 (N_25561,N_22828,N_22163);
or U25562 (N_25562,N_23007,N_23615);
and U25563 (N_25563,N_22533,N_22590);
xnor U25564 (N_25564,N_23763,N_23886);
or U25565 (N_25565,N_22708,N_22495);
nand U25566 (N_25566,N_22717,N_22683);
or U25567 (N_25567,N_22290,N_23633);
and U25568 (N_25568,N_23140,N_22361);
nand U25569 (N_25569,N_23559,N_22804);
and U25570 (N_25570,N_22590,N_22414);
xnor U25571 (N_25571,N_23842,N_22098);
nor U25572 (N_25572,N_22674,N_22097);
nand U25573 (N_25573,N_22453,N_23064);
and U25574 (N_25574,N_23283,N_23725);
and U25575 (N_25575,N_22850,N_22437);
and U25576 (N_25576,N_22312,N_23624);
or U25577 (N_25577,N_22793,N_23766);
or U25578 (N_25578,N_23115,N_23558);
nor U25579 (N_25579,N_23419,N_23256);
xnor U25580 (N_25580,N_23442,N_23907);
nor U25581 (N_25581,N_22867,N_22591);
nand U25582 (N_25582,N_23951,N_23983);
or U25583 (N_25583,N_22282,N_22481);
or U25584 (N_25584,N_22994,N_22423);
and U25585 (N_25585,N_22404,N_22826);
or U25586 (N_25586,N_22026,N_22117);
xor U25587 (N_25587,N_23156,N_22234);
nor U25588 (N_25588,N_23671,N_22668);
nand U25589 (N_25589,N_23501,N_22845);
nor U25590 (N_25590,N_23467,N_23060);
nor U25591 (N_25591,N_22715,N_22879);
xor U25592 (N_25592,N_23295,N_22234);
nor U25593 (N_25593,N_22352,N_23145);
nor U25594 (N_25594,N_23147,N_22560);
or U25595 (N_25595,N_23597,N_23464);
xnor U25596 (N_25596,N_23884,N_22565);
or U25597 (N_25597,N_22267,N_23208);
nor U25598 (N_25598,N_23359,N_23700);
nand U25599 (N_25599,N_22753,N_23117);
and U25600 (N_25600,N_23285,N_23306);
and U25601 (N_25601,N_22389,N_22005);
nand U25602 (N_25602,N_22380,N_23481);
xor U25603 (N_25603,N_22512,N_22846);
nand U25604 (N_25604,N_22284,N_23747);
or U25605 (N_25605,N_23371,N_23978);
or U25606 (N_25606,N_23369,N_22562);
and U25607 (N_25607,N_23604,N_22473);
or U25608 (N_25608,N_23192,N_22607);
xnor U25609 (N_25609,N_23276,N_23340);
nand U25610 (N_25610,N_23397,N_22035);
and U25611 (N_25611,N_22474,N_22321);
xor U25612 (N_25612,N_22451,N_22670);
xnor U25613 (N_25613,N_22772,N_22002);
or U25614 (N_25614,N_23392,N_22665);
and U25615 (N_25615,N_22212,N_22086);
or U25616 (N_25616,N_22458,N_22735);
nor U25617 (N_25617,N_22388,N_23448);
nor U25618 (N_25618,N_22122,N_22876);
nor U25619 (N_25619,N_22036,N_23006);
or U25620 (N_25620,N_23411,N_22224);
nor U25621 (N_25621,N_23776,N_23826);
or U25622 (N_25622,N_23754,N_22827);
and U25623 (N_25623,N_22647,N_23275);
nor U25624 (N_25624,N_23070,N_22073);
nand U25625 (N_25625,N_23116,N_23697);
nor U25626 (N_25626,N_23703,N_22370);
xor U25627 (N_25627,N_23872,N_23660);
nor U25628 (N_25628,N_22045,N_22027);
or U25629 (N_25629,N_23987,N_22971);
nand U25630 (N_25630,N_23096,N_23059);
or U25631 (N_25631,N_22132,N_23605);
or U25632 (N_25632,N_23914,N_22152);
nand U25633 (N_25633,N_23183,N_22398);
nor U25634 (N_25634,N_22342,N_22273);
and U25635 (N_25635,N_23236,N_23577);
nor U25636 (N_25636,N_22454,N_22813);
and U25637 (N_25637,N_23502,N_22103);
or U25638 (N_25638,N_22922,N_23782);
or U25639 (N_25639,N_22892,N_22790);
xnor U25640 (N_25640,N_23505,N_22620);
and U25641 (N_25641,N_22391,N_23784);
nor U25642 (N_25642,N_22779,N_23953);
or U25643 (N_25643,N_22655,N_22955);
xor U25644 (N_25644,N_23321,N_22168);
nand U25645 (N_25645,N_22611,N_22840);
xor U25646 (N_25646,N_22106,N_23951);
xnor U25647 (N_25647,N_22606,N_22211);
xnor U25648 (N_25648,N_23296,N_23014);
nand U25649 (N_25649,N_23997,N_22163);
nand U25650 (N_25650,N_23695,N_23548);
and U25651 (N_25651,N_22342,N_22709);
nor U25652 (N_25652,N_23027,N_22665);
nor U25653 (N_25653,N_23117,N_22454);
nor U25654 (N_25654,N_23355,N_23814);
nand U25655 (N_25655,N_22863,N_22826);
nand U25656 (N_25656,N_22156,N_22499);
nand U25657 (N_25657,N_23444,N_22291);
and U25658 (N_25658,N_23785,N_22524);
xnor U25659 (N_25659,N_22856,N_22720);
xor U25660 (N_25660,N_22151,N_23614);
nand U25661 (N_25661,N_22795,N_23442);
or U25662 (N_25662,N_22393,N_23001);
xor U25663 (N_25663,N_22783,N_22335);
or U25664 (N_25664,N_22582,N_23161);
nor U25665 (N_25665,N_23642,N_22673);
or U25666 (N_25666,N_23321,N_22009);
and U25667 (N_25667,N_22215,N_23977);
nand U25668 (N_25668,N_23778,N_22364);
or U25669 (N_25669,N_23791,N_22696);
xor U25670 (N_25670,N_22589,N_23265);
or U25671 (N_25671,N_22120,N_23608);
xor U25672 (N_25672,N_23930,N_22769);
and U25673 (N_25673,N_23812,N_23823);
or U25674 (N_25674,N_23395,N_22373);
xnor U25675 (N_25675,N_22751,N_23505);
xnor U25676 (N_25676,N_22667,N_23836);
nand U25677 (N_25677,N_23947,N_22962);
nor U25678 (N_25678,N_22561,N_23940);
xor U25679 (N_25679,N_22152,N_23153);
xor U25680 (N_25680,N_22879,N_22865);
xor U25681 (N_25681,N_22498,N_22022);
nand U25682 (N_25682,N_23358,N_23233);
xor U25683 (N_25683,N_22857,N_22057);
xor U25684 (N_25684,N_23932,N_23235);
and U25685 (N_25685,N_23200,N_22550);
and U25686 (N_25686,N_22122,N_22497);
nand U25687 (N_25687,N_22800,N_23992);
nand U25688 (N_25688,N_22985,N_23283);
xor U25689 (N_25689,N_23088,N_23073);
xor U25690 (N_25690,N_23484,N_23973);
or U25691 (N_25691,N_23820,N_23083);
or U25692 (N_25692,N_22003,N_23531);
or U25693 (N_25693,N_22347,N_23507);
nor U25694 (N_25694,N_22638,N_22043);
and U25695 (N_25695,N_22170,N_23013);
nand U25696 (N_25696,N_23059,N_22706);
nor U25697 (N_25697,N_23434,N_22715);
or U25698 (N_25698,N_22477,N_23261);
or U25699 (N_25699,N_22849,N_23146);
xor U25700 (N_25700,N_22112,N_23854);
nand U25701 (N_25701,N_22920,N_22806);
nor U25702 (N_25702,N_22391,N_23404);
nor U25703 (N_25703,N_23610,N_23487);
nor U25704 (N_25704,N_22670,N_22501);
and U25705 (N_25705,N_22007,N_22519);
nor U25706 (N_25706,N_23730,N_23102);
nor U25707 (N_25707,N_23519,N_23601);
nor U25708 (N_25708,N_22897,N_22563);
or U25709 (N_25709,N_23205,N_22541);
nand U25710 (N_25710,N_23064,N_22682);
or U25711 (N_25711,N_23275,N_22383);
xnor U25712 (N_25712,N_23708,N_23648);
nor U25713 (N_25713,N_23213,N_23463);
or U25714 (N_25714,N_22710,N_23111);
nor U25715 (N_25715,N_22662,N_22609);
nor U25716 (N_25716,N_23134,N_22392);
nand U25717 (N_25717,N_22353,N_23882);
nand U25718 (N_25718,N_22542,N_22499);
nand U25719 (N_25719,N_22462,N_22955);
and U25720 (N_25720,N_22619,N_22343);
and U25721 (N_25721,N_23024,N_23163);
or U25722 (N_25722,N_22305,N_23316);
and U25723 (N_25723,N_22505,N_22540);
or U25724 (N_25724,N_22643,N_23772);
nor U25725 (N_25725,N_23408,N_22436);
nor U25726 (N_25726,N_23930,N_23198);
nor U25727 (N_25727,N_22031,N_22749);
nor U25728 (N_25728,N_22752,N_22511);
nand U25729 (N_25729,N_23290,N_23469);
or U25730 (N_25730,N_22048,N_23784);
nor U25731 (N_25731,N_23424,N_23007);
and U25732 (N_25732,N_23248,N_22488);
and U25733 (N_25733,N_22911,N_22781);
or U25734 (N_25734,N_22916,N_22260);
and U25735 (N_25735,N_23798,N_23055);
nor U25736 (N_25736,N_23791,N_23505);
nor U25737 (N_25737,N_23923,N_23584);
or U25738 (N_25738,N_22924,N_22156);
nor U25739 (N_25739,N_22878,N_22880);
or U25740 (N_25740,N_22388,N_23934);
nand U25741 (N_25741,N_23710,N_23394);
or U25742 (N_25742,N_22767,N_23983);
nand U25743 (N_25743,N_23678,N_22733);
nor U25744 (N_25744,N_23507,N_22207);
xnor U25745 (N_25745,N_23731,N_23467);
nand U25746 (N_25746,N_22159,N_22903);
or U25747 (N_25747,N_22181,N_23391);
xnor U25748 (N_25748,N_23377,N_23639);
and U25749 (N_25749,N_23036,N_23434);
or U25750 (N_25750,N_23771,N_23764);
xnor U25751 (N_25751,N_23544,N_22555);
nand U25752 (N_25752,N_22929,N_23155);
and U25753 (N_25753,N_23522,N_23991);
nor U25754 (N_25754,N_22917,N_23028);
nor U25755 (N_25755,N_23306,N_22308);
nor U25756 (N_25756,N_23015,N_23825);
nor U25757 (N_25757,N_22663,N_23931);
xor U25758 (N_25758,N_22678,N_23061);
nand U25759 (N_25759,N_23091,N_22625);
or U25760 (N_25760,N_22292,N_22626);
xnor U25761 (N_25761,N_22802,N_22112);
or U25762 (N_25762,N_23657,N_23116);
xor U25763 (N_25763,N_22250,N_22923);
xnor U25764 (N_25764,N_23705,N_22360);
nor U25765 (N_25765,N_23851,N_23199);
nor U25766 (N_25766,N_23633,N_23607);
and U25767 (N_25767,N_22020,N_22786);
or U25768 (N_25768,N_22284,N_23916);
nand U25769 (N_25769,N_23173,N_22228);
nor U25770 (N_25770,N_22826,N_23773);
xor U25771 (N_25771,N_23069,N_23548);
xnor U25772 (N_25772,N_22092,N_22015);
or U25773 (N_25773,N_22044,N_22186);
nor U25774 (N_25774,N_23377,N_22885);
nand U25775 (N_25775,N_22805,N_23109);
nor U25776 (N_25776,N_23614,N_22689);
nor U25777 (N_25777,N_23507,N_23708);
and U25778 (N_25778,N_23099,N_23080);
and U25779 (N_25779,N_23055,N_22910);
nor U25780 (N_25780,N_22211,N_22046);
xnor U25781 (N_25781,N_23791,N_23262);
or U25782 (N_25782,N_22021,N_23166);
or U25783 (N_25783,N_23292,N_23454);
or U25784 (N_25784,N_22088,N_22109);
nand U25785 (N_25785,N_23446,N_22199);
nor U25786 (N_25786,N_23977,N_23858);
or U25787 (N_25787,N_23387,N_22617);
xor U25788 (N_25788,N_22059,N_22129);
nand U25789 (N_25789,N_23456,N_23379);
xor U25790 (N_25790,N_23185,N_22806);
and U25791 (N_25791,N_22719,N_22262);
and U25792 (N_25792,N_22441,N_23425);
nand U25793 (N_25793,N_22185,N_23820);
nor U25794 (N_25794,N_23969,N_23050);
and U25795 (N_25795,N_22117,N_23160);
nand U25796 (N_25796,N_22188,N_23172);
nand U25797 (N_25797,N_22233,N_23261);
and U25798 (N_25798,N_22948,N_22628);
and U25799 (N_25799,N_22315,N_23039);
xnor U25800 (N_25800,N_22291,N_23083);
xnor U25801 (N_25801,N_22156,N_23259);
and U25802 (N_25802,N_22165,N_23472);
nand U25803 (N_25803,N_22219,N_22105);
or U25804 (N_25804,N_23998,N_23874);
nor U25805 (N_25805,N_22879,N_23860);
and U25806 (N_25806,N_22288,N_22293);
nor U25807 (N_25807,N_23768,N_22639);
xor U25808 (N_25808,N_22423,N_22132);
nand U25809 (N_25809,N_22195,N_22086);
nand U25810 (N_25810,N_23196,N_22040);
xor U25811 (N_25811,N_22590,N_22508);
xor U25812 (N_25812,N_22884,N_23170);
nand U25813 (N_25813,N_22229,N_23090);
xor U25814 (N_25814,N_23358,N_23284);
nand U25815 (N_25815,N_22230,N_22309);
nand U25816 (N_25816,N_22692,N_23315);
nor U25817 (N_25817,N_22840,N_22819);
or U25818 (N_25818,N_23410,N_22637);
and U25819 (N_25819,N_22503,N_23347);
and U25820 (N_25820,N_23273,N_23102);
and U25821 (N_25821,N_22122,N_22055);
nand U25822 (N_25822,N_22736,N_22982);
xor U25823 (N_25823,N_22271,N_23864);
xor U25824 (N_25824,N_22498,N_23798);
or U25825 (N_25825,N_23295,N_23903);
nor U25826 (N_25826,N_23371,N_23402);
nand U25827 (N_25827,N_23553,N_23163);
nor U25828 (N_25828,N_22564,N_22209);
nand U25829 (N_25829,N_22401,N_23642);
xor U25830 (N_25830,N_23874,N_23573);
xnor U25831 (N_25831,N_22722,N_23777);
nand U25832 (N_25832,N_23326,N_23651);
or U25833 (N_25833,N_23238,N_22763);
nand U25834 (N_25834,N_23172,N_22113);
and U25835 (N_25835,N_22264,N_23341);
and U25836 (N_25836,N_22128,N_22930);
or U25837 (N_25837,N_23835,N_23044);
nand U25838 (N_25838,N_22043,N_22592);
nor U25839 (N_25839,N_22045,N_22634);
nor U25840 (N_25840,N_22611,N_23397);
or U25841 (N_25841,N_23885,N_23036);
and U25842 (N_25842,N_22791,N_23694);
nor U25843 (N_25843,N_23797,N_23740);
and U25844 (N_25844,N_23811,N_23639);
and U25845 (N_25845,N_23628,N_22096);
or U25846 (N_25846,N_22204,N_23647);
xor U25847 (N_25847,N_22705,N_22119);
nand U25848 (N_25848,N_23139,N_23981);
nor U25849 (N_25849,N_22866,N_23201);
and U25850 (N_25850,N_22831,N_23828);
nand U25851 (N_25851,N_22178,N_22346);
and U25852 (N_25852,N_22368,N_22877);
or U25853 (N_25853,N_22936,N_23790);
nand U25854 (N_25854,N_23593,N_22017);
and U25855 (N_25855,N_22248,N_23196);
nand U25856 (N_25856,N_22506,N_22370);
xor U25857 (N_25857,N_23260,N_22633);
or U25858 (N_25858,N_22407,N_22424);
xor U25859 (N_25859,N_22771,N_22510);
nor U25860 (N_25860,N_23560,N_23847);
nand U25861 (N_25861,N_22464,N_23390);
nor U25862 (N_25862,N_22117,N_23214);
nand U25863 (N_25863,N_22500,N_23022);
and U25864 (N_25864,N_23188,N_23331);
nand U25865 (N_25865,N_23898,N_22579);
or U25866 (N_25866,N_23339,N_23193);
xnor U25867 (N_25867,N_23974,N_23343);
nor U25868 (N_25868,N_23446,N_22963);
and U25869 (N_25869,N_23189,N_23782);
and U25870 (N_25870,N_23706,N_23429);
and U25871 (N_25871,N_23342,N_22336);
nor U25872 (N_25872,N_22558,N_23284);
or U25873 (N_25873,N_22503,N_23281);
and U25874 (N_25874,N_23640,N_22731);
or U25875 (N_25875,N_22103,N_22985);
xor U25876 (N_25876,N_22161,N_23534);
nand U25877 (N_25877,N_23713,N_23323);
or U25878 (N_25878,N_22182,N_22449);
nand U25879 (N_25879,N_23325,N_22300);
nand U25880 (N_25880,N_22116,N_23098);
and U25881 (N_25881,N_22801,N_22323);
xnor U25882 (N_25882,N_23240,N_23632);
nand U25883 (N_25883,N_23784,N_23989);
or U25884 (N_25884,N_23083,N_22779);
and U25885 (N_25885,N_23708,N_23863);
and U25886 (N_25886,N_23832,N_23946);
xnor U25887 (N_25887,N_22855,N_23038);
nand U25888 (N_25888,N_23999,N_22914);
or U25889 (N_25889,N_22622,N_23925);
nor U25890 (N_25890,N_23212,N_22399);
and U25891 (N_25891,N_23066,N_23555);
nand U25892 (N_25892,N_23978,N_22141);
xor U25893 (N_25893,N_22641,N_22344);
nand U25894 (N_25894,N_22112,N_23746);
nor U25895 (N_25895,N_22456,N_22639);
or U25896 (N_25896,N_22166,N_22498);
nand U25897 (N_25897,N_22353,N_23464);
nor U25898 (N_25898,N_23913,N_22086);
nand U25899 (N_25899,N_23132,N_23717);
and U25900 (N_25900,N_23583,N_23070);
or U25901 (N_25901,N_23515,N_23075);
xnor U25902 (N_25902,N_23586,N_22405);
or U25903 (N_25903,N_22535,N_22836);
and U25904 (N_25904,N_22262,N_23606);
nand U25905 (N_25905,N_22616,N_23147);
or U25906 (N_25906,N_22247,N_23728);
nand U25907 (N_25907,N_23259,N_22692);
xnor U25908 (N_25908,N_22530,N_23523);
nand U25909 (N_25909,N_23806,N_23662);
nor U25910 (N_25910,N_22899,N_22965);
xnor U25911 (N_25911,N_22318,N_23447);
nand U25912 (N_25912,N_22355,N_23867);
nand U25913 (N_25913,N_22739,N_23158);
xnor U25914 (N_25914,N_22258,N_22998);
nor U25915 (N_25915,N_22981,N_22014);
nor U25916 (N_25916,N_22567,N_22207);
or U25917 (N_25917,N_23429,N_22680);
xnor U25918 (N_25918,N_22433,N_23268);
xor U25919 (N_25919,N_22996,N_22659);
xor U25920 (N_25920,N_23752,N_22271);
and U25921 (N_25921,N_22856,N_23080);
nor U25922 (N_25922,N_23320,N_22615);
and U25923 (N_25923,N_23922,N_23848);
nor U25924 (N_25924,N_23920,N_23826);
and U25925 (N_25925,N_23883,N_23487);
xor U25926 (N_25926,N_23279,N_23439);
xor U25927 (N_25927,N_22785,N_22297);
xor U25928 (N_25928,N_23192,N_22914);
or U25929 (N_25929,N_22585,N_22307);
nor U25930 (N_25930,N_23668,N_22592);
xnor U25931 (N_25931,N_22313,N_23337);
nand U25932 (N_25932,N_23598,N_23904);
and U25933 (N_25933,N_22776,N_22299);
xor U25934 (N_25934,N_22994,N_23310);
and U25935 (N_25935,N_23293,N_22313);
or U25936 (N_25936,N_22113,N_22508);
and U25937 (N_25937,N_22594,N_22476);
or U25938 (N_25938,N_23845,N_22982);
nand U25939 (N_25939,N_23593,N_22924);
nor U25940 (N_25940,N_22651,N_22112);
nor U25941 (N_25941,N_23717,N_23817);
or U25942 (N_25942,N_23892,N_23732);
nor U25943 (N_25943,N_22043,N_23588);
nor U25944 (N_25944,N_22497,N_23623);
and U25945 (N_25945,N_23345,N_22206);
nor U25946 (N_25946,N_22780,N_23872);
xnor U25947 (N_25947,N_22975,N_23512);
or U25948 (N_25948,N_22890,N_22546);
nand U25949 (N_25949,N_22006,N_22569);
and U25950 (N_25950,N_22973,N_23142);
or U25951 (N_25951,N_22231,N_22934);
xor U25952 (N_25952,N_22047,N_22297);
or U25953 (N_25953,N_22530,N_23195);
xor U25954 (N_25954,N_22467,N_23368);
nand U25955 (N_25955,N_23997,N_23526);
xor U25956 (N_25956,N_22360,N_22612);
and U25957 (N_25957,N_22932,N_23986);
and U25958 (N_25958,N_23188,N_22670);
nand U25959 (N_25959,N_22700,N_22799);
nor U25960 (N_25960,N_23360,N_22812);
and U25961 (N_25961,N_22994,N_23892);
nand U25962 (N_25962,N_22890,N_23790);
and U25963 (N_25963,N_22169,N_23111);
nand U25964 (N_25964,N_22153,N_23948);
xnor U25965 (N_25965,N_23450,N_22465);
xnor U25966 (N_25966,N_22733,N_23801);
xnor U25967 (N_25967,N_23628,N_22424);
nor U25968 (N_25968,N_23541,N_22461);
and U25969 (N_25969,N_23462,N_23777);
nor U25970 (N_25970,N_22347,N_22833);
and U25971 (N_25971,N_22870,N_23807);
or U25972 (N_25972,N_22811,N_23395);
nand U25973 (N_25973,N_22043,N_22371);
xor U25974 (N_25974,N_22397,N_23356);
xnor U25975 (N_25975,N_22834,N_22365);
nand U25976 (N_25976,N_23273,N_22813);
or U25977 (N_25977,N_22062,N_22591);
nor U25978 (N_25978,N_23252,N_23836);
or U25979 (N_25979,N_22286,N_23962);
nor U25980 (N_25980,N_22156,N_23510);
or U25981 (N_25981,N_23949,N_22595);
or U25982 (N_25982,N_22035,N_23945);
and U25983 (N_25983,N_23475,N_22281);
and U25984 (N_25984,N_23111,N_22193);
or U25985 (N_25985,N_23345,N_23625);
or U25986 (N_25986,N_22866,N_22580);
nor U25987 (N_25987,N_23094,N_22508);
or U25988 (N_25988,N_23311,N_22127);
nand U25989 (N_25989,N_23828,N_23619);
nand U25990 (N_25990,N_23898,N_23171);
nand U25991 (N_25991,N_23085,N_22471);
nor U25992 (N_25992,N_23693,N_22422);
or U25993 (N_25993,N_23174,N_23401);
nand U25994 (N_25994,N_23398,N_23132);
or U25995 (N_25995,N_23444,N_23261);
or U25996 (N_25996,N_23138,N_23921);
nand U25997 (N_25997,N_23838,N_23728);
and U25998 (N_25998,N_22561,N_22076);
or U25999 (N_25999,N_22651,N_22035);
nand U26000 (N_26000,N_25340,N_24064);
nand U26001 (N_26001,N_24238,N_25088);
or U26002 (N_26002,N_25395,N_25744);
nor U26003 (N_26003,N_24744,N_25595);
or U26004 (N_26004,N_24709,N_25157);
and U26005 (N_26005,N_24502,N_24379);
and U26006 (N_26006,N_24743,N_24694);
and U26007 (N_26007,N_24752,N_25324);
nand U26008 (N_26008,N_24407,N_25499);
xnor U26009 (N_26009,N_25934,N_24318);
xnor U26010 (N_26010,N_24184,N_25161);
nand U26011 (N_26011,N_24125,N_25545);
and U26012 (N_26012,N_24313,N_25087);
nand U26013 (N_26013,N_25315,N_24721);
xor U26014 (N_26014,N_24289,N_24567);
and U26015 (N_26015,N_24371,N_24685);
nor U26016 (N_26016,N_25299,N_25065);
nand U26017 (N_26017,N_24814,N_24011);
or U26018 (N_26018,N_24996,N_24732);
and U26019 (N_26019,N_25678,N_24299);
and U26020 (N_26020,N_25443,N_24373);
or U26021 (N_26021,N_24903,N_25307);
nor U26022 (N_26022,N_24703,N_24839);
xnor U26023 (N_26023,N_25929,N_24550);
xnor U26024 (N_26024,N_24932,N_25982);
xnor U26025 (N_26025,N_24157,N_24649);
and U26026 (N_26026,N_25612,N_24468);
nand U26027 (N_26027,N_24033,N_24673);
xnor U26028 (N_26028,N_24155,N_24335);
xor U26029 (N_26029,N_24739,N_25142);
or U26030 (N_26030,N_24599,N_25243);
nor U26031 (N_26031,N_24866,N_25713);
and U26032 (N_26032,N_24799,N_25216);
or U26033 (N_26033,N_25298,N_25444);
nand U26034 (N_26034,N_25392,N_24279);
nand U26035 (N_26035,N_25331,N_25658);
xnor U26036 (N_26036,N_24041,N_25925);
nor U26037 (N_26037,N_24728,N_24178);
nor U26038 (N_26038,N_25946,N_25091);
or U26039 (N_26039,N_25450,N_24327);
xnor U26040 (N_26040,N_25851,N_24907);
or U26041 (N_26041,N_25090,N_25190);
and U26042 (N_26042,N_25952,N_25778);
or U26043 (N_26043,N_25940,N_25950);
xnor U26044 (N_26044,N_24225,N_24232);
or U26045 (N_26045,N_24344,N_24759);
and U26046 (N_26046,N_24042,N_25777);
or U26047 (N_26047,N_25588,N_25866);
xnor U26048 (N_26048,N_25743,N_25017);
or U26049 (N_26049,N_25659,N_25417);
nand U26050 (N_26050,N_24431,N_25811);
and U26051 (N_26051,N_25664,N_25715);
xor U26052 (N_26052,N_25108,N_25148);
and U26053 (N_26053,N_24332,N_24241);
and U26054 (N_26054,N_25020,N_24603);
nand U26055 (N_26055,N_24016,N_25810);
or U26056 (N_26056,N_25211,N_24227);
and U26057 (N_26057,N_25820,N_24142);
or U26058 (N_26058,N_24760,N_25379);
xnor U26059 (N_26059,N_24828,N_24756);
or U26060 (N_26060,N_24972,N_24219);
or U26061 (N_26061,N_25366,N_25766);
and U26062 (N_26062,N_25618,N_25297);
xnor U26063 (N_26063,N_25284,N_24798);
nor U26064 (N_26064,N_25604,N_25453);
or U26065 (N_26065,N_25310,N_25923);
xor U26066 (N_26066,N_25523,N_24205);
or U26067 (N_26067,N_24944,N_24326);
or U26068 (N_26068,N_25617,N_25122);
and U26069 (N_26069,N_25046,N_24931);
xnor U26070 (N_26070,N_24590,N_24625);
or U26071 (N_26071,N_25740,N_24441);
nand U26072 (N_26072,N_25003,N_24078);
nor U26073 (N_26073,N_24872,N_24937);
and U26074 (N_26074,N_25265,N_25847);
nor U26075 (N_26075,N_24876,N_24681);
nor U26076 (N_26076,N_25974,N_25596);
and U26077 (N_26077,N_25170,N_25972);
nand U26078 (N_26078,N_25041,N_24809);
or U26079 (N_26079,N_24242,N_24408);
nand U26080 (N_26080,N_25219,N_24719);
nor U26081 (N_26081,N_24063,N_24663);
xnor U26082 (N_26082,N_25933,N_25374);
or U26083 (N_26083,N_25369,N_25285);
xor U26084 (N_26084,N_25311,N_25371);
nand U26085 (N_26085,N_24981,N_25571);
nand U26086 (N_26086,N_24447,N_25720);
xnor U26087 (N_26087,N_24234,N_24109);
or U26088 (N_26088,N_24347,N_25802);
xor U26089 (N_26089,N_25501,N_24203);
xor U26090 (N_26090,N_24493,N_25730);
or U26091 (N_26091,N_25725,N_25312);
xor U26092 (N_26092,N_24482,N_25500);
nor U26093 (N_26093,N_25408,N_24473);
or U26094 (N_26094,N_24152,N_25842);
xor U26095 (N_26095,N_25860,N_25516);
nand U26096 (N_26096,N_24708,N_25060);
xor U26097 (N_26097,N_24171,N_25416);
and U26098 (N_26098,N_25336,N_24231);
and U26099 (N_26099,N_25313,N_24588);
nand U26100 (N_26100,N_25471,N_24149);
nand U26101 (N_26101,N_24504,N_25603);
xnor U26102 (N_26102,N_24702,N_24605);
nand U26103 (N_26103,N_24212,N_25370);
or U26104 (N_26104,N_24049,N_24018);
xnor U26105 (N_26105,N_25225,N_25449);
and U26106 (N_26106,N_25788,N_25859);
nor U26107 (N_26107,N_24677,N_24137);
or U26108 (N_26108,N_25242,N_25077);
xor U26109 (N_26109,N_25152,N_25189);
nand U26110 (N_26110,N_24644,N_24767);
nand U26111 (N_26111,N_24691,N_24501);
nand U26112 (N_26112,N_25632,N_25463);
xnor U26113 (N_26113,N_24773,N_24188);
or U26114 (N_26114,N_25249,N_24396);
nand U26115 (N_26115,N_24177,N_24031);
and U26116 (N_26116,N_25023,N_25263);
and U26117 (N_26117,N_25633,N_25487);
nor U26118 (N_26118,N_25620,N_25668);
nand U26119 (N_26119,N_24880,N_24240);
or U26120 (N_26120,N_24917,N_25911);
or U26121 (N_26121,N_25044,N_25915);
xnor U26122 (N_26122,N_24869,N_24637);
or U26123 (N_26123,N_25082,N_25614);
nor U26124 (N_26124,N_25329,N_25566);
xor U26125 (N_26125,N_25159,N_24215);
or U26126 (N_26126,N_25657,N_25261);
or U26127 (N_26127,N_24411,N_24618);
nand U26128 (N_26128,N_25845,N_25586);
nor U26129 (N_26129,N_25575,N_25355);
xor U26130 (N_26130,N_24863,N_25640);
nand U26131 (N_26131,N_25132,N_25998);
and U26132 (N_26132,N_25941,N_24005);
and U26133 (N_26133,N_25838,N_25025);
nor U26134 (N_26134,N_25746,N_24782);
and U26135 (N_26135,N_24862,N_25365);
or U26136 (N_26136,N_24337,N_25931);
nor U26137 (N_26137,N_25634,N_25455);
nor U26138 (N_26138,N_25147,N_24355);
xnor U26139 (N_26139,N_25100,N_24951);
xnor U26140 (N_26140,N_25670,N_25858);
nand U26141 (N_26141,N_24631,N_25853);
nor U26142 (N_26142,N_24805,N_25994);
and U26143 (N_26143,N_25581,N_25210);
xnor U26144 (N_26144,N_25026,N_25856);
nand U26145 (N_26145,N_25102,N_25883);
xnor U26146 (N_26146,N_24827,N_25987);
nor U26147 (N_26147,N_24024,N_25172);
and U26148 (N_26148,N_24679,N_25828);
nor U26149 (N_26149,N_24896,N_24919);
or U26150 (N_26150,N_25240,N_24870);
nand U26151 (N_26151,N_24901,N_24058);
and U26152 (N_26152,N_24097,N_24518);
and U26153 (N_26153,N_24107,N_24133);
xnor U26154 (N_26154,N_25737,N_24521);
nor U26155 (N_26155,N_24988,N_24733);
nor U26156 (N_26156,N_25874,N_24400);
or U26157 (N_26157,N_24265,N_25547);
or U26158 (N_26158,N_25275,N_25949);
or U26159 (N_26159,N_24906,N_25576);
xor U26160 (N_26160,N_25729,N_24409);
or U26161 (N_26161,N_25062,N_24922);
nand U26162 (N_26162,N_24731,N_24218);
nor U26163 (N_26163,N_24338,N_25484);
nand U26164 (N_26164,N_24004,N_24170);
and U26165 (N_26165,N_25754,N_24865);
xnor U26166 (N_26166,N_25609,N_24217);
or U26167 (N_26167,N_25273,N_25409);
and U26168 (N_26168,N_24556,N_25441);
nand U26169 (N_26169,N_24079,N_24385);
nor U26170 (N_26170,N_24878,N_25610);
nor U26171 (N_26171,N_25565,N_25555);
xnor U26172 (N_26172,N_24310,N_25767);
nand U26173 (N_26173,N_24260,N_25956);
and U26174 (N_26174,N_25120,N_25178);
and U26175 (N_26175,N_24958,N_24961);
nor U26176 (N_26176,N_25019,N_24261);
xor U26177 (N_26177,N_24264,N_25623);
nand U26178 (N_26178,N_24111,N_25153);
and U26179 (N_26179,N_25817,N_25872);
nor U26180 (N_26180,N_24669,N_24384);
xor U26181 (N_26181,N_24979,N_24623);
nand U26182 (N_26182,N_24390,N_24082);
or U26183 (N_26183,N_25004,N_25474);
xnor U26184 (N_26184,N_24275,N_24948);
and U26185 (N_26185,N_25676,N_24019);
and U26186 (N_26186,N_25671,N_25378);
nand U26187 (N_26187,N_24822,N_24969);
xor U26188 (N_26188,N_25745,N_25990);
nor U26189 (N_26189,N_24689,N_25421);
nand U26190 (N_26190,N_24941,N_24817);
or U26191 (N_26191,N_25958,N_24140);
or U26192 (N_26192,N_24580,N_24300);
nor U26193 (N_26193,N_24734,N_24965);
xnor U26194 (N_26194,N_24553,N_24168);
and U26195 (N_26195,N_25930,N_24766);
and U26196 (N_26196,N_25826,N_24340);
xor U26197 (N_26197,N_25112,N_25070);
and U26198 (N_26198,N_24528,N_25738);
nor U26199 (N_26199,N_24353,N_25475);
xor U26200 (N_26200,N_24076,N_24268);
nor U26201 (N_26201,N_24304,N_25661);
or U26202 (N_26202,N_25698,N_25599);
and U26203 (N_26203,N_25751,N_25427);
xor U26204 (N_26204,N_24596,N_24469);
nand U26205 (N_26205,N_24987,N_24593);
or U26206 (N_26206,N_24592,N_25058);
xor U26207 (N_26207,N_24443,N_25871);
or U26208 (N_26208,N_25177,N_25741);
nor U26209 (N_26209,N_24266,N_24173);
nand U26210 (N_26210,N_24035,N_24290);
or U26211 (N_26211,N_25359,N_25906);
xor U26212 (N_26212,N_25413,N_25585);
nand U26213 (N_26213,N_24710,N_25419);
nor U26214 (N_26214,N_24239,N_24027);
nor U26215 (N_26215,N_24933,N_24388);
and U26216 (N_26216,N_24888,N_24722);
and U26217 (N_26217,N_25945,N_24280);
nor U26218 (N_26218,N_24800,N_25008);
nand U26219 (N_26219,N_24450,N_25106);
xnor U26220 (N_26220,N_24640,N_25005);
nor U26221 (N_26221,N_25393,N_24886);
or U26222 (N_26222,N_24601,N_24455);
nor U26223 (N_26223,N_25719,N_25038);
or U26224 (N_26224,N_24973,N_25049);
nor U26225 (N_26225,N_24635,N_25823);
xor U26226 (N_26226,N_24258,N_25259);
xor U26227 (N_26227,N_24651,N_25289);
or U26228 (N_26228,N_25418,N_24475);
nor U26229 (N_26229,N_24253,N_25056);
or U26230 (N_26230,N_25390,N_24398);
xor U26231 (N_26231,N_24538,N_24096);
or U26232 (N_26232,N_24466,N_25988);
nor U26233 (N_26233,N_24477,N_25051);
nor U26234 (N_26234,N_24272,N_25677);
and U26235 (N_26235,N_24202,N_25066);
nand U26236 (N_26236,N_25101,N_24984);
nor U26237 (N_26237,N_24083,N_25232);
and U26238 (N_26238,N_24119,N_25063);
xnor U26239 (N_26239,N_24189,N_25895);
nand U26240 (N_26240,N_25696,N_25939);
or U26241 (N_26241,N_24707,N_25030);
and U26242 (N_26242,N_25384,N_25466);
xor U26243 (N_26243,N_24439,N_24874);
nor U26244 (N_26244,N_24832,N_24423);
nand U26245 (N_26245,N_25126,N_24855);
nand U26246 (N_26246,N_25513,N_25721);
or U26247 (N_26247,N_24252,N_24758);
xnor U26248 (N_26248,N_25837,N_24853);
nor U26249 (N_26249,N_25793,N_24309);
and U26250 (N_26250,N_24693,N_25804);
and U26251 (N_26251,N_25482,N_24893);
nor U26252 (N_26252,N_24167,N_25451);
xor U26253 (N_26253,N_24717,N_24174);
nand U26254 (N_26254,N_24500,N_25795);
nor U26255 (N_26255,N_24882,N_24437);
or U26256 (N_26256,N_25966,N_24002);
nor U26257 (N_26257,N_25024,N_24613);
nand U26258 (N_26258,N_24416,N_24511);
xnor U26259 (N_26259,N_25167,N_24522);
xor U26260 (N_26260,N_25918,N_25229);
nand U26261 (N_26261,N_25353,N_24871);
nand U26262 (N_26262,N_25684,N_25625);
xnor U26263 (N_26263,N_24576,N_25013);
nand U26264 (N_26264,N_25339,N_24611);
nand U26265 (N_26265,N_25697,N_24881);
and U26266 (N_26266,N_24051,N_24285);
or U26267 (N_26267,N_25753,N_25690);
nand U26268 (N_26268,N_24496,N_24532);
and U26269 (N_26269,N_24793,N_24248);
xor U26270 (N_26270,N_25563,N_24319);
or U26271 (N_26271,N_24386,N_25727);
and U26272 (N_26272,N_24432,N_24141);
nor U26273 (N_26273,N_24414,N_24746);
xnor U26274 (N_26274,N_24768,N_25173);
and U26275 (N_26275,N_25262,N_24790);
xor U26276 (N_26276,N_25878,N_25053);
xor U26277 (N_26277,N_25402,N_24478);
and U26278 (N_26278,N_24505,N_24271);
nand U26279 (N_26279,N_24824,N_25174);
xor U26280 (N_26280,N_25747,N_24276);
and U26281 (N_26281,N_25989,N_24247);
xnor U26282 (N_26282,N_24487,N_25672);
or U26283 (N_26283,N_24970,N_25061);
xnor U26284 (N_26284,N_25735,N_25924);
nand U26285 (N_26285,N_25042,N_24867);
nor U26286 (N_26286,N_25459,N_24484);
nand U26287 (N_26287,N_24176,N_24544);
nand U26288 (N_26288,N_25276,N_24283);
xnor U26289 (N_26289,N_24349,N_24040);
nand U26290 (N_26290,N_25202,N_24753);
and U26291 (N_26291,N_25888,N_24124);
or U26292 (N_26292,N_24868,N_25636);
or U26293 (N_26293,N_25538,N_24991);
nor U26294 (N_26294,N_25704,N_24006);
or U26295 (N_26295,N_24415,N_25430);
or U26296 (N_26296,N_25032,N_24840);
and U26297 (N_26297,N_24525,N_25304);
xor U26298 (N_26298,N_25607,N_24410);
or U26299 (N_26299,N_25695,N_25015);
or U26300 (N_26300,N_24950,N_25234);
nor U26301 (N_26301,N_25176,N_25398);
and U26302 (N_26302,N_25196,N_24401);
nor U26303 (N_26303,N_25350,N_25722);
and U26304 (N_26304,N_25305,N_25927);
and U26305 (N_26305,N_24350,N_25997);
nor U26306 (N_26306,N_24092,N_25809);
or U26307 (N_26307,N_24181,N_25151);
xnor U26308 (N_26308,N_24724,N_24150);
nor U26309 (N_26309,N_24315,N_25054);
or U26310 (N_26310,N_25943,N_24454);
or U26311 (N_26311,N_24130,N_25981);
nand U26312 (N_26312,N_24998,N_24134);
xnor U26313 (N_26313,N_24974,N_24449);
and U26314 (N_26314,N_25750,N_25278);
and U26315 (N_26315,N_24297,N_24552);
or U26316 (N_26316,N_24053,N_24578);
nand U26317 (N_26317,N_25528,N_25277);
nor U26318 (N_26318,N_25639,N_25321);
nor U26319 (N_26319,N_24296,N_25770);
and U26320 (N_26320,N_24164,N_25028);
and U26321 (N_26321,N_25055,N_25509);
and U26322 (N_26322,N_25573,N_25682);
nand U26323 (N_26323,N_24320,N_25389);
nand U26324 (N_26324,N_24186,N_25097);
nand U26325 (N_26325,N_25957,N_24526);
or U26326 (N_26326,N_25591,N_24467);
and U26327 (N_26327,N_25960,N_24259);
nor U26328 (N_26328,N_25037,N_25251);
or U26329 (N_26329,N_25436,N_25119);
nor U26330 (N_26330,N_24755,N_24025);
and U26331 (N_26331,N_25212,N_25819);
nor U26332 (N_26332,N_24928,N_24975);
or U26333 (N_26333,N_25540,N_24897);
xor U26334 (N_26334,N_25805,N_25470);
nand U26335 (N_26335,N_24531,N_24529);
xnor U26336 (N_26336,N_24547,N_25602);
nand U26337 (N_26337,N_25977,N_25085);
and U26338 (N_26338,N_25412,N_24671);
and U26339 (N_26339,N_24668,N_24001);
nor U26340 (N_26340,N_24233,N_24488);
nor U26341 (N_26341,N_24055,N_25011);
and U26342 (N_26342,N_24780,N_24038);
or U26343 (N_26343,N_25363,N_24541);
nand U26344 (N_26344,N_25855,N_24844);
nand U26345 (N_26345,N_25154,N_24345);
and U26346 (N_26346,N_25396,N_24406);
or U26347 (N_26347,N_24343,N_25193);
and U26348 (N_26348,N_24960,N_24581);
nand U26349 (N_26349,N_25308,N_24116);
xnor U26350 (N_26350,N_25424,N_25524);
xnor U26351 (N_26351,N_25179,N_25440);
and U26352 (N_26352,N_25282,N_24847);
nor U26353 (N_26353,N_25635,N_25897);
or U26354 (N_26354,N_24524,N_24517);
and U26355 (N_26355,N_25083,N_24391);
nand U26356 (N_26356,N_24682,N_24235);
xnor U26357 (N_26357,N_24192,N_24678);
and U26358 (N_26358,N_24495,N_25283);
nor U26359 (N_26359,N_25884,N_24357);
xnor U26360 (N_26360,N_24628,N_25246);
and U26361 (N_26361,N_25961,N_24595);
xor U26362 (N_26362,N_24543,N_25787);
or U26363 (N_26363,N_24270,N_25048);
and U26364 (N_26364,N_25293,N_24044);
nor U26365 (N_26365,N_24052,N_25118);
nand U26366 (N_26366,N_25605,N_24894);
and U26367 (N_26367,N_24204,N_25169);
xnor U26368 (N_26368,N_24220,N_24510);
and U26369 (N_26369,N_24925,N_25869);
and U26370 (N_26370,N_24818,N_25587);
xnor U26371 (N_26371,N_25456,N_24359);
nor U26372 (N_26372,N_25533,N_25292);
xnor U26373 (N_26373,N_25504,N_25944);
and U26374 (N_26374,N_25345,N_25914);
and U26375 (N_26375,N_25185,N_24062);
or U26376 (N_26376,N_25868,N_24546);
nand U26377 (N_26377,N_24751,N_25964);
xnor U26378 (N_26378,N_25759,N_24774);
xnor U26379 (N_26379,N_25515,N_24311);
nor U26380 (N_26380,N_25792,N_25707);
nor U26381 (N_26381,N_25397,N_25881);
nand U26382 (N_26382,N_25731,N_25899);
and U26383 (N_26383,N_25846,N_24598);
and U26384 (N_26384,N_25437,N_25537);
nor U26385 (N_26385,N_24479,N_24395);
and U26386 (N_26386,N_25546,N_25665);
nor U26387 (N_26387,N_25386,N_25291);
nor U26388 (N_26388,N_24537,N_25006);
and U26389 (N_26389,N_25887,N_24440);
and U26390 (N_26390,N_25644,N_25709);
nor U26391 (N_26391,N_24688,N_24069);
and U26392 (N_26392,N_24132,N_25579);
xnor U26393 (N_26393,N_24936,N_25903);
nand U26394 (N_26394,N_24690,N_24383);
or U26395 (N_26395,N_24336,N_24489);
and U26396 (N_26396,N_24514,N_24738);
nor U26397 (N_26397,N_24093,N_24539);
or U26398 (N_26398,N_24619,N_25733);
or U26399 (N_26399,N_25479,N_24796);
or U26400 (N_26400,N_25830,N_24230);
xor U26401 (N_26401,N_25919,N_25163);
xnor U26402 (N_26402,N_25520,N_24328);
nor U26403 (N_26403,N_25687,N_25047);
nor U26404 (N_26404,N_24426,N_24995);
xor U26405 (N_26405,N_24348,N_25531);
nand U26406 (N_26406,N_25227,N_25016);
and U26407 (N_26407,N_25476,N_24675);
xor U26408 (N_26408,N_24711,N_25765);
nor U26409 (N_26409,N_25824,N_25226);
or U26410 (N_26410,N_24013,N_24159);
xor U26411 (N_26411,N_25932,N_24540);
or U26412 (N_26412,N_25836,N_24175);
or U26413 (N_26413,N_25410,N_24959);
or U26414 (N_26414,N_25175,N_24913);
xnor U26415 (N_26415,N_24575,N_24803);
or U26416 (N_26416,N_25626,N_25271);
nand U26417 (N_26417,N_24399,N_25592);
xor U26418 (N_26418,N_25200,N_25896);
or U26419 (N_26419,N_24389,N_24968);
nand U26420 (N_26420,N_25983,N_24962);
xor U26421 (N_26421,N_24008,N_25156);
xor U26422 (N_26422,N_24577,N_25146);
xor U26423 (N_26423,N_24108,N_25429);
and U26424 (N_26424,N_25786,N_25995);
nor U26425 (N_26425,N_24191,N_24615);
xnor U26426 (N_26426,N_24148,N_25322);
and U26427 (N_26427,N_25627,N_24939);
nor U26428 (N_26428,N_25667,N_25512);
xnor U26429 (N_26429,N_24307,N_24037);
xnor U26430 (N_26430,N_25904,N_25748);
or U26431 (N_26431,N_24620,N_25926);
and U26432 (N_26432,N_25236,N_25567);
nand U26433 (N_26433,N_25680,N_24655);
nor U26434 (N_26434,N_24366,N_24459);
xor U26435 (N_26435,N_24207,N_25848);
and U26436 (N_26436,N_24823,N_25040);
nand U26437 (N_26437,N_24295,N_24249);
xnor U26438 (N_26438,N_25420,N_25223);
xnor U26439 (N_26439,N_24161,N_24956);
xnor U26440 (N_26440,N_25752,N_24445);
and U26441 (N_26441,N_24308,N_24007);
and U26442 (N_26442,N_24000,N_24610);
xor U26443 (N_26443,N_25075,N_24834);
nand U26444 (N_26444,N_24471,N_25300);
nand U26445 (N_26445,N_24117,N_25235);
xor U26446 (N_26446,N_24193,N_25529);
and U26447 (N_26447,N_24302,N_25757);
or U26448 (N_26448,N_24520,N_24314);
nor U26449 (N_26449,N_25320,N_25844);
nand U26450 (N_26450,N_25947,N_25191);
nand U26451 (N_26451,N_25959,N_25254);
nand U26452 (N_26452,N_24564,N_24138);
nand U26453 (N_26453,N_25464,N_25985);
or U26454 (N_26454,N_25404,N_25433);
nor U26455 (N_26455,N_25666,N_25431);
nand U26456 (N_26456,N_25825,N_25485);
xor U26457 (N_26457,N_24883,N_24617);
nand U26458 (N_26458,N_25314,N_25428);
and U26459 (N_26459,N_25139,N_25045);
or U26460 (N_26460,N_24555,N_25594);
and U26461 (N_26461,N_25922,N_25873);
xnor U26462 (N_26462,N_24372,N_25507);
xnor U26463 (N_26463,N_25773,N_24705);
or U26464 (N_26464,N_25891,N_25203);
nand U26465 (N_26465,N_24094,N_25822);
nor U26466 (N_26466,N_25968,N_24830);
nor U26467 (N_26467,N_24201,N_24807);
xnor U26468 (N_26468,N_25699,N_25550);
or U26469 (N_26469,N_25833,N_25791);
nand U26470 (N_26470,N_25086,N_25078);
nand U26471 (N_26471,N_25768,N_25646);
or U26472 (N_26472,N_25549,N_24068);
or U26473 (N_26473,N_25674,N_25882);
nand U26474 (N_26474,N_24930,N_24370);
xnor U26475 (N_26475,N_25728,N_25807);
or U26476 (N_26476,N_24813,N_24209);
nor U26477 (N_26477,N_25036,N_25508);
and U26478 (N_26478,N_24010,N_24503);
and U26479 (N_26479,N_24404,N_24562);
nand U26480 (N_26480,N_25840,N_25580);
nand U26481 (N_26481,N_25917,N_25708);
xnor U26482 (N_26482,N_25149,N_25162);
nand U26483 (N_26483,N_25208,N_24638);
and U26484 (N_26484,N_25701,N_24513);
and U26485 (N_26485,N_25525,N_25486);
or U26486 (N_26486,N_24387,N_24490);
nor U26487 (N_26487,N_25562,N_24061);
or U26488 (N_26488,N_25886,N_24533);
nor U26489 (N_26489,N_25279,N_25905);
and U26490 (N_26490,N_24147,N_25813);
and U26491 (N_26491,N_25467,N_25361);
or U26492 (N_26492,N_25776,N_24452);
or U26493 (N_26493,N_24953,N_24067);
nor U26494 (N_26494,N_25774,N_24735);
and U26495 (N_26495,N_24726,N_24321);
xor U26496 (N_26496,N_25237,N_25517);
and U26497 (N_26497,N_25539,N_24569);
nand U26498 (N_26498,N_24185,N_24160);
xor U26499 (N_26499,N_24187,N_24566);
nor U26500 (N_26500,N_24034,N_24425);
nand U26501 (N_26501,N_24136,N_25724);
xor U26502 (N_26502,N_24460,N_25438);
nor U26503 (N_26503,N_24403,N_25734);
xnor U26504 (N_26504,N_25492,N_24015);
or U26505 (N_26505,N_25095,N_25221);
nand U26506 (N_26506,N_25286,N_24073);
nand U26507 (N_26507,N_25104,N_25326);
or U26508 (N_26508,N_24563,N_24574);
xnor U26509 (N_26509,N_24551,N_24129);
xor U26510 (N_26510,N_25043,N_24485);
nand U26511 (N_26511,N_24875,N_25192);
nor U26512 (N_26512,N_25717,N_24394);
and U26513 (N_26513,N_25970,N_25955);
nor U26514 (N_26514,N_24761,N_24523);
or U26515 (N_26515,N_25681,N_25255);
or U26516 (N_26516,N_25526,N_25877);
and U26517 (N_26517,N_25080,N_25407);
or U26518 (N_26518,N_24199,N_25800);
and U26519 (N_26519,N_25018,N_25534);
or U26520 (N_26520,N_25783,N_25600);
xor U26521 (N_26521,N_25511,N_25779);
nand U26522 (N_26522,N_24256,N_25207);
and U26523 (N_26523,N_25478,N_25852);
nand U26524 (N_26524,N_24778,N_25264);
and U26525 (N_26525,N_25799,N_24812);
nand U26526 (N_26526,N_24582,N_25522);
and U26527 (N_26527,N_25818,N_24997);
xnor U26528 (N_26528,N_24572,N_25651);
xnor U26529 (N_26529,N_25506,N_25756);
or U26530 (N_26530,N_24022,N_25606);
nor U26531 (N_26531,N_24647,N_25991);
nand U26532 (N_26532,N_24197,N_24085);
nand U26533 (N_26533,N_25383,N_24648);
nand U26534 (N_26534,N_24317,N_24480);
xnor U26535 (N_26535,N_25483,N_24105);
and U26536 (N_26536,N_24943,N_24747);
nor U26537 (N_26537,N_24650,N_24071);
or U26538 (N_26538,N_24811,N_25892);
or U26539 (N_26539,N_25510,N_24325);
or U26540 (N_26540,N_25447,N_24499);
xnor U26541 (N_26541,N_24986,N_24208);
nor U26542 (N_26542,N_25902,N_24392);
xor U26543 (N_26543,N_25401,N_24559);
nand U26544 (N_26544,N_25205,N_25434);
xor U26545 (N_26545,N_25260,N_25505);
and U26546 (N_26546,N_25803,N_25241);
nand U26547 (N_26547,N_24128,N_24286);
or U26548 (N_26548,N_24312,N_24806);
nor U26549 (N_26549,N_25953,N_24095);
nor U26550 (N_26550,N_25494,N_25875);
nor U26551 (N_26551,N_24065,N_25295);
xor U26552 (N_26552,N_25488,N_24993);
and U26553 (N_26553,N_24213,N_24424);
and U26554 (N_26554,N_24420,N_25993);
nor U26555 (N_26555,N_24632,N_25349);
nor U26556 (N_26556,N_24393,N_25541);
nor U26557 (N_26557,N_25107,N_24785);
or U26558 (N_26558,N_24664,N_25685);
nor U26559 (N_26559,N_25736,N_24236);
nor U26560 (N_26560,N_24463,N_24451);
xor U26561 (N_26561,N_24099,N_25071);
xnor U26562 (N_26562,N_24419,N_24633);
or U26563 (N_26563,N_25689,N_25328);
xnor U26564 (N_26564,N_25710,N_24534);
xnor U26565 (N_26565,N_24946,N_25098);
nor U26566 (N_26566,N_25198,N_25472);
nor U26567 (N_26567,N_25999,N_24697);
nor U26568 (N_26568,N_25780,N_24154);
nand U26569 (N_26569,N_25360,N_24643);
xor U26570 (N_26570,N_25131,N_24624);
xnor U26571 (N_26571,N_24594,N_25835);
nand U26572 (N_26572,N_24354,N_25281);
nor U26573 (N_26573,N_24560,N_25423);
xnor U26574 (N_26574,N_24736,N_24433);
nand U26575 (N_26575,N_24331,N_24926);
nand U26576 (N_26576,N_24900,N_24123);
nand U26577 (N_26577,N_24103,N_24737);
or U26578 (N_26578,N_24548,N_25910);
xor U26579 (N_26579,N_25568,N_24453);
nor U26580 (N_26580,N_24683,N_24627);
nand U26581 (N_26581,N_25165,N_25052);
nand U26582 (N_26582,N_25554,N_24196);
and U26583 (N_26583,N_25951,N_25411);
or U26584 (N_26584,N_24497,N_25937);
nor U26585 (N_26585,N_24026,N_24706);
or U26586 (N_26586,N_25790,N_25213);
or U26587 (N_26587,N_25302,N_24229);
or U26588 (N_26588,N_24742,N_24836);
nor U26589 (N_26589,N_25624,N_24602);
nor U26590 (N_26590,N_25663,N_24162);
nor U26591 (N_26591,N_24291,N_25439);
nor U26592 (N_26592,N_25309,N_25782);
and U26593 (N_26593,N_25867,N_25031);
and U26594 (N_26594,N_25014,N_24542);
xor U26595 (N_26595,N_24330,N_25448);
nand U26596 (N_26596,N_25916,N_25976);
and U26597 (N_26597,N_24763,N_25405);
or U26598 (N_26598,N_24934,N_25590);
nand U26599 (N_26599,N_24293,N_25399);
or U26600 (N_26600,N_24879,N_24519);
nor U26601 (N_26601,N_25978,N_25168);
nor U26602 (N_26602,N_24145,N_25021);
or U26603 (N_26603,N_25469,N_25356);
xnor U26604 (N_26604,N_24228,N_25280);
or U26605 (N_26605,N_24088,N_24849);
or U26606 (N_26606,N_25150,N_24850);
xor U26607 (N_26607,N_24910,N_24156);
xor U26608 (N_26608,N_25621,N_25364);
xnor U26609 (N_26609,N_25303,N_25619);
xnor U26610 (N_26610,N_25099,N_25973);
nand U26611 (N_26611,N_24687,N_25258);
xor U26612 (N_26612,N_25067,N_25815);
and U26613 (N_26613,N_24114,N_25876);
nor U26614 (N_26614,N_25114,N_24029);
or U26615 (N_26615,N_25693,N_25201);
xnor U26616 (N_26616,N_25834,N_24070);
or U26617 (N_26617,N_25771,N_25454);
xnor U26618 (N_26618,N_25022,N_25141);
or U26619 (N_26619,N_24023,N_25079);
nor U26620 (N_26620,N_25332,N_25343);
xnor U26621 (N_26621,N_24754,N_24587);
and U26622 (N_26622,N_25908,N_24368);
and U26623 (N_26623,N_24586,N_24438);
or U26624 (N_26624,N_24195,N_24741);
nand U26625 (N_26625,N_25266,N_25457);
nand U26626 (N_26626,N_24179,N_25652);
nand U26627 (N_26627,N_25111,N_24859);
and U26628 (N_26628,N_25763,N_24444);
nor U26629 (N_26629,N_24351,N_24804);
and U26630 (N_26630,N_24791,N_25480);
xnor U26631 (N_26631,N_25481,N_25007);
nand U26632 (N_26632,N_24665,N_25244);
nor U26633 (N_26633,N_25465,N_25376);
xnor U26634 (N_26634,N_24654,N_24557);
nand U26635 (N_26635,N_25253,N_24750);
nand U26636 (N_26636,N_25702,N_25781);
and U26637 (N_26637,N_25986,N_24957);
nand U26638 (N_26638,N_24971,N_25900);
or U26639 (N_26639,N_25116,N_24629);
or U26640 (N_26640,N_24151,N_25084);
nor U26641 (N_26641,N_24591,N_24783);
nor U26642 (N_26642,N_25553,N_25337);
and U26643 (N_26643,N_25643,N_24924);
xor U26644 (N_26644,N_24481,N_24104);
xor U26645 (N_26645,N_24110,N_25327);
or U26646 (N_26646,N_25921,N_25814);
nor U26647 (N_26647,N_24686,N_24074);
or U26648 (N_26648,N_24512,N_24716);
nor U26649 (N_26649,N_25718,N_24210);
or U26650 (N_26650,N_24621,N_25789);
xnor U26651 (N_26651,N_24269,N_25849);
or U26652 (N_26652,N_24911,N_24530);
or U26653 (N_26653,N_25195,N_24045);
xnor U26654 (N_26654,N_25556,N_25181);
nand U26655 (N_26655,N_24054,N_24698);
nand U26656 (N_26656,N_24367,N_25843);
xor U26657 (N_26657,N_25352,N_25629);
xor U26658 (N_26658,N_25027,N_24825);
nand U26659 (N_26659,N_24947,N_24606);
nand U26660 (N_26660,N_25033,N_24856);
nor U26661 (N_26661,N_24153,N_24891);
nand U26662 (N_26662,N_24908,N_25854);
and U26663 (N_26663,N_25103,N_24277);
xor U26664 (N_26664,N_24106,N_24039);
nand U26665 (N_26665,N_25446,N_25552);
and U26666 (N_26666,N_24967,N_25649);
nor U26667 (N_26667,N_25073,N_25560);
and U26668 (N_26668,N_25761,N_24826);
nor U26669 (N_26669,N_24089,N_24720);
or U26670 (N_26670,N_25589,N_25250);
nand U26671 (N_26671,N_24714,N_25319);
nand U26672 (N_26672,N_24486,N_25094);
nand U26673 (N_26673,N_24674,N_25130);
or U26674 (N_26674,N_24604,N_25110);
xnor U26675 (N_26675,N_25323,N_25732);
or U26676 (N_26676,N_24057,N_25452);
nand U26677 (N_26677,N_25980,N_24226);
nand U26678 (N_26678,N_24221,N_24776);
or U26679 (N_26679,N_24434,N_25035);
and U26680 (N_26680,N_25214,N_25140);
or U26681 (N_26681,N_25920,N_24749);
or U26682 (N_26682,N_25683,N_25551);
xnor U26683 (N_26683,N_25010,N_24561);
xor U26684 (N_26684,N_24841,N_25391);
nand U26685 (N_26685,N_24009,N_24056);
and U26686 (N_26686,N_24614,N_24216);
or U26687 (N_26687,N_25694,N_25572);
nor U26688 (N_26688,N_24342,N_25880);
nand U26689 (N_26689,N_25109,N_24642);
nand U26690 (N_26690,N_24172,N_24098);
xnor U26691 (N_26691,N_24912,N_24346);
and U26692 (N_26692,N_24458,N_25654);
or U26693 (N_26693,N_24166,N_24781);
nor U26694 (N_26694,N_24245,N_24237);
and U26695 (N_26695,N_25582,N_25233);
or U26696 (N_26696,N_24589,N_24554);
xnor U26697 (N_26697,N_25829,N_25962);
and U26698 (N_26698,N_24784,N_24402);
and U26699 (N_26699,N_24244,N_24352);
nor U26700 (N_26700,N_24333,N_24169);
or U26701 (N_26701,N_25544,N_24456);
or U26702 (N_26702,N_24360,N_24935);
nor U26703 (N_26703,N_24413,N_24718);
and U26704 (N_26704,N_25377,N_24964);
and U26705 (N_26705,N_24890,N_24457);
or U26706 (N_26706,N_25388,N_24570);
and U26707 (N_26707,N_24659,N_24977);
and U26708 (N_26708,N_25769,N_25984);
nor U26709 (N_26709,N_25217,N_25971);
nor U26710 (N_26710,N_25269,N_25495);
nor U26711 (N_26711,N_25821,N_25267);
or U26712 (N_26712,N_24498,N_25317);
or U26713 (N_26713,N_24422,N_25561);
nand U26714 (N_26714,N_24080,N_24701);
or U26715 (N_26715,N_24243,N_25493);
nand U26716 (N_26716,N_24483,N_24989);
nand U26717 (N_26717,N_25532,N_25188);
nor U26718 (N_26718,N_25268,N_24448);
xnor U26719 (N_26719,N_25850,N_25182);
nor U26720 (N_26720,N_25498,N_24797);
nand U26721 (N_26721,N_25296,N_24081);
and U26722 (N_26722,N_25338,N_25415);
or U26723 (N_26723,N_24808,N_25368);
or U26724 (N_26724,N_25372,N_25992);
nand U26725 (N_26725,N_24845,N_24833);
nand U26726 (N_26726,N_24012,N_24375);
xor U26727 (N_26727,N_24047,N_25394);
nor U26728 (N_26728,N_24322,N_24163);
xnor U26729 (N_26729,N_24945,N_24075);
and U26730 (N_26730,N_25442,N_25583);
or U26731 (N_26731,N_25215,N_25714);
and U26732 (N_26732,N_25965,N_24667);
or U26733 (N_26733,N_25655,N_25622);
or U26734 (N_26734,N_25301,N_24978);
xnor U26735 (N_26735,N_25863,N_24608);
xnor U26736 (N_26736,N_24585,N_25224);
nand U26737 (N_26737,N_24666,N_25468);
nor U26738 (N_26738,N_24374,N_24418);
nand U26739 (N_26739,N_24729,N_24086);
xor U26740 (N_26740,N_24397,N_24646);
nor U26741 (N_26741,N_24113,N_25584);
and U26742 (N_26742,N_25115,N_24298);
or U26743 (N_26743,N_24316,N_25133);
nor U26744 (N_26744,N_24568,N_24662);
nand U26745 (N_26745,N_25601,N_25385);
and U26746 (N_26746,N_24476,N_25290);
nand U26747 (N_26747,N_25462,N_25230);
xnor U26748 (N_26748,N_24101,N_24288);
nor U26749 (N_26749,N_25831,N_25631);
or U26750 (N_26750,N_25686,N_24474);
or U26751 (N_26751,N_24622,N_24036);
or U26752 (N_26752,N_25491,N_25723);
xor U26753 (N_26753,N_25460,N_25209);
nand U26754 (N_26754,N_24748,N_24257);
nand U26755 (N_26755,N_25535,N_24772);
nand U26756 (N_26756,N_25245,N_25197);
xnor U26757 (N_26757,N_24942,N_24898);
nor U26758 (N_26758,N_25064,N_24158);
nand U26759 (N_26759,N_25912,N_24306);
or U26760 (N_26760,N_25473,N_25865);
or U26761 (N_26761,N_24764,N_25775);
and U26762 (N_26762,N_25403,N_24672);
and U26763 (N_26763,N_25117,N_24334);
and U26764 (N_26764,N_25124,N_25890);
nor U26765 (N_26765,N_25975,N_24380);
xnor U26766 (N_26766,N_24725,N_25967);
and U26767 (N_26767,N_25716,N_25375);
or U26768 (N_26768,N_24043,N_24442);
nand U26769 (N_26769,N_24194,N_24369);
xnor U26770 (N_26770,N_25613,N_24884);
xnor U26771 (N_26771,N_24940,N_24364);
nor U26772 (N_26772,N_25218,N_24515);
xor U26773 (N_26773,N_24378,N_24508);
or U26774 (N_26774,N_25490,N_24821);
nor U26775 (N_26775,N_25333,N_25406);
or U26776 (N_26776,N_25785,N_24829);
and U26777 (N_26777,N_24362,N_25705);
nor U26778 (N_26778,N_25797,N_24182);
or U26779 (N_26779,N_24436,N_24634);
and U26780 (N_26780,N_25432,N_25954);
nor U26781 (N_26781,N_24506,N_25496);
and U26782 (N_26782,N_24222,N_25318);
or U26783 (N_26783,N_24641,N_25256);
and U26784 (N_26784,N_25186,N_25942);
and U26785 (N_26785,N_25628,N_25839);
nand U26786 (N_26786,N_24949,N_24028);
and U26787 (N_26787,N_24661,N_25164);
nor U26788 (N_26788,N_24857,N_25382);
nor U26789 (N_26789,N_24695,N_25206);
xnor U26790 (N_26790,N_24014,N_24920);
nor U26791 (N_26791,N_25400,N_24771);
and U26792 (N_26792,N_24143,N_24904);
nand U26793 (N_26793,N_24381,N_25057);
xor U26794 (N_26794,N_25105,N_24607);
nand U26795 (N_26795,N_25204,N_24121);
xor U26796 (N_26796,N_24255,N_25089);
or U26797 (N_26797,N_25616,N_25816);
xor U26798 (N_26798,N_24223,N_24571);
nand U26799 (N_26799,N_25641,N_24630);
and U26800 (N_26800,N_25578,N_25334);
or U26801 (N_26801,N_25808,N_25519);
nor U26802 (N_26802,N_24146,N_24966);
and U26803 (N_26803,N_24060,N_25238);
and U26804 (N_26804,N_24819,N_24990);
or U26805 (N_26805,N_24902,N_25138);
xnor U26806 (N_26806,N_24918,N_24787);
and U26807 (N_26807,N_24626,N_24837);
and U26808 (N_26808,N_24281,N_24100);
and U26809 (N_26809,N_24639,N_25125);
nor U26810 (N_26810,N_24684,N_25166);
and U26811 (N_26811,N_25559,N_25726);
and U26812 (N_26812,N_24777,N_24816);
and U26813 (N_26813,N_24183,N_25199);
xnor U26814 (N_26814,N_25074,N_24852);
nand U26815 (N_26815,N_25611,N_24795);
nand U26816 (N_26816,N_24430,N_24858);
and U26817 (N_26817,N_24535,N_25367);
xor U26818 (N_26818,N_25001,N_25489);
nand U26819 (N_26819,N_25907,N_25673);
nor U26820 (N_26820,N_25794,N_24769);
nor U26821 (N_26821,N_24429,N_25527);
or U26822 (N_26822,N_25096,N_24696);
and U26823 (N_26823,N_25669,N_25344);
xnor U26824 (N_26824,N_24600,N_24909);
nand U26825 (N_26825,N_24802,N_25593);
and U26826 (N_26826,N_25287,N_25059);
and U26827 (N_26827,N_24017,N_25143);
and U26828 (N_26828,N_24066,N_25093);
and U26829 (N_26829,N_24810,N_25445);
nor U26830 (N_26830,N_25885,N_24303);
and U26831 (N_26831,N_24657,N_25348);
and U26832 (N_26832,N_25969,N_24020);
nor U26833 (N_26833,N_24435,N_25739);
and U26834 (N_26834,N_25231,N_24274);
or U26835 (N_26835,N_24670,N_25502);
nor U26836 (N_26836,N_25180,N_24021);
nor U26837 (N_26837,N_24365,N_24120);
nor U26838 (N_26838,N_25288,N_25712);
xor U26839 (N_26839,N_24091,N_24745);
and U26840 (N_26840,N_25137,N_25187);
nand U26841 (N_26841,N_25145,N_24770);
xnor U26842 (N_26842,N_25514,N_24127);
or U26843 (N_26843,N_25893,N_24786);
nand U26844 (N_26844,N_25039,N_25012);
and U26845 (N_26845,N_25688,N_24994);
and U26846 (N_26846,N_24549,N_24102);
nor U26847 (N_26847,N_24843,N_25270);
or U26848 (N_26848,N_25144,N_25557);
or U26849 (N_26849,N_24835,N_24992);
nand U26850 (N_26850,N_24860,N_24363);
nor U26851 (N_26851,N_24788,N_25798);
xnor U26852 (N_26852,N_24329,N_24916);
xor U26853 (N_26853,N_25711,N_24428);
nand U26854 (N_26854,N_24122,N_24609);
or U26855 (N_26855,N_25679,N_25862);
nand U26856 (N_26856,N_24112,N_25762);
and U26857 (N_26857,N_24851,N_25362);
or U26858 (N_26858,N_24877,N_24704);
or U26859 (N_26859,N_24294,N_25183);
nor U26860 (N_26860,N_25948,N_25136);
or U26861 (N_26861,N_24775,N_25650);
or U26862 (N_26862,N_24254,N_24224);
nor U26863 (N_26863,N_25239,N_24135);
xor U26864 (N_26864,N_25700,N_24077);
and U26865 (N_26865,N_24757,N_24692);
and U26866 (N_26866,N_25127,N_24072);
and U26867 (N_26867,N_25220,N_25426);
or U26868 (N_26868,N_24376,N_25784);
nor U26869 (N_26869,N_25435,N_25648);
nor U26870 (N_26870,N_24358,N_25380);
or U26871 (N_26871,N_25692,N_25347);
nor U26872 (N_26872,N_25002,N_24636);
or U26873 (N_26873,N_25503,N_25000);
and U26874 (N_26874,N_25801,N_24792);
or U26875 (N_26875,N_24723,N_24465);
xor U26876 (N_26876,N_24653,N_25577);
or U26877 (N_26877,N_25029,N_24214);
or U26878 (N_26878,N_24211,N_25642);
nand U26879 (N_26879,N_24727,N_24616);
or U26880 (N_26880,N_24301,N_25656);
nor U26881 (N_26881,N_25160,N_25806);
xnor U26882 (N_26882,N_24801,N_25341);
or U26883 (N_26883,N_25889,N_24198);
nand U26884 (N_26884,N_24873,N_24715);
or U26885 (N_26885,N_24494,N_24864);
or U26886 (N_26886,N_24921,N_24246);
xnor U26887 (N_26887,N_24206,N_24954);
nand U26888 (N_26888,N_25135,N_25760);
nand U26889 (N_26889,N_24030,N_25373);
or U26890 (N_26890,N_24115,N_25158);
nand U26891 (N_26891,N_24323,N_25548);
or U26892 (N_26892,N_24583,N_25458);
nor U26893 (N_26893,N_25358,N_24507);
and U26894 (N_26894,N_24794,N_24861);
nor U26895 (N_26895,N_24190,N_25050);
nand U26896 (N_26896,N_25034,N_24165);
and U26897 (N_26897,N_25935,N_24660);
nor U26898 (N_26898,N_24126,N_24324);
and U26899 (N_26899,N_25381,N_25653);
nand U26900 (N_26900,N_24405,N_24284);
xnor U26901 (N_26901,N_25901,N_25645);
xor U26902 (N_26902,N_25068,N_24509);
xor U26903 (N_26903,N_24446,N_25857);
or U26904 (N_26904,N_24652,N_25542);
nand U26905 (N_26905,N_25113,N_25598);
and U26906 (N_26906,N_24516,N_24656);
or U26907 (N_26907,N_24267,N_24131);
and U26908 (N_26908,N_25134,N_25543);
or U26909 (N_26909,N_24003,N_24838);
xor U26910 (N_26910,N_25518,N_25306);
or U26911 (N_26911,N_24292,N_24712);
or U26912 (N_26912,N_24356,N_25272);
xor U26913 (N_26913,N_25530,N_24305);
or U26914 (N_26914,N_25832,N_25316);
and U26915 (N_26915,N_25647,N_25184);
or U26916 (N_26916,N_25841,N_24382);
xor U26917 (N_26917,N_24645,N_24905);
and U26918 (N_26918,N_24491,N_24464);
nor U26919 (N_26919,N_25742,N_25477);
nor U26920 (N_26920,N_24536,N_24046);
nand U26921 (N_26921,N_24470,N_24815);
nand U26922 (N_26922,N_24885,N_24341);
or U26923 (N_26923,N_24472,N_25351);
nor U26924 (N_26924,N_25248,N_24982);
nor U26925 (N_26925,N_25354,N_24282);
nor U26926 (N_26926,N_24417,N_25706);
and U26927 (N_26927,N_25963,N_25069);
or U26928 (N_26928,N_24287,N_24427);
or U26929 (N_26929,N_25938,N_24545);
and U26930 (N_26930,N_24899,N_24059);
nand U26931 (N_26931,N_24914,N_25171);
xor U26932 (N_26932,N_25422,N_24278);
nand U26933 (N_26933,N_25637,N_24579);
nor U26934 (N_26934,N_25155,N_24118);
xnor U26935 (N_26935,N_25936,N_25194);
or U26936 (N_26936,N_24892,N_25294);
xor U26937 (N_26937,N_25357,N_25564);
nand U26938 (N_26938,N_24699,N_25081);
nor U26939 (N_26939,N_25228,N_25335);
nor U26940 (N_26940,N_24842,N_24938);
nor U26941 (N_26941,N_25346,N_25247);
and U26942 (N_26942,N_24139,N_25638);
or U26943 (N_26943,N_24339,N_24462);
and U26944 (N_26944,N_25996,N_24412);
xor U26945 (N_26945,N_25630,N_25121);
nand U26946 (N_26946,N_25898,N_24779);
nor U26947 (N_26947,N_25827,N_25615);
or U26948 (N_26948,N_24527,N_24612);
nand U26949 (N_26949,N_24730,N_25461);
or U26950 (N_26950,N_24273,N_25812);
nand U26951 (N_26951,N_25703,N_24584);
nand U26952 (N_26952,N_25660,N_24762);
and U26953 (N_26953,N_25009,N_25274);
or U26954 (N_26954,N_24740,N_24820);
xnor U26955 (N_26955,N_25691,N_24983);
nand U26956 (N_26956,N_24377,N_25257);
nand U26957 (N_26957,N_24927,N_24854);
and U26958 (N_26958,N_24952,N_24461);
or U26959 (N_26959,N_25123,N_24846);
nor U26960 (N_26960,N_24831,N_25608);
xor U26961 (N_26961,N_24573,N_25913);
and U26962 (N_26962,N_25928,N_24180);
nor U26963 (N_26963,N_25414,N_25870);
xnor U26964 (N_26964,N_24980,N_25076);
nor U26965 (N_26965,N_24889,N_25879);
or U26966 (N_26966,N_25675,N_24680);
xor U26967 (N_26967,N_25222,N_24084);
and U26968 (N_26968,N_24848,N_25342);
nor U26969 (N_26969,N_25758,N_25497);
or U26970 (N_26970,N_24251,N_25092);
and U26971 (N_26971,N_25864,N_24700);
and U26972 (N_26972,N_24789,N_24262);
nor U26973 (N_26973,N_24929,N_25662);
nor U26974 (N_26974,N_24976,N_25597);
and U26975 (N_26975,N_25129,N_24263);
and U26976 (N_26976,N_25909,N_24597);
xor U26977 (N_26977,N_25252,N_25755);
and U26978 (N_26978,N_24985,N_25749);
nand U26979 (N_26979,N_24361,N_25764);
nand U26980 (N_26980,N_24915,N_24963);
nand U26981 (N_26981,N_25521,N_24144);
or U26982 (N_26982,N_25979,N_24200);
nor U26983 (N_26983,N_24713,N_25330);
nor U26984 (N_26984,N_24558,N_24032);
nor U26985 (N_26985,N_24087,N_24923);
and U26986 (N_26986,N_24658,N_25425);
and U26987 (N_26987,N_25570,N_24492);
or U26988 (N_26988,N_25894,N_25072);
xor U26989 (N_26989,N_24955,N_25574);
nand U26990 (N_26990,N_25569,N_24048);
nor U26991 (N_26991,N_25128,N_25558);
nand U26992 (N_26992,N_24765,N_25387);
nand U26993 (N_26993,N_25796,N_24887);
nor U26994 (N_26994,N_25536,N_24895);
nor U26995 (N_26995,N_25861,N_24676);
nor U26996 (N_26996,N_24999,N_24565);
xnor U26997 (N_26997,N_24090,N_25325);
nand U26998 (N_26998,N_24421,N_24250);
and U26999 (N_26999,N_24050,N_25772);
nand U27000 (N_27000,N_25970,N_25869);
or U27001 (N_27001,N_24438,N_25129);
xor U27002 (N_27002,N_24585,N_24821);
nand U27003 (N_27003,N_24137,N_25993);
nor U27004 (N_27004,N_24152,N_24903);
nand U27005 (N_27005,N_25369,N_25474);
xor U27006 (N_27006,N_24103,N_25912);
and U27007 (N_27007,N_25852,N_24925);
and U27008 (N_27008,N_24470,N_24013);
xor U27009 (N_27009,N_25055,N_24661);
xor U27010 (N_27010,N_24853,N_25606);
xor U27011 (N_27011,N_25460,N_24059);
and U27012 (N_27012,N_24294,N_25277);
nor U27013 (N_27013,N_24150,N_25346);
nand U27014 (N_27014,N_25289,N_24153);
nand U27015 (N_27015,N_24843,N_24714);
and U27016 (N_27016,N_24825,N_25098);
or U27017 (N_27017,N_24207,N_24967);
and U27018 (N_27018,N_24770,N_24625);
nor U27019 (N_27019,N_24136,N_24028);
nor U27020 (N_27020,N_25027,N_24803);
nor U27021 (N_27021,N_24175,N_24712);
xnor U27022 (N_27022,N_25845,N_25941);
and U27023 (N_27023,N_25054,N_24196);
xor U27024 (N_27024,N_24320,N_24316);
and U27025 (N_27025,N_25123,N_25914);
nor U27026 (N_27026,N_25389,N_24356);
and U27027 (N_27027,N_24787,N_25696);
xor U27028 (N_27028,N_24042,N_25848);
xnor U27029 (N_27029,N_24977,N_25417);
nor U27030 (N_27030,N_25779,N_24936);
or U27031 (N_27031,N_24403,N_25248);
and U27032 (N_27032,N_24701,N_25148);
nand U27033 (N_27033,N_25519,N_25743);
or U27034 (N_27034,N_25303,N_25201);
nor U27035 (N_27035,N_24997,N_25632);
nor U27036 (N_27036,N_24756,N_25669);
and U27037 (N_27037,N_25409,N_24445);
nor U27038 (N_27038,N_24273,N_25846);
xnor U27039 (N_27039,N_25442,N_25485);
xnor U27040 (N_27040,N_25002,N_25886);
and U27041 (N_27041,N_25390,N_24250);
nand U27042 (N_27042,N_24051,N_24128);
nor U27043 (N_27043,N_24128,N_25187);
nor U27044 (N_27044,N_25949,N_24469);
and U27045 (N_27045,N_24269,N_24677);
or U27046 (N_27046,N_25042,N_25175);
nand U27047 (N_27047,N_25324,N_25095);
xnor U27048 (N_27048,N_24225,N_25292);
nand U27049 (N_27049,N_25466,N_24733);
and U27050 (N_27050,N_24751,N_24458);
nor U27051 (N_27051,N_25442,N_24634);
nand U27052 (N_27052,N_24787,N_24274);
xnor U27053 (N_27053,N_25077,N_24630);
xnor U27054 (N_27054,N_25097,N_25243);
or U27055 (N_27055,N_25619,N_24356);
xnor U27056 (N_27056,N_24787,N_24942);
nand U27057 (N_27057,N_25781,N_24752);
nor U27058 (N_27058,N_24595,N_25502);
or U27059 (N_27059,N_25117,N_25892);
xor U27060 (N_27060,N_24024,N_25075);
or U27061 (N_27061,N_25076,N_24321);
xnor U27062 (N_27062,N_24233,N_25938);
nand U27063 (N_27063,N_24558,N_25524);
and U27064 (N_27064,N_24123,N_25813);
xor U27065 (N_27065,N_25249,N_24845);
or U27066 (N_27066,N_24538,N_25768);
or U27067 (N_27067,N_25945,N_24635);
nor U27068 (N_27068,N_25560,N_25972);
and U27069 (N_27069,N_25652,N_24270);
nand U27070 (N_27070,N_24619,N_25003);
nand U27071 (N_27071,N_25385,N_25424);
or U27072 (N_27072,N_25918,N_25198);
xor U27073 (N_27073,N_24097,N_24541);
or U27074 (N_27074,N_24095,N_24684);
xor U27075 (N_27075,N_25206,N_25893);
nor U27076 (N_27076,N_25461,N_25989);
or U27077 (N_27077,N_25391,N_24565);
and U27078 (N_27078,N_24983,N_25813);
and U27079 (N_27079,N_24903,N_24386);
nor U27080 (N_27080,N_24821,N_25413);
or U27081 (N_27081,N_25806,N_24739);
xnor U27082 (N_27082,N_25856,N_25519);
or U27083 (N_27083,N_25176,N_25189);
nand U27084 (N_27084,N_24744,N_25318);
and U27085 (N_27085,N_25182,N_25588);
and U27086 (N_27086,N_24740,N_25363);
xnor U27087 (N_27087,N_24031,N_25149);
nor U27088 (N_27088,N_24374,N_24729);
and U27089 (N_27089,N_24385,N_24018);
xnor U27090 (N_27090,N_25195,N_24457);
nand U27091 (N_27091,N_25638,N_25443);
xnor U27092 (N_27092,N_24606,N_24000);
nand U27093 (N_27093,N_24250,N_25617);
xor U27094 (N_27094,N_24480,N_24748);
and U27095 (N_27095,N_25859,N_25974);
or U27096 (N_27096,N_25847,N_24723);
nor U27097 (N_27097,N_25076,N_24060);
xor U27098 (N_27098,N_25501,N_25737);
nand U27099 (N_27099,N_24337,N_24193);
and U27100 (N_27100,N_25664,N_25892);
or U27101 (N_27101,N_24675,N_24638);
nor U27102 (N_27102,N_24037,N_24708);
and U27103 (N_27103,N_25235,N_24604);
or U27104 (N_27104,N_25919,N_24252);
or U27105 (N_27105,N_24179,N_25224);
nor U27106 (N_27106,N_24919,N_24293);
xor U27107 (N_27107,N_24059,N_25363);
or U27108 (N_27108,N_24181,N_24327);
and U27109 (N_27109,N_25826,N_25070);
xnor U27110 (N_27110,N_24662,N_25625);
nor U27111 (N_27111,N_24217,N_25676);
and U27112 (N_27112,N_24909,N_25374);
nor U27113 (N_27113,N_25283,N_25755);
and U27114 (N_27114,N_25900,N_25234);
nand U27115 (N_27115,N_25923,N_25451);
nor U27116 (N_27116,N_25647,N_24387);
nand U27117 (N_27117,N_25817,N_24954);
and U27118 (N_27118,N_25425,N_25085);
nand U27119 (N_27119,N_25271,N_24692);
and U27120 (N_27120,N_25550,N_25204);
nand U27121 (N_27121,N_25688,N_25318);
xor U27122 (N_27122,N_25552,N_24870);
nand U27123 (N_27123,N_24404,N_25216);
nand U27124 (N_27124,N_24424,N_24716);
and U27125 (N_27125,N_24180,N_24793);
or U27126 (N_27126,N_24265,N_25548);
xnor U27127 (N_27127,N_24783,N_25948);
xnor U27128 (N_27128,N_24913,N_24297);
xor U27129 (N_27129,N_24258,N_25741);
xor U27130 (N_27130,N_25754,N_24608);
nor U27131 (N_27131,N_25135,N_25974);
and U27132 (N_27132,N_25104,N_25650);
or U27133 (N_27133,N_24700,N_25734);
or U27134 (N_27134,N_24313,N_24853);
and U27135 (N_27135,N_25651,N_24217);
nand U27136 (N_27136,N_25951,N_25982);
xnor U27137 (N_27137,N_25164,N_24380);
nor U27138 (N_27138,N_24283,N_25697);
xor U27139 (N_27139,N_25977,N_25601);
or U27140 (N_27140,N_25336,N_24070);
nor U27141 (N_27141,N_24424,N_25345);
nand U27142 (N_27142,N_24426,N_25400);
or U27143 (N_27143,N_25995,N_25857);
and U27144 (N_27144,N_24812,N_25894);
nand U27145 (N_27145,N_25137,N_25622);
and U27146 (N_27146,N_24600,N_24659);
nand U27147 (N_27147,N_25026,N_24557);
nand U27148 (N_27148,N_24772,N_25053);
and U27149 (N_27149,N_24304,N_24374);
or U27150 (N_27150,N_25766,N_25016);
xnor U27151 (N_27151,N_24156,N_25950);
nand U27152 (N_27152,N_24144,N_25162);
nand U27153 (N_27153,N_24070,N_24922);
and U27154 (N_27154,N_24797,N_24398);
or U27155 (N_27155,N_25697,N_24375);
or U27156 (N_27156,N_25328,N_25651);
nand U27157 (N_27157,N_24774,N_25885);
xor U27158 (N_27158,N_25871,N_25729);
xor U27159 (N_27159,N_25113,N_25460);
and U27160 (N_27160,N_25903,N_25588);
nor U27161 (N_27161,N_25525,N_24314);
nor U27162 (N_27162,N_25110,N_24039);
xor U27163 (N_27163,N_24166,N_24276);
and U27164 (N_27164,N_24671,N_25263);
and U27165 (N_27165,N_24750,N_24445);
xor U27166 (N_27166,N_25370,N_24693);
or U27167 (N_27167,N_25412,N_25740);
nand U27168 (N_27168,N_25009,N_24116);
and U27169 (N_27169,N_24125,N_25935);
and U27170 (N_27170,N_25704,N_25111);
nor U27171 (N_27171,N_25400,N_24732);
and U27172 (N_27172,N_25970,N_25174);
or U27173 (N_27173,N_24300,N_25938);
nand U27174 (N_27174,N_25019,N_24029);
or U27175 (N_27175,N_25969,N_24381);
nor U27176 (N_27176,N_24201,N_24923);
nand U27177 (N_27177,N_24131,N_24278);
nand U27178 (N_27178,N_24419,N_24597);
nand U27179 (N_27179,N_25415,N_25634);
or U27180 (N_27180,N_24143,N_25335);
or U27181 (N_27181,N_24901,N_25539);
and U27182 (N_27182,N_24522,N_24417);
xnor U27183 (N_27183,N_25130,N_24385);
nand U27184 (N_27184,N_25928,N_24988);
nor U27185 (N_27185,N_24348,N_25828);
xnor U27186 (N_27186,N_24638,N_24850);
and U27187 (N_27187,N_24996,N_24452);
nand U27188 (N_27188,N_24463,N_24390);
and U27189 (N_27189,N_24965,N_25553);
nor U27190 (N_27190,N_25951,N_25323);
and U27191 (N_27191,N_25912,N_25374);
and U27192 (N_27192,N_25068,N_25599);
or U27193 (N_27193,N_24513,N_25545);
and U27194 (N_27194,N_24857,N_25292);
nor U27195 (N_27195,N_25715,N_24465);
and U27196 (N_27196,N_25918,N_25434);
and U27197 (N_27197,N_25784,N_24726);
xnor U27198 (N_27198,N_25347,N_24191);
nor U27199 (N_27199,N_24046,N_25282);
or U27200 (N_27200,N_24268,N_24571);
xor U27201 (N_27201,N_25706,N_25947);
nand U27202 (N_27202,N_24162,N_25009);
and U27203 (N_27203,N_24620,N_25788);
or U27204 (N_27204,N_24070,N_25569);
or U27205 (N_27205,N_25127,N_24152);
nand U27206 (N_27206,N_25138,N_25934);
nor U27207 (N_27207,N_24726,N_25426);
xnor U27208 (N_27208,N_25743,N_25474);
nor U27209 (N_27209,N_25172,N_24503);
and U27210 (N_27210,N_24580,N_25229);
or U27211 (N_27211,N_25234,N_25769);
or U27212 (N_27212,N_25103,N_25080);
nor U27213 (N_27213,N_24909,N_24241);
xor U27214 (N_27214,N_25273,N_24102);
or U27215 (N_27215,N_25589,N_24140);
nor U27216 (N_27216,N_24513,N_25762);
nand U27217 (N_27217,N_25926,N_25145);
nand U27218 (N_27218,N_24587,N_24842);
xnor U27219 (N_27219,N_25720,N_24162);
or U27220 (N_27220,N_24657,N_25308);
xor U27221 (N_27221,N_25221,N_24267);
nand U27222 (N_27222,N_25411,N_25436);
or U27223 (N_27223,N_25747,N_24989);
xnor U27224 (N_27224,N_25561,N_25174);
xnor U27225 (N_27225,N_25697,N_25369);
and U27226 (N_27226,N_24470,N_25757);
and U27227 (N_27227,N_24277,N_24261);
xnor U27228 (N_27228,N_24788,N_25897);
nand U27229 (N_27229,N_24859,N_25362);
nand U27230 (N_27230,N_25127,N_25322);
nor U27231 (N_27231,N_25750,N_24785);
nand U27232 (N_27232,N_25133,N_24017);
nor U27233 (N_27233,N_24029,N_25172);
and U27234 (N_27234,N_25896,N_24829);
nor U27235 (N_27235,N_24798,N_24720);
nand U27236 (N_27236,N_25978,N_24092);
or U27237 (N_27237,N_25609,N_25074);
nand U27238 (N_27238,N_24095,N_24819);
or U27239 (N_27239,N_25602,N_25498);
nor U27240 (N_27240,N_25214,N_25342);
nor U27241 (N_27241,N_25738,N_25430);
nand U27242 (N_27242,N_25578,N_25263);
nor U27243 (N_27243,N_25165,N_24862);
nand U27244 (N_27244,N_25765,N_25823);
nand U27245 (N_27245,N_25261,N_25259);
xnor U27246 (N_27246,N_25910,N_25640);
and U27247 (N_27247,N_25592,N_25004);
nor U27248 (N_27248,N_25197,N_25647);
nand U27249 (N_27249,N_25483,N_25992);
nor U27250 (N_27250,N_24279,N_24007);
nand U27251 (N_27251,N_25928,N_24547);
or U27252 (N_27252,N_24243,N_25246);
or U27253 (N_27253,N_24994,N_24069);
nor U27254 (N_27254,N_25529,N_24805);
and U27255 (N_27255,N_24026,N_24825);
xor U27256 (N_27256,N_24254,N_24801);
nor U27257 (N_27257,N_25566,N_24300);
xnor U27258 (N_27258,N_25671,N_25739);
nor U27259 (N_27259,N_25697,N_25018);
nand U27260 (N_27260,N_25145,N_25319);
nor U27261 (N_27261,N_24365,N_24975);
xor U27262 (N_27262,N_25454,N_24867);
nor U27263 (N_27263,N_25013,N_24901);
and U27264 (N_27264,N_25268,N_25874);
or U27265 (N_27265,N_25197,N_24390);
xor U27266 (N_27266,N_24806,N_25659);
and U27267 (N_27267,N_24690,N_24083);
and U27268 (N_27268,N_25582,N_25884);
or U27269 (N_27269,N_24652,N_24035);
nand U27270 (N_27270,N_24797,N_25886);
nand U27271 (N_27271,N_25766,N_25042);
nand U27272 (N_27272,N_24104,N_25287);
nand U27273 (N_27273,N_24488,N_24642);
and U27274 (N_27274,N_25303,N_25854);
nand U27275 (N_27275,N_24593,N_25236);
nand U27276 (N_27276,N_25305,N_24774);
and U27277 (N_27277,N_25623,N_24058);
nor U27278 (N_27278,N_25150,N_25769);
or U27279 (N_27279,N_25312,N_24371);
or U27280 (N_27280,N_25769,N_24330);
nand U27281 (N_27281,N_24779,N_25363);
xor U27282 (N_27282,N_24319,N_24770);
nand U27283 (N_27283,N_24193,N_24070);
xor U27284 (N_27284,N_24228,N_24337);
xor U27285 (N_27285,N_25783,N_25988);
nor U27286 (N_27286,N_24070,N_25241);
or U27287 (N_27287,N_24418,N_24380);
and U27288 (N_27288,N_25498,N_25798);
nand U27289 (N_27289,N_24131,N_24646);
xnor U27290 (N_27290,N_24154,N_25422);
nand U27291 (N_27291,N_24108,N_24375);
nor U27292 (N_27292,N_24161,N_25454);
or U27293 (N_27293,N_25624,N_25325);
nand U27294 (N_27294,N_25682,N_24552);
nor U27295 (N_27295,N_25985,N_25027);
or U27296 (N_27296,N_24520,N_24274);
xor U27297 (N_27297,N_25144,N_24643);
xor U27298 (N_27298,N_24929,N_25262);
nor U27299 (N_27299,N_25930,N_24272);
nor U27300 (N_27300,N_25063,N_25011);
xor U27301 (N_27301,N_24954,N_25389);
or U27302 (N_27302,N_24845,N_25107);
nand U27303 (N_27303,N_24965,N_25870);
xnor U27304 (N_27304,N_24914,N_24450);
and U27305 (N_27305,N_24422,N_24129);
xnor U27306 (N_27306,N_25969,N_25006);
xnor U27307 (N_27307,N_25113,N_24354);
nor U27308 (N_27308,N_25242,N_24395);
and U27309 (N_27309,N_24036,N_24895);
and U27310 (N_27310,N_25386,N_24616);
or U27311 (N_27311,N_25508,N_24510);
and U27312 (N_27312,N_25736,N_25460);
nand U27313 (N_27313,N_25399,N_25513);
nor U27314 (N_27314,N_25698,N_25335);
nand U27315 (N_27315,N_25725,N_25942);
xnor U27316 (N_27316,N_25377,N_25097);
nand U27317 (N_27317,N_25356,N_25530);
nor U27318 (N_27318,N_25112,N_24518);
nand U27319 (N_27319,N_24863,N_25869);
or U27320 (N_27320,N_24318,N_24955);
nor U27321 (N_27321,N_24370,N_24905);
or U27322 (N_27322,N_24100,N_25020);
or U27323 (N_27323,N_24181,N_24082);
and U27324 (N_27324,N_24277,N_24599);
nand U27325 (N_27325,N_24541,N_25357);
or U27326 (N_27326,N_25182,N_25657);
and U27327 (N_27327,N_24685,N_24567);
xnor U27328 (N_27328,N_25104,N_25434);
xor U27329 (N_27329,N_24588,N_25950);
and U27330 (N_27330,N_24958,N_25400);
and U27331 (N_27331,N_24899,N_25795);
nor U27332 (N_27332,N_24916,N_24618);
nor U27333 (N_27333,N_24407,N_25436);
nor U27334 (N_27334,N_24706,N_24409);
xor U27335 (N_27335,N_24751,N_25749);
nand U27336 (N_27336,N_25155,N_25563);
and U27337 (N_27337,N_24690,N_25488);
and U27338 (N_27338,N_25924,N_24636);
nor U27339 (N_27339,N_24804,N_25460);
or U27340 (N_27340,N_24414,N_24571);
nor U27341 (N_27341,N_24165,N_25565);
nor U27342 (N_27342,N_24206,N_25190);
nor U27343 (N_27343,N_24512,N_24598);
nand U27344 (N_27344,N_25737,N_25687);
or U27345 (N_27345,N_25127,N_24490);
xor U27346 (N_27346,N_24722,N_25767);
nand U27347 (N_27347,N_24738,N_24793);
or U27348 (N_27348,N_24933,N_25584);
and U27349 (N_27349,N_24706,N_25077);
nor U27350 (N_27350,N_25134,N_25392);
xnor U27351 (N_27351,N_24431,N_25852);
nand U27352 (N_27352,N_25865,N_25858);
nand U27353 (N_27353,N_25193,N_24502);
nand U27354 (N_27354,N_25424,N_24036);
or U27355 (N_27355,N_25604,N_25584);
or U27356 (N_27356,N_25390,N_25968);
nor U27357 (N_27357,N_24975,N_25085);
or U27358 (N_27358,N_25202,N_24335);
and U27359 (N_27359,N_25939,N_25756);
and U27360 (N_27360,N_25469,N_25299);
or U27361 (N_27361,N_24060,N_25443);
xnor U27362 (N_27362,N_25873,N_24533);
xnor U27363 (N_27363,N_24436,N_24767);
or U27364 (N_27364,N_24933,N_25464);
and U27365 (N_27365,N_25981,N_24402);
and U27366 (N_27366,N_24883,N_24036);
and U27367 (N_27367,N_25239,N_24229);
nor U27368 (N_27368,N_24565,N_25801);
and U27369 (N_27369,N_24291,N_25794);
nor U27370 (N_27370,N_24923,N_25050);
and U27371 (N_27371,N_24894,N_25753);
and U27372 (N_27372,N_24556,N_24781);
or U27373 (N_27373,N_25211,N_25392);
nand U27374 (N_27374,N_25253,N_24968);
xnor U27375 (N_27375,N_25120,N_25549);
and U27376 (N_27376,N_25713,N_24901);
or U27377 (N_27377,N_24620,N_24904);
nor U27378 (N_27378,N_25874,N_24612);
nor U27379 (N_27379,N_24018,N_24275);
or U27380 (N_27380,N_24561,N_25096);
xnor U27381 (N_27381,N_25047,N_24531);
or U27382 (N_27382,N_24718,N_24444);
or U27383 (N_27383,N_24675,N_25908);
nor U27384 (N_27384,N_25232,N_25581);
nand U27385 (N_27385,N_24946,N_25067);
and U27386 (N_27386,N_24393,N_25146);
or U27387 (N_27387,N_24134,N_25883);
and U27388 (N_27388,N_25222,N_25714);
xor U27389 (N_27389,N_24014,N_25777);
xor U27390 (N_27390,N_25452,N_24054);
nor U27391 (N_27391,N_25775,N_25473);
xnor U27392 (N_27392,N_24285,N_25131);
xor U27393 (N_27393,N_25914,N_25902);
and U27394 (N_27394,N_25175,N_25004);
xor U27395 (N_27395,N_24609,N_24301);
or U27396 (N_27396,N_25022,N_25145);
and U27397 (N_27397,N_24126,N_25425);
and U27398 (N_27398,N_25298,N_24351);
and U27399 (N_27399,N_24159,N_24114);
nor U27400 (N_27400,N_24538,N_24200);
nand U27401 (N_27401,N_24796,N_25208);
nand U27402 (N_27402,N_24447,N_24048);
nand U27403 (N_27403,N_24287,N_24220);
nor U27404 (N_27404,N_25998,N_25212);
and U27405 (N_27405,N_25963,N_24157);
and U27406 (N_27406,N_24201,N_25815);
and U27407 (N_27407,N_25915,N_24795);
xor U27408 (N_27408,N_25277,N_24341);
and U27409 (N_27409,N_24744,N_24669);
xnor U27410 (N_27410,N_25169,N_24117);
nand U27411 (N_27411,N_24252,N_25259);
or U27412 (N_27412,N_24077,N_25477);
xnor U27413 (N_27413,N_25244,N_24215);
nor U27414 (N_27414,N_24623,N_25537);
xnor U27415 (N_27415,N_24192,N_24430);
and U27416 (N_27416,N_25805,N_24190);
or U27417 (N_27417,N_25980,N_24108);
nand U27418 (N_27418,N_24315,N_25497);
nor U27419 (N_27419,N_25795,N_24334);
and U27420 (N_27420,N_25277,N_24539);
and U27421 (N_27421,N_24065,N_24644);
xnor U27422 (N_27422,N_24822,N_25448);
nor U27423 (N_27423,N_24987,N_24096);
nor U27424 (N_27424,N_25491,N_24820);
nand U27425 (N_27425,N_25192,N_24436);
and U27426 (N_27426,N_25847,N_25819);
or U27427 (N_27427,N_24451,N_25000);
and U27428 (N_27428,N_24320,N_25253);
or U27429 (N_27429,N_24553,N_24982);
or U27430 (N_27430,N_25494,N_25445);
and U27431 (N_27431,N_25490,N_25606);
nand U27432 (N_27432,N_24799,N_24034);
xor U27433 (N_27433,N_24532,N_24619);
and U27434 (N_27434,N_25249,N_24770);
and U27435 (N_27435,N_24614,N_24576);
nor U27436 (N_27436,N_24904,N_25901);
or U27437 (N_27437,N_25586,N_24638);
and U27438 (N_27438,N_25121,N_25412);
nor U27439 (N_27439,N_24444,N_24768);
nand U27440 (N_27440,N_24608,N_24486);
nor U27441 (N_27441,N_25712,N_25936);
nor U27442 (N_27442,N_25142,N_25331);
or U27443 (N_27443,N_24662,N_24238);
nand U27444 (N_27444,N_25058,N_24660);
or U27445 (N_27445,N_24843,N_24111);
nor U27446 (N_27446,N_25249,N_24843);
nand U27447 (N_27447,N_25441,N_25631);
or U27448 (N_27448,N_24020,N_24891);
xnor U27449 (N_27449,N_25173,N_25201);
and U27450 (N_27450,N_25808,N_25909);
or U27451 (N_27451,N_24791,N_24342);
nor U27452 (N_27452,N_24709,N_25683);
or U27453 (N_27453,N_25756,N_24126);
nor U27454 (N_27454,N_25539,N_24192);
or U27455 (N_27455,N_25875,N_25708);
nor U27456 (N_27456,N_25365,N_24390);
nor U27457 (N_27457,N_24609,N_24204);
nor U27458 (N_27458,N_25803,N_25702);
nand U27459 (N_27459,N_24614,N_24310);
xor U27460 (N_27460,N_25503,N_25696);
and U27461 (N_27461,N_25557,N_24473);
and U27462 (N_27462,N_25275,N_25240);
or U27463 (N_27463,N_25099,N_24541);
nand U27464 (N_27464,N_24427,N_25548);
nor U27465 (N_27465,N_24679,N_25684);
nand U27466 (N_27466,N_25264,N_24534);
and U27467 (N_27467,N_25673,N_25569);
nand U27468 (N_27468,N_25811,N_24959);
xor U27469 (N_27469,N_25223,N_25095);
and U27470 (N_27470,N_25699,N_25736);
and U27471 (N_27471,N_25251,N_24474);
or U27472 (N_27472,N_24786,N_24661);
and U27473 (N_27473,N_25608,N_25442);
or U27474 (N_27474,N_24309,N_25056);
or U27475 (N_27475,N_25266,N_25359);
xor U27476 (N_27476,N_25015,N_24278);
and U27477 (N_27477,N_24990,N_25787);
and U27478 (N_27478,N_25990,N_25593);
xor U27479 (N_27479,N_25954,N_24896);
or U27480 (N_27480,N_24016,N_25080);
nand U27481 (N_27481,N_25263,N_25424);
or U27482 (N_27482,N_25176,N_25909);
nor U27483 (N_27483,N_24310,N_25117);
nor U27484 (N_27484,N_24031,N_25407);
nor U27485 (N_27485,N_24561,N_24727);
and U27486 (N_27486,N_25440,N_25206);
or U27487 (N_27487,N_25461,N_24546);
xnor U27488 (N_27488,N_25142,N_24689);
or U27489 (N_27489,N_24485,N_24586);
and U27490 (N_27490,N_24829,N_25479);
xnor U27491 (N_27491,N_24025,N_25264);
nand U27492 (N_27492,N_25444,N_25532);
xor U27493 (N_27493,N_25671,N_24810);
xnor U27494 (N_27494,N_25547,N_24734);
or U27495 (N_27495,N_25567,N_25743);
and U27496 (N_27496,N_25640,N_25099);
nand U27497 (N_27497,N_25980,N_24531);
or U27498 (N_27498,N_24983,N_25076);
nand U27499 (N_27499,N_24097,N_24466);
nor U27500 (N_27500,N_24851,N_24743);
nor U27501 (N_27501,N_25619,N_24256);
and U27502 (N_27502,N_24212,N_25685);
nor U27503 (N_27503,N_25191,N_24286);
nor U27504 (N_27504,N_25585,N_24895);
nor U27505 (N_27505,N_24603,N_25920);
or U27506 (N_27506,N_25674,N_24399);
xor U27507 (N_27507,N_25885,N_24128);
xor U27508 (N_27508,N_25098,N_25022);
nand U27509 (N_27509,N_25415,N_24361);
and U27510 (N_27510,N_24037,N_24167);
or U27511 (N_27511,N_25255,N_24135);
nand U27512 (N_27512,N_25309,N_24206);
or U27513 (N_27513,N_24631,N_24682);
xnor U27514 (N_27514,N_24587,N_25133);
nand U27515 (N_27515,N_25700,N_25614);
or U27516 (N_27516,N_24286,N_24956);
or U27517 (N_27517,N_24114,N_25280);
or U27518 (N_27518,N_25358,N_25055);
and U27519 (N_27519,N_25954,N_24683);
nand U27520 (N_27520,N_25465,N_24735);
nand U27521 (N_27521,N_25290,N_25329);
or U27522 (N_27522,N_25813,N_24307);
nand U27523 (N_27523,N_24063,N_25436);
xnor U27524 (N_27524,N_24209,N_24717);
xnor U27525 (N_27525,N_24883,N_25398);
or U27526 (N_27526,N_25292,N_25927);
nor U27527 (N_27527,N_24146,N_24665);
nand U27528 (N_27528,N_24236,N_24475);
nand U27529 (N_27529,N_25399,N_24472);
nand U27530 (N_27530,N_24985,N_24261);
nand U27531 (N_27531,N_24818,N_24374);
and U27532 (N_27532,N_25899,N_25718);
or U27533 (N_27533,N_25022,N_25348);
and U27534 (N_27534,N_25491,N_24669);
xor U27535 (N_27535,N_24612,N_24294);
nor U27536 (N_27536,N_24762,N_25254);
nor U27537 (N_27537,N_25884,N_24262);
or U27538 (N_27538,N_24087,N_25029);
xor U27539 (N_27539,N_24634,N_25761);
and U27540 (N_27540,N_24165,N_24611);
nand U27541 (N_27541,N_24491,N_24856);
nor U27542 (N_27542,N_25541,N_24378);
or U27543 (N_27543,N_25025,N_25985);
nand U27544 (N_27544,N_25156,N_25861);
nor U27545 (N_27545,N_24978,N_25398);
and U27546 (N_27546,N_25665,N_24502);
nor U27547 (N_27547,N_24893,N_24582);
nor U27548 (N_27548,N_24475,N_25368);
nand U27549 (N_27549,N_25197,N_25577);
nor U27550 (N_27550,N_24938,N_24869);
nand U27551 (N_27551,N_25517,N_24759);
and U27552 (N_27552,N_24993,N_24496);
nand U27553 (N_27553,N_25006,N_24363);
or U27554 (N_27554,N_25838,N_25038);
or U27555 (N_27555,N_25832,N_25406);
xnor U27556 (N_27556,N_25949,N_25396);
or U27557 (N_27557,N_24648,N_24521);
xnor U27558 (N_27558,N_24160,N_25547);
and U27559 (N_27559,N_25192,N_24983);
or U27560 (N_27560,N_25179,N_25041);
xnor U27561 (N_27561,N_25614,N_24240);
and U27562 (N_27562,N_24831,N_24649);
or U27563 (N_27563,N_24128,N_25575);
nand U27564 (N_27564,N_25079,N_25579);
nand U27565 (N_27565,N_24693,N_25294);
nor U27566 (N_27566,N_25805,N_25272);
or U27567 (N_27567,N_25839,N_25379);
nand U27568 (N_27568,N_24494,N_25175);
nor U27569 (N_27569,N_25449,N_24376);
nor U27570 (N_27570,N_24424,N_25324);
nor U27571 (N_27571,N_24800,N_25393);
or U27572 (N_27572,N_25445,N_24936);
nand U27573 (N_27573,N_25913,N_24990);
nor U27574 (N_27574,N_25384,N_25382);
or U27575 (N_27575,N_24146,N_25674);
xnor U27576 (N_27576,N_25516,N_25290);
nand U27577 (N_27577,N_25197,N_24051);
nor U27578 (N_27578,N_24675,N_25347);
xnor U27579 (N_27579,N_25013,N_24953);
nand U27580 (N_27580,N_25988,N_24025);
nor U27581 (N_27581,N_25279,N_25664);
xnor U27582 (N_27582,N_25271,N_24162);
and U27583 (N_27583,N_25841,N_24463);
nand U27584 (N_27584,N_24837,N_25143);
xnor U27585 (N_27585,N_24990,N_25179);
xnor U27586 (N_27586,N_25702,N_25160);
xor U27587 (N_27587,N_24811,N_25798);
nand U27588 (N_27588,N_24576,N_25450);
and U27589 (N_27589,N_24422,N_24874);
and U27590 (N_27590,N_24085,N_25360);
or U27591 (N_27591,N_24270,N_24088);
or U27592 (N_27592,N_24130,N_24198);
nor U27593 (N_27593,N_25798,N_24590);
xnor U27594 (N_27594,N_24670,N_25293);
nand U27595 (N_27595,N_25834,N_24248);
nor U27596 (N_27596,N_25963,N_24767);
nand U27597 (N_27597,N_25050,N_25523);
nand U27598 (N_27598,N_24800,N_24494);
nand U27599 (N_27599,N_24196,N_24172);
and U27600 (N_27600,N_25202,N_25019);
and U27601 (N_27601,N_25172,N_25038);
and U27602 (N_27602,N_25305,N_24534);
nor U27603 (N_27603,N_25852,N_24820);
nor U27604 (N_27604,N_25854,N_25039);
xnor U27605 (N_27605,N_24327,N_25049);
and U27606 (N_27606,N_25989,N_25962);
nand U27607 (N_27607,N_24278,N_25524);
and U27608 (N_27608,N_25452,N_24546);
or U27609 (N_27609,N_25299,N_24589);
nand U27610 (N_27610,N_24628,N_25551);
nor U27611 (N_27611,N_24662,N_25180);
or U27612 (N_27612,N_24974,N_25947);
nor U27613 (N_27613,N_24484,N_24849);
nor U27614 (N_27614,N_25491,N_25197);
xor U27615 (N_27615,N_25608,N_24658);
nand U27616 (N_27616,N_24521,N_24642);
nand U27617 (N_27617,N_25892,N_24776);
nand U27618 (N_27618,N_25911,N_24562);
or U27619 (N_27619,N_25918,N_24182);
and U27620 (N_27620,N_25616,N_24107);
or U27621 (N_27621,N_24072,N_24753);
xnor U27622 (N_27622,N_25202,N_24684);
nor U27623 (N_27623,N_25156,N_25747);
or U27624 (N_27624,N_25058,N_25096);
or U27625 (N_27625,N_24917,N_25720);
nor U27626 (N_27626,N_24428,N_25904);
or U27627 (N_27627,N_24849,N_25618);
or U27628 (N_27628,N_25596,N_24597);
nor U27629 (N_27629,N_24985,N_25527);
and U27630 (N_27630,N_25902,N_24693);
xnor U27631 (N_27631,N_24469,N_24550);
xor U27632 (N_27632,N_25826,N_24438);
nor U27633 (N_27633,N_25799,N_24231);
or U27634 (N_27634,N_25142,N_24004);
nand U27635 (N_27635,N_25922,N_24431);
nor U27636 (N_27636,N_24071,N_25491);
nand U27637 (N_27637,N_25035,N_25041);
nand U27638 (N_27638,N_24015,N_25188);
or U27639 (N_27639,N_25107,N_24331);
nor U27640 (N_27640,N_25766,N_24096);
nor U27641 (N_27641,N_25356,N_25211);
nor U27642 (N_27642,N_24665,N_24064);
nand U27643 (N_27643,N_25074,N_25351);
nor U27644 (N_27644,N_24520,N_24047);
and U27645 (N_27645,N_25108,N_24318);
nand U27646 (N_27646,N_25088,N_24929);
or U27647 (N_27647,N_24286,N_25228);
and U27648 (N_27648,N_24235,N_24102);
xnor U27649 (N_27649,N_25200,N_24994);
nor U27650 (N_27650,N_24837,N_24834);
nand U27651 (N_27651,N_25758,N_24104);
nand U27652 (N_27652,N_24355,N_25233);
and U27653 (N_27653,N_25017,N_25550);
nor U27654 (N_27654,N_25038,N_24886);
nand U27655 (N_27655,N_25415,N_25309);
xnor U27656 (N_27656,N_24777,N_25386);
nand U27657 (N_27657,N_24710,N_25847);
or U27658 (N_27658,N_24851,N_24634);
nand U27659 (N_27659,N_25302,N_25857);
xor U27660 (N_27660,N_25428,N_24487);
or U27661 (N_27661,N_25754,N_25681);
xor U27662 (N_27662,N_25787,N_24012);
nor U27663 (N_27663,N_25598,N_24786);
and U27664 (N_27664,N_24452,N_24608);
nand U27665 (N_27665,N_24543,N_25563);
or U27666 (N_27666,N_24790,N_25244);
nor U27667 (N_27667,N_24416,N_24596);
and U27668 (N_27668,N_24275,N_25442);
or U27669 (N_27669,N_25736,N_25669);
xnor U27670 (N_27670,N_24838,N_24573);
and U27671 (N_27671,N_25106,N_24068);
xnor U27672 (N_27672,N_25758,N_24684);
and U27673 (N_27673,N_25531,N_25413);
xnor U27674 (N_27674,N_24005,N_25204);
nor U27675 (N_27675,N_25544,N_25821);
or U27676 (N_27676,N_24935,N_24534);
and U27677 (N_27677,N_24047,N_25964);
and U27678 (N_27678,N_25452,N_24015);
xnor U27679 (N_27679,N_24411,N_24047);
or U27680 (N_27680,N_25695,N_24460);
xor U27681 (N_27681,N_25390,N_25590);
xor U27682 (N_27682,N_25279,N_24104);
xor U27683 (N_27683,N_24457,N_24408);
or U27684 (N_27684,N_24944,N_24916);
and U27685 (N_27685,N_24887,N_24021);
and U27686 (N_27686,N_24296,N_24267);
nand U27687 (N_27687,N_24467,N_24853);
and U27688 (N_27688,N_25129,N_24919);
nor U27689 (N_27689,N_24002,N_24003);
nor U27690 (N_27690,N_25368,N_25953);
nand U27691 (N_27691,N_24435,N_25173);
or U27692 (N_27692,N_25281,N_25545);
nor U27693 (N_27693,N_24592,N_24415);
nor U27694 (N_27694,N_24513,N_25252);
nor U27695 (N_27695,N_24652,N_25128);
and U27696 (N_27696,N_24264,N_24717);
or U27697 (N_27697,N_25080,N_25690);
nand U27698 (N_27698,N_24120,N_25489);
nor U27699 (N_27699,N_24596,N_24084);
nand U27700 (N_27700,N_24672,N_24799);
nor U27701 (N_27701,N_25181,N_25491);
nand U27702 (N_27702,N_25368,N_24707);
or U27703 (N_27703,N_24109,N_25093);
nand U27704 (N_27704,N_25481,N_24654);
nand U27705 (N_27705,N_24468,N_24551);
nor U27706 (N_27706,N_24154,N_24622);
or U27707 (N_27707,N_25434,N_25223);
xor U27708 (N_27708,N_25655,N_24716);
nor U27709 (N_27709,N_25648,N_24100);
xor U27710 (N_27710,N_24606,N_24027);
xnor U27711 (N_27711,N_25468,N_25394);
nor U27712 (N_27712,N_24028,N_24084);
nor U27713 (N_27713,N_24887,N_24536);
or U27714 (N_27714,N_24690,N_25123);
and U27715 (N_27715,N_24805,N_24882);
and U27716 (N_27716,N_25266,N_24069);
nor U27717 (N_27717,N_24145,N_25246);
nand U27718 (N_27718,N_25061,N_25425);
nand U27719 (N_27719,N_24097,N_24125);
xnor U27720 (N_27720,N_24948,N_25886);
xor U27721 (N_27721,N_25075,N_24112);
and U27722 (N_27722,N_25403,N_24804);
xor U27723 (N_27723,N_25215,N_24610);
xnor U27724 (N_27724,N_24507,N_25144);
and U27725 (N_27725,N_24031,N_24733);
nand U27726 (N_27726,N_24253,N_25717);
and U27727 (N_27727,N_24769,N_24137);
nor U27728 (N_27728,N_24673,N_24360);
xnor U27729 (N_27729,N_25550,N_25542);
or U27730 (N_27730,N_24018,N_24988);
or U27731 (N_27731,N_25851,N_24766);
xor U27732 (N_27732,N_24129,N_25657);
nor U27733 (N_27733,N_25346,N_25133);
and U27734 (N_27734,N_24198,N_25637);
nor U27735 (N_27735,N_25644,N_24085);
and U27736 (N_27736,N_24685,N_24177);
nor U27737 (N_27737,N_24370,N_25035);
nand U27738 (N_27738,N_24133,N_25650);
nand U27739 (N_27739,N_25737,N_25822);
nor U27740 (N_27740,N_24685,N_25809);
xnor U27741 (N_27741,N_25592,N_25050);
nor U27742 (N_27742,N_24969,N_25314);
xor U27743 (N_27743,N_25740,N_25363);
nand U27744 (N_27744,N_24951,N_24594);
xor U27745 (N_27745,N_24012,N_24291);
or U27746 (N_27746,N_25352,N_24167);
xnor U27747 (N_27747,N_25383,N_25446);
or U27748 (N_27748,N_25496,N_25346);
and U27749 (N_27749,N_25745,N_24028);
or U27750 (N_27750,N_25951,N_24331);
nand U27751 (N_27751,N_25144,N_24875);
nor U27752 (N_27752,N_24097,N_25713);
xnor U27753 (N_27753,N_24575,N_24911);
nor U27754 (N_27754,N_25964,N_25328);
xnor U27755 (N_27755,N_25934,N_25217);
or U27756 (N_27756,N_25951,N_25384);
and U27757 (N_27757,N_25406,N_25341);
xnor U27758 (N_27758,N_24580,N_24498);
or U27759 (N_27759,N_24399,N_25555);
or U27760 (N_27760,N_24646,N_24665);
or U27761 (N_27761,N_25261,N_25960);
xnor U27762 (N_27762,N_25301,N_24990);
and U27763 (N_27763,N_25794,N_24073);
xor U27764 (N_27764,N_25816,N_24236);
nor U27765 (N_27765,N_24644,N_24244);
or U27766 (N_27766,N_24283,N_24254);
nor U27767 (N_27767,N_24771,N_25614);
nand U27768 (N_27768,N_24105,N_25999);
nand U27769 (N_27769,N_24378,N_24359);
xnor U27770 (N_27770,N_24269,N_24178);
and U27771 (N_27771,N_24523,N_24195);
xnor U27772 (N_27772,N_25827,N_24542);
or U27773 (N_27773,N_24340,N_25774);
nand U27774 (N_27774,N_24093,N_24003);
and U27775 (N_27775,N_25224,N_24499);
nor U27776 (N_27776,N_25015,N_25031);
nor U27777 (N_27777,N_24909,N_24412);
and U27778 (N_27778,N_25377,N_24345);
nor U27779 (N_27779,N_24058,N_25058);
nand U27780 (N_27780,N_25994,N_25104);
xnor U27781 (N_27781,N_24058,N_25850);
xor U27782 (N_27782,N_25732,N_25505);
or U27783 (N_27783,N_24837,N_25638);
xor U27784 (N_27784,N_24540,N_24245);
nor U27785 (N_27785,N_25105,N_25948);
nor U27786 (N_27786,N_25943,N_24801);
and U27787 (N_27787,N_25812,N_24260);
and U27788 (N_27788,N_24764,N_25521);
and U27789 (N_27789,N_24780,N_24599);
nand U27790 (N_27790,N_25762,N_24698);
nor U27791 (N_27791,N_24303,N_25566);
nor U27792 (N_27792,N_25259,N_25758);
or U27793 (N_27793,N_24789,N_25133);
nand U27794 (N_27794,N_24369,N_24760);
nor U27795 (N_27795,N_25327,N_24409);
or U27796 (N_27796,N_24378,N_24068);
xor U27797 (N_27797,N_25499,N_24276);
or U27798 (N_27798,N_24124,N_24374);
nor U27799 (N_27799,N_25204,N_25562);
and U27800 (N_27800,N_24947,N_24461);
xor U27801 (N_27801,N_25361,N_24725);
or U27802 (N_27802,N_24005,N_24248);
or U27803 (N_27803,N_25133,N_25124);
nor U27804 (N_27804,N_24876,N_24091);
nand U27805 (N_27805,N_25360,N_24021);
nand U27806 (N_27806,N_25187,N_25393);
xnor U27807 (N_27807,N_24643,N_25381);
and U27808 (N_27808,N_25350,N_24635);
xor U27809 (N_27809,N_25889,N_25273);
xor U27810 (N_27810,N_24925,N_24318);
nand U27811 (N_27811,N_25737,N_24747);
and U27812 (N_27812,N_24720,N_25220);
nand U27813 (N_27813,N_25734,N_25504);
xnor U27814 (N_27814,N_25262,N_25238);
xnor U27815 (N_27815,N_24513,N_24006);
or U27816 (N_27816,N_25170,N_25980);
nor U27817 (N_27817,N_25525,N_24545);
or U27818 (N_27818,N_25081,N_24427);
nand U27819 (N_27819,N_24553,N_24231);
or U27820 (N_27820,N_24000,N_24629);
or U27821 (N_27821,N_25746,N_24777);
or U27822 (N_27822,N_25331,N_24155);
xor U27823 (N_27823,N_25722,N_24342);
xnor U27824 (N_27824,N_24220,N_24578);
and U27825 (N_27825,N_24392,N_25661);
and U27826 (N_27826,N_25063,N_24906);
or U27827 (N_27827,N_25317,N_24954);
nand U27828 (N_27828,N_24213,N_25276);
or U27829 (N_27829,N_24684,N_25153);
or U27830 (N_27830,N_25177,N_25416);
or U27831 (N_27831,N_25255,N_25574);
and U27832 (N_27832,N_24252,N_24646);
and U27833 (N_27833,N_25504,N_25937);
nand U27834 (N_27834,N_24367,N_25777);
xnor U27835 (N_27835,N_24296,N_25457);
and U27836 (N_27836,N_24663,N_25578);
xnor U27837 (N_27837,N_24610,N_24011);
or U27838 (N_27838,N_24215,N_24477);
nor U27839 (N_27839,N_24836,N_25398);
or U27840 (N_27840,N_25744,N_24022);
and U27841 (N_27841,N_25893,N_25237);
nor U27842 (N_27842,N_25220,N_24144);
nor U27843 (N_27843,N_25004,N_25384);
or U27844 (N_27844,N_24566,N_24444);
nand U27845 (N_27845,N_25063,N_24602);
nand U27846 (N_27846,N_24151,N_25622);
or U27847 (N_27847,N_24966,N_24486);
nor U27848 (N_27848,N_24743,N_25566);
or U27849 (N_27849,N_24011,N_25578);
and U27850 (N_27850,N_24191,N_25218);
or U27851 (N_27851,N_24031,N_24602);
and U27852 (N_27852,N_25031,N_24385);
and U27853 (N_27853,N_25131,N_25299);
and U27854 (N_27854,N_25456,N_25384);
or U27855 (N_27855,N_24935,N_25225);
or U27856 (N_27856,N_25100,N_24184);
xnor U27857 (N_27857,N_25057,N_24189);
and U27858 (N_27858,N_25182,N_24300);
nand U27859 (N_27859,N_25676,N_24976);
xnor U27860 (N_27860,N_25518,N_24543);
nand U27861 (N_27861,N_25790,N_25131);
nand U27862 (N_27862,N_25844,N_25107);
or U27863 (N_27863,N_24796,N_24819);
or U27864 (N_27864,N_25202,N_25513);
or U27865 (N_27865,N_25757,N_24118);
nand U27866 (N_27866,N_24043,N_25828);
or U27867 (N_27867,N_25957,N_25178);
and U27868 (N_27868,N_24750,N_25230);
and U27869 (N_27869,N_24772,N_25715);
xor U27870 (N_27870,N_24053,N_24872);
and U27871 (N_27871,N_24569,N_24691);
or U27872 (N_27872,N_25955,N_24195);
nand U27873 (N_27873,N_25927,N_25030);
xnor U27874 (N_27874,N_24360,N_25529);
xor U27875 (N_27875,N_25150,N_24634);
nor U27876 (N_27876,N_24397,N_24240);
nor U27877 (N_27877,N_24053,N_25235);
xor U27878 (N_27878,N_25946,N_25954);
or U27879 (N_27879,N_25235,N_25696);
nand U27880 (N_27880,N_25453,N_24066);
nor U27881 (N_27881,N_24526,N_25564);
or U27882 (N_27882,N_24948,N_24199);
xor U27883 (N_27883,N_25201,N_24906);
nor U27884 (N_27884,N_25840,N_24873);
and U27885 (N_27885,N_25609,N_25282);
nor U27886 (N_27886,N_25492,N_24745);
nand U27887 (N_27887,N_25589,N_24273);
nor U27888 (N_27888,N_24726,N_24371);
nor U27889 (N_27889,N_24640,N_24316);
nor U27890 (N_27890,N_25759,N_25429);
nor U27891 (N_27891,N_24787,N_25901);
and U27892 (N_27892,N_25743,N_24070);
or U27893 (N_27893,N_25948,N_25067);
nor U27894 (N_27894,N_24930,N_24888);
nand U27895 (N_27895,N_24604,N_25737);
or U27896 (N_27896,N_25119,N_25362);
xor U27897 (N_27897,N_24973,N_25256);
nand U27898 (N_27898,N_25250,N_24008);
or U27899 (N_27899,N_24032,N_25119);
nor U27900 (N_27900,N_25192,N_25402);
or U27901 (N_27901,N_25117,N_25403);
nor U27902 (N_27902,N_24767,N_24761);
nand U27903 (N_27903,N_25184,N_25669);
or U27904 (N_27904,N_25434,N_25505);
xnor U27905 (N_27905,N_24967,N_24932);
or U27906 (N_27906,N_25070,N_24599);
nor U27907 (N_27907,N_25000,N_25240);
and U27908 (N_27908,N_25827,N_24747);
and U27909 (N_27909,N_24460,N_24492);
xor U27910 (N_27910,N_24612,N_24344);
or U27911 (N_27911,N_24761,N_25193);
nand U27912 (N_27912,N_25021,N_24961);
and U27913 (N_27913,N_25835,N_24475);
xor U27914 (N_27914,N_24758,N_25334);
and U27915 (N_27915,N_25781,N_24040);
or U27916 (N_27916,N_25610,N_24823);
nand U27917 (N_27917,N_25839,N_25581);
or U27918 (N_27918,N_25009,N_25926);
and U27919 (N_27919,N_24131,N_25619);
nand U27920 (N_27920,N_24371,N_25696);
nand U27921 (N_27921,N_24187,N_24532);
and U27922 (N_27922,N_25235,N_24448);
nor U27923 (N_27923,N_24397,N_25652);
and U27924 (N_27924,N_25378,N_25596);
or U27925 (N_27925,N_24357,N_25650);
or U27926 (N_27926,N_25222,N_25976);
nor U27927 (N_27927,N_24519,N_25686);
nand U27928 (N_27928,N_24324,N_25390);
xnor U27929 (N_27929,N_25763,N_24039);
xor U27930 (N_27930,N_24605,N_24054);
xnor U27931 (N_27931,N_25129,N_24693);
nand U27932 (N_27932,N_25340,N_24712);
nand U27933 (N_27933,N_25020,N_24137);
and U27934 (N_27934,N_25237,N_25467);
or U27935 (N_27935,N_25769,N_24580);
and U27936 (N_27936,N_24101,N_25349);
or U27937 (N_27937,N_24133,N_24681);
nand U27938 (N_27938,N_24084,N_25896);
xnor U27939 (N_27939,N_25936,N_24551);
and U27940 (N_27940,N_24840,N_24715);
or U27941 (N_27941,N_25851,N_24672);
xnor U27942 (N_27942,N_25569,N_25913);
and U27943 (N_27943,N_25896,N_24846);
or U27944 (N_27944,N_24867,N_25580);
xnor U27945 (N_27945,N_25556,N_24288);
xnor U27946 (N_27946,N_24414,N_24984);
nor U27947 (N_27947,N_24292,N_25540);
and U27948 (N_27948,N_24821,N_24665);
and U27949 (N_27949,N_24864,N_25331);
nor U27950 (N_27950,N_25901,N_25840);
or U27951 (N_27951,N_24586,N_25548);
nor U27952 (N_27952,N_25230,N_24464);
nand U27953 (N_27953,N_25307,N_25627);
xnor U27954 (N_27954,N_24858,N_24662);
or U27955 (N_27955,N_25075,N_25767);
and U27956 (N_27956,N_24092,N_24106);
and U27957 (N_27957,N_25560,N_24808);
and U27958 (N_27958,N_25953,N_25318);
nor U27959 (N_27959,N_25815,N_25000);
nand U27960 (N_27960,N_24905,N_25476);
or U27961 (N_27961,N_24577,N_24157);
and U27962 (N_27962,N_24453,N_25877);
or U27963 (N_27963,N_24514,N_24574);
nor U27964 (N_27964,N_25889,N_24459);
nor U27965 (N_27965,N_25805,N_24298);
nand U27966 (N_27966,N_25717,N_24583);
or U27967 (N_27967,N_25045,N_25521);
and U27968 (N_27968,N_24370,N_25007);
nand U27969 (N_27969,N_25315,N_25988);
and U27970 (N_27970,N_25887,N_24677);
and U27971 (N_27971,N_24786,N_24063);
and U27972 (N_27972,N_24199,N_24619);
and U27973 (N_27973,N_25523,N_24395);
or U27974 (N_27974,N_24481,N_24764);
xnor U27975 (N_27975,N_25028,N_25413);
and U27976 (N_27976,N_25039,N_25682);
nor U27977 (N_27977,N_24069,N_24195);
nand U27978 (N_27978,N_25560,N_24824);
nor U27979 (N_27979,N_24808,N_25666);
xnor U27980 (N_27980,N_24885,N_24394);
nor U27981 (N_27981,N_25747,N_24209);
and U27982 (N_27982,N_25728,N_25162);
nor U27983 (N_27983,N_24002,N_25325);
xnor U27984 (N_27984,N_25255,N_24936);
nor U27985 (N_27985,N_24295,N_25578);
xor U27986 (N_27986,N_24196,N_24089);
xnor U27987 (N_27987,N_25357,N_24074);
nor U27988 (N_27988,N_24161,N_24852);
and U27989 (N_27989,N_25204,N_24895);
xor U27990 (N_27990,N_24129,N_25545);
nand U27991 (N_27991,N_24470,N_24886);
xor U27992 (N_27992,N_24150,N_24508);
xor U27993 (N_27993,N_24978,N_24043);
nor U27994 (N_27994,N_25135,N_25918);
nor U27995 (N_27995,N_24073,N_24947);
or U27996 (N_27996,N_24408,N_25946);
and U27997 (N_27997,N_24394,N_25476);
xor U27998 (N_27998,N_25351,N_25517);
xnor U27999 (N_27999,N_24265,N_25912);
nor U28000 (N_28000,N_26716,N_26322);
nand U28001 (N_28001,N_26890,N_27058);
or U28002 (N_28002,N_27625,N_27849);
nor U28003 (N_28003,N_27372,N_26630);
or U28004 (N_28004,N_26966,N_26458);
and U28005 (N_28005,N_27801,N_26598);
nand U28006 (N_28006,N_26617,N_27867);
or U28007 (N_28007,N_27773,N_27127);
or U28008 (N_28008,N_26806,N_26596);
xor U28009 (N_28009,N_27772,N_27906);
and U28010 (N_28010,N_27959,N_27286);
and U28011 (N_28011,N_27542,N_27548);
or U28012 (N_28012,N_27438,N_26225);
and U28013 (N_28013,N_26505,N_27236);
nand U28014 (N_28014,N_26571,N_27211);
xnor U28015 (N_28015,N_26165,N_26488);
nand U28016 (N_28016,N_27272,N_27770);
xnor U28017 (N_28017,N_26888,N_26507);
or U28018 (N_28018,N_27683,N_26320);
nor U28019 (N_28019,N_27055,N_26096);
nor U28020 (N_28020,N_26411,N_26574);
xnor U28021 (N_28021,N_26293,N_26399);
or U28022 (N_28022,N_26764,N_27454);
nor U28023 (N_28023,N_27147,N_27176);
nand U28024 (N_28024,N_27866,N_27191);
or U28025 (N_28025,N_26438,N_26331);
xnor U28026 (N_28026,N_27513,N_27616);
nand U28027 (N_28027,N_27148,N_26634);
and U28028 (N_28028,N_26498,N_26773);
and U28029 (N_28029,N_27208,N_26242);
xnor U28030 (N_28030,N_27641,N_26703);
or U28031 (N_28031,N_27075,N_27786);
and U28032 (N_28032,N_26779,N_27314);
xnor U28033 (N_28033,N_26661,N_27134);
nor U28034 (N_28034,N_26190,N_27675);
and U28035 (N_28035,N_27511,N_26025);
nand U28036 (N_28036,N_27806,N_27120);
xor U28037 (N_28037,N_26277,N_27471);
or U28038 (N_28038,N_26052,N_27455);
nor U28039 (N_28039,N_26284,N_27682);
xnor U28040 (N_28040,N_27881,N_26099);
nand U28041 (N_28041,N_26317,N_26881);
xnor U28042 (N_28042,N_27718,N_27585);
nand U28043 (N_28043,N_27941,N_27026);
and U28044 (N_28044,N_27578,N_26326);
or U28045 (N_28045,N_26927,N_27606);
and U28046 (N_28046,N_27823,N_26971);
and U28047 (N_28047,N_26163,N_27348);
nand U28048 (N_28048,N_27168,N_27267);
and U28049 (N_28049,N_27684,N_27488);
nor U28050 (N_28050,N_26704,N_27430);
or U28051 (N_28051,N_26552,N_26409);
xor U28052 (N_28052,N_27185,N_26583);
nor U28053 (N_28053,N_27240,N_27069);
nand U28054 (N_28054,N_27978,N_27672);
nand U28055 (N_28055,N_26378,N_27186);
nand U28056 (N_28056,N_27593,N_26524);
xnor U28057 (N_28057,N_27986,N_26270);
nand U28058 (N_28058,N_27564,N_26041);
nand U28059 (N_28059,N_26914,N_27184);
xor U28060 (N_28060,N_26218,N_26919);
nor U28061 (N_28061,N_26297,N_27189);
or U28062 (N_28062,N_26417,N_27251);
xnor U28063 (N_28063,N_26369,N_26875);
nor U28064 (N_28064,N_27465,N_27802);
nor U28065 (N_28065,N_26291,N_26368);
or U28066 (N_28066,N_26726,N_27627);
and U28067 (N_28067,N_27632,N_27311);
and U28068 (N_28068,N_26090,N_27595);
or U28069 (N_28069,N_27618,N_27373);
or U28070 (N_28070,N_26037,N_26950);
xor U28071 (N_28071,N_26472,N_26846);
nor U28072 (N_28072,N_27633,N_27164);
or U28073 (N_28073,N_27581,N_27889);
nand U28074 (N_28074,N_26449,N_27829);
or U28075 (N_28075,N_27762,N_26861);
nor U28076 (N_28076,N_27729,N_26354);
nand U28077 (N_28077,N_26851,N_26942);
nand U28078 (N_28078,N_26850,N_26391);
xor U28079 (N_28079,N_27545,N_26053);
nor U28080 (N_28080,N_27358,N_26961);
nor U28081 (N_28081,N_27587,N_27294);
and U28082 (N_28082,N_27580,N_26016);
nor U28083 (N_28083,N_27811,N_26602);
or U28084 (N_28084,N_27025,N_27153);
xor U28085 (N_28085,N_27111,N_26975);
and U28086 (N_28086,N_26511,N_27064);
nand U28087 (N_28087,N_26601,N_27139);
or U28088 (N_28088,N_26509,N_27766);
or U28089 (N_28089,N_27397,N_26652);
nor U28090 (N_28090,N_27951,N_26822);
nor U28091 (N_28091,N_27239,N_27601);
or U28092 (N_28092,N_26107,N_27280);
xor U28093 (N_28093,N_26414,N_27495);
or U28094 (N_28094,N_26710,N_26976);
nor U28095 (N_28095,N_27349,N_26852);
or U28096 (N_28096,N_26227,N_27426);
nor U28097 (N_28097,N_27434,N_27491);
or U28098 (N_28098,N_27868,N_27083);
nand U28099 (N_28099,N_26420,N_26038);
nand U28100 (N_28100,N_27344,N_26140);
nand U28101 (N_28101,N_27494,N_26489);
xnor U28102 (N_28102,N_27370,N_26821);
nand U28103 (N_28103,N_26813,N_27099);
xnor U28104 (N_28104,N_26441,N_26097);
xor U28105 (N_28105,N_26389,N_27066);
nand U28106 (N_28106,N_26567,N_26569);
and U28107 (N_28107,N_27350,N_26913);
xor U28108 (N_28108,N_27173,N_26922);
and U28109 (N_28109,N_26694,N_27567);
xnor U28110 (N_28110,N_26578,N_26046);
and U28111 (N_28111,N_26130,N_26250);
and U28112 (N_28112,N_27318,N_27261);
xor U28113 (N_28113,N_27096,N_27553);
nor U28114 (N_28114,N_26374,N_26801);
xor U28115 (N_28115,N_26103,N_27077);
nand U28116 (N_28116,N_26945,N_26864);
or U28117 (N_28117,N_27044,N_27484);
xnor U28118 (N_28118,N_26908,N_27343);
nand U28119 (N_28119,N_26957,N_27988);
nand U28120 (N_28120,N_26595,N_27022);
and U28121 (N_28121,N_26618,N_27639);
or U28122 (N_28122,N_26471,N_27283);
xor U28123 (N_28123,N_27427,N_27338);
or U28124 (N_28124,N_26461,N_27258);
nor U28125 (N_28125,N_26358,N_26713);
nor U28126 (N_28126,N_27228,N_27737);
nand U28127 (N_28127,N_26196,N_26651);
nor U28128 (N_28128,N_26810,N_26626);
and U28129 (N_28129,N_26093,N_27420);
and U28130 (N_28130,N_26772,N_27056);
and U28131 (N_28131,N_27512,N_26030);
or U28132 (N_28132,N_27469,N_27447);
nand U28133 (N_28133,N_26874,N_26403);
xor U28134 (N_28134,N_27699,N_26905);
nor U28135 (N_28135,N_27681,N_27034);
and U28136 (N_28136,N_26363,N_27203);
and U28137 (N_28137,N_27886,N_27725);
nor U28138 (N_28138,N_27500,N_27655);
nor U28139 (N_28139,N_27615,N_27245);
or U28140 (N_28140,N_27603,N_27863);
and U28141 (N_28141,N_27741,N_27523);
xor U28142 (N_28142,N_27793,N_26055);
nor U28143 (N_28143,N_26701,N_26169);
nand U28144 (N_28144,N_26241,N_27654);
nor U28145 (N_28145,N_27411,N_27162);
or U28146 (N_28146,N_26659,N_27705);
and U28147 (N_28147,N_26148,N_26972);
or U28148 (N_28148,N_26612,N_26818);
or U28149 (N_28149,N_26337,N_27316);
xnor U28150 (N_28150,N_27144,N_27649);
nand U28151 (N_28151,N_26004,N_26167);
xnor U28152 (N_28152,N_27588,N_26156);
nand U28153 (N_28153,N_26644,N_27380);
nand U28154 (N_28154,N_27010,N_27758);
nor U28155 (N_28155,N_27453,N_27650);
xor U28156 (N_28156,N_27014,N_27932);
nor U28157 (N_28157,N_26166,N_27930);
nor U28158 (N_28158,N_26380,N_26530);
nor U28159 (N_28159,N_26677,N_27944);
xor U28160 (N_28160,N_26994,N_27417);
or U28161 (N_28161,N_26355,N_26010);
nand U28162 (N_28162,N_27233,N_27385);
or U28163 (N_28163,N_27861,N_27326);
nor U28164 (N_28164,N_27563,N_27156);
nor U28165 (N_28165,N_26514,N_27924);
and U28166 (N_28166,N_27652,N_27409);
xnor U28167 (N_28167,N_27320,N_26546);
and U28168 (N_28168,N_26269,N_26879);
xor U28169 (N_28169,N_26620,N_27755);
and U28170 (N_28170,N_27394,N_27717);
nor U28171 (N_28171,N_27333,N_26762);
xor U28172 (N_28172,N_27598,N_27323);
and U28173 (N_28173,N_26480,N_27808);
nand U28174 (N_28174,N_27329,N_26732);
or U28175 (N_28175,N_26792,N_26256);
nand U28176 (N_28176,N_27727,N_27855);
nor U28177 (N_28177,N_27017,N_26907);
or U28178 (N_28178,N_26862,N_26221);
nor U28179 (N_28179,N_27850,N_26342);
or U28180 (N_28180,N_27573,N_27676);
or U28181 (N_28181,N_26777,N_26537);
xnor U28182 (N_28182,N_26641,N_27537);
nand U28183 (N_28183,N_27442,N_26629);
and U28184 (N_28184,N_27230,N_26272);
or U28185 (N_28185,N_27334,N_27276);
nand U28186 (N_28186,N_27508,N_27118);
nand U28187 (N_28187,N_27554,N_27253);
or U28188 (N_28188,N_26512,N_27835);
and U28189 (N_28189,N_26068,N_27817);
and U28190 (N_28190,N_26171,N_27327);
and U28191 (N_28191,N_26201,N_27589);
xor U28192 (N_28192,N_26551,N_26457);
nor U28193 (N_28193,N_26521,N_26247);
xnor U28194 (N_28194,N_26903,N_27163);
and U28195 (N_28195,N_26650,N_27592);
and U28196 (N_28196,N_26717,N_27630);
xnor U28197 (N_28197,N_26889,N_27094);
xor U28198 (N_28198,N_27072,N_26559);
or U28199 (N_28199,N_26078,N_26120);
xnor U28200 (N_28200,N_27306,N_27828);
nand U28201 (N_28201,N_26199,N_27489);
xor U28202 (N_28202,N_27605,N_27460);
and U28203 (N_28203,N_27146,N_27353);
and U28204 (N_28204,N_27408,N_27112);
nor U28205 (N_28205,N_27799,N_26310);
nand U28206 (N_28206,N_27975,N_27266);
xor U28207 (N_28207,N_27635,N_26178);
nand U28208 (N_28208,N_27027,N_27486);
and U28209 (N_28209,N_27923,N_27966);
xnor U28210 (N_28210,N_27254,N_26083);
nor U28211 (N_28211,N_27621,N_26588);
xnor U28212 (N_28212,N_26614,N_27840);
xor U28213 (N_28213,N_27694,N_27088);
xnor U28214 (N_28214,N_26820,N_27328);
nand U28215 (N_28215,N_27401,N_27858);
xor U28216 (N_28216,N_26314,N_27535);
xor U28217 (N_28217,N_26315,N_27352);
or U28218 (N_28218,N_27207,N_27070);
and U28219 (N_28219,N_27956,N_27872);
nor U28220 (N_28220,N_26640,N_27960);
nand U28221 (N_28221,N_26406,N_26878);
nor U28222 (N_28222,N_26579,N_26695);
and U28223 (N_28223,N_26676,N_27935);
xor U28224 (N_28224,N_27238,N_27541);
nor U28225 (N_28225,N_26566,N_27857);
xnor U28226 (N_28226,N_26575,N_26767);
or U28227 (N_28227,N_27085,N_27478);
nand U28228 (N_28228,N_27883,N_27464);
and U28229 (N_28229,N_26295,N_26476);
and U28230 (N_28230,N_26607,N_27730);
and U28231 (N_28231,N_27955,N_26024);
or U28232 (N_28232,N_26141,N_27183);
or U28233 (N_28233,N_26536,N_26527);
xnor U28234 (N_28234,N_27325,N_26510);
nand U28235 (N_28235,N_26137,N_27086);
and U28236 (N_28236,N_26970,N_27476);
nor U28237 (N_28237,N_26371,N_26868);
nor U28238 (N_28238,N_26439,N_27629);
nand U28239 (N_28239,N_27876,N_27499);
or U28240 (N_28240,N_27778,N_27984);
xnor U28241 (N_28241,N_27104,N_27706);
and U28242 (N_28242,N_26381,N_26817);
nand U28243 (N_28243,N_26664,N_27378);
nor U28244 (N_28244,N_26238,N_27043);
or U28245 (N_28245,N_26871,N_27670);
or U28246 (N_28246,N_27403,N_26340);
and U28247 (N_28247,N_27151,N_26430);
or U28248 (N_28248,N_26036,N_27748);
xnor U28249 (N_28249,N_26958,N_26398);
nand U28250 (N_28250,N_26249,N_26056);
xor U28251 (N_28251,N_27519,N_27768);
nand U28252 (N_28252,N_27971,N_26947);
nand U28253 (N_28253,N_26145,N_27040);
and U28254 (N_28254,N_26553,N_26134);
nand U28255 (N_28255,N_27902,N_26361);
nand U28256 (N_28256,N_26386,N_27747);
and U28257 (N_28257,N_26487,N_27792);
and U28258 (N_28258,N_26836,N_26799);
nor U28259 (N_28259,N_27375,N_27475);
nor U28260 (N_28260,N_27662,N_27011);
or U28261 (N_28261,N_27561,N_26518);
nand U28262 (N_28262,N_27695,N_26916);
and U28263 (N_28263,N_26076,N_27636);
nor U28264 (N_28264,N_26302,N_27062);
or U28265 (N_28265,N_26485,N_27733);
or U28266 (N_28266,N_26265,N_26832);
and U28267 (N_28267,N_27371,N_26177);
or U28268 (N_28268,N_26312,N_27550);
and U28269 (N_28269,N_27594,N_27451);
and U28270 (N_28270,N_27379,N_26721);
nor U28271 (N_28271,N_26666,N_26203);
and U28272 (N_28272,N_27692,N_27666);
and U28273 (N_28273,N_26711,N_26727);
nand U28274 (N_28274,N_27340,N_27903);
nor U28275 (N_28275,N_26720,N_26435);
xor U28276 (N_28276,N_27260,N_26637);
nor U28277 (N_28277,N_26548,N_26131);
or U28278 (N_28278,N_26188,N_27977);
or U28279 (N_28279,N_27999,N_26775);
or U28280 (N_28280,N_26741,N_27090);
nand U28281 (N_28281,N_26503,N_26978);
and U28282 (N_28282,N_27078,N_27160);
xor U28283 (N_28283,N_26197,N_27698);
or U28284 (N_28284,N_26979,N_27399);
or U28285 (N_28285,N_27376,N_26660);
xnor U28286 (N_28286,N_27387,N_26572);
nand U28287 (N_28287,N_27171,N_26969);
nand U28288 (N_28288,N_27031,N_27949);
nand U28289 (N_28289,N_26054,N_26885);
and U28290 (N_28290,N_27783,N_27982);
nand U28291 (N_28291,N_27067,N_26086);
nand U28292 (N_28292,N_26364,N_26747);
nor U28293 (N_28293,N_27958,N_27538);
nor U28294 (N_28294,N_26653,N_27877);
xor U28295 (N_28295,N_27215,N_26211);
or U28296 (N_28296,N_27507,N_27967);
and U28297 (N_28297,N_27771,N_26467);
or U28298 (N_28298,N_26463,N_27012);
or U28299 (N_28299,N_27405,N_27888);
or U28300 (N_28300,N_27925,N_27800);
and U28301 (N_28301,N_27287,N_27223);
and U28302 (N_28302,N_27421,N_26622);
or U28303 (N_28303,N_27838,N_27911);
or U28304 (N_28304,N_26985,N_27292);
xor U28305 (N_28305,N_27987,N_26195);
and U28306 (N_28306,N_26639,N_26847);
nand U28307 (N_28307,N_26800,N_26251);
nand U28308 (N_28308,N_26491,N_26643);
xnor U28309 (N_28309,N_27165,N_27624);
nand U28310 (N_28310,N_26765,N_27243);
nand U28311 (N_28311,N_26421,N_27103);
xor U28312 (N_28312,N_27887,N_27049);
xnor U28313 (N_28313,N_26980,N_26845);
or U28314 (N_28314,N_27824,N_26700);
xnor U28315 (N_28315,N_27305,N_26264);
nand U28316 (N_28316,N_26327,N_26949);
or U28317 (N_28317,N_26789,N_26345);
or U28318 (N_28318,N_26044,N_26606);
xor U28319 (N_28319,N_27042,N_27780);
and U28320 (N_28320,N_26252,N_27302);
or U28321 (N_28321,N_26645,N_27929);
or U28322 (N_28322,N_27119,N_26910);
nand U28323 (N_28323,N_26943,N_26873);
xor U28324 (N_28324,N_26712,N_26128);
xnor U28325 (N_28325,N_27712,N_26132);
nor U28326 (N_28326,N_27374,N_26756);
or U28327 (N_28327,N_27281,N_26045);
nor U28328 (N_28328,N_26493,N_27115);
or U28329 (N_28329,N_27710,N_26731);
xor U28330 (N_28330,N_27029,N_27347);
xor U28331 (N_28331,N_27277,N_27345);
or U28332 (N_28332,N_26589,N_26819);
nor U28333 (N_28333,N_26605,N_27051);
and U28334 (N_28334,N_26642,N_26164);
nor U28335 (N_28335,N_27407,N_26805);
and U28336 (N_28336,N_26465,N_27809);
or U28337 (N_28337,N_27954,N_27021);
or U28338 (N_28338,N_26259,N_27895);
xor U28339 (N_28339,N_27023,N_27722);
xor U28340 (N_28340,N_26469,N_27235);
and U28341 (N_28341,N_26080,N_27300);
and U28342 (N_28342,N_26347,N_27504);
or U28343 (N_28343,N_27496,N_27897);
nor U28344 (N_28344,N_26370,N_27101);
nor U28345 (N_28345,N_26603,N_26675);
or U28346 (N_28346,N_26941,N_26321);
nand U28347 (N_28347,N_27679,N_26181);
nor U28348 (N_28348,N_26307,N_26515);
and U28349 (N_28349,N_27013,N_26112);
or U28350 (N_28350,N_27413,N_26900);
and U28351 (N_28351,N_27844,N_26023);
or U28352 (N_28352,N_26740,N_26586);
nor U28353 (N_28353,N_27531,N_27576);
xnor U28354 (N_28354,N_27392,N_26582);
or U28355 (N_28355,N_26474,N_27524);
xnor U28356 (N_28356,N_26110,N_27830);
nor U28357 (N_28357,N_27610,N_27206);
or U28358 (N_28358,N_27979,N_27480);
nor U28359 (N_28359,N_27781,N_26468);
or U28360 (N_28360,N_27668,N_26904);
or U28361 (N_28361,N_26176,N_27776);
and U28362 (N_28362,N_26475,N_26754);
or U28363 (N_28363,N_26960,N_26229);
and U28364 (N_28364,N_27398,N_27452);
or U28365 (N_28365,N_26007,N_27948);
xnor U28366 (N_28366,N_27961,N_26301);
and U28367 (N_28367,N_27377,N_26212);
and U28368 (N_28368,N_26804,N_27572);
nand U28369 (N_28369,N_26988,N_27249);
nor U28370 (N_28370,N_26431,N_27321);
nor U28371 (N_28371,N_27822,N_26451);
nand U28372 (N_28372,N_27130,N_27790);
and U28373 (N_28373,N_27275,N_26982);
nor U28374 (N_28374,N_26253,N_27273);
nor U28375 (N_28375,N_27487,N_26624);
nor U28376 (N_28376,N_27634,N_27319);
and U28377 (N_28377,N_26285,N_26745);
and U28378 (N_28378,N_26547,N_27746);
nor U28379 (N_28379,N_26830,N_26434);
xor U28380 (N_28380,N_26814,N_27785);
nand U28381 (N_28381,N_27367,N_26593);
xnor U28382 (N_28382,N_27418,N_26452);
xor U28383 (N_28383,N_26022,N_27068);
xnor U28384 (N_28384,N_27509,N_27631);
nand U28385 (N_28385,N_26135,N_27059);
and U28386 (N_28386,N_26048,N_27301);
nor U28387 (N_28387,N_27751,N_27647);
nor U28388 (N_28388,N_27693,N_27004);
nor U28389 (N_28389,N_26304,N_27931);
nand U28390 (N_28390,N_27179,N_27591);
or U28391 (N_28391,N_26738,N_27315);
xnor U28392 (N_28392,N_26224,N_27231);
nand U28393 (N_28393,N_26357,N_26170);
nor U28394 (N_28394,N_27404,N_26428);
or U28395 (N_28395,N_27878,N_26194);
and U28396 (N_28396,N_26060,N_26108);
nor U28397 (N_28397,N_27938,N_27896);
nand U28398 (N_28398,N_26788,N_26244);
or U28399 (N_28399,N_26802,N_26013);
xor U28400 (N_28400,N_27845,N_27423);
nor U28401 (N_28401,N_27574,N_27514);
or U28402 (N_28402,N_27933,N_27336);
and U28403 (N_28403,N_26373,N_26394);
xor U28404 (N_28404,N_27007,N_26892);
nand U28405 (N_28405,N_27255,N_27312);
and U28406 (N_28406,N_26999,N_26808);
nor U28407 (N_28407,N_26590,N_27658);
xnor U28408 (N_28408,N_27226,N_27458);
nor U28409 (N_28409,N_27357,N_26816);
or U28410 (N_28410,N_26213,N_27142);
or U28411 (N_28411,N_27674,N_26299);
nor U28412 (N_28412,N_27020,N_27145);
xor U28413 (N_28413,N_27356,N_26860);
nand U28414 (N_28414,N_27685,N_26228);
and U28415 (N_28415,N_27310,N_27981);
xor U28416 (N_28416,N_26182,N_27920);
xor U28417 (N_28417,N_26412,N_27415);
and U28418 (N_28418,N_26027,N_26549);
and U28419 (N_28419,N_27885,N_26967);
nand U28420 (N_28420,N_27194,N_26750);
and U28421 (N_28421,N_27530,N_26499);
xnor U28422 (N_28422,N_26619,N_26993);
or U28423 (N_28423,N_26944,N_26884);
nor U28424 (N_28424,N_26125,N_27082);
nand U28425 (N_28425,N_27091,N_26334);
or U28426 (N_28426,N_27282,N_26419);
xnor U28427 (N_28427,N_26183,N_26723);
or U28428 (N_28428,N_26555,N_26372);
xor U28429 (N_28429,N_26952,N_26193);
xnor U28430 (N_28430,N_27993,N_27623);
or U28431 (N_28431,N_26996,N_27432);
and U28432 (N_28432,N_26191,N_27506);
and U28433 (N_28433,N_26094,N_27937);
nand U28434 (N_28434,N_27905,N_26989);
or U28435 (N_28435,N_27539,N_26150);
and U28436 (N_28436,N_27490,N_27225);
nand U28437 (N_28437,N_27178,N_26008);
nor U28438 (N_28438,N_27536,N_27291);
xnor U28439 (N_28439,N_27973,N_27308);
nand U28440 (N_28440,N_26275,N_26787);
and U28441 (N_28441,N_27980,N_27284);
and U28442 (N_28442,N_26206,N_26689);
or U28443 (N_28443,N_26233,N_27199);
nand U28444 (N_28444,N_27969,N_27175);
and U28445 (N_28445,N_26351,N_27743);
nor U28446 (N_28446,N_27383,N_26184);
and U28447 (N_28447,N_27113,N_27678);
or U28448 (N_28448,N_26387,N_27503);
and U28449 (N_28449,N_26833,N_26826);
xor U28450 (N_28450,N_26311,N_26872);
xor U28451 (N_28451,N_27669,N_27522);
nand U28452 (N_28452,N_26562,N_26823);
nand U28453 (N_28453,N_26162,N_27934);
or U28454 (N_28454,N_26724,N_26113);
nor U28455 (N_28455,N_27568,N_26216);
or U28456 (N_28456,N_26939,N_27181);
nand U28457 (N_28457,N_26730,N_26180);
and U28458 (N_28458,N_27213,N_27818);
or U28459 (N_28459,N_27540,N_26636);
xor U28460 (N_28460,N_27721,N_27299);
or U28461 (N_28461,N_27293,N_26528);
and U28462 (N_28462,N_26353,N_26283);
or U28463 (N_28463,N_27219,N_27505);
xor U28464 (N_28464,N_26848,N_26974);
nand U28465 (N_28465,N_26274,N_27138);
nor U28466 (N_28466,N_26159,N_26743);
nor U28467 (N_28467,N_26114,N_26621);
nor U28468 (N_28468,N_26714,N_26172);
nor U28469 (N_28469,N_27424,N_26494);
and U28470 (N_28470,N_27856,N_26139);
nand U28471 (N_28471,N_26576,N_26674);
or U28472 (N_28472,N_26858,N_26425);
nand U28473 (N_28473,N_27346,N_26043);
nor U28474 (N_28474,N_26123,N_26550);
nand U28475 (N_28475,N_27149,N_27673);
nand U28476 (N_28476,N_26867,N_26525);
or U28477 (N_28477,N_27141,N_27073);
xnor U28478 (N_28478,N_27677,N_27355);
xor U28479 (N_28479,N_27117,N_26174);
nor U28480 (N_28480,N_26759,N_26077);
xnor U28481 (N_28481,N_26392,N_27363);
and U28482 (N_28482,N_26794,N_27812);
xnor U28483 (N_28483,N_26091,N_26028);
nor U28484 (N_28484,N_27874,N_27779);
nand U28485 (N_28485,N_26279,N_27656);
xnor U28486 (N_28486,N_27614,N_26897);
or U28487 (N_28487,N_26124,N_27110);
and U28488 (N_28488,N_26443,N_26936);
xnor U28489 (N_28489,N_27202,N_26896);
nand U28490 (N_28490,N_27767,N_27754);
nor U28491 (N_28491,N_26835,N_26121);
xnor U28492 (N_28492,N_27076,N_26854);
nor U28493 (N_28493,N_27739,N_26210);
or U28494 (N_28494,N_27671,N_27834);
and U28495 (N_28495,N_26255,N_26151);
or U28496 (N_28496,N_27661,N_26360);
and U28497 (N_28497,N_26529,N_27093);
or U28498 (N_28498,N_27234,N_27192);
xnor U28499 (N_28499,N_26445,N_27241);
xor U28500 (N_28500,N_27763,N_26179);
nand U28501 (N_28501,N_26440,N_27789);
xor U28502 (N_28502,N_26516,N_27557);
xor U28503 (N_28503,N_26869,N_26519);
nand U28504 (N_28504,N_27498,N_26116);
or U28505 (N_28505,N_27229,N_26407);
nand U28506 (N_28506,N_26992,N_27998);
nand U28507 (N_28507,N_27008,N_27726);
nand U28508 (N_28508,N_27342,N_26230);
xor U28509 (N_28509,N_27259,N_26019);
nor U28510 (N_28510,N_26938,N_27483);
nor U28511 (N_28511,N_26069,N_26073);
or U28512 (N_28512,N_26753,N_26332);
nand U28513 (N_28513,N_26880,N_26433);
and U28514 (N_28514,N_26349,N_26654);
and U28515 (N_28515,N_27382,N_26672);
and U28516 (N_28516,N_26234,N_26774);
nor U28517 (N_28517,N_26065,N_26681);
and U28518 (N_28518,N_26838,N_27892);
nor U28519 (N_28519,N_27989,N_26613);
or U28520 (N_28520,N_27190,N_26138);
nor U28521 (N_28521,N_26563,N_27893);
or U28522 (N_28522,N_27821,N_27640);
xnor U28523 (N_28523,N_27201,N_26333);
or U28524 (N_28524,N_26239,N_27009);
nor U28525 (N_28525,N_27852,N_26815);
nand U28526 (N_28526,N_27079,N_26436);
and U28527 (N_28527,N_26902,N_26405);
and U28528 (N_28528,N_26236,N_26215);
or U28529 (N_28529,N_27657,N_26719);
and U28530 (N_28530,N_26670,N_26981);
xor U28531 (N_28531,N_27604,N_27990);
nand U28532 (N_28532,N_27166,N_26564);
or U28533 (N_28533,N_27386,N_27204);
or U28534 (N_28534,N_27307,N_27109);
or U28535 (N_28535,N_27728,N_27298);
nand U28536 (N_28536,N_26082,N_27232);
and U28537 (N_28537,N_26697,N_27922);
xor U28538 (N_28538,N_26152,N_26404);
or U28539 (N_28539,N_26359,N_27061);
and U28540 (N_28540,N_26101,N_26338);
nor U28541 (N_28541,N_27041,N_26350);
and U28542 (N_28542,N_27736,N_27196);
and U28543 (N_28543,N_27048,N_27365);
xnor U28544 (N_28544,N_26119,N_27384);
xor U28545 (N_28545,N_27927,N_27814);
xor U28546 (N_28546,N_27575,N_26956);
xnor U28547 (N_28547,N_27596,N_26470);
xor U28548 (N_28548,N_26611,N_26278);
nand U28549 (N_28549,N_27182,N_26281);
and U28550 (N_28550,N_27688,N_26538);
nor U28551 (N_28551,N_26928,N_26231);
xor U28552 (N_28552,N_26725,N_26017);
nor U28553 (N_28553,N_27943,N_26446);
and U28554 (N_28554,N_26649,N_26751);
and U28555 (N_28555,N_26540,N_27250);
or U28556 (N_28556,N_27177,N_27626);
xnor U28557 (N_28557,N_27244,N_27445);
and U28558 (N_28558,N_27221,N_26015);
or U28559 (N_28559,N_27659,N_27644);
and U28560 (N_28560,N_26154,N_27528);
nand U28561 (N_28561,N_26508,N_27412);
and U28562 (N_28562,N_26133,N_27869);
or U28563 (N_28563,N_27797,N_26683);
nand U28564 (N_28564,N_27582,N_27744);
nand U28565 (N_28565,N_27687,N_26346);
and U28566 (N_28566,N_27719,N_26168);
and U28567 (N_28567,N_27170,N_26663);
and U28568 (N_28568,N_27123,N_27697);
xor U28569 (N_28569,N_27188,N_27612);
xor U28570 (N_28570,N_27481,N_26973);
or U28571 (N_28571,N_27713,N_27533);
or U28572 (N_28572,N_27047,N_26014);
nand U28573 (N_28573,N_27807,N_26161);
nand U28574 (N_28574,N_26929,N_27036);
and U28575 (N_28575,N_26450,N_26155);
and U28576 (N_28576,N_27965,N_26796);
xnor U28577 (N_28577,N_27332,N_27032);
xor U28578 (N_28578,N_27831,N_27463);
nand U28579 (N_28579,N_26615,N_27197);
nor U28580 (N_28580,N_27714,N_26534);
nor U28581 (N_28581,N_27105,N_27089);
or U28582 (N_28582,N_27092,N_26667);
nand U28583 (N_28583,N_27841,N_27894);
nand U28584 (N_28584,N_27095,N_27777);
nand U28585 (N_28585,N_26021,N_26006);
or U28586 (N_28586,N_27665,N_26539);
nand U28587 (N_28587,N_27124,N_26931);
xnor U28588 (N_28588,N_26959,N_26002);
and U28589 (N_28589,N_26877,N_27926);
or U28590 (N_28590,N_27071,N_26003);
nand U28591 (N_28591,N_27436,N_26894);
and U28592 (N_28592,N_26362,N_26208);
nand U28593 (N_28593,N_26300,N_26329);
and U28594 (N_28594,N_27129,N_27637);
and U28595 (N_28595,N_26098,N_27571);
nand U28596 (N_28596,N_26581,N_27843);
xor U28597 (N_28597,N_26631,N_27709);
nor U28598 (N_28598,N_26289,N_27909);
or U28599 (N_28599,N_26662,N_26923);
nand U28600 (N_28600,N_26330,N_26655);
and U28601 (N_28601,N_26761,N_26051);
nand U28602 (N_28602,N_27914,N_27054);
or U28603 (N_28603,N_27468,N_27133);
or U28604 (N_28604,N_26084,N_26997);
nand U28605 (N_28605,N_27784,N_27520);
nor U28606 (N_28606,N_26160,N_26616);
xnor U28607 (N_28607,N_26444,N_27278);
nor U28608 (N_28608,N_27648,N_26012);
xor U28609 (N_28609,N_27419,N_26102);
and U28610 (N_28610,N_26587,N_26205);
nor U28611 (N_28611,N_26964,N_27485);
nor U28612 (N_28612,N_26842,N_26839);
nand U28613 (N_28613,N_26066,N_27795);
nand U28614 (N_28614,N_26886,N_26286);
or U28615 (N_28615,N_26189,N_26965);
nor U28616 (N_28616,N_26456,N_27155);
or U28617 (N_28617,N_26390,N_26632);
xor U28618 (N_28618,N_26580,N_27599);
xor U28619 (N_28619,N_26647,N_27686);
xor U28620 (N_28620,N_26638,N_26106);
nor U28621 (N_28621,N_26735,N_26882);
or U28622 (N_28622,N_27608,N_27939);
xor U28623 (N_28623,N_26402,N_27516);
and U28624 (N_28624,N_26287,N_26408);
or U28625 (N_28625,N_27477,N_26497);
and U28626 (N_28626,N_26143,N_27388);
and U28627 (N_28627,N_27583,N_26778);
nor U28628 (N_28628,N_27912,N_26232);
or U28629 (N_28629,N_26837,N_27053);
nand U28630 (N_28630,N_27446,N_26324);
nand U28631 (N_28631,N_26876,N_27870);
or U28632 (N_28632,N_27459,N_27081);
xnor U28633 (N_28633,N_27035,N_26925);
xnor U28634 (N_28634,N_27891,N_26585);
nor U28635 (N_28635,N_27472,N_26803);
xnor U28636 (N_28636,N_26142,N_26245);
nand U28637 (N_28637,N_27220,N_27172);
xnor U28638 (N_28638,N_26033,N_27359);
or U28639 (N_28639,N_27429,N_26688);
nor U28640 (N_28640,N_27450,N_27351);
or U28641 (N_28641,N_26481,N_27016);
nand U28642 (N_28642,N_27660,N_27195);
nor U28643 (N_28643,N_27562,N_27174);
nor U28644 (N_28644,N_26926,N_27050);
xor U28645 (N_28645,N_26009,N_26600);
xnor U28646 (N_28646,N_27964,N_26556);
and U28647 (N_28647,N_26733,N_27457);
nor U28648 (N_28648,N_26786,N_27205);
nand U28649 (N_28649,N_26442,N_27501);
or U28650 (N_28650,N_27544,N_26698);
nor U28651 (N_28651,N_27667,N_27826);
or U28652 (N_28652,N_26990,N_27529);
nand U28653 (N_28653,N_26737,N_26087);
or U28654 (N_28654,N_26827,N_27269);
or U28655 (N_28655,N_26520,N_26887);
nand U28656 (N_28656,N_26490,N_27791);
xor U28657 (N_28657,N_26448,N_27745);
nor U28658 (N_28658,N_27579,N_27901);
and U28659 (N_28659,N_26824,N_27638);
nand U28660 (N_28660,N_26035,N_26863);
xnor U28661 (N_28661,N_26365,N_27732);
or U28662 (N_28662,N_27337,N_26153);
or U28663 (N_28663,N_26034,N_26429);
nand U28664 (N_28664,N_26857,N_26781);
xor U28665 (N_28665,N_26855,N_26267);
or U28666 (N_28666,N_27787,N_27159);
nor U28667 (N_28667,N_27518,N_26692);
or U28668 (N_28668,N_27854,N_27248);
nor U28669 (N_28669,N_26328,N_26722);
nor U28670 (N_28670,N_27600,N_27502);
xor U28671 (N_28671,N_27565,N_26204);
or U28672 (N_28672,N_27102,N_26339);
xnor U28673 (N_28673,N_27703,N_26462);
nand U28674 (N_28674,N_27723,N_27613);
nand U28675 (N_28675,N_27804,N_26158);
nor U28676 (N_28676,N_27128,N_27335);
and U28677 (N_28677,N_26940,N_26437);
nand U28678 (N_28678,N_27700,N_26496);
nand U28679 (N_28679,N_26734,N_26366);
nor U28680 (N_28680,N_26026,N_26316);
xnor U28681 (N_28681,N_27525,N_26776);
and U28682 (N_28682,N_26209,N_26628);
or U28683 (N_28683,N_27414,N_26319);
nor U28684 (N_28684,N_26807,N_27493);
nand U28685 (N_28685,N_27296,N_26506);
nor U28686 (N_28686,N_27216,N_27642);
xor U28687 (N_28687,N_27534,N_27559);
or U28688 (N_28688,N_26062,N_26811);
nand U28689 (N_28689,N_26793,N_27366);
nor U28690 (N_28690,N_26109,N_27402);
xor U28691 (N_28691,N_27038,N_26367);
nand U28692 (N_28692,N_26671,N_26577);
xor U28693 (N_28693,N_27782,N_26899);
nor U28694 (N_28694,N_26500,N_26757);
or U28695 (N_28695,N_26257,N_26313);
or U28696 (N_28696,N_27974,N_26031);
or U28697 (N_28697,N_26050,N_26175);
nand U28698 (N_28698,N_26280,N_27997);
and U28699 (N_28699,N_27303,N_27910);
and U28700 (N_28700,N_26933,N_27262);
or U28701 (N_28701,N_26746,N_27448);
and U28702 (N_28702,N_27209,N_27837);
and U28703 (N_28703,N_26273,N_26400);
or U28704 (N_28704,N_27295,N_27680);
and U28705 (N_28705,N_27847,N_27701);
nand U28706 (N_28706,N_26702,N_26220);
nand U28707 (N_28707,N_26995,N_27521);
or U28708 (N_28708,N_27976,N_26728);
nor U28709 (N_28709,N_27242,N_27846);
or U28710 (N_28710,N_26870,N_26258);
nor U28711 (N_28711,N_27290,N_27473);
nand U28712 (N_28712,N_26453,N_26071);
nor U28713 (N_28713,N_26597,N_26410);
or U28714 (N_28714,N_26111,N_26679);
and U28715 (N_28715,N_27304,N_26447);
nand U28716 (N_28716,N_26535,N_26454);
xor U28717 (N_28717,N_26937,N_27470);
and U28718 (N_28718,N_26752,N_27441);
xnor U28719 (N_28719,N_27515,N_27690);
nor U28720 (N_28720,N_26570,N_26523);
or U28721 (N_28721,N_26797,N_27437);
nand U28722 (N_28722,N_27157,N_26235);
or U28723 (N_28723,N_26187,N_27560);
and U28724 (N_28724,N_27039,N_26665);
xor U28725 (N_28725,N_27963,N_26893);
xnor U28726 (N_28726,N_26282,N_27707);
or U28727 (N_28727,N_26415,N_27193);
or U28728 (N_28728,N_27918,N_27002);
xor U28729 (N_28729,N_27030,N_26318);
xnor U28730 (N_28730,N_26769,N_26785);
and U28731 (N_28731,N_26768,N_27052);
nand U28732 (N_28732,N_26543,N_27552);
and U28733 (N_28733,N_26504,N_27628);
or U28734 (N_28734,N_27921,N_27431);
nor U28735 (N_28735,N_26533,N_27788);
or U28736 (N_28736,N_26901,N_26825);
or U28737 (N_28737,N_26948,N_26325);
xor U28738 (N_28738,N_27775,N_26748);
xor U28739 (N_28739,N_26513,N_27125);
xor U28740 (N_28740,N_26591,N_26696);
nand U28741 (N_28741,N_26292,N_26780);
nor U28742 (N_28742,N_26542,N_26397);
and U28743 (N_28743,N_26915,N_26930);
and U28744 (N_28744,N_27246,N_26610);
xnor U28745 (N_28745,N_27864,N_27161);
xor U28746 (N_28746,N_27003,N_26382);
or U28747 (N_28747,N_27449,N_26401);
xnor U28748 (N_28748,N_26343,N_27558);
nor U28749 (N_28749,N_26464,N_26763);
and U28750 (N_28750,N_26384,N_27555);
or U28751 (N_28751,N_26984,N_26067);
nor U28752 (N_28752,N_26736,N_26998);
and U28753 (N_28753,N_27617,N_26473);
nand U28754 (N_28754,N_26147,N_27247);
nand U28755 (N_28755,N_27945,N_26531);
and U28756 (N_28756,N_27389,N_26185);
nor U28757 (N_28757,N_26248,N_27907);
nor U28758 (N_28758,N_27853,N_26517);
nand U28759 (N_28759,N_26739,N_27983);
and U28760 (N_28760,N_27121,N_27871);
xor U28761 (N_28761,N_26117,N_27716);
nor U28762 (N_28762,N_27532,N_27735);
and U28763 (N_28763,N_27339,N_27264);
nand U28764 (N_28764,N_26946,N_26783);
or U28765 (N_28765,N_26557,N_26744);
xnor U28766 (N_28766,N_27391,N_27060);
nand U28767 (N_28767,N_26379,N_27663);
and U28768 (N_28768,N_26207,N_27526);
nor U28769 (N_28769,N_27970,N_26136);
xnor U28770 (N_28770,N_27274,N_27842);
and U28771 (N_28771,N_26924,N_27479);
nor U28772 (N_28772,N_27996,N_26968);
and U28773 (N_28773,N_27439,N_27024);
xor U28774 (N_28774,N_27018,N_27180);
and U28775 (N_28775,N_26912,N_26290);
or U28776 (N_28776,N_26898,N_26260);
or U28777 (N_28777,N_26426,N_27440);
nand U28778 (N_28778,N_26385,N_26243);
xor U28779 (N_28779,N_27884,N_26126);
and U28780 (N_28780,N_27428,N_27271);
and U28781 (N_28781,N_27882,N_27753);
nand U28782 (N_28782,N_26657,N_26466);
and U28783 (N_28783,N_26623,N_26920);
nand U28784 (N_28784,N_26486,N_27097);
xor U28785 (N_28785,N_27015,N_26356);
xor U28786 (N_28786,N_27317,N_26834);
and U28787 (N_28787,N_26214,N_27764);
nor U28788 (N_28788,N_27001,N_26323);
nand U28789 (N_28789,N_26395,N_27551);
nor U28790 (N_28790,N_27362,N_27899);
and U28791 (N_28791,N_26705,N_27796);
nand U28792 (N_28792,N_27080,N_26782);
xnor U28793 (N_28793,N_26104,N_27313);
xnor U28794 (N_28794,N_26375,N_26416);
nand U28795 (N_28795,N_26592,N_27132);
and U28796 (N_28796,N_26522,N_27360);
or U28797 (N_28797,N_27731,N_26656);
xor U28798 (N_28798,N_27734,N_27341);
nand U28799 (N_28799,N_27691,N_27759);
nand U28800 (N_28800,N_27136,N_26758);
nor U28801 (N_28801,N_26072,N_26266);
xnor U28802 (N_28802,N_26011,N_27620);
and U28803 (N_28803,N_26795,N_27354);
and U28804 (N_28804,N_26545,N_26831);
nand U28805 (N_28805,N_26853,N_27279);
nand U28806 (N_28806,N_26770,N_26095);
or U28807 (N_28807,N_26039,N_27265);
or U28808 (N_28808,N_26983,N_26977);
and U28809 (N_28809,N_26895,N_26790);
or U28810 (N_28810,N_26459,N_27851);
nor U28811 (N_28811,N_27815,N_27543);
nor U28812 (N_28812,N_27474,N_26955);
nand U28813 (N_28813,N_26627,N_27711);
and U28814 (N_28814,N_26658,N_27456);
xnor U28815 (N_28815,N_27873,N_26760);
xnor U28816 (N_28816,N_27769,N_26268);
xor U28817 (N_28817,N_27510,N_27005);
nand U28818 (N_28818,N_26085,N_26771);
nor U28819 (N_28819,N_27761,N_27750);
nor U28820 (N_28820,N_27361,N_26483);
or U28821 (N_28821,N_26202,N_27752);
nand U28822 (N_28822,N_26906,N_27406);
nand U28823 (N_28823,N_27033,N_27756);
xnor U28824 (N_28824,N_27803,N_27724);
nor U28825 (N_28825,N_27651,N_26059);
or U28826 (N_28826,N_27738,N_26891);
or U28827 (N_28827,N_27396,N_26856);
xor U28828 (N_28828,N_27322,N_26186);
xor U28829 (N_28829,N_26079,N_27435);
and U28830 (N_28830,N_26953,N_26495);
and U28831 (N_28831,N_27000,N_27390);
or U28832 (N_28832,N_27860,N_26479);
nand U28833 (N_28833,N_26484,N_27749);
or U28834 (N_28834,N_27037,N_27381);
or U28835 (N_28835,N_26376,N_26276);
nand U28836 (N_28836,N_27065,N_26115);
nor U28837 (N_28837,N_27331,N_27740);
nand U28838 (N_28838,N_26427,N_26418);
xnor U28839 (N_28839,N_27482,N_26198);
nor U28840 (N_28840,N_26335,N_26223);
or U28841 (N_28841,N_27212,N_27643);
and U28842 (N_28842,N_27497,N_27904);
nand U28843 (N_28843,N_27653,N_27400);
nand U28844 (N_28844,N_27098,N_27057);
nand U28845 (N_28845,N_26584,N_27517);
and U28846 (N_28846,N_26129,N_27862);
xnor U28847 (N_28847,N_27946,N_26633);
nor U28848 (N_28848,N_27288,N_26560);
xor U28849 (N_28849,N_27898,N_26478);
nand U28850 (N_28850,N_26422,N_27816);
xor U28851 (N_28851,N_27546,N_26691);
or U28852 (N_28852,N_26089,N_27720);
or U28853 (N_28853,N_27972,N_26263);
nor U28854 (N_28854,N_26844,N_26918);
nor U28855 (N_28855,N_27227,N_26987);
and U28856 (N_28856,N_27607,N_27045);
nand U28857 (N_28857,N_26246,N_27819);
nand U28858 (N_28858,N_26070,N_27952);
and U28859 (N_28859,N_27991,N_26057);
and U28860 (N_28860,N_27433,N_27765);
nand U28861 (N_28861,N_27268,N_26951);
nand U28862 (N_28862,N_27570,N_26594);
nor U28863 (N_28863,N_27919,N_26699);
nand U28864 (N_28864,N_27995,N_26766);
xnor U28865 (N_28865,N_27256,N_26460);
nor U28866 (N_28866,N_27270,N_27198);
xor U28867 (N_28867,N_26226,N_26173);
or U28868 (N_28868,N_27936,N_27126);
xnor U28869 (N_28869,N_26081,N_27466);
xor U28870 (N_28870,N_27810,N_26909);
and U28871 (N_28871,N_27839,N_26064);
nor U28872 (N_28872,N_26669,N_26678);
nand U28873 (N_28873,N_26455,N_26047);
and U28874 (N_28874,N_27330,N_27742);
nand U28875 (N_28875,N_27805,N_26309);
nor U28876 (N_28876,N_26061,N_27140);
nor U28877 (N_28877,N_26122,N_27702);
xnor U28878 (N_28878,N_26859,N_26565);
or U28879 (N_28879,N_27425,N_26262);
xor U28880 (N_28880,N_27622,N_26482);
and U28881 (N_28881,N_27422,N_27917);
xnor U28882 (N_28882,N_26502,N_27985);
xor U28883 (N_28883,N_26866,N_27122);
nand U28884 (N_28884,N_27992,N_26840);
and U28885 (N_28885,N_26029,N_27708);
nand U28886 (N_28886,N_26798,N_26063);
xnor U28887 (N_28887,N_27957,N_26217);
xor U28888 (N_28888,N_27410,N_26532);
or U28889 (N_28889,N_26841,N_26625);
nor U28890 (N_28890,N_26558,N_27556);
or U28891 (N_28891,N_26348,N_27214);
nand U28892 (N_28892,N_26042,N_26100);
nor U28893 (N_28893,N_27848,N_26828);
xnor U28894 (N_28894,N_27760,N_27950);
xor U28895 (N_28895,N_27324,N_27006);
nor U28896 (N_28896,N_26684,N_27028);
nor U28897 (N_28897,N_26917,N_27116);
nand U28898 (N_28898,N_27689,N_27566);
xnor U28899 (N_28899,N_26646,N_26424);
nor U28900 (N_28900,N_27879,N_26849);
and U28901 (N_28901,N_27364,N_26934);
or U28902 (N_28902,N_27947,N_26306);
or U28903 (N_28903,N_26568,N_26001);
xnor U28904 (N_28904,N_26935,N_26288);
or U28905 (N_28905,N_26709,N_27444);
and U28906 (N_28906,N_27158,N_26261);
nand U28907 (N_28907,N_26192,N_26609);
xor U28908 (N_28908,N_27237,N_26049);
or U28909 (N_28909,N_26911,N_26075);
nand U28910 (N_28910,N_26396,N_27462);
xor U28911 (N_28911,N_26388,N_26296);
xor U28912 (N_28912,N_27664,N_26308);
nor U28913 (N_28913,N_27953,N_27928);
or U28914 (N_28914,N_27890,N_26599);
xnor U28915 (N_28915,N_27169,N_26554);
or U28916 (N_28916,N_27222,N_26000);
or U28917 (N_28917,N_26298,N_26921);
nand U28918 (N_28918,N_27200,N_26680);
or U28919 (N_28919,N_27940,N_26200);
xnor U28920 (N_28920,N_27131,N_27263);
xnor U28921 (N_28921,N_26393,N_27257);
xor U28922 (N_28922,N_26058,N_27368);
nor U28923 (N_28923,N_27609,N_26294);
xnor U28924 (N_28924,N_26686,N_27467);
and U28925 (N_28925,N_27602,N_27836);
nor U28926 (N_28926,N_26706,N_26271);
xnor U28927 (N_28927,N_26865,N_27492);
and U28928 (N_28928,N_27825,N_26749);
or U28929 (N_28929,N_26573,N_26020);
or U28930 (N_28930,N_27827,N_26105);
and U28931 (N_28931,N_27100,N_27084);
or U28932 (N_28932,N_26687,N_27913);
nor U28933 (N_28933,N_27137,N_26829);
nor U28934 (N_28934,N_26755,N_26791);
and U28935 (N_28935,N_26222,N_26219);
and U28936 (N_28936,N_27167,N_27547);
xnor U28937 (N_28937,N_27154,N_26157);
nand U28938 (N_28938,N_27549,N_26341);
nand U28939 (N_28939,N_27289,N_26608);
nand U28940 (N_28940,N_27217,N_27597);
and U28941 (N_28941,N_27611,N_26074);
xnor U28942 (N_28942,N_27416,N_26648);
and U28943 (N_28943,N_26718,N_27019);
xor U28944 (N_28944,N_26729,N_27645);
and U28945 (N_28945,N_27619,N_27586);
or U28946 (N_28946,N_27224,N_27915);
or U28947 (N_28947,N_26501,N_27880);
or U28948 (N_28948,N_27135,N_26092);
and U28949 (N_28949,N_26693,N_26352);
xor U28950 (N_28950,N_27715,N_26544);
nand U28951 (N_28951,N_27590,N_27569);
or U28952 (N_28952,N_26305,N_27794);
or U28953 (N_28953,N_27114,N_26954);
or U28954 (N_28954,N_26377,N_27875);
nor U28955 (N_28955,N_26673,N_27813);
nand U28956 (N_28956,N_27285,N_27187);
or U28957 (N_28957,N_27774,N_26682);
xor U28958 (N_28958,N_26336,N_26018);
xnor U28959 (N_28959,N_26413,N_27252);
nand U28960 (N_28960,N_26088,N_26492);
nor U28961 (N_28961,N_26963,N_27696);
xnor U28962 (N_28962,N_27900,N_26423);
nand U28963 (N_28963,N_26118,N_26809);
and U28964 (N_28964,N_26144,N_26237);
nor U28965 (N_28965,N_26146,N_26708);
xnor U28966 (N_28966,N_26383,N_26254);
nor U28967 (N_28967,N_27908,N_26784);
and U28968 (N_28968,N_26635,N_26685);
nand U28969 (N_28969,N_27577,N_26432);
nand U28970 (N_28970,N_26715,N_27218);
and U28971 (N_28971,N_27443,N_27832);
nor U28972 (N_28972,N_26526,N_27150);
nand U28973 (N_28973,N_27859,N_26127);
xor U28974 (N_28974,N_27820,N_27369);
xnor U28975 (N_28975,N_27108,N_27106);
xor U28976 (N_28976,N_27143,N_27757);
and U28977 (N_28977,N_26005,N_26344);
xnor U28978 (N_28978,N_26843,N_27994);
nand U28979 (N_28979,N_26812,N_27461);
or U28980 (N_28980,N_26690,N_27942);
or U28981 (N_28981,N_27297,N_26883);
nor U28982 (N_28982,N_26040,N_27395);
nand U28983 (N_28983,N_27962,N_26604);
or U28984 (N_28984,N_26986,N_26668);
nand U28985 (N_28985,N_26149,N_27074);
nor U28986 (N_28986,N_27393,N_26303);
or U28987 (N_28987,N_27107,N_27087);
nor U28988 (N_28988,N_27968,N_27704);
nand U28989 (N_28989,N_27833,N_26477);
nand U28990 (N_28990,N_27152,N_26541);
nand U28991 (N_28991,N_26991,N_27646);
or U28992 (N_28992,N_26932,N_27798);
nor U28993 (N_28993,N_27527,N_27309);
or U28994 (N_28994,N_27916,N_26742);
and U28995 (N_28995,N_27865,N_26240);
nand U28996 (N_28996,N_26962,N_27210);
nand U28997 (N_28997,N_27046,N_26707);
or U28998 (N_28998,N_26561,N_27584);
or U28999 (N_28999,N_27063,N_26032);
and U29000 (N_29000,N_26017,N_27748);
and U29001 (N_29001,N_27381,N_27029);
nor U29002 (N_29002,N_27979,N_27109);
nand U29003 (N_29003,N_27986,N_27755);
nor U29004 (N_29004,N_27358,N_27384);
or U29005 (N_29005,N_27489,N_26293);
and U29006 (N_29006,N_27643,N_26173);
nand U29007 (N_29007,N_26360,N_26620);
or U29008 (N_29008,N_26236,N_26297);
xnor U29009 (N_29009,N_26516,N_27692);
or U29010 (N_29010,N_27295,N_27285);
nor U29011 (N_29011,N_26272,N_27823);
or U29012 (N_29012,N_26556,N_26521);
and U29013 (N_29013,N_26148,N_27369);
or U29014 (N_29014,N_26055,N_27805);
xnor U29015 (N_29015,N_26503,N_26152);
or U29016 (N_29016,N_27926,N_27810);
nand U29017 (N_29017,N_27160,N_27244);
xnor U29018 (N_29018,N_26671,N_26780);
nor U29019 (N_29019,N_27162,N_26321);
xnor U29020 (N_29020,N_26164,N_26076);
nand U29021 (N_29021,N_27705,N_27853);
nor U29022 (N_29022,N_27138,N_27236);
nand U29023 (N_29023,N_27387,N_27236);
nor U29024 (N_29024,N_27667,N_26102);
nor U29025 (N_29025,N_27239,N_26986);
nand U29026 (N_29026,N_27426,N_26341);
and U29027 (N_29027,N_26928,N_26708);
nor U29028 (N_29028,N_27303,N_27997);
nor U29029 (N_29029,N_26423,N_26471);
nor U29030 (N_29030,N_26683,N_27271);
and U29031 (N_29031,N_27013,N_26768);
xor U29032 (N_29032,N_26152,N_27692);
and U29033 (N_29033,N_26169,N_27523);
nor U29034 (N_29034,N_26376,N_26992);
and U29035 (N_29035,N_27519,N_27666);
or U29036 (N_29036,N_27160,N_27746);
nor U29037 (N_29037,N_27561,N_26615);
nand U29038 (N_29038,N_26700,N_27337);
and U29039 (N_29039,N_27381,N_27771);
nor U29040 (N_29040,N_26419,N_27809);
xnor U29041 (N_29041,N_26835,N_27364);
xnor U29042 (N_29042,N_26863,N_26833);
nor U29043 (N_29043,N_27227,N_26424);
and U29044 (N_29044,N_26811,N_26369);
nor U29045 (N_29045,N_27678,N_26547);
and U29046 (N_29046,N_26851,N_27438);
nor U29047 (N_29047,N_26204,N_27839);
or U29048 (N_29048,N_26590,N_26346);
nand U29049 (N_29049,N_26220,N_26744);
nand U29050 (N_29050,N_27269,N_27190);
and U29051 (N_29051,N_26038,N_26204);
xnor U29052 (N_29052,N_27427,N_27009);
nand U29053 (N_29053,N_27070,N_26047);
or U29054 (N_29054,N_27100,N_27713);
xnor U29055 (N_29055,N_26397,N_26731);
and U29056 (N_29056,N_27348,N_27292);
nor U29057 (N_29057,N_27345,N_26192);
xor U29058 (N_29058,N_27703,N_27720);
nor U29059 (N_29059,N_27651,N_26313);
nor U29060 (N_29060,N_27810,N_26996);
or U29061 (N_29061,N_26256,N_27018);
and U29062 (N_29062,N_27883,N_26059);
nor U29063 (N_29063,N_27928,N_27636);
nor U29064 (N_29064,N_26393,N_27343);
or U29065 (N_29065,N_26132,N_27554);
and U29066 (N_29066,N_27870,N_26970);
nor U29067 (N_29067,N_26876,N_27533);
nor U29068 (N_29068,N_26202,N_26971);
nand U29069 (N_29069,N_27862,N_26578);
nor U29070 (N_29070,N_26944,N_26959);
and U29071 (N_29071,N_27463,N_27023);
or U29072 (N_29072,N_26656,N_27360);
nand U29073 (N_29073,N_26768,N_26999);
nor U29074 (N_29074,N_26258,N_26781);
nand U29075 (N_29075,N_27682,N_26562);
and U29076 (N_29076,N_26187,N_26658);
nand U29077 (N_29077,N_26242,N_27316);
xnor U29078 (N_29078,N_27716,N_26923);
and U29079 (N_29079,N_27343,N_27249);
or U29080 (N_29080,N_26384,N_27174);
nor U29081 (N_29081,N_26534,N_27923);
nand U29082 (N_29082,N_27678,N_26969);
or U29083 (N_29083,N_27842,N_26466);
and U29084 (N_29084,N_26529,N_27611);
nor U29085 (N_29085,N_27081,N_27858);
and U29086 (N_29086,N_27824,N_26541);
nor U29087 (N_29087,N_27834,N_27998);
and U29088 (N_29088,N_27934,N_27312);
xnor U29089 (N_29089,N_26683,N_27406);
xnor U29090 (N_29090,N_26741,N_26322);
and U29091 (N_29091,N_27256,N_26376);
nor U29092 (N_29092,N_26697,N_27370);
xnor U29093 (N_29093,N_27944,N_26777);
nand U29094 (N_29094,N_27970,N_27253);
and U29095 (N_29095,N_26977,N_26147);
nor U29096 (N_29096,N_27469,N_27152);
xnor U29097 (N_29097,N_27284,N_26224);
nor U29098 (N_29098,N_26705,N_26694);
or U29099 (N_29099,N_27343,N_27485);
nor U29100 (N_29100,N_27001,N_26002);
or U29101 (N_29101,N_27031,N_27700);
nand U29102 (N_29102,N_27328,N_27377);
or U29103 (N_29103,N_27698,N_27891);
or U29104 (N_29104,N_26111,N_27438);
or U29105 (N_29105,N_26109,N_27866);
and U29106 (N_29106,N_26249,N_27978);
xnor U29107 (N_29107,N_27607,N_26745);
nand U29108 (N_29108,N_26144,N_26777);
or U29109 (N_29109,N_26317,N_27741);
nor U29110 (N_29110,N_27996,N_27083);
and U29111 (N_29111,N_27593,N_26597);
nand U29112 (N_29112,N_27933,N_27983);
and U29113 (N_29113,N_27127,N_27407);
nor U29114 (N_29114,N_27058,N_26438);
xnor U29115 (N_29115,N_27754,N_26694);
nand U29116 (N_29116,N_27519,N_26784);
xnor U29117 (N_29117,N_27108,N_26423);
nor U29118 (N_29118,N_27504,N_27839);
or U29119 (N_29119,N_26050,N_26838);
nand U29120 (N_29120,N_27649,N_26613);
nor U29121 (N_29121,N_27347,N_27702);
nor U29122 (N_29122,N_27260,N_26412);
xor U29123 (N_29123,N_26255,N_27897);
nor U29124 (N_29124,N_27794,N_26994);
nor U29125 (N_29125,N_26265,N_27367);
nand U29126 (N_29126,N_26882,N_27960);
nand U29127 (N_29127,N_27490,N_26130);
nand U29128 (N_29128,N_27467,N_26250);
nand U29129 (N_29129,N_26117,N_26637);
nand U29130 (N_29130,N_26101,N_27338);
and U29131 (N_29131,N_26000,N_27269);
or U29132 (N_29132,N_26126,N_27169);
and U29133 (N_29133,N_26760,N_27390);
nor U29134 (N_29134,N_27315,N_26345);
nand U29135 (N_29135,N_26829,N_26014);
and U29136 (N_29136,N_26988,N_26709);
xnor U29137 (N_29137,N_26434,N_26968);
or U29138 (N_29138,N_26351,N_27113);
nor U29139 (N_29139,N_26426,N_27382);
nor U29140 (N_29140,N_27232,N_26062);
nand U29141 (N_29141,N_26567,N_27039);
xor U29142 (N_29142,N_26219,N_26111);
nand U29143 (N_29143,N_26787,N_27468);
nand U29144 (N_29144,N_26030,N_26476);
xnor U29145 (N_29145,N_27292,N_26095);
and U29146 (N_29146,N_26814,N_26749);
nor U29147 (N_29147,N_26444,N_26192);
and U29148 (N_29148,N_26027,N_26051);
or U29149 (N_29149,N_26938,N_26264);
xor U29150 (N_29150,N_27459,N_26753);
nor U29151 (N_29151,N_26205,N_27916);
nand U29152 (N_29152,N_26365,N_26235);
xor U29153 (N_29153,N_26250,N_26413);
nand U29154 (N_29154,N_27069,N_27511);
and U29155 (N_29155,N_27004,N_27179);
xor U29156 (N_29156,N_26399,N_27992);
nor U29157 (N_29157,N_26937,N_26955);
nor U29158 (N_29158,N_26719,N_27926);
or U29159 (N_29159,N_26460,N_26006);
nand U29160 (N_29160,N_27497,N_26977);
and U29161 (N_29161,N_26731,N_27839);
nor U29162 (N_29162,N_26872,N_27957);
or U29163 (N_29163,N_27349,N_27677);
nor U29164 (N_29164,N_26075,N_26512);
xnor U29165 (N_29165,N_26072,N_27333);
and U29166 (N_29166,N_27095,N_26927);
nand U29167 (N_29167,N_26810,N_26620);
xor U29168 (N_29168,N_26492,N_27156);
and U29169 (N_29169,N_27754,N_27712);
nand U29170 (N_29170,N_26307,N_26280);
nor U29171 (N_29171,N_27104,N_27897);
nand U29172 (N_29172,N_27145,N_26518);
or U29173 (N_29173,N_27454,N_27819);
nand U29174 (N_29174,N_26515,N_26768);
xnor U29175 (N_29175,N_26078,N_26542);
and U29176 (N_29176,N_26504,N_26079);
xor U29177 (N_29177,N_27263,N_26610);
nor U29178 (N_29178,N_26551,N_26313);
or U29179 (N_29179,N_26220,N_27554);
or U29180 (N_29180,N_26487,N_26866);
nor U29181 (N_29181,N_27047,N_26468);
or U29182 (N_29182,N_26736,N_27542);
or U29183 (N_29183,N_27250,N_26552);
xnor U29184 (N_29184,N_26704,N_27809);
and U29185 (N_29185,N_27553,N_26546);
nor U29186 (N_29186,N_27849,N_26111);
nor U29187 (N_29187,N_26036,N_27313);
nor U29188 (N_29188,N_26395,N_27020);
xnor U29189 (N_29189,N_27756,N_27309);
nand U29190 (N_29190,N_27395,N_26519);
and U29191 (N_29191,N_27795,N_27521);
xnor U29192 (N_29192,N_26858,N_26754);
xnor U29193 (N_29193,N_26809,N_27801);
and U29194 (N_29194,N_27386,N_27037);
and U29195 (N_29195,N_26088,N_26629);
nor U29196 (N_29196,N_27674,N_27804);
xor U29197 (N_29197,N_27017,N_26222);
nand U29198 (N_29198,N_27621,N_27097);
xnor U29199 (N_29199,N_26486,N_27401);
nand U29200 (N_29200,N_27022,N_27802);
nand U29201 (N_29201,N_27641,N_27905);
xnor U29202 (N_29202,N_27247,N_27328);
nor U29203 (N_29203,N_26447,N_26422);
or U29204 (N_29204,N_26547,N_26890);
nor U29205 (N_29205,N_26056,N_26969);
and U29206 (N_29206,N_27738,N_26655);
nand U29207 (N_29207,N_26356,N_27286);
and U29208 (N_29208,N_27694,N_26018);
xor U29209 (N_29209,N_27868,N_27323);
nor U29210 (N_29210,N_27384,N_27409);
nor U29211 (N_29211,N_27800,N_26715);
and U29212 (N_29212,N_27573,N_27331);
or U29213 (N_29213,N_26071,N_27579);
xor U29214 (N_29214,N_27346,N_26485);
or U29215 (N_29215,N_26878,N_26941);
and U29216 (N_29216,N_27210,N_26288);
or U29217 (N_29217,N_27324,N_27725);
nand U29218 (N_29218,N_27981,N_27201);
nor U29219 (N_29219,N_26931,N_27453);
and U29220 (N_29220,N_27192,N_26113);
and U29221 (N_29221,N_27552,N_27638);
or U29222 (N_29222,N_27766,N_27074);
xor U29223 (N_29223,N_27207,N_26738);
and U29224 (N_29224,N_26624,N_26907);
or U29225 (N_29225,N_26273,N_26872);
or U29226 (N_29226,N_26642,N_27397);
or U29227 (N_29227,N_27236,N_26575);
nand U29228 (N_29228,N_26246,N_26239);
or U29229 (N_29229,N_26448,N_26316);
nand U29230 (N_29230,N_26717,N_26029);
or U29231 (N_29231,N_27337,N_27792);
xor U29232 (N_29232,N_26888,N_27565);
or U29233 (N_29233,N_27334,N_27394);
or U29234 (N_29234,N_26499,N_27650);
xor U29235 (N_29235,N_26524,N_27786);
and U29236 (N_29236,N_27067,N_26878);
and U29237 (N_29237,N_26021,N_26601);
or U29238 (N_29238,N_27601,N_26999);
xor U29239 (N_29239,N_27988,N_26385);
xnor U29240 (N_29240,N_27692,N_27986);
or U29241 (N_29241,N_26233,N_27137);
xor U29242 (N_29242,N_27909,N_26497);
nand U29243 (N_29243,N_27157,N_26121);
and U29244 (N_29244,N_27948,N_26229);
nand U29245 (N_29245,N_26264,N_26209);
nand U29246 (N_29246,N_26588,N_27170);
xor U29247 (N_29247,N_27161,N_27361);
and U29248 (N_29248,N_27033,N_27804);
nand U29249 (N_29249,N_27416,N_27394);
nor U29250 (N_29250,N_27067,N_26563);
nand U29251 (N_29251,N_26163,N_27054);
and U29252 (N_29252,N_26025,N_27525);
xnor U29253 (N_29253,N_27044,N_26603);
and U29254 (N_29254,N_26383,N_26298);
nor U29255 (N_29255,N_27019,N_27774);
or U29256 (N_29256,N_27904,N_26860);
xor U29257 (N_29257,N_27728,N_26138);
and U29258 (N_29258,N_27121,N_26007);
and U29259 (N_29259,N_26706,N_27980);
nor U29260 (N_29260,N_26862,N_27007);
nand U29261 (N_29261,N_26988,N_27207);
xor U29262 (N_29262,N_27950,N_26238);
xnor U29263 (N_29263,N_26696,N_26300);
xnor U29264 (N_29264,N_27470,N_27542);
nor U29265 (N_29265,N_26969,N_26148);
nand U29266 (N_29266,N_27895,N_26521);
nor U29267 (N_29267,N_26076,N_26254);
or U29268 (N_29268,N_27181,N_27387);
nor U29269 (N_29269,N_27110,N_26206);
xor U29270 (N_29270,N_27505,N_26167);
nand U29271 (N_29271,N_26188,N_26661);
xor U29272 (N_29272,N_26077,N_27235);
xnor U29273 (N_29273,N_27062,N_27194);
nand U29274 (N_29274,N_26981,N_26742);
xnor U29275 (N_29275,N_27930,N_27432);
nor U29276 (N_29276,N_27174,N_26488);
xor U29277 (N_29277,N_27170,N_27342);
or U29278 (N_29278,N_27965,N_27917);
nand U29279 (N_29279,N_27415,N_27737);
and U29280 (N_29280,N_26119,N_27403);
nand U29281 (N_29281,N_26798,N_26184);
and U29282 (N_29282,N_26934,N_26044);
xnor U29283 (N_29283,N_27425,N_26775);
nor U29284 (N_29284,N_27705,N_26965);
xor U29285 (N_29285,N_27842,N_27882);
and U29286 (N_29286,N_27831,N_27100);
or U29287 (N_29287,N_27697,N_26571);
xnor U29288 (N_29288,N_26921,N_27157);
nor U29289 (N_29289,N_27155,N_27578);
or U29290 (N_29290,N_27794,N_27464);
nor U29291 (N_29291,N_27939,N_26496);
and U29292 (N_29292,N_27397,N_26355);
and U29293 (N_29293,N_27091,N_26664);
xnor U29294 (N_29294,N_26172,N_26185);
nand U29295 (N_29295,N_27896,N_26433);
and U29296 (N_29296,N_26585,N_27759);
nor U29297 (N_29297,N_27670,N_27407);
xnor U29298 (N_29298,N_27201,N_26960);
or U29299 (N_29299,N_27167,N_26398);
and U29300 (N_29300,N_26611,N_26110);
nand U29301 (N_29301,N_27194,N_27497);
or U29302 (N_29302,N_26637,N_26162);
xnor U29303 (N_29303,N_26803,N_27763);
xor U29304 (N_29304,N_27303,N_26125);
xnor U29305 (N_29305,N_26181,N_26682);
xnor U29306 (N_29306,N_26351,N_26651);
nor U29307 (N_29307,N_26940,N_26310);
or U29308 (N_29308,N_27340,N_27370);
and U29309 (N_29309,N_26531,N_26752);
and U29310 (N_29310,N_26777,N_26666);
xor U29311 (N_29311,N_26197,N_26889);
xnor U29312 (N_29312,N_26392,N_27649);
nand U29313 (N_29313,N_26911,N_27725);
or U29314 (N_29314,N_26248,N_27234);
or U29315 (N_29315,N_27790,N_26611);
nor U29316 (N_29316,N_26716,N_26939);
or U29317 (N_29317,N_26959,N_26811);
xnor U29318 (N_29318,N_27187,N_26998);
nor U29319 (N_29319,N_27393,N_26447);
xor U29320 (N_29320,N_27431,N_27789);
nor U29321 (N_29321,N_26234,N_26302);
and U29322 (N_29322,N_27386,N_26604);
and U29323 (N_29323,N_27035,N_26236);
and U29324 (N_29324,N_27941,N_26078);
nand U29325 (N_29325,N_26673,N_26079);
nor U29326 (N_29326,N_26555,N_26444);
and U29327 (N_29327,N_26513,N_26875);
or U29328 (N_29328,N_26626,N_27349);
nor U29329 (N_29329,N_26346,N_27507);
nand U29330 (N_29330,N_27636,N_27182);
and U29331 (N_29331,N_27465,N_27407);
xor U29332 (N_29332,N_26532,N_26593);
and U29333 (N_29333,N_27591,N_27710);
nor U29334 (N_29334,N_26963,N_26540);
nor U29335 (N_29335,N_27038,N_27311);
nand U29336 (N_29336,N_26106,N_27128);
or U29337 (N_29337,N_26669,N_26751);
nand U29338 (N_29338,N_27073,N_27962);
xnor U29339 (N_29339,N_26208,N_27030);
nor U29340 (N_29340,N_27060,N_27222);
nand U29341 (N_29341,N_27371,N_27361);
nor U29342 (N_29342,N_26566,N_27258);
and U29343 (N_29343,N_27212,N_26545);
nor U29344 (N_29344,N_27459,N_27143);
nor U29345 (N_29345,N_26435,N_26222);
nand U29346 (N_29346,N_26542,N_26950);
nor U29347 (N_29347,N_27790,N_26997);
nand U29348 (N_29348,N_27488,N_26276);
nand U29349 (N_29349,N_26623,N_27662);
xor U29350 (N_29350,N_26717,N_27853);
and U29351 (N_29351,N_26780,N_27622);
or U29352 (N_29352,N_27097,N_27745);
nand U29353 (N_29353,N_26020,N_27353);
nor U29354 (N_29354,N_26625,N_26602);
nand U29355 (N_29355,N_26967,N_26217);
and U29356 (N_29356,N_27747,N_26705);
and U29357 (N_29357,N_27722,N_27603);
and U29358 (N_29358,N_27692,N_27402);
xnor U29359 (N_29359,N_27165,N_26004);
nor U29360 (N_29360,N_26449,N_27846);
and U29361 (N_29361,N_26181,N_26089);
nand U29362 (N_29362,N_27311,N_27657);
nand U29363 (N_29363,N_26023,N_27864);
or U29364 (N_29364,N_26730,N_27727);
nand U29365 (N_29365,N_27432,N_27760);
and U29366 (N_29366,N_27638,N_27126);
nor U29367 (N_29367,N_27512,N_26860);
xor U29368 (N_29368,N_26904,N_27184);
nor U29369 (N_29369,N_27349,N_26913);
or U29370 (N_29370,N_27084,N_26147);
nor U29371 (N_29371,N_26703,N_27899);
xor U29372 (N_29372,N_26991,N_26539);
xnor U29373 (N_29373,N_26846,N_27838);
nor U29374 (N_29374,N_27956,N_27874);
nand U29375 (N_29375,N_27851,N_27143);
nor U29376 (N_29376,N_26938,N_27680);
xnor U29377 (N_29377,N_26815,N_27609);
xnor U29378 (N_29378,N_26978,N_27060);
xor U29379 (N_29379,N_27057,N_26345);
nand U29380 (N_29380,N_27009,N_26580);
nor U29381 (N_29381,N_26514,N_27036);
nand U29382 (N_29382,N_27908,N_26213);
or U29383 (N_29383,N_27303,N_26649);
or U29384 (N_29384,N_26078,N_27255);
and U29385 (N_29385,N_26489,N_26191);
nand U29386 (N_29386,N_27141,N_27904);
nor U29387 (N_29387,N_26406,N_27278);
and U29388 (N_29388,N_27148,N_27873);
or U29389 (N_29389,N_27384,N_27239);
nand U29390 (N_29390,N_26430,N_27044);
nor U29391 (N_29391,N_27432,N_27709);
or U29392 (N_29392,N_26306,N_26474);
or U29393 (N_29393,N_27298,N_27006);
xnor U29394 (N_29394,N_26069,N_26066);
or U29395 (N_29395,N_26091,N_26408);
and U29396 (N_29396,N_26406,N_26712);
nand U29397 (N_29397,N_27456,N_26056);
or U29398 (N_29398,N_26884,N_27372);
nand U29399 (N_29399,N_27791,N_27169);
and U29400 (N_29400,N_27407,N_26442);
or U29401 (N_29401,N_26708,N_27115);
nor U29402 (N_29402,N_26076,N_27676);
and U29403 (N_29403,N_26386,N_26401);
or U29404 (N_29404,N_26015,N_27763);
or U29405 (N_29405,N_26686,N_26168);
nor U29406 (N_29406,N_27675,N_26709);
or U29407 (N_29407,N_27203,N_27225);
or U29408 (N_29408,N_27782,N_27825);
xor U29409 (N_29409,N_26555,N_26809);
or U29410 (N_29410,N_27924,N_27478);
and U29411 (N_29411,N_27118,N_27221);
nand U29412 (N_29412,N_26531,N_26249);
nor U29413 (N_29413,N_26503,N_26723);
xor U29414 (N_29414,N_27742,N_26902);
xor U29415 (N_29415,N_26331,N_27430);
and U29416 (N_29416,N_26014,N_26452);
or U29417 (N_29417,N_27666,N_27548);
nand U29418 (N_29418,N_27037,N_27733);
nand U29419 (N_29419,N_26584,N_26165);
xnor U29420 (N_29420,N_27827,N_26630);
nor U29421 (N_29421,N_26530,N_27050);
xnor U29422 (N_29422,N_27357,N_27425);
nand U29423 (N_29423,N_26714,N_27584);
xor U29424 (N_29424,N_26902,N_27268);
or U29425 (N_29425,N_27071,N_26821);
or U29426 (N_29426,N_27880,N_26859);
or U29427 (N_29427,N_27337,N_27543);
nand U29428 (N_29428,N_26120,N_26931);
nand U29429 (N_29429,N_26955,N_27235);
nand U29430 (N_29430,N_27831,N_27012);
xor U29431 (N_29431,N_27223,N_26163);
or U29432 (N_29432,N_26526,N_27574);
nor U29433 (N_29433,N_27311,N_27049);
nor U29434 (N_29434,N_27814,N_26627);
or U29435 (N_29435,N_27811,N_27348);
xor U29436 (N_29436,N_26213,N_26661);
or U29437 (N_29437,N_26959,N_26401);
nor U29438 (N_29438,N_27734,N_27952);
and U29439 (N_29439,N_27871,N_26063);
nand U29440 (N_29440,N_27124,N_27316);
nor U29441 (N_29441,N_26995,N_26870);
nor U29442 (N_29442,N_27576,N_26923);
nand U29443 (N_29443,N_26409,N_26028);
or U29444 (N_29444,N_27074,N_27608);
and U29445 (N_29445,N_27277,N_26313);
or U29446 (N_29446,N_27264,N_26900);
and U29447 (N_29447,N_27183,N_27489);
nand U29448 (N_29448,N_26930,N_27288);
or U29449 (N_29449,N_26430,N_27624);
xor U29450 (N_29450,N_26448,N_27096);
and U29451 (N_29451,N_26582,N_26772);
nor U29452 (N_29452,N_27196,N_27146);
and U29453 (N_29453,N_27835,N_27074);
nand U29454 (N_29454,N_27890,N_26080);
or U29455 (N_29455,N_26088,N_26006);
or U29456 (N_29456,N_27139,N_27176);
nor U29457 (N_29457,N_26287,N_26599);
nand U29458 (N_29458,N_26249,N_27770);
nor U29459 (N_29459,N_26287,N_27919);
xor U29460 (N_29460,N_26056,N_27797);
or U29461 (N_29461,N_27547,N_27691);
or U29462 (N_29462,N_26080,N_27217);
and U29463 (N_29463,N_26400,N_27017);
nor U29464 (N_29464,N_27239,N_26909);
nor U29465 (N_29465,N_27028,N_27486);
or U29466 (N_29466,N_26660,N_27181);
nor U29467 (N_29467,N_27963,N_27634);
or U29468 (N_29468,N_26894,N_27985);
or U29469 (N_29469,N_27826,N_27399);
and U29470 (N_29470,N_26724,N_27891);
nand U29471 (N_29471,N_27325,N_27777);
nand U29472 (N_29472,N_26801,N_27109);
nor U29473 (N_29473,N_26970,N_26921);
or U29474 (N_29474,N_26600,N_27555);
xnor U29475 (N_29475,N_26204,N_26973);
and U29476 (N_29476,N_26266,N_27517);
or U29477 (N_29477,N_27561,N_26951);
or U29478 (N_29478,N_26110,N_27591);
and U29479 (N_29479,N_26372,N_27415);
or U29480 (N_29480,N_26651,N_27672);
and U29481 (N_29481,N_27674,N_27846);
xnor U29482 (N_29482,N_26501,N_26396);
nand U29483 (N_29483,N_26243,N_26811);
and U29484 (N_29484,N_27970,N_26077);
nand U29485 (N_29485,N_26467,N_26533);
nand U29486 (N_29486,N_26368,N_26724);
or U29487 (N_29487,N_26777,N_26767);
nor U29488 (N_29488,N_27445,N_26525);
or U29489 (N_29489,N_27090,N_27665);
xor U29490 (N_29490,N_26872,N_27891);
nand U29491 (N_29491,N_27636,N_27594);
nor U29492 (N_29492,N_26995,N_27119);
nand U29493 (N_29493,N_27892,N_27842);
xnor U29494 (N_29494,N_26039,N_27184);
and U29495 (N_29495,N_27166,N_27207);
and U29496 (N_29496,N_27779,N_26462);
nand U29497 (N_29497,N_26279,N_26459);
and U29498 (N_29498,N_26331,N_26779);
and U29499 (N_29499,N_27520,N_26423);
and U29500 (N_29500,N_27553,N_26658);
or U29501 (N_29501,N_26057,N_26552);
xnor U29502 (N_29502,N_27089,N_27473);
or U29503 (N_29503,N_27055,N_27232);
xor U29504 (N_29504,N_26316,N_27157);
or U29505 (N_29505,N_26705,N_27079);
or U29506 (N_29506,N_26765,N_27925);
nor U29507 (N_29507,N_27538,N_26907);
and U29508 (N_29508,N_27960,N_27905);
and U29509 (N_29509,N_27257,N_27579);
nand U29510 (N_29510,N_27261,N_27243);
or U29511 (N_29511,N_27611,N_27359);
or U29512 (N_29512,N_26803,N_26052);
xor U29513 (N_29513,N_27503,N_26888);
nor U29514 (N_29514,N_27215,N_26805);
or U29515 (N_29515,N_27388,N_27457);
or U29516 (N_29516,N_26696,N_27551);
nor U29517 (N_29517,N_26714,N_26785);
xnor U29518 (N_29518,N_27885,N_26344);
nand U29519 (N_29519,N_26839,N_27016);
and U29520 (N_29520,N_26508,N_26385);
nand U29521 (N_29521,N_26047,N_27809);
nand U29522 (N_29522,N_27614,N_26843);
nor U29523 (N_29523,N_26192,N_27664);
nor U29524 (N_29524,N_27555,N_27408);
nand U29525 (N_29525,N_26496,N_27609);
or U29526 (N_29526,N_26158,N_27895);
and U29527 (N_29527,N_26823,N_26883);
nand U29528 (N_29528,N_27687,N_27409);
and U29529 (N_29529,N_26200,N_26644);
and U29530 (N_29530,N_26872,N_27265);
nor U29531 (N_29531,N_27690,N_27818);
xnor U29532 (N_29532,N_26362,N_26571);
nor U29533 (N_29533,N_26443,N_27067);
and U29534 (N_29534,N_26203,N_27120);
and U29535 (N_29535,N_27356,N_26173);
nor U29536 (N_29536,N_26129,N_27357);
or U29537 (N_29537,N_26073,N_27718);
nand U29538 (N_29538,N_26162,N_26594);
nand U29539 (N_29539,N_27762,N_26365);
or U29540 (N_29540,N_26442,N_27246);
or U29541 (N_29541,N_26448,N_26283);
nand U29542 (N_29542,N_27356,N_26927);
nor U29543 (N_29543,N_27341,N_26723);
or U29544 (N_29544,N_26177,N_27542);
or U29545 (N_29545,N_26055,N_27606);
nor U29546 (N_29546,N_27132,N_27552);
nand U29547 (N_29547,N_27615,N_26104);
nor U29548 (N_29548,N_27528,N_27045);
or U29549 (N_29549,N_26991,N_27873);
or U29550 (N_29550,N_27685,N_27519);
or U29551 (N_29551,N_26669,N_27064);
nand U29552 (N_29552,N_27670,N_26931);
nor U29553 (N_29553,N_26828,N_26035);
and U29554 (N_29554,N_26395,N_27495);
and U29555 (N_29555,N_26081,N_26190);
and U29556 (N_29556,N_27203,N_26525);
xnor U29557 (N_29557,N_27677,N_27208);
xnor U29558 (N_29558,N_27649,N_26531);
nor U29559 (N_29559,N_26113,N_26914);
nand U29560 (N_29560,N_26245,N_27309);
xnor U29561 (N_29561,N_26709,N_26498);
xor U29562 (N_29562,N_27574,N_26063);
nor U29563 (N_29563,N_27704,N_27798);
xnor U29564 (N_29564,N_26247,N_27087);
nand U29565 (N_29565,N_27017,N_26518);
xor U29566 (N_29566,N_26222,N_27192);
xnor U29567 (N_29567,N_26034,N_27601);
or U29568 (N_29568,N_26371,N_26324);
nor U29569 (N_29569,N_26757,N_26264);
and U29570 (N_29570,N_27038,N_27499);
or U29571 (N_29571,N_27562,N_27389);
or U29572 (N_29572,N_26032,N_26199);
xnor U29573 (N_29573,N_26780,N_27093);
nor U29574 (N_29574,N_27642,N_26439);
or U29575 (N_29575,N_27617,N_27950);
or U29576 (N_29576,N_26068,N_26182);
nand U29577 (N_29577,N_26251,N_26195);
and U29578 (N_29578,N_26878,N_26410);
xor U29579 (N_29579,N_27365,N_27835);
nor U29580 (N_29580,N_26589,N_27671);
xor U29581 (N_29581,N_27876,N_27678);
and U29582 (N_29582,N_27629,N_26418);
or U29583 (N_29583,N_27038,N_27754);
xnor U29584 (N_29584,N_26959,N_26563);
xnor U29585 (N_29585,N_26295,N_27139);
or U29586 (N_29586,N_26168,N_27618);
nand U29587 (N_29587,N_27788,N_27949);
or U29588 (N_29588,N_27392,N_27375);
nand U29589 (N_29589,N_26469,N_26860);
xnor U29590 (N_29590,N_26138,N_26137);
xor U29591 (N_29591,N_26032,N_27740);
or U29592 (N_29592,N_26933,N_26384);
nor U29593 (N_29593,N_26717,N_27900);
nor U29594 (N_29594,N_26834,N_26992);
and U29595 (N_29595,N_26072,N_27053);
nor U29596 (N_29596,N_27576,N_26051);
xnor U29597 (N_29597,N_27016,N_27349);
nand U29598 (N_29598,N_26711,N_27225);
or U29599 (N_29599,N_27082,N_26223);
or U29600 (N_29600,N_27568,N_26538);
nand U29601 (N_29601,N_27908,N_26669);
nor U29602 (N_29602,N_26149,N_27161);
and U29603 (N_29603,N_26463,N_27292);
nor U29604 (N_29604,N_26868,N_26152);
xnor U29605 (N_29605,N_26745,N_26858);
or U29606 (N_29606,N_26826,N_26917);
xnor U29607 (N_29607,N_27721,N_26467);
or U29608 (N_29608,N_26787,N_27020);
xnor U29609 (N_29609,N_27702,N_27079);
nor U29610 (N_29610,N_27836,N_27742);
and U29611 (N_29611,N_26377,N_27570);
nand U29612 (N_29612,N_27828,N_27299);
or U29613 (N_29613,N_27581,N_27047);
xor U29614 (N_29614,N_26940,N_26091);
or U29615 (N_29615,N_26236,N_26273);
or U29616 (N_29616,N_26491,N_27834);
nand U29617 (N_29617,N_26557,N_26645);
xnor U29618 (N_29618,N_26504,N_27981);
and U29619 (N_29619,N_26287,N_26297);
or U29620 (N_29620,N_27556,N_27631);
or U29621 (N_29621,N_27523,N_27336);
xnor U29622 (N_29622,N_26148,N_26901);
or U29623 (N_29623,N_26451,N_26341);
or U29624 (N_29624,N_27557,N_27224);
xnor U29625 (N_29625,N_27188,N_27322);
xnor U29626 (N_29626,N_26003,N_27800);
nand U29627 (N_29627,N_26741,N_26371);
nor U29628 (N_29628,N_27272,N_27950);
or U29629 (N_29629,N_26923,N_26261);
nand U29630 (N_29630,N_27380,N_27981);
nand U29631 (N_29631,N_26882,N_27060);
nand U29632 (N_29632,N_27259,N_27178);
xor U29633 (N_29633,N_27973,N_26319);
nor U29634 (N_29634,N_27107,N_26596);
nand U29635 (N_29635,N_27980,N_27788);
nand U29636 (N_29636,N_26580,N_27447);
nor U29637 (N_29637,N_26334,N_27823);
or U29638 (N_29638,N_27254,N_26980);
and U29639 (N_29639,N_26407,N_27214);
and U29640 (N_29640,N_26925,N_27438);
nor U29641 (N_29641,N_26836,N_27274);
nor U29642 (N_29642,N_27174,N_26141);
or U29643 (N_29643,N_27945,N_27612);
and U29644 (N_29644,N_27507,N_26004);
or U29645 (N_29645,N_27744,N_26825);
xnor U29646 (N_29646,N_26619,N_27677);
and U29647 (N_29647,N_26216,N_26013);
and U29648 (N_29648,N_27870,N_27901);
and U29649 (N_29649,N_27286,N_26305);
xnor U29650 (N_29650,N_26773,N_26718);
xor U29651 (N_29651,N_27864,N_26153);
nor U29652 (N_29652,N_26856,N_27369);
nor U29653 (N_29653,N_26757,N_27052);
nor U29654 (N_29654,N_27560,N_27970);
and U29655 (N_29655,N_26175,N_27131);
xnor U29656 (N_29656,N_27619,N_27419);
or U29657 (N_29657,N_26476,N_26683);
xor U29658 (N_29658,N_26222,N_26771);
and U29659 (N_29659,N_26290,N_26882);
xnor U29660 (N_29660,N_27751,N_27673);
nand U29661 (N_29661,N_26938,N_27415);
and U29662 (N_29662,N_26182,N_27741);
nand U29663 (N_29663,N_26197,N_26534);
nand U29664 (N_29664,N_26797,N_26329);
or U29665 (N_29665,N_27698,N_26169);
or U29666 (N_29666,N_26327,N_26408);
or U29667 (N_29667,N_26808,N_27142);
or U29668 (N_29668,N_26860,N_27667);
and U29669 (N_29669,N_26809,N_27590);
and U29670 (N_29670,N_26736,N_27041);
or U29671 (N_29671,N_27060,N_26690);
and U29672 (N_29672,N_26792,N_26485);
xor U29673 (N_29673,N_27101,N_26038);
or U29674 (N_29674,N_26857,N_27305);
xor U29675 (N_29675,N_27340,N_26233);
or U29676 (N_29676,N_26481,N_26060);
nand U29677 (N_29677,N_27783,N_27492);
or U29678 (N_29678,N_27231,N_26703);
nor U29679 (N_29679,N_27911,N_26064);
and U29680 (N_29680,N_26297,N_27712);
nand U29681 (N_29681,N_26579,N_26917);
xor U29682 (N_29682,N_26276,N_27413);
nor U29683 (N_29683,N_27635,N_27886);
nor U29684 (N_29684,N_26913,N_26364);
or U29685 (N_29685,N_27760,N_27001);
nand U29686 (N_29686,N_27987,N_26970);
and U29687 (N_29687,N_27853,N_27625);
nand U29688 (N_29688,N_27369,N_27537);
and U29689 (N_29689,N_26279,N_27637);
nor U29690 (N_29690,N_27330,N_26914);
xor U29691 (N_29691,N_27065,N_26797);
xor U29692 (N_29692,N_27864,N_26411);
nand U29693 (N_29693,N_27118,N_26223);
and U29694 (N_29694,N_27663,N_27546);
xor U29695 (N_29695,N_26008,N_27385);
nor U29696 (N_29696,N_26729,N_26358);
xnor U29697 (N_29697,N_27333,N_26341);
xnor U29698 (N_29698,N_27444,N_27835);
or U29699 (N_29699,N_26986,N_27791);
nor U29700 (N_29700,N_26158,N_27811);
or U29701 (N_29701,N_27016,N_26660);
and U29702 (N_29702,N_26975,N_27422);
nor U29703 (N_29703,N_27380,N_27204);
nand U29704 (N_29704,N_26973,N_27107);
xor U29705 (N_29705,N_26592,N_26588);
nand U29706 (N_29706,N_27121,N_27224);
and U29707 (N_29707,N_27423,N_27207);
and U29708 (N_29708,N_27284,N_26175);
nand U29709 (N_29709,N_26032,N_26245);
nor U29710 (N_29710,N_26837,N_26114);
or U29711 (N_29711,N_27771,N_26848);
and U29712 (N_29712,N_27390,N_26781);
nor U29713 (N_29713,N_27055,N_26191);
nor U29714 (N_29714,N_27504,N_27859);
and U29715 (N_29715,N_26360,N_26458);
or U29716 (N_29716,N_26927,N_27446);
xor U29717 (N_29717,N_26771,N_27398);
nand U29718 (N_29718,N_26432,N_27116);
and U29719 (N_29719,N_26302,N_27639);
nand U29720 (N_29720,N_27666,N_26233);
nor U29721 (N_29721,N_27714,N_26064);
or U29722 (N_29722,N_26451,N_26519);
xnor U29723 (N_29723,N_26271,N_27562);
and U29724 (N_29724,N_26860,N_27479);
nand U29725 (N_29725,N_26693,N_26137);
nand U29726 (N_29726,N_26437,N_27721);
or U29727 (N_29727,N_26723,N_27736);
xor U29728 (N_29728,N_26190,N_27935);
xor U29729 (N_29729,N_27054,N_26362);
or U29730 (N_29730,N_27147,N_26501);
nor U29731 (N_29731,N_26140,N_27332);
nor U29732 (N_29732,N_26862,N_26634);
nand U29733 (N_29733,N_26532,N_26142);
nor U29734 (N_29734,N_27449,N_27017);
and U29735 (N_29735,N_27980,N_27710);
nand U29736 (N_29736,N_27941,N_27100);
and U29737 (N_29737,N_26567,N_27832);
xnor U29738 (N_29738,N_26534,N_27268);
nand U29739 (N_29739,N_26227,N_27044);
xor U29740 (N_29740,N_26386,N_26497);
and U29741 (N_29741,N_26904,N_27337);
and U29742 (N_29742,N_27834,N_27280);
xor U29743 (N_29743,N_26906,N_27585);
or U29744 (N_29744,N_27042,N_27985);
and U29745 (N_29745,N_27614,N_26360);
and U29746 (N_29746,N_26178,N_27861);
xor U29747 (N_29747,N_26686,N_27525);
nor U29748 (N_29748,N_27468,N_26282);
or U29749 (N_29749,N_26705,N_26162);
or U29750 (N_29750,N_27121,N_26193);
nor U29751 (N_29751,N_27802,N_27912);
nand U29752 (N_29752,N_26320,N_26831);
or U29753 (N_29753,N_26680,N_27604);
nand U29754 (N_29754,N_27077,N_26102);
and U29755 (N_29755,N_27964,N_27038);
nand U29756 (N_29756,N_26959,N_26827);
nor U29757 (N_29757,N_27449,N_27731);
xnor U29758 (N_29758,N_27071,N_27981);
nand U29759 (N_29759,N_26571,N_27545);
nor U29760 (N_29760,N_26820,N_26466);
xor U29761 (N_29761,N_27465,N_26793);
xnor U29762 (N_29762,N_26024,N_27545);
or U29763 (N_29763,N_26488,N_27922);
nor U29764 (N_29764,N_26393,N_27259);
xnor U29765 (N_29765,N_26995,N_27906);
nand U29766 (N_29766,N_26307,N_27492);
xor U29767 (N_29767,N_26463,N_27036);
or U29768 (N_29768,N_27105,N_27874);
xnor U29769 (N_29769,N_27630,N_26886);
nand U29770 (N_29770,N_27816,N_26805);
nor U29771 (N_29771,N_26661,N_27322);
xnor U29772 (N_29772,N_26107,N_26051);
and U29773 (N_29773,N_26465,N_27870);
and U29774 (N_29774,N_27477,N_27167);
xor U29775 (N_29775,N_26529,N_26472);
or U29776 (N_29776,N_27512,N_26369);
or U29777 (N_29777,N_27091,N_26479);
nor U29778 (N_29778,N_27427,N_27790);
or U29779 (N_29779,N_26693,N_27471);
xor U29780 (N_29780,N_27115,N_27838);
nor U29781 (N_29781,N_27023,N_27499);
nor U29782 (N_29782,N_26892,N_27148);
and U29783 (N_29783,N_26754,N_27897);
nand U29784 (N_29784,N_27445,N_27091);
nor U29785 (N_29785,N_26429,N_26359);
and U29786 (N_29786,N_26904,N_26226);
nand U29787 (N_29787,N_27960,N_27788);
nand U29788 (N_29788,N_26844,N_27499);
and U29789 (N_29789,N_27238,N_26559);
and U29790 (N_29790,N_26896,N_26526);
nor U29791 (N_29791,N_27606,N_27360);
or U29792 (N_29792,N_26026,N_26184);
nor U29793 (N_29793,N_26313,N_27383);
nand U29794 (N_29794,N_27630,N_26044);
or U29795 (N_29795,N_27613,N_27084);
and U29796 (N_29796,N_27108,N_26936);
xnor U29797 (N_29797,N_26961,N_27661);
xnor U29798 (N_29798,N_27130,N_26546);
nand U29799 (N_29799,N_26812,N_27776);
or U29800 (N_29800,N_26092,N_27005);
nor U29801 (N_29801,N_27996,N_27062);
and U29802 (N_29802,N_26337,N_26552);
nor U29803 (N_29803,N_26423,N_26779);
and U29804 (N_29804,N_26053,N_27090);
nand U29805 (N_29805,N_27468,N_26742);
and U29806 (N_29806,N_26420,N_27584);
and U29807 (N_29807,N_26762,N_27926);
nor U29808 (N_29808,N_26695,N_27244);
and U29809 (N_29809,N_26375,N_27592);
nor U29810 (N_29810,N_26145,N_26565);
and U29811 (N_29811,N_26963,N_26629);
nand U29812 (N_29812,N_27965,N_26045);
or U29813 (N_29813,N_26267,N_26895);
and U29814 (N_29814,N_26338,N_27651);
or U29815 (N_29815,N_27658,N_27961);
xor U29816 (N_29816,N_26042,N_26510);
nand U29817 (N_29817,N_26084,N_27614);
and U29818 (N_29818,N_26089,N_27484);
xnor U29819 (N_29819,N_27244,N_26726);
and U29820 (N_29820,N_26805,N_26202);
xnor U29821 (N_29821,N_26135,N_26499);
or U29822 (N_29822,N_27022,N_27596);
nand U29823 (N_29823,N_27890,N_27241);
nor U29824 (N_29824,N_27735,N_26006);
nor U29825 (N_29825,N_26271,N_26529);
nor U29826 (N_29826,N_26329,N_26723);
or U29827 (N_29827,N_26289,N_27647);
xor U29828 (N_29828,N_26229,N_27615);
or U29829 (N_29829,N_27339,N_26360);
and U29830 (N_29830,N_26346,N_27934);
xor U29831 (N_29831,N_26569,N_27578);
nor U29832 (N_29832,N_27336,N_26290);
nand U29833 (N_29833,N_27417,N_27316);
or U29834 (N_29834,N_27932,N_27603);
or U29835 (N_29835,N_26562,N_27861);
or U29836 (N_29836,N_26384,N_27001);
and U29837 (N_29837,N_27392,N_27227);
or U29838 (N_29838,N_27238,N_27431);
or U29839 (N_29839,N_27016,N_27683);
and U29840 (N_29840,N_26064,N_26998);
nor U29841 (N_29841,N_26434,N_27057);
or U29842 (N_29842,N_27549,N_27968);
or U29843 (N_29843,N_27627,N_26532);
or U29844 (N_29844,N_26738,N_27923);
xor U29845 (N_29845,N_27921,N_26842);
or U29846 (N_29846,N_27120,N_27254);
nor U29847 (N_29847,N_26036,N_27121);
nand U29848 (N_29848,N_27852,N_26979);
xnor U29849 (N_29849,N_27350,N_26368);
or U29850 (N_29850,N_26363,N_27135);
xor U29851 (N_29851,N_26533,N_26296);
or U29852 (N_29852,N_26448,N_27790);
or U29853 (N_29853,N_27780,N_27260);
or U29854 (N_29854,N_27037,N_26188);
nand U29855 (N_29855,N_27312,N_26627);
nor U29856 (N_29856,N_26309,N_27821);
nand U29857 (N_29857,N_27052,N_26474);
xnor U29858 (N_29858,N_26683,N_26087);
or U29859 (N_29859,N_26709,N_27540);
nand U29860 (N_29860,N_27157,N_27707);
nor U29861 (N_29861,N_27461,N_26054);
xnor U29862 (N_29862,N_27128,N_26695);
nor U29863 (N_29863,N_27076,N_27965);
xnor U29864 (N_29864,N_27843,N_27901);
and U29865 (N_29865,N_27611,N_26271);
nand U29866 (N_29866,N_26352,N_26967);
or U29867 (N_29867,N_27564,N_27047);
nand U29868 (N_29868,N_26962,N_27253);
xnor U29869 (N_29869,N_26460,N_26224);
nand U29870 (N_29870,N_27981,N_27946);
nor U29871 (N_29871,N_26208,N_27156);
and U29872 (N_29872,N_26794,N_26378);
and U29873 (N_29873,N_26450,N_27850);
xnor U29874 (N_29874,N_26774,N_26487);
nand U29875 (N_29875,N_27234,N_26338);
nand U29876 (N_29876,N_26361,N_26858);
xnor U29877 (N_29877,N_27686,N_26410);
and U29878 (N_29878,N_27851,N_27223);
and U29879 (N_29879,N_26878,N_26480);
xor U29880 (N_29880,N_27238,N_26301);
and U29881 (N_29881,N_26569,N_27184);
nor U29882 (N_29882,N_26312,N_27678);
and U29883 (N_29883,N_26099,N_26712);
and U29884 (N_29884,N_27761,N_27333);
and U29885 (N_29885,N_27831,N_27262);
nand U29886 (N_29886,N_27199,N_27018);
and U29887 (N_29887,N_27829,N_27090);
nor U29888 (N_29888,N_27820,N_27825);
nor U29889 (N_29889,N_27396,N_27546);
or U29890 (N_29890,N_27001,N_26174);
or U29891 (N_29891,N_27464,N_26006);
or U29892 (N_29892,N_27250,N_26361);
xnor U29893 (N_29893,N_26976,N_27983);
and U29894 (N_29894,N_27772,N_27179);
xor U29895 (N_29895,N_27524,N_27966);
nor U29896 (N_29896,N_26693,N_27669);
or U29897 (N_29897,N_27528,N_27257);
nor U29898 (N_29898,N_26080,N_27599);
nand U29899 (N_29899,N_27140,N_27174);
or U29900 (N_29900,N_27055,N_26484);
nand U29901 (N_29901,N_27554,N_26868);
nor U29902 (N_29902,N_27999,N_27892);
nand U29903 (N_29903,N_26510,N_26997);
or U29904 (N_29904,N_26173,N_26530);
or U29905 (N_29905,N_26242,N_27183);
or U29906 (N_29906,N_26923,N_27545);
and U29907 (N_29907,N_27679,N_26770);
and U29908 (N_29908,N_26477,N_27747);
nand U29909 (N_29909,N_27379,N_26561);
nor U29910 (N_29910,N_26198,N_27379);
or U29911 (N_29911,N_26911,N_26633);
nand U29912 (N_29912,N_27135,N_27802);
nor U29913 (N_29913,N_26893,N_27009);
xor U29914 (N_29914,N_26057,N_27446);
and U29915 (N_29915,N_26452,N_26540);
xor U29916 (N_29916,N_27178,N_26749);
or U29917 (N_29917,N_27484,N_26746);
xnor U29918 (N_29918,N_27909,N_26057);
or U29919 (N_29919,N_27838,N_26391);
nor U29920 (N_29920,N_26119,N_26812);
xnor U29921 (N_29921,N_26054,N_26395);
nand U29922 (N_29922,N_27403,N_26215);
or U29923 (N_29923,N_26524,N_27574);
nand U29924 (N_29924,N_26963,N_27811);
or U29925 (N_29925,N_27088,N_26468);
and U29926 (N_29926,N_26030,N_27267);
and U29927 (N_29927,N_26578,N_27959);
or U29928 (N_29928,N_27752,N_27268);
xnor U29929 (N_29929,N_26564,N_26101);
nand U29930 (N_29930,N_26764,N_27274);
xnor U29931 (N_29931,N_27324,N_26593);
nor U29932 (N_29932,N_26166,N_26794);
or U29933 (N_29933,N_27846,N_26902);
or U29934 (N_29934,N_26353,N_27781);
nor U29935 (N_29935,N_27314,N_27731);
and U29936 (N_29936,N_26215,N_27591);
nor U29937 (N_29937,N_26234,N_27628);
or U29938 (N_29938,N_26191,N_27771);
nand U29939 (N_29939,N_27249,N_26619);
or U29940 (N_29940,N_27919,N_27865);
xor U29941 (N_29941,N_26219,N_27616);
xnor U29942 (N_29942,N_26246,N_26094);
or U29943 (N_29943,N_27444,N_27724);
or U29944 (N_29944,N_27548,N_26033);
nand U29945 (N_29945,N_27032,N_26703);
or U29946 (N_29946,N_27992,N_26803);
or U29947 (N_29947,N_27980,N_27883);
nor U29948 (N_29948,N_27502,N_27624);
xnor U29949 (N_29949,N_26962,N_27409);
and U29950 (N_29950,N_27062,N_27699);
nand U29951 (N_29951,N_26329,N_27506);
xor U29952 (N_29952,N_26928,N_27743);
xor U29953 (N_29953,N_26093,N_26508);
nand U29954 (N_29954,N_27257,N_27230);
and U29955 (N_29955,N_26492,N_27078);
xor U29956 (N_29956,N_26645,N_27182);
nand U29957 (N_29957,N_26962,N_26825);
nand U29958 (N_29958,N_27010,N_27755);
and U29959 (N_29959,N_27524,N_26207);
nor U29960 (N_29960,N_26681,N_26056);
or U29961 (N_29961,N_27357,N_27508);
or U29962 (N_29962,N_26845,N_26560);
nand U29963 (N_29963,N_26288,N_27154);
nor U29964 (N_29964,N_27148,N_27336);
xor U29965 (N_29965,N_27571,N_26890);
and U29966 (N_29966,N_27791,N_26348);
nand U29967 (N_29967,N_27007,N_26445);
and U29968 (N_29968,N_27185,N_26490);
xor U29969 (N_29969,N_27269,N_27645);
xnor U29970 (N_29970,N_26231,N_26511);
xor U29971 (N_29971,N_26127,N_27283);
xnor U29972 (N_29972,N_26836,N_26186);
or U29973 (N_29973,N_27396,N_26125);
or U29974 (N_29974,N_26724,N_27595);
xnor U29975 (N_29975,N_27515,N_27979);
nor U29976 (N_29976,N_27687,N_27989);
nor U29977 (N_29977,N_26796,N_26406);
or U29978 (N_29978,N_26228,N_27253);
or U29979 (N_29979,N_26159,N_26960);
or U29980 (N_29980,N_27771,N_27774);
nand U29981 (N_29981,N_27673,N_27073);
nor U29982 (N_29982,N_27159,N_26231);
nor U29983 (N_29983,N_26664,N_27433);
nor U29984 (N_29984,N_26310,N_27541);
or U29985 (N_29985,N_26844,N_26624);
nor U29986 (N_29986,N_26073,N_27665);
nor U29987 (N_29987,N_26441,N_27603);
nor U29988 (N_29988,N_26568,N_27835);
nand U29989 (N_29989,N_27331,N_26814);
and U29990 (N_29990,N_26772,N_26147);
and U29991 (N_29991,N_26331,N_26851);
or U29992 (N_29992,N_26022,N_27710);
nor U29993 (N_29993,N_26901,N_26686);
nand U29994 (N_29994,N_26178,N_27680);
and U29995 (N_29995,N_27573,N_26804);
xnor U29996 (N_29996,N_27063,N_26484);
or U29997 (N_29997,N_27461,N_26342);
xor U29998 (N_29998,N_26330,N_26910);
and U29999 (N_29999,N_26668,N_26040);
and U30000 (N_30000,N_29776,N_29587);
and U30001 (N_30001,N_28687,N_28526);
nand U30002 (N_30002,N_29270,N_28021);
xor U30003 (N_30003,N_28277,N_28648);
nor U30004 (N_30004,N_28613,N_28897);
and U30005 (N_30005,N_28864,N_29672);
xnor U30006 (N_30006,N_28690,N_28436);
nand U30007 (N_30007,N_29530,N_29262);
nand U30008 (N_30008,N_28343,N_29446);
or U30009 (N_30009,N_29615,N_28312);
nand U30010 (N_30010,N_29766,N_28336);
nor U30011 (N_30011,N_29410,N_29884);
or U30012 (N_30012,N_28699,N_28433);
or U30013 (N_30013,N_29283,N_29735);
or U30014 (N_30014,N_28276,N_28786);
nand U30015 (N_30015,N_29662,N_28210);
or U30016 (N_30016,N_29279,N_28377);
and U30017 (N_30017,N_28647,N_28297);
xor U30018 (N_30018,N_29678,N_29609);
or U30019 (N_30019,N_29496,N_29962);
or U30020 (N_30020,N_28726,N_28386);
nor U30021 (N_30021,N_28176,N_28400);
or U30022 (N_30022,N_29408,N_28670);
xor U30023 (N_30023,N_28351,N_29225);
xnor U30024 (N_30024,N_28104,N_29995);
or U30025 (N_30025,N_28225,N_29327);
nand U30026 (N_30026,N_29689,N_28906);
or U30027 (N_30027,N_29006,N_29764);
xnor U30028 (N_30028,N_28322,N_29429);
and U30029 (N_30029,N_28121,N_29793);
nor U30030 (N_30030,N_28619,N_28829);
xnor U30031 (N_30031,N_29010,N_28468);
nor U30032 (N_30032,N_29625,N_28941);
and U30033 (N_30033,N_28744,N_29065);
nand U30034 (N_30034,N_29636,N_28843);
or U30035 (N_30035,N_29140,N_28541);
and U30036 (N_30036,N_29059,N_28542);
and U30037 (N_30037,N_28175,N_28732);
nor U30038 (N_30038,N_29497,N_28066);
xor U30039 (N_30039,N_28618,N_29513);
and U30040 (N_30040,N_28678,N_29778);
or U30041 (N_30041,N_28862,N_28053);
and U30042 (N_30042,N_29405,N_29382);
and U30043 (N_30043,N_28527,N_29946);
and U30044 (N_30044,N_29618,N_29610);
and U30045 (N_30045,N_28701,N_29545);
and U30046 (N_30046,N_28376,N_28331);
nand U30047 (N_30047,N_28034,N_28500);
or U30048 (N_30048,N_29812,N_29559);
xor U30049 (N_30049,N_28410,N_28092);
or U30050 (N_30050,N_28890,N_28237);
nor U30051 (N_30051,N_28146,N_28991);
xor U30052 (N_30052,N_29244,N_29440);
nor U30053 (N_30053,N_28911,N_29990);
and U30054 (N_30054,N_29451,N_29192);
nor U30055 (N_30055,N_28586,N_29288);
or U30056 (N_30056,N_29874,N_29835);
nor U30057 (N_30057,N_29369,N_28992);
xnor U30058 (N_30058,N_28020,N_29544);
xor U30059 (N_30059,N_29997,N_28965);
nor U30060 (N_30060,N_29677,N_28528);
nor U30061 (N_30061,N_29871,N_29373);
and U30062 (N_30062,N_29450,N_28576);
or U30063 (N_30063,N_29774,N_29794);
nor U30064 (N_30064,N_28651,N_28951);
nor U30065 (N_30065,N_29121,N_29388);
nor U30066 (N_30066,N_28698,N_28620);
nor U30067 (N_30067,N_28616,N_29036);
and U30068 (N_30068,N_28804,N_29500);
and U30069 (N_30069,N_28523,N_29313);
and U30070 (N_30070,N_29744,N_29681);
and U30071 (N_30071,N_28221,N_29414);
or U30072 (N_30072,N_29630,N_29222);
nand U30073 (N_30073,N_28264,N_28043);
xnor U30074 (N_30074,N_28957,N_28011);
nor U30075 (N_30075,N_29576,N_28534);
nor U30076 (N_30076,N_28899,N_28877);
xnor U30077 (N_30077,N_29436,N_28524);
or U30078 (N_30078,N_29475,N_29135);
nand U30079 (N_30079,N_28742,N_28398);
nor U30080 (N_30080,N_28779,N_29391);
xnor U30081 (N_30081,N_28996,N_29887);
xor U30082 (N_30082,N_29643,N_28704);
or U30083 (N_30083,N_29307,N_29113);
nand U30084 (N_30084,N_29593,N_29136);
or U30085 (N_30085,N_29740,N_28999);
nor U30086 (N_30086,N_28590,N_28131);
xor U30087 (N_30087,N_28977,N_28230);
or U30088 (N_30088,N_28054,N_28000);
nand U30089 (N_30089,N_28943,N_29931);
xor U30090 (N_30090,N_28956,N_29782);
xor U30091 (N_30091,N_28925,N_28729);
nor U30092 (N_30092,N_28371,N_29914);
xor U30093 (N_30093,N_29138,N_28674);
nand U30094 (N_30094,N_29196,N_29152);
and U30095 (N_30095,N_28640,N_28617);
nor U30096 (N_30096,N_28988,N_28505);
and U30097 (N_30097,N_28681,N_29855);
nor U30098 (N_30098,N_28115,N_28511);
nand U30099 (N_30099,N_28167,N_29842);
nand U30100 (N_30100,N_29016,N_29597);
nor U30101 (N_30101,N_29772,N_29302);
nand U30102 (N_30102,N_28318,N_29404);
and U30103 (N_30103,N_29329,N_28994);
and U30104 (N_30104,N_29711,N_29721);
or U30105 (N_30105,N_28326,N_29015);
nor U30106 (N_30106,N_28555,N_29599);
or U30107 (N_30107,N_29110,N_29910);
nand U30108 (N_30108,N_29119,N_29312);
nand U30109 (N_30109,N_29868,N_29722);
or U30110 (N_30110,N_28027,N_29582);
nor U30111 (N_30111,N_28472,N_28782);
nand U30112 (N_30112,N_29822,N_28261);
nand U30113 (N_30113,N_29748,N_28350);
and U30114 (N_30114,N_28163,N_29657);
nand U30115 (N_30115,N_29202,N_28208);
xor U30116 (N_30116,N_29737,N_28112);
xor U30117 (N_30117,N_29653,N_29938);
nand U30118 (N_30118,N_29233,N_28224);
or U30119 (N_30119,N_29347,N_29998);
nand U30120 (N_30120,N_28026,N_28735);
xnor U30121 (N_30121,N_28520,N_28970);
and U30122 (N_30122,N_29965,N_28425);
nor U30123 (N_30123,N_28407,N_29558);
nor U30124 (N_30124,N_29453,N_29023);
nand U30125 (N_30125,N_29017,N_29700);
xor U30126 (N_30126,N_28592,N_29590);
and U30127 (N_30127,N_29331,N_28724);
nor U30128 (N_30128,N_29728,N_28588);
nor U30129 (N_30129,N_29183,N_28234);
nor U30130 (N_30130,N_28900,N_29889);
xor U30131 (N_30131,N_28033,N_29758);
xor U30132 (N_30132,N_28861,N_29201);
and U30133 (N_30133,N_29349,N_29725);
nor U30134 (N_30134,N_28204,N_28283);
nand U30135 (N_30135,N_28579,N_28253);
and U30136 (N_30136,N_29668,N_29033);
nand U30137 (N_30137,N_29466,N_28295);
or U30138 (N_30138,N_28789,N_29102);
xnor U30139 (N_30139,N_29571,N_28244);
and U30140 (N_30140,N_29512,N_29295);
and U30141 (N_30141,N_28095,N_29546);
xor U30142 (N_30142,N_28537,N_29528);
nand U30143 (N_30143,N_28978,N_29939);
xor U30144 (N_30144,N_28337,N_29894);
nor U30145 (N_30145,N_28335,N_29480);
nor U30146 (N_30146,N_29134,N_29975);
nand U30147 (N_30147,N_28898,N_28573);
and U30148 (N_30148,N_28867,N_28869);
and U30149 (N_30149,N_28814,N_29375);
xnor U30150 (N_30150,N_28076,N_29370);
nand U30151 (N_30151,N_29114,N_28580);
xnor U30152 (N_30152,N_29223,N_29490);
xor U30153 (N_30153,N_28258,N_28438);
nor U30154 (N_30154,N_28418,N_29959);
or U30155 (N_30155,N_28111,N_29961);
and U30156 (N_30156,N_29434,N_29338);
xor U30157 (N_30157,N_29981,N_29991);
and U30158 (N_30158,N_28117,N_28968);
nor U30159 (N_30159,N_28915,N_29292);
xor U30160 (N_30160,N_28695,N_28952);
and U30161 (N_30161,N_29577,N_28480);
nor U30162 (N_30162,N_28945,N_29923);
or U30163 (N_30163,N_28649,N_28046);
xor U30164 (N_30164,N_28139,N_28296);
xnor U30165 (N_30165,N_29235,N_28305);
and U30166 (N_30166,N_29316,N_28625);
xor U30167 (N_30167,N_29780,N_28487);
xnor U30168 (N_30168,N_28160,N_29692);
or U30169 (N_30169,N_28199,N_29832);
nor U30170 (N_30170,N_29260,N_28345);
xor U30171 (N_30171,N_28072,N_29562);
xnor U30172 (N_30172,N_29258,N_29168);
and U30173 (N_30173,N_28990,N_29541);
nor U30174 (N_30174,N_29853,N_29819);
nor U30175 (N_30175,N_29104,N_29415);
nand U30176 (N_30176,N_28792,N_28203);
and U30177 (N_30177,N_29605,N_29698);
xor U30178 (N_30178,N_29272,N_28554);
and U30179 (N_30179,N_29207,N_28820);
and U30180 (N_30180,N_29483,N_29580);
and U30181 (N_30181,N_29108,N_29730);
xnor U30182 (N_30182,N_28212,N_29515);
xor U30183 (N_30183,N_28668,N_29120);
nand U30184 (N_30184,N_28406,N_29351);
and U30185 (N_30185,N_29775,N_28135);
nand U30186 (N_30186,N_28389,N_29919);
or U30187 (N_30187,N_28215,N_28173);
nor U30188 (N_30188,N_29841,N_29826);
nor U30189 (N_30189,N_28872,N_28071);
xor U30190 (N_30190,N_29458,N_29204);
and U30191 (N_30191,N_29824,N_29200);
nand U30192 (N_30192,N_29642,N_28161);
and U30193 (N_30193,N_29073,N_29374);
nor U30194 (N_30194,N_29718,N_28762);
or U30195 (N_30195,N_29821,N_28508);
nor U30196 (N_30196,N_29090,N_29875);
nand U30197 (N_30197,N_28063,N_28091);
nor U30198 (N_30198,N_28257,N_29701);
and U30199 (N_30199,N_28781,N_28561);
or U30200 (N_30200,N_29960,N_28720);
xor U30201 (N_30201,N_28645,N_28662);
nand U30202 (N_30202,N_28486,N_29484);
nand U30203 (N_30203,N_29825,N_29703);
nand U30204 (N_30204,N_28304,N_29333);
nor U30205 (N_30205,N_29237,N_29989);
or U30206 (N_30206,N_29663,N_29573);
nand U30207 (N_30207,N_28876,N_29680);
nor U30208 (N_30208,N_29257,N_29300);
xnor U30209 (N_30209,N_28439,N_29879);
xor U30210 (N_30210,N_28315,N_29697);
xnor U30211 (N_30211,N_29308,N_28181);
xnor U30212 (N_30212,N_28214,N_29465);
or U30213 (N_30213,N_29569,N_28064);
nand U30214 (N_30214,N_29034,N_29251);
nor U30215 (N_30215,N_28207,N_28078);
nand U30216 (N_30216,N_29175,N_29967);
nand U30217 (N_30217,N_28251,N_28856);
nor U30218 (N_30218,N_29218,N_28341);
or U30219 (N_30219,N_28529,N_29087);
and U30220 (N_30220,N_28910,N_28327);
nand U30221 (N_30221,N_28197,N_28395);
nor U30222 (N_30222,N_28044,N_28416);
nand U30223 (N_30223,N_29238,N_29340);
nor U30224 (N_30224,N_29078,N_29284);
nor U30225 (N_30225,N_29620,N_28597);
and U30226 (N_30226,N_29935,N_28634);
or U30227 (N_30227,N_28007,N_28706);
and U30228 (N_30228,N_29651,N_29430);
nand U30229 (N_30229,N_29655,N_28414);
and U30230 (N_30230,N_28452,N_29658);
nor U30231 (N_30231,N_28552,N_28666);
nand U30232 (N_30232,N_28308,N_28464);
nand U30233 (N_30233,N_29901,N_29427);
and U30234 (N_30234,N_28434,N_29845);
and U30235 (N_30235,N_29971,N_29049);
or U30236 (N_30236,N_28947,N_28714);
xor U30237 (N_30237,N_28495,N_29877);
nor U30238 (N_30238,N_28226,N_28417);
and U30239 (N_30239,N_28822,N_29263);
or U30240 (N_30240,N_28819,N_29491);
nand U30241 (N_30241,N_28928,N_28473);
nor U30242 (N_30242,N_29153,N_29506);
nor U30243 (N_30243,N_29507,N_29456);
nand U30244 (N_30244,N_28694,N_29792);
and U30245 (N_30245,N_28293,N_28460);
nand U30246 (N_30246,N_29406,N_28703);
and U30247 (N_30247,N_28641,N_29221);
and U30248 (N_30248,N_28094,N_28873);
or U30249 (N_30249,N_28909,N_28477);
xnor U30250 (N_30250,N_28006,N_28231);
or U30251 (N_30251,N_29710,N_28469);
and U30252 (N_30252,N_29656,N_28980);
or U30253 (N_30253,N_29892,N_29171);
nor U30254 (N_30254,N_29984,N_29638);
nor U30255 (N_30255,N_29753,N_28461);
nor U30256 (N_30256,N_29525,N_28858);
or U30257 (N_30257,N_29293,N_29372);
nand U30258 (N_30258,N_28525,N_29085);
and U30259 (N_30259,N_29676,N_28321);
and U30260 (N_30260,N_29008,N_29908);
nor U30261 (N_30261,N_29442,N_29585);
nor U30262 (N_30262,N_29798,N_28466);
and U30263 (N_30263,N_28615,N_28362);
nor U30264 (N_30264,N_28474,N_29359);
or U30265 (N_30265,N_28778,N_28136);
nand U30266 (N_30266,N_28018,N_29531);
nor U30267 (N_30267,N_28841,N_29286);
nand U30268 (N_30268,N_28810,N_28358);
nand U30269 (N_30269,N_28577,N_29188);
xor U30270 (N_30270,N_28894,N_28169);
nor U30271 (N_30271,N_29075,N_28730);
and U30272 (N_30272,N_28828,N_28939);
nor U30273 (N_30273,N_29021,N_29122);
nor U30274 (N_30274,N_29791,N_28973);
xnor U30275 (N_30275,N_29360,N_28278);
or U30276 (N_30276,N_29907,N_28451);
nand U30277 (N_30277,N_28140,N_28935);
nand U30278 (N_30278,N_28959,N_28445);
nand U30279 (N_30279,N_29502,N_29169);
and U30280 (N_30280,N_28752,N_29481);
and U30281 (N_30281,N_29301,N_28549);
nand U30282 (N_30282,N_29335,N_29452);
and U30283 (N_30283,N_28349,N_29886);
xor U30284 (N_30284,N_28252,N_29918);
nor U30285 (N_30285,N_28675,N_29880);
nand U30286 (N_30286,N_29294,N_29371);
xnor U30287 (N_30287,N_28731,N_29448);
or U30288 (N_30288,N_29915,N_29714);
xor U30289 (N_30289,N_28799,N_29147);
nand U30290 (N_30290,N_29176,N_29733);
or U30291 (N_30291,N_28288,N_29786);
xnor U30292 (N_30292,N_28340,N_28557);
or U30293 (N_30293,N_28771,N_28837);
nor U30294 (N_30294,N_29437,N_28008);
and U30295 (N_30295,N_28272,N_28854);
xor U30296 (N_30296,N_29635,N_28891);
nand U30297 (N_30297,N_29649,N_29039);
or U30298 (N_30298,N_29851,N_28403);
xnor U30299 (N_30299,N_29232,N_28476);
or U30300 (N_30300,N_28815,N_29478);
xnor U30301 (N_30301,N_29724,N_28038);
and U30302 (N_30302,N_29505,N_28491);
or U30303 (N_30303,N_28462,N_29071);
xnor U30304 (N_30304,N_29203,N_28096);
and U30305 (N_30305,N_28880,N_28086);
xnor U30306 (N_30306,N_29029,N_29926);
xnor U30307 (N_30307,N_29584,N_28922);
xor U30308 (N_30308,N_29986,N_28133);
and U30309 (N_30309,N_28602,N_28800);
nand U30310 (N_30310,N_29604,N_28702);
or U30311 (N_30311,N_28423,N_28733);
nor U30312 (N_30312,N_29290,N_28926);
nand U30313 (N_30313,N_28187,N_29675);
and U30314 (N_30314,N_29191,N_28598);
nand U30315 (N_30315,N_28982,N_29025);
or U30316 (N_30316,N_29161,N_29905);
xor U30317 (N_30317,N_28431,N_28806);
xor U30318 (N_30318,N_28156,N_28718);
and U30319 (N_30319,N_28188,N_28089);
xor U30320 (N_30320,N_29241,N_29217);
nand U30321 (N_30321,N_28757,N_28656);
and U30322 (N_30322,N_29332,N_28249);
and U30323 (N_30323,N_28429,N_28986);
and U30324 (N_30324,N_29432,N_28369);
or U30325 (N_30325,N_28587,N_29801);
xor U30326 (N_30326,N_28422,N_28964);
nor U30327 (N_30327,N_28332,N_28931);
or U30328 (N_30328,N_28242,N_28784);
or U30329 (N_30329,N_28608,N_29457);
nor U30330 (N_30330,N_29158,N_29588);
and U30331 (N_30331,N_28756,N_29166);
or U30332 (N_30332,N_28193,N_28420);
nand U30333 (N_30333,N_29020,N_29230);
nand U30334 (N_30334,N_29291,N_29930);
and U30335 (N_30335,N_28059,N_28192);
nand U30336 (N_30336,N_29190,N_29616);
or U30337 (N_30337,N_28907,N_28005);
and U30338 (N_30338,N_28798,N_28736);
and U30339 (N_30339,N_29115,N_28844);
nor U30340 (N_30340,N_29704,N_28938);
or U30341 (N_30341,N_28081,N_29142);
xor U30342 (N_30342,N_29389,N_28217);
nand U30343 (N_30343,N_28453,N_28606);
xor U30344 (N_30344,N_29395,N_28213);
xor U30345 (N_30345,N_28067,N_29848);
or U30346 (N_30346,N_29362,N_29355);
or U30347 (N_30347,N_28611,N_29807);
nor U30348 (N_30348,N_28709,N_29210);
xor U30349 (N_30349,N_28504,N_28470);
nand U30350 (N_30350,N_29575,N_28725);
nor U30351 (N_30351,N_29857,N_29354);
or U30352 (N_30352,N_29948,N_28863);
and U30353 (N_30353,N_28412,N_29045);
xor U30354 (N_30354,N_29631,N_28075);
nor U30355 (N_30355,N_29823,N_29240);
nand U30356 (N_30356,N_29149,N_28028);
or U30357 (N_30357,N_28463,N_28574);
or U30358 (N_30358,N_28825,N_29194);
nor U30359 (N_30359,N_29357,N_28239);
nor U30360 (N_30360,N_28785,N_29883);
nand U30361 (N_30361,N_29785,N_29518);
and U30362 (N_30362,N_28220,N_29846);
nand U30363 (N_30363,N_28275,N_29081);
and U30364 (N_30364,N_28818,N_29393);
nand U30365 (N_30365,N_28759,N_28955);
and U30366 (N_30366,N_29834,N_29053);
nor U30367 (N_30367,N_28683,N_29486);
and U30368 (N_30368,N_29925,N_28682);
and U30369 (N_30369,N_28969,N_28428);
or U30370 (N_30370,N_28155,N_29623);
xor U30371 (N_30371,N_28514,N_29399);
xnor U30372 (N_30372,N_29208,N_29271);
nor U30373 (N_30373,N_28179,N_29729);
nand U30374 (N_30374,N_29719,N_28359);
or U30375 (N_30375,N_28878,N_29024);
nor U30376 (N_30376,N_29064,N_28510);
xnor U30377 (N_30377,N_28874,N_29645);
nor U30378 (N_30378,N_29873,N_28077);
and U30379 (N_30379,N_28962,N_28390);
or U30380 (N_30380,N_28855,N_28129);
nand U30381 (N_30381,N_29754,N_28001);
or U30382 (N_30382,N_29337,N_29172);
and U30383 (N_30383,N_28454,N_28022);
or U30384 (N_30384,N_29982,N_28334);
or U30385 (N_30385,N_29330,N_29561);
nand U30386 (N_30386,N_29983,N_28562);
or U30387 (N_30387,N_28811,N_28055);
xor U30388 (N_30388,N_28110,N_28793);
or U30389 (N_30389,N_28328,N_28248);
or U30390 (N_30390,N_29156,N_29159);
xor U30391 (N_30391,N_28605,N_28780);
nand U30392 (N_30392,N_28367,N_28062);
and U30393 (N_30393,N_29003,N_29274);
and U30394 (N_30394,N_29468,N_29072);
nor U30395 (N_30395,N_29574,N_29199);
xnor U30396 (N_30396,N_29077,N_29787);
nor U30397 (N_30397,N_28347,N_28853);
or U30398 (N_30398,N_28488,N_29057);
xor U30399 (N_30399,N_29702,N_29195);
nor U30400 (N_30400,N_28908,N_28817);
nor U30401 (N_30401,N_28109,N_28623);
and U30402 (N_30402,N_28707,N_29379);
nand U30403 (N_30403,N_29963,N_28612);
and U30404 (N_30404,N_28747,N_29570);
xor U30405 (N_30405,N_29250,N_28141);
and U30406 (N_30406,N_29058,N_29428);
xor U30407 (N_30407,N_29304,N_29617);
xnor U30408 (N_30408,N_28513,N_29056);
and U30409 (N_30409,N_29596,N_29184);
xor U30410 (N_30410,N_28556,N_29103);
nand U30411 (N_30411,N_29511,N_29859);
or U30412 (N_30412,N_29671,N_28498);
xnor U30413 (N_30413,N_28457,N_29863);
or U30414 (N_30414,N_29278,N_29581);
nand U30415 (N_30415,N_28809,N_28484);
xor U30416 (N_30416,N_28539,N_28255);
nor U30417 (N_30417,N_29276,N_28560);
nor U30418 (N_30418,N_29236,N_29591);
xor U30419 (N_30419,N_29193,N_28551);
and U30420 (N_30420,N_28478,N_29131);
nor U30421 (N_30421,N_28421,N_28721);
nor U30422 (N_30422,N_28243,N_28449);
nand U30423 (N_30423,N_28961,N_29177);
and U30424 (N_30424,N_29390,N_29298);
and U30425 (N_30425,N_29629,N_28993);
and U30426 (N_30426,N_29876,N_29326);
and U30427 (N_30427,N_29186,N_28794);
or U30428 (N_30428,N_29900,N_29779);
or U30429 (N_30429,N_28069,N_28538);
and U30430 (N_30430,N_29885,N_29137);
and U30431 (N_30431,N_28128,N_29533);
nand U30432 (N_30432,N_28303,N_29896);
or U30433 (N_30433,N_28316,N_28583);
xnor U30434 (N_30434,N_29999,N_29070);
xor U30435 (N_30435,N_28717,N_28045);
xor U30436 (N_30436,N_29245,N_28132);
nor U30437 (N_30437,N_28821,N_29556);
or U30438 (N_30438,N_29867,N_28593);
and U30439 (N_30439,N_29150,N_28205);
nand U30440 (N_30440,N_29957,N_29647);
xnor U30441 (N_30441,N_28233,N_28165);
nor U30442 (N_30442,N_29055,N_29673);
nand U30443 (N_30443,N_29891,N_28715);
and U30444 (N_30444,N_28402,N_29659);
or U30445 (N_30445,N_28665,N_28074);
or U30446 (N_30446,N_29974,N_28535);
nor U30447 (N_30447,N_28924,N_28546);
xnor U30448 (N_30448,N_29943,N_28629);
nor U30449 (N_30449,N_29454,N_28536);
xnor U30450 (N_30450,N_29189,N_28677);
and U30451 (N_30451,N_28388,N_29992);
nand U30452 (N_30452,N_29637,N_28170);
xnor U30453 (N_30453,N_29028,N_29209);
or U30454 (N_30454,N_29564,N_29560);
xor U30455 (N_30455,N_28404,N_29091);
nor U30456 (N_30456,N_28875,N_29685);
or U30457 (N_30457,N_29401,N_29109);
or U30458 (N_30458,N_28937,N_29802);
nand U30459 (N_30459,N_29280,N_28148);
or U30460 (N_30460,N_29309,N_29770);
or U30461 (N_30461,N_29317,N_28851);
xnor U30462 (N_30462,N_29557,N_28361);
nand U30463 (N_30463,N_29828,N_29922);
and U30464 (N_30464,N_28692,N_29985);
and U30465 (N_30465,N_29094,N_29384);
nor U30466 (N_30466,N_28553,N_28314);
and U30467 (N_30467,N_28570,N_28578);
nor U30468 (N_30468,N_28773,N_28201);
nand U30469 (N_30469,N_28627,N_28265);
nand U30470 (N_30470,N_29473,N_29510);
nand U30471 (N_30471,N_28599,N_28979);
and U30472 (N_30472,N_28079,N_29912);
nand U30473 (N_30473,N_29157,N_29380);
nor U30474 (N_30474,N_28300,N_29916);
or U30475 (N_30475,N_29501,N_29829);
and U30476 (N_30476,N_29606,N_29443);
nor U30477 (N_30477,N_28025,N_28440);
xnor U30478 (N_30478,N_28151,N_28659);
or U30479 (N_30479,N_29482,N_29690);
xnor U30480 (N_30480,N_28567,N_28373);
and U30481 (N_30481,N_29259,N_29540);
or U30482 (N_30482,N_28284,N_29987);
nor U30483 (N_30483,N_28370,N_28672);
and U30484 (N_30484,N_29040,N_29743);
or U30485 (N_30485,N_28738,N_28745);
nor U30486 (N_30486,N_29773,N_29937);
nand U30487 (N_30487,N_29958,N_29348);
and U30488 (N_30488,N_28516,N_29862);
nand U30489 (N_30489,N_29589,N_28688);
nor U30490 (N_30490,N_28895,N_28739);
xnor U30491 (N_30491,N_28116,N_28885);
or U30492 (N_30492,N_29022,N_28413);
nand U30493 (N_30493,N_29519,N_28060);
or U30494 (N_30494,N_28705,N_28680);
xor U30495 (N_30495,N_29164,N_29143);
nor U30496 (N_30496,N_28492,N_28219);
xor U30497 (N_30497,N_29368,N_29322);
nor U30498 (N_30498,N_29048,N_29079);
and U30499 (N_30499,N_29767,N_28519);
or U30500 (N_30500,N_29532,N_29350);
nor U30501 (N_30501,N_29578,N_28240);
or U30502 (N_30502,N_28879,N_29394);
or U30503 (N_30503,N_28805,N_29459);
nor U30504 (N_30504,N_29341,N_28051);
or U30505 (N_30505,N_28262,N_28375);
xor U30506 (N_30506,N_28235,N_29179);
xnor U30507 (N_30507,N_28522,N_28712);
nand U30508 (N_30508,N_29398,N_29165);
and U30509 (N_30509,N_28636,N_29433);
xor U30510 (N_30510,N_28016,N_29539);
and U30511 (N_30511,N_28285,N_29083);
nand U30512 (N_30512,N_28566,N_29601);
nand U30513 (N_30513,N_29383,N_28381);
nor U30514 (N_30514,N_28787,N_29594);
or U30515 (N_30515,N_28585,N_28352);
nor U30516 (N_30516,N_28643,N_29691);
xor U30517 (N_30517,N_29650,N_29069);
and U30518 (N_30518,N_28178,N_29185);
nand U30519 (N_30519,N_28775,N_28975);
or U30520 (N_30520,N_28184,N_29795);
and U30521 (N_30521,N_29757,N_29460);
xor U30522 (N_30522,N_29552,N_28405);
and U30523 (N_30523,N_28056,N_28684);
and U30524 (N_30524,N_29682,N_29723);
nand U30525 (N_30525,N_28642,N_29132);
or U30526 (N_30526,N_28569,N_29750);
nand U30527 (N_30527,N_28443,N_28273);
or U30528 (N_30528,N_28090,N_29878);
xor U30529 (N_30529,N_28143,N_28385);
xnor U30530 (N_30530,N_28030,N_28147);
and U30531 (N_30531,N_29426,N_29044);
nor U30532 (N_30532,N_28600,N_28097);
nand U30533 (N_30533,N_28465,N_29032);
and U30534 (N_30534,N_28323,N_29941);
nand U30535 (N_30535,N_28048,N_29756);
nor U30536 (N_30536,N_28686,N_29396);
xor U30537 (N_30537,N_28357,N_28889);
or U30538 (N_30538,N_29129,N_29897);
and U30539 (N_30539,N_29139,N_28250);
and U30540 (N_30540,N_29227,N_28543);
or U30541 (N_30541,N_28896,N_28189);
nor U30542 (N_30542,N_29479,N_29683);
xor U30543 (N_30543,N_28737,N_29813);
nand U30544 (N_30544,N_29872,N_28150);
nand U30545 (N_30545,N_29717,N_28456);
nor U30546 (N_30546,N_28444,N_28307);
nor U30547 (N_30547,N_28353,N_29524);
and U30548 (N_30548,N_28741,N_29097);
and U30549 (N_30549,N_29765,N_28946);
xnor U30550 (N_30550,N_28263,N_28247);
or U30551 (N_30551,N_29281,N_29082);
nor U30552 (N_30552,N_29843,N_28236);
nand U30553 (N_30553,N_28036,N_29741);
or U30554 (N_30554,N_28292,N_28628);
nor U30555 (N_30555,N_29864,N_29840);
or U30556 (N_30556,N_29760,N_28790);
nor U30557 (N_30557,N_29799,N_28144);
nor U30558 (N_30558,N_28471,N_29462);
and U30559 (N_30559,N_28164,N_28545);
nor U30560 (N_30560,N_28073,N_28483);
nand U30561 (N_30561,N_28040,N_29932);
xnor U30562 (N_30562,N_28995,N_29839);
or U30563 (N_30563,N_28696,N_29904);
or U30564 (N_30564,N_28758,N_29365);
or U30565 (N_30565,N_29543,N_28974);
xnor U30566 (N_30566,N_29838,N_29198);
nor U30567 (N_30567,N_29535,N_28037);
xnor U30568 (N_30568,N_28766,N_29043);
nor U30569 (N_30569,N_28106,N_29567);
nor U30570 (N_30570,N_29027,N_28245);
or U30571 (N_30571,N_29303,N_29167);
nand U30572 (N_30572,N_29893,N_29988);
nand U30573 (N_30573,N_28882,N_28691);
nand U30574 (N_30574,N_28227,N_29956);
nand U30575 (N_30575,N_28654,N_29376);
nand U30576 (N_30576,N_29220,N_28166);
xor U30577 (N_30577,N_28664,N_29516);
and U30578 (N_30578,N_28499,N_28568);
and U30579 (N_30579,N_29861,N_28259);
nor U30580 (N_30580,N_29624,N_29612);
xor U30581 (N_30581,N_29417,N_28154);
or U30582 (N_30582,N_28653,N_28824);
nand U30583 (N_30583,N_28269,N_29890);
nand U30584 (N_30584,N_29523,N_28796);
nand U30585 (N_30585,N_28004,N_28497);
xor U30586 (N_30586,N_29555,N_29269);
xnor U30587 (N_30587,N_28835,N_29738);
xor U30588 (N_30588,N_28228,N_28533);
nand U30589 (N_30589,N_29709,N_28320);
xnor U30590 (N_30590,N_28325,N_28865);
nand U30591 (N_30591,N_28830,N_29949);
or U30592 (N_30592,N_29749,N_29924);
nor U30593 (N_30593,N_28396,N_29726);
nand U30594 (N_30594,N_28881,N_29499);
nor U30595 (N_30595,N_29005,N_29127);
nand U30596 (N_30596,N_29699,N_29996);
or U30597 (N_30597,N_29854,N_29945);
xnor U30598 (N_30598,N_29229,N_29447);
nor U30599 (N_30599,N_28658,N_29224);
xnor U30600 (N_30600,N_28087,N_29409);
or U30601 (N_30601,N_29211,N_28774);
and U30602 (N_30602,N_28260,N_28019);
and U30603 (N_30603,N_29031,N_29144);
xor U30604 (N_30604,N_28107,N_28042);
xnor U30605 (N_30605,N_29130,N_29494);
nand U30606 (N_30606,N_29148,N_28838);
nor U30607 (N_30607,N_28339,N_28013);
or U30608 (N_30608,N_29856,N_28816);
xor U30609 (N_30609,N_29181,N_29378);
or U30610 (N_30610,N_28860,N_28981);
and U30611 (N_30611,N_29219,N_28765);
and U30612 (N_30612,N_29820,N_29522);
nand U30613 (N_30613,N_28857,N_29187);
nand U30614 (N_30614,N_28082,N_29969);
nand U30615 (N_30615,N_29425,N_29009);
nor U30616 (N_30616,N_28009,N_29377);
or U30617 (N_30617,N_29627,N_29315);
nand U30618 (N_30618,N_29979,N_28223);
nand U30619 (N_30619,N_28813,N_28984);
or U30620 (N_30620,N_29583,N_28014);
nand U30621 (N_30621,N_29007,N_28850);
nand U30622 (N_30622,N_29954,N_28581);
and U30623 (N_30623,N_28174,N_28382);
nand U30624 (N_30624,N_28502,N_29439);
nor U30625 (N_30625,N_28333,N_28041);
or U30626 (N_30626,N_28650,N_29716);
or U30627 (N_30627,N_28254,N_28971);
and U30628 (N_30628,N_28031,N_29572);
and U30629 (N_30629,N_28002,N_29755);
or U30630 (N_30630,N_29881,N_28409);
or U30631 (N_30631,N_28595,N_28485);
and U30632 (N_30632,N_29063,N_29955);
xor U30633 (N_30633,N_29903,N_29936);
and U30634 (N_30634,N_28558,N_29554);
nor U30635 (N_30635,N_28419,N_28290);
nor U30636 (N_30636,N_28610,N_29520);
and U30637 (N_30637,N_29062,N_29118);
nor U30638 (N_30638,N_29666,N_29869);
nand U30639 (N_30639,N_29215,N_29266);
or U30640 (N_30640,N_29768,N_28185);
nand U30641 (N_30641,N_29632,N_28503);
nand U30642 (N_30642,N_28088,N_28392);
nor U30643 (N_30643,N_28142,N_28447);
and U30644 (N_30644,N_28768,N_29226);
nand U30645 (N_30645,N_28289,N_28070);
or U30646 (N_30646,N_28515,N_28944);
or U30647 (N_30647,N_28017,N_28200);
nor U30648 (N_30648,N_29469,N_28202);
or U30649 (N_30649,N_28826,N_29088);
nand U30650 (N_30650,N_29622,N_29781);
nor U30651 (N_30651,N_28776,N_28271);
nand U30652 (N_30652,N_28827,N_29387);
and U30653 (N_30653,N_28622,N_29012);
or U30654 (N_30654,N_29212,N_29947);
nand U30655 (N_30655,N_28356,N_28518);
xor U30656 (N_30656,N_28049,N_29099);
or U30657 (N_30657,N_28479,N_29254);
nor U30658 (N_30658,N_29253,N_29827);
xnor U30659 (N_30659,N_29579,N_29777);
xnor U30660 (N_30660,N_29669,N_29865);
and U30661 (N_30661,N_29463,N_29117);
nor U30662 (N_30662,N_29051,N_29246);
and U30663 (N_30663,N_28563,N_29763);
xnor U30664 (N_30664,N_29514,N_28697);
nor U30665 (N_30665,N_29654,N_28904);
or U30666 (N_30666,N_29921,N_28113);
nor U30667 (N_30667,N_29731,N_29407);
or U30668 (N_30668,N_28750,N_29180);
nand U30669 (N_30669,N_28932,N_28966);
or U30670 (N_30670,N_29679,N_28933);
nand U30671 (N_30671,N_28099,N_28669);
and U30672 (N_30672,N_28481,N_29353);
xnor U30673 (N_30673,N_29477,N_28050);
and U30674 (N_30674,N_28032,N_29361);
or U30675 (N_30675,N_29899,N_29105);
nor U30676 (N_30676,N_28761,N_28366);
xnor U30677 (N_30677,N_29684,N_28490);
nor U30678 (N_30678,N_28842,N_28626);
xor U30679 (N_30679,N_28716,N_29818);
nand U30680 (N_30680,N_29068,N_28916);
and U30681 (N_30681,N_28760,N_28108);
and U30682 (N_30682,N_29687,N_29600);
or U30683 (N_30683,N_28211,N_28102);
nand U30684 (N_30684,N_28727,N_29247);
or U30685 (N_30685,N_29870,N_28949);
xnor U30686 (N_30686,N_29381,N_29934);
nor U30687 (N_30687,N_28609,N_29004);
and U30688 (N_30688,N_29472,N_28427);
and U30689 (N_30689,N_29444,N_28084);
and U30690 (N_30690,N_29548,N_28145);
nand U30691 (N_30691,N_28571,N_28646);
xor U30692 (N_30692,N_28159,N_29906);
nand U30693 (N_30693,N_28644,N_29951);
and U30694 (N_30694,N_29141,N_28719);
xor U30695 (N_30695,N_29013,N_28130);
nor U30696 (N_30696,N_29325,N_29736);
or U30697 (N_30697,N_29563,N_28103);
or U30698 (N_30698,N_29050,N_29849);
or U30699 (N_30699,N_28229,N_28216);
or U30700 (N_30700,N_29001,N_28118);
nand U30701 (N_30701,N_29809,N_28845);
or U30702 (N_30702,N_28918,N_28364);
xnor U30703 (N_30703,N_28936,N_29641);
nand U30704 (N_30704,N_28530,N_28997);
xor U30705 (N_30705,N_29282,N_29422);
xnor U30706 (N_30706,N_29116,N_28512);
xor U30707 (N_30707,N_29553,N_28194);
xor U30708 (N_30708,N_29566,N_29242);
nand U30709 (N_30709,N_28755,N_28455);
xor U30710 (N_30710,N_29762,N_28689);
or U30711 (N_30711,N_29431,N_29107);
or U30712 (N_30712,N_28840,N_28190);
nor U30713 (N_30713,N_29860,N_29608);
nand U30714 (N_30714,N_28280,N_28496);
or U30715 (N_30715,N_29850,N_29445);
nor U30716 (N_30716,N_28550,N_29614);
nand U30717 (N_30717,N_29968,N_28122);
or U30718 (N_30718,N_28589,N_29476);
nand U30719 (N_30719,N_29492,N_28630);
and U30720 (N_30720,N_28065,N_29953);
and U30721 (N_30721,N_28521,N_28638);
and U30722 (N_30722,N_28080,N_29311);
nand U30723 (N_30723,N_29000,N_28948);
nand U30724 (N_30724,N_29328,N_29154);
nor U30725 (N_30725,N_29994,N_28859);
nor U30726 (N_30726,N_28158,N_29461);
and U30727 (N_30727,N_28888,N_28886);
nand U30728 (N_30728,N_29306,N_28346);
xor U30729 (N_30729,N_29742,N_29917);
or U30730 (N_30730,N_29550,N_28138);
xnor U30731 (N_30731,N_29814,N_28673);
and U30732 (N_30732,N_28544,N_28105);
nand U30733 (N_30733,N_29493,N_29804);
xor U30734 (N_30734,N_29667,N_29323);
nand U30735 (N_30735,N_28934,N_29706);
nor U30736 (N_30736,N_29435,N_28268);
nor U30737 (N_30737,N_29978,N_29633);
nor U30738 (N_30738,N_29611,N_29902);
xnor U30739 (N_30739,N_28921,N_28360);
and U30740 (N_30740,N_29321,N_29252);
nor U30741 (N_30741,N_28963,N_28061);
nand U30742 (N_30742,N_29940,N_29086);
nand U30743 (N_30743,N_29400,N_29898);
xnor U30744 (N_30744,N_29162,N_28430);
nand U30745 (N_30745,N_29670,N_29054);
or U30746 (N_30746,N_29112,N_28930);
or U30747 (N_30747,N_29509,N_28344);
nor U30748 (N_30748,N_28424,N_28772);
xor U30749 (N_30749,N_28124,N_28363);
nor U30750 (N_30750,N_29640,N_29866);
xnor U30751 (N_30751,N_29837,N_29950);
nor U30752 (N_30752,N_29784,N_28489);
nor U30753 (N_30753,N_28989,N_28432);
xor U30754 (N_30754,N_29299,N_29942);
nor U30755 (N_30755,N_28125,N_29026);
or U30756 (N_30756,N_28126,N_29123);
and U30757 (N_30757,N_28802,N_29002);
and U30758 (N_30758,N_29747,N_29052);
nand U30759 (N_30759,N_28068,N_28196);
xor U30760 (N_30760,N_29273,N_29076);
or U30761 (N_30761,N_28209,N_29011);
xor U30762 (N_30762,N_29660,N_28833);
and U30763 (N_30763,N_28532,N_29037);
xnor U30764 (N_30764,N_29789,N_28299);
nor U30765 (N_30765,N_28100,N_29810);
nand U30766 (N_30766,N_29534,N_28372);
nand U30767 (N_30767,N_28506,N_28329);
or U30768 (N_30768,N_29928,N_29030);
nor U30769 (N_30769,N_28603,N_29441);
xor U30770 (N_30770,N_28808,N_29909);
nand U30771 (N_30771,N_28852,N_29602);
nor U30772 (N_30772,N_28575,N_29549);
xnor U30773 (N_30773,N_29106,N_28313);
and U30774 (N_30774,N_29745,N_29538);
or U30775 (N_30775,N_29089,N_29146);
nand U30776 (N_30776,N_28746,N_28940);
nand U30777 (N_30777,N_29504,N_28448);
and U30778 (N_30778,N_29586,N_29708);
nand U30779 (N_30779,N_28442,N_29019);
xor U30780 (N_30780,N_28942,N_29715);
and U30781 (N_30781,N_29844,N_29339);
nand U30782 (N_30782,N_28378,N_29438);
xnor U30783 (N_30783,N_29385,N_28348);
or U30784 (N_30784,N_28632,N_28493);
nor U30785 (N_30785,N_28324,N_28058);
nor U30786 (N_30786,N_29858,N_28435);
nor U30787 (N_30787,N_29095,N_29320);
nand U30788 (N_30788,N_28770,N_28401);
xor U30789 (N_30789,N_29619,N_28301);
nand U30790 (N_30790,N_28238,N_29264);
or U30791 (N_30791,N_29093,N_29489);
and U30792 (N_30792,N_29173,N_29096);
nand U30793 (N_30793,N_29261,N_28191);
nor U30794 (N_30794,N_29920,N_28083);
nor U30795 (N_30795,N_29933,N_28241);
and U30796 (N_30796,N_28823,N_29334);
and U30797 (N_30797,N_28098,N_28355);
xnor U30798 (N_30798,N_29100,N_29688);
or U30799 (N_30799,N_28003,N_28270);
and U30800 (N_30800,N_28591,N_28958);
or U30801 (N_30801,N_28180,N_29346);
and U30802 (N_30802,N_29830,N_29972);
xor U30803 (N_30803,N_28029,N_29363);
or U30804 (N_30804,N_29206,N_29613);
nand U30805 (N_30805,N_29145,N_29713);
nor U30806 (N_30806,N_28246,N_29358);
nand U30807 (N_30807,N_29205,N_29817);
nand U30808 (N_30808,N_28795,N_28172);
and U30809 (N_30809,N_28222,N_28769);
nand U30810 (N_30810,N_28903,N_29014);
or U30811 (N_30811,N_29595,N_28868);
and U30812 (N_30812,N_28572,N_29216);
nor U30813 (N_30813,N_29806,N_29536);
nand U30814 (N_30814,N_28950,N_28713);
xnor U30815 (N_30815,N_29803,N_29485);
xnor U30816 (N_30816,N_29098,N_29503);
nor U30817 (N_30817,N_29927,N_28010);
nand U30818 (N_30818,N_29178,N_28655);
nor U30819 (N_30819,N_29314,N_28330);
xor U30820 (N_30820,N_29759,N_28657);
nor U30821 (N_30821,N_28803,N_29977);
nand U30822 (N_30822,N_28475,N_29498);
and U30823 (N_30823,N_28415,N_29344);
nand U30824 (N_30824,N_29343,N_28848);
or U30825 (N_30825,N_29761,N_29796);
nand U30826 (N_30826,N_29607,N_29970);
or U30827 (N_30827,N_29707,N_28920);
and U30828 (N_30828,N_28437,N_29603);
or U30829 (N_30829,N_29913,N_28287);
nand U30830 (N_30830,N_29424,N_29296);
xnor U30831 (N_30831,N_28866,N_29508);
xnor U30832 (N_30832,N_28559,N_29345);
and U30833 (N_30833,N_29626,N_29277);
and U30834 (N_30834,N_28338,N_28887);
nor U30835 (N_30835,N_28596,N_28291);
and U30836 (N_30836,N_28846,N_29686);
nand U30837 (N_30837,N_28614,N_28834);
nand U30838 (N_30838,N_28047,N_29418);
or U30839 (N_30839,N_28374,N_29243);
nor U30840 (N_30840,N_29474,N_29833);
or U30841 (N_30841,N_29598,N_29976);
or U30842 (N_30842,N_28847,N_29980);
and U30843 (N_30843,N_28983,N_28749);
xor U30844 (N_30844,N_28954,N_29771);
and U30845 (N_30845,N_29836,N_29412);
nand U30846 (N_30846,N_28849,N_28302);
nor U30847 (N_30847,N_29287,N_28700);
nand U30848 (N_30848,N_29170,N_29751);
and U30849 (N_30849,N_28494,N_29882);
xor U30850 (N_30850,N_28604,N_29526);
and U30851 (N_30851,N_28411,N_29366);
nor U30852 (N_30852,N_28801,N_28317);
or U30853 (N_30853,N_29592,N_29783);
nor U30854 (N_30854,N_29694,N_28788);
and U30855 (N_30855,N_29471,N_29182);
nand U30856 (N_30856,N_29752,N_28310);
and U30857 (N_30857,N_29495,N_29467);
nand U30858 (N_30858,N_28384,N_29364);
or U30859 (N_30859,N_29419,N_29808);
or U30860 (N_30860,N_29423,N_29035);
or U30861 (N_30861,N_28279,N_28182);
or U30862 (N_30862,N_28426,N_29815);
or U30863 (N_30863,N_28153,N_29788);
nor U30864 (N_30864,N_28601,N_28391);
and U30865 (N_30865,N_29712,N_29018);
and U30866 (N_30866,N_29769,N_29060);
nand U30867 (N_30867,N_29285,N_29464);
nor U30868 (N_30868,N_29228,N_29811);
xnor U30869 (N_30869,N_28267,N_28342);
nand U30870 (N_30870,N_28157,N_28913);
or U30871 (N_30871,N_29739,N_28286);
or U30872 (N_30872,N_29944,N_29816);
nand U30873 (N_30873,N_28232,N_29852);
nand U30874 (N_30874,N_28186,N_29041);
or U30875 (N_30875,N_28871,N_28976);
or U30876 (N_30876,N_29929,N_28183);
xor U30877 (N_30877,N_28306,N_29319);
nand U30878 (N_30878,N_29042,N_28408);
nor U30879 (N_30879,N_29805,N_29973);
nand U30880 (N_30880,N_28914,N_29646);
nor U30881 (N_30881,N_28507,N_28917);
nand U30882 (N_30882,N_28763,N_29746);
nor U30883 (N_30883,N_28274,N_28972);
nor U30884 (N_30884,N_28728,N_29797);
xor U30885 (N_30885,N_28753,N_29342);
nor U30886 (N_30886,N_29084,N_28902);
or U30887 (N_30887,N_28998,N_28685);
and U30888 (N_30888,N_28093,N_29111);
xor U30889 (N_30889,N_28901,N_28256);
and U30890 (N_30890,N_29255,N_28266);
and U30891 (N_30891,N_29403,N_28905);
nor U30892 (N_30892,N_29537,N_28927);
nor U30893 (N_30893,N_28171,N_28387);
or U30894 (N_30894,N_29413,N_29074);
xnor U30895 (N_30895,N_29634,N_29648);
or U30896 (N_30896,N_28639,N_29966);
nand U30897 (N_30897,N_29066,N_29397);
or U30898 (N_30898,N_28621,N_28206);
nor U30899 (N_30899,N_29644,N_29197);
or U30900 (N_30900,N_29542,N_28710);
or U30901 (N_30901,N_28777,N_29449);
nor U30902 (N_30902,N_28134,N_29067);
nor U30903 (N_30903,N_29275,N_28711);
nor U30904 (N_30904,N_28149,N_29310);
and U30905 (N_30905,N_28754,N_29800);
nand U30906 (N_30906,N_28052,N_28311);
nand U30907 (N_30907,N_28564,N_28635);
xor U30908 (N_30908,N_28399,N_28024);
xor U30909 (N_30909,N_29367,N_29174);
xor U30910 (N_30910,N_28831,N_28743);
and U30911 (N_30911,N_28633,N_29487);
nand U30912 (N_30912,N_29402,N_28354);
xnor U30913 (N_30913,N_28547,N_28137);
nand U30914 (N_30914,N_28797,N_28368);
nand U30915 (N_30915,N_28531,N_29517);
and U30916 (N_30916,N_28751,N_29734);
xor U30917 (N_30917,N_28953,N_28594);
xor U30918 (N_30918,N_28023,N_29046);
and U30919 (N_30919,N_28807,N_28467);
or U30920 (N_30920,N_28929,N_29124);
xnor U30921 (N_30921,N_28085,N_29336);
nor U30922 (N_30922,N_29133,N_29665);
xnor U30923 (N_30923,N_28120,N_29911);
and U30924 (N_30924,N_28919,N_28517);
xnor U30925 (N_30925,N_28282,N_29061);
or U30926 (N_30926,N_28832,N_28836);
xnor U30927 (N_30927,N_29421,N_29831);
xor U30928 (N_30928,N_29038,N_28114);
or U30929 (N_30929,N_28893,N_28458);
xnor U30930 (N_30930,N_29790,N_29151);
and U30931 (N_30931,N_29727,N_28394);
and U30932 (N_30932,N_28892,N_28884);
nor U30933 (N_30933,N_28035,N_28380);
and U30934 (N_30934,N_29267,N_29214);
nand U30935 (N_30935,N_28624,N_29318);
or U30936 (N_30936,N_29993,N_29297);
or U30937 (N_30937,N_28152,N_29527);
or U30938 (N_30938,N_28127,N_28584);
nor U30939 (N_30939,N_28967,N_28168);
or U30940 (N_30940,N_28459,N_29488);
and U30941 (N_30941,N_28565,N_28661);
xor U30942 (N_30942,N_28723,N_28708);
and U30943 (N_30943,N_28195,N_29628);
or U30944 (N_30944,N_28667,N_28218);
and U30945 (N_30945,N_29289,N_28582);
and U30946 (N_30946,N_28482,N_28309);
xor U30947 (N_30947,N_28734,N_28839);
nor U30948 (N_30948,N_28101,N_28548);
or U30949 (N_30949,N_28660,N_29248);
xnor U30950 (N_30950,N_29411,N_28379);
nor U30951 (N_30951,N_28365,N_29047);
and U30952 (N_30952,N_29231,N_29356);
and U30953 (N_30953,N_28923,N_29239);
and U30954 (N_30954,N_29234,N_29249);
nor U30955 (N_30955,N_28123,N_29952);
xnor U30956 (N_30956,N_28671,N_29416);
or U30957 (N_30957,N_28281,N_28509);
nor U30958 (N_30958,N_28607,N_29268);
or U30959 (N_30959,N_28679,N_28012);
nor U30960 (N_30960,N_29092,N_28631);
and U30961 (N_30961,N_29847,N_28870);
and U30962 (N_30962,N_29888,N_29256);
and U30963 (N_30963,N_28791,N_29125);
or U30964 (N_30964,N_29101,N_29213);
and U30965 (N_30965,N_29392,N_29732);
xnor U30966 (N_30966,N_29521,N_29324);
xnor U30967 (N_30967,N_28039,N_28294);
and U30968 (N_30968,N_28912,N_29160);
xor U30969 (N_30969,N_29964,N_29155);
nand U30970 (N_30970,N_28198,N_28397);
nor U30971 (N_30971,N_29695,N_28663);
xnor U30972 (N_30972,N_28177,N_29305);
nand U30973 (N_30973,N_29265,N_28319);
or U30974 (N_30974,N_28383,N_29565);
nand U30975 (N_30975,N_29720,N_29674);
nand U30976 (N_30976,N_29621,N_29664);
xor U30977 (N_30977,N_28676,N_29547);
and U30978 (N_30978,N_28987,N_28162);
and U30979 (N_30979,N_29455,N_29568);
or U30980 (N_30980,N_28015,N_29386);
or U30981 (N_30981,N_28501,N_28740);
or U30982 (N_30982,N_28693,N_28540);
nor U30983 (N_30983,N_29080,N_29163);
nand U30984 (N_30984,N_28652,N_28441);
or U30985 (N_30985,N_29895,N_29529);
nand U30986 (N_30986,N_28119,N_29639);
nand U30987 (N_30987,N_28748,N_29693);
or U30988 (N_30988,N_28783,N_28393);
and U30989 (N_30989,N_29652,N_28057);
and U30990 (N_30990,N_29126,N_28450);
nand U30991 (N_30991,N_28985,N_28722);
and U30992 (N_30992,N_29352,N_28960);
or U30993 (N_30993,N_29420,N_29705);
or U30994 (N_30994,N_28764,N_29661);
or U30995 (N_30995,N_29696,N_29551);
and U30996 (N_30996,N_28637,N_29470);
or U30997 (N_30997,N_28767,N_28812);
and U30998 (N_30998,N_28446,N_29128);
or U30999 (N_30999,N_28298,N_28883);
nor U31000 (N_31000,N_28985,N_29079);
and U31001 (N_31001,N_28632,N_28828);
xor U31002 (N_31002,N_29919,N_29581);
nor U31003 (N_31003,N_29549,N_28343);
nand U31004 (N_31004,N_28623,N_28487);
nand U31005 (N_31005,N_28475,N_29930);
xnor U31006 (N_31006,N_29225,N_29312);
or U31007 (N_31007,N_28840,N_29720);
nor U31008 (N_31008,N_28147,N_29990);
and U31009 (N_31009,N_28704,N_29382);
xor U31010 (N_31010,N_28790,N_29362);
and U31011 (N_31011,N_28853,N_29949);
or U31012 (N_31012,N_29154,N_28890);
or U31013 (N_31013,N_29507,N_29399);
and U31014 (N_31014,N_29657,N_29663);
xnor U31015 (N_31015,N_29666,N_28526);
nor U31016 (N_31016,N_29148,N_28203);
or U31017 (N_31017,N_29432,N_28063);
nor U31018 (N_31018,N_28151,N_29967);
and U31019 (N_31019,N_28701,N_29304);
or U31020 (N_31020,N_28027,N_28523);
or U31021 (N_31021,N_28736,N_28903);
nor U31022 (N_31022,N_28061,N_28707);
xnor U31023 (N_31023,N_28947,N_28375);
and U31024 (N_31024,N_28150,N_29792);
and U31025 (N_31025,N_28464,N_29781);
xor U31026 (N_31026,N_28136,N_28129);
nand U31027 (N_31027,N_28581,N_29373);
xor U31028 (N_31028,N_28853,N_28362);
nand U31029 (N_31029,N_28566,N_29906);
or U31030 (N_31030,N_29516,N_28010);
or U31031 (N_31031,N_29361,N_28771);
nand U31032 (N_31032,N_28108,N_28074);
xor U31033 (N_31033,N_28901,N_28683);
and U31034 (N_31034,N_28032,N_29675);
or U31035 (N_31035,N_29309,N_29134);
nor U31036 (N_31036,N_29853,N_29396);
xor U31037 (N_31037,N_29086,N_29826);
and U31038 (N_31038,N_28259,N_29025);
nand U31039 (N_31039,N_29012,N_28944);
xnor U31040 (N_31040,N_29471,N_29773);
and U31041 (N_31041,N_29332,N_28791);
or U31042 (N_31042,N_28211,N_29526);
xor U31043 (N_31043,N_29215,N_28499);
nand U31044 (N_31044,N_29807,N_29542);
or U31045 (N_31045,N_28378,N_28904);
xor U31046 (N_31046,N_29843,N_29336);
or U31047 (N_31047,N_29125,N_28304);
nand U31048 (N_31048,N_29150,N_28800);
or U31049 (N_31049,N_29089,N_29481);
nand U31050 (N_31050,N_29488,N_29201);
or U31051 (N_31051,N_28705,N_28644);
xor U31052 (N_31052,N_28437,N_29819);
nand U31053 (N_31053,N_28420,N_29101);
nand U31054 (N_31054,N_29644,N_28168);
nand U31055 (N_31055,N_29917,N_29341);
and U31056 (N_31056,N_29327,N_29509);
nor U31057 (N_31057,N_28698,N_29247);
and U31058 (N_31058,N_29657,N_28858);
nor U31059 (N_31059,N_28198,N_28886);
or U31060 (N_31060,N_29891,N_29212);
or U31061 (N_31061,N_28611,N_28327);
nand U31062 (N_31062,N_29872,N_28492);
nor U31063 (N_31063,N_28698,N_28813);
or U31064 (N_31064,N_28992,N_29237);
and U31065 (N_31065,N_28075,N_29644);
and U31066 (N_31066,N_28695,N_28307);
xnor U31067 (N_31067,N_28681,N_29131);
and U31068 (N_31068,N_28218,N_29837);
or U31069 (N_31069,N_28241,N_28541);
xnor U31070 (N_31070,N_28682,N_28790);
or U31071 (N_31071,N_29111,N_29221);
nor U31072 (N_31072,N_29584,N_28371);
xor U31073 (N_31073,N_29839,N_28979);
and U31074 (N_31074,N_29870,N_29597);
or U31075 (N_31075,N_29356,N_28283);
nor U31076 (N_31076,N_29388,N_28990);
and U31077 (N_31077,N_29538,N_28294);
or U31078 (N_31078,N_29565,N_29046);
or U31079 (N_31079,N_28509,N_28371);
and U31080 (N_31080,N_28463,N_28293);
xor U31081 (N_31081,N_29885,N_29447);
nand U31082 (N_31082,N_29940,N_29677);
and U31083 (N_31083,N_29335,N_28777);
and U31084 (N_31084,N_29435,N_28661);
nor U31085 (N_31085,N_28478,N_28392);
xnor U31086 (N_31086,N_28127,N_28338);
or U31087 (N_31087,N_29691,N_28782);
nor U31088 (N_31088,N_28269,N_28149);
nand U31089 (N_31089,N_29998,N_28113);
nand U31090 (N_31090,N_28724,N_28174);
nor U31091 (N_31091,N_28517,N_29183);
nor U31092 (N_31092,N_28671,N_28710);
nor U31093 (N_31093,N_29212,N_29201);
nand U31094 (N_31094,N_29759,N_29430);
xor U31095 (N_31095,N_29455,N_28799);
nor U31096 (N_31096,N_29293,N_29924);
nor U31097 (N_31097,N_29903,N_28023);
nor U31098 (N_31098,N_29277,N_28274);
nand U31099 (N_31099,N_28813,N_29567);
and U31100 (N_31100,N_28730,N_29260);
and U31101 (N_31101,N_29443,N_29616);
xnor U31102 (N_31102,N_28959,N_28257);
and U31103 (N_31103,N_28474,N_28864);
xnor U31104 (N_31104,N_28797,N_28612);
xor U31105 (N_31105,N_28586,N_29650);
or U31106 (N_31106,N_28690,N_29334);
or U31107 (N_31107,N_29840,N_28069);
or U31108 (N_31108,N_29905,N_29142);
xnor U31109 (N_31109,N_29885,N_28011);
nor U31110 (N_31110,N_28644,N_28222);
nor U31111 (N_31111,N_28248,N_29130);
or U31112 (N_31112,N_29204,N_28636);
nor U31113 (N_31113,N_28757,N_28994);
xnor U31114 (N_31114,N_28696,N_29876);
and U31115 (N_31115,N_28399,N_28480);
and U31116 (N_31116,N_29816,N_28237);
xnor U31117 (N_31117,N_28315,N_28610);
nand U31118 (N_31118,N_28472,N_28990);
or U31119 (N_31119,N_28379,N_29490);
nand U31120 (N_31120,N_29476,N_29089);
nand U31121 (N_31121,N_29161,N_28762);
or U31122 (N_31122,N_29448,N_29018);
nand U31123 (N_31123,N_29291,N_29721);
and U31124 (N_31124,N_28614,N_29602);
or U31125 (N_31125,N_29312,N_29836);
nor U31126 (N_31126,N_29543,N_28220);
and U31127 (N_31127,N_29205,N_29235);
nand U31128 (N_31128,N_28782,N_28083);
or U31129 (N_31129,N_29498,N_29361);
or U31130 (N_31130,N_29880,N_28255);
or U31131 (N_31131,N_29173,N_29163);
and U31132 (N_31132,N_29941,N_29463);
nand U31133 (N_31133,N_28280,N_28162);
and U31134 (N_31134,N_29971,N_28993);
nor U31135 (N_31135,N_28179,N_29751);
and U31136 (N_31136,N_28707,N_28305);
or U31137 (N_31137,N_28509,N_28291);
nor U31138 (N_31138,N_28792,N_29136);
nor U31139 (N_31139,N_29206,N_29471);
nor U31140 (N_31140,N_28228,N_29036);
xor U31141 (N_31141,N_29869,N_28428);
or U31142 (N_31142,N_28305,N_29623);
xor U31143 (N_31143,N_28704,N_28365);
nand U31144 (N_31144,N_29118,N_28189);
nor U31145 (N_31145,N_28517,N_28095);
xnor U31146 (N_31146,N_28540,N_29875);
and U31147 (N_31147,N_28014,N_29654);
nor U31148 (N_31148,N_28377,N_29822);
xnor U31149 (N_31149,N_29808,N_28268);
and U31150 (N_31150,N_28349,N_29191);
nand U31151 (N_31151,N_28497,N_29579);
xor U31152 (N_31152,N_29616,N_29981);
or U31153 (N_31153,N_28920,N_29313);
or U31154 (N_31154,N_29036,N_29653);
and U31155 (N_31155,N_29872,N_29963);
nor U31156 (N_31156,N_29157,N_28921);
and U31157 (N_31157,N_29576,N_29912);
nand U31158 (N_31158,N_29923,N_29086);
xor U31159 (N_31159,N_29864,N_29905);
xor U31160 (N_31160,N_29335,N_29340);
and U31161 (N_31161,N_29560,N_29951);
xnor U31162 (N_31162,N_28013,N_29046);
nor U31163 (N_31163,N_29498,N_29778);
xnor U31164 (N_31164,N_29047,N_29086);
nand U31165 (N_31165,N_29172,N_28615);
or U31166 (N_31166,N_29437,N_29096);
or U31167 (N_31167,N_28889,N_29787);
nor U31168 (N_31168,N_28438,N_29258);
nor U31169 (N_31169,N_29086,N_29165);
and U31170 (N_31170,N_29080,N_28745);
and U31171 (N_31171,N_29633,N_29186);
or U31172 (N_31172,N_29969,N_29046);
or U31173 (N_31173,N_29230,N_28317);
xor U31174 (N_31174,N_29110,N_29811);
and U31175 (N_31175,N_28188,N_29407);
or U31176 (N_31176,N_28702,N_29717);
nand U31177 (N_31177,N_28053,N_29018);
nand U31178 (N_31178,N_29277,N_28284);
and U31179 (N_31179,N_28361,N_28054);
or U31180 (N_31180,N_28681,N_29314);
and U31181 (N_31181,N_29194,N_29468);
nand U31182 (N_31182,N_28216,N_28800);
or U31183 (N_31183,N_28404,N_28444);
nor U31184 (N_31184,N_28250,N_28929);
and U31185 (N_31185,N_28482,N_29702);
nand U31186 (N_31186,N_28021,N_29871);
xnor U31187 (N_31187,N_28190,N_28976);
nand U31188 (N_31188,N_28582,N_29069);
nand U31189 (N_31189,N_29535,N_29057);
and U31190 (N_31190,N_28390,N_29757);
nand U31191 (N_31191,N_29496,N_29973);
or U31192 (N_31192,N_28911,N_28788);
and U31193 (N_31193,N_29973,N_28561);
or U31194 (N_31194,N_28680,N_28480);
nor U31195 (N_31195,N_29959,N_28872);
nand U31196 (N_31196,N_28186,N_28256);
or U31197 (N_31197,N_29923,N_28122);
xor U31198 (N_31198,N_29845,N_29430);
nand U31199 (N_31199,N_29468,N_28669);
nand U31200 (N_31200,N_28768,N_29356);
or U31201 (N_31201,N_29808,N_29192);
or U31202 (N_31202,N_28161,N_28401);
nand U31203 (N_31203,N_28206,N_29471);
nor U31204 (N_31204,N_29770,N_29564);
or U31205 (N_31205,N_29539,N_28730);
nand U31206 (N_31206,N_29134,N_28504);
nor U31207 (N_31207,N_28029,N_29307);
xor U31208 (N_31208,N_29671,N_29000);
xnor U31209 (N_31209,N_29270,N_28921);
and U31210 (N_31210,N_29238,N_28112);
xor U31211 (N_31211,N_28970,N_29027);
nand U31212 (N_31212,N_28992,N_28729);
and U31213 (N_31213,N_29729,N_29931);
and U31214 (N_31214,N_28969,N_29750);
and U31215 (N_31215,N_29396,N_28182);
nor U31216 (N_31216,N_28255,N_28287);
xnor U31217 (N_31217,N_28783,N_28789);
nand U31218 (N_31218,N_28219,N_29813);
nor U31219 (N_31219,N_28392,N_29613);
or U31220 (N_31220,N_29898,N_29159);
nor U31221 (N_31221,N_28800,N_28679);
xnor U31222 (N_31222,N_29888,N_28777);
nand U31223 (N_31223,N_29560,N_28904);
and U31224 (N_31224,N_28200,N_29539);
or U31225 (N_31225,N_29185,N_29506);
and U31226 (N_31226,N_29703,N_29746);
nor U31227 (N_31227,N_28272,N_29065);
nor U31228 (N_31228,N_29969,N_29359);
nor U31229 (N_31229,N_29384,N_28004);
xnor U31230 (N_31230,N_29033,N_28367);
nand U31231 (N_31231,N_29578,N_29598);
nor U31232 (N_31232,N_28831,N_28703);
nor U31233 (N_31233,N_29504,N_29760);
nor U31234 (N_31234,N_28820,N_29738);
or U31235 (N_31235,N_28639,N_28655);
nand U31236 (N_31236,N_28941,N_29941);
and U31237 (N_31237,N_29891,N_29133);
and U31238 (N_31238,N_29181,N_28456);
and U31239 (N_31239,N_28247,N_28726);
and U31240 (N_31240,N_29631,N_28336);
xnor U31241 (N_31241,N_29247,N_28461);
xor U31242 (N_31242,N_29010,N_29821);
nor U31243 (N_31243,N_28526,N_28224);
and U31244 (N_31244,N_28734,N_28938);
nor U31245 (N_31245,N_29453,N_28841);
and U31246 (N_31246,N_28594,N_28430);
or U31247 (N_31247,N_28253,N_28266);
and U31248 (N_31248,N_29047,N_29200);
or U31249 (N_31249,N_28026,N_28545);
and U31250 (N_31250,N_29363,N_29047);
xnor U31251 (N_31251,N_28788,N_28342);
or U31252 (N_31252,N_29261,N_28607);
and U31253 (N_31253,N_28994,N_28922);
xnor U31254 (N_31254,N_29242,N_29581);
xor U31255 (N_31255,N_29468,N_28976);
nand U31256 (N_31256,N_29027,N_28911);
nor U31257 (N_31257,N_28714,N_28753);
nand U31258 (N_31258,N_29504,N_29830);
and U31259 (N_31259,N_29347,N_28153);
xnor U31260 (N_31260,N_28306,N_28734);
nand U31261 (N_31261,N_28408,N_28434);
or U31262 (N_31262,N_29407,N_29654);
and U31263 (N_31263,N_28200,N_29883);
or U31264 (N_31264,N_29426,N_29903);
or U31265 (N_31265,N_29445,N_29326);
or U31266 (N_31266,N_28474,N_29194);
xnor U31267 (N_31267,N_29324,N_29344);
xor U31268 (N_31268,N_29438,N_29968);
and U31269 (N_31269,N_29925,N_28947);
nor U31270 (N_31270,N_28519,N_29014);
nor U31271 (N_31271,N_28156,N_29643);
or U31272 (N_31272,N_29467,N_28910);
xor U31273 (N_31273,N_28831,N_29494);
and U31274 (N_31274,N_28357,N_29431);
xnor U31275 (N_31275,N_28897,N_28582);
xor U31276 (N_31276,N_28842,N_29085);
or U31277 (N_31277,N_28527,N_28623);
nand U31278 (N_31278,N_28862,N_28728);
xor U31279 (N_31279,N_28830,N_29292);
and U31280 (N_31280,N_29910,N_29522);
nor U31281 (N_31281,N_28083,N_29878);
and U31282 (N_31282,N_28382,N_29640);
nor U31283 (N_31283,N_29382,N_29477);
and U31284 (N_31284,N_28113,N_28970);
or U31285 (N_31285,N_29048,N_28404);
nor U31286 (N_31286,N_28025,N_28826);
or U31287 (N_31287,N_28263,N_28033);
and U31288 (N_31288,N_29368,N_28138);
nand U31289 (N_31289,N_28860,N_29002);
or U31290 (N_31290,N_28021,N_28252);
nand U31291 (N_31291,N_28419,N_29174);
nor U31292 (N_31292,N_28787,N_29162);
nor U31293 (N_31293,N_29116,N_28184);
or U31294 (N_31294,N_28236,N_28850);
nand U31295 (N_31295,N_28402,N_29837);
and U31296 (N_31296,N_29987,N_29299);
nor U31297 (N_31297,N_28884,N_28150);
xnor U31298 (N_31298,N_29584,N_28422);
xnor U31299 (N_31299,N_29811,N_28666);
and U31300 (N_31300,N_29259,N_29859);
nor U31301 (N_31301,N_28361,N_29640);
nand U31302 (N_31302,N_28484,N_28068);
nor U31303 (N_31303,N_28164,N_28396);
or U31304 (N_31304,N_28126,N_29594);
and U31305 (N_31305,N_29955,N_29495);
nor U31306 (N_31306,N_29660,N_29830);
or U31307 (N_31307,N_28035,N_29655);
nand U31308 (N_31308,N_28088,N_29314);
and U31309 (N_31309,N_28252,N_29643);
and U31310 (N_31310,N_28103,N_29128);
nand U31311 (N_31311,N_29408,N_29584);
nand U31312 (N_31312,N_28413,N_29897);
and U31313 (N_31313,N_28726,N_28539);
and U31314 (N_31314,N_29926,N_29091);
nor U31315 (N_31315,N_28667,N_28462);
nor U31316 (N_31316,N_29076,N_29222);
or U31317 (N_31317,N_28993,N_28851);
nand U31318 (N_31318,N_28614,N_28417);
xnor U31319 (N_31319,N_28763,N_29559);
nor U31320 (N_31320,N_29452,N_28578);
nor U31321 (N_31321,N_28688,N_28548);
xor U31322 (N_31322,N_29142,N_29821);
nor U31323 (N_31323,N_29271,N_29494);
nand U31324 (N_31324,N_28495,N_28396);
and U31325 (N_31325,N_28861,N_28973);
xnor U31326 (N_31326,N_28127,N_29766);
nor U31327 (N_31327,N_28864,N_28799);
or U31328 (N_31328,N_28627,N_28611);
nand U31329 (N_31329,N_29631,N_28046);
nand U31330 (N_31330,N_28687,N_28814);
or U31331 (N_31331,N_28815,N_29140);
xor U31332 (N_31332,N_29183,N_29196);
or U31333 (N_31333,N_29712,N_28275);
nor U31334 (N_31334,N_28898,N_28553);
and U31335 (N_31335,N_29419,N_28444);
or U31336 (N_31336,N_28982,N_29599);
xnor U31337 (N_31337,N_28316,N_29616);
or U31338 (N_31338,N_28460,N_29914);
and U31339 (N_31339,N_29008,N_29288);
nor U31340 (N_31340,N_28745,N_28139);
nor U31341 (N_31341,N_29047,N_28377);
nor U31342 (N_31342,N_28387,N_28491);
nand U31343 (N_31343,N_29113,N_28043);
nor U31344 (N_31344,N_28687,N_29529);
xnor U31345 (N_31345,N_28024,N_28174);
nor U31346 (N_31346,N_29985,N_29185);
or U31347 (N_31347,N_29684,N_29461);
xnor U31348 (N_31348,N_28061,N_29157);
xnor U31349 (N_31349,N_28288,N_28895);
nand U31350 (N_31350,N_29026,N_28933);
or U31351 (N_31351,N_29190,N_28760);
nand U31352 (N_31352,N_28326,N_29737);
xor U31353 (N_31353,N_28460,N_28735);
or U31354 (N_31354,N_29046,N_28332);
nor U31355 (N_31355,N_29003,N_29472);
and U31356 (N_31356,N_29515,N_28854);
nor U31357 (N_31357,N_28191,N_29953);
xnor U31358 (N_31358,N_29773,N_28165);
nand U31359 (N_31359,N_28638,N_28294);
xor U31360 (N_31360,N_29039,N_29273);
and U31361 (N_31361,N_29781,N_28636);
and U31362 (N_31362,N_29851,N_28380);
nand U31363 (N_31363,N_28787,N_29321);
and U31364 (N_31364,N_29395,N_29933);
and U31365 (N_31365,N_29705,N_28424);
and U31366 (N_31366,N_28077,N_28199);
xnor U31367 (N_31367,N_28349,N_29555);
nor U31368 (N_31368,N_29813,N_29404);
or U31369 (N_31369,N_29031,N_29282);
nand U31370 (N_31370,N_29512,N_28455);
nor U31371 (N_31371,N_29091,N_28207);
xor U31372 (N_31372,N_28777,N_29254);
nand U31373 (N_31373,N_29796,N_29638);
and U31374 (N_31374,N_29519,N_28874);
and U31375 (N_31375,N_29124,N_28871);
or U31376 (N_31376,N_28191,N_29754);
nor U31377 (N_31377,N_28370,N_28515);
and U31378 (N_31378,N_28375,N_28323);
and U31379 (N_31379,N_29361,N_28998);
and U31380 (N_31380,N_28230,N_28284);
and U31381 (N_31381,N_28249,N_28831);
and U31382 (N_31382,N_29526,N_28286);
or U31383 (N_31383,N_29607,N_29005);
or U31384 (N_31384,N_28694,N_28015);
xor U31385 (N_31385,N_28748,N_29845);
nor U31386 (N_31386,N_28346,N_28905);
and U31387 (N_31387,N_28688,N_29294);
and U31388 (N_31388,N_29011,N_29394);
xnor U31389 (N_31389,N_28351,N_29088);
or U31390 (N_31390,N_29115,N_29786);
or U31391 (N_31391,N_28531,N_29438);
nor U31392 (N_31392,N_28016,N_29756);
and U31393 (N_31393,N_28132,N_28991);
nand U31394 (N_31394,N_29227,N_28385);
nor U31395 (N_31395,N_29985,N_29775);
nor U31396 (N_31396,N_28753,N_29973);
nor U31397 (N_31397,N_28796,N_28384);
nand U31398 (N_31398,N_28381,N_29432);
nor U31399 (N_31399,N_28723,N_29449);
nor U31400 (N_31400,N_28188,N_28763);
or U31401 (N_31401,N_29808,N_29159);
or U31402 (N_31402,N_29263,N_29785);
and U31403 (N_31403,N_29721,N_28419);
nand U31404 (N_31404,N_29272,N_28986);
and U31405 (N_31405,N_29230,N_28959);
nand U31406 (N_31406,N_28835,N_29296);
nand U31407 (N_31407,N_28742,N_29489);
nor U31408 (N_31408,N_29906,N_28617);
and U31409 (N_31409,N_29708,N_28345);
nor U31410 (N_31410,N_28081,N_28609);
nand U31411 (N_31411,N_28547,N_29066);
nand U31412 (N_31412,N_28819,N_28508);
or U31413 (N_31413,N_29646,N_28336);
xor U31414 (N_31414,N_29397,N_28497);
or U31415 (N_31415,N_28176,N_28528);
xor U31416 (N_31416,N_29721,N_29428);
nor U31417 (N_31417,N_29172,N_28511);
nand U31418 (N_31418,N_28802,N_29164);
and U31419 (N_31419,N_29814,N_29901);
or U31420 (N_31420,N_29616,N_29437);
nor U31421 (N_31421,N_28646,N_29948);
nand U31422 (N_31422,N_28229,N_28400);
and U31423 (N_31423,N_29235,N_28113);
and U31424 (N_31424,N_29606,N_28339);
nand U31425 (N_31425,N_29280,N_28281);
nor U31426 (N_31426,N_28895,N_28180);
nand U31427 (N_31427,N_28297,N_28819);
and U31428 (N_31428,N_29863,N_28641);
and U31429 (N_31429,N_28619,N_28741);
or U31430 (N_31430,N_28477,N_28699);
nand U31431 (N_31431,N_29975,N_29087);
nor U31432 (N_31432,N_28751,N_29334);
nand U31433 (N_31433,N_29337,N_28885);
nor U31434 (N_31434,N_28551,N_29474);
and U31435 (N_31435,N_29539,N_28335);
nand U31436 (N_31436,N_29629,N_29689);
xnor U31437 (N_31437,N_28388,N_29253);
and U31438 (N_31438,N_28849,N_28482);
or U31439 (N_31439,N_29581,N_29964);
nand U31440 (N_31440,N_29252,N_29808);
or U31441 (N_31441,N_29422,N_28402);
and U31442 (N_31442,N_28988,N_29839);
xor U31443 (N_31443,N_29085,N_29952);
and U31444 (N_31444,N_29399,N_29563);
or U31445 (N_31445,N_29003,N_29709);
nor U31446 (N_31446,N_28680,N_28155);
nand U31447 (N_31447,N_28460,N_29032);
and U31448 (N_31448,N_28626,N_28180);
nor U31449 (N_31449,N_29591,N_29257);
or U31450 (N_31450,N_29224,N_29743);
xor U31451 (N_31451,N_29420,N_29625);
or U31452 (N_31452,N_29625,N_28236);
or U31453 (N_31453,N_29376,N_28694);
and U31454 (N_31454,N_29150,N_29840);
or U31455 (N_31455,N_29376,N_29399);
xor U31456 (N_31456,N_29879,N_28928);
and U31457 (N_31457,N_28412,N_29494);
nor U31458 (N_31458,N_28381,N_28752);
nand U31459 (N_31459,N_29729,N_28871);
xor U31460 (N_31460,N_29336,N_28642);
xor U31461 (N_31461,N_28171,N_29055);
and U31462 (N_31462,N_28639,N_29157);
nand U31463 (N_31463,N_29807,N_29434);
nand U31464 (N_31464,N_28815,N_28463);
nor U31465 (N_31465,N_29787,N_28542);
xnor U31466 (N_31466,N_29330,N_29887);
nand U31467 (N_31467,N_29454,N_28969);
nor U31468 (N_31468,N_28458,N_28812);
xnor U31469 (N_31469,N_28237,N_28472);
nand U31470 (N_31470,N_29388,N_28363);
xnor U31471 (N_31471,N_28810,N_28910);
and U31472 (N_31472,N_29971,N_29396);
nor U31473 (N_31473,N_28940,N_28459);
xor U31474 (N_31474,N_29921,N_28461);
nor U31475 (N_31475,N_28391,N_29173);
and U31476 (N_31476,N_28754,N_28755);
xor U31477 (N_31477,N_29362,N_29932);
and U31478 (N_31478,N_28429,N_28655);
or U31479 (N_31479,N_28830,N_29984);
nand U31480 (N_31480,N_28058,N_28293);
nand U31481 (N_31481,N_29344,N_28591);
xor U31482 (N_31482,N_28797,N_29498);
or U31483 (N_31483,N_28547,N_28265);
nand U31484 (N_31484,N_28719,N_29296);
nand U31485 (N_31485,N_28384,N_29883);
xnor U31486 (N_31486,N_29151,N_28914);
xor U31487 (N_31487,N_29359,N_29159);
or U31488 (N_31488,N_28762,N_29898);
or U31489 (N_31489,N_29229,N_29694);
and U31490 (N_31490,N_28246,N_29249);
nor U31491 (N_31491,N_28743,N_29474);
xor U31492 (N_31492,N_28854,N_28534);
xnor U31493 (N_31493,N_29131,N_28326);
nor U31494 (N_31494,N_28609,N_29656);
nor U31495 (N_31495,N_29190,N_29063);
xor U31496 (N_31496,N_29643,N_29003);
or U31497 (N_31497,N_28065,N_28513);
nor U31498 (N_31498,N_29945,N_28647);
nor U31499 (N_31499,N_28164,N_28540);
and U31500 (N_31500,N_28276,N_29043);
nor U31501 (N_31501,N_29107,N_28085);
nor U31502 (N_31502,N_29788,N_28041);
nor U31503 (N_31503,N_28654,N_28397);
xnor U31504 (N_31504,N_29839,N_28566);
or U31505 (N_31505,N_29688,N_28850);
xor U31506 (N_31506,N_29974,N_29020);
nand U31507 (N_31507,N_28913,N_28059);
nor U31508 (N_31508,N_28315,N_28174);
or U31509 (N_31509,N_29204,N_28436);
nand U31510 (N_31510,N_29324,N_28273);
and U31511 (N_31511,N_29445,N_29897);
and U31512 (N_31512,N_29360,N_28883);
or U31513 (N_31513,N_28940,N_29393);
or U31514 (N_31514,N_28756,N_28763);
or U31515 (N_31515,N_29150,N_28660);
and U31516 (N_31516,N_29959,N_28533);
xor U31517 (N_31517,N_28397,N_28730);
nor U31518 (N_31518,N_29700,N_28710);
or U31519 (N_31519,N_29574,N_28106);
or U31520 (N_31520,N_29947,N_29007);
nor U31521 (N_31521,N_28131,N_29137);
and U31522 (N_31522,N_28717,N_29267);
nand U31523 (N_31523,N_28762,N_29757);
nor U31524 (N_31524,N_28014,N_28612);
xor U31525 (N_31525,N_29504,N_28163);
and U31526 (N_31526,N_28997,N_28504);
nor U31527 (N_31527,N_28148,N_28011);
nand U31528 (N_31528,N_28357,N_29300);
nor U31529 (N_31529,N_29256,N_28123);
and U31530 (N_31530,N_28593,N_28867);
xnor U31531 (N_31531,N_28508,N_28602);
or U31532 (N_31532,N_29780,N_28532);
xor U31533 (N_31533,N_29080,N_28280);
xnor U31534 (N_31534,N_29493,N_29858);
nand U31535 (N_31535,N_28576,N_29626);
nand U31536 (N_31536,N_28602,N_29134);
and U31537 (N_31537,N_29181,N_28830);
nor U31538 (N_31538,N_29662,N_28203);
nand U31539 (N_31539,N_29996,N_28622);
or U31540 (N_31540,N_28785,N_29147);
or U31541 (N_31541,N_28056,N_29093);
or U31542 (N_31542,N_28456,N_29815);
nor U31543 (N_31543,N_28156,N_29759);
or U31544 (N_31544,N_28760,N_28471);
nand U31545 (N_31545,N_28632,N_28908);
or U31546 (N_31546,N_29274,N_28538);
or U31547 (N_31547,N_29269,N_28325);
xnor U31548 (N_31548,N_29170,N_28327);
nand U31549 (N_31549,N_28233,N_29065);
nor U31550 (N_31550,N_29522,N_29169);
nor U31551 (N_31551,N_28286,N_28490);
nand U31552 (N_31552,N_28730,N_28162);
xor U31553 (N_31553,N_29862,N_29533);
and U31554 (N_31554,N_28402,N_29060);
nor U31555 (N_31555,N_28427,N_28253);
xor U31556 (N_31556,N_29710,N_28651);
or U31557 (N_31557,N_28114,N_29203);
nand U31558 (N_31558,N_28072,N_28870);
nand U31559 (N_31559,N_29147,N_29392);
xor U31560 (N_31560,N_28091,N_29848);
or U31561 (N_31561,N_28266,N_28426);
xnor U31562 (N_31562,N_29075,N_29227);
nand U31563 (N_31563,N_29516,N_29177);
xnor U31564 (N_31564,N_28485,N_28597);
nand U31565 (N_31565,N_29928,N_29303);
xor U31566 (N_31566,N_28215,N_29784);
or U31567 (N_31567,N_28937,N_29965);
and U31568 (N_31568,N_29235,N_29010);
xnor U31569 (N_31569,N_29005,N_28297);
nor U31570 (N_31570,N_28141,N_28643);
and U31571 (N_31571,N_28573,N_29203);
nor U31572 (N_31572,N_29481,N_29233);
nand U31573 (N_31573,N_28440,N_28253);
nand U31574 (N_31574,N_28382,N_29948);
xor U31575 (N_31575,N_28398,N_29143);
nand U31576 (N_31576,N_28727,N_29388);
xnor U31577 (N_31577,N_29050,N_28077);
nand U31578 (N_31578,N_29035,N_29607);
and U31579 (N_31579,N_29272,N_28130);
or U31580 (N_31580,N_29921,N_28826);
or U31581 (N_31581,N_29800,N_28098);
nand U31582 (N_31582,N_29841,N_28417);
and U31583 (N_31583,N_29795,N_29086);
xor U31584 (N_31584,N_28303,N_29844);
nand U31585 (N_31585,N_29045,N_29753);
nand U31586 (N_31586,N_28386,N_28807);
and U31587 (N_31587,N_28240,N_28200);
and U31588 (N_31588,N_29643,N_28790);
nand U31589 (N_31589,N_29101,N_29366);
and U31590 (N_31590,N_28363,N_28931);
nor U31591 (N_31591,N_28120,N_28771);
xor U31592 (N_31592,N_29930,N_28132);
nand U31593 (N_31593,N_29658,N_28637);
nand U31594 (N_31594,N_28372,N_29391);
or U31595 (N_31595,N_29773,N_28740);
and U31596 (N_31596,N_28295,N_29627);
nand U31597 (N_31597,N_28030,N_28235);
or U31598 (N_31598,N_29904,N_29889);
nand U31599 (N_31599,N_28705,N_28621);
or U31600 (N_31600,N_29795,N_29709);
nor U31601 (N_31601,N_29321,N_29286);
and U31602 (N_31602,N_28220,N_28135);
and U31603 (N_31603,N_28535,N_29261);
nand U31604 (N_31604,N_29539,N_28099);
or U31605 (N_31605,N_28352,N_29262);
and U31606 (N_31606,N_28591,N_28327);
and U31607 (N_31607,N_28548,N_29941);
xnor U31608 (N_31608,N_28360,N_28049);
xor U31609 (N_31609,N_29689,N_28309);
xor U31610 (N_31610,N_29895,N_29912);
or U31611 (N_31611,N_29612,N_29401);
nand U31612 (N_31612,N_29743,N_29657);
nand U31613 (N_31613,N_28147,N_29022);
nand U31614 (N_31614,N_28088,N_28635);
nand U31615 (N_31615,N_29208,N_28354);
xor U31616 (N_31616,N_29749,N_29342);
or U31617 (N_31617,N_29585,N_28861);
xor U31618 (N_31618,N_29798,N_29988);
nand U31619 (N_31619,N_28892,N_28745);
or U31620 (N_31620,N_28883,N_28084);
xnor U31621 (N_31621,N_29763,N_28139);
and U31622 (N_31622,N_29617,N_29118);
xor U31623 (N_31623,N_29942,N_28592);
and U31624 (N_31624,N_28982,N_28244);
or U31625 (N_31625,N_29125,N_28257);
nor U31626 (N_31626,N_29543,N_28958);
and U31627 (N_31627,N_29175,N_28024);
nor U31628 (N_31628,N_28401,N_28725);
or U31629 (N_31629,N_29952,N_29516);
nor U31630 (N_31630,N_28500,N_28217);
xnor U31631 (N_31631,N_28534,N_28527);
or U31632 (N_31632,N_29488,N_29043);
and U31633 (N_31633,N_28541,N_29443);
nand U31634 (N_31634,N_28092,N_28238);
nand U31635 (N_31635,N_28938,N_28209);
nand U31636 (N_31636,N_29782,N_28143);
nor U31637 (N_31637,N_28602,N_29582);
nor U31638 (N_31638,N_28527,N_28428);
or U31639 (N_31639,N_28723,N_29924);
or U31640 (N_31640,N_29531,N_29692);
or U31641 (N_31641,N_28102,N_28631);
xnor U31642 (N_31642,N_29181,N_28603);
nand U31643 (N_31643,N_29970,N_29051);
nor U31644 (N_31644,N_29108,N_28635);
xnor U31645 (N_31645,N_29838,N_29951);
nor U31646 (N_31646,N_29121,N_29979);
nand U31647 (N_31647,N_28286,N_28878);
or U31648 (N_31648,N_28995,N_28161);
xor U31649 (N_31649,N_29830,N_28446);
nand U31650 (N_31650,N_28895,N_28377);
nor U31651 (N_31651,N_29960,N_28634);
nand U31652 (N_31652,N_29291,N_28788);
xnor U31653 (N_31653,N_29800,N_29835);
and U31654 (N_31654,N_29446,N_28194);
nor U31655 (N_31655,N_28358,N_28677);
nand U31656 (N_31656,N_28719,N_29326);
and U31657 (N_31657,N_28795,N_28340);
xor U31658 (N_31658,N_29519,N_29295);
nor U31659 (N_31659,N_28348,N_29089);
nor U31660 (N_31660,N_28896,N_29332);
or U31661 (N_31661,N_29447,N_28181);
nand U31662 (N_31662,N_29945,N_29069);
nor U31663 (N_31663,N_28945,N_28934);
xnor U31664 (N_31664,N_29027,N_28637);
xor U31665 (N_31665,N_28365,N_29895);
or U31666 (N_31666,N_28648,N_28730);
nor U31667 (N_31667,N_28558,N_29470);
nand U31668 (N_31668,N_29172,N_28012);
nand U31669 (N_31669,N_28418,N_28058);
or U31670 (N_31670,N_28867,N_28117);
xor U31671 (N_31671,N_28261,N_28108);
nor U31672 (N_31672,N_29441,N_28022);
nor U31673 (N_31673,N_28974,N_28040);
nor U31674 (N_31674,N_29887,N_29204);
nor U31675 (N_31675,N_29484,N_29244);
and U31676 (N_31676,N_28288,N_29976);
xnor U31677 (N_31677,N_28051,N_28703);
nor U31678 (N_31678,N_28821,N_29487);
nand U31679 (N_31679,N_28009,N_28409);
or U31680 (N_31680,N_29582,N_29440);
nand U31681 (N_31681,N_28819,N_29247);
or U31682 (N_31682,N_28315,N_29405);
nor U31683 (N_31683,N_28480,N_29273);
or U31684 (N_31684,N_29168,N_29300);
and U31685 (N_31685,N_28562,N_29736);
or U31686 (N_31686,N_28284,N_28246);
and U31687 (N_31687,N_28987,N_28917);
nand U31688 (N_31688,N_28685,N_28925);
nand U31689 (N_31689,N_28933,N_28255);
nor U31690 (N_31690,N_28628,N_29144);
or U31691 (N_31691,N_29158,N_28585);
or U31692 (N_31692,N_29447,N_28827);
nor U31693 (N_31693,N_29875,N_28186);
or U31694 (N_31694,N_29942,N_29966);
xor U31695 (N_31695,N_28290,N_28552);
nand U31696 (N_31696,N_29476,N_29817);
and U31697 (N_31697,N_29455,N_28872);
xnor U31698 (N_31698,N_29352,N_28021);
or U31699 (N_31699,N_29882,N_29182);
xnor U31700 (N_31700,N_29254,N_29703);
xnor U31701 (N_31701,N_29981,N_28304);
or U31702 (N_31702,N_28485,N_29496);
xor U31703 (N_31703,N_29684,N_28486);
and U31704 (N_31704,N_29638,N_29027);
and U31705 (N_31705,N_29296,N_28119);
xor U31706 (N_31706,N_28658,N_28177);
or U31707 (N_31707,N_29650,N_29690);
or U31708 (N_31708,N_28347,N_28530);
nand U31709 (N_31709,N_28201,N_28948);
xnor U31710 (N_31710,N_28605,N_29187);
nand U31711 (N_31711,N_29894,N_28918);
nor U31712 (N_31712,N_28830,N_28235);
nand U31713 (N_31713,N_29329,N_29690);
nor U31714 (N_31714,N_29605,N_28110);
and U31715 (N_31715,N_28209,N_29835);
and U31716 (N_31716,N_28222,N_28525);
and U31717 (N_31717,N_29461,N_29750);
xnor U31718 (N_31718,N_28352,N_29074);
or U31719 (N_31719,N_28407,N_29049);
nand U31720 (N_31720,N_28500,N_29390);
nor U31721 (N_31721,N_28570,N_28552);
xnor U31722 (N_31722,N_28787,N_28978);
or U31723 (N_31723,N_28896,N_29563);
and U31724 (N_31724,N_28829,N_28964);
and U31725 (N_31725,N_29713,N_29694);
and U31726 (N_31726,N_28634,N_28842);
nand U31727 (N_31727,N_28004,N_29584);
and U31728 (N_31728,N_29994,N_28632);
and U31729 (N_31729,N_28883,N_28192);
nor U31730 (N_31730,N_29322,N_28333);
xor U31731 (N_31731,N_28336,N_28724);
xnor U31732 (N_31732,N_29314,N_29062);
nand U31733 (N_31733,N_29545,N_28848);
or U31734 (N_31734,N_28336,N_28802);
nand U31735 (N_31735,N_28594,N_28306);
nand U31736 (N_31736,N_29210,N_29275);
nand U31737 (N_31737,N_28651,N_29767);
or U31738 (N_31738,N_28380,N_28946);
xor U31739 (N_31739,N_28142,N_29186);
and U31740 (N_31740,N_29101,N_28523);
nand U31741 (N_31741,N_29335,N_29719);
and U31742 (N_31742,N_29788,N_29308);
xor U31743 (N_31743,N_28688,N_28147);
nor U31744 (N_31744,N_28540,N_28548);
or U31745 (N_31745,N_28991,N_28613);
and U31746 (N_31746,N_29941,N_28315);
xor U31747 (N_31747,N_28744,N_29323);
and U31748 (N_31748,N_29734,N_29531);
and U31749 (N_31749,N_29582,N_28067);
xnor U31750 (N_31750,N_28473,N_29808);
or U31751 (N_31751,N_28366,N_29870);
and U31752 (N_31752,N_29172,N_29456);
nor U31753 (N_31753,N_29236,N_28242);
nor U31754 (N_31754,N_28019,N_29137);
and U31755 (N_31755,N_29726,N_29574);
and U31756 (N_31756,N_28348,N_28201);
or U31757 (N_31757,N_29025,N_29379);
nand U31758 (N_31758,N_28767,N_28896);
xor U31759 (N_31759,N_28435,N_28934);
nand U31760 (N_31760,N_28528,N_29183);
or U31761 (N_31761,N_28036,N_29862);
or U31762 (N_31762,N_28991,N_29054);
nor U31763 (N_31763,N_28447,N_28369);
xnor U31764 (N_31764,N_28217,N_29243);
or U31765 (N_31765,N_29133,N_29710);
nand U31766 (N_31766,N_28294,N_28255);
nand U31767 (N_31767,N_28376,N_28691);
or U31768 (N_31768,N_29191,N_29664);
or U31769 (N_31769,N_29422,N_28913);
and U31770 (N_31770,N_29348,N_28265);
or U31771 (N_31771,N_29699,N_29826);
xnor U31772 (N_31772,N_29436,N_29659);
xnor U31773 (N_31773,N_28998,N_28036);
xor U31774 (N_31774,N_29952,N_28984);
nor U31775 (N_31775,N_28899,N_29831);
or U31776 (N_31776,N_28641,N_29030);
nor U31777 (N_31777,N_29474,N_28356);
and U31778 (N_31778,N_28648,N_28060);
or U31779 (N_31779,N_29858,N_29103);
and U31780 (N_31780,N_28766,N_29633);
nand U31781 (N_31781,N_29868,N_29402);
xnor U31782 (N_31782,N_28609,N_29393);
or U31783 (N_31783,N_28749,N_28946);
nand U31784 (N_31784,N_29311,N_28667);
nand U31785 (N_31785,N_29846,N_29171);
nor U31786 (N_31786,N_29188,N_28498);
or U31787 (N_31787,N_28379,N_28708);
xnor U31788 (N_31788,N_29768,N_28223);
xnor U31789 (N_31789,N_28884,N_29186);
xnor U31790 (N_31790,N_29299,N_28255);
nand U31791 (N_31791,N_29996,N_28952);
nand U31792 (N_31792,N_28670,N_28346);
and U31793 (N_31793,N_29151,N_28461);
or U31794 (N_31794,N_28577,N_29939);
and U31795 (N_31795,N_28600,N_28726);
and U31796 (N_31796,N_28030,N_28213);
or U31797 (N_31797,N_29767,N_28181);
nand U31798 (N_31798,N_28940,N_28332);
nand U31799 (N_31799,N_28916,N_28227);
xor U31800 (N_31800,N_28289,N_29670);
xor U31801 (N_31801,N_28503,N_29788);
or U31802 (N_31802,N_29457,N_29857);
xnor U31803 (N_31803,N_28402,N_29851);
xnor U31804 (N_31804,N_28006,N_28683);
nor U31805 (N_31805,N_29902,N_28903);
xor U31806 (N_31806,N_29340,N_29723);
nor U31807 (N_31807,N_28193,N_29267);
and U31808 (N_31808,N_29373,N_28610);
nand U31809 (N_31809,N_28425,N_28075);
or U31810 (N_31810,N_29249,N_28452);
or U31811 (N_31811,N_29923,N_29892);
nor U31812 (N_31812,N_29501,N_28027);
nor U31813 (N_31813,N_29431,N_28832);
or U31814 (N_31814,N_29937,N_28044);
nor U31815 (N_31815,N_29219,N_28858);
and U31816 (N_31816,N_29337,N_28480);
nand U31817 (N_31817,N_28194,N_29167);
nand U31818 (N_31818,N_29460,N_29414);
nor U31819 (N_31819,N_28868,N_28423);
nand U31820 (N_31820,N_29755,N_28837);
and U31821 (N_31821,N_29893,N_29501);
xnor U31822 (N_31822,N_28802,N_29600);
xor U31823 (N_31823,N_28271,N_28299);
xor U31824 (N_31824,N_29498,N_28477);
xor U31825 (N_31825,N_29346,N_28740);
xor U31826 (N_31826,N_28763,N_29681);
or U31827 (N_31827,N_29129,N_28732);
nand U31828 (N_31828,N_28112,N_29587);
nor U31829 (N_31829,N_29105,N_29783);
xor U31830 (N_31830,N_29602,N_29275);
nor U31831 (N_31831,N_28340,N_29301);
xnor U31832 (N_31832,N_29827,N_29834);
and U31833 (N_31833,N_28061,N_29431);
nor U31834 (N_31834,N_29453,N_28207);
nor U31835 (N_31835,N_29576,N_29771);
xor U31836 (N_31836,N_29754,N_28520);
nand U31837 (N_31837,N_29826,N_29602);
and U31838 (N_31838,N_29260,N_29357);
nor U31839 (N_31839,N_28452,N_28086);
xnor U31840 (N_31840,N_28802,N_28229);
xnor U31841 (N_31841,N_28904,N_28310);
and U31842 (N_31842,N_29075,N_28546);
nor U31843 (N_31843,N_28004,N_28569);
or U31844 (N_31844,N_28408,N_29550);
or U31845 (N_31845,N_29300,N_29220);
xnor U31846 (N_31846,N_29873,N_29785);
and U31847 (N_31847,N_28964,N_29239);
and U31848 (N_31848,N_29030,N_29075);
xnor U31849 (N_31849,N_29791,N_29360);
nand U31850 (N_31850,N_29874,N_28149);
xnor U31851 (N_31851,N_29425,N_28749);
nand U31852 (N_31852,N_28371,N_28139);
or U31853 (N_31853,N_28622,N_29625);
nand U31854 (N_31854,N_28496,N_28450);
and U31855 (N_31855,N_28778,N_28086);
nand U31856 (N_31856,N_29343,N_28231);
nand U31857 (N_31857,N_28829,N_28021);
nand U31858 (N_31858,N_29704,N_29168);
nor U31859 (N_31859,N_28800,N_28920);
nand U31860 (N_31860,N_28206,N_29235);
or U31861 (N_31861,N_29865,N_28480);
and U31862 (N_31862,N_29442,N_29736);
nand U31863 (N_31863,N_29836,N_29856);
and U31864 (N_31864,N_29965,N_28199);
nor U31865 (N_31865,N_28033,N_28253);
and U31866 (N_31866,N_29307,N_29524);
nand U31867 (N_31867,N_28273,N_29445);
xnor U31868 (N_31868,N_28580,N_29875);
and U31869 (N_31869,N_28296,N_29803);
nor U31870 (N_31870,N_28504,N_29560);
nor U31871 (N_31871,N_28299,N_28072);
nand U31872 (N_31872,N_28289,N_29003);
nor U31873 (N_31873,N_29121,N_29097);
or U31874 (N_31874,N_29817,N_28537);
nor U31875 (N_31875,N_29313,N_28774);
xnor U31876 (N_31876,N_29118,N_29066);
nand U31877 (N_31877,N_29472,N_28331);
xor U31878 (N_31878,N_28505,N_29589);
nand U31879 (N_31879,N_28706,N_29692);
nor U31880 (N_31880,N_28718,N_28684);
xnor U31881 (N_31881,N_28755,N_28464);
and U31882 (N_31882,N_29791,N_29183);
or U31883 (N_31883,N_28820,N_28260);
or U31884 (N_31884,N_28297,N_29260);
nand U31885 (N_31885,N_28601,N_28809);
xnor U31886 (N_31886,N_28124,N_28504);
nand U31887 (N_31887,N_28018,N_29627);
nand U31888 (N_31888,N_28981,N_28098);
xor U31889 (N_31889,N_28522,N_28651);
or U31890 (N_31890,N_29895,N_29661);
and U31891 (N_31891,N_29896,N_29242);
or U31892 (N_31892,N_28845,N_28873);
nor U31893 (N_31893,N_28242,N_29803);
xor U31894 (N_31894,N_29137,N_28205);
xor U31895 (N_31895,N_28412,N_29242);
and U31896 (N_31896,N_29010,N_28204);
nand U31897 (N_31897,N_28601,N_29709);
nand U31898 (N_31898,N_29553,N_29353);
or U31899 (N_31899,N_28112,N_29514);
nand U31900 (N_31900,N_28269,N_28610);
nand U31901 (N_31901,N_29853,N_28833);
xnor U31902 (N_31902,N_28941,N_28622);
or U31903 (N_31903,N_29071,N_28714);
nor U31904 (N_31904,N_28685,N_29415);
and U31905 (N_31905,N_28885,N_29775);
nand U31906 (N_31906,N_29231,N_29274);
nand U31907 (N_31907,N_28218,N_28319);
and U31908 (N_31908,N_28298,N_29528);
and U31909 (N_31909,N_29005,N_29575);
or U31910 (N_31910,N_28192,N_29969);
or U31911 (N_31911,N_28827,N_28380);
and U31912 (N_31912,N_29408,N_29698);
or U31913 (N_31913,N_28063,N_29961);
and U31914 (N_31914,N_29768,N_28704);
nor U31915 (N_31915,N_28629,N_29253);
nand U31916 (N_31916,N_28471,N_29250);
nand U31917 (N_31917,N_29234,N_28171);
and U31918 (N_31918,N_29871,N_28024);
nor U31919 (N_31919,N_29216,N_28336);
or U31920 (N_31920,N_28159,N_29644);
nor U31921 (N_31921,N_28944,N_29717);
nor U31922 (N_31922,N_29510,N_29801);
nand U31923 (N_31923,N_28931,N_29337);
nor U31924 (N_31924,N_28036,N_28690);
nand U31925 (N_31925,N_29122,N_28689);
nor U31926 (N_31926,N_29406,N_28382);
xnor U31927 (N_31927,N_28824,N_28368);
xor U31928 (N_31928,N_29879,N_28476);
nor U31929 (N_31929,N_28396,N_28645);
or U31930 (N_31930,N_28697,N_29471);
nor U31931 (N_31931,N_29260,N_29442);
or U31932 (N_31932,N_28335,N_28218);
xnor U31933 (N_31933,N_29482,N_29524);
or U31934 (N_31934,N_29815,N_29667);
nand U31935 (N_31935,N_28177,N_29104);
nor U31936 (N_31936,N_29462,N_29170);
or U31937 (N_31937,N_29390,N_28184);
and U31938 (N_31938,N_29132,N_28434);
xnor U31939 (N_31939,N_29661,N_29247);
and U31940 (N_31940,N_28406,N_29453);
nand U31941 (N_31941,N_28729,N_28484);
nor U31942 (N_31942,N_29593,N_29139);
nor U31943 (N_31943,N_29925,N_29473);
nor U31944 (N_31944,N_28739,N_28291);
nand U31945 (N_31945,N_29845,N_29729);
and U31946 (N_31946,N_28566,N_29815);
xnor U31947 (N_31947,N_29286,N_28679);
and U31948 (N_31948,N_28347,N_29102);
nand U31949 (N_31949,N_29849,N_29164);
xor U31950 (N_31950,N_29762,N_28306);
nor U31951 (N_31951,N_29529,N_28699);
xnor U31952 (N_31952,N_28353,N_28377);
nand U31953 (N_31953,N_29489,N_29045);
nand U31954 (N_31954,N_28796,N_29239);
xnor U31955 (N_31955,N_29527,N_29901);
or U31956 (N_31956,N_29231,N_28996);
or U31957 (N_31957,N_28917,N_29611);
and U31958 (N_31958,N_29085,N_28387);
nor U31959 (N_31959,N_28812,N_29217);
and U31960 (N_31960,N_29685,N_29236);
xor U31961 (N_31961,N_29495,N_28318);
nand U31962 (N_31962,N_28154,N_29663);
and U31963 (N_31963,N_29043,N_29368);
or U31964 (N_31964,N_28575,N_28504);
or U31965 (N_31965,N_28371,N_29045);
nor U31966 (N_31966,N_29107,N_29574);
nor U31967 (N_31967,N_28892,N_29972);
and U31968 (N_31968,N_29854,N_28105);
xnor U31969 (N_31969,N_28148,N_28514);
nand U31970 (N_31970,N_28902,N_28785);
xnor U31971 (N_31971,N_29559,N_28801);
xnor U31972 (N_31972,N_29063,N_29833);
or U31973 (N_31973,N_28441,N_29214);
xor U31974 (N_31974,N_29093,N_29743);
nand U31975 (N_31975,N_29746,N_29730);
nand U31976 (N_31976,N_29313,N_29190);
and U31977 (N_31977,N_28747,N_28445);
or U31978 (N_31978,N_29668,N_28805);
nor U31979 (N_31979,N_29033,N_28871);
nor U31980 (N_31980,N_29696,N_29936);
nand U31981 (N_31981,N_29824,N_28121);
xnor U31982 (N_31982,N_29670,N_29589);
or U31983 (N_31983,N_29062,N_28496);
nor U31984 (N_31984,N_29911,N_29418);
nand U31985 (N_31985,N_29767,N_28351);
nand U31986 (N_31986,N_29886,N_28494);
and U31987 (N_31987,N_28546,N_28498);
nor U31988 (N_31988,N_29652,N_29821);
and U31989 (N_31989,N_29138,N_28797);
xor U31990 (N_31990,N_28567,N_29409);
and U31991 (N_31991,N_29188,N_29637);
nor U31992 (N_31992,N_29146,N_29398);
nor U31993 (N_31993,N_29339,N_28642);
xor U31994 (N_31994,N_28625,N_29876);
xnor U31995 (N_31995,N_28925,N_29874);
nand U31996 (N_31996,N_28396,N_29609);
nor U31997 (N_31997,N_28248,N_28451);
and U31998 (N_31998,N_28965,N_28209);
and U31999 (N_31999,N_28110,N_28122);
nor U32000 (N_32000,N_30978,N_31490);
nor U32001 (N_32001,N_30533,N_31926);
xnor U32002 (N_32002,N_31523,N_30448);
nand U32003 (N_32003,N_31911,N_31456);
and U32004 (N_32004,N_30436,N_31977);
and U32005 (N_32005,N_30074,N_30262);
or U32006 (N_32006,N_30101,N_30960);
nor U32007 (N_32007,N_31001,N_31649);
and U32008 (N_32008,N_30626,N_31793);
nor U32009 (N_32009,N_31244,N_31408);
and U32010 (N_32010,N_30623,N_30048);
xor U32011 (N_32011,N_31288,N_30974);
nand U32012 (N_32012,N_31352,N_31894);
nand U32013 (N_32013,N_30182,N_30096);
and U32014 (N_32014,N_30830,N_31849);
nand U32015 (N_32015,N_31133,N_30965);
xor U32016 (N_32016,N_31810,N_31417);
nand U32017 (N_32017,N_31956,N_31949);
nand U32018 (N_32018,N_30632,N_30019);
xor U32019 (N_32019,N_31897,N_30037);
xor U32020 (N_32020,N_30038,N_31064);
xnor U32021 (N_32021,N_30153,N_31188);
nor U32022 (N_32022,N_31636,N_30762);
nand U32023 (N_32023,N_30730,N_31454);
nand U32024 (N_32024,N_31983,N_31089);
nand U32025 (N_32025,N_30144,N_31913);
or U32026 (N_32026,N_31449,N_30158);
nor U32027 (N_32027,N_31340,N_31403);
or U32028 (N_32028,N_30909,N_31836);
nand U32029 (N_32029,N_31960,N_31997);
nor U32030 (N_32030,N_31317,N_31726);
nor U32031 (N_32031,N_30968,N_31308);
xor U32032 (N_32032,N_30699,N_31973);
nor U32033 (N_32033,N_31604,N_31896);
xnor U32034 (N_32034,N_31728,N_31758);
and U32035 (N_32035,N_31295,N_31821);
nor U32036 (N_32036,N_30201,N_31218);
xor U32037 (N_32037,N_31424,N_31119);
and U32038 (N_32038,N_31080,N_30889);
or U32039 (N_32039,N_31768,N_30484);
nand U32040 (N_32040,N_30069,N_30439);
nand U32041 (N_32041,N_31666,N_31933);
and U32042 (N_32042,N_31816,N_30270);
xor U32043 (N_32043,N_31060,N_30597);
nor U32044 (N_32044,N_31304,N_30024);
nand U32045 (N_32045,N_31615,N_31274);
xnor U32046 (N_32046,N_31923,N_31412);
xnor U32047 (N_32047,N_30177,N_31260);
xor U32048 (N_32048,N_30726,N_30209);
or U32049 (N_32049,N_31632,N_31290);
xor U32050 (N_32050,N_31463,N_30156);
nor U32051 (N_32051,N_31267,N_31455);
or U32052 (N_32052,N_31738,N_30339);
or U32053 (N_32053,N_31177,N_31660);
xnor U32054 (N_32054,N_30149,N_31785);
nand U32055 (N_32055,N_31679,N_30513);
and U32056 (N_32056,N_31322,N_30652);
nor U32057 (N_32057,N_31185,N_30694);
xor U32058 (N_32058,N_31556,N_30303);
nand U32059 (N_32059,N_30160,N_30495);
and U32060 (N_32060,N_30592,N_31062);
and U32061 (N_32061,N_30518,N_30396);
and U32062 (N_32062,N_30725,N_31837);
nand U32063 (N_32063,N_30264,N_30105);
or U32064 (N_32064,N_31381,N_31867);
nor U32065 (N_32065,N_30346,N_31864);
and U32066 (N_32066,N_31413,N_30745);
xor U32067 (N_32067,N_31259,N_31674);
nor U32068 (N_32068,N_30213,N_31780);
or U32069 (N_32069,N_31311,N_31238);
nor U32070 (N_32070,N_30918,N_31655);
nand U32071 (N_32071,N_30471,N_30344);
xnor U32072 (N_32072,N_30366,N_31646);
nand U32073 (N_32073,N_30738,N_30550);
or U32074 (N_32074,N_30227,N_31959);
xnor U32075 (N_32075,N_30296,N_31221);
and U32076 (N_32076,N_30211,N_31234);
or U32077 (N_32077,N_31709,N_31981);
and U32078 (N_32078,N_30145,N_31915);
and U32079 (N_32079,N_30335,N_31103);
nand U32080 (N_32080,N_31982,N_31801);
nand U32081 (N_32081,N_30140,N_30188);
or U32082 (N_32082,N_31624,N_30406);
nand U32083 (N_32083,N_31710,N_31204);
and U32084 (N_32084,N_31426,N_30364);
or U32085 (N_32085,N_30655,N_31727);
nor U32086 (N_32086,N_30580,N_31325);
nor U32087 (N_32087,N_30208,N_31677);
and U32088 (N_32088,N_31979,N_30404);
and U32089 (N_32089,N_30467,N_31819);
xnor U32090 (N_32090,N_30287,N_30685);
nor U32091 (N_32091,N_30068,N_30020);
and U32092 (N_32092,N_31741,N_31106);
nor U32093 (N_32093,N_30435,N_30141);
nand U32094 (N_32094,N_31831,N_30875);
or U32095 (N_32095,N_30542,N_31430);
nor U32096 (N_32096,N_31049,N_30767);
and U32097 (N_32097,N_31158,N_30292);
and U32098 (N_32098,N_30848,N_30373);
nor U32099 (N_32099,N_30446,N_30713);
or U32100 (N_32100,N_31642,N_30319);
nand U32101 (N_32101,N_31714,N_30840);
nand U32102 (N_32102,N_30253,N_30554);
nor U32103 (N_32103,N_30825,N_31282);
nand U32104 (N_32104,N_30108,N_30982);
xnor U32105 (N_32105,N_30089,N_31358);
and U32106 (N_32106,N_30415,N_30214);
nand U32107 (N_32107,N_31687,N_30739);
xor U32108 (N_32108,N_31372,N_30804);
xor U32109 (N_32109,N_30747,N_30817);
nand U32110 (N_32110,N_31688,N_31483);
and U32111 (N_32111,N_31929,N_31800);
xor U32112 (N_32112,N_31077,N_31389);
and U32113 (N_32113,N_31100,N_30838);
or U32114 (N_32114,N_31740,N_30806);
nand U32115 (N_32115,N_30734,N_31895);
or U32116 (N_32116,N_31623,N_31941);
xor U32117 (N_32117,N_30285,N_30330);
and U32118 (N_32118,N_31429,N_31385);
and U32119 (N_32119,N_31198,N_30576);
or U32120 (N_32120,N_31494,N_31190);
nor U32121 (N_32121,N_30980,N_31347);
and U32122 (N_32122,N_31685,N_31083);
xor U32123 (N_32123,N_31892,N_30322);
xor U32124 (N_32124,N_31086,N_31349);
and U32125 (N_32125,N_30640,N_30937);
nor U32126 (N_32126,N_31310,N_30206);
and U32127 (N_32127,N_30923,N_31153);
and U32128 (N_32128,N_30361,N_30511);
and U32129 (N_32129,N_31675,N_30677);
or U32130 (N_32130,N_31191,N_30774);
nor U32131 (N_32131,N_30260,N_30827);
and U32132 (N_32132,N_30055,N_30263);
nand U32133 (N_32133,N_30083,N_31551);
or U32134 (N_32134,N_30220,N_31113);
xnor U32135 (N_32135,N_31067,N_31240);
xor U32136 (N_32136,N_30246,N_31420);
and U32137 (N_32137,N_31447,N_30579);
and U32138 (N_32138,N_31134,N_30133);
nand U32139 (N_32139,N_30901,N_31070);
or U32140 (N_32140,N_30168,N_31374);
xor U32141 (N_32141,N_30539,N_30028);
nand U32142 (N_32142,N_30801,N_30023);
nand U32143 (N_32143,N_31559,N_30199);
or U32144 (N_32144,N_30823,N_30075);
or U32145 (N_32145,N_31453,N_31535);
xor U32146 (N_32146,N_30919,N_30894);
xnor U32147 (N_32147,N_30218,N_31508);
or U32148 (N_32148,N_31414,N_31847);
or U32149 (N_32149,N_31465,N_31283);
and U32150 (N_32150,N_30805,N_31316);
and U32151 (N_32151,N_31052,N_31418);
nand U32152 (N_32152,N_30625,N_31937);
or U32153 (N_32153,N_31013,N_30914);
and U32154 (N_32154,N_31572,N_30050);
and U32155 (N_32155,N_31826,N_31396);
and U32156 (N_32156,N_31015,N_31691);
xor U32157 (N_32157,N_31294,N_30631);
nor U32158 (N_32158,N_30957,N_30298);
nor U32159 (N_32159,N_31686,N_30671);
or U32160 (N_32160,N_30190,N_30131);
xnor U32161 (N_32161,N_30546,N_31910);
and U32162 (N_32162,N_30724,N_31205);
nor U32163 (N_32163,N_30035,N_30305);
nand U32164 (N_32164,N_31628,N_31024);
xor U32165 (N_32165,N_30086,N_31605);
nor U32166 (N_32166,N_31442,N_30485);
xnor U32167 (N_32167,N_30594,N_30920);
nor U32168 (N_32168,N_30947,N_30200);
xor U32169 (N_32169,N_30519,N_31183);
nor U32170 (N_32170,N_30252,N_30810);
xor U32171 (N_32171,N_30112,N_30723);
nor U32172 (N_32172,N_30635,N_31008);
nand U32173 (N_32173,N_31293,N_31504);
nand U32174 (N_32174,N_31730,N_30565);
or U32175 (N_32175,N_31359,N_31634);
or U32176 (N_32176,N_31265,N_31107);
nor U32177 (N_32177,N_31639,N_31795);
nand U32178 (N_32178,N_30386,N_30783);
nor U32179 (N_32179,N_31850,N_30202);
xor U32180 (N_32180,N_31635,N_30824);
nand U32181 (N_32181,N_31068,N_30135);
xnor U32182 (N_32182,N_30499,N_30629);
and U32183 (N_32183,N_30690,N_30512);
xnor U32184 (N_32184,N_30167,N_31613);
nand U32185 (N_32185,N_30721,N_31650);
nand U32186 (N_32186,N_31278,N_31767);
xnor U32187 (N_32187,N_30039,N_31472);
and U32188 (N_32188,N_30047,N_30682);
or U32189 (N_32189,N_30052,N_31287);
xnor U32190 (N_32190,N_31232,N_31373);
xor U32191 (N_32191,N_30977,N_31644);
xor U32192 (N_32192,N_31787,N_31326);
nand U32193 (N_32193,N_30586,N_30938);
and U32194 (N_32194,N_31763,N_31314);
nor U32195 (N_32195,N_31380,N_31841);
or U32196 (N_32196,N_30714,N_30362);
and U32197 (N_32197,N_30867,N_31735);
nand U32198 (N_32198,N_30608,N_31757);
and U32199 (N_32199,N_30456,N_31048);
and U32200 (N_32200,N_31952,N_31434);
nor U32201 (N_32201,N_30462,N_31502);
and U32202 (N_32202,N_31118,N_30116);
or U32203 (N_32203,N_30704,N_31222);
or U32204 (N_32204,N_30399,N_30136);
xor U32205 (N_32205,N_31269,N_31227);
or U32206 (N_32206,N_30084,N_31762);
nor U32207 (N_32207,N_31264,N_31174);
nand U32208 (N_32208,N_31032,N_31362);
or U32209 (N_32209,N_30314,N_31560);
xnor U32210 (N_32210,N_30290,N_31654);
nand U32211 (N_32211,N_30870,N_30618);
xnor U32212 (N_32212,N_31808,N_31945);
xnor U32213 (N_32213,N_30316,N_30814);
nor U32214 (N_32214,N_30186,N_30115);
or U32215 (N_32215,N_30033,N_31891);
nand U32216 (N_32216,N_30321,N_31866);
nor U32217 (N_32217,N_31579,N_31301);
nand U32218 (N_32218,N_30871,N_31046);
and U32219 (N_32219,N_31631,N_30152);
nor U32220 (N_32220,N_31939,N_31718);
xnor U32221 (N_32221,N_31824,N_31725);
nand U32222 (N_32222,N_30216,N_31590);
nor U32223 (N_32223,N_31815,N_31073);
and U32224 (N_32224,N_30660,N_31307);
nand U32225 (N_32225,N_30737,N_31868);
and U32226 (N_32226,N_30657,N_30056);
or U32227 (N_32227,N_30798,N_30663);
xnor U32228 (N_32228,N_31415,N_31263);
and U32229 (N_32229,N_31803,N_31286);
or U32230 (N_32230,N_30256,N_31582);
nand U32231 (N_32231,N_30482,N_31909);
or U32232 (N_32232,N_30654,N_31402);
nand U32233 (N_32233,N_30999,N_30046);
and U32234 (N_32234,N_30861,N_30778);
nor U32235 (N_32235,N_30526,N_31102);
nand U32236 (N_32236,N_31899,N_30772);
and U32237 (N_32237,N_31625,N_30754);
nand U32238 (N_32238,N_30181,N_31395);
and U32239 (N_32239,N_31859,N_31392);
and U32240 (N_32240,N_31746,N_31000);
nor U32241 (N_32241,N_31390,N_31026);
and U32242 (N_32242,N_31769,N_31781);
nand U32243 (N_32243,N_31647,N_31432);
nor U32244 (N_32244,N_30045,N_31441);
or U32245 (N_32245,N_30839,N_31883);
nand U32246 (N_32246,N_30548,N_31886);
and U32247 (N_32247,N_31607,N_31275);
or U32248 (N_32248,N_30588,N_31079);
nand U32249 (N_32249,N_30222,N_30241);
nor U32250 (N_32250,N_30890,N_31266);
or U32251 (N_32251,N_30493,N_30800);
nand U32252 (N_32252,N_31898,N_30882);
and U32253 (N_32253,N_30098,N_30317);
xnor U32254 (N_32254,N_30537,N_31236);
and U32255 (N_32255,N_30329,N_30434);
and U32256 (N_32256,N_30427,N_31843);
xnor U32257 (N_32257,N_31142,N_30172);
or U32258 (N_32258,N_31594,N_30555);
nand U32259 (N_32259,N_31854,N_31323);
and U32260 (N_32260,N_30297,N_31262);
xor U32261 (N_32261,N_31518,N_30433);
nor U32262 (N_32262,N_31969,N_30194);
or U32263 (N_32263,N_31419,N_31863);
or U32264 (N_32264,N_30197,N_31182);
or U32265 (N_32265,N_31680,N_30233);
or U32266 (N_32266,N_31889,N_31703);
or U32267 (N_32267,N_31571,N_30771);
nor U32268 (N_32268,N_30275,N_30575);
nor U32269 (N_32269,N_31245,N_31798);
nand U32270 (N_32270,N_30650,N_31870);
and U32271 (N_32271,N_31497,N_31099);
or U32272 (N_32272,N_31862,N_30443);
nand U32273 (N_32273,N_31509,N_31890);
nand U32274 (N_32274,N_31489,N_31360);
or U32275 (N_32275,N_30232,N_30185);
xnor U32276 (N_32276,N_30180,N_30864);
nor U32277 (N_32277,N_31276,N_31367);
xor U32278 (N_32278,N_30378,N_30568);
xnor U32279 (N_32279,N_31742,N_31382);
nor U32280 (N_32280,N_31452,N_30418);
nor U32281 (N_32281,N_30081,N_30114);
nor U32282 (N_32282,N_30274,N_30766);
and U32283 (N_32283,N_31733,N_30929);
nor U32284 (N_32284,N_30178,N_30480);
xor U32285 (N_32285,N_30627,N_31593);
nand U32286 (N_32286,N_30502,N_30731);
or U32287 (N_32287,N_31467,N_31657);
or U32288 (N_32288,N_30470,N_31566);
and U32289 (N_32289,N_31313,N_31496);
xnor U32290 (N_32290,N_31169,N_30506);
nor U32291 (N_32291,N_30312,N_31194);
and U32292 (N_32292,N_30641,N_31531);
xor U32293 (N_32293,N_31331,N_31123);
or U32294 (N_32294,N_30769,N_30904);
or U32295 (N_32295,N_30230,N_31946);
xnor U32296 (N_32296,N_30390,N_30010);
or U32297 (N_32297,N_31547,N_31124);
or U32298 (N_32298,N_30529,N_31541);
or U32299 (N_32299,N_30916,N_30358);
or U32300 (N_32300,N_30925,N_31516);
or U32301 (N_32301,N_31958,N_31027);
and U32302 (N_32302,N_30455,N_30868);
nor U32303 (N_32303,N_30082,N_30698);
xnor U32304 (N_32304,N_30057,N_30637);
and U32305 (N_32305,N_30796,N_30066);
and U32306 (N_32306,N_31629,N_30647);
or U32307 (N_32307,N_30602,N_30828);
xor U32308 (N_32308,N_31967,N_31054);
and U32309 (N_32309,N_30041,N_30736);
or U32310 (N_32310,N_30788,N_31476);
and U32311 (N_32311,N_31672,N_30858);
nor U32312 (N_32312,N_30006,N_31962);
and U32313 (N_32313,N_31019,N_31552);
nand U32314 (N_32314,N_30989,N_30667);
nand U32315 (N_32315,N_31342,N_31659);
and U32316 (N_32316,N_30459,N_30031);
nor U32317 (N_32317,N_31643,N_30496);
xnor U32318 (N_32318,N_30844,N_30874);
or U32319 (N_32319,N_30077,N_30915);
and U32320 (N_32320,N_30616,N_31700);
nor U32321 (N_32321,N_31935,N_31005);
xor U32322 (N_32322,N_31018,N_31706);
and U32323 (N_32323,N_30291,N_30430);
and U32324 (N_32324,N_30271,N_30681);
or U32325 (N_32325,N_31464,N_31876);
xnor U32326 (N_32326,N_30976,N_30374);
xor U32327 (N_32327,N_31619,N_30000);
xnor U32328 (N_32328,N_30951,N_30254);
and U32329 (N_32329,N_31736,N_31737);
and U32330 (N_32330,N_30478,N_30582);
xnor U32331 (N_32331,N_31284,N_31989);
nand U32332 (N_32332,N_31957,N_31242);
or U32333 (N_32333,N_30567,N_31428);
xor U32334 (N_32334,N_31694,N_31806);
nand U32335 (N_32335,N_31580,N_30943);
and U32336 (N_32336,N_30338,N_31586);
nor U32337 (N_32337,N_31012,N_31906);
or U32338 (N_32338,N_31431,N_30166);
nor U32339 (N_32339,N_30451,N_30595);
and U32340 (N_32340,N_30469,N_30237);
and U32341 (N_32341,N_30097,N_31754);
xnor U32342 (N_32342,N_30577,N_30611);
or U32343 (N_32343,N_31823,N_30878);
and U32344 (N_32344,N_30793,N_31129);
or U32345 (N_32345,N_31163,N_30300);
and U32346 (N_32346,N_31011,N_31549);
xnor U32347 (N_32347,N_30591,N_31003);
xor U32348 (N_32348,N_30016,N_31411);
xor U32349 (N_32349,N_31893,N_31976);
nand U32350 (N_32350,N_31492,N_31528);
nand U32351 (N_32351,N_30022,N_30802);
and U32352 (N_32352,N_31161,N_31160);
or U32353 (N_32353,N_31475,N_31788);
nand U32354 (N_32354,N_31792,N_31789);
nor U32355 (N_32355,N_31592,N_30643);
or U32356 (N_32356,N_30383,N_31056);
and U32357 (N_32357,N_30773,N_30728);
nor U32358 (N_32358,N_30924,N_30856);
xor U32359 (N_32359,N_30696,N_30102);
nor U32360 (N_32360,N_30600,N_31157);
and U32361 (N_32361,N_30012,N_30425);
and U32362 (N_32362,N_31950,N_30104);
or U32363 (N_32363,N_31394,N_31671);
nand U32364 (N_32364,N_31712,N_30155);
xnor U32365 (N_32365,N_30281,N_31042);
and U32366 (N_32366,N_30409,N_30389);
nor U32367 (N_32367,N_31618,N_31022);
nand U32368 (N_32368,N_31638,N_31330);
nor U32369 (N_32369,N_30922,N_30125);
and U32370 (N_32370,N_31912,N_31213);
or U32371 (N_32371,N_31884,N_31127);
xor U32372 (N_32372,N_31637,N_31542);
nand U32373 (N_32373,N_30255,N_30426);
xor U32374 (N_32374,N_31830,N_30040);
or U32375 (N_32375,N_31350,N_31925);
and U32376 (N_32376,N_31148,N_30106);
nor U32377 (N_32377,N_30768,N_31553);
nand U32378 (N_32378,N_31096,N_31128);
and U32379 (N_32379,N_31948,N_31799);
and U32380 (N_32380,N_31953,N_31627);
xor U32381 (N_32381,N_31423,N_31341);
nor U32382 (N_32382,N_30051,N_31887);
xor U32383 (N_32383,N_30605,N_30950);
or U32384 (N_32384,N_31963,N_31369);
or U32385 (N_32385,N_30421,N_31510);
nor U32386 (N_32386,N_30424,N_31150);
nand U32387 (N_32387,N_30092,N_31930);
xor U32388 (N_32388,N_31201,N_30552);
xor U32389 (N_32389,N_30808,N_30109);
xor U32390 (N_32390,N_30941,N_31702);
and U32391 (N_32391,N_31332,N_30189);
nor U32392 (N_32392,N_31764,N_31045);
and U32393 (N_32393,N_30231,N_30722);
and U32394 (N_32394,N_30692,N_31802);
xor U32395 (N_32395,N_31784,N_30137);
nor U32396 (N_32396,N_31155,N_30958);
nor U32397 (N_32397,N_31406,N_31527);
and U32398 (N_32398,N_31777,N_31857);
nor U32399 (N_32399,N_31732,N_31482);
nor U32400 (N_32400,N_31546,N_31832);
or U32401 (N_32401,N_30452,N_30873);
or U32402 (N_32402,N_30787,N_30405);
xor U32403 (N_32403,N_31495,N_31507);
nand U32404 (N_32404,N_30818,N_30372);
xor U32405 (N_32405,N_30417,N_30184);
nand U32406 (N_32406,N_30763,N_31842);
or U32407 (N_32407,N_30423,N_30672);
nand U32408 (N_32408,N_30130,N_30743);
nand U32409 (N_32409,N_30388,N_30833);
or U32410 (N_32410,N_30797,N_31916);
or U32411 (N_32411,N_30176,N_30520);
nand U32412 (N_32412,N_30545,N_31924);
nor U32413 (N_32413,N_30187,N_30850);
xor U32414 (N_32414,N_31066,N_31606);
nand U32415 (N_32415,N_31357,N_31995);
and U32416 (N_32416,N_30441,N_30604);
or U32417 (N_32417,N_31231,N_30063);
and U32418 (N_32418,N_31755,N_30282);
or U32419 (N_32419,N_31036,N_31111);
nand U32420 (N_32420,N_30750,N_31147);
or U32421 (N_32421,N_30741,N_31713);
xor U32422 (N_32422,N_30174,N_31711);
xor U32423 (N_32423,N_30375,N_30170);
and U32424 (N_32424,N_30460,N_30669);
nand U32425 (N_32425,N_31548,N_30440);
and U32426 (N_32426,N_31166,N_30912);
nand U32427 (N_32427,N_31254,N_31991);
nand U32428 (N_32428,N_31524,N_30638);
xnor U32429 (N_32429,N_31663,N_30815);
nand U32430 (N_32430,N_30444,N_30352);
xor U32431 (N_32431,N_30183,N_30946);
nand U32432 (N_32432,N_30080,N_31578);
nand U32433 (N_32433,N_31202,N_30619);
or U32434 (N_32434,N_31141,N_30265);
xnor U32435 (N_32435,N_31440,N_31258);
nor U32436 (N_32436,N_30558,N_30151);
xor U32437 (N_32437,N_31599,N_31651);
nand U32438 (N_32438,N_31591,N_31211);
xor U32439 (N_32439,N_31834,N_31817);
nand U32440 (N_32440,N_30720,N_30986);
nor U32441 (N_32441,N_30442,N_31104);
xor U32442 (N_32442,N_31031,N_30705);
xnor U32443 (N_32443,N_30644,N_30500);
nand U32444 (N_32444,N_30969,N_30569);
or U32445 (N_32445,N_31130,N_31391);
nand U32446 (N_32446,N_31486,N_30009);
and U32447 (N_32447,N_31365,N_30341);
xor U32448 (N_32448,N_31555,N_31587);
nand U32449 (N_32449,N_31466,N_30892);
nand U32450 (N_32450,N_31460,N_31137);
or U32451 (N_32451,N_30782,N_31731);
and U32452 (N_32452,N_31116,N_31028);
xor U32453 (N_32453,N_31230,N_30953);
xor U32454 (N_32454,N_30295,N_31273);
or U32455 (N_32455,N_31829,N_31088);
nor U32456 (N_32456,N_31645,N_30356);
or U32457 (N_32457,N_31280,N_30359);
nor U32458 (N_32458,N_30323,N_31739);
and U32459 (N_32459,N_31164,N_31058);
nand U32460 (N_32460,N_30204,N_30221);
or U32461 (N_32461,N_31573,N_31302);
or U32462 (N_32462,N_30278,N_31470);
xnor U32463 (N_32463,N_31985,N_31577);
and U32464 (N_32464,N_31353,N_30684);
nand U32465 (N_32465,N_30304,N_31506);
xor U32466 (N_32466,N_30508,N_31968);
nor U32467 (N_32467,N_31820,N_30393);
or U32468 (N_32468,N_30972,N_31480);
xnor U32469 (N_32469,N_31255,N_30571);
nand U32470 (N_32470,N_30887,N_30053);
and U32471 (N_32471,N_31597,N_30985);
xor U32472 (N_32472,N_31807,N_30991);
and U32473 (N_32473,N_31383,N_30553);
xor U32474 (N_32474,N_30085,N_31557);
or U32475 (N_32475,N_31707,N_31378);
and U32476 (N_32476,N_30994,N_31143);
or U32477 (N_32477,N_31641,N_31779);
or U32478 (N_32478,N_30507,N_30707);
nor U32479 (N_32479,N_31309,N_31297);
nand U32480 (N_32480,N_31471,N_30289);
or U32481 (N_32481,N_30585,N_31856);
or U32482 (N_32482,N_31477,N_31132);
nand U32483 (N_32483,N_31699,N_31206);
nand U32484 (N_32484,N_30132,N_30210);
and U32485 (N_32485,N_30908,N_31498);
and U32486 (N_32486,N_30497,N_30636);
nand U32487 (N_32487,N_30348,N_31241);
nor U32488 (N_32488,N_31030,N_30261);
nor U32489 (N_32489,N_31519,N_31596);
nor U32490 (N_32490,N_30107,N_31626);
xnor U32491 (N_32491,N_31296,N_30995);
or U32492 (N_32492,N_31292,N_30891);
or U32493 (N_32493,N_30932,N_31261);
or U32494 (N_32494,N_30207,N_31035);
nor U32495 (N_32495,N_30601,N_31151);
nor U32496 (N_32496,N_31656,N_31878);
or U32497 (N_32497,N_30492,N_31180);
xor U32498 (N_32498,N_30228,N_30729);
xor U32499 (N_32499,N_31881,N_30535);
nor U32500 (N_32500,N_31667,N_30477);
and U32501 (N_32501,N_31229,N_31844);
or U32502 (N_32502,N_30382,N_31620);
or U32503 (N_32503,N_31662,N_31653);
nor U32504 (N_32504,N_30821,N_31822);
nand U32505 (N_32505,N_30973,N_30791);
xnor U32506 (N_32506,N_31074,N_31697);
and U32507 (N_32507,N_30258,N_31305);
and U32508 (N_32508,N_31225,N_30927);
xor U32509 (N_32509,N_30071,N_31942);
or U32510 (N_32510,N_31536,N_30633);
xor U32511 (N_32511,N_30103,N_31053);
nor U32512 (N_32512,N_31772,N_30679);
or U32513 (N_32513,N_30379,N_31996);
xnor U32514 (N_32514,N_31345,N_31794);
or U32515 (N_32515,N_31485,N_31955);
xnor U32516 (N_32516,N_31315,N_31371);
nor U32517 (N_32517,N_30624,N_31811);
or U32518 (N_32518,N_31927,N_31840);
or U32519 (N_32519,N_30573,N_30325);
and U32520 (N_32520,N_30517,N_31877);
and U32521 (N_32521,N_31689,N_31581);
and U32522 (N_32522,N_31149,N_31529);
and U32523 (N_32523,N_30324,N_31377);
or U32524 (N_32524,N_30161,N_30536);
xor U32525 (N_32525,N_30437,N_31721);
nor U32526 (N_32526,N_31270,N_30299);
and U32527 (N_32527,N_30992,N_30391);
or U32528 (N_32528,N_30385,N_31187);
nand U32529 (N_32529,N_31563,N_30527);
xor U32530 (N_32530,N_31907,N_30693);
or U32531 (N_32531,N_30716,N_31348);
xnor U32532 (N_32532,N_30004,N_30464);
nand U32533 (N_32533,N_30780,N_31513);
xor U32534 (N_32534,N_31920,N_30002);
nor U32535 (N_32535,N_30398,N_30205);
or U32536 (N_32536,N_30664,N_30883);
and U32537 (N_32537,N_30283,N_30979);
or U32538 (N_32538,N_30607,N_31055);
and U32539 (N_32539,N_31300,N_30394);
nand U32540 (N_32540,N_31162,N_31608);
and U32541 (N_32541,N_31622,N_30907);
xor U32542 (N_32542,N_30163,N_31729);
or U32543 (N_32543,N_31468,N_30381);
xor U32544 (N_32544,N_31253,N_30756);
and U32545 (N_32545,N_31771,N_30070);
nand U32546 (N_32546,N_31298,N_31335);
nand U32547 (N_32547,N_31386,N_30964);
and U32548 (N_32548,N_31354,N_31917);
nand U32549 (N_32549,N_31610,N_31681);
or U32550 (N_32550,N_31521,N_30574);
nor U32551 (N_32551,N_31775,N_31168);
xor U32552 (N_32552,N_30030,N_30357);
or U32553 (N_32553,N_31338,N_31023);
xnor U32554 (N_32554,N_30143,N_30622);
nand U32555 (N_32555,N_30809,N_30678);
xor U32556 (N_32556,N_31034,N_31683);
or U32557 (N_32557,N_30011,N_31569);
or U32558 (N_32558,N_31715,N_31478);
or U32559 (N_32559,N_30770,N_30229);
nand U32560 (N_32560,N_31445,N_31828);
xor U32561 (N_32561,N_30367,N_30428);
xnor U32562 (N_32562,N_31797,N_30333);
or U32563 (N_32563,N_30279,N_30532);
xor U32564 (N_32564,N_30159,N_31747);
and U32565 (N_32565,N_30369,N_30313);
and U32566 (N_32566,N_31175,N_30834);
nand U32567 (N_32567,N_30363,N_30934);
xor U32568 (N_32568,N_30005,N_31838);
xnor U32569 (N_32569,N_31743,N_31176);
nand U32570 (N_32570,N_31813,N_31940);
or U32571 (N_32571,N_31670,N_31115);
and U32572 (N_32572,N_30665,N_31093);
nor U32573 (N_32573,N_30447,N_30494);
xor U32574 (N_32574,N_31882,N_31009);
nor U32575 (N_32575,N_30549,N_31848);
and U32576 (N_32576,N_31328,N_31658);
nor U32577 (N_32577,N_31210,N_31159);
or U32578 (N_32578,N_30267,N_30733);
or U32579 (N_32579,N_31904,N_30100);
and U32580 (N_32580,N_30851,N_30859);
nand U32581 (N_32581,N_31200,N_30008);
or U32582 (N_32582,N_30058,N_30122);
nand U32583 (N_32583,N_31585,N_30674);
nand U32584 (N_32584,N_30014,N_31094);
nor U32585 (N_32585,N_31193,N_30355);
and U32586 (N_32586,N_30473,N_31401);
nand U32587 (N_32587,N_30583,N_30365);
nor U32588 (N_32588,N_31312,N_30195);
nand U32589 (N_32589,N_30302,N_31246);
or U32590 (N_32590,N_31682,N_30501);
nand U32591 (N_32591,N_30906,N_30881);
xnor U32592 (N_32592,N_31217,N_31481);
or U32593 (N_32593,N_30504,N_31833);
nand U32594 (N_32594,N_30735,N_30110);
and U32595 (N_32595,N_30942,N_31749);
nand U32596 (N_32596,N_30472,N_31522);
xnor U32597 (N_32597,N_30093,N_30123);
and U32598 (N_32598,N_31901,N_31146);
or U32599 (N_32599,N_31717,N_30785);
and U32600 (N_32600,N_31487,N_31818);
xor U32601 (N_32601,N_31277,N_31783);
or U32602 (N_32602,N_31208,N_31765);
nor U32603 (N_32603,N_30683,N_30560);
xor U32604 (N_32604,N_31461,N_31366);
or U32605 (N_32605,N_30842,N_30732);
nand U32606 (N_32606,N_31384,N_31051);
nor U32607 (N_32607,N_30245,N_30407);
xor U32608 (N_32608,N_31846,N_30347);
nor U32609 (N_32609,N_31122,N_31987);
nor U32610 (N_32610,N_31692,N_30411);
xnor U32611 (N_32611,N_30259,N_31235);
or U32612 (N_32612,N_30826,N_30503);
nor U32613 (N_32613,N_30795,N_31195);
or U32614 (N_32614,N_30043,N_30196);
nand U32615 (N_32615,N_31433,N_31364);
and U32616 (N_32616,N_30165,N_30847);
or U32617 (N_32617,N_31545,N_30171);
or U32618 (N_32618,N_30127,N_30689);
and U32619 (N_32619,N_31853,N_30849);
and U32620 (N_32620,N_31938,N_30746);
and U32621 (N_32621,N_30813,N_30792);
and U32622 (N_32622,N_30073,N_30710);
or U32623 (N_32623,N_30955,N_30146);
xor U32624 (N_32624,N_30896,N_30845);
nor U32625 (N_32625,N_30410,N_30564);
or U32626 (N_32626,N_31203,N_31398);
nand U32627 (N_32627,N_31601,N_30831);
or U32628 (N_32628,N_30111,N_30587);
xnor U32629 (N_32629,N_31285,N_30653);
and U32630 (N_32630,N_30727,N_31534);
xnor U32631 (N_32631,N_30243,N_31914);
and U32632 (N_32632,N_30566,N_31538);
and U32633 (N_32633,N_30129,N_30998);
nand U32634 (N_32634,N_31724,N_30543);
nand U32635 (N_32635,N_30308,N_30117);
nand U32636 (N_32636,N_30286,N_30764);
nand U32637 (N_32637,N_31493,N_31069);
xor U32638 (N_32638,N_31156,N_30087);
or U32639 (N_32639,N_30776,N_31570);
or U32640 (N_32640,N_30079,N_30354);
nand U32641 (N_32641,N_30118,N_31439);
nand U32642 (N_32642,N_30266,N_30687);
and U32643 (N_32643,N_30029,N_31603);
nor U32644 (N_32644,N_31900,N_30544);
xor U32645 (N_32645,N_31319,N_30897);
nand U32646 (N_32646,N_31750,N_31970);
nor U32647 (N_32647,N_30781,N_30634);
and U32648 (N_32648,N_30983,N_31407);
nand U32649 (N_32649,N_30236,N_30794);
nor U32650 (N_32650,N_31279,N_31082);
nand U32651 (N_32651,N_30987,N_30490);
nand U32652 (N_32652,N_30419,N_31994);
nand U32653 (N_32653,N_31379,N_31589);
nand U32654 (N_32654,N_31701,N_30940);
or U32655 (N_32655,N_31172,N_31216);
xor U32656 (N_32656,N_31514,N_31219);
xnor U32657 (N_32657,N_31855,N_31170);
nor U32658 (N_32658,N_31091,N_30126);
nor U32659 (N_32659,N_30457,N_30990);
nor U32660 (N_32660,N_30412,N_30670);
nand U32661 (N_32661,N_30509,N_31084);
and U32662 (N_32662,N_31138,N_30697);
and U32663 (N_32663,N_30350,N_31108);
or U32664 (N_32664,N_31479,N_31984);
and U32665 (N_32665,N_31567,N_31633);
and U32666 (N_32666,N_31761,N_31568);
nor U32667 (N_32667,N_30119,N_31558);
xor U32668 (N_32668,N_30886,N_30402);
or U32669 (N_32669,N_31562,N_31690);
nor U32670 (N_32670,N_30025,N_30026);
and U32671 (N_32671,N_30812,N_30981);
or U32672 (N_32672,N_30095,N_30179);
and U32673 (N_32673,N_30673,N_31661);
nor U32674 (N_32674,N_30191,N_30173);
nor U32675 (N_32675,N_31532,N_30238);
or U32676 (N_32676,N_31021,N_31520);
and U32677 (N_32677,N_31752,N_31427);
and U32678 (N_32678,N_30888,N_30531);
or U32679 (N_32679,N_31179,N_31459);
nand U32680 (N_32680,N_31393,N_30445);
nor U32681 (N_32681,N_30561,N_31075);
nand U32682 (N_32682,N_31410,N_30377);
nor U32683 (N_32683,N_30307,N_31600);
and U32684 (N_32684,N_31517,N_30169);
or U32685 (N_32685,N_30525,N_31247);
nor U32686 (N_32686,N_31167,N_30807);
nand U32687 (N_32687,N_31760,N_31790);
xnor U32688 (N_32688,N_31609,N_31289);
nor U32689 (N_32689,N_30403,N_31165);
xnor U32690 (N_32690,N_31243,N_31630);
and U32691 (N_32691,N_30522,N_30540);
and U32692 (N_32692,N_30392,N_30789);
nand U32693 (N_32693,N_30113,N_30784);
or U32694 (N_32694,N_30276,N_30884);
nor U32695 (N_32695,N_30018,N_31324);
nand U32696 (N_32696,N_31745,N_30563);
nand U32697 (N_32697,N_30301,N_30803);
nand U32698 (N_32698,N_31782,N_31918);
nand U32699 (N_32699,N_31303,N_31215);
nor U32700 (N_32700,N_30971,N_30257);
or U32701 (N_32701,N_30003,N_31751);
nor U32702 (N_32702,N_31248,N_31537);
nor U32703 (N_32703,N_30528,N_30835);
nor U32704 (N_32704,N_30612,N_31072);
nor U32705 (N_32705,N_31044,N_31154);
or U32706 (N_32706,N_30524,N_30150);
and U32707 (N_32707,N_30836,N_31087);
nor U32708 (N_32708,N_31698,N_30368);
and U32709 (N_32709,N_30970,N_30474);
nand U32710 (N_32710,N_30755,N_30744);
or U32711 (N_32711,N_30688,N_31250);
nor U32712 (N_32712,N_30021,N_31327);
xor U32713 (N_32713,N_30175,N_30855);
nand U32714 (N_32714,N_31063,N_31693);
nand U32715 (N_32715,N_31515,N_31291);
or U32716 (N_32716,N_30975,N_30498);
and U32717 (N_32717,N_31748,N_31852);
nor U32718 (N_32718,N_31251,N_30709);
xor U32719 (N_32719,N_30956,N_30846);
and U32720 (N_32720,N_31773,N_31583);
xnor U32721 (N_32721,N_30148,N_31306);
or U32722 (N_32722,N_30719,N_30138);
and U32723 (N_32723,N_30651,N_31616);
and U32724 (N_32724,N_30036,N_30076);
xor U32725 (N_32725,N_30799,N_30277);
and U32726 (N_32726,N_30059,N_30646);
and U32727 (N_32727,N_31770,N_31002);
xnor U32728 (N_32728,N_30869,N_30936);
nor U32729 (N_32729,N_30370,N_31112);
xor U32730 (N_32730,N_31705,N_31491);
nand U32731 (N_32731,N_31759,N_30450);
or U32732 (N_32732,N_31043,N_30401);
xor U32733 (N_32733,N_30481,N_31404);
and U32734 (N_32734,N_31902,N_31090);
and U32735 (N_32735,N_30534,N_30609);
nand U32736 (N_32736,N_30931,N_30212);
or U32737 (N_32737,N_30147,N_30091);
or U32738 (N_32738,N_30203,N_31007);
nand U32739 (N_32739,N_30589,N_30860);
xor U32740 (N_32740,N_30639,N_31010);
or U32741 (N_32741,N_30476,N_30610);
nor U32742 (N_32742,N_31774,N_31530);
and U32743 (N_32743,N_31076,N_31503);
nor U32744 (N_32744,N_30326,N_30251);
or U32745 (N_32745,N_30718,N_30613);
or U32746 (N_32746,N_31575,N_31004);
xor U32747 (N_32747,N_31696,N_31865);
nor U32748 (N_32748,N_31256,N_30913);
xor U32749 (N_32749,N_30617,N_31121);
or U32750 (N_32750,N_30328,N_30064);
nand U32751 (N_32751,N_30007,N_30676);
and U32752 (N_32752,N_30422,N_31951);
and U32753 (N_32753,N_30121,N_31131);
nand U32754 (N_32754,N_31448,N_30225);
nor U32755 (N_32755,N_31041,N_31117);
nor U32756 (N_32756,N_30065,N_31954);
nor U32757 (N_32757,N_30458,N_30340);
nand U32758 (N_32758,N_30215,N_30748);
nand U32759 (N_32759,N_30072,N_30661);
or U32760 (N_32760,N_30930,N_31804);
nor U32761 (N_32761,N_30642,N_30706);
nor U32762 (N_32762,N_30898,N_31057);
and U32763 (N_32763,N_31533,N_31526);
xor U32764 (N_32764,N_31336,N_31861);
and U32765 (N_32765,N_30547,N_30310);
xor U32766 (N_32766,N_31980,N_31888);
or U32767 (N_32767,N_30680,N_31978);
nor U32768 (N_32768,N_31257,N_31565);
xor U32769 (N_32769,N_30420,N_31214);
nand U32770 (N_32770,N_31450,N_31421);
or U32771 (N_32771,N_30088,N_30562);
xor U32772 (N_32772,N_31186,N_30749);
and U32773 (N_32773,N_30854,N_30269);
and U32774 (N_32774,N_31664,N_31588);
xor U32775 (N_32775,N_31908,N_31617);
and U32776 (N_32776,N_30820,N_31972);
nand U32777 (N_32777,N_31451,N_31271);
xnor U32778 (N_32778,N_30905,N_31554);
xor U32779 (N_32779,N_31178,N_31016);
and U32780 (N_32780,N_31961,N_30668);
xnor U32781 (N_32781,N_31719,N_31363);
nor U32782 (N_32782,N_30993,N_30094);
xnor U32783 (N_32783,N_31974,N_30606);
and U32784 (N_32784,N_31252,N_31339);
nor U32785 (N_32785,N_30630,N_31665);
xnor U32786 (N_32786,N_31321,N_30910);
nand U32787 (N_32787,N_31550,N_31020);
nand U32788 (N_32788,N_30061,N_31207);
nor U32789 (N_32789,N_30162,N_30899);
xor U32790 (N_32790,N_31126,N_30360);
xor U32791 (N_32791,N_31092,N_30939);
xor U32792 (N_32792,N_30572,N_30060);
nand U32793 (N_32793,N_31766,N_30487);
nand U32794 (N_32794,N_31614,N_30510);
nor U32795 (N_32795,N_31880,N_30139);
or U32796 (N_32796,N_31988,N_31437);
nor U32797 (N_32797,N_31399,N_30345);
nor U32798 (N_32798,N_30963,N_30120);
xor U32799 (N_32799,N_31135,N_30917);
and U32800 (N_32800,N_30880,N_31268);
nor U32801 (N_32801,N_30505,N_31574);
nor U32802 (N_32802,N_31333,N_30514);
or U32803 (N_32803,N_31668,N_31173);
nor U32804 (N_32804,N_30293,N_30628);
nand U32805 (N_32805,N_31858,N_30811);
or U32806 (N_32806,N_31576,N_30234);
or U32807 (N_32807,N_31756,N_31648);
xor U32808 (N_32808,N_30614,N_31081);
xor U32809 (N_32809,N_31602,N_30235);
and U32810 (N_32810,N_31903,N_30584);
xnor U32811 (N_32811,N_31006,N_31171);
or U32812 (N_32812,N_30596,N_30318);
or U32813 (N_32813,N_31101,N_30996);
nand U32814 (N_32814,N_31845,N_30751);
nand U32815 (N_32815,N_30603,N_30691);
or U32816 (N_32816,N_31753,N_30311);
nor U32817 (N_32817,N_30032,N_30438);
or U32818 (N_32818,N_30702,N_31140);
xnor U32819 (N_32819,N_30740,N_30034);
and U32820 (N_32820,N_31473,N_31197);
nand U32821 (N_32821,N_30715,N_30593);
nand U32822 (N_32822,N_31337,N_30523);
nor U32823 (N_32823,N_30866,N_31474);
and U32824 (N_32824,N_30384,N_31500);
or U32825 (N_32825,N_30128,N_31814);
nor U32826 (N_32826,N_30337,N_30928);
nor U32827 (N_32827,N_30666,N_31446);
and U32828 (N_32828,N_31228,N_30001);
and U32829 (N_32829,N_30416,N_30491);
nor U32830 (N_32830,N_31189,N_30959);
nand U32831 (N_32831,N_31975,N_31669);
nor U32832 (N_32832,N_30753,N_31038);
xor U32833 (N_32833,N_30885,N_31965);
or U32834 (N_32834,N_30468,N_30658);
xnor U32835 (N_32835,N_31584,N_30465);
nand U32836 (N_32836,N_31397,N_31061);
or U32837 (N_32837,N_31233,N_31869);
or U32838 (N_32838,N_31776,N_30268);
nor U32839 (N_32839,N_31114,N_31105);
or U32840 (N_32840,N_30832,N_31125);
or U32841 (N_32841,N_31422,N_31921);
nor U32842 (N_32842,N_30759,N_30752);
or U32843 (N_32843,N_30217,N_30049);
or U32844 (N_32844,N_30288,N_31543);
nor U32845 (N_32845,N_31695,N_31223);
and U32846 (N_32846,N_31919,N_31722);
or U32847 (N_32847,N_31356,N_30134);
nor U32848 (N_32848,N_30758,N_30017);
nor U32849 (N_32849,N_30343,N_31875);
or U32850 (N_32850,N_31484,N_30224);
nand U32851 (N_32851,N_30538,N_31059);
nand U32852 (N_32852,N_31986,N_30570);
or U32853 (N_32853,N_31744,N_30879);
nand U32854 (N_32854,N_30273,N_30911);
nand U32855 (N_32855,N_31033,N_30841);
or U32856 (N_32856,N_30695,N_30461);
nor U32857 (N_32857,N_30620,N_31716);
nor U32858 (N_32858,N_30044,N_30837);
and U32859 (N_32859,N_30397,N_31085);
nand U32860 (N_32860,N_31640,N_31932);
nand U32861 (N_32861,N_30961,N_31564);
nand U32862 (N_32862,N_31039,N_31595);
nand U32863 (N_32863,N_30342,N_30054);
xnor U32864 (N_32864,N_31873,N_30376);
nor U32865 (N_32865,N_30142,N_30648);
xor U32866 (N_32866,N_30400,N_30353);
nor U32867 (N_32867,N_31734,N_31944);
xor U32868 (N_32868,N_30272,N_30902);
xor U32869 (N_32869,N_31029,N_30765);
or U32870 (N_32870,N_30380,N_30219);
nor U32871 (N_32871,N_31809,N_30988);
or U32872 (N_32872,N_30872,N_30193);
and U32873 (N_32873,N_31078,N_31351);
or U32874 (N_32874,N_30944,N_31723);
and U32875 (N_32875,N_31438,N_30790);
nor U32876 (N_32876,N_30712,N_31409);
or U32877 (N_32877,N_30757,N_30843);
or U32878 (N_32878,N_30154,N_30349);
and U32879 (N_32879,N_30488,N_30336);
xor U32880 (N_32880,N_31544,N_30775);
and U32881 (N_32881,N_30949,N_30862);
or U32882 (N_32882,N_31778,N_31370);
or U32883 (N_32883,N_30541,N_31458);
or U32884 (N_32884,N_31505,N_30334);
and U32885 (N_32885,N_30449,N_31239);
xnor U32886 (N_32886,N_31425,N_30240);
nor U32887 (N_32887,N_31299,N_30351);
nand U32888 (N_32888,N_31320,N_31318);
nand U32889 (N_32889,N_30516,N_31040);
and U32890 (N_32890,N_31885,N_30662);
xor U32891 (N_32891,N_30966,N_30413);
and U32892 (N_32892,N_30432,N_31612);
xnor U32893 (N_32893,N_31435,N_30309);
nor U32894 (N_32894,N_31851,N_31098);
nor U32895 (N_32895,N_30954,N_31871);
nand U32896 (N_32896,N_30192,N_30829);
and U32897 (N_32897,N_31922,N_31457);
nand U32898 (N_32898,N_31825,N_31561);
or U32899 (N_32899,N_30711,N_30157);
xnor U32900 (N_32900,N_30590,N_31355);
or U32901 (N_32901,N_31704,N_31539);
nor U32902 (N_32902,N_31827,N_30284);
nand U32903 (N_32903,N_30223,N_30099);
nor U32904 (N_32904,N_30515,N_31329);
or U32905 (N_32905,N_30226,N_31281);
nor U32906 (N_32906,N_31525,N_31934);
xor U32907 (N_32907,N_30248,N_31905);
or U32908 (N_32908,N_31652,N_31839);
nand U32909 (N_32909,N_31416,N_31065);
xor U32910 (N_32910,N_31462,N_31860);
nor U32911 (N_32911,N_30703,N_30280);
and U32912 (N_32912,N_30249,N_31872);
xnor U32913 (N_32913,N_30408,N_30779);
nor U32914 (N_32914,N_30853,N_30475);
and U32915 (N_32915,N_30786,N_30395);
or U32916 (N_32916,N_31110,N_31344);
and U32917 (N_32917,N_31376,N_31966);
nor U32918 (N_32918,N_30952,N_31249);
and U32919 (N_32919,N_30700,N_31220);
nand U32920 (N_32920,N_31928,N_31192);
xor U32921 (N_32921,N_30581,N_30777);
xor U32922 (N_32922,N_30903,N_30414);
xnor U32923 (N_32923,N_30331,N_30893);
xnor U32924 (N_32924,N_30239,N_30078);
nor U32925 (N_32925,N_30242,N_31796);
nand U32926 (N_32926,N_31109,N_31343);
xor U32927 (N_32927,N_30645,N_31488);
nand U32928 (N_32928,N_30967,N_30042);
nor U32929 (N_32929,N_30962,N_30198);
and U32930 (N_32930,N_31540,N_31443);
nand U32931 (N_32931,N_30315,N_30701);
nor U32932 (N_32932,N_30164,N_30649);
xor U32933 (N_32933,N_31025,N_30530);
xnor U32934 (N_32934,N_31144,N_30521);
xor U32935 (N_32935,N_31212,N_31184);
xor U32936 (N_32936,N_30578,N_31444);
or U32937 (N_32937,N_31621,N_30819);
nor U32938 (N_32938,N_31993,N_30933);
and U32939 (N_32939,N_31874,N_31152);
nor U32940 (N_32940,N_30559,N_30327);
nor U32941 (N_32941,N_30453,N_30945);
or U32942 (N_32942,N_31050,N_30876);
xnor U32943 (N_32943,N_31095,N_31684);
or U32944 (N_32944,N_31037,N_31361);
and U32945 (N_32945,N_31237,N_31676);
nand U32946 (N_32946,N_31791,N_31931);
or U32947 (N_32947,N_31999,N_30877);
or U32948 (N_32948,N_30294,N_30250);
or U32949 (N_32949,N_31678,N_31469);
nor U32950 (N_32950,N_30895,N_30244);
xnor U32951 (N_32951,N_31334,N_31071);
nand U32952 (N_32952,N_30247,N_30857);
and U32953 (N_32953,N_30320,N_30556);
xor U32954 (N_32954,N_31708,N_30852);
and U32955 (N_32955,N_31346,N_30717);
nand U32956 (N_32956,N_30062,N_31387);
nand U32957 (N_32957,N_31199,N_30013);
nand U32958 (N_32958,N_31405,N_31835);
and U32959 (N_32959,N_31512,N_30948);
nor U32960 (N_32960,N_30659,N_31209);
xnor U32961 (N_32961,N_30921,N_30615);
and U32962 (N_32962,N_30742,N_31196);
and U32963 (N_32963,N_30489,N_30486);
nand U32964 (N_32964,N_30863,N_31499);
or U32965 (N_32965,N_30984,N_31943);
xor U32966 (N_32966,N_31136,N_31272);
xnor U32967 (N_32967,N_31120,N_31971);
or U32968 (N_32968,N_31964,N_30371);
and U32969 (N_32969,N_30935,N_30463);
and U32970 (N_32970,N_30621,N_31224);
nand U32971 (N_32971,N_31998,N_30926);
nor U32972 (N_32972,N_30387,N_30816);
nor U32973 (N_32973,N_30306,N_31720);
nand U32974 (N_32974,N_31436,N_31388);
nor U32975 (N_32975,N_31786,N_31014);
nor U32976 (N_32976,N_30997,N_31181);
nor U32977 (N_32977,N_30454,N_31879);
or U32978 (N_32978,N_31139,N_31990);
xnor U32979 (N_32979,N_31611,N_30466);
and U32980 (N_32980,N_31805,N_31375);
nand U32981 (N_32981,N_30067,N_30599);
xnor U32982 (N_32982,N_31511,N_30027);
and U32983 (N_32983,N_30760,N_30865);
or U32984 (N_32984,N_31400,N_31947);
nand U32985 (N_32985,N_31097,N_30598);
xnor U32986 (N_32986,N_30557,N_31145);
and U32987 (N_32987,N_31047,N_30431);
xnor U32988 (N_32988,N_30675,N_30124);
and U32989 (N_32989,N_30900,N_30761);
nor U32990 (N_32990,N_31812,N_31017);
or U32991 (N_32991,N_30686,N_30822);
or U32992 (N_32992,N_31368,N_30429);
nand U32993 (N_32993,N_31673,N_30656);
and U32994 (N_32994,N_30015,N_30708);
or U32995 (N_32995,N_31992,N_30483);
and U32996 (N_32996,N_30332,N_31598);
nand U32997 (N_32997,N_30551,N_31501);
nor U32998 (N_32998,N_30090,N_31936);
xor U32999 (N_32999,N_31226,N_30479);
nor U33000 (N_33000,N_30658,N_30145);
and U33001 (N_33001,N_31993,N_31142);
nand U33002 (N_33002,N_31017,N_30798);
and U33003 (N_33003,N_31773,N_30661);
nor U33004 (N_33004,N_30837,N_30664);
or U33005 (N_33005,N_31933,N_31163);
nand U33006 (N_33006,N_31970,N_30259);
xnor U33007 (N_33007,N_31632,N_31382);
xnor U33008 (N_33008,N_31529,N_30799);
xnor U33009 (N_33009,N_31636,N_31691);
nand U33010 (N_33010,N_31142,N_30619);
nand U33011 (N_33011,N_31399,N_30104);
and U33012 (N_33012,N_31250,N_31541);
and U33013 (N_33013,N_31333,N_31547);
and U33014 (N_33014,N_31894,N_30310);
nand U33015 (N_33015,N_30614,N_30260);
or U33016 (N_33016,N_31037,N_31557);
xnor U33017 (N_33017,N_31856,N_31045);
and U33018 (N_33018,N_31928,N_31128);
and U33019 (N_33019,N_30596,N_31548);
nand U33020 (N_33020,N_31084,N_30768);
or U33021 (N_33021,N_30641,N_30935);
xnor U33022 (N_33022,N_31547,N_30435);
nor U33023 (N_33023,N_30430,N_31063);
and U33024 (N_33024,N_31488,N_30383);
nor U33025 (N_33025,N_31070,N_31783);
and U33026 (N_33026,N_31300,N_30142);
xnor U33027 (N_33027,N_31243,N_31428);
xnor U33028 (N_33028,N_31683,N_30631);
or U33029 (N_33029,N_30874,N_31142);
nor U33030 (N_33030,N_31639,N_30163);
nor U33031 (N_33031,N_30788,N_30256);
nor U33032 (N_33032,N_30151,N_31264);
xor U33033 (N_33033,N_31999,N_31715);
or U33034 (N_33034,N_31362,N_31233);
xor U33035 (N_33035,N_30880,N_31156);
xor U33036 (N_33036,N_31828,N_30986);
nor U33037 (N_33037,N_31501,N_30259);
and U33038 (N_33038,N_31245,N_31956);
nor U33039 (N_33039,N_31906,N_31274);
nor U33040 (N_33040,N_31586,N_31728);
nor U33041 (N_33041,N_30390,N_30066);
nor U33042 (N_33042,N_30810,N_30318);
nand U33043 (N_33043,N_30500,N_31331);
xor U33044 (N_33044,N_30440,N_31212);
xor U33045 (N_33045,N_30306,N_31134);
or U33046 (N_33046,N_31881,N_30177);
and U33047 (N_33047,N_30673,N_31822);
and U33048 (N_33048,N_31541,N_31602);
xnor U33049 (N_33049,N_31500,N_31488);
nand U33050 (N_33050,N_31944,N_31297);
xor U33051 (N_33051,N_30517,N_30262);
nor U33052 (N_33052,N_30839,N_30794);
xor U33053 (N_33053,N_31228,N_30568);
nand U33054 (N_33054,N_30367,N_30608);
nand U33055 (N_33055,N_31858,N_30672);
nor U33056 (N_33056,N_31621,N_30349);
nand U33057 (N_33057,N_30833,N_31774);
and U33058 (N_33058,N_30265,N_31825);
or U33059 (N_33059,N_30735,N_30169);
and U33060 (N_33060,N_31317,N_31541);
nand U33061 (N_33061,N_30212,N_30423);
nor U33062 (N_33062,N_30352,N_30962);
and U33063 (N_33063,N_30214,N_31447);
or U33064 (N_33064,N_31063,N_31252);
nand U33065 (N_33065,N_30171,N_31002);
or U33066 (N_33066,N_31319,N_31682);
xor U33067 (N_33067,N_30154,N_31719);
xnor U33068 (N_33068,N_31543,N_31951);
nor U33069 (N_33069,N_31692,N_31726);
or U33070 (N_33070,N_31502,N_30779);
and U33071 (N_33071,N_30136,N_31050);
and U33072 (N_33072,N_31364,N_31565);
and U33073 (N_33073,N_31510,N_31994);
or U33074 (N_33074,N_30617,N_31542);
xor U33075 (N_33075,N_31017,N_30852);
xor U33076 (N_33076,N_31860,N_31907);
nor U33077 (N_33077,N_31898,N_30450);
and U33078 (N_33078,N_31476,N_30761);
or U33079 (N_33079,N_30564,N_31472);
or U33080 (N_33080,N_30363,N_30221);
and U33081 (N_33081,N_31132,N_31000);
or U33082 (N_33082,N_30057,N_31280);
nor U33083 (N_33083,N_31625,N_30525);
and U33084 (N_33084,N_30944,N_30990);
and U33085 (N_33085,N_30350,N_30217);
nor U33086 (N_33086,N_30429,N_30761);
or U33087 (N_33087,N_31377,N_30899);
nand U33088 (N_33088,N_31000,N_31358);
nand U33089 (N_33089,N_31917,N_31454);
nor U33090 (N_33090,N_31962,N_30422);
or U33091 (N_33091,N_30308,N_30768);
or U33092 (N_33092,N_30563,N_30567);
xnor U33093 (N_33093,N_30272,N_30412);
or U33094 (N_33094,N_31995,N_31843);
or U33095 (N_33095,N_30036,N_31975);
xor U33096 (N_33096,N_30540,N_31444);
nand U33097 (N_33097,N_31481,N_31733);
and U33098 (N_33098,N_30461,N_30107);
nand U33099 (N_33099,N_30723,N_30760);
nand U33100 (N_33100,N_30047,N_31535);
nor U33101 (N_33101,N_31990,N_30240);
or U33102 (N_33102,N_31511,N_31519);
xor U33103 (N_33103,N_30260,N_30645);
xnor U33104 (N_33104,N_31498,N_31260);
or U33105 (N_33105,N_30564,N_31059);
nand U33106 (N_33106,N_30214,N_31789);
xor U33107 (N_33107,N_30859,N_31466);
nand U33108 (N_33108,N_31174,N_30429);
nand U33109 (N_33109,N_30908,N_31138);
xnor U33110 (N_33110,N_30997,N_30944);
nor U33111 (N_33111,N_31533,N_30751);
xor U33112 (N_33112,N_31320,N_30794);
xor U33113 (N_33113,N_31547,N_30602);
xnor U33114 (N_33114,N_30519,N_30373);
or U33115 (N_33115,N_31529,N_30602);
or U33116 (N_33116,N_31220,N_30115);
and U33117 (N_33117,N_30468,N_31237);
xnor U33118 (N_33118,N_30436,N_30863);
or U33119 (N_33119,N_31626,N_30913);
and U33120 (N_33120,N_30596,N_30885);
or U33121 (N_33121,N_31391,N_30071);
and U33122 (N_33122,N_31283,N_30858);
nand U33123 (N_33123,N_31631,N_30548);
and U33124 (N_33124,N_30574,N_31288);
nand U33125 (N_33125,N_30136,N_30770);
xor U33126 (N_33126,N_30099,N_31753);
xor U33127 (N_33127,N_31404,N_30003);
and U33128 (N_33128,N_31831,N_31923);
xor U33129 (N_33129,N_31587,N_31798);
nor U33130 (N_33130,N_31845,N_30575);
and U33131 (N_33131,N_30614,N_31350);
and U33132 (N_33132,N_31096,N_30072);
nand U33133 (N_33133,N_30204,N_30659);
and U33134 (N_33134,N_30856,N_30757);
xor U33135 (N_33135,N_31238,N_31283);
and U33136 (N_33136,N_30856,N_31747);
xor U33137 (N_33137,N_30975,N_30235);
nor U33138 (N_33138,N_31587,N_31962);
nand U33139 (N_33139,N_31419,N_31729);
xor U33140 (N_33140,N_31649,N_30841);
nand U33141 (N_33141,N_31407,N_31347);
or U33142 (N_33142,N_30583,N_31362);
nor U33143 (N_33143,N_30413,N_30115);
xor U33144 (N_33144,N_31959,N_30322);
nor U33145 (N_33145,N_31614,N_30498);
nor U33146 (N_33146,N_30484,N_30243);
nand U33147 (N_33147,N_30749,N_31967);
nor U33148 (N_33148,N_31458,N_30505);
or U33149 (N_33149,N_30193,N_30329);
or U33150 (N_33150,N_31558,N_31974);
and U33151 (N_33151,N_31158,N_30269);
xnor U33152 (N_33152,N_31368,N_30655);
and U33153 (N_33153,N_31716,N_31294);
nor U33154 (N_33154,N_30852,N_31819);
xnor U33155 (N_33155,N_30349,N_31838);
nor U33156 (N_33156,N_30755,N_31960);
or U33157 (N_33157,N_31933,N_30448);
nor U33158 (N_33158,N_30645,N_31671);
nor U33159 (N_33159,N_31552,N_30342);
nor U33160 (N_33160,N_30178,N_30597);
and U33161 (N_33161,N_31824,N_31651);
nor U33162 (N_33162,N_30141,N_31537);
xnor U33163 (N_33163,N_30024,N_31012);
nand U33164 (N_33164,N_30544,N_31162);
and U33165 (N_33165,N_31332,N_30936);
and U33166 (N_33166,N_30653,N_31086);
nand U33167 (N_33167,N_30788,N_30631);
and U33168 (N_33168,N_31822,N_31320);
nor U33169 (N_33169,N_31460,N_30973);
or U33170 (N_33170,N_30090,N_31739);
and U33171 (N_33171,N_31523,N_30209);
and U33172 (N_33172,N_30042,N_30181);
and U33173 (N_33173,N_30639,N_31114);
and U33174 (N_33174,N_30767,N_31731);
nor U33175 (N_33175,N_31199,N_31311);
xnor U33176 (N_33176,N_31906,N_31208);
or U33177 (N_33177,N_30991,N_31350);
xor U33178 (N_33178,N_30464,N_31760);
or U33179 (N_33179,N_30899,N_30675);
nor U33180 (N_33180,N_30623,N_30333);
and U33181 (N_33181,N_30714,N_31678);
xnor U33182 (N_33182,N_31004,N_31329);
nand U33183 (N_33183,N_31354,N_30298);
xor U33184 (N_33184,N_30550,N_30745);
or U33185 (N_33185,N_30352,N_31523);
nor U33186 (N_33186,N_30898,N_30760);
nor U33187 (N_33187,N_31072,N_31688);
nand U33188 (N_33188,N_30256,N_30897);
nor U33189 (N_33189,N_31095,N_30821);
and U33190 (N_33190,N_30255,N_30284);
and U33191 (N_33191,N_30749,N_31084);
nor U33192 (N_33192,N_31582,N_30675);
or U33193 (N_33193,N_31554,N_30894);
nand U33194 (N_33194,N_31186,N_31230);
or U33195 (N_33195,N_31563,N_31172);
and U33196 (N_33196,N_30934,N_31499);
and U33197 (N_33197,N_30988,N_30066);
xnor U33198 (N_33198,N_30749,N_31741);
and U33199 (N_33199,N_31989,N_30691);
and U33200 (N_33200,N_30123,N_31190);
xnor U33201 (N_33201,N_30542,N_31333);
or U33202 (N_33202,N_31582,N_30487);
nor U33203 (N_33203,N_30042,N_31192);
or U33204 (N_33204,N_31808,N_30978);
or U33205 (N_33205,N_31694,N_30647);
or U33206 (N_33206,N_31192,N_30518);
and U33207 (N_33207,N_31370,N_31313);
or U33208 (N_33208,N_30706,N_30236);
and U33209 (N_33209,N_31082,N_31198);
and U33210 (N_33210,N_30828,N_30738);
or U33211 (N_33211,N_31020,N_31205);
xor U33212 (N_33212,N_30353,N_31051);
nand U33213 (N_33213,N_30064,N_30239);
xnor U33214 (N_33214,N_31184,N_31132);
nand U33215 (N_33215,N_31799,N_30220);
and U33216 (N_33216,N_31756,N_31356);
or U33217 (N_33217,N_30417,N_30220);
and U33218 (N_33218,N_30570,N_30460);
or U33219 (N_33219,N_31465,N_30302);
and U33220 (N_33220,N_30881,N_30596);
or U33221 (N_33221,N_30865,N_31641);
and U33222 (N_33222,N_30709,N_30457);
and U33223 (N_33223,N_31679,N_30694);
or U33224 (N_33224,N_30740,N_31527);
nand U33225 (N_33225,N_30763,N_31334);
or U33226 (N_33226,N_31134,N_31953);
nor U33227 (N_33227,N_30184,N_30982);
xnor U33228 (N_33228,N_31874,N_30416);
and U33229 (N_33229,N_30099,N_31524);
and U33230 (N_33230,N_31863,N_30817);
nand U33231 (N_33231,N_31284,N_31371);
nor U33232 (N_33232,N_31750,N_30344);
or U33233 (N_33233,N_30753,N_30482);
xnor U33234 (N_33234,N_31556,N_31381);
nand U33235 (N_33235,N_31451,N_31487);
and U33236 (N_33236,N_30884,N_31039);
nand U33237 (N_33237,N_31601,N_30436);
and U33238 (N_33238,N_31190,N_31885);
nor U33239 (N_33239,N_30148,N_30269);
nor U33240 (N_33240,N_30400,N_31944);
nand U33241 (N_33241,N_30897,N_30689);
and U33242 (N_33242,N_31172,N_30043);
nor U33243 (N_33243,N_31649,N_31471);
or U33244 (N_33244,N_30802,N_30532);
nor U33245 (N_33245,N_31621,N_31828);
xnor U33246 (N_33246,N_31092,N_30417);
nor U33247 (N_33247,N_31336,N_30255);
xor U33248 (N_33248,N_31646,N_30430);
and U33249 (N_33249,N_31118,N_31148);
nand U33250 (N_33250,N_31989,N_31341);
and U33251 (N_33251,N_30631,N_30153);
xor U33252 (N_33252,N_30681,N_30655);
xnor U33253 (N_33253,N_31314,N_31484);
nor U33254 (N_33254,N_30767,N_30983);
or U33255 (N_33255,N_30965,N_31221);
and U33256 (N_33256,N_31623,N_31565);
and U33257 (N_33257,N_31296,N_30286);
nand U33258 (N_33258,N_31423,N_31515);
xnor U33259 (N_33259,N_30220,N_31355);
or U33260 (N_33260,N_31587,N_30392);
nor U33261 (N_33261,N_30200,N_31552);
xor U33262 (N_33262,N_31013,N_30910);
and U33263 (N_33263,N_31837,N_30970);
xor U33264 (N_33264,N_30111,N_30751);
or U33265 (N_33265,N_31143,N_30832);
or U33266 (N_33266,N_31220,N_31488);
xor U33267 (N_33267,N_31487,N_30961);
xor U33268 (N_33268,N_31133,N_30390);
or U33269 (N_33269,N_30447,N_31207);
and U33270 (N_33270,N_31519,N_31214);
nor U33271 (N_33271,N_30828,N_30448);
nand U33272 (N_33272,N_31929,N_30891);
nor U33273 (N_33273,N_30600,N_31446);
nor U33274 (N_33274,N_31634,N_31940);
nand U33275 (N_33275,N_31940,N_30501);
and U33276 (N_33276,N_30356,N_30450);
and U33277 (N_33277,N_30684,N_30781);
and U33278 (N_33278,N_30739,N_31325);
xnor U33279 (N_33279,N_31804,N_31340);
nand U33280 (N_33280,N_30434,N_31592);
or U33281 (N_33281,N_30667,N_31661);
nor U33282 (N_33282,N_31164,N_31671);
and U33283 (N_33283,N_31547,N_30963);
xor U33284 (N_33284,N_31754,N_31392);
xor U33285 (N_33285,N_30531,N_31907);
nor U33286 (N_33286,N_31868,N_30788);
xor U33287 (N_33287,N_31435,N_30836);
nand U33288 (N_33288,N_31851,N_31528);
xor U33289 (N_33289,N_30139,N_30304);
xor U33290 (N_33290,N_30904,N_31183);
and U33291 (N_33291,N_31323,N_31610);
or U33292 (N_33292,N_30948,N_30616);
nor U33293 (N_33293,N_30039,N_30140);
nor U33294 (N_33294,N_31553,N_30208);
xnor U33295 (N_33295,N_30388,N_30212);
nor U33296 (N_33296,N_30302,N_31067);
nor U33297 (N_33297,N_31495,N_30172);
and U33298 (N_33298,N_31328,N_31036);
or U33299 (N_33299,N_31610,N_31749);
or U33300 (N_33300,N_30001,N_31546);
xor U33301 (N_33301,N_31654,N_30034);
xnor U33302 (N_33302,N_30216,N_31641);
nor U33303 (N_33303,N_30609,N_30573);
nand U33304 (N_33304,N_31084,N_30518);
xor U33305 (N_33305,N_31927,N_30139);
and U33306 (N_33306,N_31487,N_31443);
xnor U33307 (N_33307,N_31939,N_30736);
or U33308 (N_33308,N_31420,N_30692);
xor U33309 (N_33309,N_30320,N_31047);
nand U33310 (N_33310,N_31663,N_31802);
nand U33311 (N_33311,N_31048,N_30018);
nor U33312 (N_33312,N_31643,N_30075);
and U33313 (N_33313,N_30987,N_31653);
nor U33314 (N_33314,N_31077,N_30801);
nand U33315 (N_33315,N_30396,N_31573);
nor U33316 (N_33316,N_30431,N_31594);
xnor U33317 (N_33317,N_30128,N_30342);
nand U33318 (N_33318,N_31500,N_31810);
xnor U33319 (N_33319,N_30075,N_31848);
or U33320 (N_33320,N_30983,N_30131);
or U33321 (N_33321,N_30126,N_30692);
or U33322 (N_33322,N_30090,N_30393);
nand U33323 (N_33323,N_31342,N_30955);
or U33324 (N_33324,N_31066,N_31531);
and U33325 (N_33325,N_30428,N_30880);
xor U33326 (N_33326,N_30568,N_31852);
or U33327 (N_33327,N_31623,N_31855);
or U33328 (N_33328,N_30278,N_30649);
nor U33329 (N_33329,N_30430,N_31350);
and U33330 (N_33330,N_31217,N_30296);
or U33331 (N_33331,N_30984,N_31211);
xor U33332 (N_33332,N_30456,N_30867);
xor U33333 (N_33333,N_30401,N_30369);
xor U33334 (N_33334,N_30692,N_30004);
nand U33335 (N_33335,N_30488,N_31605);
or U33336 (N_33336,N_31400,N_30923);
nand U33337 (N_33337,N_31424,N_31291);
xor U33338 (N_33338,N_30508,N_31041);
or U33339 (N_33339,N_30146,N_31567);
nand U33340 (N_33340,N_30385,N_30065);
nor U33341 (N_33341,N_31107,N_30145);
xnor U33342 (N_33342,N_30090,N_31236);
nand U33343 (N_33343,N_31522,N_30214);
or U33344 (N_33344,N_31886,N_31977);
xnor U33345 (N_33345,N_31157,N_30098);
nand U33346 (N_33346,N_30889,N_30767);
xnor U33347 (N_33347,N_30507,N_30227);
or U33348 (N_33348,N_31730,N_30259);
and U33349 (N_33349,N_31435,N_31452);
and U33350 (N_33350,N_31327,N_31932);
and U33351 (N_33351,N_30231,N_30363);
nand U33352 (N_33352,N_30114,N_31233);
nand U33353 (N_33353,N_30981,N_31119);
xnor U33354 (N_33354,N_30831,N_30364);
xnor U33355 (N_33355,N_30164,N_30252);
and U33356 (N_33356,N_31847,N_31185);
and U33357 (N_33357,N_31633,N_30144);
and U33358 (N_33358,N_30371,N_31059);
and U33359 (N_33359,N_31111,N_30932);
and U33360 (N_33360,N_31695,N_30513);
or U33361 (N_33361,N_31321,N_30235);
xnor U33362 (N_33362,N_30305,N_31046);
or U33363 (N_33363,N_31128,N_31884);
or U33364 (N_33364,N_30868,N_30043);
nand U33365 (N_33365,N_30206,N_31536);
or U33366 (N_33366,N_31457,N_31203);
nor U33367 (N_33367,N_30977,N_30881);
and U33368 (N_33368,N_30640,N_31496);
nor U33369 (N_33369,N_30724,N_30282);
and U33370 (N_33370,N_31814,N_31778);
or U33371 (N_33371,N_31401,N_30390);
nor U33372 (N_33372,N_30163,N_30575);
or U33373 (N_33373,N_31139,N_30893);
nand U33374 (N_33374,N_31335,N_30652);
nand U33375 (N_33375,N_31846,N_31356);
and U33376 (N_33376,N_30847,N_31269);
nand U33377 (N_33377,N_30021,N_30885);
nor U33378 (N_33378,N_30519,N_31806);
nand U33379 (N_33379,N_30010,N_31658);
and U33380 (N_33380,N_30698,N_31977);
xor U33381 (N_33381,N_30506,N_30999);
nor U33382 (N_33382,N_31753,N_31285);
nor U33383 (N_33383,N_30263,N_30064);
nor U33384 (N_33384,N_30918,N_31410);
nor U33385 (N_33385,N_31949,N_31317);
xnor U33386 (N_33386,N_31594,N_31063);
or U33387 (N_33387,N_31871,N_31694);
and U33388 (N_33388,N_30491,N_30339);
nor U33389 (N_33389,N_30824,N_31441);
or U33390 (N_33390,N_31873,N_30589);
nor U33391 (N_33391,N_31013,N_30760);
or U33392 (N_33392,N_30066,N_30408);
or U33393 (N_33393,N_31475,N_31321);
nor U33394 (N_33394,N_31614,N_31322);
or U33395 (N_33395,N_30033,N_30464);
nand U33396 (N_33396,N_30756,N_30837);
xnor U33397 (N_33397,N_31172,N_31072);
nor U33398 (N_33398,N_31238,N_30199);
nor U33399 (N_33399,N_31636,N_30632);
nand U33400 (N_33400,N_30081,N_30637);
nor U33401 (N_33401,N_31495,N_30858);
nand U33402 (N_33402,N_30682,N_30502);
xor U33403 (N_33403,N_31861,N_30382);
nor U33404 (N_33404,N_30604,N_30780);
or U33405 (N_33405,N_31057,N_31965);
nor U33406 (N_33406,N_30962,N_31979);
and U33407 (N_33407,N_31821,N_31371);
or U33408 (N_33408,N_31097,N_30177);
or U33409 (N_33409,N_30025,N_31697);
and U33410 (N_33410,N_31551,N_31154);
nor U33411 (N_33411,N_31907,N_30478);
xnor U33412 (N_33412,N_30146,N_30936);
or U33413 (N_33413,N_31028,N_30849);
and U33414 (N_33414,N_31729,N_30919);
or U33415 (N_33415,N_30949,N_30047);
nor U33416 (N_33416,N_30970,N_30696);
or U33417 (N_33417,N_31246,N_31148);
or U33418 (N_33418,N_31931,N_30881);
nor U33419 (N_33419,N_30812,N_30236);
and U33420 (N_33420,N_31066,N_31465);
and U33421 (N_33421,N_31741,N_31819);
and U33422 (N_33422,N_31229,N_31963);
and U33423 (N_33423,N_30057,N_30235);
and U33424 (N_33424,N_30264,N_31430);
nand U33425 (N_33425,N_31497,N_30582);
nor U33426 (N_33426,N_31750,N_31941);
nand U33427 (N_33427,N_31278,N_31997);
or U33428 (N_33428,N_30624,N_30630);
xor U33429 (N_33429,N_30747,N_31384);
and U33430 (N_33430,N_31470,N_31660);
xor U33431 (N_33431,N_30409,N_31725);
nor U33432 (N_33432,N_30271,N_30031);
and U33433 (N_33433,N_30522,N_30282);
or U33434 (N_33434,N_30232,N_31456);
and U33435 (N_33435,N_31142,N_31435);
and U33436 (N_33436,N_31537,N_31588);
or U33437 (N_33437,N_31714,N_31374);
nand U33438 (N_33438,N_30680,N_30600);
nor U33439 (N_33439,N_31016,N_30465);
nand U33440 (N_33440,N_30025,N_30987);
nand U33441 (N_33441,N_30186,N_30195);
xnor U33442 (N_33442,N_31508,N_30125);
xnor U33443 (N_33443,N_31676,N_31413);
xnor U33444 (N_33444,N_30999,N_31520);
or U33445 (N_33445,N_30529,N_31277);
nand U33446 (N_33446,N_30956,N_30301);
or U33447 (N_33447,N_31216,N_30607);
xor U33448 (N_33448,N_31347,N_31645);
and U33449 (N_33449,N_30412,N_30957);
and U33450 (N_33450,N_30155,N_30396);
or U33451 (N_33451,N_31297,N_31924);
or U33452 (N_33452,N_30519,N_31456);
and U33453 (N_33453,N_30780,N_31276);
nor U33454 (N_33454,N_31052,N_30503);
and U33455 (N_33455,N_31598,N_30625);
nor U33456 (N_33456,N_30128,N_31399);
or U33457 (N_33457,N_31359,N_30187);
nand U33458 (N_33458,N_31898,N_31354);
nand U33459 (N_33459,N_30443,N_31214);
nand U33460 (N_33460,N_31739,N_31927);
nor U33461 (N_33461,N_31319,N_31441);
or U33462 (N_33462,N_31026,N_31515);
nand U33463 (N_33463,N_31549,N_31679);
or U33464 (N_33464,N_31594,N_30495);
nor U33465 (N_33465,N_30491,N_30157);
nor U33466 (N_33466,N_31146,N_31766);
nand U33467 (N_33467,N_30901,N_30883);
or U33468 (N_33468,N_31208,N_30087);
nor U33469 (N_33469,N_31588,N_31595);
or U33470 (N_33470,N_31378,N_31143);
xnor U33471 (N_33471,N_30585,N_30640);
and U33472 (N_33472,N_31919,N_31397);
nand U33473 (N_33473,N_31329,N_30991);
and U33474 (N_33474,N_31838,N_31385);
nor U33475 (N_33475,N_31405,N_31514);
nor U33476 (N_33476,N_30064,N_30146);
nand U33477 (N_33477,N_30884,N_30106);
or U33478 (N_33478,N_31012,N_31596);
xor U33479 (N_33479,N_30578,N_31722);
nand U33480 (N_33480,N_31088,N_30721);
or U33481 (N_33481,N_31354,N_30213);
or U33482 (N_33482,N_30720,N_30641);
xnor U33483 (N_33483,N_30034,N_30065);
nor U33484 (N_33484,N_30954,N_31429);
and U33485 (N_33485,N_31431,N_30960);
or U33486 (N_33486,N_30841,N_31454);
nor U33487 (N_33487,N_30539,N_31093);
nor U33488 (N_33488,N_31300,N_30978);
xor U33489 (N_33489,N_30957,N_31314);
and U33490 (N_33490,N_31180,N_31225);
and U33491 (N_33491,N_30967,N_30127);
nand U33492 (N_33492,N_30620,N_30313);
and U33493 (N_33493,N_30393,N_30890);
or U33494 (N_33494,N_31272,N_30965);
and U33495 (N_33495,N_30619,N_30577);
nand U33496 (N_33496,N_30786,N_31094);
and U33497 (N_33497,N_30238,N_31264);
and U33498 (N_33498,N_30397,N_31401);
and U33499 (N_33499,N_30526,N_31466);
nand U33500 (N_33500,N_31111,N_31358);
and U33501 (N_33501,N_30472,N_30759);
nand U33502 (N_33502,N_30591,N_30317);
and U33503 (N_33503,N_31724,N_31867);
xor U33504 (N_33504,N_30114,N_30939);
xor U33505 (N_33505,N_31284,N_30405);
nand U33506 (N_33506,N_31549,N_30751);
xnor U33507 (N_33507,N_31987,N_30333);
and U33508 (N_33508,N_30819,N_31479);
and U33509 (N_33509,N_30774,N_30175);
nand U33510 (N_33510,N_30297,N_31193);
and U33511 (N_33511,N_31101,N_30017);
xor U33512 (N_33512,N_30029,N_31715);
or U33513 (N_33513,N_31695,N_30790);
or U33514 (N_33514,N_30290,N_31145);
xor U33515 (N_33515,N_31909,N_31279);
and U33516 (N_33516,N_30493,N_30234);
nor U33517 (N_33517,N_30003,N_31290);
and U33518 (N_33518,N_31018,N_31466);
nor U33519 (N_33519,N_30407,N_30090);
nand U33520 (N_33520,N_30987,N_30281);
xnor U33521 (N_33521,N_30897,N_31052);
and U33522 (N_33522,N_30871,N_30213);
xnor U33523 (N_33523,N_31194,N_31916);
nor U33524 (N_33524,N_30506,N_31109);
and U33525 (N_33525,N_31166,N_31098);
or U33526 (N_33526,N_31637,N_31461);
xnor U33527 (N_33527,N_30236,N_30783);
xnor U33528 (N_33528,N_31348,N_31093);
or U33529 (N_33529,N_31413,N_30835);
xnor U33530 (N_33530,N_31892,N_31035);
xnor U33531 (N_33531,N_30147,N_30946);
and U33532 (N_33532,N_31601,N_30421);
or U33533 (N_33533,N_30629,N_31290);
and U33534 (N_33534,N_30859,N_30099);
and U33535 (N_33535,N_31702,N_31296);
and U33536 (N_33536,N_30876,N_31577);
and U33537 (N_33537,N_31389,N_31298);
nand U33538 (N_33538,N_30254,N_31585);
and U33539 (N_33539,N_30098,N_31078);
nand U33540 (N_33540,N_31461,N_31256);
or U33541 (N_33541,N_31520,N_30195);
nand U33542 (N_33542,N_30274,N_30621);
and U33543 (N_33543,N_30565,N_31502);
xnor U33544 (N_33544,N_31733,N_31380);
xnor U33545 (N_33545,N_31969,N_31962);
nor U33546 (N_33546,N_30190,N_31549);
nor U33547 (N_33547,N_30246,N_30676);
or U33548 (N_33548,N_31081,N_30188);
nor U33549 (N_33549,N_31527,N_31408);
nand U33550 (N_33550,N_30272,N_31001);
nand U33551 (N_33551,N_30753,N_31073);
and U33552 (N_33552,N_31812,N_30812);
xnor U33553 (N_33553,N_30928,N_31681);
nor U33554 (N_33554,N_31696,N_30126);
xor U33555 (N_33555,N_31265,N_31770);
nand U33556 (N_33556,N_31704,N_31762);
nor U33557 (N_33557,N_30978,N_30341);
nand U33558 (N_33558,N_31802,N_31863);
xor U33559 (N_33559,N_30470,N_30710);
nor U33560 (N_33560,N_30021,N_31112);
nor U33561 (N_33561,N_30038,N_30705);
or U33562 (N_33562,N_30582,N_31035);
or U33563 (N_33563,N_30584,N_31661);
xor U33564 (N_33564,N_30040,N_30235);
nand U33565 (N_33565,N_30668,N_31669);
nor U33566 (N_33566,N_31001,N_31548);
nand U33567 (N_33567,N_30876,N_31354);
or U33568 (N_33568,N_30265,N_30322);
nor U33569 (N_33569,N_30014,N_31881);
xor U33570 (N_33570,N_31903,N_31774);
or U33571 (N_33571,N_31443,N_31011);
or U33572 (N_33572,N_31498,N_31983);
xnor U33573 (N_33573,N_30256,N_31406);
nand U33574 (N_33574,N_31942,N_30877);
nor U33575 (N_33575,N_30174,N_31333);
nand U33576 (N_33576,N_31931,N_30308);
or U33577 (N_33577,N_31959,N_30566);
nand U33578 (N_33578,N_31980,N_30092);
or U33579 (N_33579,N_30233,N_30556);
nand U33580 (N_33580,N_30801,N_31739);
nand U33581 (N_33581,N_31186,N_30608);
nand U33582 (N_33582,N_31411,N_30270);
nand U33583 (N_33583,N_30399,N_31402);
nor U33584 (N_33584,N_31981,N_30698);
nor U33585 (N_33585,N_31915,N_31129);
and U33586 (N_33586,N_30276,N_31410);
or U33587 (N_33587,N_31021,N_30736);
xor U33588 (N_33588,N_31931,N_30557);
nor U33589 (N_33589,N_31469,N_31711);
nand U33590 (N_33590,N_31681,N_30268);
and U33591 (N_33591,N_30858,N_30416);
nand U33592 (N_33592,N_30395,N_30558);
nor U33593 (N_33593,N_31223,N_31080);
nor U33594 (N_33594,N_30492,N_31188);
xnor U33595 (N_33595,N_31927,N_31769);
and U33596 (N_33596,N_31994,N_31786);
and U33597 (N_33597,N_30010,N_31292);
nand U33598 (N_33598,N_31604,N_31771);
and U33599 (N_33599,N_30571,N_30486);
and U33600 (N_33600,N_30881,N_31732);
nor U33601 (N_33601,N_30569,N_31139);
or U33602 (N_33602,N_30581,N_31790);
xnor U33603 (N_33603,N_30536,N_30709);
nor U33604 (N_33604,N_31558,N_30228);
nand U33605 (N_33605,N_30162,N_31137);
or U33606 (N_33606,N_30132,N_31482);
nor U33607 (N_33607,N_30332,N_30875);
and U33608 (N_33608,N_30842,N_30779);
and U33609 (N_33609,N_30615,N_31200);
nor U33610 (N_33610,N_31492,N_30913);
xnor U33611 (N_33611,N_31947,N_30804);
nor U33612 (N_33612,N_31155,N_30341);
or U33613 (N_33613,N_31359,N_30689);
and U33614 (N_33614,N_31556,N_31724);
and U33615 (N_33615,N_30137,N_31362);
xor U33616 (N_33616,N_30335,N_31487);
xor U33617 (N_33617,N_30933,N_30883);
nand U33618 (N_33618,N_30663,N_30089);
nand U33619 (N_33619,N_30491,N_31147);
and U33620 (N_33620,N_30779,N_31186);
or U33621 (N_33621,N_30925,N_31542);
nor U33622 (N_33622,N_30852,N_30778);
xor U33623 (N_33623,N_31359,N_30226);
nand U33624 (N_33624,N_30600,N_30551);
nor U33625 (N_33625,N_30881,N_31877);
nor U33626 (N_33626,N_30440,N_31885);
or U33627 (N_33627,N_31751,N_31327);
and U33628 (N_33628,N_30516,N_30936);
xnor U33629 (N_33629,N_30334,N_31082);
xnor U33630 (N_33630,N_30207,N_30042);
or U33631 (N_33631,N_30730,N_31456);
nor U33632 (N_33632,N_30165,N_30166);
nor U33633 (N_33633,N_31068,N_30188);
or U33634 (N_33634,N_30281,N_30881);
and U33635 (N_33635,N_30398,N_31596);
or U33636 (N_33636,N_30805,N_30019);
and U33637 (N_33637,N_31678,N_30521);
or U33638 (N_33638,N_30909,N_30654);
nand U33639 (N_33639,N_31759,N_31625);
and U33640 (N_33640,N_30207,N_31617);
nand U33641 (N_33641,N_30275,N_31145);
or U33642 (N_33642,N_30501,N_30999);
nand U33643 (N_33643,N_30508,N_30790);
xnor U33644 (N_33644,N_31916,N_31460);
nand U33645 (N_33645,N_31862,N_31855);
or U33646 (N_33646,N_30279,N_31663);
xnor U33647 (N_33647,N_31554,N_31897);
nor U33648 (N_33648,N_30000,N_30067);
and U33649 (N_33649,N_30027,N_30635);
or U33650 (N_33650,N_30577,N_31520);
and U33651 (N_33651,N_30230,N_31092);
nor U33652 (N_33652,N_30997,N_31981);
xnor U33653 (N_33653,N_31671,N_31749);
xnor U33654 (N_33654,N_30036,N_31788);
or U33655 (N_33655,N_30243,N_31711);
or U33656 (N_33656,N_30268,N_31279);
or U33657 (N_33657,N_30881,N_31986);
or U33658 (N_33658,N_31993,N_31797);
nand U33659 (N_33659,N_31387,N_30738);
nor U33660 (N_33660,N_31351,N_30145);
xor U33661 (N_33661,N_30099,N_31804);
nand U33662 (N_33662,N_31612,N_30440);
nor U33663 (N_33663,N_31849,N_31666);
and U33664 (N_33664,N_30293,N_30629);
nand U33665 (N_33665,N_31607,N_30888);
xnor U33666 (N_33666,N_31139,N_31525);
xor U33667 (N_33667,N_30554,N_31980);
xor U33668 (N_33668,N_31217,N_30301);
and U33669 (N_33669,N_30388,N_31745);
or U33670 (N_33670,N_30001,N_31852);
or U33671 (N_33671,N_30756,N_30019);
xnor U33672 (N_33672,N_30866,N_30776);
nand U33673 (N_33673,N_31993,N_30230);
xor U33674 (N_33674,N_30655,N_31744);
nand U33675 (N_33675,N_30423,N_30649);
nand U33676 (N_33676,N_31248,N_31165);
or U33677 (N_33677,N_30542,N_31049);
nor U33678 (N_33678,N_30996,N_31638);
nor U33679 (N_33679,N_31617,N_30793);
nand U33680 (N_33680,N_31464,N_31407);
and U33681 (N_33681,N_31879,N_31657);
nand U33682 (N_33682,N_31009,N_30529);
xor U33683 (N_33683,N_31059,N_30574);
nand U33684 (N_33684,N_30172,N_30134);
xor U33685 (N_33685,N_30748,N_31420);
nand U33686 (N_33686,N_31586,N_31914);
and U33687 (N_33687,N_30141,N_31033);
and U33688 (N_33688,N_31309,N_31184);
nor U33689 (N_33689,N_30830,N_30574);
nand U33690 (N_33690,N_31485,N_31093);
xnor U33691 (N_33691,N_31552,N_30666);
nand U33692 (N_33692,N_31345,N_30371);
nand U33693 (N_33693,N_31397,N_30661);
xor U33694 (N_33694,N_30561,N_31836);
or U33695 (N_33695,N_31561,N_30544);
nand U33696 (N_33696,N_30023,N_30137);
or U33697 (N_33697,N_31950,N_31162);
nor U33698 (N_33698,N_30645,N_31019);
and U33699 (N_33699,N_30739,N_31029);
xnor U33700 (N_33700,N_31905,N_30517);
and U33701 (N_33701,N_31886,N_30442);
xor U33702 (N_33702,N_30566,N_31932);
xor U33703 (N_33703,N_30862,N_30604);
or U33704 (N_33704,N_30016,N_31026);
and U33705 (N_33705,N_30822,N_30567);
xor U33706 (N_33706,N_31487,N_31071);
nand U33707 (N_33707,N_30491,N_30478);
or U33708 (N_33708,N_31937,N_30377);
nor U33709 (N_33709,N_31014,N_30089);
nor U33710 (N_33710,N_30375,N_30005);
nand U33711 (N_33711,N_30813,N_30364);
xnor U33712 (N_33712,N_30420,N_31772);
nor U33713 (N_33713,N_31712,N_30601);
and U33714 (N_33714,N_30670,N_30843);
or U33715 (N_33715,N_30803,N_30000);
xnor U33716 (N_33716,N_30854,N_30711);
xor U33717 (N_33717,N_30697,N_30315);
nor U33718 (N_33718,N_30227,N_30799);
and U33719 (N_33719,N_30811,N_31225);
nor U33720 (N_33720,N_31385,N_30693);
or U33721 (N_33721,N_31255,N_30663);
nand U33722 (N_33722,N_31191,N_31918);
xor U33723 (N_33723,N_31847,N_31557);
or U33724 (N_33724,N_31252,N_31354);
and U33725 (N_33725,N_31294,N_30391);
xor U33726 (N_33726,N_31203,N_31100);
or U33727 (N_33727,N_31032,N_31211);
nand U33728 (N_33728,N_31175,N_30828);
and U33729 (N_33729,N_30992,N_31299);
and U33730 (N_33730,N_30020,N_30975);
nand U33731 (N_33731,N_30418,N_30095);
xnor U33732 (N_33732,N_30256,N_30120);
or U33733 (N_33733,N_31388,N_30911);
nor U33734 (N_33734,N_31376,N_31832);
xor U33735 (N_33735,N_30314,N_31377);
or U33736 (N_33736,N_30928,N_31905);
xor U33737 (N_33737,N_30663,N_31415);
xor U33738 (N_33738,N_31172,N_31711);
or U33739 (N_33739,N_30355,N_30360);
nor U33740 (N_33740,N_30951,N_31313);
and U33741 (N_33741,N_31397,N_30138);
nand U33742 (N_33742,N_31966,N_31317);
xnor U33743 (N_33743,N_30689,N_30418);
or U33744 (N_33744,N_31686,N_30625);
and U33745 (N_33745,N_30367,N_31296);
and U33746 (N_33746,N_31034,N_30604);
and U33747 (N_33747,N_30989,N_31147);
nand U33748 (N_33748,N_30747,N_31932);
or U33749 (N_33749,N_31564,N_31323);
nand U33750 (N_33750,N_31509,N_30089);
nand U33751 (N_33751,N_30564,N_30195);
xor U33752 (N_33752,N_31903,N_30143);
and U33753 (N_33753,N_31896,N_31541);
nor U33754 (N_33754,N_31021,N_30614);
or U33755 (N_33755,N_31820,N_31117);
and U33756 (N_33756,N_30367,N_30831);
and U33757 (N_33757,N_30916,N_30103);
nand U33758 (N_33758,N_31875,N_30595);
and U33759 (N_33759,N_31326,N_31294);
or U33760 (N_33760,N_31061,N_31999);
nor U33761 (N_33761,N_30612,N_30466);
and U33762 (N_33762,N_30681,N_30627);
xor U33763 (N_33763,N_31759,N_30145);
xor U33764 (N_33764,N_30851,N_31497);
xor U33765 (N_33765,N_31926,N_30177);
or U33766 (N_33766,N_31390,N_30681);
nand U33767 (N_33767,N_31671,N_30655);
nand U33768 (N_33768,N_31392,N_31855);
nor U33769 (N_33769,N_31343,N_31841);
and U33770 (N_33770,N_31936,N_30611);
xnor U33771 (N_33771,N_31947,N_30674);
nand U33772 (N_33772,N_30431,N_31593);
xor U33773 (N_33773,N_31093,N_31692);
xor U33774 (N_33774,N_30402,N_31451);
and U33775 (N_33775,N_31464,N_30822);
xor U33776 (N_33776,N_31966,N_31472);
nand U33777 (N_33777,N_30075,N_30929);
and U33778 (N_33778,N_30201,N_30312);
nor U33779 (N_33779,N_31331,N_31694);
nand U33780 (N_33780,N_31837,N_31265);
xor U33781 (N_33781,N_30017,N_31366);
nand U33782 (N_33782,N_31439,N_31748);
nor U33783 (N_33783,N_30849,N_30347);
nor U33784 (N_33784,N_30191,N_31511);
nand U33785 (N_33785,N_31350,N_31677);
nand U33786 (N_33786,N_30513,N_30907);
nand U33787 (N_33787,N_31338,N_31214);
and U33788 (N_33788,N_30507,N_30312);
nor U33789 (N_33789,N_31080,N_30773);
or U33790 (N_33790,N_31167,N_31757);
xnor U33791 (N_33791,N_31083,N_31979);
nor U33792 (N_33792,N_31660,N_30820);
nand U33793 (N_33793,N_30699,N_31681);
or U33794 (N_33794,N_31335,N_31127);
nor U33795 (N_33795,N_30195,N_31845);
nor U33796 (N_33796,N_31751,N_30460);
nor U33797 (N_33797,N_31902,N_31662);
or U33798 (N_33798,N_30478,N_31511);
nand U33799 (N_33799,N_31399,N_31132);
xor U33800 (N_33800,N_31593,N_30230);
and U33801 (N_33801,N_30950,N_31445);
or U33802 (N_33802,N_31838,N_31257);
nor U33803 (N_33803,N_30247,N_31072);
nor U33804 (N_33804,N_31367,N_30687);
nand U33805 (N_33805,N_31035,N_31847);
nand U33806 (N_33806,N_31650,N_30795);
and U33807 (N_33807,N_31646,N_30678);
nor U33808 (N_33808,N_30253,N_30681);
or U33809 (N_33809,N_30058,N_31709);
xor U33810 (N_33810,N_30818,N_30063);
xnor U33811 (N_33811,N_31227,N_31585);
and U33812 (N_33812,N_30832,N_30465);
or U33813 (N_33813,N_30434,N_31898);
or U33814 (N_33814,N_31725,N_31074);
and U33815 (N_33815,N_30744,N_31919);
xnor U33816 (N_33816,N_31301,N_30366);
or U33817 (N_33817,N_31476,N_31498);
nand U33818 (N_33818,N_31507,N_30922);
nor U33819 (N_33819,N_30476,N_30670);
or U33820 (N_33820,N_30082,N_30074);
and U33821 (N_33821,N_31574,N_30269);
xnor U33822 (N_33822,N_31127,N_30675);
nand U33823 (N_33823,N_31533,N_30091);
nor U33824 (N_33824,N_30472,N_30336);
and U33825 (N_33825,N_30081,N_30190);
or U33826 (N_33826,N_30889,N_30945);
nor U33827 (N_33827,N_30453,N_30350);
nor U33828 (N_33828,N_30229,N_30615);
nand U33829 (N_33829,N_30249,N_31758);
nand U33830 (N_33830,N_31688,N_30473);
xnor U33831 (N_33831,N_31228,N_30356);
or U33832 (N_33832,N_31931,N_30023);
xor U33833 (N_33833,N_31042,N_31418);
and U33834 (N_33834,N_31256,N_30624);
xnor U33835 (N_33835,N_30583,N_30331);
or U33836 (N_33836,N_30430,N_30822);
nand U33837 (N_33837,N_30710,N_31776);
and U33838 (N_33838,N_30123,N_30896);
nand U33839 (N_33839,N_30657,N_30440);
or U33840 (N_33840,N_30313,N_30843);
and U33841 (N_33841,N_31896,N_30904);
xnor U33842 (N_33842,N_31862,N_30435);
nor U33843 (N_33843,N_31704,N_30835);
nand U33844 (N_33844,N_30110,N_31586);
xor U33845 (N_33845,N_30811,N_30892);
xnor U33846 (N_33846,N_30898,N_31953);
and U33847 (N_33847,N_31267,N_30247);
nor U33848 (N_33848,N_30683,N_31618);
nand U33849 (N_33849,N_30094,N_31713);
or U33850 (N_33850,N_31153,N_31071);
and U33851 (N_33851,N_30167,N_30745);
nor U33852 (N_33852,N_31328,N_30732);
and U33853 (N_33853,N_30077,N_30550);
nand U33854 (N_33854,N_31804,N_30074);
and U33855 (N_33855,N_31003,N_31707);
nand U33856 (N_33856,N_31958,N_30580);
nor U33857 (N_33857,N_30620,N_31793);
nor U33858 (N_33858,N_31973,N_31169);
nor U33859 (N_33859,N_31338,N_31053);
nor U33860 (N_33860,N_30380,N_31896);
nand U33861 (N_33861,N_31304,N_31263);
xor U33862 (N_33862,N_31681,N_30470);
nor U33863 (N_33863,N_30765,N_30146);
and U33864 (N_33864,N_31449,N_31053);
or U33865 (N_33865,N_30216,N_30675);
xor U33866 (N_33866,N_31390,N_30300);
nor U33867 (N_33867,N_30315,N_30999);
nand U33868 (N_33868,N_31628,N_30825);
nor U33869 (N_33869,N_31708,N_30071);
or U33870 (N_33870,N_31776,N_31187);
and U33871 (N_33871,N_31656,N_30434);
or U33872 (N_33872,N_31375,N_30722);
and U33873 (N_33873,N_30702,N_30336);
or U33874 (N_33874,N_30266,N_31561);
nor U33875 (N_33875,N_31752,N_30927);
nor U33876 (N_33876,N_31981,N_31277);
nor U33877 (N_33877,N_30813,N_31489);
nand U33878 (N_33878,N_31322,N_31569);
or U33879 (N_33879,N_31141,N_30576);
nor U33880 (N_33880,N_30274,N_31108);
and U33881 (N_33881,N_30710,N_30353);
nand U33882 (N_33882,N_31249,N_30569);
xnor U33883 (N_33883,N_30771,N_30039);
or U33884 (N_33884,N_30169,N_30456);
or U33885 (N_33885,N_30648,N_30919);
or U33886 (N_33886,N_30968,N_31764);
nand U33887 (N_33887,N_31874,N_30127);
and U33888 (N_33888,N_30437,N_30807);
xor U33889 (N_33889,N_30253,N_31721);
xnor U33890 (N_33890,N_31375,N_30175);
xor U33891 (N_33891,N_31113,N_31432);
nor U33892 (N_33892,N_31373,N_30288);
nor U33893 (N_33893,N_30279,N_31564);
nand U33894 (N_33894,N_30132,N_30926);
and U33895 (N_33895,N_30267,N_30659);
nand U33896 (N_33896,N_31935,N_31368);
or U33897 (N_33897,N_31192,N_30492);
xor U33898 (N_33898,N_30810,N_30357);
nand U33899 (N_33899,N_31125,N_31231);
and U33900 (N_33900,N_30824,N_30490);
xor U33901 (N_33901,N_30565,N_30943);
or U33902 (N_33902,N_31584,N_30585);
xnor U33903 (N_33903,N_31785,N_31988);
nand U33904 (N_33904,N_31709,N_30294);
xnor U33905 (N_33905,N_31176,N_30601);
or U33906 (N_33906,N_31110,N_30671);
nor U33907 (N_33907,N_31473,N_31582);
xor U33908 (N_33908,N_30774,N_30043);
and U33909 (N_33909,N_31764,N_31118);
nand U33910 (N_33910,N_30959,N_31760);
nand U33911 (N_33911,N_31388,N_30449);
or U33912 (N_33912,N_30797,N_30665);
nor U33913 (N_33913,N_31035,N_30472);
and U33914 (N_33914,N_30251,N_31733);
nor U33915 (N_33915,N_30364,N_31690);
or U33916 (N_33916,N_30412,N_30787);
or U33917 (N_33917,N_31385,N_31225);
nand U33918 (N_33918,N_31013,N_31579);
nand U33919 (N_33919,N_30761,N_31455);
nor U33920 (N_33920,N_31702,N_31184);
and U33921 (N_33921,N_31757,N_31788);
and U33922 (N_33922,N_31773,N_30552);
xor U33923 (N_33923,N_30658,N_30500);
nor U33924 (N_33924,N_31749,N_30722);
and U33925 (N_33925,N_31761,N_31878);
or U33926 (N_33926,N_30355,N_31017);
and U33927 (N_33927,N_31651,N_30611);
nand U33928 (N_33928,N_31771,N_31683);
xor U33929 (N_33929,N_30618,N_31485);
nor U33930 (N_33930,N_31790,N_31411);
or U33931 (N_33931,N_30787,N_31988);
nand U33932 (N_33932,N_31571,N_31427);
nor U33933 (N_33933,N_31688,N_30144);
nor U33934 (N_33934,N_31110,N_31649);
nand U33935 (N_33935,N_30400,N_31836);
nand U33936 (N_33936,N_30004,N_30966);
or U33937 (N_33937,N_30227,N_30989);
nor U33938 (N_33938,N_30821,N_30748);
nand U33939 (N_33939,N_30149,N_30246);
nor U33940 (N_33940,N_31279,N_31738);
nor U33941 (N_33941,N_31420,N_31819);
nor U33942 (N_33942,N_30225,N_31880);
nor U33943 (N_33943,N_30318,N_31413);
or U33944 (N_33944,N_31585,N_31484);
and U33945 (N_33945,N_31813,N_31244);
nand U33946 (N_33946,N_30395,N_31932);
xnor U33947 (N_33947,N_31560,N_31991);
or U33948 (N_33948,N_31029,N_30795);
nor U33949 (N_33949,N_30858,N_30404);
nor U33950 (N_33950,N_30617,N_30139);
or U33951 (N_33951,N_30371,N_31151);
and U33952 (N_33952,N_30149,N_31506);
nand U33953 (N_33953,N_30820,N_31407);
nand U33954 (N_33954,N_30378,N_30756);
nand U33955 (N_33955,N_31423,N_31960);
or U33956 (N_33956,N_31068,N_31366);
and U33957 (N_33957,N_30234,N_30045);
nor U33958 (N_33958,N_31913,N_30847);
xnor U33959 (N_33959,N_30583,N_31212);
and U33960 (N_33960,N_30035,N_31860);
nand U33961 (N_33961,N_30084,N_30790);
nand U33962 (N_33962,N_31820,N_31889);
xor U33963 (N_33963,N_30884,N_31703);
xnor U33964 (N_33964,N_30689,N_31281);
and U33965 (N_33965,N_30319,N_30827);
xor U33966 (N_33966,N_30881,N_31025);
nor U33967 (N_33967,N_31451,N_30567);
nand U33968 (N_33968,N_30084,N_31415);
or U33969 (N_33969,N_30803,N_31773);
nand U33970 (N_33970,N_31214,N_31384);
xor U33971 (N_33971,N_30003,N_31835);
or U33972 (N_33972,N_31969,N_31952);
xor U33973 (N_33973,N_30096,N_31908);
nor U33974 (N_33974,N_30067,N_31775);
or U33975 (N_33975,N_30839,N_31671);
nand U33976 (N_33976,N_31268,N_31077);
nand U33977 (N_33977,N_30022,N_31156);
xnor U33978 (N_33978,N_30714,N_31216);
or U33979 (N_33979,N_31894,N_30210);
and U33980 (N_33980,N_30548,N_31971);
and U33981 (N_33981,N_31146,N_31060);
or U33982 (N_33982,N_31226,N_31477);
nand U33983 (N_33983,N_30661,N_31308);
and U33984 (N_33984,N_30852,N_30441);
nor U33985 (N_33985,N_30271,N_31847);
nor U33986 (N_33986,N_31642,N_30737);
nand U33987 (N_33987,N_30498,N_31379);
nor U33988 (N_33988,N_30784,N_30204);
and U33989 (N_33989,N_30509,N_30443);
and U33990 (N_33990,N_31464,N_30047);
xor U33991 (N_33991,N_31771,N_30974);
nand U33992 (N_33992,N_31057,N_30138);
xnor U33993 (N_33993,N_31348,N_31153);
nand U33994 (N_33994,N_31364,N_31314);
or U33995 (N_33995,N_30953,N_30795);
nand U33996 (N_33996,N_30289,N_30294);
nor U33997 (N_33997,N_30872,N_30374);
and U33998 (N_33998,N_30614,N_31210);
nor U33999 (N_33999,N_31012,N_30013);
nand U34000 (N_34000,N_32356,N_33958);
nand U34001 (N_34001,N_32607,N_32447);
and U34002 (N_34002,N_32796,N_32702);
nand U34003 (N_34003,N_33813,N_32912);
and U34004 (N_34004,N_33763,N_32347);
and U34005 (N_34005,N_32267,N_32830);
nand U34006 (N_34006,N_32513,N_32493);
or U34007 (N_34007,N_32373,N_33653);
xor U34008 (N_34008,N_32235,N_33745);
or U34009 (N_34009,N_33833,N_33038);
and U34010 (N_34010,N_33872,N_32247);
or U34011 (N_34011,N_33969,N_33750);
xor U34012 (N_34012,N_33448,N_33214);
or U34013 (N_34013,N_32305,N_32108);
xnor U34014 (N_34014,N_32670,N_33353);
or U34015 (N_34015,N_32226,N_33447);
or U34016 (N_34016,N_33183,N_33823);
or U34017 (N_34017,N_33385,N_33485);
and U34018 (N_34018,N_33998,N_33379);
or U34019 (N_34019,N_33061,N_33382);
and U34020 (N_34020,N_33370,N_33034);
and U34021 (N_34021,N_32189,N_33595);
nor U34022 (N_34022,N_33192,N_32540);
nand U34023 (N_34023,N_33285,N_33155);
xnor U34024 (N_34024,N_32681,N_32041);
nand U34025 (N_34025,N_32823,N_32369);
nor U34026 (N_34026,N_32906,N_32875);
nand U34027 (N_34027,N_33014,N_33083);
and U34028 (N_34028,N_33340,N_33298);
nand U34029 (N_34029,N_32421,N_32606);
or U34030 (N_34030,N_32709,N_32654);
nor U34031 (N_34031,N_33310,N_32029);
nor U34032 (N_34032,N_32116,N_33035);
or U34033 (N_34033,N_33159,N_33466);
or U34034 (N_34034,N_33737,N_32904);
and U34035 (N_34035,N_33207,N_33578);
or U34036 (N_34036,N_33198,N_33897);
and U34037 (N_34037,N_32896,N_32802);
and U34038 (N_34038,N_32468,N_33074);
xnor U34039 (N_34039,N_32067,N_32657);
or U34040 (N_34040,N_32626,N_33131);
and U34041 (N_34041,N_33363,N_32095);
nor U34042 (N_34042,N_33108,N_32053);
xor U34043 (N_34043,N_32722,N_33654);
nor U34044 (N_34044,N_32455,N_32159);
nor U34045 (N_34045,N_32308,N_32649);
and U34046 (N_34046,N_33919,N_33966);
and U34047 (N_34047,N_32523,N_33455);
and U34048 (N_34048,N_33105,N_32564);
nand U34049 (N_34049,N_33381,N_33586);
nor U34050 (N_34050,N_33484,N_32557);
and U34051 (N_34051,N_33293,N_32725);
nand U34052 (N_34052,N_33650,N_32089);
or U34053 (N_34053,N_32525,N_33140);
nor U34054 (N_34054,N_32700,N_32418);
and U34055 (N_34055,N_33180,N_32056);
or U34056 (N_34056,N_32266,N_33994);
or U34057 (N_34057,N_32218,N_32847);
xnor U34058 (N_34058,N_32798,N_33028);
nor U34059 (N_34059,N_32175,N_32771);
xnor U34060 (N_34060,N_33608,N_32080);
xnor U34061 (N_34061,N_33288,N_32931);
nor U34062 (N_34062,N_33817,N_33716);
or U34063 (N_34063,N_33304,N_33200);
nand U34064 (N_34064,N_32664,N_32027);
and U34065 (N_34065,N_32742,N_33889);
nand U34066 (N_34066,N_32715,N_33844);
xnor U34067 (N_34067,N_33011,N_33594);
nor U34068 (N_34068,N_32495,N_32737);
or U34069 (N_34069,N_33753,N_33409);
or U34070 (N_34070,N_32419,N_33352);
and U34071 (N_34071,N_32211,N_32276);
xnor U34072 (N_34072,N_32905,N_32255);
nor U34073 (N_34073,N_32142,N_32332);
or U34074 (N_34074,N_33579,N_33515);
or U34075 (N_34075,N_33880,N_33627);
or U34076 (N_34076,N_32337,N_32102);
xnor U34077 (N_34077,N_33252,N_33431);
nor U34078 (N_34078,N_33975,N_32708);
and U34079 (N_34079,N_33169,N_32683);
nand U34080 (N_34080,N_33973,N_32443);
nand U34081 (N_34081,N_33477,N_33981);
nand U34082 (N_34082,N_33452,N_33333);
and U34083 (N_34083,N_32705,N_33176);
or U34084 (N_34084,N_32789,N_32836);
nand U34085 (N_34085,N_32158,N_33164);
nand U34086 (N_34086,N_32204,N_32376);
and U34087 (N_34087,N_32751,N_33989);
xnor U34088 (N_34088,N_33827,N_33396);
and U34089 (N_34089,N_32516,N_33341);
or U34090 (N_34090,N_33540,N_33179);
and U34091 (N_34091,N_32587,N_33980);
nand U34092 (N_34092,N_32182,N_33806);
xor U34093 (N_34093,N_33680,N_32582);
xnor U34094 (N_34094,N_32778,N_32932);
nand U34095 (N_34095,N_32133,N_32660);
or U34096 (N_34096,N_33072,N_32225);
xor U34097 (N_34097,N_33896,N_32922);
or U34098 (N_34098,N_32819,N_32925);
or U34099 (N_34099,N_33326,N_32231);
and U34100 (N_34100,N_33644,N_32992);
and U34101 (N_34101,N_33033,N_32219);
nand U34102 (N_34102,N_33555,N_33646);
xnor U34103 (N_34103,N_33849,N_33281);
or U34104 (N_34104,N_33442,N_33243);
or U34105 (N_34105,N_32001,N_33300);
nand U34106 (N_34106,N_33191,N_33612);
nor U34107 (N_34107,N_32471,N_32038);
or U34108 (N_34108,N_32147,N_32300);
and U34109 (N_34109,N_32791,N_33251);
xnor U34110 (N_34110,N_32155,N_33007);
nand U34111 (N_34111,N_33054,N_32193);
and U34112 (N_34112,N_33699,N_32094);
nand U34113 (N_34113,N_33532,N_32604);
xor U34114 (N_34114,N_33622,N_32489);
nand U34115 (N_34115,N_32192,N_32026);
nor U34116 (N_34116,N_32938,N_32854);
nor U34117 (N_34117,N_32698,N_32458);
or U34118 (N_34118,N_32595,N_32676);
nor U34119 (N_34119,N_33487,N_32908);
xor U34120 (N_34120,N_32409,N_32766);
nand U34121 (N_34121,N_32849,N_32336);
xor U34122 (N_34122,N_33456,N_32633);
and U34123 (N_34123,N_33803,N_32974);
nand U34124 (N_34124,N_32949,N_32130);
and U34125 (N_34125,N_33138,N_32696);
or U34126 (N_34126,N_33031,N_32392);
nand U34127 (N_34127,N_32872,N_33562);
nand U34128 (N_34128,N_32551,N_33649);
xor U34129 (N_34129,N_32031,N_33267);
or U34130 (N_34130,N_32240,N_32128);
or U34131 (N_34131,N_33686,N_33939);
or U34132 (N_34132,N_33205,N_32375);
nand U34133 (N_34133,N_32400,N_32030);
and U34134 (N_34134,N_33797,N_33717);
nor U34135 (N_34135,N_32120,N_33589);
nand U34136 (N_34136,N_32697,N_33694);
or U34137 (N_34137,N_33242,N_33808);
xor U34138 (N_34138,N_33365,N_32253);
nor U34139 (N_34139,N_33773,N_33538);
xor U34140 (N_34140,N_32691,N_33469);
or U34141 (N_34141,N_32799,N_33906);
xor U34142 (N_34142,N_33316,N_33162);
or U34143 (N_34143,N_32188,N_32416);
nor U34144 (N_34144,N_32893,N_32618);
xor U34145 (N_34145,N_32257,N_33483);
nor U34146 (N_34146,N_33768,N_32517);
nor U34147 (N_34147,N_33493,N_33701);
nand U34148 (N_34148,N_32174,N_33729);
nor U34149 (N_34149,N_32762,N_32134);
nand U34150 (N_34150,N_32976,N_32273);
nand U34151 (N_34151,N_33926,N_32731);
nor U34152 (N_34152,N_33438,N_33344);
nand U34153 (N_34153,N_33204,N_32674);
or U34154 (N_34154,N_32752,N_33317);
xor U34155 (N_34155,N_33818,N_32341);
and U34156 (N_34156,N_32601,N_33367);
xnor U34157 (N_34157,N_33741,N_33387);
nand U34158 (N_34158,N_33463,N_33807);
or U34159 (N_34159,N_33507,N_33721);
and U34160 (N_34160,N_32474,N_33368);
and U34161 (N_34161,N_33790,N_32093);
or U34162 (N_34162,N_32815,N_32748);
or U34163 (N_34163,N_32754,N_32741);
or U34164 (N_34164,N_32572,N_33949);
and U34165 (N_34165,N_32804,N_33467);
and U34166 (N_34166,N_32014,N_32459);
nand U34167 (N_34167,N_32853,N_32101);
nor U34168 (N_34168,N_33581,N_32999);
nand U34169 (N_34169,N_32704,N_33247);
nand U34170 (N_34170,N_32449,N_33858);
nor U34171 (N_34171,N_32294,N_32363);
nor U34172 (N_34172,N_32206,N_33834);
or U34173 (N_34173,N_32977,N_32321);
and U34174 (N_34174,N_32502,N_32575);
and U34175 (N_34175,N_33158,N_32947);
nor U34176 (N_34176,N_32055,N_32738);
nand U34177 (N_34177,N_33016,N_33836);
or U34178 (N_34178,N_33677,N_33777);
or U34179 (N_34179,N_33319,N_32726);
nor U34180 (N_34180,N_33023,N_33787);
xnor U34181 (N_34181,N_32615,N_32956);
xor U34182 (N_34182,N_33505,N_32993);
nand U34183 (N_34183,N_32484,N_33462);
nor U34184 (N_34184,N_32934,N_32724);
or U34185 (N_34185,N_32839,N_32883);
xor U34186 (N_34186,N_32229,N_32028);
and U34187 (N_34187,N_33795,N_32512);
and U34188 (N_34188,N_32597,N_33566);
nand U34189 (N_34189,N_33044,N_32359);
or U34190 (N_34190,N_33454,N_32773);
and U34191 (N_34191,N_33284,N_33419);
and U34192 (N_34192,N_32610,N_33804);
xor U34193 (N_34193,N_32728,N_33755);
and U34194 (N_34194,N_32611,N_33395);
or U34195 (N_34195,N_33372,N_32184);
nand U34196 (N_34196,N_33953,N_32667);
or U34197 (N_34197,N_33090,N_32536);
xor U34198 (N_34198,N_33552,N_33758);
xnor U34199 (N_34199,N_32509,N_33119);
or U34200 (N_34200,N_33881,N_33071);
nor U34201 (N_34201,N_33286,N_33605);
nand U34202 (N_34202,N_33748,N_33099);
nor U34203 (N_34203,N_33743,N_33219);
nor U34204 (N_34204,N_33342,N_32650);
xor U34205 (N_34205,N_32281,N_33160);
nor U34206 (N_34206,N_32861,N_33514);
xor U34207 (N_34207,N_32609,N_32537);
or U34208 (N_34208,N_32625,N_33468);
xnor U34209 (N_34209,N_33635,N_33020);
nand U34210 (N_34210,N_33910,N_32916);
nor U34211 (N_34211,N_33390,N_32214);
or U34212 (N_34212,N_33272,N_33705);
nand U34213 (N_34213,N_33700,N_32552);
nand U34214 (N_34214,N_32427,N_32790);
nor U34215 (N_34215,N_32948,N_33837);
and U34216 (N_34216,N_33757,N_33026);
nor U34217 (N_34217,N_32085,N_32213);
nand U34218 (N_34218,N_32807,N_32630);
and U34219 (N_34219,N_33315,N_32437);
and U34220 (N_34220,N_33545,N_32812);
or U34221 (N_34221,N_32593,N_33141);
nand U34222 (N_34222,N_32221,N_32432);
and U34223 (N_34223,N_33908,N_32886);
xnor U34224 (N_34224,N_33436,N_33561);
and U34225 (N_34225,N_33056,N_32648);
xnor U34226 (N_34226,N_33118,N_33921);
and U34227 (N_34227,N_33793,N_33551);
xor U34228 (N_34228,N_33410,N_32361);
or U34229 (N_34229,N_33959,N_33230);
or U34230 (N_34230,N_32640,N_32685);
xnor U34231 (N_34231,N_32342,N_32758);
nand U34232 (N_34232,N_33574,N_33256);
nand U34233 (N_34233,N_33868,N_32672);
nand U34234 (N_34234,N_33450,N_33525);
and U34235 (N_34235,N_32478,N_32656);
nor U34236 (N_34236,N_32844,N_32260);
nand U34237 (N_34237,N_33309,N_33691);
or U34238 (N_34238,N_33312,N_32797);
or U34239 (N_34239,N_33327,N_32786);
xnor U34240 (N_34240,N_32091,N_33335);
xnor U34241 (N_34241,N_33893,N_32431);
and U34242 (N_34242,N_32370,N_33898);
and U34243 (N_34243,N_33259,N_33990);
and U34244 (N_34244,N_33541,N_33572);
xnor U34245 (N_34245,N_32312,N_33511);
or U34246 (N_34246,N_32122,N_33723);
and U34247 (N_34247,N_33671,N_33979);
nor U34248 (N_34248,N_32242,N_32970);
and U34249 (N_34249,N_32486,N_32497);
and U34250 (N_34250,N_33003,N_32968);
nand U34251 (N_34251,N_33345,N_32613);
or U34252 (N_34252,N_32494,N_33962);
or U34253 (N_34253,N_33628,N_32288);
xnor U34254 (N_34254,N_33197,N_33651);
or U34255 (N_34255,N_32313,N_33132);
xor U34256 (N_34256,N_33775,N_32360);
nand U34257 (N_34257,N_33134,N_32510);
or U34258 (N_34258,N_33934,N_33185);
nor U34259 (N_34259,N_32258,N_32243);
or U34260 (N_34260,N_32951,N_32394);
nor U34261 (N_34261,N_32515,N_32903);
xor U34262 (N_34262,N_33604,N_33583);
xnor U34263 (N_34263,N_32061,N_33135);
and U34264 (N_34264,N_32869,N_33528);
xor U34265 (N_34265,N_33708,N_33550);
xnor U34266 (N_34266,N_33839,N_32435);
and U34267 (N_34267,N_33967,N_33210);
xor U34268 (N_34268,N_33856,N_33883);
nand U34269 (N_34269,N_33482,N_32961);
nor U34270 (N_34270,N_32851,N_33346);
and U34271 (N_34271,N_32612,N_33472);
nand U34272 (N_34272,N_32631,N_32000);
nand U34273 (N_34273,N_32713,N_33864);
and U34274 (N_34274,N_33626,N_33960);
nand U34275 (N_34275,N_32901,N_32840);
and U34276 (N_34276,N_32075,N_33394);
xor U34277 (N_34277,N_33992,N_33978);
nor U34278 (N_34278,N_32309,N_33789);
nand U34279 (N_34279,N_32450,N_33283);
nand U34280 (N_34280,N_33587,N_32441);
or U34281 (N_34281,N_32902,N_33430);
nand U34282 (N_34282,N_32334,N_33718);
and U34283 (N_34283,N_32928,N_33322);
and U34284 (N_34284,N_32350,N_32177);
and U34285 (N_34285,N_32153,N_33064);
and U34286 (N_34286,N_32396,N_33079);
nand U34287 (N_34287,N_33599,N_33142);
xnor U34288 (N_34288,N_32910,N_32793);
and U34289 (N_34289,N_32296,N_32256);
or U34290 (N_34290,N_32720,N_32451);
and U34291 (N_34291,N_33576,N_32139);
nand U34292 (N_34292,N_33117,N_33930);
or U34293 (N_34293,N_32248,N_32271);
nand U34294 (N_34294,N_32554,N_32149);
nor U34295 (N_34295,N_33995,N_32436);
and U34296 (N_34296,N_32306,N_32892);
or U34297 (N_34297,N_33631,N_32605);
nor U34298 (N_34298,N_33114,N_33903);
or U34299 (N_34299,N_33328,N_33674);
nand U34300 (N_34300,N_32740,N_33682);
xor U34301 (N_34301,N_32366,N_32472);
xor U34302 (N_34302,N_32614,N_33776);
and U34303 (N_34303,N_33121,N_33325);
and U34304 (N_34304,N_32803,N_32052);
xor U34305 (N_34305,N_33879,N_32475);
and U34306 (N_34306,N_32556,N_32216);
or U34307 (N_34307,N_33662,N_33434);
and U34308 (N_34308,N_33222,N_33656);
nor U34309 (N_34309,N_33684,N_32957);
or U34310 (N_34310,N_33867,N_32870);
and U34311 (N_34311,N_33560,N_32924);
nor U34312 (N_34312,N_32212,N_33404);
nand U34313 (N_34313,N_33095,N_32131);
or U34314 (N_34314,N_32716,N_33475);
nand U34315 (N_34315,N_32818,N_33542);
nor U34316 (N_34316,N_33902,N_33280);
nand U34317 (N_34317,N_32003,N_32152);
xnor U34318 (N_34318,N_33843,N_32379);
and U34319 (N_34319,N_32719,N_33660);
and U34320 (N_34320,N_33888,N_33218);
or U34321 (N_34321,N_33266,N_33544);
nor U34322 (N_34322,N_32317,N_33749);
nor U34323 (N_34323,N_33403,N_32592);
or U34324 (N_34324,N_33740,N_32616);
and U34325 (N_34325,N_32580,N_32507);
nor U34326 (N_34326,N_32721,N_32531);
and U34327 (N_34327,N_33152,N_33202);
and U34328 (N_34328,N_32011,N_33968);
and U34329 (N_34329,N_32286,N_33624);
nand U34330 (N_34330,N_32107,N_33799);
nand U34331 (N_34331,N_33711,N_32989);
or U34332 (N_34332,N_32774,N_33276);
nand U34333 (N_34333,N_33416,N_33109);
xnor U34334 (N_34334,N_32487,N_33539);
and U34335 (N_34335,N_32064,N_32062);
and U34336 (N_34336,N_33330,N_33527);
nor U34337 (N_34337,N_32636,N_32937);
nand U34338 (N_34338,N_33821,N_33490);
nor U34339 (N_34339,N_33417,N_32542);
nand U34340 (N_34340,N_32561,N_33678);
nor U34341 (N_34341,N_32743,N_32909);
nand U34342 (N_34342,N_32960,N_33010);
or U34343 (N_34343,N_32167,N_33318);
nor U34344 (N_34344,N_33041,N_32401);
or U34345 (N_34345,N_32996,N_32405);
or U34346 (N_34346,N_33000,N_33983);
nor U34347 (N_34347,N_32945,N_32828);
nand U34348 (N_34348,N_32251,N_33851);
and U34349 (N_34349,N_32860,N_33929);
nor U34350 (N_34350,N_33015,N_33715);
or U34351 (N_34351,N_33943,N_33106);
or U34352 (N_34352,N_32759,N_32821);
or U34353 (N_34353,N_33767,N_32862);
and U34354 (N_34354,N_32339,N_33945);
nand U34355 (N_34355,N_33569,N_33443);
nor U34356 (N_34356,N_32824,N_32374);
xor U34357 (N_34357,N_33565,N_33977);
xor U34358 (N_34358,N_33005,N_32162);
or U34359 (N_34359,N_33629,N_32440);
nand U34360 (N_34360,N_32287,N_33263);
nand U34361 (N_34361,N_32596,N_32746);
and U34362 (N_34362,N_32569,N_32749);
nor U34363 (N_34363,N_33186,N_33916);
xnor U34364 (N_34364,N_32984,N_33642);
or U34365 (N_34365,N_33290,N_32635);
xor U34366 (N_34366,N_32780,N_32422);
and U34367 (N_34367,N_33955,N_33151);
xor U34368 (N_34368,N_33088,N_32254);
or U34369 (N_34369,N_33647,N_33941);
or U34370 (N_34370,N_32378,N_32975);
nand U34371 (N_34371,N_32492,N_32051);
and U34372 (N_34372,N_32498,N_32393);
or U34373 (N_34373,N_32602,N_33947);
or U34374 (N_34374,N_32987,N_33963);
xnor U34375 (N_34375,N_33603,N_32732);
nand U34376 (N_34376,N_32567,N_33332);
or U34377 (N_34377,N_32942,N_32384);
nand U34378 (N_34378,N_32263,N_32600);
and U34379 (N_34379,N_33040,N_33128);
xnor U34380 (N_34380,N_33925,N_32426);
and U34381 (N_34381,N_32010,N_33254);
xor U34382 (N_34382,N_32025,N_33004);
xnor U34383 (N_34383,N_33497,N_33761);
nand U34384 (N_34384,N_33349,N_33418);
and U34385 (N_34385,N_32890,N_32663);
or U34386 (N_34386,N_33167,N_33009);
nor U34387 (N_34387,N_32558,N_33065);
and U34388 (N_34388,N_33092,N_33593);
nand U34389 (N_34389,N_32086,N_33194);
and U34390 (N_34390,N_32164,N_32461);
xnor U34391 (N_34391,N_33725,N_32855);
or U34392 (N_34392,N_32388,N_33492);
and U34393 (N_34393,N_32320,N_33607);
and U34394 (N_34394,N_32037,N_32929);
nand U34395 (N_34395,N_33537,N_32382);
or U34396 (N_34396,N_33397,N_33504);
or U34397 (N_34397,N_32168,N_33832);
nand U34398 (N_34398,N_32303,N_33361);
and U34399 (N_34399,N_33081,N_33580);
or U34400 (N_34400,N_32476,N_33917);
or U34401 (N_34401,N_33950,N_32148);
xnor U34402 (N_34402,N_33148,N_33047);
xor U34403 (N_34403,N_32060,N_32012);
nand U34404 (N_34404,N_32163,N_32816);
nor U34405 (N_34405,N_32639,N_32289);
xor U34406 (N_34406,N_32386,N_32081);
nor U34407 (N_34407,N_32203,N_33306);
xor U34408 (N_34408,N_32228,N_33369);
xor U34409 (N_34409,N_32842,N_32036);
or U34410 (N_34410,N_33356,N_33841);
or U34411 (N_34411,N_33411,N_32940);
and U34412 (N_34412,N_33445,N_33029);
xnor U34413 (N_34413,N_32326,N_32009);
nand U34414 (N_34414,N_32668,N_33274);
nor U34415 (N_34415,N_32881,N_33291);
and U34416 (N_34416,N_32680,N_32763);
xor U34417 (N_34417,N_32907,N_33224);
and U34418 (N_34418,N_32621,N_33264);
nand U34419 (N_34419,N_32146,N_33089);
nor U34420 (N_34420,N_32735,N_33865);
xnor U34421 (N_34421,N_33078,N_33559);
or U34422 (N_34422,N_32785,N_33122);
xnor U34423 (N_34423,N_32546,N_33812);
and U34424 (N_34424,N_33652,N_33408);
and U34425 (N_34425,N_33766,N_33261);
and U34426 (N_34426,N_33951,N_33944);
xor U34427 (N_34427,N_32215,N_33533);
xor U34428 (N_34428,N_33428,N_33172);
nor U34429 (N_34429,N_33780,N_33124);
nand U34430 (N_34430,N_33859,N_32776);
xnor U34431 (N_34431,N_33704,N_32895);
nor U34432 (N_34432,N_33297,N_33842);
nand U34433 (N_34433,N_32187,N_32760);
nand U34434 (N_34434,N_32328,N_32047);
and U34435 (N_34435,N_32661,N_32325);
or U34436 (N_34436,N_32527,N_33268);
xnor U34437 (N_34437,N_32747,N_32559);
xor U34438 (N_34438,N_33190,N_32562);
or U34439 (N_34439,N_33911,N_33573);
nor U34440 (N_34440,N_33618,N_32808);
and U34441 (N_34441,N_32550,N_32997);
or U34442 (N_34442,N_33722,N_33805);
nand U34443 (N_34443,N_33695,N_33156);
nor U34444 (N_34444,N_32397,N_33553);
nand U34445 (N_34445,N_33894,N_32125);
or U34446 (N_34446,N_33055,N_33771);
nor U34447 (N_34447,N_33228,N_32470);
nor U34448 (N_34448,N_33378,N_32353);
nand U34449 (N_34449,N_32829,N_33696);
or U34450 (N_34450,N_33783,N_32730);
or U34451 (N_34451,N_32180,N_32831);
or U34452 (N_34452,N_33847,N_32016);
and U34453 (N_34453,N_32245,N_32481);
and U34454 (N_34454,N_33223,N_33498);
nor U34455 (N_34455,N_33076,N_32383);
or U34456 (N_34456,N_32327,N_32669);
or U34457 (N_34457,N_33855,N_32822);
and U34458 (N_34458,N_32008,N_32946);
xnor U34459 (N_34459,N_32980,N_32826);
nand U34460 (N_34460,N_33157,N_32467);
or U34461 (N_34461,N_32377,N_33425);
xnor U34462 (N_34462,N_33059,N_33829);
or U34463 (N_34463,N_33042,N_32514);
nor U34464 (N_34464,N_33495,N_32573);
nor U34465 (N_34465,N_32577,N_33008);
nor U34466 (N_34466,N_32814,N_32117);
or U34467 (N_34467,N_32677,N_33248);
xnor U34468 (N_34468,N_33439,N_33024);
or U34469 (N_34469,N_32688,N_32852);
nor U34470 (N_34470,N_32183,N_32298);
nand U34471 (N_34471,N_33509,N_32845);
or U34472 (N_34472,N_32015,N_33073);
or U34473 (N_34473,N_32410,N_33937);
or U34474 (N_34474,N_33125,N_33873);
nor U34475 (N_34475,N_33305,N_33129);
or U34476 (N_34476,N_33501,N_32408);
nand U34477 (N_34477,N_33918,N_32295);
xnor U34478 (N_34478,N_32671,N_33739);
nor U34479 (N_34479,N_33681,N_32230);
and U34480 (N_34480,N_32132,N_33970);
xor U34481 (N_34481,N_33444,N_32054);
nand U34482 (N_34482,N_33993,N_32072);
xnor U34483 (N_34483,N_32395,N_32693);
nand U34484 (N_34484,N_32355,N_33423);
xnor U34485 (N_34485,N_32768,N_33100);
xnor U34486 (N_34486,N_33102,N_33640);
or U34487 (N_34487,N_32265,N_32491);
and U34488 (N_34488,N_32863,N_32269);
nand U34489 (N_34489,N_33240,N_32590);
xnor U34490 (N_34490,N_33137,N_32927);
nor U34491 (N_34491,N_33554,N_33273);
and U34492 (N_34492,N_33277,N_33320);
or U34493 (N_34493,N_33257,N_33299);
or U34494 (N_34494,N_33449,N_33478);
or U34495 (N_34495,N_33853,N_32501);
nand U34496 (N_34496,N_33380,N_33216);
xor U34497 (N_34497,N_33457,N_33810);
nand U34498 (N_34498,N_33706,N_33130);
xor U34499 (N_34499,N_33698,N_33519);
nand U34500 (N_34500,N_33002,N_32714);
or U34501 (N_34501,N_32083,N_32197);
nor U34502 (N_34502,N_32617,N_32865);
nor U34503 (N_34503,N_33195,N_33249);
or U34504 (N_34504,N_32898,N_33809);
and U34505 (N_34505,N_33057,N_32136);
xnor U34506 (N_34506,N_32238,N_32119);
nor U34507 (N_34507,N_32191,N_32889);
or U34508 (N_34508,N_32917,N_32239);
nand U34509 (N_34509,N_32035,N_32770);
and U34510 (N_34510,N_33710,N_32439);
xor U34511 (N_34511,N_32711,N_32402);
nor U34512 (N_34512,N_32448,N_32643);
nor U34513 (N_34513,N_32706,N_32057);
xor U34514 (N_34514,N_32227,N_32800);
and U34515 (N_34515,N_33602,N_33590);
and U34516 (N_34516,N_32259,N_33143);
xnor U34517 (N_34517,N_32998,N_33289);
nor U34518 (N_34518,N_33976,N_33208);
and U34519 (N_34519,N_33049,N_32348);
nor U34520 (N_34520,N_32876,N_33175);
or U34521 (N_34521,N_32703,N_32483);
and U34522 (N_34522,N_32420,N_33168);
or U34523 (N_34523,N_33523,N_33080);
xor U34524 (N_34524,N_33494,N_32331);
xor U34525 (N_34525,N_32857,N_33066);
or U34526 (N_34526,N_32586,N_32659);
xnor U34527 (N_34527,N_32871,N_33150);
nor U34528 (N_34528,N_33295,N_33203);
xor U34529 (N_34529,N_32172,N_33211);
or U34530 (N_34530,N_32873,N_33791);
nand U34531 (N_34531,N_33366,N_33928);
xnor U34532 (N_34532,N_32106,N_33006);
and U34533 (N_34533,N_32202,N_33302);
nand U34534 (N_34534,N_32835,N_33638);
and U34535 (N_34535,N_33427,N_32662);
or U34536 (N_34536,N_33426,N_33549);
or U34537 (N_34537,N_33407,N_32505);
nor U34538 (N_34538,N_32404,N_33012);
or U34539 (N_34539,N_33857,N_32354);
nor U34540 (N_34540,N_32301,N_33909);
or U34541 (N_34541,N_33630,N_33401);
nand U34542 (N_34542,N_32335,N_32710);
or U34543 (N_34543,N_33013,N_33253);
nor U34544 (N_34544,N_32456,N_32566);
nor U34545 (N_34545,N_32687,N_32526);
nand U34546 (N_34546,N_33389,N_33846);
and U34547 (N_34547,N_32707,N_32170);
xor U34548 (N_34548,N_32039,N_32365);
nor U34549 (N_34549,N_33719,N_32319);
xor U34550 (N_34550,N_33601,N_32877);
nand U34551 (N_34551,N_33189,N_33661);
or U34552 (N_34552,N_33161,N_33094);
nand U34553 (N_34553,N_33616,N_33920);
nand U34554 (N_34554,N_33728,N_33474);
xnor U34555 (N_34555,N_32264,N_33258);
nor U34556 (N_34556,N_32438,N_32433);
xor U34557 (N_34557,N_32113,N_33524);
and U34558 (N_34558,N_32233,N_33051);
or U34559 (N_34559,N_32198,N_33611);
xor U34560 (N_34560,N_32411,N_33437);
or U34561 (N_34561,N_33563,N_32530);
xnor U34562 (N_34562,N_33085,N_33956);
nand U34563 (N_34563,N_32900,N_32651);
xor U34564 (N_34564,N_33091,N_33933);
nor U34565 (N_34565,N_33227,N_32966);
nand U34566 (N_34566,N_32430,N_33927);
nor U34567 (N_34567,N_32518,N_32841);
and U34568 (N_34568,N_32788,N_33900);
xnor U34569 (N_34569,N_33531,N_32499);
xor U34570 (N_34570,N_32407,N_33421);
or U34571 (N_34571,N_33720,N_32040);
nand U34572 (N_34572,N_32480,N_32272);
nand U34573 (N_34573,N_33954,N_33193);
nand U34574 (N_34574,N_32958,N_33802);
nand U34575 (N_34575,N_32002,N_32368);
nand U34576 (N_34576,N_33371,N_32563);
or U34577 (N_34577,N_32315,N_32699);
or U34578 (N_34578,N_33052,N_32535);
xor U34579 (N_34579,N_32465,N_33619);
nor U34580 (N_34580,N_33575,N_33491);
nand U34581 (N_34581,N_33932,N_32071);
and U34582 (N_34582,N_32316,N_32764);
xnor U34583 (N_34583,N_33557,N_32775);
nor U34584 (N_34584,N_32105,N_32232);
or U34585 (N_34585,N_32205,N_33101);
xor U34586 (N_34586,N_33952,N_33582);
xor U34587 (N_34587,N_33591,N_32123);
xor U34588 (N_34588,N_33759,N_32583);
and U34589 (N_34589,N_32866,N_33357);
and U34590 (N_34590,N_32810,N_33679);
or U34591 (N_34591,N_32181,N_32969);
nor U34592 (N_34592,N_32059,N_32695);
nand U34593 (N_34593,N_32506,N_32293);
and U34594 (N_34594,N_33331,N_32990);
nand U34595 (N_34595,N_32528,N_32270);
nor U34596 (N_34596,N_32952,N_32837);
and U34597 (N_34597,N_32466,N_32200);
nor U34598 (N_34598,N_32073,N_32813);
nor U34599 (N_34599,N_33584,N_33350);
nor U34600 (N_34600,N_32371,N_32078);
xor U34601 (N_34601,N_33237,N_33375);
and U34602 (N_34602,N_33988,N_32750);
xor U34603 (N_34603,N_32504,N_33279);
nand U34604 (N_34604,N_33828,N_32241);
and U34605 (N_34605,N_32063,N_33781);
nand U34606 (N_34606,N_33785,N_33875);
nor U34607 (N_34607,N_33018,N_33307);
nand U34608 (N_34608,N_33120,N_32261);
nor U34609 (N_34609,N_33096,N_33641);
xor U34610 (N_34610,N_33053,N_33348);
xor U34611 (N_34611,N_32971,N_33458);
or U34612 (N_34612,N_33196,N_32129);
xor U34613 (N_34613,N_33282,N_32521);
and U34614 (N_34614,N_32208,N_32171);
nand U34615 (N_34615,N_32915,N_32460);
or U34616 (N_34616,N_33275,N_33201);
or U34617 (N_34617,N_33792,N_33835);
xnor U34618 (N_34618,N_33386,N_32756);
and U34619 (N_34619,N_33985,N_33811);
or U34620 (N_34620,N_33337,N_32868);
nor U34621 (N_34621,N_32846,N_32285);
xnor U34622 (N_34622,N_32644,N_32684);
nand U34623 (N_34623,N_33481,N_32004);
nor U34624 (N_34624,N_32389,N_33025);
nor U34625 (N_34625,N_32283,N_33665);
and U34626 (N_34626,N_32352,N_33136);
xnor U34627 (N_34627,N_33163,N_33473);
nor U34628 (N_34628,N_32729,N_33139);
and U34629 (N_34629,N_33255,N_33769);
nor U34630 (N_34630,N_32745,N_32920);
xnor U34631 (N_34631,N_32959,N_32292);
and U34632 (N_34632,N_33429,N_33212);
xnor U34633 (N_34633,N_33039,N_33948);
xor U34634 (N_34634,N_33178,N_32811);
and U34635 (N_34635,N_32343,N_33571);
or U34636 (N_34636,N_33621,N_33779);
and U34637 (N_34637,N_33982,N_33633);
and U34638 (N_34638,N_33278,N_32185);
xnor U34639 (N_34639,N_33987,N_33354);
xnor U34640 (N_34640,N_32346,N_32985);
nand U34641 (N_34641,N_32833,N_33940);
xnor U34642 (N_34642,N_32673,N_32282);
xnor U34643 (N_34643,N_32150,N_33082);
nor U34644 (N_34644,N_33413,N_32013);
xnor U34645 (N_34645,N_33782,N_32645);
or U34646 (N_34646,N_32385,N_32549);
xnor U34647 (N_34647,N_32372,N_32100);
nor U34648 (N_34648,N_33184,N_32769);
nand U34649 (N_34649,N_32783,N_32911);
xor U34650 (N_34650,N_32568,N_33019);
and U34651 (N_34651,N_33270,N_33234);
nand U34652 (N_34652,N_32290,N_32324);
nand U34653 (N_34653,N_33377,N_32115);
nand U34654 (N_34654,N_32275,N_33850);
and U34655 (N_34655,N_33314,N_32744);
and U34656 (N_34656,N_33503,N_33713);
nor U34657 (N_34657,N_33685,N_33383);
xor U34658 (N_34658,N_32541,N_33664);
and U34659 (N_34659,N_33145,N_32415);
nand U34660 (N_34660,N_32357,N_32658);
or U34661 (N_34661,N_32121,N_33225);
xor U34662 (N_34662,N_33174,N_33321);
or U34663 (N_34663,N_32362,N_33600);
xor U34664 (N_34664,N_33738,N_33965);
xor U34665 (N_34665,N_33420,N_32399);
xor U34666 (N_34666,N_32017,N_33816);
nand U34667 (N_34667,N_32310,N_33615);
nor U34668 (N_34668,N_32723,N_33824);
or U34669 (N_34669,N_32249,N_32686);
nor U34670 (N_34670,N_33744,N_33637);
or U34671 (N_34671,N_33676,N_33360);
and U34672 (N_34672,N_33522,N_33355);
nand U34673 (N_34673,N_33311,N_32953);
nor U34674 (N_34674,N_33464,N_32144);
nor U34675 (N_34675,N_32490,N_32140);
and U34676 (N_34676,N_33294,N_33712);
and U34677 (N_34677,N_33166,N_32544);
nor U34678 (N_34678,N_32539,N_33825);
nor U34679 (N_34679,N_33113,N_33246);
xnor U34680 (N_34680,N_32141,N_33432);
xnor U34681 (N_34681,N_32878,N_32496);
nand U34682 (N_34682,N_32859,N_32154);
or U34683 (N_34683,N_32717,N_33236);
and U34684 (N_34684,N_33440,N_33060);
and U34685 (N_34685,N_33453,N_33206);
xor U34686 (N_34686,N_32262,N_32820);
and U34687 (N_34687,N_32160,N_32972);
xor U34688 (N_34688,N_33127,N_32340);
xor U34689 (N_34689,N_32024,N_33689);
and U34690 (N_34690,N_33517,N_33265);
and U34691 (N_34691,N_32045,N_32454);
nor U34692 (N_34692,N_32066,N_32199);
nand U34693 (N_34693,N_33675,N_32817);
nor U34694 (N_34694,N_32457,N_32642);
nand U34695 (N_34695,N_33021,N_32224);
or U34696 (N_34696,N_32692,N_33862);
nand U34697 (N_34697,N_33414,N_33964);
or U34698 (N_34698,N_32477,N_32210);
and U34699 (N_34699,N_33343,N_32220);
nand U34700 (N_34700,N_32165,N_33424);
xnor U34701 (N_34701,N_33149,N_32864);
nand U34702 (N_34702,N_32209,N_32500);
nor U34703 (N_34703,N_32579,N_33822);
xnor U34704 (N_34704,N_32096,N_33577);
nor U34705 (N_34705,N_33754,N_33422);
or U34706 (N_34706,N_33226,N_32065);
or U34707 (N_34707,N_33188,N_33070);
nand U34708 (N_34708,N_33232,N_33935);
nor U34709 (N_34709,N_33942,N_32381);
and U34710 (N_34710,N_32114,N_33133);
and U34711 (N_34711,N_33732,N_33338);
and U34712 (N_34712,N_32157,N_33530);
nand U34713 (N_34713,N_33736,N_32417);
nor U34714 (N_34714,N_33546,N_33751);
xnor U34715 (N_34715,N_32338,N_33339);
or U34716 (N_34716,N_33734,N_33521);
nand U34717 (N_34717,N_33688,N_33506);
or U34718 (N_34718,N_32936,N_32179);
nor U34719 (N_34719,N_33489,N_32843);
and U34720 (N_34720,N_32941,N_32237);
or U34721 (N_34721,N_33996,N_33666);
nand U34722 (N_34722,N_33568,N_33400);
nor U34723 (N_34723,N_33670,N_33126);
nand U34724 (N_34724,N_33891,N_32646);
nand U34725 (N_34725,N_32423,N_33433);
nand U34726 (N_34726,N_33221,N_33870);
xor U34727 (N_34727,N_32806,N_32576);
or U34728 (N_34728,N_33643,N_32986);
xnor U34729 (N_34729,N_32508,N_32682);
or U34730 (N_34730,N_33376,N_33620);
xnor U34731 (N_34731,N_33614,N_33351);
or U34732 (N_34732,N_32446,N_32196);
nor U34733 (N_34733,N_32570,N_32022);
or U34734 (N_34734,N_32734,N_33045);
nand U34735 (N_34735,N_33788,N_32689);
nor U34736 (N_34736,N_32553,N_32795);
and U34737 (N_34737,N_33609,N_33046);
xnor U34738 (N_34738,N_33648,N_32979);
nor U34739 (N_34739,N_32145,N_33324);
nand U34740 (N_34740,N_32983,N_33658);
or U34741 (N_34741,N_32574,N_32329);
xnor U34742 (N_34742,N_32588,N_33373);
nor U34743 (N_34743,N_33470,N_32097);
nand U34744 (N_34744,N_33075,N_33912);
nand U34745 (N_34745,N_33235,N_32805);
nand U34746 (N_34746,N_33885,N_33874);
nand U34747 (N_34747,N_32598,N_32923);
or U34748 (N_34748,N_32899,N_32520);
and U34749 (N_34749,N_32794,N_33746);
or U34750 (N_34750,N_33742,N_33036);
and U34751 (N_34751,N_32006,N_33598);
xnor U34752 (N_34752,N_33050,N_32511);
nor U34753 (N_34753,N_33534,N_33840);
nand U34754 (N_34754,N_32111,N_32594);
nand U34755 (N_34755,N_32718,N_33882);
nand U34756 (N_34756,N_32195,N_33451);
nand U34757 (N_34757,N_33084,N_33597);
or U34758 (N_34758,N_32074,N_33488);
nand U34759 (N_34759,N_33262,N_33461);
nand U34760 (N_34760,N_32406,N_33831);
and U34761 (N_34761,N_32018,N_32832);
nor U34762 (N_34762,N_32885,N_33177);
or U34763 (N_34763,N_32207,N_32739);
nand U34764 (N_34764,N_32049,N_33890);
or U34765 (N_34765,N_32109,N_33465);
xnor U34766 (N_34766,N_32578,N_32755);
and U34767 (N_34767,N_33229,N_33231);
xor U34768 (N_34768,N_33518,N_33499);
or U34769 (N_34769,N_32079,N_33733);
xnor U34770 (N_34770,N_33323,N_32727);
and U34771 (N_34771,N_32299,N_33460);
nor U34772 (N_34772,N_32641,N_33871);
and U34773 (N_34773,N_33077,N_33876);
nor U34774 (N_34774,N_33625,N_33860);
nand U34775 (N_34775,N_33170,N_32981);
nand U34776 (N_34776,N_32268,N_32234);
or U34777 (N_34777,N_32867,N_33901);
and U34778 (N_34778,N_32761,N_33668);
xor U34779 (N_34779,N_32978,N_32973);
or U34780 (N_34780,N_32277,N_32442);
or U34781 (N_34781,N_33814,N_33358);
and U34782 (N_34782,N_32201,N_32629);
xnor U34783 (N_34783,N_33543,N_32623);
nand U34784 (N_34784,N_32652,N_32965);
and U34785 (N_34785,N_33623,N_32801);
or U34786 (N_34786,N_32124,N_32894);
xor U34787 (N_34787,N_33709,N_33730);
or U34788 (N_34788,N_33098,N_33946);
nand U34789 (N_34789,N_32364,N_32280);
nand U34790 (N_34790,N_33703,N_33657);
xnor U34791 (N_34791,N_32584,N_32143);
or U34792 (N_34792,N_33861,N_32522);
xnor U34793 (N_34793,N_33535,N_33111);
or U34794 (N_34794,N_33144,N_32007);
nor U34795 (N_34795,N_32880,N_33244);
xor U34796 (N_34796,N_32519,N_33786);
nor U34797 (N_34797,N_33774,N_33392);
and U34798 (N_34798,N_32884,N_32178);
xnor U34799 (N_34799,N_32244,N_33800);
nor U34800 (N_34800,N_33923,N_33913);
xor U34801 (N_34801,N_33147,N_32462);
and U34802 (N_34802,N_33724,N_33022);
xor U34803 (N_34803,N_32046,N_32913);
xor U34804 (N_34804,N_33063,N_33770);
nor U34805 (N_34805,N_32021,N_32127);
nor U34806 (N_34806,N_32624,N_32891);
or U34807 (N_34807,N_32784,N_33087);
and U34808 (N_34808,N_32463,N_32042);
xnor U34809 (N_34809,N_32781,N_32485);
or U34810 (N_34810,N_32874,N_32274);
xnor U34811 (N_34811,N_32186,N_32619);
and U34812 (N_34812,N_32311,N_33069);
or U34813 (N_34813,N_32302,N_32137);
and U34814 (N_34814,N_32856,N_32391);
nand U34815 (N_34815,N_32424,N_32882);
nand U34816 (N_34816,N_33391,N_33508);
and U34817 (N_34817,N_32387,N_32538);
or U34818 (N_34818,N_33707,N_32236);
nand U34819 (N_34819,N_32297,N_33347);
and U34820 (N_34820,N_33606,N_33697);
or U34821 (N_34821,N_32380,N_32452);
nand U34822 (N_34822,N_32020,N_33502);
nor U34823 (N_34823,N_33999,N_33512);
or U34824 (N_34824,N_33819,N_32967);
and U34825 (N_34825,N_33838,N_33123);
or U34826 (N_34826,N_33852,N_33220);
and U34827 (N_34827,N_32307,N_32991);
or U34828 (N_34828,N_32850,N_33972);
and U34829 (N_34829,N_32291,N_32943);
and U34830 (N_34830,N_33520,N_33287);
nor U34831 (N_34831,N_32250,N_32782);
and U34832 (N_34832,N_33669,N_32914);
and U34833 (N_34833,N_33984,N_32138);
nor U34834 (N_34834,N_32398,N_33068);
nor U34835 (N_34835,N_33914,N_33364);
nand U34836 (N_34836,N_33673,N_32926);
nor U34837 (N_34837,N_32627,N_33778);
or U34838 (N_34838,N_33260,N_33690);
xor U34839 (N_34839,N_33588,N_33564);
or U34840 (N_34840,N_32964,N_33104);
nor U34841 (N_34841,N_33765,N_32653);
nand U34842 (N_34842,N_33645,N_33215);
nor U34843 (N_34843,N_33884,N_32092);
and U34844 (N_34844,N_32571,N_33895);
or U34845 (N_34845,N_33037,N_33112);
nor U34846 (N_34846,N_32412,N_33058);
and U34847 (N_34847,N_32647,N_33570);
nand U34848 (N_34848,N_32921,N_32753);
nand U34849 (N_34849,N_32349,N_33659);
nand U34850 (N_34850,N_32675,N_33292);
and U34851 (N_34851,N_33526,N_32955);
xnor U34852 (N_34852,N_33727,N_33655);
nand U34853 (N_34853,N_33412,N_32792);
or U34854 (N_34854,N_32473,N_32176);
nor U34855 (N_34855,N_32879,N_32736);
xnor U34856 (N_34856,N_33567,N_32005);
nand U34857 (N_34857,N_33826,N_33250);
or U34858 (N_34858,N_32453,N_33854);
xnor U34859 (N_34859,N_33936,N_32772);
nor U34860 (N_34860,N_33296,N_33714);
nand U34861 (N_34861,N_32166,N_32190);
xnor U34862 (N_34862,N_33548,N_32838);
and U34863 (N_34863,N_32413,N_33107);
xnor U34864 (N_34864,N_32532,N_33672);
nand U34865 (N_34865,N_33702,N_32919);
nand U34866 (N_34866,N_32534,N_33904);
or U34867 (N_34867,N_32589,N_33271);
xnor U34868 (N_34868,N_33476,N_32033);
and U34869 (N_34869,N_33801,N_32304);
and U34870 (N_34870,N_33762,N_33406);
xor U34871 (N_34871,N_32414,N_33632);
nand U34872 (N_34872,N_32246,N_32962);
or U34873 (N_34873,N_33301,N_33513);
nor U34874 (N_34874,N_32733,N_33794);
and U34875 (N_34875,N_32628,N_32767);
or U34876 (N_34876,N_32252,N_33359);
and U34877 (N_34877,N_33116,N_32994);
xnor U34878 (N_34878,N_32524,N_32757);
or U34879 (N_34879,N_32545,N_32069);
nor U34880 (N_34880,N_33182,N_33585);
or U34881 (N_34881,N_33398,N_32077);
xnor U34882 (N_34882,N_32548,N_33887);
nor U34883 (N_34883,N_33115,N_33017);
and U34884 (N_34884,N_32345,N_32779);
nor U34885 (N_34885,N_32019,N_32678);
xor U34886 (N_34886,N_33233,N_32939);
and U34887 (N_34887,N_33869,N_32110);
or U34888 (N_34888,N_33154,N_33845);
nor U34889 (N_34889,N_33399,N_33610);
and U34890 (N_34890,N_33329,N_32565);
nand U34891 (N_34891,N_33986,N_32344);
nor U34892 (N_34892,N_32622,N_33747);
xnor U34893 (N_34893,N_32690,N_33796);
xor U34894 (N_34894,N_33153,N_32023);
nor U34895 (N_34895,N_33510,N_32701);
xor U34896 (N_34896,N_32118,N_32428);
or U34897 (N_34897,N_32825,N_33760);
or U34898 (N_34898,N_32543,N_32318);
xnor U34899 (N_34899,N_33415,N_33772);
xor U34900 (N_34900,N_33030,N_33093);
and U34901 (N_34901,N_33815,N_33213);
and U34902 (N_34902,N_32777,N_33032);
nor U34903 (N_34903,N_32043,N_33516);
nor U34904 (N_34904,N_33886,N_32809);
or U34905 (N_34905,N_33558,N_32222);
xor U34906 (N_34906,N_33500,N_33446);
nor U34907 (N_34907,N_33617,N_33001);
xnor U34908 (N_34908,N_32944,N_33878);
nand U34909 (N_34909,N_33556,N_33097);
and U34910 (N_34910,N_32173,N_33915);
xor U34911 (N_34911,N_33209,N_33308);
xor U34912 (N_34912,N_32314,N_32076);
and U34913 (N_34913,N_33336,N_33043);
and U34914 (N_34914,N_32284,N_33171);
or U34915 (N_34915,N_32351,N_33692);
or U34916 (N_34916,N_33241,N_33731);
nor U34917 (N_34917,N_33027,N_33435);
nor U34918 (N_34918,N_32560,N_33269);
xor U34919 (N_34919,N_32827,N_32533);
nor U34920 (N_34920,N_32084,N_33735);
xor U34921 (N_34921,N_33639,N_32887);
and U34922 (N_34922,N_32103,N_33405);
nand U34923 (N_34923,N_32135,N_32638);
nand U34924 (N_34924,N_32930,N_32367);
nor U34925 (N_34925,N_32390,N_33199);
nand U34926 (N_34926,N_32634,N_33997);
nand U34927 (N_34927,N_33924,N_32322);
nand U34928 (N_34928,N_33877,N_33830);
nand U34929 (N_34929,N_32954,N_33899);
or U34930 (N_34930,N_32603,N_32995);
xnor U34931 (N_34931,N_33048,N_33479);
or U34932 (N_34932,N_33067,N_32935);
and U34933 (N_34933,N_33388,N_32217);
and U34934 (N_34934,N_33726,N_32278);
xor U34935 (N_34935,N_33922,N_32637);
or U34936 (N_34936,N_32444,N_33496);
nand U34937 (N_34937,N_32787,N_33110);
and U34938 (N_34938,N_33961,N_33848);
and U34939 (N_34939,N_32112,N_32425);
or U34940 (N_34940,N_33784,N_33971);
xor U34941 (N_34941,N_33471,N_32963);
nor U34942 (N_34942,N_32464,N_32503);
and U34943 (N_34943,N_33663,N_32591);
xor U34944 (N_34944,N_32897,N_32888);
and U34945 (N_34945,N_32050,N_33486);
nor U34946 (N_34946,N_33217,N_32482);
xnor U34947 (N_34947,N_32982,N_33667);
and U34948 (N_34948,N_32665,N_32599);
nor U34949 (N_34949,N_32098,N_33239);
xor U34950 (N_34950,N_33866,N_32156);
or U34951 (N_34951,N_33165,N_33863);
nor U34952 (N_34952,N_32358,N_33173);
nor U34953 (N_34953,N_32429,N_32434);
nand U34954 (N_34954,N_33393,N_32070);
or U34955 (N_34955,N_33245,N_33687);
or U34956 (N_34956,N_32088,N_32194);
or U34957 (N_34957,N_33683,N_32333);
nor U34958 (N_34958,N_33334,N_32479);
or U34959 (N_34959,N_32666,N_32555);
and U34960 (N_34960,N_32090,N_32279);
nand U34961 (N_34961,N_32469,N_33536);
or U34962 (N_34962,N_32529,N_33529);
and U34963 (N_34963,N_32858,N_33693);
and U34964 (N_34964,N_33764,N_32712);
and U34965 (N_34965,N_33402,N_32034);
nor U34966 (N_34966,N_33957,N_32848);
nand U34967 (N_34967,N_32323,N_32161);
xnor U34968 (N_34968,N_32058,N_32655);
or U34969 (N_34969,N_33752,N_33187);
and U34970 (N_34970,N_32104,N_32933);
nor U34971 (N_34971,N_33931,N_32044);
nor U34972 (N_34972,N_33303,N_32223);
and U34973 (N_34973,N_32950,N_32445);
or U34974 (N_34974,N_33974,N_33592);
and U34975 (N_34975,N_32585,N_32488);
nor U34976 (N_34976,N_32834,N_33636);
xor U34977 (N_34977,N_33907,N_32032);
xnor U34978 (N_34978,N_33146,N_33596);
nand U34979 (N_34979,N_32151,N_33798);
xor U34980 (N_34980,N_32082,N_32765);
nor U34981 (N_34981,N_33374,N_32581);
nor U34982 (N_34982,N_32330,N_32608);
or U34983 (N_34983,N_33892,N_32126);
and U34984 (N_34984,N_33103,N_32403);
or U34985 (N_34985,N_32087,N_33362);
nand U34986 (N_34986,N_33991,N_32988);
nand U34987 (N_34987,N_33238,N_33384);
or U34988 (N_34988,N_33480,N_33181);
or U34989 (N_34989,N_33756,N_32169);
nand U34990 (N_34990,N_32068,N_33905);
or U34991 (N_34991,N_32694,N_32620);
nand U34992 (N_34992,N_32099,N_33086);
nor U34993 (N_34993,N_33613,N_33634);
xor U34994 (N_34994,N_32632,N_32918);
xnor U34995 (N_34995,N_33441,N_32048);
nor U34996 (N_34996,N_33938,N_33313);
xor U34997 (N_34997,N_33062,N_33820);
nor U34998 (N_34998,N_33459,N_32547);
xor U34999 (N_34999,N_32679,N_33547);
and U35000 (N_35000,N_33599,N_33958);
and U35001 (N_35001,N_33673,N_33534);
xnor U35002 (N_35002,N_33150,N_32368);
xnor U35003 (N_35003,N_33383,N_32407);
or U35004 (N_35004,N_33292,N_33181);
nor U35005 (N_35005,N_32982,N_33646);
xor U35006 (N_35006,N_33355,N_32589);
xor U35007 (N_35007,N_32049,N_33038);
nor U35008 (N_35008,N_32060,N_32018);
or U35009 (N_35009,N_33743,N_33734);
or U35010 (N_35010,N_32246,N_33827);
and U35011 (N_35011,N_33780,N_32259);
or U35012 (N_35012,N_32964,N_32081);
nor U35013 (N_35013,N_33503,N_33459);
and U35014 (N_35014,N_32799,N_32316);
nand U35015 (N_35015,N_33027,N_33826);
xnor U35016 (N_35016,N_33452,N_33027);
nor U35017 (N_35017,N_32844,N_32610);
and U35018 (N_35018,N_33738,N_32812);
nor U35019 (N_35019,N_33553,N_32697);
nor U35020 (N_35020,N_33369,N_33868);
and U35021 (N_35021,N_33950,N_33797);
or U35022 (N_35022,N_32307,N_32576);
or U35023 (N_35023,N_32111,N_33546);
nand U35024 (N_35024,N_32058,N_32506);
nor U35025 (N_35025,N_32837,N_33994);
or U35026 (N_35026,N_32036,N_32367);
xnor U35027 (N_35027,N_32781,N_33234);
and U35028 (N_35028,N_33700,N_32398);
nor U35029 (N_35029,N_33406,N_33024);
nor U35030 (N_35030,N_33970,N_33184);
nand U35031 (N_35031,N_33504,N_33494);
nor U35032 (N_35032,N_33081,N_33484);
nor U35033 (N_35033,N_32992,N_32753);
nand U35034 (N_35034,N_33872,N_33338);
or U35035 (N_35035,N_33176,N_33088);
and U35036 (N_35036,N_33757,N_32182);
nand U35037 (N_35037,N_32723,N_32048);
nor U35038 (N_35038,N_32955,N_32455);
and U35039 (N_35039,N_33610,N_33111);
nand U35040 (N_35040,N_32653,N_33364);
xnor U35041 (N_35041,N_33251,N_33410);
and U35042 (N_35042,N_32060,N_33988);
nor U35043 (N_35043,N_32779,N_33209);
and U35044 (N_35044,N_32031,N_33945);
nor U35045 (N_35045,N_33790,N_32705);
nand U35046 (N_35046,N_33483,N_33953);
nor U35047 (N_35047,N_33398,N_32953);
xnor U35048 (N_35048,N_33662,N_32507);
or U35049 (N_35049,N_33550,N_33575);
nand U35050 (N_35050,N_33080,N_32798);
xnor U35051 (N_35051,N_32874,N_32929);
nor U35052 (N_35052,N_33688,N_32600);
and U35053 (N_35053,N_33764,N_32648);
or U35054 (N_35054,N_32809,N_32337);
or U35055 (N_35055,N_32831,N_33148);
nand U35056 (N_35056,N_32015,N_33779);
nand U35057 (N_35057,N_32491,N_32442);
nor U35058 (N_35058,N_33358,N_32231);
or U35059 (N_35059,N_32504,N_32491);
and U35060 (N_35060,N_33164,N_33271);
or U35061 (N_35061,N_32583,N_33219);
or U35062 (N_35062,N_32127,N_32999);
nand U35063 (N_35063,N_33045,N_33560);
or U35064 (N_35064,N_32965,N_33297);
xnor U35065 (N_35065,N_33862,N_33760);
nor U35066 (N_35066,N_33056,N_33505);
nand U35067 (N_35067,N_33414,N_32428);
nand U35068 (N_35068,N_33770,N_32750);
nor U35069 (N_35069,N_32758,N_33474);
nor U35070 (N_35070,N_33226,N_33719);
nand U35071 (N_35071,N_33248,N_32997);
and U35072 (N_35072,N_33622,N_32848);
nor U35073 (N_35073,N_33196,N_32556);
or U35074 (N_35074,N_33605,N_32895);
or U35075 (N_35075,N_33979,N_32050);
xor U35076 (N_35076,N_32474,N_32087);
or U35077 (N_35077,N_33157,N_32044);
and U35078 (N_35078,N_32465,N_32624);
xor U35079 (N_35079,N_32962,N_32978);
xnor U35080 (N_35080,N_33668,N_33792);
nand U35081 (N_35081,N_33644,N_33766);
nand U35082 (N_35082,N_32991,N_33463);
or U35083 (N_35083,N_33595,N_33918);
or U35084 (N_35084,N_32807,N_33653);
and U35085 (N_35085,N_32125,N_32486);
or U35086 (N_35086,N_32492,N_33657);
and U35087 (N_35087,N_33584,N_33882);
nor U35088 (N_35088,N_33522,N_32098);
xor U35089 (N_35089,N_32925,N_33212);
xor U35090 (N_35090,N_32206,N_33036);
nand U35091 (N_35091,N_33864,N_33637);
nand U35092 (N_35092,N_32472,N_32430);
xnor U35093 (N_35093,N_33349,N_33132);
or U35094 (N_35094,N_33302,N_33411);
or U35095 (N_35095,N_33838,N_32902);
nand U35096 (N_35096,N_33277,N_33621);
or U35097 (N_35097,N_32187,N_32113);
and U35098 (N_35098,N_33691,N_32768);
xor U35099 (N_35099,N_32578,N_33346);
and U35100 (N_35100,N_32406,N_32474);
xor U35101 (N_35101,N_32406,N_32916);
and U35102 (N_35102,N_33117,N_32322);
and U35103 (N_35103,N_32331,N_32492);
xor U35104 (N_35104,N_33364,N_33120);
nor U35105 (N_35105,N_33703,N_32164);
and U35106 (N_35106,N_32103,N_33874);
or U35107 (N_35107,N_33407,N_33526);
nor U35108 (N_35108,N_32864,N_32914);
or U35109 (N_35109,N_33082,N_32464);
nor U35110 (N_35110,N_33648,N_33902);
or U35111 (N_35111,N_33441,N_32898);
and U35112 (N_35112,N_33884,N_32151);
xor U35113 (N_35113,N_32947,N_33115);
nand U35114 (N_35114,N_32831,N_32712);
or U35115 (N_35115,N_32101,N_33522);
nand U35116 (N_35116,N_32139,N_32704);
xnor U35117 (N_35117,N_32630,N_32195);
and U35118 (N_35118,N_32978,N_32731);
nand U35119 (N_35119,N_32112,N_33230);
xor U35120 (N_35120,N_33280,N_32329);
xor U35121 (N_35121,N_32247,N_32157);
or U35122 (N_35122,N_33422,N_32587);
xor U35123 (N_35123,N_32507,N_33793);
xnor U35124 (N_35124,N_33345,N_32974);
nand U35125 (N_35125,N_33685,N_33668);
xnor U35126 (N_35126,N_33731,N_32303);
and U35127 (N_35127,N_32818,N_32085);
nand U35128 (N_35128,N_33625,N_32840);
xor U35129 (N_35129,N_32941,N_32220);
or U35130 (N_35130,N_32980,N_32472);
nand U35131 (N_35131,N_32264,N_32435);
and U35132 (N_35132,N_33568,N_33562);
nand U35133 (N_35133,N_33197,N_32504);
xnor U35134 (N_35134,N_32637,N_32626);
and U35135 (N_35135,N_33796,N_33561);
and U35136 (N_35136,N_33152,N_32667);
and U35137 (N_35137,N_33173,N_32648);
or U35138 (N_35138,N_32405,N_33346);
and U35139 (N_35139,N_32663,N_33410);
or U35140 (N_35140,N_33798,N_33189);
and U35141 (N_35141,N_32105,N_33965);
and U35142 (N_35142,N_32479,N_33683);
xnor U35143 (N_35143,N_32607,N_33200);
or U35144 (N_35144,N_33010,N_32945);
nand U35145 (N_35145,N_32893,N_32163);
or U35146 (N_35146,N_32969,N_32265);
nor U35147 (N_35147,N_32580,N_32318);
nor U35148 (N_35148,N_32997,N_32747);
nand U35149 (N_35149,N_32667,N_33529);
nand U35150 (N_35150,N_32147,N_32821);
xnor U35151 (N_35151,N_32573,N_32034);
xor U35152 (N_35152,N_33996,N_32032);
nor U35153 (N_35153,N_33329,N_32455);
nand U35154 (N_35154,N_33989,N_33319);
nand U35155 (N_35155,N_32925,N_32007);
nor U35156 (N_35156,N_32226,N_32119);
nand U35157 (N_35157,N_32779,N_33253);
nor U35158 (N_35158,N_33303,N_32155);
nand U35159 (N_35159,N_32124,N_33108);
and U35160 (N_35160,N_32730,N_33535);
and U35161 (N_35161,N_32679,N_32583);
xor U35162 (N_35162,N_32454,N_33926);
nor U35163 (N_35163,N_32529,N_32090);
nand U35164 (N_35164,N_32545,N_33036);
nor U35165 (N_35165,N_33358,N_33798);
nor U35166 (N_35166,N_33751,N_32453);
nand U35167 (N_35167,N_32709,N_32305);
or U35168 (N_35168,N_32206,N_33326);
or U35169 (N_35169,N_32442,N_32235);
nor U35170 (N_35170,N_32511,N_33889);
and U35171 (N_35171,N_32995,N_33447);
xnor U35172 (N_35172,N_33517,N_33169);
nand U35173 (N_35173,N_33919,N_33292);
nor U35174 (N_35174,N_33018,N_33612);
xor U35175 (N_35175,N_33910,N_33618);
nand U35176 (N_35176,N_32300,N_33114);
and U35177 (N_35177,N_33553,N_33426);
nand U35178 (N_35178,N_32525,N_33334);
xor U35179 (N_35179,N_33737,N_33547);
or U35180 (N_35180,N_33534,N_32307);
nand U35181 (N_35181,N_33419,N_33048);
and U35182 (N_35182,N_32009,N_33672);
and U35183 (N_35183,N_33095,N_33500);
nor U35184 (N_35184,N_32663,N_32757);
nor U35185 (N_35185,N_32679,N_33358);
or U35186 (N_35186,N_33778,N_33566);
and U35187 (N_35187,N_32905,N_32586);
nor U35188 (N_35188,N_33298,N_32311);
or U35189 (N_35189,N_32073,N_33508);
or U35190 (N_35190,N_33470,N_32580);
nor U35191 (N_35191,N_32439,N_32922);
xnor U35192 (N_35192,N_33227,N_33287);
or U35193 (N_35193,N_32713,N_32177);
xor U35194 (N_35194,N_32869,N_32447);
nor U35195 (N_35195,N_33011,N_33165);
nand U35196 (N_35196,N_33020,N_32062);
nor U35197 (N_35197,N_32948,N_33153);
xnor U35198 (N_35198,N_33267,N_32125);
xnor U35199 (N_35199,N_33571,N_33582);
nand U35200 (N_35200,N_32933,N_32425);
xnor U35201 (N_35201,N_32113,N_32641);
and U35202 (N_35202,N_33488,N_33973);
nand U35203 (N_35203,N_32038,N_32697);
or U35204 (N_35204,N_33861,N_32146);
xor U35205 (N_35205,N_32257,N_32576);
xnor U35206 (N_35206,N_32599,N_33211);
and U35207 (N_35207,N_33966,N_32000);
nand U35208 (N_35208,N_33816,N_33829);
xnor U35209 (N_35209,N_33286,N_33317);
xnor U35210 (N_35210,N_33296,N_33175);
or U35211 (N_35211,N_32136,N_32889);
or U35212 (N_35212,N_32814,N_32089);
or U35213 (N_35213,N_33256,N_33036);
and U35214 (N_35214,N_32013,N_32885);
or U35215 (N_35215,N_33074,N_32738);
nand U35216 (N_35216,N_33251,N_32742);
nor U35217 (N_35217,N_32414,N_33332);
xor U35218 (N_35218,N_33257,N_32564);
and U35219 (N_35219,N_32058,N_32921);
or U35220 (N_35220,N_32954,N_32754);
and U35221 (N_35221,N_33848,N_32907);
and U35222 (N_35222,N_32880,N_32777);
or U35223 (N_35223,N_32549,N_32145);
nand U35224 (N_35224,N_33816,N_32302);
xor U35225 (N_35225,N_33700,N_32751);
and U35226 (N_35226,N_32136,N_32981);
or U35227 (N_35227,N_33068,N_32850);
nand U35228 (N_35228,N_32666,N_33604);
and U35229 (N_35229,N_33458,N_33649);
or U35230 (N_35230,N_33573,N_33417);
nand U35231 (N_35231,N_33834,N_33523);
or U35232 (N_35232,N_32028,N_32189);
and U35233 (N_35233,N_33428,N_32710);
nand U35234 (N_35234,N_32025,N_32443);
and U35235 (N_35235,N_32618,N_32274);
nor U35236 (N_35236,N_33614,N_32633);
nor U35237 (N_35237,N_32483,N_33738);
xnor U35238 (N_35238,N_33407,N_33776);
or U35239 (N_35239,N_33703,N_32778);
and U35240 (N_35240,N_32892,N_32978);
and U35241 (N_35241,N_32919,N_32894);
nand U35242 (N_35242,N_33033,N_33565);
nor U35243 (N_35243,N_32117,N_32409);
nor U35244 (N_35244,N_32703,N_32169);
and U35245 (N_35245,N_32095,N_33529);
or U35246 (N_35246,N_33199,N_33781);
nand U35247 (N_35247,N_33945,N_33349);
or U35248 (N_35248,N_32049,N_32945);
nand U35249 (N_35249,N_33592,N_33387);
nand U35250 (N_35250,N_32565,N_33520);
nor U35251 (N_35251,N_33732,N_33431);
xor U35252 (N_35252,N_33963,N_33765);
xor U35253 (N_35253,N_32266,N_32683);
nand U35254 (N_35254,N_33746,N_32433);
or U35255 (N_35255,N_33452,N_32929);
xnor U35256 (N_35256,N_32149,N_32315);
or U35257 (N_35257,N_32990,N_32625);
nand U35258 (N_35258,N_32524,N_32037);
and U35259 (N_35259,N_32128,N_33300);
and U35260 (N_35260,N_32767,N_33869);
xnor U35261 (N_35261,N_32662,N_33041);
xnor U35262 (N_35262,N_32630,N_33357);
nand U35263 (N_35263,N_32322,N_32398);
xor U35264 (N_35264,N_33511,N_33167);
or U35265 (N_35265,N_32933,N_32946);
nand U35266 (N_35266,N_32372,N_32123);
nor U35267 (N_35267,N_33764,N_33067);
xor U35268 (N_35268,N_33379,N_32221);
nor U35269 (N_35269,N_33093,N_33723);
nor U35270 (N_35270,N_32178,N_32008);
and U35271 (N_35271,N_32896,N_33257);
nand U35272 (N_35272,N_33345,N_33281);
nor U35273 (N_35273,N_32809,N_33079);
nor U35274 (N_35274,N_33898,N_33378);
or U35275 (N_35275,N_33892,N_32755);
or U35276 (N_35276,N_33995,N_32679);
or U35277 (N_35277,N_33547,N_33972);
and U35278 (N_35278,N_33534,N_33480);
nor U35279 (N_35279,N_33513,N_32497);
nand U35280 (N_35280,N_33870,N_32054);
xor U35281 (N_35281,N_32674,N_32089);
nand U35282 (N_35282,N_33723,N_33980);
nor U35283 (N_35283,N_33009,N_32180);
or U35284 (N_35284,N_32419,N_32588);
nor U35285 (N_35285,N_32748,N_33858);
or U35286 (N_35286,N_33880,N_32026);
and U35287 (N_35287,N_32392,N_32002);
xnor U35288 (N_35288,N_32594,N_32134);
and U35289 (N_35289,N_33530,N_32131);
nand U35290 (N_35290,N_32001,N_32086);
nor U35291 (N_35291,N_32561,N_33371);
or U35292 (N_35292,N_32095,N_32041);
and U35293 (N_35293,N_33241,N_32747);
and U35294 (N_35294,N_33320,N_33443);
nand U35295 (N_35295,N_32412,N_32021);
or U35296 (N_35296,N_33912,N_33557);
nor U35297 (N_35297,N_32268,N_32508);
xnor U35298 (N_35298,N_33672,N_32073);
nor U35299 (N_35299,N_33768,N_32694);
and U35300 (N_35300,N_32681,N_32468);
and U35301 (N_35301,N_33876,N_33416);
nand U35302 (N_35302,N_32567,N_32882);
and U35303 (N_35303,N_32621,N_32019);
and U35304 (N_35304,N_33757,N_32379);
and U35305 (N_35305,N_33057,N_32371);
xnor U35306 (N_35306,N_32484,N_33670);
nor U35307 (N_35307,N_32988,N_32014);
or U35308 (N_35308,N_33108,N_32349);
xor U35309 (N_35309,N_32534,N_33473);
xor U35310 (N_35310,N_33801,N_32148);
nand U35311 (N_35311,N_33146,N_33594);
nor U35312 (N_35312,N_32741,N_33628);
nor U35313 (N_35313,N_33772,N_33275);
and U35314 (N_35314,N_33292,N_33366);
and U35315 (N_35315,N_32299,N_33353);
and U35316 (N_35316,N_32314,N_32940);
xnor U35317 (N_35317,N_33865,N_32197);
nor U35318 (N_35318,N_33044,N_32033);
xnor U35319 (N_35319,N_33944,N_32513);
xnor U35320 (N_35320,N_33473,N_32515);
or U35321 (N_35321,N_33817,N_33845);
nor U35322 (N_35322,N_33363,N_33817);
and U35323 (N_35323,N_33254,N_32454);
xnor U35324 (N_35324,N_32279,N_32444);
nor U35325 (N_35325,N_32216,N_33565);
nand U35326 (N_35326,N_32216,N_33291);
and U35327 (N_35327,N_33624,N_33083);
nor U35328 (N_35328,N_32007,N_32231);
and U35329 (N_35329,N_33057,N_33203);
nand U35330 (N_35330,N_32843,N_33356);
or U35331 (N_35331,N_32559,N_33815);
nor U35332 (N_35332,N_33148,N_33720);
and U35333 (N_35333,N_32594,N_32998);
xnor U35334 (N_35334,N_33086,N_32609);
or U35335 (N_35335,N_33607,N_33224);
nand U35336 (N_35336,N_33825,N_33979);
or U35337 (N_35337,N_32350,N_33889);
nor U35338 (N_35338,N_32715,N_33751);
xor U35339 (N_35339,N_33652,N_33585);
xnor U35340 (N_35340,N_33812,N_32247);
xor U35341 (N_35341,N_32272,N_32764);
nor U35342 (N_35342,N_32728,N_32092);
and U35343 (N_35343,N_32492,N_32478);
nand U35344 (N_35344,N_33946,N_33291);
and U35345 (N_35345,N_33833,N_32054);
nand U35346 (N_35346,N_33769,N_33727);
and U35347 (N_35347,N_32944,N_32634);
nand U35348 (N_35348,N_32660,N_32286);
nand U35349 (N_35349,N_32684,N_32401);
nand U35350 (N_35350,N_33463,N_32033);
or U35351 (N_35351,N_33780,N_32102);
nor U35352 (N_35352,N_33873,N_33818);
xor U35353 (N_35353,N_32392,N_33008);
xnor U35354 (N_35354,N_32976,N_33353);
nand U35355 (N_35355,N_32285,N_33020);
xor U35356 (N_35356,N_32337,N_32724);
nand U35357 (N_35357,N_32622,N_32096);
xnor U35358 (N_35358,N_32798,N_32181);
or U35359 (N_35359,N_33402,N_32870);
nand U35360 (N_35360,N_32439,N_32499);
and U35361 (N_35361,N_32638,N_33439);
or U35362 (N_35362,N_32591,N_32537);
nor U35363 (N_35363,N_33859,N_32210);
nand U35364 (N_35364,N_33131,N_32616);
and U35365 (N_35365,N_33819,N_32780);
and U35366 (N_35366,N_33450,N_32870);
nand U35367 (N_35367,N_33869,N_33334);
nand U35368 (N_35368,N_32637,N_32912);
nand U35369 (N_35369,N_32416,N_32424);
and U35370 (N_35370,N_33885,N_32345);
nand U35371 (N_35371,N_32562,N_33946);
and U35372 (N_35372,N_33582,N_32220);
nand U35373 (N_35373,N_33304,N_32872);
and U35374 (N_35374,N_32676,N_32352);
or U35375 (N_35375,N_32752,N_33259);
or U35376 (N_35376,N_33195,N_33664);
xnor U35377 (N_35377,N_32049,N_32157);
nor U35378 (N_35378,N_33536,N_33153);
nand U35379 (N_35379,N_33916,N_33776);
nand U35380 (N_35380,N_32535,N_33654);
nor U35381 (N_35381,N_33111,N_32366);
nor U35382 (N_35382,N_33090,N_33027);
or U35383 (N_35383,N_32692,N_32082);
and U35384 (N_35384,N_33650,N_33426);
and U35385 (N_35385,N_32646,N_33204);
nor U35386 (N_35386,N_32071,N_32283);
nand U35387 (N_35387,N_33090,N_32225);
xor U35388 (N_35388,N_33801,N_33346);
nand U35389 (N_35389,N_32547,N_33484);
and U35390 (N_35390,N_32894,N_32860);
nor U35391 (N_35391,N_33664,N_33341);
nor U35392 (N_35392,N_32237,N_32093);
and U35393 (N_35393,N_32772,N_33263);
or U35394 (N_35394,N_32261,N_32783);
xnor U35395 (N_35395,N_32673,N_33892);
nand U35396 (N_35396,N_32006,N_33920);
and U35397 (N_35397,N_33087,N_32676);
xor U35398 (N_35398,N_33493,N_33661);
nand U35399 (N_35399,N_32690,N_33792);
nand U35400 (N_35400,N_33972,N_33863);
and U35401 (N_35401,N_32835,N_32715);
nand U35402 (N_35402,N_33425,N_32584);
xor U35403 (N_35403,N_33263,N_33606);
xor U35404 (N_35404,N_32246,N_33251);
nor U35405 (N_35405,N_32301,N_32555);
nand U35406 (N_35406,N_33166,N_32669);
nand U35407 (N_35407,N_33266,N_32075);
and U35408 (N_35408,N_33790,N_32006);
nand U35409 (N_35409,N_33179,N_32097);
nor U35410 (N_35410,N_33861,N_33485);
xnor U35411 (N_35411,N_33966,N_33155);
xor U35412 (N_35412,N_32563,N_33310);
nor U35413 (N_35413,N_32630,N_33761);
xor U35414 (N_35414,N_33592,N_33085);
xor U35415 (N_35415,N_32495,N_33195);
nand U35416 (N_35416,N_33477,N_33280);
and U35417 (N_35417,N_32241,N_33162);
nand U35418 (N_35418,N_33148,N_32829);
nor U35419 (N_35419,N_32422,N_32652);
or U35420 (N_35420,N_33725,N_33409);
or U35421 (N_35421,N_32584,N_32038);
nor U35422 (N_35422,N_32138,N_32023);
nand U35423 (N_35423,N_32984,N_32337);
and U35424 (N_35424,N_32559,N_32749);
xor U35425 (N_35425,N_33348,N_32727);
and U35426 (N_35426,N_32212,N_33804);
xnor U35427 (N_35427,N_33017,N_32830);
or U35428 (N_35428,N_32582,N_32123);
xor U35429 (N_35429,N_32021,N_32294);
xor U35430 (N_35430,N_32654,N_32737);
nand U35431 (N_35431,N_33664,N_32607);
nor U35432 (N_35432,N_33923,N_33983);
nand U35433 (N_35433,N_33952,N_32081);
xnor U35434 (N_35434,N_33701,N_32551);
and U35435 (N_35435,N_32650,N_33211);
or U35436 (N_35436,N_32044,N_33093);
nand U35437 (N_35437,N_32820,N_32652);
xor U35438 (N_35438,N_33629,N_32648);
nor U35439 (N_35439,N_32190,N_32513);
nand U35440 (N_35440,N_32563,N_33141);
or U35441 (N_35441,N_33937,N_33578);
nand U35442 (N_35442,N_33510,N_32842);
xor U35443 (N_35443,N_33565,N_33104);
nor U35444 (N_35444,N_33673,N_33628);
and U35445 (N_35445,N_33648,N_32318);
nor U35446 (N_35446,N_33523,N_32084);
nor U35447 (N_35447,N_32931,N_32438);
nand U35448 (N_35448,N_33768,N_33621);
xor U35449 (N_35449,N_32452,N_32949);
or U35450 (N_35450,N_32853,N_33575);
xor U35451 (N_35451,N_33257,N_33928);
xnor U35452 (N_35452,N_33921,N_33395);
or U35453 (N_35453,N_33231,N_33558);
xnor U35454 (N_35454,N_32243,N_33140);
xnor U35455 (N_35455,N_33104,N_32850);
nor U35456 (N_35456,N_32720,N_32116);
xor U35457 (N_35457,N_32156,N_32756);
nand U35458 (N_35458,N_33838,N_32471);
and U35459 (N_35459,N_33618,N_33357);
xor U35460 (N_35460,N_33596,N_32302);
nor U35461 (N_35461,N_33064,N_33188);
nand U35462 (N_35462,N_33385,N_32534);
or U35463 (N_35463,N_32507,N_32957);
nor U35464 (N_35464,N_33967,N_33074);
nor U35465 (N_35465,N_32782,N_32280);
nor U35466 (N_35466,N_33265,N_32188);
nand U35467 (N_35467,N_33754,N_32253);
and U35468 (N_35468,N_32278,N_32607);
xor U35469 (N_35469,N_32411,N_33888);
nor U35470 (N_35470,N_33705,N_32899);
or U35471 (N_35471,N_33531,N_32694);
nor U35472 (N_35472,N_33522,N_32506);
and U35473 (N_35473,N_33859,N_32031);
xor U35474 (N_35474,N_33179,N_32120);
xor U35475 (N_35475,N_32012,N_33902);
nor U35476 (N_35476,N_32183,N_32198);
nand U35477 (N_35477,N_33297,N_32977);
nor U35478 (N_35478,N_32126,N_33565);
xnor U35479 (N_35479,N_33764,N_33505);
or U35480 (N_35480,N_33293,N_33344);
and U35481 (N_35481,N_32203,N_32133);
and U35482 (N_35482,N_33751,N_33449);
xnor U35483 (N_35483,N_33360,N_32196);
or U35484 (N_35484,N_33352,N_33929);
and U35485 (N_35485,N_32257,N_33855);
or U35486 (N_35486,N_33288,N_32066);
nor U35487 (N_35487,N_32430,N_32450);
and U35488 (N_35488,N_32187,N_33055);
xnor U35489 (N_35489,N_32986,N_32282);
nand U35490 (N_35490,N_33165,N_33778);
and U35491 (N_35491,N_33019,N_33808);
nand U35492 (N_35492,N_32288,N_33471);
xor U35493 (N_35493,N_33876,N_32029);
nand U35494 (N_35494,N_32458,N_32557);
xnor U35495 (N_35495,N_32247,N_33765);
nor U35496 (N_35496,N_32851,N_32587);
and U35497 (N_35497,N_32128,N_33036);
or U35498 (N_35498,N_32592,N_32067);
or U35499 (N_35499,N_33881,N_32391);
or U35500 (N_35500,N_32397,N_33700);
xor U35501 (N_35501,N_33176,N_33653);
and U35502 (N_35502,N_33627,N_33781);
or U35503 (N_35503,N_32640,N_32429);
or U35504 (N_35504,N_32405,N_32233);
nor U35505 (N_35505,N_33850,N_33023);
or U35506 (N_35506,N_32883,N_33659);
or U35507 (N_35507,N_33470,N_33629);
nand U35508 (N_35508,N_33061,N_33146);
or U35509 (N_35509,N_33571,N_33728);
nand U35510 (N_35510,N_32792,N_32666);
or U35511 (N_35511,N_32551,N_33822);
xor U35512 (N_35512,N_33261,N_33398);
nor U35513 (N_35513,N_33299,N_33325);
and U35514 (N_35514,N_33580,N_32038);
xnor U35515 (N_35515,N_32304,N_33431);
nand U35516 (N_35516,N_33309,N_33931);
or U35517 (N_35517,N_33998,N_32658);
xor U35518 (N_35518,N_33897,N_33506);
nand U35519 (N_35519,N_33615,N_32808);
xor U35520 (N_35520,N_33650,N_33068);
nand U35521 (N_35521,N_32415,N_32476);
and U35522 (N_35522,N_33970,N_33131);
or U35523 (N_35523,N_33028,N_32353);
xor U35524 (N_35524,N_33780,N_32055);
nand U35525 (N_35525,N_33410,N_32150);
xor U35526 (N_35526,N_33592,N_32970);
xnor U35527 (N_35527,N_33668,N_32039);
nand U35528 (N_35528,N_32018,N_33756);
and U35529 (N_35529,N_33792,N_32397);
xor U35530 (N_35530,N_32902,N_32921);
xor U35531 (N_35531,N_33476,N_33458);
or U35532 (N_35532,N_32082,N_32166);
or U35533 (N_35533,N_33717,N_33251);
nor U35534 (N_35534,N_33290,N_32120);
or U35535 (N_35535,N_32718,N_33983);
nand U35536 (N_35536,N_32520,N_32005);
nand U35537 (N_35537,N_32799,N_32004);
and U35538 (N_35538,N_32077,N_33065);
nor U35539 (N_35539,N_32652,N_32734);
or U35540 (N_35540,N_33762,N_32772);
nor U35541 (N_35541,N_32572,N_33870);
nor U35542 (N_35542,N_32298,N_33324);
nor U35543 (N_35543,N_33437,N_33655);
xor U35544 (N_35544,N_33475,N_32423);
and U35545 (N_35545,N_32567,N_33122);
xor U35546 (N_35546,N_33212,N_33069);
nand U35547 (N_35547,N_32972,N_33971);
and U35548 (N_35548,N_33952,N_33261);
or U35549 (N_35549,N_32522,N_32489);
and U35550 (N_35550,N_33661,N_33272);
nor U35551 (N_35551,N_32470,N_32349);
or U35552 (N_35552,N_33838,N_32456);
nand U35553 (N_35553,N_33702,N_33027);
and U35554 (N_35554,N_33506,N_32393);
xor U35555 (N_35555,N_32971,N_32007);
and U35556 (N_35556,N_32344,N_33192);
xnor U35557 (N_35557,N_32939,N_32766);
and U35558 (N_35558,N_32083,N_33222);
and U35559 (N_35559,N_33252,N_33888);
xnor U35560 (N_35560,N_33484,N_32629);
nand U35561 (N_35561,N_32024,N_33453);
nand U35562 (N_35562,N_32154,N_33889);
xor U35563 (N_35563,N_33892,N_33198);
or U35564 (N_35564,N_32791,N_32459);
nand U35565 (N_35565,N_32880,N_33156);
nand U35566 (N_35566,N_33258,N_32076);
or U35567 (N_35567,N_32580,N_33433);
and U35568 (N_35568,N_32126,N_32759);
and U35569 (N_35569,N_32845,N_32712);
or U35570 (N_35570,N_32739,N_32514);
and U35571 (N_35571,N_33917,N_32426);
nor U35572 (N_35572,N_32368,N_32159);
and U35573 (N_35573,N_32391,N_32953);
nor U35574 (N_35574,N_33063,N_33839);
or U35575 (N_35575,N_33786,N_33173);
xor U35576 (N_35576,N_32560,N_33702);
nand U35577 (N_35577,N_32553,N_33690);
or U35578 (N_35578,N_32952,N_33463);
or U35579 (N_35579,N_32376,N_32836);
nor U35580 (N_35580,N_33603,N_32465);
xnor U35581 (N_35581,N_33727,N_32209);
xor U35582 (N_35582,N_33302,N_32573);
or U35583 (N_35583,N_33302,N_32096);
nand U35584 (N_35584,N_32624,N_33342);
or U35585 (N_35585,N_33513,N_33087);
and U35586 (N_35586,N_32092,N_32633);
nand U35587 (N_35587,N_33957,N_32849);
nand U35588 (N_35588,N_32948,N_33140);
xor U35589 (N_35589,N_33469,N_32185);
or U35590 (N_35590,N_32526,N_32351);
or U35591 (N_35591,N_33783,N_33445);
or U35592 (N_35592,N_33504,N_33833);
or U35593 (N_35593,N_33917,N_33655);
nand U35594 (N_35594,N_33308,N_32099);
or U35595 (N_35595,N_32801,N_32023);
nor U35596 (N_35596,N_32413,N_32906);
xor U35597 (N_35597,N_33363,N_32305);
nand U35598 (N_35598,N_33623,N_32144);
and U35599 (N_35599,N_33555,N_33346);
and U35600 (N_35600,N_33022,N_32855);
xor U35601 (N_35601,N_33050,N_33566);
and U35602 (N_35602,N_33389,N_33916);
and U35603 (N_35603,N_33004,N_32249);
xnor U35604 (N_35604,N_32042,N_33050);
or U35605 (N_35605,N_33382,N_33247);
and U35606 (N_35606,N_32965,N_33876);
and U35607 (N_35607,N_32559,N_33870);
xnor U35608 (N_35608,N_32412,N_33867);
xnor U35609 (N_35609,N_33134,N_33522);
or U35610 (N_35610,N_33957,N_33897);
xnor U35611 (N_35611,N_33159,N_32537);
nand U35612 (N_35612,N_33474,N_33239);
nor U35613 (N_35613,N_33991,N_32043);
or U35614 (N_35614,N_32704,N_33572);
nand U35615 (N_35615,N_32157,N_33194);
and U35616 (N_35616,N_32436,N_33645);
or U35617 (N_35617,N_32450,N_33153);
nor U35618 (N_35618,N_33770,N_33000);
nand U35619 (N_35619,N_32749,N_33607);
xor U35620 (N_35620,N_33800,N_33730);
or U35621 (N_35621,N_32936,N_32255);
xor U35622 (N_35622,N_33934,N_33566);
nor U35623 (N_35623,N_32715,N_32498);
nor U35624 (N_35624,N_32531,N_32994);
or U35625 (N_35625,N_32674,N_32169);
xnor U35626 (N_35626,N_33255,N_33508);
nand U35627 (N_35627,N_33686,N_33273);
or U35628 (N_35628,N_33963,N_33067);
nand U35629 (N_35629,N_33669,N_32680);
or U35630 (N_35630,N_33274,N_33698);
nor U35631 (N_35631,N_32489,N_33293);
nand U35632 (N_35632,N_33237,N_32185);
xnor U35633 (N_35633,N_33665,N_33790);
or U35634 (N_35634,N_33906,N_33193);
nor U35635 (N_35635,N_33774,N_33473);
or U35636 (N_35636,N_33559,N_32924);
nand U35637 (N_35637,N_32082,N_33338);
nand U35638 (N_35638,N_32259,N_32198);
xnor U35639 (N_35639,N_32819,N_32128);
nand U35640 (N_35640,N_33087,N_33163);
xnor U35641 (N_35641,N_32675,N_33608);
and U35642 (N_35642,N_33212,N_32870);
nor U35643 (N_35643,N_32253,N_32873);
or U35644 (N_35644,N_32272,N_32963);
xor U35645 (N_35645,N_33379,N_33622);
xnor U35646 (N_35646,N_33554,N_33055);
nor U35647 (N_35647,N_32487,N_33724);
and U35648 (N_35648,N_33891,N_33016);
nor U35649 (N_35649,N_33229,N_32569);
nor U35650 (N_35650,N_33882,N_32693);
and U35651 (N_35651,N_32385,N_33437);
and U35652 (N_35652,N_33692,N_33753);
xor U35653 (N_35653,N_33773,N_33173);
nor U35654 (N_35654,N_32440,N_33367);
and U35655 (N_35655,N_32384,N_33578);
or U35656 (N_35656,N_32310,N_33555);
nand U35657 (N_35657,N_32238,N_33193);
xnor U35658 (N_35658,N_32821,N_32134);
nand U35659 (N_35659,N_32794,N_33805);
or U35660 (N_35660,N_33129,N_32463);
nor U35661 (N_35661,N_32546,N_33728);
or U35662 (N_35662,N_32587,N_33359);
or U35663 (N_35663,N_32720,N_33023);
nand U35664 (N_35664,N_33622,N_33657);
xnor U35665 (N_35665,N_32245,N_33070);
nor U35666 (N_35666,N_32818,N_32991);
and U35667 (N_35667,N_33544,N_32859);
xnor U35668 (N_35668,N_32293,N_33328);
xor U35669 (N_35669,N_33252,N_32075);
and U35670 (N_35670,N_32056,N_33255);
and U35671 (N_35671,N_32119,N_32342);
xor U35672 (N_35672,N_32033,N_33517);
xor U35673 (N_35673,N_32920,N_32524);
nor U35674 (N_35674,N_32358,N_33201);
nor U35675 (N_35675,N_33937,N_33859);
xnor U35676 (N_35676,N_33136,N_33751);
xor U35677 (N_35677,N_33449,N_33951);
and U35678 (N_35678,N_33394,N_33420);
or U35679 (N_35679,N_33081,N_33634);
and U35680 (N_35680,N_32277,N_32533);
nand U35681 (N_35681,N_33546,N_32647);
nor U35682 (N_35682,N_33172,N_32698);
or U35683 (N_35683,N_33665,N_33050);
xnor U35684 (N_35684,N_33536,N_32766);
xor U35685 (N_35685,N_32588,N_32848);
nand U35686 (N_35686,N_32299,N_32507);
and U35687 (N_35687,N_33862,N_33813);
nor U35688 (N_35688,N_33555,N_33470);
nor U35689 (N_35689,N_32322,N_32164);
and U35690 (N_35690,N_33190,N_32499);
xnor U35691 (N_35691,N_33285,N_33378);
nand U35692 (N_35692,N_32835,N_32736);
or U35693 (N_35693,N_32590,N_33986);
or U35694 (N_35694,N_33342,N_32191);
or U35695 (N_35695,N_32448,N_32820);
nand U35696 (N_35696,N_33128,N_33073);
or U35697 (N_35697,N_33432,N_33854);
or U35698 (N_35698,N_33226,N_33567);
or U35699 (N_35699,N_32872,N_33262);
nand U35700 (N_35700,N_33075,N_32288);
nor U35701 (N_35701,N_32827,N_33708);
and U35702 (N_35702,N_33366,N_32233);
nand U35703 (N_35703,N_32948,N_33711);
or U35704 (N_35704,N_33283,N_33227);
xnor U35705 (N_35705,N_32033,N_32455);
nor U35706 (N_35706,N_32261,N_32831);
nand U35707 (N_35707,N_33937,N_32983);
xnor U35708 (N_35708,N_32469,N_32622);
nand U35709 (N_35709,N_32852,N_33199);
nor U35710 (N_35710,N_32364,N_32358);
xnor U35711 (N_35711,N_32583,N_32639);
nor U35712 (N_35712,N_32151,N_33685);
nand U35713 (N_35713,N_33622,N_33790);
xor U35714 (N_35714,N_32086,N_33969);
xnor U35715 (N_35715,N_32010,N_33658);
or U35716 (N_35716,N_32877,N_32730);
nor U35717 (N_35717,N_32363,N_33006);
nand U35718 (N_35718,N_32368,N_33066);
nand U35719 (N_35719,N_33894,N_33595);
xnor U35720 (N_35720,N_33199,N_33684);
nor U35721 (N_35721,N_32721,N_32114);
nand U35722 (N_35722,N_33635,N_33100);
and U35723 (N_35723,N_32608,N_33408);
nand U35724 (N_35724,N_33470,N_32272);
nand U35725 (N_35725,N_32724,N_33949);
xnor U35726 (N_35726,N_32824,N_32008);
nand U35727 (N_35727,N_33325,N_32078);
nand U35728 (N_35728,N_33074,N_33326);
nor U35729 (N_35729,N_32749,N_32214);
or U35730 (N_35730,N_33514,N_33393);
and U35731 (N_35731,N_32019,N_33631);
nor U35732 (N_35732,N_33106,N_32744);
xor U35733 (N_35733,N_33121,N_32693);
and U35734 (N_35734,N_33736,N_33991);
nor U35735 (N_35735,N_32065,N_32779);
or U35736 (N_35736,N_33084,N_32792);
or U35737 (N_35737,N_32680,N_33786);
nor U35738 (N_35738,N_33621,N_32074);
xor U35739 (N_35739,N_32146,N_32831);
xnor U35740 (N_35740,N_33010,N_32583);
xnor U35741 (N_35741,N_33330,N_32044);
nand U35742 (N_35742,N_32417,N_32870);
xor U35743 (N_35743,N_32807,N_32468);
xor U35744 (N_35744,N_33676,N_32736);
nand U35745 (N_35745,N_32856,N_32449);
xor U35746 (N_35746,N_32697,N_33859);
nor U35747 (N_35747,N_32865,N_32723);
and U35748 (N_35748,N_32385,N_32695);
or U35749 (N_35749,N_33910,N_32603);
nand U35750 (N_35750,N_33528,N_32878);
and U35751 (N_35751,N_32676,N_33104);
and U35752 (N_35752,N_33225,N_32869);
nor U35753 (N_35753,N_32589,N_32411);
nand U35754 (N_35754,N_32668,N_32821);
or U35755 (N_35755,N_33690,N_33723);
and U35756 (N_35756,N_33774,N_33451);
nand U35757 (N_35757,N_32831,N_32253);
and U35758 (N_35758,N_33760,N_32492);
or U35759 (N_35759,N_33052,N_32506);
and U35760 (N_35760,N_33342,N_33831);
xor U35761 (N_35761,N_32833,N_32060);
and U35762 (N_35762,N_33809,N_32347);
or U35763 (N_35763,N_33493,N_33121);
and U35764 (N_35764,N_32514,N_32125);
and U35765 (N_35765,N_32980,N_32744);
or U35766 (N_35766,N_33461,N_32097);
or U35767 (N_35767,N_33216,N_32338);
and U35768 (N_35768,N_33489,N_33204);
xor U35769 (N_35769,N_33251,N_33173);
nand U35770 (N_35770,N_33065,N_32976);
or U35771 (N_35771,N_33051,N_33479);
and U35772 (N_35772,N_33415,N_33723);
or U35773 (N_35773,N_32691,N_33119);
xor U35774 (N_35774,N_32625,N_32454);
xnor U35775 (N_35775,N_33575,N_32363);
nand U35776 (N_35776,N_32339,N_32628);
and U35777 (N_35777,N_32676,N_33030);
or U35778 (N_35778,N_33492,N_33389);
xor U35779 (N_35779,N_32620,N_32301);
xnor U35780 (N_35780,N_33791,N_32391);
nand U35781 (N_35781,N_33838,N_33321);
or U35782 (N_35782,N_33070,N_33933);
xnor U35783 (N_35783,N_32401,N_33729);
and U35784 (N_35784,N_33587,N_33420);
xnor U35785 (N_35785,N_33140,N_32672);
nand U35786 (N_35786,N_33827,N_32286);
and U35787 (N_35787,N_33756,N_32142);
nand U35788 (N_35788,N_33153,N_33043);
or U35789 (N_35789,N_33890,N_33472);
or U35790 (N_35790,N_33640,N_32462);
or U35791 (N_35791,N_33135,N_32493);
or U35792 (N_35792,N_33235,N_32543);
nor U35793 (N_35793,N_33046,N_33881);
nand U35794 (N_35794,N_32339,N_32436);
nor U35795 (N_35795,N_33731,N_32210);
nand U35796 (N_35796,N_33132,N_33894);
or U35797 (N_35797,N_33749,N_33715);
or U35798 (N_35798,N_32468,N_32013);
or U35799 (N_35799,N_33832,N_32169);
nor U35800 (N_35800,N_32170,N_32296);
xnor U35801 (N_35801,N_33160,N_32497);
and U35802 (N_35802,N_32475,N_32348);
nand U35803 (N_35803,N_33561,N_33537);
xor U35804 (N_35804,N_33902,N_33442);
nor U35805 (N_35805,N_32519,N_33610);
nor U35806 (N_35806,N_33968,N_33473);
xor U35807 (N_35807,N_33465,N_33357);
nor U35808 (N_35808,N_32427,N_33279);
nor U35809 (N_35809,N_32638,N_33656);
nor U35810 (N_35810,N_33892,N_32420);
and U35811 (N_35811,N_33384,N_32189);
xnor U35812 (N_35812,N_32513,N_33847);
or U35813 (N_35813,N_32772,N_32652);
or U35814 (N_35814,N_33900,N_33041);
or U35815 (N_35815,N_32059,N_32463);
and U35816 (N_35816,N_33620,N_33806);
nor U35817 (N_35817,N_33317,N_33624);
or U35818 (N_35818,N_32078,N_33774);
nand U35819 (N_35819,N_32756,N_33692);
or U35820 (N_35820,N_33200,N_33288);
nor U35821 (N_35821,N_33694,N_32624);
nand U35822 (N_35822,N_33838,N_33081);
nand U35823 (N_35823,N_33839,N_32876);
and U35824 (N_35824,N_32141,N_32535);
nor U35825 (N_35825,N_32141,N_32990);
xnor U35826 (N_35826,N_33673,N_32486);
xor U35827 (N_35827,N_32053,N_33587);
nor U35828 (N_35828,N_33300,N_33693);
nand U35829 (N_35829,N_33218,N_32063);
nand U35830 (N_35830,N_32504,N_32709);
and U35831 (N_35831,N_33762,N_33710);
nand U35832 (N_35832,N_33279,N_33201);
xor U35833 (N_35833,N_33350,N_33814);
xor U35834 (N_35834,N_32921,N_32509);
or U35835 (N_35835,N_33067,N_32309);
or U35836 (N_35836,N_32728,N_33384);
nand U35837 (N_35837,N_33716,N_33875);
or U35838 (N_35838,N_33762,N_32113);
nand U35839 (N_35839,N_32174,N_32044);
nor U35840 (N_35840,N_33274,N_33974);
xnor U35841 (N_35841,N_33775,N_32732);
nor U35842 (N_35842,N_32964,N_32604);
or U35843 (N_35843,N_32257,N_33658);
nor U35844 (N_35844,N_33017,N_33199);
nor U35845 (N_35845,N_33845,N_32639);
nor U35846 (N_35846,N_33902,N_33244);
nand U35847 (N_35847,N_33813,N_33421);
or U35848 (N_35848,N_33753,N_33959);
xor U35849 (N_35849,N_32011,N_33256);
xor U35850 (N_35850,N_32816,N_32071);
xor U35851 (N_35851,N_33118,N_32146);
or U35852 (N_35852,N_33377,N_32338);
and U35853 (N_35853,N_33589,N_32101);
nor U35854 (N_35854,N_32336,N_32324);
or U35855 (N_35855,N_33571,N_33743);
and U35856 (N_35856,N_33798,N_33433);
and U35857 (N_35857,N_33878,N_33874);
xnor U35858 (N_35858,N_33516,N_32542);
or U35859 (N_35859,N_33496,N_32276);
nor U35860 (N_35860,N_32880,N_33252);
and U35861 (N_35861,N_32497,N_33047);
or U35862 (N_35862,N_32664,N_33525);
nor U35863 (N_35863,N_32455,N_32015);
or U35864 (N_35864,N_32897,N_32247);
nand U35865 (N_35865,N_33539,N_33263);
nor U35866 (N_35866,N_32369,N_33272);
and U35867 (N_35867,N_32084,N_33111);
xnor U35868 (N_35868,N_33306,N_32803);
and U35869 (N_35869,N_33593,N_32735);
and U35870 (N_35870,N_32569,N_32720);
or U35871 (N_35871,N_33353,N_33179);
xor U35872 (N_35872,N_33025,N_33541);
nand U35873 (N_35873,N_32762,N_32187);
nor U35874 (N_35874,N_32113,N_32014);
nand U35875 (N_35875,N_33297,N_32570);
xor U35876 (N_35876,N_32918,N_33081);
nand U35877 (N_35877,N_32769,N_33392);
xnor U35878 (N_35878,N_33083,N_32493);
xor U35879 (N_35879,N_32004,N_33762);
or U35880 (N_35880,N_33826,N_33099);
and U35881 (N_35881,N_33344,N_33474);
and U35882 (N_35882,N_32208,N_33851);
or U35883 (N_35883,N_33951,N_32195);
or U35884 (N_35884,N_32605,N_32695);
nand U35885 (N_35885,N_32528,N_33513);
nor U35886 (N_35886,N_33475,N_32314);
and U35887 (N_35887,N_33285,N_33322);
xnor U35888 (N_35888,N_33132,N_33805);
xor U35889 (N_35889,N_33715,N_32526);
nand U35890 (N_35890,N_33147,N_33018);
and U35891 (N_35891,N_32259,N_33245);
or U35892 (N_35892,N_32075,N_32855);
nor U35893 (N_35893,N_33843,N_32430);
and U35894 (N_35894,N_33075,N_32843);
or U35895 (N_35895,N_33046,N_32049);
xnor U35896 (N_35896,N_32191,N_33201);
nor U35897 (N_35897,N_32860,N_32698);
xnor U35898 (N_35898,N_33045,N_32079);
or U35899 (N_35899,N_32829,N_32168);
nor U35900 (N_35900,N_32120,N_32582);
and U35901 (N_35901,N_33883,N_32429);
or U35902 (N_35902,N_32938,N_33289);
xnor U35903 (N_35903,N_33222,N_33708);
or U35904 (N_35904,N_32887,N_33034);
xor U35905 (N_35905,N_32683,N_32709);
xor U35906 (N_35906,N_33620,N_33449);
and U35907 (N_35907,N_32077,N_33232);
and U35908 (N_35908,N_33973,N_33969);
xnor U35909 (N_35909,N_32625,N_33383);
nand U35910 (N_35910,N_33016,N_32472);
and U35911 (N_35911,N_32885,N_32075);
nand U35912 (N_35912,N_33660,N_33445);
xnor U35913 (N_35913,N_33761,N_32345);
xnor U35914 (N_35914,N_33891,N_33165);
or U35915 (N_35915,N_32792,N_32842);
and U35916 (N_35916,N_32594,N_33949);
or U35917 (N_35917,N_32949,N_32911);
and U35918 (N_35918,N_33823,N_33338);
and U35919 (N_35919,N_33902,N_33389);
xor U35920 (N_35920,N_33039,N_33771);
nor U35921 (N_35921,N_33116,N_32408);
or U35922 (N_35922,N_32298,N_32973);
nand U35923 (N_35923,N_33260,N_33647);
or U35924 (N_35924,N_32520,N_32655);
nor U35925 (N_35925,N_32124,N_33682);
or U35926 (N_35926,N_33597,N_32523);
or U35927 (N_35927,N_33570,N_32197);
xor U35928 (N_35928,N_32654,N_32389);
and U35929 (N_35929,N_32353,N_33905);
nand U35930 (N_35930,N_33846,N_32998);
nor U35931 (N_35931,N_32688,N_33310);
or U35932 (N_35932,N_32309,N_33593);
nand U35933 (N_35933,N_32263,N_33511);
and U35934 (N_35934,N_33640,N_32561);
or U35935 (N_35935,N_33980,N_32373);
nand U35936 (N_35936,N_33924,N_33978);
or U35937 (N_35937,N_32190,N_33753);
nor U35938 (N_35938,N_33802,N_33195);
nor U35939 (N_35939,N_33241,N_32789);
xnor U35940 (N_35940,N_33692,N_33116);
or U35941 (N_35941,N_33611,N_32005);
nor U35942 (N_35942,N_32520,N_33906);
nand U35943 (N_35943,N_33597,N_33145);
nor U35944 (N_35944,N_32425,N_33954);
and U35945 (N_35945,N_33771,N_32656);
and U35946 (N_35946,N_32472,N_33415);
or U35947 (N_35947,N_32596,N_32953);
xnor U35948 (N_35948,N_33512,N_32146);
and U35949 (N_35949,N_32439,N_32917);
and U35950 (N_35950,N_33519,N_33829);
nor U35951 (N_35951,N_33144,N_32771);
and U35952 (N_35952,N_32046,N_32335);
or U35953 (N_35953,N_33777,N_33717);
nor U35954 (N_35954,N_33456,N_32897);
or U35955 (N_35955,N_33551,N_33983);
xnor U35956 (N_35956,N_32304,N_33263);
nor U35957 (N_35957,N_32175,N_33498);
nand U35958 (N_35958,N_32944,N_32807);
nand U35959 (N_35959,N_33802,N_33948);
or U35960 (N_35960,N_32009,N_32187);
and U35961 (N_35961,N_33970,N_32166);
nand U35962 (N_35962,N_32571,N_33779);
nand U35963 (N_35963,N_32352,N_33704);
and U35964 (N_35964,N_32712,N_33107);
and U35965 (N_35965,N_32305,N_32866);
xor U35966 (N_35966,N_33977,N_33249);
xor U35967 (N_35967,N_33645,N_33170);
nand U35968 (N_35968,N_32565,N_32076);
nor U35969 (N_35969,N_33876,N_33627);
nor U35970 (N_35970,N_32761,N_32049);
or U35971 (N_35971,N_33929,N_32566);
nand U35972 (N_35972,N_32694,N_33207);
and U35973 (N_35973,N_33785,N_33758);
xnor U35974 (N_35974,N_32253,N_33244);
or U35975 (N_35975,N_32488,N_32621);
and U35976 (N_35976,N_32901,N_33189);
and U35977 (N_35977,N_32323,N_32983);
or U35978 (N_35978,N_33640,N_33964);
xnor U35979 (N_35979,N_32031,N_32677);
xnor U35980 (N_35980,N_33189,N_33841);
nand U35981 (N_35981,N_33356,N_33481);
xor U35982 (N_35982,N_33367,N_33306);
nor U35983 (N_35983,N_32572,N_32656);
xor U35984 (N_35984,N_33780,N_32303);
and U35985 (N_35985,N_32231,N_33261);
and U35986 (N_35986,N_33914,N_33394);
nand U35987 (N_35987,N_32372,N_33355);
nor U35988 (N_35988,N_32113,N_32448);
xnor U35989 (N_35989,N_33267,N_33548);
or U35990 (N_35990,N_32741,N_33163);
and U35991 (N_35991,N_33438,N_32606);
nand U35992 (N_35992,N_33062,N_33777);
and U35993 (N_35993,N_32642,N_32235);
and U35994 (N_35994,N_32842,N_32363);
nor U35995 (N_35995,N_32618,N_33440);
and U35996 (N_35996,N_32890,N_33712);
and U35997 (N_35997,N_32812,N_33209);
or U35998 (N_35998,N_32647,N_33648);
nor U35999 (N_35999,N_32172,N_33066);
nand U36000 (N_36000,N_35692,N_34793);
nand U36001 (N_36001,N_35454,N_35456);
nor U36002 (N_36002,N_34589,N_35082);
or U36003 (N_36003,N_35283,N_34180);
and U36004 (N_36004,N_35187,N_34039);
nor U36005 (N_36005,N_34247,N_34116);
or U36006 (N_36006,N_35872,N_35934);
or U36007 (N_36007,N_35693,N_34009);
xnor U36008 (N_36008,N_35084,N_34171);
or U36009 (N_36009,N_35570,N_35834);
xnor U36010 (N_36010,N_34233,N_35806);
or U36011 (N_36011,N_35359,N_35729);
xor U36012 (N_36012,N_35053,N_34702);
xor U36013 (N_36013,N_35541,N_34572);
or U36014 (N_36014,N_35509,N_35211);
xnor U36015 (N_36015,N_34908,N_34129);
or U36016 (N_36016,N_35478,N_34272);
and U36017 (N_36017,N_34303,N_34024);
nand U36018 (N_36018,N_34723,N_35195);
xor U36019 (N_36019,N_34652,N_34422);
nand U36020 (N_36020,N_34077,N_35214);
nor U36021 (N_36021,N_35865,N_35320);
nand U36022 (N_36022,N_34862,N_34537);
and U36023 (N_36023,N_35831,N_35114);
xor U36024 (N_36024,N_34395,N_34670);
or U36025 (N_36025,N_34201,N_34837);
nand U36026 (N_36026,N_34642,N_34256);
nand U36027 (N_36027,N_34358,N_34415);
nor U36028 (N_36028,N_35725,N_35614);
or U36029 (N_36029,N_35567,N_34444);
nand U36030 (N_36030,N_35916,N_34665);
xor U36031 (N_36031,N_34337,N_34559);
or U36032 (N_36032,N_35315,N_34248);
or U36033 (N_36033,N_35559,N_34599);
xnor U36034 (N_36034,N_34551,N_34547);
or U36035 (N_36035,N_34174,N_34743);
nand U36036 (N_36036,N_35455,N_35892);
and U36037 (N_36037,N_34015,N_35005);
and U36038 (N_36038,N_35905,N_34825);
or U36039 (N_36039,N_35293,N_35881);
xnor U36040 (N_36040,N_35471,N_34838);
nor U36041 (N_36041,N_35586,N_34666);
nand U36042 (N_36042,N_34041,N_34591);
nor U36043 (N_36043,N_35982,N_35165);
xnor U36044 (N_36044,N_35024,N_35687);
and U36045 (N_36045,N_35357,N_34208);
and U36046 (N_36046,N_35378,N_35969);
xor U36047 (N_36047,N_35135,N_34413);
nand U36048 (N_36048,N_35757,N_34001);
nand U36049 (N_36049,N_34404,N_35812);
nand U36050 (N_36050,N_35708,N_34586);
and U36051 (N_36051,N_35001,N_35664);
or U36052 (N_36052,N_35741,N_34219);
nand U36053 (N_36053,N_35717,N_35893);
or U36054 (N_36054,N_35353,N_34207);
and U36055 (N_36055,N_35434,N_35032);
or U36056 (N_36056,N_35610,N_35801);
nand U36057 (N_36057,N_35700,N_35154);
xor U36058 (N_36058,N_34524,N_35677);
nand U36059 (N_36059,N_34013,N_34382);
xor U36060 (N_36060,N_35047,N_35612);
or U36061 (N_36061,N_34437,N_34979);
nor U36062 (N_36062,N_35854,N_35852);
nand U36063 (N_36063,N_34084,N_34312);
nand U36064 (N_36064,N_35274,N_35156);
xnor U36065 (N_36065,N_34896,N_34265);
and U36066 (N_36066,N_34562,N_35759);
and U36067 (N_36067,N_34257,N_34785);
and U36068 (N_36068,N_35185,N_34392);
and U36069 (N_36069,N_35799,N_34971);
xnor U36070 (N_36070,N_35606,N_35948);
nor U36071 (N_36071,N_34092,N_35894);
nand U36072 (N_36072,N_34611,N_35367);
and U36073 (N_36073,N_35262,N_35583);
xnor U36074 (N_36074,N_35520,N_34700);
or U36075 (N_36075,N_35221,N_35105);
nand U36076 (N_36076,N_34860,N_35292);
nor U36077 (N_36077,N_35825,N_34450);
nor U36078 (N_36078,N_34117,N_34906);
or U36079 (N_36079,N_35575,N_35295);
nor U36080 (N_36080,N_34465,N_35668);
nand U36081 (N_36081,N_34922,N_34058);
and U36082 (N_36082,N_34717,N_34606);
nor U36083 (N_36083,N_34806,N_35231);
nand U36084 (N_36084,N_34703,N_35415);
or U36085 (N_36085,N_35038,N_35213);
and U36086 (N_36086,N_34495,N_35818);
nor U36087 (N_36087,N_34302,N_34133);
nor U36088 (N_36088,N_34503,N_34255);
nor U36089 (N_36089,N_35383,N_35308);
nand U36090 (N_36090,N_34430,N_35448);
and U36091 (N_36091,N_35226,N_35273);
and U36092 (N_36092,N_35630,N_34683);
xnor U36093 (N_36093,N_35751,N_35322);
nand U36094 (N_36094,N_34060,N_34391);
or U36095 (N_36095,N_35793,N_34941);
nand U36096 (N_36096,N_35596,N_35469);
xor U36097 (N_36097,N_34294,N_34138);
and U36098 (N_36098,N_35390,N_34622);
nor U36099 (N_36099,N_35473,N_34780);
nand U36100 (N_36100,N_35549,N_35632);
and U36101 (N_36101,N_35666,N_35403);
nand U36102 (N_36102,N_35451,N_34992);
or U36103 (N_36103,N_35023,N_34890);
or U36104 (N_36104,N_35622,N_35754);
nand U36105 (N_36105,N_34710,N_35323);
and U36106 (N_36106,N_34200,N_34976);
nor U36107 (N_36107,N_35885,N_34298);
nand U36108 (N_36108,N_35765,N_35095);
or U36109 (N_36109,N_35843,N_35527);
xnor U36110 (N_36110,N_34831,N_35072);
xnor U36111 (N_36111,N_34584,N_35984);
or U36112 (N_36112,N_35564,N_34159);
or U36113 (N_36113,N_35774,N_34716);
xor U36114 (N_36114,N_34292,N_34891);
nand U36115 (N_36115,N_35930,N_34799);
nor U36116 (N_36116,N_34000,N_34148);
nor U36117 (N_36117,N_34915,N_35420);
nor U36118 (N_36118,N_35925,N_35137);
nor U36119 (N_36119,N_35873,N_35395);
nor U36120 (N_36120,N_35251,N_34545);
or U36121 (N_36121,N_34453,N_35974);
xnor U36122 (N_36122,N_34763,N_35887);
nor U36123 (N_36123,N_34898,N_34705);
nor U36124 (N_36124,N_34033,N_35372);
xor U36125 (N_36125,N_35380,N_34616);
or U36126 (N_36126,N_35722,N_35052);
nor U36127 (N_36127,N_35216,N_35310);
or U36128 (N_36128,N_34658,N_34140);
and U36129 (N_36129,N_35710,N_35627);
and U36130 (N_36130,N_35965,N_34446);
nand U36131 (N_36131,N_35270,N_34252);
xor U36132 (N_36132,N_35588,N_35162);
xnor U36133 (N_36133,N_34181,N_34509);
nand U36134 (N_36134,N_34045,N_35938);
nor U36135 (N_36135,N_35504,N_35025);
and U36136 (N_36136,N_34680,N_35712);
and U36137 (N_36137,N_34516,N_34070);
nand U36138 (N_36138,N_34428,N_34685);
or U36139 (N_36139,N_34850,N_34003);
nand U36140 (N_36140,N_35337,N_35816);
or U36141 (N_36141,N_34938,N_35261);
and U36142 (N_36142,N_34594,N_34724);
xor U36143 (N_36143,N_35497,N_35903);
nor U36144 (N_36144,N_35902,N_34903);
xor U36145 (N_36145,N_34955,N_34401);
nor U36146 (N_36146,N_35417,N_34089);
and U36147 (N_36147,N_34739,N_35747);
xor U36148 (N_36148,N_35506,N_34028);
xor U36149 (N_36149,N_34919,N_34281);
xnor U36150 (N_36150,N_34223,N_35134);
and U36151 (N_36151,N_34355,N_35371);
nand U36152 (N_36152,N_34911,N_34317);
nor U36153 (N_36153,N_35241,N_34918);
nor U36154 (N_36154,N_35858,N_34244);
xor U36155 (N_36155,N_34188,N_35242);
nand U36156 (N_36156,N_34985,N_34556);
xor U36157 (N_36157,N_34479,N_35699);
xor U36158 (N_36158,N_35142,N_35617);
and U36159 (N_36159,N_34369,N_34651);
or U36160 (N_36160,N_34823,N_34367);
xor U36161 (N_36161,N_35795,N_35602);
nor U36162 (N_36162,N_34502,N_35387);
or U36163 (N_36163,N_35492,N_35169);
or U36164 (N_36164,N_34494,N_34820);
xor U36165 (N_36165,N_35484,N_35418);
or U36166 (N_36166,N_35136,N_35198);
xnor U36167 (N_36167,N_35212,N_34674);
and U36168 (N_36168,N_34696,N_34101);
nor U36169 (N_36169,N_34788,N_35869);
or U36170 (N_36170,N_35091,N_35150);
and U36171 (N_36171,N_35821,N_35794);
or U36172 (N_36172,N_35393,N_34935);
and U36173 (N_36173,N_34929,N_35440);
and U36174 (N_36174,N_35408,N_34832);
xor U36175 (N_36175,N_35953,N_35155);
and U36176 (N_36176,N_34859,N_34673);
nor U36177 (N_36177,N_35963,N_35516);
nand U36178 (N_36178,N_34669,N_34974);
xor U36179 (N_36179,N_35370,N_35083);
xor U36180 (N_36180,N_35051,N_34924);
or U36181 (N_36181,N_34197,N_35642);
nor U36182 (N_36182,N_35254,N_34814);
or U36183 (N_36183,N_34688,N_35167);
and U36184 (N_36184,N_35446,N_35303);
and U36185 (N_36185,N_35714,N_34151);
nand U36186 (N_36186,N_34725,N_35979);
xnor U36187 (N_36187,N_35592,N_34283);
nor U36188 (N_36188,N_35442,N_34517);
and U36189 (N_36189,N_34709,N_35316);
xor U36190 (N_36190,N_35724,N_34243);
nand U36191 (N_36191,N_34293,N_35581);
or U36192 (N_36192,N_34533,N_34712);
or U36193 (N_36193,N_35635,N_34552);
and U36194 (N_36194,N_34774,N_35042);
nor U36195 (N_36195,N_34754,N_34889);
nor U36196 (N_36196,N_35686,N_34393);
or U36197 (N_36197,N_34612,N_34273);
xnor U36198 (N_36198,N_35886,N_35347);
nor U36199 (N_36199,N_35284,N_34377);
or U36200 (N_36200,N_35628,N_35603);
xor U36201 (N_36201,N_35066,N_35998);
xor U36202 (N_36202,N_35229,N_34407);
xnor U36203 (N_36203,N_35120,N_35048);
nand U36204 (N_36204,N_35595,N_35059);
or U36205 (N_36205,N_35561,N_34948);
nand U36206 (N_36206,N_34105,N_35553);
nand U36207 (N_36207,N_35133,N_34930);
nor U36208 (N_36208,N_35576,N_34098);
nand U36209 (N_36209,N_34123,N_35736);
nand U36210 (N_36210,N_35220,N_34681);
xnor U36211 (N_36211,N_35030,N_35179);
nor U36212 (N_36212,N_34500,N_34878);
xor U36213 (N_36213,N_35463,N_34328);
and U36214 (N_36214,N_34693,N_34203);
xnor U36215 (N_36215,N_34557,N_35917);
and U36216 (N_36216,N_35003,N_35379);
nor U36217 (N_36217,N_34625,N_35591);
or U36218 (N_36218,N_35494,N_34514);
and U36219 (N_36219,N_35349,N_34964);
and U36220 (N_36220,N_35600,N_34234);
or U36221 (N_36221,N_35698,N_35870);
or U36222 (N_36222,N_35897,N_35111);
nand U36223 (N_36223,N_35180,N_35148);
xor U36224 (N_36224,N_34141,N_35788);
and U36225 (N_36225,N_34664,N_35577);
nor U36226 (N_36226,N_34711,N_34677);
nand U36227 (N_36227,N_34068,N_34759);
and U36228 (N_36228,N_35287,N_34425);
nor U36229 (N_36229,N_35046,N_34966);
nand U36230 (N_36230,N_34018,N_35988);
nand U36231 (N_36231,N_35809,N_35425);
and U36232 (N_36232,N_34866,N_35620);
nor U36233 (N_36233,N_34132,N_34854);
xnor U36234 (N_36234,N_34370,N_34322);
xor U36235 (N_36235,N_35493,N_35312);
nand U36236 (N_36236,N_35459,N_34513);
or U36237 (N_36237,N_35803,N_35594);
and U36238 (N_36238,N_34926,N_35785);
and U36239 (N_36239,N_34816,N_35512);
xnor U36240 (N_36240,N_34157,N_35758);
nor U36241 (N_36241,N_35110,N_34353);
and U36242 (N_36242,N_35715,N_35720);
and U36243 (N_36243,N_34289,N_34999);
nor U36244 (N_36244,N_34176,N_35407);
and U36245 (N_36245,N_34629,N_34508);
nor U36246 (N_36246,N_34639,N_35298);
and U36247 (N_36247,N_35108,N_35129);
or U36248 (N_36248,N_35099,N_35615);
xor U36249 (N_36249,N_35234,N_34541);
and U36250 (N_36250,N_35695,N_35365);
or U36251 (N_36251,N_35299,N_35483);
xnor U36252 (N_36252,N_35962,N_34732);
and U36253 (N_36253,N_34021,N_35264);
nor U36254 (N_36254,N_34419,N_35074);
nor U36255 (N_36255,N_34183,N_34139);
or U36256 (N_36256,N_35524,N_34268);
and U36257 (N_36257,N_35486,N_35311);
and U36258 (N_36258,N_34744,N_34359);
nand U36259 (N_36259,N_34817,N_34905);
or U36260 (N_36260,N_34083,N_34834);
nor U36261 (N_36261,N_34261,N_34950);
and U36262 (N_36262,N_34477,N_34094);
xnor U36263 (N_36263,N_34363,N_35054);
nor U36264 (N_36264,N_34645,N_35625);
and U36265 (N_36265,N_34279,N_34080);
and U36266 (N_36266,N_35513,N_35236);
or U36267 (N_36267,N_34145,N_35992);
or U36268 (N_36268,N_35205,N_34102);
or U36269 (N_36269,N_34323,N_35530);
and U36270 (N_36270,N_35944,N_35662);
or U36271 (N_36271,N_34338,N_35374);
or U36272 (N_36272,N_35288,N_35723);
nor U36273 (N_36273,N_35611,N_34857);
xnor U36274 (N_36274,N_35325,N_34287);
nor U36275 (N_36275,N_34345,N_35884);
xor U36276 (N_36276,N_35652,N_35853);
or U36277 (N_36277,N_35739,N_34120);
xor U36278 (N_36278,N_35866,N_35279);
nand U36279 (N_36279,N_35272,N_35608);
nor U36280 (N_36280,N_34959,N_35623);
or U36281 (N_36281,N_34427,N_34871);
or U36282 (N_36282,N_34153,N_35871);
xor U36283 (N_36283,N_34779,N_34927);
nor U36284 (N_36284,N_34168,N_35546);
or U36285 (N_36285,N_34987,N_34472);
nor U36286 (N_36286,N_35305,N_34262);
xor U36287 (N_36287,N_35186,N_34628);
nand U36288 (N_36288,N_35840,N_35034);
and U36289 (N_36289,N_35369,N_34191);
or U36290 (N_36290,N_34086,N_34598);
and U36291 (N_36291,N_34571,N_34037);
nor U36292 (N_36292,N_34436,N_35659);
nor U36293 (N_36293,N_34631,N_34947);
xnor U36294 (N_36294,N_35833,N_35647);
nand U36295 (N_36295,N_35939,N_34142);
or U36296 (N_36296,N_35629,N_34373);
nand U36297 (N_36297,N_34886,N_34755);
or U36298 (N_36298,N_34592,N_35731);
xor U36299 (N_36299,N_34331,N_34112);
nor U36300 (N_36300,N_34035,N_35452);
or U36301 (N_36301,N_34726,N_34136);
nor U36302 (N_36302,N_34242,N_34555);
or U36303 (N_36303,N_34963,N_35718);
nor U36304 (N_36304,N_35200,N_35604);
nand U36305 (N_36305,N_35580,N_34747);
xnor U36306 (N_36306,N_34879,N_35055);
xor U36307 (N_36307,N_35680,N_34036);
or U36308 (N_36308,N_35007,N_34752);
nand U36309 (N_36309,N_35118,N_35783);
nor U36310 (N_36310,N_35981,N_35020);
nor U36311 (N_36311,N_34280,N_34127);
xnor U36312 (N_36312,N_35923,N_34249);
or U36313 (N_36313,N_35745,N_35972);
and U36314 (N_36314,N_34314,N_35521);
nand U36315 (N_36315,N_34577,N_35268);
xnor U36316 (N_36316,N_34967,N_34489);
nand U36317 (N_36317,N_35314,N_35073);
or U36318 (N_36318,N_34520,N_34231);
nor U36319 (N_36319,N_34167,N_34376);
nor U36320 (N_36320,N_35946,N_34789);
or U36321 (N_36321,N_35648,N_34528);
or U36322 (N_36322,N_35249,N_35276);
and U36323 (N_36323,N_35289,N_34291);
or U36324 (N_36324,N_34569,N_35368);
nand U36325 (N_36325,N_35624,N_35384);
nor U36326 (N_36326,N_35940,N_34729);
or U36327 (N_36327,N_35814,N_34097);
or U36328 (N_36328,N_34025,N_34321);
and U36329 (N_36329,N_34232,N_34305);
and U36330 (N_36330,N_35343,N_35574);
xnor U36331 (N_36331,N_35883,N_35499);
xnor U36332 (N_36332,N_34384,N_35050);
xor U36333 (N_36333,N_35790,N_34530);
nor U36334 (N_36334,N_34689,N_34196);
and U36335 (N_36335,N_34354,N_35784);
and U36336 (N_36336,N_34307,N_34390);
nand U36337 (N_36337,N_35550,N_35081);
and U36338 (N_36338,N_35485,N_35970);
xnor U36339 (N_36339,N_35014,N_35752);
and U36340 (N_36340,N_35037,N_35457);
and U36341 (N_36341,N_35829,N_35145);
or U36342 (N_36342,N_34497,N_35004);
nand U36343 (N_36343,N_35470,N_34099);
nand U36344 (N_36344,N_34435,N_34982);
nor U36345 (N_36345,N_34676,N_34748);
or U36346 (N_36346,N_34017,N_34381);
nand U36347 (N_36347,N_34897,N_34205);
xnor U36348 (N_36348,N_34412,N_34893);
xnor U36349 (N_36349,N_35479,N_34449);
and U36350 (N_36350,N_34357,N_34753);
nand U36351 (N_36351,N_34065,N_34177);
nand U36352 (N_36352,N_34276,N_34184);
and U36353 (N_36353,N_34568,N_35542);
nor U36354 (N_36354,N_35565,N_35787);
xor U36355 (N_36355,N_34202,N_34684);
and U36356 (N_36356,N_35356,N_34483);
and U36357 (N_36357,N_35011,N_34836);
and U36358 (N_36358,N_34316,N_34301);
and U36359 (N_36359,N_34643,N_35445);
nand U36360 (N_36360,N_35225,N_35002);
xor U36361 (N_36361,N_35453,N_35507);
and U36362 (N_36362,N_35296,N_35245);
and U36363 (N_36363,N_35411,N_35980);
nor U36364 (N_36364,N_34030,N_35531);
and U36365 (N_36365,N_34944,N_34870);
or U36366 (N_36366,N_34124,N_35913);
or U36367 (N_36367,N_35820,N_34697);
nand U36368 (N_36368,N_34469,N_35100);
nand U36369 (N_36369,N_34061,N_34968);
nor U36370 (N_36370,N_34518,N_34965);
nor U36371 (N_36371,N_35404,N_34226);
xor U36372 (N_36372,N_34274,N_35027);
nor U36373 (N_36373,N_35830,N_34805);
nor U36374 (N_36374,N_34904,N_34161);
nor U36375 (N_36375,N_35703,N_34221);
xor U36376 (N_36376,N_34016,N_35915);
and U36377 (N_36377,N_34179,N_34601);
nand U36378 (N_36378,N_34750,N_34588);
nor U36379 (N_36379,N_35092,N_34423);
and U36380 (N_36380,N_34678,N_34459);
nand U36381 (N_36381,N_35300,N_34564);
nand U36382 (N_36382,N_35545,N_35430);
or U36383 (N_36383,N_35709,N_35235);
xor U36384 (N_36384,N_35875,N_34051);
and U36385 (N_36385,N_34214,N_34728);
nand U36386 (N_36386,N_34366,N_35243);
nand U36387 (N_36387,N_34844,N_35432);
nand U36388 (N_36388,N_34064,N_34330);
or U36389 (N_36389,N_35975,N_35436);
xnor U36390 (N_36390,N_35260,N_34341);
and U36391 (N_36391,N_34198,N_35317);
nand U36392 (N_36392,N_35267,N_35888);
and U36393 (N_36393,N_34309,N_35044);
nor U36394 (N_36394,N_35090,N_35398);
or U36395 (N_36395,N_35966,N_35598);
or U36396 (N_36396,N_35360,N_35748);
or U36397 (N_36397,N_34576,N_35294);
nor U36398 (N_36398,N_34027,N_35836);
nand U36399 (N_36399,N_34109,N_35321);
or U36400 (N_36400,N_34544,N_35067);
xor U36401 (N_36401,N_34956,N_35086);
and U36402 (N_36402,N_35345,N_34325);
and U36403 (N_36403,N_34641,N_34949);
nand U36404 (N_36404,N_35579,N_34672);
and U36405 (N_36405,N_34761,N_35339);
xnor U36406 (N_36406,N_34189,N_34119);
nor U36407 (N_36407,N_35889,N_34902);
nand U36408 (N_36408,N_35706,N_34154);
nor U36409 (N_36409,N_35775,N_34451);
and U36410 (N_36410,N_35307,N_35015);
xnor U36411 (N_36411,N_35319,N_34909);
nand U36412 (N_36412,N_35914,N_35688);
xnor U36413 (N_36413,N_34111,N_34736);
nand U36414 (N_36414,N_35450,N_34484);
or U36415 (N_36415,N_35558,N_34914);
xnor U36416 (N_36416,N_35522,N_34636);
or U36417 (N_36417,N_34554,N_34861);
nand U36418 (N_36418,N_34319,N_35846);
xnor U36419 (N_36419,N_35824,N_34285);
nand U36420 (N_36420,N_34720,N_34237);
xnor U36421 (N_36421,N_34361,N_34146);
or U36422 (N_36422,N_35904,N_35727);
or U36423 (N_36423,N_35743,N_35767);
nand U36424 (N_36424,N_35266,N_35665);
nand U36425 (N_36425,N_34011,N_34055);
nor U36426 (N_36426,N_34730,N_34867);
and U36427 (N_36427,N_34082,N_35153);
nor U36428 (N_36428,N_34858,N_35125);
or U36429 (N_36429,N_34187,N_35679);
nor U36430 (N_36430,N_34646,N_34130);
nand U36431 (N_36431,N_34199,N_35514);
and U36432 (N_36432,N_34057,N_35143);
nor U36433 (N_36433,N_34596,N_34063);
and U36434 (N_36434,N_35800,N_35638);
xnor U36435 (N_36435,N_35016,N_35589);
and U36436 (N_36436,N_34883,N_35518);
xnor U36437 (N_36437,N_34795,N_35676);
nor U36438 (N_36438,N_35076,N_35945);
and U36439 (N_36439,N_34595,N_34721);
and U36440 (N_36440,N_35204,N_35949);
and U36441 (N_36441,N_34880,N_34784);
xnor U36442 (N_36442,N_35912,N_35756);
and U36443 (N_36443,N_34856,N_35104);
nand U36444 (N_36444,N_35855,N_35728);
nor U36445 (N_36445,N_35070,N_34560);
nand U36446 (N_36446,N_35957,N_34931);
and U36447 (N_36447,N_34951,N_34888);
or U36448 (N_36448,N_35246,N_35193);
xor U36449 (N_36449,N_34843,N_34884);
nor U36450 (N_36450,N_35943,N_34627);
nor U36451 (N_36451,N_34110,N_34212);
and U36452 (N_36452,N_35428,N_35275);
or U36453 (N_36453,N_34458,N_34473);
nor U36454 (N_36454,N_35472,N_35797);
xnor U36455 (N_36455,N_35536,N_34031);
and U36456 (N_36456,N_35619,N_35286);
nor U36457 (N_36457,N_34398,N_35977);
nand U36458 (N_36458,N_34770,N_34192);
nor U36459 (N_36459,N_35828,N_34983);
nand U36460 (N_36460,N_35633,N_35909);
and U36461 (N_36461,N_35777,N_35540);
and U36462 (N_36462,N_35621,N_35626);
nand U36463 (N_36463,N_35569,N_34523);
and U36464 (N_36464,N_35281,N_35094);
and U36465 (N_36465,N_34839,N_34254);
nor U36466 (N_36466,N_34481,N_34173);
and U36467 (N_36467,N_34447,N_35995);
and U36468 (N_36468,N_34998,N_35529);
and U36469 (N_36469,N_35764,N_35402);
nand U36470 (N_36470,N_35146,N_35474);
xnor U36471 (N_36471,N_35851,N_35489);
or U36472 (N_36472,N_35358,N_35999);
nand U36473 (N_36473,N_34213,N_34186);
nand U36474 (N_36474,N_34848,N_35978);
and U36475 (N_36475,N_34371,N_34618);
xnor U36476 (N_36476,N_34434,N_34215);
xnor U36477 (N_36477,N_35132,N_34026);
nand U36478 (N_36478,N_34981,N_35753);
xnor U36479 (N_36479,N_34808,N_34326);
nor U36480 (N_36480,N_34769,N_35646);
or U36481 (N_36481,N_34813,N_34881);
xnor U36482 (N_36482,N_35056,N_35952);
nor U36483 (N_36483,N_34579,N_34029);
nor U36484 (N_36484,N_35309,N_35126);
nand U36485 (N_36485,N_34131,N_34863);
xnor U36486 (N_36486,N_35528,N_35707);
or U36487 (N_36487,N_35151,N_35557);
nand U36488 (N_36488,N_34515,N_35461);
and U36489 (N_36489,N_34454,N_34166);
xor U36490 (N_36490,N_35927,N_34091);
nand U36491 (N_36491,N_34803,N_34574);
or U36492 (N_36492,N_34038,N_34977);
nor U36493 (N_36493,N_34416,N_34360);
or U36494 (N_36494,N_35416,N_35460);
xnor U36495 (N_36495,N_34010,N_34776);
and U36496 (N_36496,N_34538,N_35163);
nor U36497 (N_36497,N_34662,N_35421);
nand U36498 (N_36498,N_34308,N_34505);
xor U36499 (N_36499,N_34442,N_35063);
nand U36500 (N_36500,N_35424,N_34235);
xnor U36501 (N_36501,N_34715,N_34827);
nand U36502 (N_36502,N_34263,N_34733);
and U36503 (N_36503,N_34845,N_35786);
xnor U36504 (N_36504,N_35227,N_34104);
nor U36505 (N_36505,N_34811,N_34869);
or U36506 (N_36506,N_35077,N_34540);
and U36507 (N_36507,N_34277,N_34757);
and U36508 (N_36508,N_35832,N_34735);
nor U36509 (N_36509,N_35218,N_34762);
or U36510 (N_36510,N_35862,N_34580);
and U36511 (N_36511,N_35819,N_35035);
nand U36512 (N_36512,N_35410,N_34046);
nor U36513 (N_36513,N_35901,N_35924);
nor U36514 (N_36514,N_34342,N_35822);
xnor U36515 (N_36515,N_34071,N_35396);
nand U36516 (N_36516,N_34614,N_35209);
nand U36517 (N_36517,N_35742,N_35304);
and U36518 (N_36518,N_34892,N_34002);
nor U36519 (N_36519,N_35324,N_34405);
or U36520 (N_36520,N_34417,N_34240);
or U36521 (N_36521,N_34096,N_35839);
or U36522 (N_36522,N_34228,N_35823);
or U36523 (N_36523,N_34841,N_34224);
xnor U36524 (N_36524,N_35192,N_34510);
xor U36525 (N_36525,N_34334,N_34954);
xor U36526 (N_36526,N_34582,N_34916);
and U36527 (N_36527,N_34164,N_34040);
nor U36528 (N_36528,N_34313,N_35386);
and U36529 (N_36529,N_34418,N_35964);
or U36530 (N_36530,N_35805,N_35942);
or U36531 (N_36531,N_35206,N_35043);
nand U36532 (N_36532,N_34085,N_34775);
xnor U36533 (N_36533,N_34553,N_35994);
nand U36534 (N_36534,N_34691,N_34828);
nand U36535 (N_36535,N_34529,N_35248);
xnor U36536 (N_36536,N_34824,N_34783);
or U36537 (N_36537,N_35439,N_34296);
or U36538 (N_36538,N_35500,N_34267);
nor U36539 (N_36539,N_34800,N_34475);
and U36540 (N_36540,N_35690,N_34193);
nand U36541 (N_36541,N_35102,N_35716);
or U36542 (N_36542,N_34374,N_35525);
xnor U36543 (N_36543,N_35616,N_35124);
and U36544 (N_36544,N_35986,N_35058);
xnor U36545 (N_36545,N_35898,N_34118);
nor U36546 (N_36546,N_34137,N_34347);
nor U36547 (N_36547,N_35848,N_34135);
or U36548 (N_36548,N_34476,N_34988);
or U36549 (N_36549,N_35475,N_34346);
nor U36550 (N_36550,N_34934,N_35908);
and U36551 (N_36551,N_34498,N_34004);
nor U36552 (N_36552,N_34657,N_34329);
and U36553 (N_36553,N_35498,N_34792);
or U36554 (N_36554,N_35019,N_34306);
xnor U36555 (N_36555,N_35993,N_34487);
or U36556 (N_36556,N_34364,N_34394);
or U36557 (N_36557,N_34012,N_35827);
or U36558 (N_36558,N_34368,N_34773);
and U36559 (N_36559,N_35427,N_35277);
and U36560 (N_36560,N_34441,N_35208);
xnor U36561 (N_36561,N_35631,N_34638);
xor U36562 (N_36562,N_35517,N_34380);
and U36563 (N_36563,N_35496,N_35060);
nor U36564 (N_36564,N_35171,N_35394);
and U36565 (N_36565,N_34932,N_34426);
or U36566 (N_36566,N_34852,N_34826);
and U36567 (N_36567,N_35278,N_35735);
xnor U36568 (N_36568,N_34807,N_35128);
or U36569 (N_36569,N_34464,N_35856);
xnor U36570 (N_36570,N_34218,N_34707);
and U36571 (N_36571,N_34053,N_35257);
nand U36572 (N_36572,N_35350,N_35363);
and U36573 (N_36573,N_35895,N_34266);
or U36574 (N_36574,N_35468,N_35449);
nor U36575 (N_36575,N_34994,N_35533);
and U36576 (N_36576,N_34007,N_34332);
or U36577 (N_36577,N_35931,N_35224);
or U36578 (N_36578,N_34694,N_34887);
or U36579 (N_36579,N_34882,N_34936);
xnor U36580 (N_36580,N_35174,N_35991);
or U36581 (N_36581,N_35896,N_34493);
nor U36582 (N_36582,N_35196,N_34343);
nor U36583 (N_36583,N_35164,N_34583);
xor U36584 (N_36584,N_34100,N_35203);
nor U36585 (N_36585,N_34150,N_34062);
or U36586 (N_36586,N_35197,N_34336);
and U36587 (N_36587,N_35364,N_34895);
or U36588 (N_36588,N_35571,N_34259);
xnor U36589 (N_36589,N_34278,N_34216);
nor U36590 (N_36590,N_34362,N_35476);
nor U36591 (N_36591,N_35560,N_35481);
and U36592 (N_36592,N_34269,N_35643);
xnor U36593 (N_36593,N_34969,N_34246);
nand U36594 (N_36594,N_34978,N_35101);
and U36595 (N_36595,N_34143,N_35910);
nor U36596 (N_36596,N_34403,N_34402);
xor U36597 (N_36597,N_35563,N_34126);
nor U36598 (N_36598,N_35392,N_35705);
nand U36599 (N_36599,N_34548,N_34833);
and U36600 (N_36600,N_34649,N_35556);
xor U36601 (N_36601,N_35194,N_35537);
or U36602 (N_36602,N_34090,N_34802);
and U36603 (N_36603,N_35333,N_34019);
or U36604 (N_36604,N_34536,N_34609);
or U36605 (N_36605,N_34438,N_34778);
or U36606 (N_36606,N_35191,N_35538);
nand U36607 (N_36607,N_35562,N_35772);
xnor U36608 (N_36608,N_34327,N_34499);
or U36609 (N_36609,N_34229,N_34005);
or U36610 (N_36610,N_35808,N_35951);
xnor U36611 (N_36611,N_34290,N_34989);
or U36612 (N_36612,N_35149,N_34535);
xnor U36613 (N_36613,N_34388,N_35173);
nor U36614 (N_36614,N_35441,N_35678);
nor U36615 (N_36615,N_35890,N_35087);
or U36616 (N_36616,N_34050,N_34840);
xor U36617 (N_36617,N_35669,N_35280);
and U36618 (N_36618,N_35510,N_34945);
xor U36619 (N_36619,N_34411,N_35259);
xnor U36620 (N_36620,N_34288,N_35107);
nand U36621 (N_36621,N_34389,N_35519);
nand U36622 (N_36622,N_34885,N_35477);
nand U36623 (N_36623,N_35302,N_34420);
nor U36624 (N_36624,N_35534,N_34375);
and U36625 (N_36625,N_34400,N_34220);
xor U36626 (N_36626,N_34095,N_34378);
xnor U36627 (N_36627,N_34953,N_34396);
nor U36628 (N_36628,N_35658,N_35237);
or U36629 (N_36629,N_35326,N_34740);
and U36630 (N_36630,N_35636,N_35645);
and U36631 (N_36631,N_35397,N_35447);
nor U36632 (N_36632,N_35250,N_35068);
xnor U36633 (N_36633,N_34457,N_34812);
nor U36634 (N_36634,N_34668,N_34692);
or U36635 (N_36635,N_35811,N_35740);
xnor U36636 (N_36636,N_34713,N_34448);
or U36637 (N_36637,N_35798,N_35649);
and U36638 (N_36638,N_34424,N_34156);
nor U36639 (N_36639,N_34864,N_34829);
or U36640 (N_36640,N_35256,N_34637);
nor U36641 (N_36641,N_35694,N_35681);
and U36642 (N_36642,N_35935,N_34573);
xnor U36643 (N_36643,N_35654,N_34340);
nor U36644 (N_36644,N_34630,N_34486);
nor U36645 (N_36645,N_34563,N_35199);
xor U36646 (N_36646,N_35726,N_34907);
or U36647 (N_36647,N_35297,N_35106);
nor U36648 (N_36648,N_34958,N_35158);
and U36649 (N_36649,N_35613,N_35921);
or U36650 (N_36650,N_35780,N_35990);
xnor U36651 (N_36651,N_34121,N_35332);
nor U36652 (N_36652,N_35989,N_35555);
and U36653 (N_36653,N_35683,N_35252);
xor U36654 (N_36654,N_35444,N_35675);
and U36655 (N_36655,N_34522,N_35340);
or U36656 (N_36656,N_34282,N_35078);
nand U36657 (N_36657,N_34491,N_35271);
nand U36658 (N_36658,N_34901,N_34431);
xor U36659 (N_36659,N_35584,N_34250);
or U36660 (N_36660,N_35548,N_34587);
and U36661 (N_36661,N_35141,N_35755);
and U36662 (N_36662,N_35290,N_34299);
xnor U36663 (N_36663,N_35926,N_34048);
nand U36664 (N_36664,N_35792,N_34115);
nand U36665 (N_36665,N_35419,N_34270);
nor U36666 (N_36666,N_34251,N_35381);
xnor U36667 (N_36667,N_34635,N_35804);
nor U36668 (N_36668,N_35013,N_35401);
or U36669 (N_36669,N_35495,N_35258);
nand U36670 (N_36670,N_35958,N_35684);
or U36671 (N_36671,N_34597,N_35713);
and U36672 (N_36672,N_35781,N_35113);
and U36673 (N_36673,N_35109,N_35230);
nand U36674 (N_36674,N_34593,N_34912);
nor U36675 (N_36675,N_34610,N_34165);
nand U36676 (N_36676,N_35508,N_35409);
or U36677 (N_36677,N_34686,N_34605);
nand U36678 (N_36678,N_35342,N_35219);
nor U36679 (N_36679,N_35188,N_35431);
or U36680 (N_36680,N_35405,N_35667);
xor U36681 (N_36681,N_35329,N_35328);
nand U36682 (N_36682,N_35670,N_34320);
or U36683 (N_36683,N_35511,N_35933);
or U36684 (N_36684,N_34633,N_34745);
nor U36685 (N_36685,N_35523,N_35069);
nor U36686 (N_36686,N_35026,N_34182);
nor U36687 (N_36687,N_35079,N_35609);
or U36688 (N_36688,N_34995,N_34650);
or U36689 (N_36689,N_34152,N_35573);
or U36690 (N_36690,N_34047,N_34008);
nand U36691 (N_36691,N_34706,N_34819);
xor U36692 (N_36692,N_34648,N_34549);
xnor U36693 (N_36693,N_34809,N_34284);
nand U36694 (N_36694,N_35776,N_34043);
nand U36695 (N_36695,N_35845,N_35351);
xnor U36696 (N_36696,N_34225,N_35433);
xor U36697 (N_36697,N_35017,N_34708);
and U36698 (N_36698,N_35177,N_35346);
nor U36699 (N_36699,N_34797,N_35202);
nand U36700 (N_36700,N_34804,N_34106);
and U36701 (N_36701,N_34718,N_34746);
and U36702 (N_36702,N_35730,N_35482);
xnor U36703 (N_36703,N_35838,N_35501);
nand U36704 (N_36704,N_35971,N_35973);
nand U36705 (N_36705,N_35691,N_35018);
xnor U36706 (N_36706,N_34865,N_35152);
or U36707 (N_36707,N_35159,N_35711);
or U36708 (N_36708,N_34561,N_35657);
xnor U36709 (N_36709,N_35587,N_35860);
and U36710 (N_36710,N_34445,N_35967);
xor U36711 (N_36711,N_35413,N_35590);
nand U36712 (N_36712,N_35779,N_34147);
nand U36713 (N_36713,N_34344,N_34134);
nand U36714 (N_36714,N_35976,N_34660);
and U36715 (N_36715,N_35093,N_35161);
xor U36716 (N_36716,N_34738,N_34300);
or U36717 (N_36717,N_35906,N_34600);
xnor U36718 (N_36718,N_34190,N_35874);
nand U36719 (N_36719,N_35762,N_35605);
nand U36720 (N_36720,N_34913,N_34607);
xnor U36721 (N_36721,N_34490,N_35115);
or U36722 (N_36722,N_34768,N_34211);
xor U36723 (N_36723,N_35139,N_34647);
or U36724 (N_36724,N_34626,N_35247);
nor U36725 (N_36725,N_35544,N_34304);
or U36726 (N_36726,N_35936,N_34452);
nand U36727 (N_36727,N_34468,N_35088);
and U36728 (N_36728,N_34787,N_35922);
nand U36729 (N_36729,N_34245,N_35769);
nor U36730 (N_36730,N_34855,N_34741);
xnor U36731 (N_36731,N_34615,N_35672);
nand U36732 (N_36732,N_35920,N_35355);
and U36733 (N_36733,N_35414,N_34339);
nand U36734 (N_36734,N_35029,N_35127);
and U36735 (N_36735,N_35696,N_35618);
nand U36736 (N_36736,N_34671,N_35233);
nor U36737 (N_36737,N_34478,N_35835);
xor U36738 (N_36738,N_34727,N_34295);
or U36739 (N_36739,N_35097,N_34653);
or U36740 (N_36740,N_35157,N_35956);
or U36741 (N_36741,N_34604,N_35334);
nand U36742 (N_36742,N_35721,N_35021);
nand U36743 (N_36743,N_34993,N_34742);
nor U36744 (N_36744,N_35467,N_34492);
nor U36745 (N_36745,N_35253,N_35634);
or U36746 (N_36746,N_34386,N_34079);
and U36747 (N_36747,N_35929,N_35487);
nand U36748 (N_36748,N_34474,N_35437);
xor U36749 (N_36749,N_34972,N_34022);
or U36750 (N_36750,N_35849,N_34103);
and U36751 (N_36751,N_35543,N_34113);
nand U36752 (N_36752,N_35732,N_35490);
or U36753 (N_36753,N_35655,N_34185);
nand U36754 (N_36754,N_35112,N_35868);
nor U36755 (N_36755,N_35997,N_34558);
or U36756 (N_36756,N_35377,N_34659);
and U36757 (N_36757,N_34059,N_35826);
nor U36758 (N_36758,N_35802,N_35847);
or U36759 (N_36759,N_34383,N_34679);
and U36760 (N_36760,N_35937,N_35176);
nor U36761 (N_36761,N_35877,N_35607);
and U36762 (N_36762,N_34566,N_35719);
nor U36763 (N_36763,N_35423,N_35429);
xor U36764 (N_36764,N_35844,N_35071);
nand U36765 (N_36765,N_35168,N_34846);
nand U36766 (N_36766,N_34067,N_34271);
nor U36767 (N_36767,N_35028,N_34771);
and U36768 (N_36768,N_35313,N_34075);
or U36769 (N_36769,N_35121,N_35426);
or U36770 (N_36770,N_34675,N_35354);
nor U36771 (N_36771,N_35031,N_34128);
or U36772 (N_36772,N_35138,N_35813);
nor U36773 (N_36773,N_35062,N_34900);
nand U36774 (N_36774,N_35255,N_35815);
xor U36775 (N_36775,N_35181,N_34765);
xnor U36776 (N_36776,N_34488,N_34456);
nand U36777 (N_36777,N_35147,N_34960);
nor U36778 (N_36778,N_35172,N_34764);
nor U36779 (N_36779,N_35918,N_34943);
or U36780 (N_36780,N_35223,N_34351);
xor U36781 (N_36781,N_35265,N_35033);
or U36782 (N_36782,N_34511,N_34722);
and U36783 (N_36783,N_34239,N_34439);
xor U36784 (N_36784,N_35215,N_34634);
nor U36785 (N_36785,N_34286,N_34786);
and U36786 (N_36786,N_34830,N_34975);
or U36787 (N_36787,N_34162,N_34460);
and U36788 (N_36788,N_35932,N_35503);
and U36789 (N_36789,N_34663,N_35491);
or U36790 (N_36790,N_34849,N_34410);
nor U36791 (N_36791,N_35593,N_34920);
and U36792 (N_36792,N_35422,N_34667);
and U36793 (N_36793,N_34910,N_34227);
or U36794 (N_36794,N_35585,N_35306);
xnor U36795 (N_36795,N_35232,N_35269);
xor U36796 (N_36796,N_35240,N_34749);
and U36797 (N_36797,N_35391,N_35065);
and U36798 (N_36798,N_35959,N_35782);
nand U36799 (N_36799,N_34758,N_34760);
xnor U36800 (N_36800,N_34081,N_35566);
nor U36801 (N_36801,N_35130,N_35352);
and U36802 (N_36802,N_35222,N_35400);
nand U36803 (N_36803,N_34175,N_34066);
xnor U36804 (N_36804,N_35685,N_34408);
nand U36805 (N_36805,N_35080,N_35773);
nand U36806 (N_36806,N_34114,N_34155);
xor U36807 (N_36807,N_34069,N_35502);
nor U36808 (N_36808,N_35864,N_34970);
nor U36809 (N_36809,N_35103,N_34087);
xnor U36810 (N_36810,N_35761,N_34125);
nor U36811 (N_36811,N_35682,N_34767);
nand U36812 (N_36812,N_35389,N_35061);
xor U36813 (N_36813,N_35412,N_35040);
xor U36814 (N_36814,N_34531,N_35919);
nand U36815 (N_36815,N_35189,N_35582);
and U36816 (N_36816,N_35228,N_35458);
or U36817 (N_36817,N_34049,N_35572);
xor U36818 (N_36818,N_34397,N_34899);
and U36819 (N_36819,N_35057,N_35462);
xnor U36820 (N_36820,N_35182,N_35704);
nand U36821 (N_36821,N_34687,N_34512);
or U36822 (N_36822,N_35911,N_35738);
or U36823 (N_36823,N_34682,N_35701);
nor U36824 (N_36824,N_35318,N_35671);
nand U36825 (N_36825,N_34894,N_34939);
nand U36826 (N_36826,N_35644,N_35170);
xnor U36827 (N_36827,N_35117,N_35098);
xnor U36828 (N_36828,N_35768,N_34525);
and U36829 (N_36829,N_34034,N_34751);
nor U36830 (N_36830,N_34310,N_35882);
nand U36831 (N_36831,N_35184,N_35863);
or U36832 (N_36832,N_34957,N_34074);
or U36833 (N_36833,N_34714,N_34952);
xnor U36834 (N_36834,N_35554,N_34624);
nor U36835 (N_36835,N_35861,N_34877);
xor U36836 (N_36836,N_35807,N_34073);
nor U36837 (N_36837,N_35650,N_34699);
or U36838 (N_36838,N_35488,N_35568);
xor U36839 (N_36839,N_35960,N_34737);
and U36840 (N_36840,N_34875,N_35551);
and U36841 (N_36841,N_34356,N_34794);
or U36842 (N_36842,N_34149,N_34230);
xor U36843 (N_36843,N_34798,N_34222);
nor U36844 (N_36844,N_34585,N_35116);
xor U36845 (N_36845,N_34654,N_34023);
nor U36846 (N_36846,N_34072,N_34698);
and U36847 (N_36847,N_35122,N_34991);
and U36848 (N_36848,N_34324,N_34937);
or U36849 (N_36849,N_35941,N_35438);
xor U36850 (N_36850,N_34917,N_35985);
and U36851 (N_36851,N_35049,N_34570);
nor U36852 (N_36852,N_34399,N_35466);
xnor U36853 (N_36853,N_34032,N_34921);
nor U36854 (N_36854,N_34925,N_35096);
or U36855 (N_36855,N_34835,N_35238);
or U36856 (N_36856,N_34443,N_35955);
or U36857 (N_36857,N_34163,N_35763);
or U36858 (N_36858,N_35653,N_35750);
xnor U36859 (N_36859,N_34506,N_35547);
xnor U36860 (N_36860,N_35366,N_34275);
nand U36861 (N_36861,N_35119,N_35330);
xor U36862 (N_36862,N_35661,N_34052);
xnor U36863 (N_36863,N_34781,N_34772);
nor U36864 (N_36864,N_34543,N_34997);
nor U36865 (N_36865,N_35282,N_35702);
nand U36866 (N_36866,N_35656,N_34756);
or U36867 (N_36867,N_35535,N_34818);
nor U36868 (N_36868,N_35464,N_35641);
nor U36869 (N_36869,N_34318,N_34429);
and U36870 (N_36870,N_34260,N_35983);
xor U36871 (N_36871,N_34690,N_34996);
and U36872 (N_36872,N_34209,N_34873);
nor U36873 (N_36873,N_35338,N_35876);
and U36874 (N_36874,N_34144,N_35012);
xnor U36875 (N_36875,N_34581,N_34782);
xor U36876 (N_36876,N_34480,N_34466);
xor U36877 (N_36877,N_34455,N_35183);
nand U36878 (N_36878,N_34076,N_34961);
nor U36879 (N_36879,N_34719,N_34620);
nor U36880 (N_36880,N_35878,N_35009);
and U36881 (N_36881,N_35791,N_35036);
or U36882 (N_36882,N_35987,N_34640);
nand U36883 (N_36883,N_35045,N_35760);
xor U36884 (N_36884,N_35660,N_34796);
nor U36885 (N_36885,N_35737,N_35131);
nor U36886 (N_36886,N_35639,N_35526);
or U36887 (N_36887,N_34632,N_34567);
or U36888 (N_36888,N_34206,N_35796);
nor U36889 (N_36889,N_35341,N_35907);
nor U36890 (N_36890,N_34496,N_35008);
and U36891 (N_36891,N_34471,N_34539);
xor U36892 (N_36892,N_34526,N_34311);
nor U36893 (N_36893,N_35842,N_35382);
nor U36894 (N_36894,N_34821,N_35891);
or U36895 (N_36895,N_34020,N_34385);
or U36896 (N_36896,N_34940,N_34946);
xnor U36897 (N_36897,N_35673,N_35140);
nand U36898 (N_36898,N_34482,N_34874);
nand U36899 (N_36899,N_34990,N_35175);
xnor U36900 (N_36900,N_34178,N_34210);
xor U36901 (N_36901,N_34791,N_35010);
nor U36902 (N_36902,N_35899,N_35178);
and U36903 (N_36903,N_34194,N_34195);
xor U36904 (N_36904,N_34238,N_34644);
and U36905 (N_36905,N_34349,N_34352);
nor U36906 (N_36906,N_35160,N_34731);
and U36907 (N_36907,N_35578,N_34521);
and U36908 (N_36908,N_34462,N_35947);
or U36909 (N_36909,N_35789,N_35285);
nor U36910 (N_36910,N_35388,N_34766);
nor U36911 (N_36911,N_34379,N_34350);
nor U36912 (N_36912,N_34406,N_35867);
nor U36913 (N_36913,N_34777,N_35961);
nand U36914 (N_36914,N_35841,N_35385);
or U36915 (N_36915,N_34078,N_34054);
and U36916 (N_36916,N_34335,N_34701);
xnor U36917 (N_36917,N_34006,N_35435);
nand U36918 (N_36918,N_34876,N_34578);
or U36919 (N_36919,N_35766,N_35263);
nor U36920 (N_36920,N_34534,N_35406);
nor U36921 (N_36921,N_35733,N_34160);
xnor U36922 (N_36922,N_35552,N_34532);
or U36923 (N_36923,N_34734,N_35376);
xor U36924 (N_36924,N_35201,N_35859);
and U36925 (N_36925,N_34550,N_34519);
xor U36926 (N_36926,N_34056,N_35778);
nand U36927 (N_36927,N_34942,N_34014);
nor U36928 (N_36928,N_34962,N_35301);
nor U36929 (N_36929,N_35000,N_34170);
or U36930 (N_36930,N_35817,N_34853);
nand U36931 (N_36931,N_35771,N_35362);
xnor U36932 (N_36932,N_34847,N_34621);
nor U36933 (N_36933,N_35749,N_34414);
or U36934 (N_36934,N_35480,N_35880);
or U36935 (N_36935,N_34387,N_34108);
xor U36936 (N_36936,N_35039,N_34467);
nand U36937 (N_36937,N_35640,N_34107);
and U36938 (N_36938,N_34365,N_35335);
nor U36939 (N_36939,N_35837,N_35089);
nor U36940 (N_36940,N_35166,N_34590);
nand U36941 (N_36941,N_34619,N_34122);
nor U36942 (N_36942,N_34868,N_34253);
and U36943 (N_36943,N_35968,N_34044);
and U36944 (N_36944,N_34822,N_34815);
nor U36945 (N_36945,N_34575,N_34258);
xor U36946 (N_36946,N_34204,N_34236);
nor U36947 (N_36947,N_34842,N_35689);
or U36948 (N_36948,N_35746,N_34432);
or U36949 (N_36949,N_34790,N_35637);
nand U36950 (N_36950,N_35465,N_34602);
and U36951 (N_36951,N_34315,N_34546);
nand U36952 (N_36952,N_34440,N_35996);
xnor U36953 (N_36953,N_34501,N_34461);
and U36954 (N_36954,N_34933,N_35361);
nor U36955 (N_36955,N_35734,N_35954);
nor U36956 (N_36956,N_35207,N_34661);
nand U36957 (N_36957,N_34928,N_34264);
or U36958 (N_36958,N_35190,N_34169);
and U36959 (N_36959,N_35850,N_35674);
xor U36960 (N_36960,N_34851,N_35443);
or U36961 (N_36961,N_34542,N_34617);
nor U36962 (N_36962,N_34565,N_35291);
xnor U36963 (N_36963,N_34507,N_35928);
nand U36964 (N_36964,N_34704,N_35651);
xor U36965 (N_36965,N_34872,N_35244);
nor U36966 (N_36966,N_35532,N_35041);
nor U36967 (N_36967,N_35123,N_34984);
xnor U36968 (N_36968,N_34973,N_35085);
nand U36969 (N_36969,N_34433,N_34348);
xnor U36970 (N_36970,N_35022,N_34923);
and U36971 (N_36971,N_34409,N_34088);
nor U36972 (N_36972,N_35597,N_35599);
nand U36973 (N_36973,N_34980,N_34608);
and U36974 (N_36974,N_34463,N_35900);
nor U36975 (N_36975,N_34485,N_35505);
or U36976 (N_36976,N_34333,N_34372);
nor U36977 (N_36977,N_35770,N_34504);
nor U36978 (N_36978,N_35344,N_34470);
nand U36979 (N_36979,N_34603,N_35663);
nand U36980 (N_36980,N_35601,N_35064);
and U36981 (N_36981,N_35857,N_34042);
xor U36982 (N_36982,N_35697,N_35144);
and U36983 (N_36983,N_35327,N_34613);
nand U36984 (N_36984,N_34527,N_35539);
nand U36985 (N_36985,N_35375,N_34241);
nor U36986 (N_36986,N_35744,N_35348);
nor U36987 (N_36987,N_34172,N_34801);
nand U36988 (N_36988,N_34623,N_34217);
nor U36989 (N_36989,N_34421,N_35336);
nor U36990 (N_36990,N_35399,N_34695);
and U36991 (N_36991,N_35515,N_34655);
and U36992 (N_36992,N_34158,N_34297);
or U36993 (N_36993,N_35239,N_35006);
or U36994 (N_36994,N_35810,N_35879);
nand U36995 (N_36995,N_34093,N_35217);
and U36996 (N_36996,N_34986,N_35373);
and U36997 (N_36997,N_35075,N_35331);
xor U36998 (N_36998,N_34810,N_35210);
or U36999 (N_36999,N_34656,N_35950);
or U37000 (N_37000,N_35869,N_34431);
nor U37001 (N_37001,N_35516,N_34197);
or U37002 (N_37002,N_34048,N_35192);
xor U37003 (N_37003,N_35402,N_34742);
and U37004 (N_37004,N_34273,N_35817);
or U37005 (N_37005,N_35703,N_35607);
xor U37006 (N_37006,N_34728,N_34443);
or U37007 (N_37007,N_34557,N_35205);
and U37008 (N_37008,N_34896,N_34024);
xnor U37009 (N_37009,N_34581,N_35423);
and U37010 (N_37010,N_35833,N_34385);
nor U37011 (N_37011,N_34436,N_34281);
xnor U37012 (N_37012,N_35153,N_35943);
nand U37013 (N_37013,N_35602,N_34860);
xnor U37014 (N_37014,N_35230,N_35254);
nand U37015 (N_37015,N_34787,N_35988);
xnor U37016 (N_37016,N_35764,N_35199);
and U37017 (N_37017,N_34721,N_35341);
xnor U37018 (N_37018,N_34096,N_34649);
nor U37019 (N_37019,N_35766,N_35194);
xor U37020 (N_37020,N_35573,N_35207);
nand U37021 (N_37021,N_34050,N_35877);
nand U37022 (N_37022,N_35744,N_34025);
nor U37023 (N_37023,N_35762,N_34415);
nand U37024 (N_37024,N_34620,N_34695);
or U37025 (N_37025,N_35301,N_35338);
and U37026 (N_37026,N_34931,N_35554);
nor U37027 (N_37027,N_34163,N_34259);
xnor U37028 (N_37028,N_35063,N_34443);
nor U37029 (N_37029,N_34548,N_34956);
nor U37030 (N_37030,N_35408,N_34129);
or U37031 (N_37031,N_34873,N_35200);
xnor U37032 (N_37032,N_35418,N_34646);
nor U37033 (N_37033,N_35815,N_35567);
xor U37034 (N_37034,N_34844,N_35083);
nand U37035 (N_37035,N_34813,N_34333);
xnor U37036 (N_37036,N_34456,N_35681);
nor U37037 (N_37037,N_35111,N_34410);
and U37038 (N_37038,N_34900,N_35168);
and U37039 (N_37039,N_34413,N_35453);
xnor U37040 (N_37040,N_35267,N_34570);
and U37041 (N_37041,N_34180,N_34030);
nand U37042 (N_37042,N_34304,N_35672);
or U37043 (N_37043,N_34747,N_34966);
nand U37044 (N_37044,N_35443,N_35350);
or U37045 (N_37045,N_35666,N_35988);
or U37046 (N_37046,N_35335,N_34241);
or U37047 (N_37047,N_34098,N_35103);
and U37048 (N_37048,N_34909,N_34118);
nand U37049 (N_37049,N_35322,N_35525);
nand U37050 (N_37050,N_34984,N_35377);
or U37051 (N_37051,N_34645,N_35526);
and U37052 (N_37052,N_34748,N_35211);
or U37053 (N_37053,N_34949,N_34613);
or U37054 (N_37054,N_34654,N_35741);
and U37055 (N_37055,N_34796,N_35624);
and U37056 (N_37056,N_35308,N_35060);
or U37057 (N_37057,N_34621,N_35902);
or U37058 (N_37058,N_34414,N_35445);
xnor U37059 (N_37059,N_34424,N_35060);
xnor U37060 (N_37060,N_34380,N_34088);
nor U37061 (N_37061,N_34434,N_35468);
xnor U37062 (N_37062,N_35050,N_35926);
xnor U37063 (N_37063,N_35321,N_35604);
nand U37064 (N_37064,N_34676,N_34393);
xor U37065 (N_37065,N_35902,N_35771);
nand U37066 (N_37066,N_34763,N_35729);
xnor U37067 (N_37067,N_35859,N_35307);
xor U37068 (N_37068,N_34667,N_34318);
xnor U37069 (N_37069,N_35024,N_34230);
or U37070 (N_37070,N_34944,N_34673);
or U37071 (N_37071,N_34178,N_35383);
and U37072 (N_37072,N_34311,N_35880);
and U37073 (N_37073,N_34064,N_34570);
nand U37074 (N_37074,N_35968,N_35217);
xnor U37075 (N_37075,N_34217,N_34970);
or U37076 (N_37076,N_34187,N_34156);
nor U37077 (N_37077,N_34885,N_34711);
or U37078 (N_37078,N_35556,N_35981);
nand U37079 (N_37079,N_35688,N_34042);
and U37080 (N_37080,N_34477,N_35591);
nor U37081 (N_37081,N_34276,N_34989);
and U37082 (N_37082,N_34434,N_34391);
or U37083 (N_37083,N_35481,N_34709);
and U37084 (N_37084,N_34010,N_34081);
or U37085 (N_37085,N_35686,N_34315);
and U37086 (N_37086,N_34974,N_35012);
xor U37087 (N_37087,N_35836,N_34433);
nand U37088 (N_37088,N_34530,N_34826);
nand U37089 (N_37089,N_34674,N_34172);
xor U37090 (N_37090,N_34179,N_35143);
nand U37091 (N_37091,N_35814,N_34953);
nand U37092 (N_37092,N_35650,N_34684);
and U37093 (N_37093,N_35524,N_35297);
or U37094 (N_37094,N_35035,N_34180);
or U37095 (N_37095,N_34385,N_34601);
nand U37096 (N_37096,N_35072,N_35095);
nor U37097 (N_37097,N_34726,N_35479);
nor U37098 (N_37098,N_35608,N_35939);
or U37099 (N_37099,N_34115,N_34451);
or U37100 (N_37100,N_35330,N_35466);
nor U37101 (N_37101,N_34190,N_35972);
nand U37102 (N_37102,N_35188,N_35363);
or U37103 (N_37103,N_34329,N_35777);
nor U37104 (N_37104,N_34520,N_34704);
and U37105 (N_37105,N_34032,N_34780);
xnor U37106 (N_37106,N_35733,N_35070);
or U37107 (N_37107,N_34204,N_35358);
nor U37108 (N_37108,N_34940,N_35441);
or U37109 (N_37109,N_34896,N_34258);
nand U37110 (N_37110,N_34491,N_34678);
nand U37111 (N_37111,N_34553,N_35953);
nand U37112 (N_37112,N_35980,N_34514);
and U37113 (N_37113,N_34315,N_35087);
and U37114 (N_37114,N_35787,N_35110);
nor U37115 (N_37115,N_35273,N_35048);
and U37116 (N_37116,N_34339,N_34568);
xnor U37117 (N_37117,N_34568,N_34172);
nand U37118 (N_37118,N_35653,N_34036);
nor U37119 (N_37119,N_35801,N_35620);
xnor U37120 (N_37120,N_34447,N_34429);
nor U37121 (N_37121,N_35313,N_35631);
xor U37122 (N_37122,N_34708,N_35592);
nor U37123 (N_37123,N_34960,N_34242);
nor U37124 (N_37124,N_34260,N_34115);
nor U37125 (N_37125,N_35846,N_34218);
and U37126 (N_37126,N_35434,N_35857);
xnor U37127 (N_37127,N_35791,N_34852);
nor U37128 (N_37128,N_34621,N_35668);
or U37129 (N_37129,N_35238,N_35101);
or U37130 (N_37130,N_34408,N_35273);
xnor U37131 (N_37131,N_34162,N_34055);
nor U37132 (N_37132,N_34277,N_35188);
nor U37133 (N_37133,N_34032,N_35286);
xnor U37134 (N_37134,N_34904,N_35697);
and U37135 (N_37135,N_34920,N_35479);
and U37136 (N_37136,N_35877,N_35976);
or U37137 (N_37137,N_35891,N_34310);
nand U37138 (N_37138,N_34825,N_34980);
nand U37139 (N_37139,N_35464,N_34311);
and U37140 (N_37140,N_35630,N_34353);
nor U37141 (N_37141,N_34601,N_35573);
and U37142 (N_37142,N_35340,N_34246);
nor U37143 (N_37143,N_34008,N_35303);
nor U37144 (N_37144,N_35219,N_35091);
nor U37145 (N_37145,N_35103,N_35148);
nand U37146 (N_37146,N_34361,N_35338);
and U37147 (N_37147,N_35649,N_34424);
or U37148 (N_37148,N_34113,N_35219);
xnor U37149 (N_37149,N_35578,N_35710);
and U37150 (N_37150,N_34531,N_34766);
nand U37151 (N_37151,N_34643,N_35910);
nor U37152 (N_37152,N_34256,N_34954);
and U37153 (N_37153,N_34423,N_34131);
nand U37154 (N_37154,N_35947,N_34500);
or U37155 (N_37155,N_35605,N_35897);
and U37156 (N_37156,N_34021,N_35865);
nor U37157 (N_37157,N_35414,N_34228);
and U37158 (N_37158,N_35053,N_34874);
and U37159 (N_37159,N_34299,N_34642);
xnor U37160 (N_37160,N_35767,N_35340);
nor U37161 (N_37161,N_34894,N_35556);
nor U37162 (N_37162,N_34780,N_34166);
or U37163 (N_37163,N_34809,N_34698);
xor U37164 (N_37164,N_35263,N_35306);
nand U37165 (N_37165,N_34262,N_35563);
nand U37166 (N_37166,N_34914,N_35802);
xnor U37167 (N_37167,N_35714,N_34136);
or U37168 (N_37168,N_35001,N_34450);
and U37169 (N_37169,N_34480,N_35327);
and U37170 (N_37170,N_34688,N_34801);
xnor U37171 (N_37171,N_35487,N_35802);
xnor U37172 (N_37172,N_35892,N_34166);
nor U37173 (N_37173,N_35371,N_34619);
nor U37174 (N_37174,N_35390,N_35967);
or U37175 (N_37175,N_34997,N_34221);
or U37176 (N_37176,N_34163,N_34086);
and U37177 (N_37177,N_34782,N_35800);
and U37178 (N_37178,N_34414,N_35471);
or U37179 (N_37179,N_34268,N_35118);
and U37180 (N_37180,N_34806,N_34831);
or U37181 (N_37181,N_34657,N_35178);
nand U37182 (N_37182,N_34603,N_35616);
nand U37183 (N_37183,N_35124,N_34367);
xnor U37184 (N_37184,N_35241,N_35510);
xnor U37185 (N_37185,N_35095,N_35639);
xnor U37186 (N_37186,N_35318,N_34170);
nor U37187 (N_37187,N_34069,N_35118);
and U37188 (N_37188,N_34217,N_34704);
xnor U37189 (N_37189,N_35160,N_35033);
nor U37190 (N_37190,N_35727,N_35731);
xor U37191 (N_37191,N_35443,N_34079);
and U37192 (N_37192,N_35761,N_35510);
and U37193 (N_37193,N_34333,N_34406);
and U37194 (N_37194,N_34057,N_35713);
and U37195 (N_37195,N_34808,N_34429);
nand U37196 (N_37196,N_34355,N_35736);
xor U37197 (N_37197,N_34391,N_35446);
nor U37198 (N_37198,N_35826,N_35504);
and U37199 (N_37199,N_34166,N_35922);
or U37200 (N_37200,N_34722,N_35130);
and U37201 (N_37201,N_34220,N_34908);
or U37202 (N_37202,N_34381,N_35148);
nor U37203 (N_37203,N_34425,N_35468);
nor U37204 (N_37204,N_35531,N_35198);
xnor U37205 (N_37205,N_35579,N_35515);
and U37206 (N_37206,N_35480,N_34157);
or U37207 (N_37207,N_35393,N_34605);
nand U37208 (N_37208,N_35533,N_35090);
nor U37209 (N_37209,N_35933,N_35349);
and U37210 (N_37210,N_35952,N_35527);
nor U37211 (N_37211,N_35061,N_34604);
nor U37212 (N_37212,N_35503,N_34442);
and U37213 (N_37213,N_35518,N_35229);
or U37214 (N_37214,N_34113,N_34112);
xor U37215 (N_37215,N_35398,N_35789);
and U37216 (N_37216,N_35249,N_34572);
nor U37217 (N_37217,N_35626,N_35551);
and U37218 (N_37218,N_35891,N_34566);
xor U37219 (N_37219,N_35447,N_35018);
nand U37220 (N_37220,N_35346,N_35101);
or U37221 (N_37221,N_35570,N_35340);
nor U37222 (N_37222,N_34856,N_34388);
or U37223 (N_37223,N_34151,N_34161);
and U37224 (N_37224,N_34155,N_35449);
or U37225 (N_37225,N_34452,N_35773);
and U37226 (N_37226,N_34806,N_34022);
nand U37227 (N_37227,N_35890,N_34075);
or U37228 (N_37228,N_34818,N_34773);
nor U37229 (N_37229,N_35152,N_35400);
and U37230 (N_37230,N_35222,N_35152);
or U37231 (N_37231,N_35303,N_35998);
xnor U37232 (N_37232,N_34814,N_35573);
or U37233 (N_37233,N_35515,N_35314);
or U37234 (N_37234,N_35477,N_35107);
nor U37235 (N_37235,N_35378,N_35275);
xnor U37236 (N_37236,N_34228,N_35166);
and U37237 (N_37237,N_35535,N_35498);
nand U37238 (N_37238,N_34901,N_35783);
nor U37239 (N_37239,N_34452,N_35436);
xor U37240 (N_37240,N_34949,N_35311);
nor U37241 (N_37241,N_35652,N_35878);
or U37242 (N_37242,N_35203,N_34185);
or U37243 (N_37243,N_35596,N_34082);
nand U37244 (N_37244,N_35884,N_34506);
nor U37245 (N_37245,N_35220,N_35659);
xnor U37246 (N_37246,N_34307,N_35952);
and U37247 (N_37247,N_35556,N_35321);
or U37248 (N_37248,N_35371,N_35773);
or U37249 (N_37249,N_35094,N_34190);
xnor U37250 (N_37250,N_35684,N_35275);
nand U37251 (N_37251,N_35053,N_34893);
or U37252 (N_37252,N_34993,N_35027);
nand U37253 (N_37253,N_34039,N_35092);
and U37254 (N_37254,N_35175,N_34230);
or U37255 (N_37255,N_35356,N_34367);
nor U37256 (N_37256,N_35925,N_34347);
or U37257 (N_37257,N_35142,N_34024);
or U37258 (N_37258,N_35702,N_35845);
nand U37259 (N_37259,N_35297,N_34737);
nand U37260 (N_37260,N_34954,N_35065);
nor U37261 (N_37261,N_34426,N_35166);
and U37262 (N_37262,N_35119,N_35866);
and U37263 (N_37263,N_35269,N_34463);
xnor U37264 (N_37264,N_35854,N_35485);
nand U37265 (N_37265,N_34220,N_35109);
and U37266 (N_37266,N_35732,N_34965);
nand U37267 (N_37267,N_34170,N_34430);
and U37268 (N_37268,N_35007,N_35850);
or U37269 (N_37269,N_34012,N_35693);
nor U37270 (N_37270,N_35708,N_35388);
and U37271 (N_37271,N_34554,N_34093);
nand U37272 (N_37272,N_34144,N_34043);
or U37273 (N_37273,N_34030,N_35651);
nor U37274 (N_37274,N_35649,N_34064);
and U37275 (N_37275,N_35877,N_35920);
nor U37276 (N_37276,N_34508,N_34098);
or U37277 (N_37277,N_34811,N_34378);
and U37278 (N_37278,N_34868,N_34848);
nand U37279 (N_37279,N_35617,N_34497);
or U37280 (N_37280,N_35290,N_34545);
xor U37281 (N_37281,N_34908,N_35151);
nand U37282 (N_37282,N_34762,N_35069);
nor U37283 (N_37283,N_34650,N_34277);
or U37284 (N_37284,N_35039,N_34400);
or U37285 (N_37285,N_35541,N_34012);
or U37286 (N_37286,N_34468,N_35527);
and U37287 (N_37287,N_35781,N_35731);
nand U37288 (N_37288,N_35485,N_35241);
xnor U37289 (N_37289,N_35570,N_34229);
or U37290 (N_37290,N_34187,N_34680);
and U37291 (N_37291,N_34467,N_34907);
nand U37292 (N_37292,N_35644,N_35867);
nor U37293 (N_37293,N_35931,N_34790);
or U37294 (N_37294,N_34416,N_34621);
or U37295 (N_37295,N_34394,N_35141);
nor U37296 (N_37296,N_34527,N_34317);
and U37297 (N_37297,N_34854,N_34252);
or U37298 (N_37298,N_34637,N_34120);
nor U37299 (N_37299,N_35716,N_35025);
or U37300 (N_37300,N_35890,N_34525);
nor U37301 (N_37301,N_35116,N_35186);
xor U37302 (N_37302,N_34908,N_34087);
nor U37303 (N_37303,N_34642,N_34667);
xnor U37304 (N_37304,N_35683,N_35317);
and U37305 (N_37305,N_34332,N_35712);
nand U37306 (N_37306,N_34300,N_34263);
nor U37307 (N_37307,N_35185,N_35484);
or U37308 (N_37308,N_35594,N_35097);
nand U37309 (N_37309,N_35526,N_35457);
xor U37310 (N_37310,N_34317,N_34732);
and U37311 (N_37311,N_35801,N_34176);
nand U37312 (N_37312,N_34195,N_34118);
or U37313 (N_37313,N_35430,N_34102);
and U37314 (N_37314,N_35706,N_35798);
nand U37315 (N_37315,N_34750,N_34359);
or U37316 (N_37316,N_34720,N_35650);
xor U37317 (N_37317,N_35235,N_34419);
nand U37318 (N_37318,N_35987,N_35608);
nand U37319 (N_37319,N_34123,N_34798);
nand U37320 (N_37320,N_34525,N_34504);
nand U37321 (N_37321,N_35261,N_34056);
and U37322 (N_37322,N_35649,N_34377);
or U37323 (N_37323,N_34203,N_34988);
nand U37324 (N_37324,N_35803,N_34272);
xor U37325 (N_37325,N_35536,N_34772);
nor U37326 (N_37326,N_35049,N_35357);
and U37327 (N_37327,N_34543,N_34081);
nand U37328 (N_37328,N_35714,N_35285);
xnor U37329 (N_37329,N_35968,N_35321);
nor U37330 (N_37330,N_35531,N_35625);
nor U37331 (N_37331,N_35656,N_34109);
xnor U37332 (N_37332,N_34600,N_34034);
xnor U37333 (N_37333,N_35914,N_35474);
or U37334 (N_37334,N_34592,N_34331);
xnor U37335 (N_37335,N_34938,N_34624);
and U37336 (N_37336,N_34918,N_34599);
xnor U37337 (N_37337,N_34930,N_35155);
nand U37338 (N_37338,N_34212,N_34053);
or U37339 (N_37339,N_34425,N_34220);
nor U37340 (N_37340,N_34947,N_34712);
xnor U37341 (N_37341,N_34670,N_34487);
and U37342 (N_37342,N_35096,N_34243);
or U37343 (N_37343,N_34958,N_35913);
and U37344 (N_37344,N_35239,N_35029);
nand U37345 (N_37345,N_35640,N_34192);
nand U37346 (N_37346,N_34638,N_34900);
xor U37347 (N_37347,N_34459,N_34107);
nand U37348 (N_37348,N_34843,N_34927);
or U37349 (N_37349,N_35929,N_35701);
nand U37350 (N_37350,N_35057,N_34745);
nand U37351 (N_37351,N_34848,N_34287);
nor U37352 (N_37352,N_34424,N_34846);
and U37353 (N_37353,N_34603,N_35035);
xor U37354 (N_37354,N_34093,N_35191);
or U37355 (N_37355,N_35821,N_34672);
nor U37356 (N_37356,N_35620,N_34921);
or U37357 (N_37357,N_35662,N_35849);
nand U37358 (N_37358,N_34360,N_34154);
nand U37359 (N_37359,N_35507,N_34393);
and U37360 (N_37360,N_35390,N_34371);
or U37361 (N_37361,N_35329,N_34292);
xnor U37362 (N_37362,N_34371,N_35466);
nand U37363 (N_37363,N_35145,N_34726);
and U37364 (N_37364,N_35688,N_34758);
or U37365 (N_37365,N_34816,N_35945);
xnor U37366 (N_37366,N_35975,N_34711);
or U37367 (N_37367,N_35554,N_35527);
xnor U37368 (N_37368,N_35931,N_34924);
xnor U37369 (N_37369,N_34379,N_35614);
xor U37370 (N_37370,N_34364,N_35063);
nor U37371 (N_37371,N_35635,N_35559);
nand U37372 (N_37372,N_34560,N_34640);
or U37373 (N_37373,N_34229,N_35736);
nand U37374 (N_37374,N_34258,N_34980);
nor U37375 (N_37375,N_34924,N_35954);
or U37376 (N_37376,N_35795,N_35039);
nand U37377 (N_37377,N_35897,N_34196);
nor U37378 (N_37378,N_34927,N_35294);
xor U37379 (N_37379,N_35042,N_35259);
nor U37380 (N_37380,N_34156,N_34752);
or U37381 (N_37381,N_35650,N_34642);
xor U37382 (N_37382,N_35786,N_35663);
nand U37383 (N_37383,N_34602,N_35860);
nor U37384 (N_37384,N_34922,N_35595);
or U37385 (N_37385,N_35153,N_34055);
or U37386 (N_37386,N_35292,N_34481);
xnor U37387 (N_37387,N_35718,N_34699);
or U37388 (N_37388,N_34858,N_35582);
nor U37389 (N_37389,N_34926,N_34284);
nand U37390 (N_37390,N_35826,N_35085);
or U37391 (N_37391,N_35313,N_34249);
and U37392 (N_37392,N_35526,N_35829);
nand U37393 (N_37393,N_34047,N_35037);
and U37394 (N_37394,N_34541,N_34107);
nor U37395 (N_37395,N_34239,N_34079);
or U37396 (N_37396,N_34415,N_34987);
nand U37397 (N_37397,N_34561,N_35122);
or U37398 (N_37398,N_35743,N_35166);
xnor U37399 (N_37399,N_34263,N_34392);
or U37400 (N_37400,N_34202,N_34855);
nand U37401 (N_37401,N_34827,N_34942);
and U37402 (N_37402,N_35200,N_35764);
nor U37403 (N_37403,N_34827,N_34805);
nand U37404 (N_37404,N_34261,N_34400);
nor U37405 (N_37405,N_34338,N_35546);
xor U37406 (N_37406,N_34785,N_35441);
nand U37407 (N_37407,N_35638,N_34329);
and U37408 (N_37408,N_34433,N_34077);
nor U37409 (N_37409,N_34727,N_35302);
and U37410 (N_37410,N_34159,N_35191);
nor U37411 (N_37411,N_34693,N_35753);
xor U37412 (N_37412,N_35995,N_34240);
xnor U37413 (N_37413,N_35404,N_34632);
nor U37414 (N_37414,N_34325,N_35650);
xnor U37415 (N_37415,N_34202,N_35450);
or U37416 (N_37416,N_35216,N_34206);
and U37417 (N_37417,N_34548,N_34501);
or U37418 (N_37418,N_35056,N_35629);
nand U37419 (N_37419,N_35001,N_34051);
nand U37420 (N_37420,N_34707,N_35854);
or U37421 (N_37421,N_35110,N_35444);
or U37422 (N_37422,N_34712,N_35387);
nand U37423 (N_37423,N_35995,N_34072);
nor U37424 (N_37424,N_34370,N_34853);
nand U37425 (N_37425,N_35720,N_35341);
nor U37426 (N_37426,N_35613,N_35606);
and U37427 (N_37427,N_34508,N_35826);
nand U37428 (N_37428,N_35540,N_34089);
or U37429 (N_37429,N_35504,N_34393);
or U37430 (N_37430,N_34708,N_34339);
nor U37431 (N_37431,N_35818,N_34675);
nor U37432 (N_37432,N_35643,N_34736);
nand U37433 (N_37433,N_34908,N_34013);
nor U37434 (N_37434,N_35230,N_35496);
and U37435 (N_37435,N_35210,N_34024);
or U37436 (N_37436,N_34058,N_34890);
or U37437 (N_37437,N_34098,N_35630);
xnor U37438 (N_37438,N_34118,N_34084);
xnor U37439 (N_37439,N_35298,N_35426);
and U37440 (N_37440,N_35595,N_34486);
nor U37441 (N_37441,N_34909,N_35993);
nand U37442 (N_37442,N_35079,N_34505);
and U37443 (N_37443,N_35603,N_34617);
nor U37444 (N_37444,N_34776,N_34584);
nand U37445 (N_37445,N_34357,N_35553);
or U37446 (N_37446,N_34467,N_35764);
nor U37447 (N_37447,N_34203,N_34637);
nor U37448 (N_37448,N_34432,N_35662);
nor U37449 (N_37449,N_35014,N_35224);
or U37450 (N_37450,N_35771,N_34294);
xor U37451 (N_37451,N_34312,N_35938);
nand U37452 (N_37452,N_35935,N_35398);
or U37453 (N_37453,N_35427,N_34966);
nor U37454 (N_37454,N_34293,N_34177);
and U37455 (N_37455,N_35747,N_35854);
nor U37456 (N_37456,N_35625,N_35276);
or U37457 (N_37457,N_34365,N_34166);
nand U37458 (N_37458,N_35944,N_34009);
nor U37459 (N_37459,N_35701,N_34298);
nand U37460 (N_37460,N_34247,N_34758);
nor U37461 (N_37461,N_34173,N_35935);
nor U37462 (N_37462,N_34158,N_34424);
xor U37463 (N_37463,N_34137,N_34168);
nand U37464 (N_37464,N_34101,N_35962);
or U37465 (N_37465,N_34452,N_35000);
and U37466 (N_37466,N_34700,N_35111);
or U37467 (N_37467,N_34147,N_35923);
xnor U37468 (N_37468,N_35906,N_34337);
nand U37469 (N_37469,N_35993,N_35253);
and U37470 (N_37470,N_34695,N_34156);
or U37471 (N_37471,N_35346,N_34893);
xor U37472 (N_37472,N_34920,N_34917);
xor U37473 (N_37473,N_35946,N_34853);
nor U37474 (N_37474,N_35631,N_34975);
and U37475 (N_37475,N_34776,N_35313);
or U37476 (N_37476,N_35297,N_34983);
nor U37477 (N_37477,N_34782,N_35351);
xor U37478 (N_37478,N_35381,N_35568);
nor U37479 (N_37479,N_35250,N_35874);
xnor U37480 (N_37480,N_34040,N_35016);
xnor U37481 (N_37481,N_35463,N_34392);
and U37482 (N_37482,N_34956,N_34482);
nand U37483 (N_37483,N_35282,N_34691);
nor U37484 (N_37484,N_34170,N_35225);
and U37485 (N_37485,N_35535,N_34422);
or U37486 (N_37486,N_34902,N_35069);
xnor U37487 (N_37487,N_35462,N_35960);
nor U37488 (N_37488,N_35289,N_34615);
and U37489 (N_37489,N_34496,N_35770);
and U37490 (N_37490,N_35552,N_35184);
nand U37491 (N_37491,N_35267,N_35979);
nand U37492 (N_37492,N_34259,N_35605);
and U37493 (N_37493,N_34243,N_35842);
xnor U37494 (N_37494,N_35963,N_34244);
nand U37495 (N_37495,N_35610,N_35803);
and U37496 (N_37496,N_35722,N_34598);
and U37497 (N_37497,N_35734,N_34708);
and U37498 (N_37498,N_34077,N_35004);
and U37499 (N_37499,N_34584,N_35096);
nor U37500 (N_37500,N_34032,N_35614);
xnor U37501 (N_37501,N_35328,N_34817);
nor U37502 (N_37502,N_35325,N_35697);
nor U37503 (N_37503,N_35919,N_35079);
nor U37504 (N_37504,N_35311,N_35853);
nor U37505 (N_37505,N_34439,N_35216);
and U37506 (N_37506,N_34260,N_35736);
or U37507 (N_37507,N_34791,N_34539);
nor U37508 (N_37508,N_35178,N_34749);
and U37509 (N_37509,N_34206,N_34059);
nand U37510 (N_37510,N_34365,N_34555);
xnor U37511 (N_37511,N_34526,N_34495);
and U37512 (N_37512,N_35378,N_34018);
xor U37513 (N_37513,N_34138,N_35301);
xor U37514 (N_37514,N_35839,N_35012);
nand U37515 (N_37515,N_35418,N_34206);
and U37516 (N_37516,N_35832,N_35720);
nor U37517 (N_37517,N_35343,N_34391);
nand U37518 (N_37518,N_34547,N_34608);
nand U37519 (N_37519,N_34649,N_34844);
nand U37520 (N_37520,N_34254,N_34241);
xnor U37521 (N_37521,N_35833,N_34419);
nand U37522 (N_37522,N_35885,N_34947);
nor U37523 (N_37523,N_34166,N_35864);
and U37524 (N_37524,N_35567,N_34415);
and U37525 (N_37525,N_35682,N_34884);
nand U37526 (N_37526,N_34157,N_34567);
and U37527 (N_37527,N_34993,N_34497);
or U37528 (N_37528,N_35563,N_34251);
nor U37529 (N_37529,N_34472,N_35416);
or U37530 (N_37530,N_35818,N_34356);
or U37531 (N_37531,N_34215,N_35439);
nand U37532 (N_37532,N_34825,N_34971);
xnor U37533 (N_37533,N_34753,N_35751);
or U37534 (N_37534,N_34139,N_35778);
nor U37535 (N_37535,N_34305,N_34003);
and U37536 (N_37536,N_35819,N_34322);
or U37537 (N_37537,N_35021,N_35731);
nor U37538 (N_37538,N_35745,N_35500);
nor U37539 (N_37539,N_35780,N_34087);
or U37540 (N_37540,N_34590,N_35710);
nand U37541 (N_37541,N_34454,N_34201);
xor U37542 (N_37542,N_35957,N_35886);
and U37543 (N_37543,N_35777,N_34677);
and U37544 (N_37544,N_34202,N_35812);
nor U37545 (N_37545,N_35348,N_35252);
xnor U37546 (N_37546,N_35905,N_35294);
xor U37547 (N_37547,N_34377,N_35588);
nor U37548 (N_37548,N_35071,N_34411);
and U37549 (N_37549,N_34090,N_35717);
and U37550 (N_37550,N_35935,N_34044);
xor U37551 (N_37551,N_34314,N_35724);
and U37552 (N_37552,N_34098,N_35982);
xor U37553 (N_37553,N_35009,N_35207);
xor U37554 (N_37554,N_34502,N_35350);
or U37555 (N_37555,N_34104,N_35707);
nor U37556 (N_37556,N_35532,N_34010);
or U37557 (N_37557,N_34068,N_34966);
nor U37558 (N_37558,N_35500,N_34907);
xnor U37559 (N_37559,N_34613,N_35721);
xor U37560 (N_37560,N_35607,N_35200);
nor U37561 (N_37561,N_34520,N_34879);
xnor U37562 (N_37562,N_34482,N_35287);
and U37563 (N_37563,N_35491,N_35911);
nor U37564 (N_37564,N_35050,N_35401);
or U37565 (N_37565,N_35248,N_35318);
or U37566 (N_37566,N_35219,N_34784);
and U37567 (N_37567,N_34455,N_34089);
or U37568 (N_37568,N_35950,N_35427);
xor U37569 (N_37569,N_34798,N_34615);
nor U37570 (N_37570,N_34487,N_35412);
nand U37571 (N_37571,N_35213,N_34780);
xor U37572 (N_37572,N_34048,N_35364);
and U37573 (N_37573,N_35011,N_34383);
nor U37574 (N_37574,N_35678,N_34959);
and U37575 (N_37575,N_34684,N_35954);
or U37576 (N_37576,N_34876,N_34160);
nor U37577 (N_37577,N_34879,N_35127);
xnor U37578 (N_37578,N_34632,N_35875);
xnor U37579 (N_37579,N_34156,N_35180);
nor U37580 (N_37580,N_35785,N_34770);
and U37581 (N_37581,N_34277,N_34160);
xor U37582 (N_37582,N_34630,N_34472);
xnor U37583 (N_37583,N_34289,N_35408);
or U37584 (N_37584,N_35117,N_34918);
or U37585 (N_37585,N_35313,N_35921);
xnor U37586 (N_37586,N_34131,N_34153);
and U37587 (N_37587,N_35295,N_35675);
xor U37588 (N_37588,N_35733,N_34453);
xor U37589 (N_37589,N_34030,N_34572);
and U37590 (N_37590,N_34788,N_35635);
and U37591 (N_37591,N_34333,N_35598);
and U37592 (N_37592,N_34587,N_35587);
nand U37593 (N_37593,N_35260,N_35763);
and U37594 (N_37594,N_34927,N_34446);
and U37595 (N_37595,N_34461,N_34274);
nor U37596 (N_37596,N_34065,N_34584);
and U37597 (N_37597,N_35678,N_35839);
or U37598 (N_37598,N_34112,N_35757);
nor U37599 (N_37599,N_34781,N_34587);
nand U37600 (N_37600,N_34638,N_34559);
nand U37601 (N_37601,N_34032,N_34190);
nand U37602 (N_37602,N_35738,N_35384);
xor U37603 (N_37603,N_35796,N_34819);
nor U37604 (N_37604,N_35839,N_34361);
nand U37605 (N_37605,N_34648,N_35455);
and U37606 (N_37606,N_35107,N_34657);
nand U37607 (N_37607,N_35572,N_35511);
and U37608 (N_37608,N_34674,N_34307);
or U37609 (N_37609,N_35956,N_34020);
nand U37610 (N_37610,N_35835,N_34294);
nor U37611 (N_37611,N_34498,N_34524);
xor U37612 (N_37612,N_34995,N_35867);
xor U37613 (N_37613,N_34000,N_35623);
xnor U37614 (N_37614,N_34138,N_35407);
nor U37615 (N_37615,N_35163,N_34209);
or U37616 (N_37616,N_35799,N_35746);
xor U37617 (N_37617,N_34337,N_35695);
nand U37618 (N_37618,N_35629,N_35461);
nor U37619 (N_37619,N_35253,N_34585);
nor U37620 (N_37620,N_35961,N_35063);
xor U37621 (N_37621,N_35805,N_35019);
xnor U37622 (N_37622,N_34941,N_34989);
nor U37623 (N_37623,N_35449,N_34190);
xnor U37624 (N_37624,N_35313,N_34649);
or U37625 (N_37625,N_34500,N_35653);
nand U37626 (N_37626,N_35523,N_34965);
nand U37627 (N_37627,N_35381,N_35148);
nand U37628 (N_37628,N_35997,N_35285);
xor U37629 (N_37629,N_35127,N_34945);
xnor U37630 (N_37630,N_35631,N_35402);
nor U37631 (N_37631,N_34264,N_34966);
nor U37632 (N_37632,N_34825,N_34942);
nor U37633 (N_37633,N_34729,N_34904);
and U37634 (N_37634,N_35988,N_34889);
and U37635 (N_37635,N_35742,N_35536);
xnor U37636 (N_37636,N_34779,N_34096);
xor U37637 (N_37637,N_35437,N_35575);
nor U37638 (N_37638,N_34950,N_35473);
nor U37639 (N_37639,N_34379,N_35168);
nand U37640 (N_37640,N_35234,N_35098);
nand U37641 (N_37641,N_35606,N_35448);
nor U37642 (N_37642,N_35099,N_34430);
or U37643 (N_37643,N_34494,N_35862);
or U37644 (N_37644,N_35558,N_34464);
nand U37645 (N_37645,N_34841,N_35096);
nand U37646 (N_37646,N_34925,N_34097);
nand U37647 (N_37647,N_35186,N_35637);
xor U37648 (N_37648,N_34525,N_35178);
or U37649 (N_37649,N_35473,N_35985);
and U37650 (N_37650,N_34245,N_35860);
and U37651 (N_37651,N_35850,N_34316);
xnor U37652 (N_37652,N_35068,N_35852);
or U37653 (N_37653,N_35671,N_34877);
nor U37654 (N_37654,N_34093,N_35792);
and U37655 (N_37655,N_34585,N_35044);
xnor U37656 (N_37656,N_35042,N_34599);
xnor U37657 (N_37657,N_34298,N_34636);
nand U37658 (N_37658,N_34744,N_35287);
nand U37659 (N_37659,N_35480,N_34369);
xnor U37660 (N_37660,N_35349,N_35524);
or U37661 (N_37661,N_34120,N_34659);
or U37662 (N_37662,N_34956,N_34188);
xor U37663 (N_37663,N_35636,N_34084);
nor U37664 (N_37664,N_35437,N_35803);
or U37665 (N_37665,N_34594,N_35572);
xor U37666 (N_37666,N_35082,N_35566);
xnor U37667 (N_37667,N_35337,N_34169);
nand U37668 (N_37668,N_34027,N_34748);
or U37669 (N_37669,N_35071,N_35990);
and U37670 (N_37670,N_34447,N_35188);
and U37671 (N_37671,N_34604,N_34061);
xnor U37672 (N_37672,N_34010,N_34084);
nand U37673 (N_37673,N_34000,N_34097);
and U37674 (N_37674,N_35312,N_35876);
nand U37675 (N_37675,N_35035,N_34221);
or U37676 (N_37676,N_34406,N_34847);
xor U37677 (N_37677,N_35047,N_35886);
and U37678 (N_37678,N_34119,N_34659);
nand U37679 (N_37679,N_35855,N_35103);
xnor U37680 (N_37680,N_35995,N_35045);
and U37681 (N_37681,N_35473,N_34896);
xor U37682 (N_37682,N_35881,N_35160);
or U37683 (N_37683,N_34985,N_34999);
and U37684 (N_37684,N_35715,N_35004);
or U37685 (N_37685,N_35896,N_35967);
xor U37686 (N_37686,N_34884,N_34887);
xor U37687 (N_37687,N_34180,N_35254);
nand U37688 (N_37688,N_34021,N_35543);
nor U37689 (N_37689,N_35500,N_35414);
nor U37690 (N_37690,N_34947,N_34503);
nor U37691 (N_37691,N_34542,N_34983);
nand U37692 (N_37692,N_34301,N_34432);
nand U37693 (N_37693,N_34538,N_34986);
nand U37694 (N_37694,N_34900,N_34359);
or U37695 (N_37695,N_34279,N_35244);
xnor U37696 (N_37696,N_34944,N_34938);
nand U37697 (N_37697,N_35500,N_34057);
or U37698 (N_37698,N_35942,N_35132);
nor U37699 (N_37699,N_34932,N_34823);
xnor U37700 (N_37700,N_35405,N_35556);
nand U37701 (N_37701,N_35346,N_34326);
and U37702 (N_37702,N_34081,N_35577);
nand U37703 (N_37703,N_35157,N_34707);
nor U37704 (N_37704,N_35528,N_34145);
or U37705 (N_37705,N_34254,N_35098);
nand U37706 (N_37706,N_34879,N_34050);
nand U37707 (N_37707,N_35924,N_35994);
xor U37708 (N_37708,N_34770,N_34584);
and U37709 (N_37709,N_35047,N_34110);
xor U37710 (N_37710,N_34114,N_35293);
nand U37711 (N_37711,N_35445,N_35302);
or U37712 (N_37712,N_34713,N_34904);
or U37713 (N_37713,N_35260,N_35333);
nor U37714 (N_37714,N_34926,N_35913);
nand U37715 (N_37715,N_34261,N_35471);
nand U37716 (N_37716,N_35246,N_34767);
and U37717 (N_37717,N_35555,N_35232);
or U37718 (N_37718,N_34514,N_34256);
or U37719 (N_37719,N_35232,N_34865);
and U37720 (N_37720,N_34261,N_34546);
xor U37721 (N_37721,N_34615,N_34980);
and U37722 (N_37722,N_35296,N_34314);
xor U37723 (N_37723,N_35855,N_34306);
or U37724 (N_37724,N_35822,N_34982);
xor U37725 (N_37725,N_35288,N_35953);
or U37726 (N_37726,N_34658,N_34959);
nor U37727 (N_37727,N_34642,N_35598);
nand U37728 (N_37728,N_34502,N_34401);
and U37729 (N_37729,N_35586,N_35676);
and U37730 (N_37730,N_34238,N_35867);
or U37731 (N_37731,N_35664,N_34372);
or U37732 (N_37732,N_34260,N_35691);
nor U37733 (N_37733,N_34026,N_34507);
xor U37734 (N_37734,N_34823,N_35313);
and U37735 (N_37735,N_35907,N_35531);
or U37736 (N_37736,N_35183,N_35907);
xor U37737 (N_37737,N_34458,N_35077);
and U37738 (N_37738,N_35607,N_35400);
nand U37739 (N_37739,N_34135,N_35450);
nand U37740 (N_37740,N_34753,N_35341);
nor U37741 (N_37741,N_34128,N_35727);
nand U37742 (N_37742,N_35142,N_34695);
nand U37743 (N_37743,N_35607,N_34738);
or U37744 (N_37744,N_35852,N_34647);
xor U37745 (N_37745,N_34660,N_34475);
nand U37746 (N_37746,N_35984,N_34957);
nor U37747 (N_37747,N_34224,N_34289);
nor U37748 (N_37748,N_35421,N_34895);
xnor U37749 (N_37749,N_35037,N_34691);
or U37750 (N_37750,N_34020,N_34672);
or U37751 (N_37751,N_35424,N_35203);
nand U37752 (N_37752,N_35000,N_35500);
or U37753 (N_37753,N_35752,N_34302);
nor U37754 (N_37754,N_34861,N_35328);
or U37755 (N_37755,N_34699,N_35328);
xnor U37756 (N_37756,N_35256,N_35039);
and U37757 (N_37757,N_34286,N_35925);
xnor U37758 (N_37758,N_34427,N_34638);
nor U37759 (N_37759,N_35120,N_34709);
or U37760 (N_37760,N_34865,N_34120);
or U37761 (N_37761,N_35225,N_35303);
xnor U37762 (N_37762,N_35138,N_34003);
nor U37763 (N_37763,N_34381,N_35466);
or U37764 (N_37764,N_35005,N_34151);
or U37765 (N_37765,N_35340,N_34240);
or U37766 (N_37766,N_35544,N_35981);
xnor U37767 (N_37767,N_34336,N_34538);
and U37768 (N_37768,N_35840,N_34493);
nand U37769 (N_37769,N_34814,N_34667);
nor U37770 (N_37770,N_34170,N_35267);
nor U37771 (N_37771,N_35289,N_35669);
xnor U37772 (N_37772,N_35463,N_34240);
nand U37773 (N_37773,N_35484,N_35538);
nand U37774 (N_37774,N_34953,N_34012);
nand U37775 (N_37775,N_34299,N_35906);
and U37776 (N_37776,N_34888,N_35000);
nand U37777 (N_37777,N_35944,N_34243);
nand U37778 (N_37778,N_35027,N_34291);
and U37779 (N_37779,N_34242,N_35991);
nor U37780 (N_37780,N_34352,N_34726);
nand U37781 (N_37781,N_35590,N_35281);
and U37782 (N_37782,N_34886,N_34545);
and U37783 (N_37783,N_35880,N_34600);
or U37784 (N_37784,N_35917,N_34776);
nand U37785 (N_37785,N_34321,N_35145);
xor U37786 (N_37786,N_35362,N_35521);
and U37787 (N_37787,N_34540,N_35973);
nor U37788 (N_37788,N_34106,N_34264);
xor U37789 (N_37789,N_35272,N_35862);
or U37790 (N_37790,N_34178,N_35550);
xnor U37791 (N_37791,N_34748,N_34646);
or U37792 (N_37792,N_34556,N_35249);
and U37793 (N_37793,N_34919,N_35692);
xor U37794 (N_37794,N_34435,N_34261);
and U37795 (N_37795,N_35521,N_34232);
xor U37796 (N_37796,N_35944,N_35823);
and U37797 (N_37797,N_35466,N_35181);
xor U37798 (N_37798,N_35076,N_35563);
nand U37799 (N_37799,N_35769,N_34155);
and U37800 (N_37800,N_35394,N_34546);
and U37801 (N_37801,N_34765,N_35018);
nand U37802 (N_37802,N_34940,N_34507);
nand U37803 (N_37803,N_35080,N_34468);
or U37804 (N_37804,N_34320,N_34956);
xor U37805 (N_37805,N_35040,N_34423);
nand U37806 (N_37806,N_34238,N_35750);
xnor U37807 (N_37807,N_34678,N_35850);
nand U37808 (N_37808,N_35017,N_34908);
nand U37809 (N_37809,N_34423,N_35489);
nor U37810 (N_37810,N_34763,N_35361);
and U37811 (N_37811,N_35677,N_35482);
or U37812 (N_37812,N_35707,N_34454);
xor U37813 (N_37813,N_35342,N_34389);
nor U37814 (N_37814,N_34720,N_34723);
nor U37815 (N_37815,N_34075,N_35930);
or U37816 (N_37816,N_34292,N_34646);
nand U37817 (N_37817,N_34439,N_35680);
or U37818 (N_37818,N_34837,N_35773);
nand U37819 (N_37819,N_35196,N_34305);
or U37820 (N_37820,N_35282,N_34874);
and U37821 (N_37821,N_35514,N_35440);
or U37822 (N_37822,N_34492,N_34196);
or U37823 (N_37823,N_35552,N_35961);
nor U37824 (N_37824,N_34187,N_35990);
nor U37825 (N_37825,N_35061,N_35435);
and U37826 (N_37826,N_34622,N_35557);
or U37827 (N_37827,N_35125,N_35467);
xnor U37828 (N_37828,N_35020,N_34171);
xnor U37829 (N_37829,N_35372,N_35621);
xor U37830 (N_37830,N_34530,N_34466);
nand U37831 (N_37831,N_35505,N_34539);
and U37832 (N_37832,N_35876,N_35592);
and U37833 (N_37833,N_35039,N_34231);
and U37834 (N_37834,N_35211,N_34074);
nor U37835 (N_37835,N_35094,N_34608);
or U37836 (N_37836,N_34616,N_35104);
or U37837 (N_37837,N_35208,N_34600);
nand U37838 (N_37838,N_35342,N_35430);
or U37839 (N_37839,N_35342,N_34927);
xnor U37840 (N_37840,N_34433,N_35438);
nand U37841 (N_37841,N_34129,N_34677);
xnor U37842 (N_37842,N_35557,N_35912);
nor U37843 (N_37843,N_35793,N_35534);
or U37844 (N_37844,N_34362,N_35903);
nand U37845 (N_37845,N_35732,N_34461);
xnor U37846 (N_37846,N_35926,N_35982);
nor U37847 (N_37847,N_34827,N_34839);
or U37848 (N_37848,N_34040,N_34195);
xnor U37849 (N_37849,N_34953,N_34689);
and U37850 (N_37850,N_35017,N_35933);
xnor U37851 (N_37851,N_35194,N_34665);
nand U37852 (N_37852,N_34447,N_34845);
or U37853 (N_37853,N_34858,N_34009);
xor U37854 (N_37854,N_34581,N_35218);
or U37855 (N_37855,N_34505,N_34027);
xor U37856 (N_37856,N_35608,N_35561);
nor U37857 (N_37857,N_35358,N_34618);
nand U37858 (N_37858,N_35304,N_34056);
and U37859 (N_37859,N_34991,N_35453);
nor U37860 (N_37860,N_34156,N_35453);
or U37861 (N_37861,N_35123,N_35335);
or U37862 (N_37862,N_34271,N_35567);
nor U37863 (N_37863,N_34529,N_34954);
and U37864 (N_37864,N_34082,N_35077);
nand U37865 (N_37865,N_35588,N_34899);
nand U37866 (N_37866,N_35580,N_35105);
xor U37867 (N_37867,N_35739,N_35767);
nor U37868 (N_37868,N_34072,N_35403);
or U37869 (N_37869,N_35423,N_35645);
xor U37870 (N_37870,N_34529,N_34760);
xnor U37871 (N_37871,N_35389,N_34896);
nor U37872 (N_37872,N_35340,N_35106);
xor U37873 (N_37873,N_34029,N_35804);
and U37874 (N_37874,N_34242,N_34641);
or U37875 (N_37875,N_34607,N_34777);
and U37876 (N_37876,N_34633,N_35551);
nand U37877 (N_37877,N_35053,N_34002);
and U37878 (N_37878,N_35071,N_34775);
nand U37879 (N_37879,N_34596,N_34268);
or U37880 (N_37880,N_34746,N_34971);
xor U37881 (N_37881,N_35096,N_34639);
or U37882 (N_37882,N_35214,N_35706);
and U37883 (N_37883,N_34696,N_35515);
nor U37884 (N_37884,N_34713,N_34765);
and U37885 (N_37885,N_34377,N_34242);
nor U37886 (N_37886,N_34016,N_35360);
nor U37887 (N_37887,N_34335,N_34004);
or U37888 (N_37888,N_35239,N_35671);
nand U37889 (N_37889,N_34810,N_35035);
xnor U37890 (N_37890,N_35694,N_35640);
xor U37891 (N_37891,N_34728,N_35282);
and U37892 (N_37892,N_34511,N_35469);
xor U37893 (N_37893,N_35877,N_34470);
nor U37894 (N_37894,N_34418,N_34647);
and U37895 (N_37895,N_35948,N_34090);
nor U37896 (N_37896,N_34212,N_35142);
nor U37897 (N_37897,N_34454,N_35100);
or U37898 (N_37898,N_34517,N_35408);
xor U37899 (N_37899,N_35180,N_34764);
nand U37900 (N_37900,N_34320,N_34061);
nand U37901 (N_37901,N_35531,N_34221);
xnor U37902 (N_37902,N_35376,N_35900);
and U37903 (N_37903,N_34392,N_34021);
xnor U37904 (N_37904,N_35693,N_34821);
nand U37905 (N_37905,N_34413,N_34401);
nand U37906 (N_37906,N_34397,N_35573);
xnor U37907 (N_37907,N_35309,N_34998);
and U37908 (N_37908,N_34625,N_34729);
nor U37909 (N_37909,N_34852,N_35503);
nor U37910 (N_37910,N_34002,N_35464);
xor U37911 (N_37911,N_34347,N_35337);
or U37912 (N_37912,N_34901,N_35428);
nor U37913 (N_37913,N_35638,N_34068);
nor U37914 (N_37914,N_34647,N_34993);
xnor U37915 (N_37915,N_34361,N_34639);
xnor U37916 (N_37916,N_34076,N_35496);
xor U37917 (N_37917,N_35073,N_34705);
xnor U37918 (N_37918,N_35005,N_35654);
nand U37919 (N_37919,N_35388,N_35920);
xnor U37920 (N_37920,N_34204,N_34968);
xor U37921 (N_37921,N_35209,N_35053);
nor U37922 (N_37922,N_35537,N_34440);
nor U37923 (N_37923,N_34751,N_35867);
or U37924 (N_37924,N_34659,N_34389);
and U37925 (N_37925,N_34381,N_34591);
xor U37926 (N_37926,N_34189,N_35276);
nor U37927 (N_37927,N_34323,N_34653);
or U37928 (N_37928,N_35455,N_34094);
and U37929 (N_37929,N_34250,N_35647);
nor U37930 (N_37930,N_34680,N_34490);
nand U37931 (N_37931,N_34694,N_34661);
nand U37932 (N_37932,N_34497,N_35026);
xor U37933 (N_37933,N_35653,N_35914);
and U37934 (N_37934,N_35107,N_35675);
xor U37935 (N_37935,N_35757,N_34948);
nor U37936 (N_37936,N_35122,N_34568);
and U37937 (N_37937,N_34123,N_34380);
xor U37938 (N_37938,N_34411,N_35892);
nand U37939 (N_37939,N_35442,N_35292);
and U37940 (N_37940,N_35757,N_35423);
nand U37941 (N_37941,N_34274,N_34265);
and U37942 (N_37942,N_35557,N_35216);
or U37943 (N_37943,N_35017,N_35862);
xor U37944 (N_37944,N_35875,N_34362);
nand U37945 (N_37945,N_34851,N_35897);
or U37946 (N_37946,N_34407,N_34465);
xor U37947 (N_37947,N_34525,N_34727);
or U37948 (N_37948,N_34626,N_35518);
nor U37949 (N_37949,N_35590,N_35067);
nand U37950 (N_37950,N_34575,N_34376);
and U37951 (N_37951,N_35678,N_35071);
nor U37952 (N_37952,N_35967,N_35163);
nand U37953 (N_37953,N_35510,N_34682);
xnor U37954 (N_37954,N_34127,N_35076);
nand U37955 (N_37955,N_34842,N_35336);
or U37956 (N_37956,N_35906,N_35854);
xor U37957 (N_37957,N_35343,N_35075);
nor U37958 (N_37958,N_35608,N_34603);
nand U37959 (N_37959,N_35701,N_34728);
and U37960 (N_37960,N_34050,N_34241);
or U37961 (N_37961,N_35934,N_35878);
and U37962 (N_37962,N_35543,N_35846);
xnor U37963 (N_37963,N_34611,N_34341);
nor U37964 (N_37964,N_34635,N_35935);
xor U37965 (N_37965,N_34930,N_34365);
nand U37966 (N_37966,N_35604,N_34728);
and U37967 (N_37967,N_34146,N_34963);
or U37968 (N_37968,N_35054,N_35924);
nand U37969 (N_37969,N_34966,N_34509);
xnor U37970 (N_37970,N_34505,N_34593);
nand U37971 (N_37971,N_34755,N_35757);
nand U37972 (N_37972,N_35176,N_35997);
and U37973 (N_37973,N_34655,N_34968);
nor U37974 (N_37974,N_34829,N_34002);
nor U37975 (N_37975,N_34831,N_35521);
xnor U37976 (N_37976,N_34447,N_34211);
and U37977 (N_37977,N_34096,N_34191);
or U37978 (N_37978,N_34969,N_34529);
xor U37979 (N_37979,N_34214,N_35601);
and U37980 (N_37980,N_35612,N_35326);
nand U37981 (N_37981,N_35612,N_34763);
nand U37982 (N_37982,N_34320,N_35178);
nand U37983 (N_37983,N_34723,N_35461);
xnor U37984 (N_37984,N_34676,N_35757);
and U37985 (N_37985,N_35879,N_35706);
nor U37986 (N_37986,N_35837,N_34855);
xnor U37987 (N_37987,N_35737,N_34162);
nor U37988 (N_37988,N_35673,N_35825);
and U37989 (N_37989,N_34609,N_35202);
and U37990 (N_37990,N_34165,N_34730);
xor U37991 (N_37991,N_34733,N_34602);
and U37992 (N_37992,N_35506,N_35638);
nand U37993 (N_37993,N_35655,N_34941);
xor U37994 (N_37994,N_34959,N_34627);
nand U37995 (N_37995,N_34028,N_34808);
and U37996 (N_37996,N_35224,N_35132);
or U37997 (N_37997,N_35422,N_34573);
and U37998 (N_37998,N_34203,N_34038);
nand U37999 (N_37999,N_34260,N_35339);
and U38000 (N_38000,N_36045,N_37261);
nand U38001 (N_38001,N_37367,N_37420);
and U38002 (N_38002,N_36637,N_37195);
xor U38003 (N_38003,N_37755,N_36756);
xnor U38004 (N_38004,N_36215,N_36999);
or U38005 (N_38005,N_36491,N_36110);
nand U38006 (N_38006,N_36681,N_36646);
nor U38007 (N_38007,N_36414,N_37984);
and U38008 (N_38008,N_36722,N_37108);
nand U38009 (N_38009,N_37128,N_36204);
xor U38010 (N_38010,N_37571,N_36453);
and U38011 (N_38011,N_36085,N_36154);
or U38012 (N_38012,N_36140,N_37980);
xnor U38013 (N_38013,N_36362,N_37930);
and U38014 (N_38014,N_37931,N_36957);
nor U38015 (N_38015,N_37474,N_37170);
nand U38016 (N_38016,N_36741,N_36977);
nor U38017 (N_38017,N_36847,N_37310);
and U38018 (N_38018,N_36946,N_36793);
or U38019 (N_38019,N_36114,N_37599);
nand U38020 (N_38020,N_36042,N_36436);
xor U38021 (N_38021,N_37694,N_37027);
xnor U38022 (N_38022,N_37024,N_36472);
nand U38023 (N_38023,N_37088,N_37965);
xor U38024 (N_38024,N_37097,N_37482);
nor U38025 (N_38025,N_36295,N_36032);
or U38026 (N_38026,N_37999,N_37381);
and U38027 (N_38027,N_36508,N_36011);
xnor U38028 (N_38028,N_37217,N_37515);
and U38029 (N_38029,N_37591,N_36787);
or U38030 (N_38030,N_36368,N_36276);
and U38031 (N_38031,N_36222,N_37629);
nand U38032 (N_38032,N_36830,N_37174);
xnor U38033 (N_38033,N_36514,N_37552);
and U38034 (N_38034,N_36408,N_37211);
nor U38035 (N_38035,N_37129,N_37787);
nand U38036 (N_38036,N_36729,N_36937);
and U38037 (N_38037,N_36172,N_36372);
or U38038 (N_38038,N_37825,N_37072);
or U38039 (N_38039,N_36310,N_36713);
nand U38040 (N_38040,N_36346,N_36071);
xnor U38041 (N_38041,N_36649,N_36993);
nand U38042 (N_38042,N_37454,N_37225);
xnor U38043 (N_38043,N_36082,N_36364);
and U38044 (N_38044,N_37146,N_37524);
xor U38045 (N_38045,N_36175,N_37455);
nand U38046 (N_38046,N_37478,N_37350);
and U38047 (N_38047,N_36583,N_37971);
and U38048 (N_38048,N_37255,N_36992);
nand U38049 (N_38049,N_37116,N_37765);
xnor U38050 (N_38050,N_37866,N_37732);
nor U38051 (N_38051,N_36885,N_36166);
and U38052 (N_38052,N_37019,N_37754);
nor U38053 (N_38053,N_37817,N_37460);
xnor U38054 (N_38054,N_37890,N_37569);
nor U38055 (N_38055,N_36487,N_36021);
and U38056 (N_38056,N_37968,N_36200);
nor U38057 (N_38057,N_36780,N_37973);
or U38058 (N_38058,N_36356,N_37775);
or U38059 (N_38059,N_36902,N_37047);
or U38060 (N_38060,N_36018,N_37561);
nor U38061 (N_38061,N_36844,N_36242);
nand U38062 (N_38062,N_36476,N_37250);
xor U38063 (N_38063,N_36568,N_36653);
or U38064 (N_38064,N_37388,N_37810);
nand U38065 (N_38065,N_36046,N_36390);
nand U38066 (N_38066,N_37864,N_36869);
xor U38067 (N_38067,N_36265,N_37034);
and U38068 (N_38068,N_37744,N_36919);
xnor U38069 (N_38069,N_37962,N_37177);
nand U38070 (N_38070,N_36790,N_37149);
xnor U38071 (N_38071,N_36828,N_37394);
xnor U38072 (N_38072,N_37313,N_37992);
nor U38073 (N_38073,N_36973,N_36402);
nor U38074 (N_38074,N_37635,N_37183);
nor U38075 (N_38075,N_37393,N_37945);
and U38076 (N_38076,N_37773,N_37716);
and U38077 (N_38077,N_37323,N_37337);
and U38078 (N_38078,N_36909,N_36229);
nand U38079 (N_38079,N_37574,N_36304);
xnor U38080 (N_38080,N_36299,N_37539);
or U38081 (N_38081,N_36639,N_36631);
xnor U38082 (N_38082,N_37402,N_36578);
xnor U38083 (N_38083,N_36227,N_36111);
xor U38084 (N_38084,N_36438,N_36289);
nand U38085 (N_38085,N_36171,N_36334);
xnor U38086 (N_38086,N_36692,N_37155);
and U38087 (N_38087,N_37481,N_37606);
nand U38088 (N_38088,N_37532,N_36572);
or U38089 (N_38089,N_36378,N_37734);
or U38090 (N_38090,N_36425,N_37054);
nand U38091 (N_38091,N_37657,N_37084);
nand U38092 (N_38092,N_37895,N_36202);
and U38093 (N_38093,N_36412,N_37256);
nand U38094 (N_38094,N_37878,N_36747);
xor U38095 (N_38095,N_36214,N_37760);
xor U38096 (N_38096,N_36084,N_36617);
nor U38097 (N_38097,N_37193,N_36479);
nand U38098 (N_38098,N_37079,N_36879);
and U38099 (N_38099,N_37485,N_37925);
or U38100 (N_38100,N_36317,N_36504);
and U38101 (N_38101,N_37022,N_36002);
nor U38102 (N_38102,N_36056,N_36484);
and U38103 (N_38103,N_37682,N_37926);
nor U38104 (N_38104,N_37633,N_37090);
and U38105 (N_38105,N_37986,N_37498);
and U38106 (N_38106,N_36252,N_36292);
or U38107 (N_38107,N_37206,N_36659);
nor U38108 (N_38108,N_37809,N_36664);
xnor U38109 (N_38109,N_37675,N_36521);
nand U38110 (N_38110,N_37615,N_36584);
nor U38111 (N_38111,N_37082,N_37366);
and U38112 (N_38112,N_37770,N_37939);
xnor U38113 (N_38113,N_37526,N_36181);
nor U38114 (N_38114,N_37351,N_37278);
nor U38115 (N_38115,N_37194,N_37182);
xor U38116 (N_38116,N_36927,N_36591);
nand U38117 (N_38117,N_37187,N_37963);
and U38118 (N_38118,N_36822,N_36314);
or U38119 (N_38119,N_36406,N_36569);
xor U38120 (N_38120,N_37840,N_36093);
xor U38121 (N_38121,N_37941,N_36718);
nor U38122 (N_38122,N_36494,N_36666);
or U38123 (N_38123,N_37602,N_37842);
xor U38124 (N_38124,N_37889,N_37265);
nor U38125 (N_38125,N_37081,N_36709);
and U38126 (N_38126,N_36734,N_36458);
nand U38127 (N_38127,N_37906,N_36636);
nor U38128 (N_38128,N_37588,N_37424);
or U38129 (N_38129,N_37821,N_37184);
xnor U38130 (N_38130,N_36766,N_37766);
nand U38131 (N_38131,N_37975,N_37300);
xor U38132 (N_38132,N_36726,N_36817);
and U38133 (N_38133,N_37336,N_36644);
and U38134 (N_38134,N_36701,N_37163);
nand U38135 (N_38135,N_37510,N_36634);
nor U38136 (N_38136,N_36095,N_37276);
nand U38137 (N_38137,N_36814,N_37859);
or U38138 (N_38138,N_37339,N_36682);
nand U38139 (N_38139,N_37514,N_36542);
and U38140 (N_38140,N_36278,N_37404);
nor U38141 (N_38141,N_36758,N_37290);
nor U38142 (N_38142,N_36001,N_37144);
and U38143 (N_38143,N_36186,N_37502);
xor U38144 (N_38144,N_37249,N_37075);
xor U38145 (N_38145,N_37333,N_36429);
or U38146 (N_38146,N_37969,N_37080);
nand U38147 (N_38147,N_36103,N_36271);
nor U38148 (N_38148,N_36629,N_37724);
nor U38149 (N_38149,N_37593,N_36036);
and U38150 (N_38150,N_37277,N_37143);
nor U38151 (N_38151,N_36336,N_37673);
nand U38152 (N_38152,N_36055,N_37953);
nor U38153 (N_38153,N_37554,N_37726);
or U38154 (N_38154,N_37383,N_37964);
nand U38155 (N_38155,N_37745,N_36164);
nand U38156 (N_38156,N_36267,N_36351);
and U38157 (N_38157,N_37888,N_37033);
nand U38158 (N_38158,N_36220,N_37348);
and U38159 (N_38159,N_36444,N_37066);
xnor U38160 (N_38160,N_36661,N_37230);
or U38161 (N_38161,N_36625,N_36353);
nand U38162 (N_38162,N_37346,N_36795);
and U38163 (N_38163,N_36211,N_36410);
xor U38164 (N_38164,N_37302,N_37352);
nand U38165 (N_38165,N_37533,N_36123);
or U38166 (N_38166,N_36467,N_36481);
and U38167 (N_38167,N_36327,N_37039);
nand U38168 (N_38168,N_37186,N_36802);
or U38169 (N_38169,N_37447,N_36761);
nand U38170 (N_38170,N_37434,N_37709);
nor U38171 (N_38171,N_36740,N_37091);
nor U38172 (N_38172,N_36370,N_36066);
nand U38173 (N_38173,N_37610,N_36539);
nor U38174 (N_38174,N_36344,N_37876);
nand U38175 (N_38175,N_37192,N_36000);
nand U38176 (N_38176,N_37909,N_37305);
and U38177 (N_38177,N_37595,N_37506);
or U38178 (N_38178,N_37518,N_36129);
xor U38179 (N_38179,N_36939,N_37156);
xnor U38180 (N_38180,N_37839,N_37123);
nand U38181 (N_38181,N_37042,N_37259);
or U38182 (N_38182,N_36587,N_36854);
nor U38183 (N_38183,N_36903,N_37897);
nand U38184 (N_38184,N_36759,N_37780);
or U38185 (N_38185,N_36142,N_36024);
and U38186 (N_38186,N_36176,N_36915);
or U38187 (N_38187,N_36030,N_37040);
or U38188 (N_38188,N_37776,N_37469);
or U38189 (N_38189,N_36579,N_37900);
nand U38190 (N_38190,N_37493,N_37213);
and U38191 (N_38191,N_37059,N_37753);
or U38192 (N_38192,N_37873,N_37446);
or U38193 (N_38193,N_36563,N_37672);
nand U38194 (N_38194,N_36449,N_37948);
nand U38195 (N_38195,N_37253,N_36513);
xor U38196 (N_38196,N_36037,N_36050);
nor U38197 (N_38197,N_36357,N_36643);
nor U38198 (N_38198,N_36109,N_36763);
or U38199 (N_38199,N_36485,N_37115);
nand U38200 (N_38200,N_37154,N_36840);
xor U38201 (N_38201,N_37646,N_36609);
xor U38202 (N_38202,N_36423,N_36038);
and U38203 (N_38203,N_37248,N_37718);
nor U38204 (N_38204,N_36654,N_37160);
nand U38205 (N_38205,N_36240,N_36595);
xor U38206 (N_38206,N_37856,N_37004);
nand U38207 (N_38207,N_36363,N_36516);
xnor U38208 (N_38208,N_37916,N_36935);
and U38209 (N_38209,N_37216,N_36034);
and U38210 (N_38210,N_37597,N_37807);
nor U38211 (N_38211,N_36621,N_37152);
or U38212 (N_38212,N_36051,N_36380);
and U38213 (N_38213,N_37911,N_37466);
nor U38214 (N_38214,N_37566,N_37670);
or U38215 (N_38215,N_37262,N_37171);
xnor U38216 (N_38216,N_37204,N_37860);
nand U38217 (N_38217,N_36197,N_37412);
or U38218 (N_38218,N_37285,N_36843);
xnor U38219 (N_38219,N_37689,N_36153);
nor U38220 (N_38220,N_37553,N_36255);
and U38221 (N_38221,N_36886,N_37055);
nand U38222 (N_38222,N_36690,N_37122);
and U38223 (N_38223,N_37391,N_36477);
xor U38224 (N_38224,N_36724,N_37801);
or U38225 (N_38225,N_36074,N_37788);
nand U38226 (N_38226,N_36942,N_36686);
or U38227 (N_38227,N_36248,N_37231);
xor U38228 (N_38228,N_36523,N_36419);
nand U38229 (N_38229,N_37288,N_36801);
and U38230 (N_38230,N_37121,N_37159);
nor U38231 (N_38231,N_36541,N_37451);
xor U38232 (N_38232,N_36850,N_37529);
and U38233 (N_38233,N_37639,N_37432);
nand U38234 (N_38234,N_37835,N_36340);
nor U38235 (N_38235,N_36259,N_36228);
nor U38236 (N_38236,N_36529,N_37795);
or U38237 (N_38237,N_36622,N_36995);
and U38238 (N_38238,N_36628,N_36319);
nor U38239 (N_38239,N_37934,N_37137);
or U38240 (N_38240,N_36023,N_36199);
nor U38241 (N_38241,N_37486,N_37609);
xnor U38242 (N_38242,N_37843,N_36512);
xor U38243 (N_38243,N_36208,N_36520);
nand U38244 (N_38244,N_37794,N_36745);
and U38245 (N_38245,N_36499,N_36096);
xnor U38246 (N_38246,N_36600,N_36088);
nand U38247 (N_38247,N_37935,N_37031);
nand U38248 (N_38248,N_37303,N_37752);
or U38249 (N_38249,N_36465,N_36400);
nor U38250 (N_38250,N_37541,N_36715);
nand U38251 (N_38251,N_36057,N_37101);
xor U38252 (N_38252,N_37737,N_36594);
xnor U38253 (N_38253,N_36656,N_37096);
or U38254 (N_38254,N_36198,N_37731);
and U38255 (N_38255,N_37007,N_37983);
or U38256 (N_38256,N_37865,N_36169);
or U38257 (N_38257,N_37756,N_36565);
xor U38258 (N_38258,N_36302,N_36960);
or U38259 (N_38259,N_37396,N_37060);
xor U38260 (N_38260,N_37601,N_37919);
nor U38261 (N_38261,N_36463,N_37377);
nand U38262 (N_38262,N_36474,N_36126);
nand U38263 (N_38263,N_36853,N_37671);
or U38264 (N_38264,N_37625,N_37407);
and U38265 (N_38265,N_37000,N_36431);
and U38266 (N_38266,N_36280,N_36016);
nand U38267 (N_38267,N_37044,N_36767);
or U38268 (N_38268,N_36501,N_36633);
or U38269 (N_38269,N_37818,N_36270);
nand U38270 (N_38270,N_36752,N_36697);
nor U38271 (N_38271,N_36522,N_37087);
or U38272 (N_38272,N_37100,N_37064);
nor U38273 (N_38273,N_37309,N_37120);
nor U38274 (N_38274,N_37239,N_37789);
and U38275 (N_38275,N_37165,N_36015);
and U38276 (N_38276,N_36810,N_36985);
and U38277 (N_38277,N_36914,N_36792);
and U38278 (N_38278,N_37228,N_36727);
nor U38279 (N_38279,N_37484,N_37470);
and U38280 (N_38280,N_36645,N_37083);
nand U38281 (N_38281,N_36687,N_36978);
and U38282 (N_38282,N_37208,N_37886);
or U38283 (N_38283,N_37373,N_36282);
xor U38284 (N_38284,N_36097,N_37882);
nor U38285 (N_38285,N_37605,N_36857);
xor U38286 (N_38286,N_36389,N_37555);
and U38287 (N_38287,N_37790,N_37497);
nand U38288 (N_38288,N_37932,N_36475);
and U38289 (N_38289,N_36800,N_36861);
nor U38290 (N_38290,N_37612,N_36660);
and U38291 (N_38291,N_36266,N_37178);
xnor U38292 (N_38292,N_37659,N_36760);
nand U38293 (N_38293,N_37589,N_36842);
nand U38294 (N_38294,N_37812,N_36489);
xnor U38295 (N_38295,N_37683,N_37409);
nand U38296 (N_38296,N_37637,N_37870);
nor U38297 (N_38297,N_37858,N_37836);
xnor U38298 (N_38298,N_36789,N_36249);
nand U38299 (N_38299,N_37631,N_36880);
xor U38300 (N_38300,N_36710,N_37769);
or U38301 (N_38301,N_37796,N_36488);
xnor U38302 (N_38302,N_37997,N_37103);
or U38303 (N_38303,N_37320,N_36236);
nand U38304 (N_38304,N_36253,N_36900);
and U38305 (N_38305,N_36768,N_37431);
nor U38306 (N_38306,N_36141,N_36662);
xor U38307 (N_38307,N_36603,N_36026);
or U38308 (N_38308,N_37205,N_36441);
nor U38309 (N_38309,N_37598,N_37862);
nand U38310 (N_38310,N_37824,N_36127);
nand U38311 (N_38311,N_36546,N_37768);
xnor U38312 (N_38312,N_37736,N_36940);
xnor U38313 (N_38313,N_36174,N_37820);
xnor U38314 (N_38314,N_36273,N_37307);
xor U38315 (N_38315,N_36545,N_37777);
and U38316 (N_38316,N_37086,N_37563);
nand U38317 (N_38317,N_36798,N_37778);
nor U38318 (N_38318,N_36531,N_37490);
and U38319 (N_38319,N_37287,N_37767);
and U38320 (N_38320,N_36899,N_36862);
xor U38321 (N_38321,N_36665,N_37219);
and U38322 (N_38322,N_36116,N_37928);
and U38323 (N_38323,N_37762,N_37564);
and U38324 (N_38324,N_37190,N_36673);
nand U38325 (N_38325,N_37480,N_37499);
nand U38326 (N_38326,N_36012,N_37439);
or U38327 (N_38327,N_36388,N_37702);
and U38328 (N_38328,N_36901,N_36401);
nand U38329 (N_38329,N_36361,N_36691);
nor U38330 (N_38330,N_37459,N_37677);
nand U38331 (N_38331,N_37293,N_37372);
xnor U38332 (N_38332,N_37967,N_37369);
nand U38333 (N_38333,N_36807,N_36232);
xnor U38334 (N_38334,N_37326,N_36365);
nor U38335 (N_38335,N_36509,N_36812);
xnor U38336 (N_38336,N_36905,N_36080);
nand U38337 (N_38337,N_36201,N_36139);
nand U38338 (N_38338,N_37981,N_37099);
or U38339 (N_38339,N_37977,N_37135);
nand U38340 (N_38340,N_37330,N_37158);
xnor U38341 (N_38341,N_37666,N_36680);
nor U38342 (N_38342,N_36330,N_36374);
nand U38343 (N_38343,N_37551,N_37511);
and U38344 (N_38344,N_36839,N_37619);
and U38345 (N_38345,N_37397,N_36619);
nor U38346 (N_38346,N_37345,N_37956);
xor U38347 (N_38347,N_36736,N_36497);
or U38348 (N_38348,N_36823,N_36627);
xor U38349 (N_38349,N_37826,N_36031);
xnor U38350 (N_38350,N_36592,N_36067);
nand U38351 (N_38351,N_37210,N_37540);
or U38352 (N_38352,N_37349,N_37245);
or U38353 (N_38353,N_37703,N_37433);
and U38354 (N_38354,N_36316,N_36770);
and U38355 (N_38355,N_37038,N_37644);
xor U38356 (N_38356,N_36290,N_36971);
xnor U38357 (N_38357,N_37133,N_37311);
nand U38358 (N_38358,N_36764,N_36156);
nor U38359 (N_38359,N_36367,N_37200);
nand U38360 (N_38360,N_36998,N_37959);
nand U38361 (N_38361,N_37203,N_36179);
and U38362 (N_38362,N_37126,N_37251);
and U38363 (N_38363,N_37329,N_37001);
xor U38364 (N_38364,N_36415,N_37740);
or U38365 (N_38365,N_36874,N_36818);
or U38366 (N_38366,N_37421,N_36816);
nand U38367 (N_38367,N_36274,N_36268);
nand U38368 (N_38368,N_37359,N_37508);
xnor U38369 (N_38369,N_36315,N_36532);
or U38370 (N_38370,N_36409,N_36205);
xor U38371 (N_38371,N_37600,N_37419);
nand U38372 (N_38372,N_36538,N_37140);
nor U38373 (N_38373,N_37189,N_37415);
and U38374 (N_38374,N_36396,N_37147);
xor U38375 (N_38375,N_36833,N_36554);
or U38376 (N_38376,N_37940,N_37885);
xor U38377 (N_38377,N_36407,N_37636);
or U38378 (N_38378,N_36552,N_37621);
xnor U38379 (N_38379,N_37721,N_37452);
nor U38380 (N_38380,N_36398,N_36948);
nand U38381 (N_38381,N_36308,N_36473);
and U38382 (N_38382,N_36859,N_36122);
nand U38383 (N_38383,N_36872,N_37746);
and U38384 (N_38384,N_36447,N_37869);
or U38385 (N_38385,N_37874,N_37085);
xor U38386 (N_38386,N_37164,N_36968);
and U38387 (N_38387,N_37861,N_36941);
or U38388 (N_38388,N_37223,N_36217);
or U38389 (N_38389,N_36492,N_37281);
xor U38390 (N_38390,N_37378,N_37487);
nor U38391 (N_38391,N_36989,N_37640);
nand U38392 (N_38392,N_36773,N_36470);
nand U38393 (N_38393,N_36178,N_37658);
and U38394 (N_38394,N_37725,N_36496);
xnor U38395 (N_38395,N_37946,N_36642);
nor U38396 (N_38396,N_37527,N_36781);
nor U38397 (N_38397,N_36456,N_37831);
nor U38398 (N_38398,N_37784,N_37802);
nand U38399 (N_38399,N_36348,N_36247);
xor U38400 (N_38400,N_37148,N_36951);
or U38401 (N_38401,N_37009,N_36047);
xnor U38402 (N_38402,N_37656,N_37627);
nor U38403 (N_38403,N_36206,N_36856);
and U38404 (N_38404,N_36029,N_36386);
xor U38405 (N_38405,N_37723,N_37893);
xnor U38406 (N_38406,N_36655,N_36526);
or U38407 (N_38407,N_36755,N_36303);
or U38408 (N_38408,N_37914,N_37834);
nor U38409 (N_38409,N_36917,N_37863);
nor U38410 (N_38410,N_36284,N_36733);
or U38411 (N_38411,N_36984,N_36834);
and U38412 (N_38412,N_36696,N_37390);
xor U38413 (N_38413,N_37500,N_36528);
nor U38414 (N_38414,N_36846,N_37557);
and U38415 (N_38415,N_37845,N_37663);
xnor U38416 (N_38416,N_37318,N_37445);
nor U38417 (N_38417,N_36098,N_36723);
nor U38418 (N_38418,N_37198,N_37476);
or U38419 (N_38419,N_36961,N_36820);
or U38420 (N_38420,N_36519,N_36459);
or U38421 (N_38421,N_36331,N_37495);
xnor U38422 (N_38422,N_37068,N_37581);
nor U38423 (N_38423,N_36525,N_36432);
and U38424 (N_38424,N_37708,N_36213);
and U38425 (N_38425,N_36072,N_37938);
nand U38426 (N_38426,N_37854,N_36451);
or U38427 (N_38427,N_36728,N_37852);
nor U38428 (N_38428,N_37379,N_37783);
and U38429 (N_38429,N_36897,N_36738);
nor U38430 (N_38430,N_37095,N_36369);
or U38431 (N_38431,N_37556,N_36683);
nand U38432 (N_38432,N_36657,N_36375);
nor U38433 (N_38433,N_37584,N_36162);
nor U38434 (N_38434,N_36924,N_36053);
nor U38435 (N_38435,N_36180,N_36354);
xnor U38436 (N_38436,N_36774,N_36866);
and U38437 (N_38437,N_37892,N_36589);
and U38438 (N_38438,N_37395,N_37705);
and U38439 (N_38439,N_36033,N_36712);
and U38440 (N_38440,N_37426,N_36689);
or U38441 (N_38441,N_37618,N_36976);
xnor U38442 (N_38442,N_36549,N_36251);
and U38443 (N_38443,N_36966,N_37757);
nand U38444 (N_38444,N_36829,N_37015);
nor U38445 (N_38445,N_37538,N_36932);
or U38446 (N_38446,N_37667,N_36212);
xnor U38447 (N_38447,N_37713,N_37063);
xor U38448 (N_38448,N_36613,N_37577);
xnor U38449 (N_38449,N_36732,N_37436);
xor U38450 (N_38450,N_36596,N_36813);
xor U38451 (N_38451,N_37803,N_36170);
nor U38452 (N_38452,N_36667,N_37697);
nand U38453 (N_38453,N_36107,N_37271);
nand U38454 (N_38454,N_36860,N_37202);
and U38455 (N_38455,N_36808,N_37234);
or U38456 (N_38456,N_36221,N_37284);
xnor U38457 (N_38457,N_36326,N_37292);
or U38458 (N_38458,N_36272,N_37105);
and U38459 (N_38459,N_37772,N_37651);
or U38460 (N_38460,N_36632,N_37008);
and U38461 (N_38461,N_37833,N_37429);
or U38462 (N_38462,N_36749,N_37544);
nor U38463 (N_38463,N_37449,N_36832);
nor U38464 (N_38464,N_37343,N_37078);
or U38465 (N_38465,N_37037,N_36183);
or U38466 (N_38466,N_37664,N_36837);
nor U38467 (N_38467,N_36720,N_36328);
nor U38468 (N_38468,N_37036,N_37207);
nand U38469 (N_38469,N_37550,N_36158);
xnor U38470 (N_38470,N_36678,N_37653);
nand U38471 (N_38471,N_36851,N_36648);
xnor U38472 (N_38472,N_37496,N_37857);
nor U38473 (N_38473,N_37611,N_36254);
and U38474 (N_38474,N_36063,N_36534);
xnor U38475 (N_38475,N_37418,N_36605);
nand U38476 (N_38476,N_37405,N_36059);
or U38477 (N_38477,N_37884,N_36502);
nor U38478 (N_38478,N_37117,N_37387);
or U38479 (N_38479,N_36865,N_36906);
or U38480 (N_38480,N_37003,N_37414);
nor U38481 (N_38481,N_36944,N_36452);
and U38482 (N_38482,N_37237,N_36742);
and U38483 (N_38483,N_37976,N_36873);
or U38484 (N_38484,N_36855,N_36196);
and U38485 (N_38485,N_36352,N_36577);
nand U38486 (N_38486,N_37173,N_37304);
nor U38487 (N_38487,N_36442,N_37425);
nor U38488 (N_38488,N_37632,N_37603);
nand U38489 (N_38489,N_37501,N_37056);
nand U38490 (N_38490,N_37645,N_37741);
xor U38491 (N_38491,N_36291,N_37844);
xnor U38492 (N_38492,N_37638,N_37920);
nor U38493 (N_38493,N_36553,N_37026);
nand U38494 (N_38494,N_37384,N_37197);
nand U38495 (N_38495,N_37572,N_37012);
and U38496 (N_38496,N_37877,N_37649);
nor U38497 (N_38497,N_36647,N_37504);
and U38498 (N_38498,N_36635,N_37727);
and U38499 (N_38499,N_37238,N_36392);
nand U38500 (N_38500,N_37907,N_37730);
nand U38501 (N_38501,N_36703,N_36604);
xnor U38502 (N_38502,N_36173,N_37848);
nor U38503 (N_38503,N_37950,N_36987);
and U38504 (N_38504,N_36468,N_36663);
and U38505 (N_38505,N_37654,N_36099);
or U38506 (N_38506,N_37815,N_36982);
nor U38507 (N_38507,N_36815,N_37850);
xnor U38508 (N_38508,N_36256,N_36893);
or U38509 (N_38509,N_37479,N_37996);
nor U38510 (N_38510,N_36574,N_37665);
or U38511 (N_38511,N_37560,N_36788);
xor U38512 (N_38512,N_36440,N_37805);
nor U38513 (N_38513,N_36007,N_37295);
and U38514 (N_38514,N_37077,N_36930);
and U38515 (N_38515,N_37542,N_36241);
and U38516 (N_38516,N_36411,N_36209);
or U38517 (N_38517,N_36305,N_36106);
and U38518 (N_38518,N_37512,N_37503);
nand U38519 (N_38519,N_36610,N_37583);
and U38520 (N_38520,N_37030,N_37505);
or U38521 (N_38521,N_36765,N_36246);
and U38522 (N_38522,N_37813,N_37132);
and U38523 (N_38523,N_37947,N_37680);
nand U38524 (N_38524,N_36224,N_36076);
xor U38525 (N_38525,N_37855,N_36791);
nor U38526 (N_38526,N_37722,N_37933);
and U38527 (N_38527,N_36500,N_37720);
nor U38528 (N_38528,N_36043,N_37062);
nand U38529 (N_38529,N_36702,N_37254);
or U38530 (N_38530,N_37578,N_37829);
nor U38531 (N_38531,N_36799,N_37687);
xor U38532 (N_38532,N_37299,N_36561);
or U38533 (N_38533,N_36836,N_37951);
or U38534 (N_38534,N_37520,N_37119);
xor U38535 (N_38535,N_37879,N_37696);
nand U38536 (N_38536,N_36286,N_37822);
or U38537 (N_38537,N_36483,N_36714);
or U38538 (N_38538,N_36347,N_36908);
nand U38539 (N_38539,N_37990,N_36313);
and U38540 (N_38540,N_37294,N_36878);
and U38541 (N_38541,N_37341,N_37240);
xnor U38542 (N_38542,N_36898,N_37715);
nand U38543 (N_38543,N_37761,N_36235);
or U38544 (N_38544,N_36132,N_36543);
or U38545 (N_38545,N_37628,N_37974);
or U38546 (N_38546,N_37018,N_36119);
xnor U38547 (N_38547,N_37525,N_37365);
xnor U38548 (N_38548,N_36730,N_37799);
and U38549 (N_38549,N_37896,N_36890);
or U38550 (N_38550,N_36005,N_37297);
xnor U38551 (N_38551,N_36786,N_37894);
or U38552 (N_38552,N_36434,N_36355);
nor U38553 (N_38553,N_37798,N_37648);
nor U38554 (N_38554,N_37161,N_36366);
or U38555 (N_38555,N_36028,N_37771);
nand U38556 (N_38556,N_36498,N_37991);
nand U38557 (N_38557,N_36339,N_36184);
and U38558 (N_38558,N_36025,N_37806);
nor U38559 (N_38559,N_37576,N_37151);
or U38560 (N_38560,N_36537,N_37347);
nor U38561 (N_38561,N_37534,N_37543);
or U38562 (N_38562,N_37565,N_36762);
and U38563 (N_38563,N_37356,N_36188);
xnor U38564 (N_38564,N_36882,N_36753);
or U38565 (N_38565,N_37389,N_37382);
nor U38566 (N_38566,N_36612,N_37273);
nor U38567 (N_38567,N_36424,N_36877);
or U38568 (N_38568,N_36573,N_37547);
xnor U38569 (N_38569,N_36382,N_37260);
and U38570 (N_38570,N_37269,N_37150);
xnor U38571 (N_38571,N_36108,N_37127);
and U38572 (N_38572,N_37613,N_36699);
xor U38573 (N_38573,N_36580,N_37435);
or U38574 (N_38574,N_37902,N_36849);
nand U38575 (N_38575,N_37558,N_36075);
xnor U38576 (N_38576,N_37399,N_37191);
and U38577 (N_38577,N_37461,N_37617);
and U38578 (N_38578,N_36652,N_37111);
xor U38579 (N_38579,N_37823,N_37489);
xnor U38580 (N_38580,N_36954,N_37181);
and U38581 (N_38581,N_37046,N_36838);
and U38582 (N_38582,N_37995,N_36044);
nand U38583 (N_38583,N_36157,N_36230);
nor U38584 (N_38584,N_37035,N_37357);
xor U38585 (N_38585,N_37188,N_37011);
nor U38586 (N_38586,N_36138,N_36969);
nand U38587 (N_38587,N_36207,N_36146);
nand U38588 (N_38588,N_37494,N_37828);
or U38589 (N_38589,N_36959,N_36490);
nor U38590 (N_38590,N_37942,N_37032);
nand U38591 (N_38591,N_37257,N_36394);
nand U38592 (N_38592,N_36298,N_36450);
nor U38593 (N_38593,N_36926,N_36101);
xor U38594 (N_38594,N_37410,N_36824);
and U38595 (N_38595,N_36991,N_36185);
and U38596 (N_38596,N_37069,N_36933);
and U38597 (N_38597,N_36945,N_36949);
nand U38598 (N_38598,N_37272,N_37408);
and U38599 (N_38599,N_36620,N_36540);
nand U38600 (N_38600,N_37224,N_37647);
nor U38601 (N_38601,N_36471,N_36448);
or U38602 (N_38602,N_37616,N_37471);
xor U38603 (N_38603,N_37041,N_36010);
and U38604 (N_38604,N_36826,N_37898);
nor U38605 (N_38605,N_36717,N_36943);
nor U38606 (N_38606,N_36040,N_37913);
xnor U38607 (N_38607,N_37226,N_36884);
or U38608 (N_38608,N_37690,N_37883);
nand U38609 (N_38609,N_36530,N_37808);
nor U38610 (N_38610,N_37960,N_36754);
nand U38611 (N_38611,N_37104,N_36006);
nand U38612 (N_38612,N_36306,N_36864);
xor U38613 (N_38613,N_36776,N_37846);
or U38614 (N_38614,N_36996,N_37785);
and U38615 (N_38615,N_37903,N_36505);
nand U38616 (N_38616,N_36669,N_36611);
and U38617 (N_38617,N_36779,N_36078);
nand U38618 (N_38618,N_36684,N_37180);
and U38619 (N_38619,N_37630,N_37185);
and U38620 (N_38620,N_37061,N_37464);
nor U38621 (N_38621,N_37328,N_37676);
or U38622 (N_38622,N_37006,N_37291);
nand U38623 (N_38623,N_36060,N_36064);
nand U38624 (N_38624,N_37332,N_36750);
nand U38625 (N_38625,N_37196,N_37908);
and U38626 (N_38626,N_37586,N_36190);
nor U38627 (N_38627,N_36716,N_37957);
and U38628 (N_38628,N_36725,N_36052);
nor U38629 (N_38629,N_36160,N_36677);
nor U38630 (N_38630,N_37523,N_36892);
or U38631 (N_38631,N_36014,N_36022);
and U38632 (N_38632,N_36518,N_37289);
nor U38633 (N_38633,N_37562,N_36708);
nand U38634 (N_38634,N_36803,N_37321);
nor U38635 (N_38635,N_37401,N_37966);
nand U38636 (N_38636,N_37463,N_37791);
or U38637 (N_38637,N_36557,N_37360);
nand U38638 (N_38638,N_37579,N_36556);
xor U38639 (N_38639,N_36626,N_36058);
nor U38640 (N_38640,N_36671,N_36867);
nand U38641 (N_38641,N_37923,N_36559);
or U38642 (N_38642,N_36443,N_36426);
xor U38643 (N_38643,N_37742,N_37441);
or U38644 (N_38644,N_36705,N_37021);
and U38645 (N_38645,N_37620,N_36430);
nor U38646 (N_38646,N_37661,N_37286);
nand U38647 (N_38647,N_37089,N_36383);
nor U38648 (N_38648,N_37342,N_36105);
nor U38649 (N_38649,N_36507,N_37710);
nor U38650 (N_38650,N_36260,N_37314);
nor U38651 (N_38651,N_36601,N_36548);
and U38652 (N_38652,N_37875,N_37222);
or U38653 (N_38653,N_37707,N_37634);
xor U38654 (N_38654,N_37107,N_37472);
xnor U38655 (N_38655,N_37594,N_36962);
and U38656 (N_38656,N_36263,N_37692);
and U38657 (N_38657,N_37747,N_36437);
nor U38658 (N_38658,N_36193,N_36870);
nand U38659 (N_38659,N_36576,N_37456);
nand U38660 (N_38660,N_36068,N_36775);
and U38661 (N_38661,N_37819,N_36145);
nor U38662 (N_38662,N_37199,N_36772);
xor U38663 (N_38663,N_37267,N_36668);
nand U38664 (N_38664,N_36404,N_37954);
or U38665 (N_38665,N_36461,N_36258);
and U38666 (N_38666,N_36182,N_36480);
and U38667 (N_38667,N_37623,N_36257);
nor U38668 (N_38668,N_37937,N_37522);
xnor U38669 (N_38669,N_37728,N_37029);
and U38670 (N_38670,N_36345,N_36135);
nor U38671 (N_38671,N_37958,N_37403);
nand U38672 (N_38672,N_36695,N_37681);
and U38673 (N_38673,N_37363,N_36194);
or U38674 (N_38674,N_36707,N_37020);
or U38675 (N_38675,N_37136,N_37025);
xor U38676 (N_38676,N_37993,N_36003);
nand U38677 (N_38677,N_37301,N_37535);
and U38678 (N_38678,N_37013,N_36420);
nor U38679 (N_38679,N_37901,N_37641);
and U38680 (N_38680,N_36163,N_37699);
or U38681 (N_38681,N_36980,N_36416);
and U38682 (N_38682,N_37134,N_37400);
nor U38683 (N_38683,N_37701,N_36131);
nor U38684 (N_38684,N_37073,N_36785);
nor U38685 (N_38685,N_36054,N_36567);
nor U38686 (N_38686,N_36149,N_36322);
or U38687 (N_38687,N_36638,N_37247);
and U38688 (N_38688,N_37537,N_37340);
nor U38689 (N_38689,N_36210,N_36435);
nand U38690 (N_38690,N_36321,N_36102);
xnor U38691 (N_38691,N_37376,N_37118);
nand U38692 (N_38692,N_37955,N_37131);
xor U38693 (N_38693,N_36936,N_37052);
nand U38694 (N_38694,N_36831,N_36675);
nor U38695 (N_38695,N_36338,N_36809);
and U38696 (N_38696,N_36203,N_37549);
nor U38697 (N_38697,N_36100,N_37918);
or U38698 (N_38698,N_36017,N_36261);
or U38699 (N_38699,N_36972,N_37614);
and U38700 (N_38700,N_37070,N_36506);
xnor U38701 (N_38701,N_37792,N_37872);
nor U38702 (N_38702,N_37043,N_36811);
and U38703 (N_38703,N_37130,N_36744);
nand U38704 (N_38704,N_36269,N_37917);
xnor U38705 (N_38705,N_36464,N_37098);
nor U38706 (N_38706,N_36511,N_37028);
or U38707 (N_38707,N_37465,N_36911);
and U38708 (N_38708,N_37985,N_36841);
and U38709 (N_38709,N_36371,N_36288);
nand U38710 (N_38710,N_37719,N_36881);
xnor U38711 (N_38711,N_37988,N_37624);
nand U38712 (N_38712,N_36337,N_36244);
xnor U38713 (N_38713,N_36349,N_37924);
xor U38714 (N_38714,N_37392,N_37467);
nand U38715 (N_38715,N_37450,N_36397);
nor U38716 (N_38716,N_36806,N_36307);
nand U38717 (N_38717,N_37051,N_36994);
and U38718 (N_38718,N_36916,N_36275);
and U38719 (N_38719,N_36737,N_37678);
and U38720 (N_38720,N_36137,N_36350);
nand U38721 (N_38721,N_37315,N_36929);
or U38722 (N_38722,N_36283,N_37519);
nand U38723 (N_38723,N_37733,N_37094);
xor U38724 (N_38724,N_36094,N_36070);
xor U38725 (N_38725,N_36387,N_36144);
nor U38726 (N_38726,N_36931,N_37910);
or U38727 (N_38727,N_36413,N_37017);
nand U38728 (N_38728,N_37622,N_36921);
or U38729 (N_38729,N_37308,N_37748);
and U38730 (N_38730,N_37509,N_36446);
or U38731 (N_38731,N_36279,N_36165);
nand U38732 (N_38732,N_36570,N_36341);
or U38733 (N_38733,N_36250,N_37982);
nand U38734 (N_38734,N_36039,N_36564);
nand U38735 (N_38735,N_36287,N_36688);
nand U38736 (N_38736,N_37282,N_36297);
nand U38737 (N_38737,N_36533,N_36896);
or U38738 (N_38738,N_37374,N_37749);
and U38739 (N_38739,N_36113,N_37738);
nor U38740 (N_38740,N_36192,N_36237);
nand U38741 (N_38741,N_37804,N_37849);
or U38742 (N_38742,N_37212,N_37331);
xor U38743 (N_38743,N_36167,N_36827);
xnor U38744 (N_38744,N_37488,N_36558);
nor U38745 (N_38745,N_37652,N_36928);
or U38746 (N_38746,N_36958,N_37521);
or U38747 (N_38747,N_37241,N_36997);
xnor U38748 (N_38748,N_37138,N_36333);
nor U38749 (N_38749,N_37319,N_37559);
and U38750 (N_38750,N_37530,N_36041);
or U38751 (N_38751,N_36120,N_36950);
or U38752 (N_38752,N_36887,N_37660);
or U38753 (N_38753,N_37643,N_36399);
nand U38754 (N_38754,N_36148,N_37430);
xor U38755 (N_38755,N_37573,N_37743);
nand U38756 (N_38756,N_37793,N_36393);
nor U38757 (N_38757,N_36225,N_37867);
and U38758 (N_38758,N_37227,N_36588);
nor U38759 (N_38759,N_36524,N_36300);
nor U38760 (N_38760,N_37786,N_36597);
xnor U38761 (N_38761,N_36599,N_37058);
nand U38762 (N_38762,N_36312,N_37545);
nor U38763 (N_38763,N_37057,N_37994);
nand U38764 (N_38764,N_37607,N_36784);
xor U38765 (N_38765,N_36147,N_37325);
and U38766 (N_38766,N_36019,N_37989);
nor U38767 (N_38767,N_36335,N_36794);
xnor U38768 (N_38768,N_36264,N_36226);
nor U38769 (N_38769,N_37354,N_36020);
or U38770 (N_38770,N_37838,N_36796);
nor U38771 (N_38771,N_36986,N_36891);
xnor U38772 (N_38772,N_36560,N_36883);
xnor U38773 (N_38773,N_37507,N_36955);
nand U38774 (N_38774,N_37067,N_37153);
nor U38775 (N_38775,N_36797,N_36925);
nor U38776 (N_38776,N_36585,N_37491);
nand U38777 (N_38777,N_37362,N_36693);
and U38778 (N_38778,N_36782,N_37201);
and U38779 (N_38779,N_36571,N_37814);
and U38780 (N_38780,N_36187,N_36641);
nand U38781 (N_38781,N_37669,N_37458);
and U38782 (N_38782,N_37139,N_37922);
nand U38783 (N_38783,N_37176,N_36965);
nor U38784 (N_38784,N_37936,N_36607);
or U38785 (N_38785,N_37949,N_37344);
nand U38786 (N_38786,N_37442,N_37797);
and U38787 (N_38787,N_36195,N_37076);
xor U38788 (N_38788,N_36698,N_37375);
and U38789 (N_38789,N_37827,N_37110);
or U38790 (N_38790,N_36777,N_36427);
or U38791 (N_38791,N_36035,N_36562);
and U38792 (N_38792,N_36547,N_37853);
nand U38793 (N_38793,N_37475,N_36602);
and U38794 (N_38794,N_36918,N_36460);
or U38795 (N_38795,N_37411,N_37626);
xnor U38796 (N_38796,N_37279,N_36825);
xor U38797 (N_38797,N_36852,N_36863);
nor U38798 (N_38798,N_37157,N_36379);
xnor U38799 (N_38799,N_37546,N_37590);
xor U38800 (N_38800,N_36704,N_36694);
or U38801 (N_38801,N_37868,N_36871);
nor U38802 (N_38802,N_37596,N_36218);
xnor U38803 (N_38803,N_37686,N_36739);
xor U38804 (N_38804,N_37582,N_36598);
or U38805 (N_38805,N_36155,N_36934);
nand U38806 (N_38806,N_37306,N_37175);
xor U38807 (N_38807,N_37168,N_36048);
nand U38808 (N_38808,N_36133,N_36482);
xnor U38809 (N_38809,N_37513,N_36385);
nand U38810 (N_38810,N_36445,N_37871);
nor U38811 (N_38811,N_37468,N_37608);
xnor U38812 (N_38812,N_37912,N_36376);
nor U38813 (N_38813,N_36309,N_37233);
nor U38814 (N_38814,N_37688,N_37243);
nand U38815 (N_38815,N_36360,N_37568);
or U38816 (N_38816,N_37221,N_36168);
nor U38817 (N_38817,N_37048,N_37704);
nor U38818 (N_38818,N_37700,N_36281);
and U38819 (N_38819,N_37444,N_36104);
or U38820 (N_38820,N_37462,N_37016);
nand U38821 (N_38821,N_36342,N_36746);
or U38822 (N_38822,N_36894,N_36952);
and U38823 (N_38823,N_36231,N_37887);
xnor U38824 (N_38824,N_36151,N_37236);
or U38825 (N_38825,N_37528,N_36418);
and U38826 (N_38826,N_37252,N_36130);
nand U38827 (N_38827,N_37172,N_36128);
nor U38828 (N_38828,N_37655,N_36403);
or U38829 (N_38829,N_36277,N_36964);
and U38830 (N_38830,N_36486,N_36670);
nor U38831 (N_38831,N_36536,N_36323);
nand U38832 (N_38832,N_36910,N_37592);
nand U38833 (N_38833,N_37364,N_36630);
and U38834 (N_38834,N_37169,N_36771);
and U38835 (N_38835,N_36783,N_36769);
and U38836 (N_38836,N_37453,N_36325);
xnor U38837 (N_38837,N_37712,N_36658);
nand U38838 (N_38838,N_37782,N_37049);
or U38839 (N_38839,N_36748,N_36301);
nor U38840 (N_38840,N_37927,N_36296);
xnor U38841 (N_38841,N_36081,N_37167);
or U38842 (N_38842,N_36778,N_37642);
nor U38843 (N_38843,N_36819,N_37847);
or U38844 (N_38844,N_36177,N_36079);
or U38845 (N_38845,N_37575,N_36821);
nor U38846 (N_38846,N_36077,N_36324);
nor U38847 (N_38847,N_36967,N_36895);
nand U38848 (N_38848,N_37714,N_36544);
and U38849 (N_38849,N_37880,N_37473);
xnor U38850 (N_38850,N_36092,N_37232);
nand U38851 (N_38851,N_36904,N_37781);
and U38852 (N_38852,N_36651,N_37275);
and U38853 (N_38853,N_37952,N_37112);
nor U38854 (N_38854,N_36606,N_36990);
xnor U38855 (N_38855,N_37915,N_37662);
and U38856 (N_38856,N_37385,N_37371);
nand U38857 (N_38857,N_37280,N_36065);
nand U38858 (N_38858,N_37422,N_37209);
or U38859 (N_38859,N_37979,N_36757);
nand U38860 (N_38860,N_37005,N_37685);
and U38861 (N_38861,N_36845,N_36868);
nor U38862 (N_38862,N_37679,N_36008);
and U38863 (N_38863,N_36115,N_37380);
and U38864 (N_38864,N_36359,N_36858);
xnor U38865 (N_38865,N_36913,N_36421);
nor U38866 (N_38866,N_37691,N_37106);
nand U38867 (N_38867,N_36118,N_36329);
nor U38868 (N_38868,N_37246,N_37215);
or U38869 (N_38869,N_37693,N_36062);
xnor U38870 (N_38870,N_36125,N_36953);
and U38871 (N_38871,N_37516,N_37071);
xor U38872 (N_38872,N_37580,N_36293);
nand U38873 (N_38873,N_37548,N_37440);
or U38874 (N_38874,N_37092,N_37263);
nand U38875 (N_38875,N_36091,N_36134);
nor U38876 (N_38876,N_37604,N_37830);
and U38877 (N_38877,N_36615,N_36083);
nor U38878 (N_38878,N_37904,N_36721);
nor U38879 (N_38879,N_37166,N_36974);
xnor U38880 (N_38880,N_37109,N_36582);
and U38881 (N_38881,N_36294,N_37711);
nor U38882 (N_38882,N_36377,N_36515);
and U38883 (N_38883,N_37220,N_37881);
nor U38884 (N_38884,N_37242,N_37477);
and U38885 (N_38885,N_37125,N_37124);
and U38886 (N_38886,N_37141,N_37102);
or U38887 (N_38887,N_36216,N_37014);
nand U38888 (N_38888,N_36888,N_37706);
xnor U38889 (N_38889,N_36089,N_36358);
nor U38890 (N_38890,N_37361,N_36009);
and U38891 (N_38891,N_36963,N_36835);
xnor U38892 (N_38892,N_37717,N_36495);
xnor U38893 (N_38893,N_36069,N_37739);
or U38894 (N_38894,N_36422,N_36112);
nor U38895 (N_38895,N_36049,N_37764);
nor U38896 (N_38896,N_36527,N_36124);
nand U38897 (N_38897,N_36238,N_37162);
and U38898 (N_38898,N_36907,N_36912);
nand U38899 (N_38899,N_36616,N_36676);
nand U38900 (N_38900,N_36243,N_37457);
nand U38901 (N_38901,N_36731,N_37800);
nand U38902 (N_38902,N_36234,N_36593);
nor U38903 (N_38903,N_37053,N_36245);
xnor U38904 (N_38904,N_37759,N_37517);
xor U38905 (N_38905,N_37338,N_37413);
nand U38906 (N_38906,N_37324,N_37274);
or U38907 (N_38907,N_37978,N_37536);
xor U38908 (N_38908,N_37353,N_37316);
and U38909 (N_38909,N_36189,N_36975);
nor U38910 (N_38910,N_36219,N_37368);
or U38911 (N_38911,N_36027,N_36233);
and U38912 (N_38912,N_36373,N_36640);
nor U38913 (N_38913,N_36575,N_36923);
nand U38914 (N_38914,N_37698,N_37416);
nor U38915 (N_38915,N_37065,N_37438);
or U38916 (N_38916,N_36086,N_36428);
nand U38917 (N_38917,N_37423,N_36439);
or U38918 (N_38918,N_36614,N_36455);
nand U38919 (N_38919,N_36805,N_37386);
or U38920 (N_38920,N_37322,N_36535);
nand U38921 (N_38921,N_37270,N_37045);
xnor U38922 (N_38922,N_37650,N_36700);
xor U38923 (N_38923,N_36938,N_37492);
and U38924 (N_38924,N_36262,N_36143);
and U38925 (N_38925,N_37258,N_36685);
nor U38926 (N_38926,N_36624,N_37905);
xnor U38927 (N_38927,N_37428,N_36586);
nor U38928 (N_38928,N_37312,N_36417);
nand U38929 (N_38929,N_36136,N_36555);
or U38930 (N_38930,N_36804,N_36947);
or U38931 (N_38931,N_36152,N_36674);
xor U38932 (N_38932,N_37816,N_36343);
and U38933 (N_38933,N_37998,N_37406);
nand U38934 (N_38934,N_36711,N_37358);
or U38935 (N_38935,N_36566,N_36061);
and U38936 (N_38936,N_36517,N_36087);
nand U38937 (N_38937,N_36623,N_37987);
nand U38938 (N_38938,N_36381,N_37570);
and U38939 (N_38939,N_37587,N_37235);
or U38940 (N_38940,N_37448,N_37145);
nor U38941 (N_38941,N_37970,N_36510);
xor U38942 (N_38942,N_37750,N_37684);
or U38943 (N_38943,N_37427,N_37296);
or U38944 (N_38944,N_37417,N_36395);
xnor U38945 (N_38945,N_37779,N_36876);
xnor U38946 (N_38946,N_37929,N_37229);
nor U38947 (N_38947,N_36384,N_36159);
nand U38948 (N_38948,N_36875,N_37266);
nand U38949 (N_38949,N_37943,N_36743);
xnor U38950 (N_38950,N_36318,N_37837);
nor U38951 (N_38951,N_37113,N_37370);
or U38952 (N_38952,N_36405,N_37763);
nor U38953 (N_38953,N_37961,N_36466);
nor U38954 (N_38954,N_36550,N_36073);
xor U38955 (N_38955,N_36848,N_36920);
xnor U38956 (N_38956,N_37010,N_37841);
and U38957 (N_38957,N_36590,N_37944);
nor U38958 (N_38958,N_36706,N_36191);
or U38959 (N_38959,N_37437,N_37972);
and U38960 (N_38960,N_36981,N_36970);
or U38961 (N_38961,N_37774,N_36672);
and U38962 (N_38962,N_37244,N_36239);
nor U38963 (N_38963,N_37023,N_36983);
nand U38964 (N_38964,N_36311,N_36922);
or U38965 (N_38965,N_36679,N_36391);
nand U38966 (N_38966,N_36223,N_36988);
and U38967 (N_38967,N_37317,N_37335);
nor U38968 (N_38968,N_37142,N_37483);
nor U38969 (N_38969,N_36493,N_36332);
xor U38970 (N_38970,N_37050,N_36956);
nor U38971 (N_38971,N_37668,N_36117);
nor U38972 (N_38972,N_37327,N_37567);
and U38973 (N_38973,N_36581,N_36469);
nand U38974 (N_38974,N_36751,N_36004);
xnor U38975 (N_38975,N_36454,N_37758);
nor U38976 (N_38976,N_37114,N_36551);
and U38977 (N_38977,N_37735,N_36650);
xor U38978 (N_38978,N_36320,N_36121);
nor U38979 (N_38979,N_37093,N_36285);
or U38980 (N_38980,N_36462,N_37283);
xor U38981 (N_38981,N_36889,N_37398);
or U38982 (N_38982,N_36503,N_36979);
nor U38983 (N_38983,N_37832,N_37218);
or U38984 (N_38984,N_36161,N_37899);
nor U38985 (N_38985,N_37214,N_37695);
nor U38986 (N_38986,N_37891,N_37585);
xor U38987 (N_38987,N_37443,N_37074);
nand U38988 (N_38988,N_36090,N_37531);
nand U38989 (N_38989,N_36735,N_37751);
and U38990 (N_38990,N_37264,N_36608);
xnor U38991 (N_38991,N_37729,N_36433);
or U38992 (N_38992,N_37674,N_37268);
or U38993 (N_38993,N_37811,N_36719);
nor U38994 (N_38994,N_36457,N_37851);
or U38995 (N_38995,N_37179,N_36478);
nand U38996 (N_38996,N_37298,N_37002);
and U38997 (N_38997,N_36618,N_36150);
xor U38998 (N_38998,N_37355,N_37921);
and U38999 (N_38999,N_37334,N_36013);
xor U39000 (N_39000,N_36294,N_36253);
or U39001 (N_39001,N_36508,N_36687);
nor U39002 (N_39002,N_36426,N_37243);
nand U39003 (N_39003,N_36254,N_37312);
nor U39004 (N_39004,N_36289,N_37882);
xor U39005 (N_39005,N_36364,N_36191);
xor U39006 (N_39006,N_36229,N_36609);
or U39007 (N_39007,N_36350,N_37773);
nand U39008 (N_39008,N_36992,N_36084);
or U39009 (N_39009,N_36181,N_36186);
xnor U39010 (N_39010,N_36984,N_37543);
or U39011 (N_39011,N_36286,N_37534);
or U39012 (N_39012,N_36878,N_37631);
or U39013 (N_39013,N_37451,N_37648);
and U39014 (N_39014,N_37013,N_36590);
or U39015 (N_39015,N_36977,N_36538);
nor U39016 (N_39016,N_37535,N_37473);
or U39017 (N_39017,N_37461,N_37046);
nor U39018 (N_39018,N_37779,N_37451);
and U39019 (N_39019,N_36128,N_37989);
xnor U39020 (N_39020,N_36806,N_37160);
or U39021 (N_39021,N_36140,N_37842);
xnor U39022 (N_39022,N_37802,N_37690);
nor U39023 (N_39023,N_36011,N_37162);
nor U39024 (N_39024,N_36479,N_37906);
nor U39025 (N_39025,N_37160,N_37649);
and U39026 (N_39026,N_36402,N_37427);
nor U39027 (N_39027,N_37145,N_36168);
nand U39028 (N_39028,N_37227,N_37573);
xnor U39029 (N_39029,N_37366,N_36090);
or U39030 (N_39030,N_36285,N_36212);
or U39031 (N_39031,N_37147,N_36264);
or U39032 (N_39032,N_36816,N_36914);
xnor U39033 (N_39033,N_36296,N_36612);
nand U39034 (N_39034,N_36766,N_36583);
nand U39035 (N_39035,N_36462,N_37040);
nor U39036 (N_39036,N_36616,N_36775);
nor U39037 (N_39037,N_36334,N_37440);
and U39038 (N_39038,N_36562,N_36679);
nand U39039 (N_39039,N_36842,N_37683);
nor U39040 (N_39040,N_37776,N_37560);
and U39041 (N_39041,N_37999,N_36167);
nor U39042 (N_39042,N_36567,N_36590);
nand U39043 (N_39043,N_37527,N_37873);
xor U39044 (N_39044,N_37212,N_37943);
nand U39045 (N_39045,N_37909,N_36080);
xnor U39046 (N_39046,N_36260,N_36529);
xnor U39047 (N_39047,N_37947,N_36230);
nor U39048 (N_39048,N_37616,N_37672);
nor U39049 (N_39049,N_37292,N_36104);
or U39050 (N_39050,N_36117,N_37284);
and U39051 (N_39051,N_37751,N_37098);
and U39052 (N_39052,N_36792,N_36907);
xnor U39053 (N_39053,N_36792,N_36860);
xnor U39054 (N_39054,N_37838,N_36635);
nand U39055 (N_39055,N_36643,N_36822);
or U39056 (N_39056,N_36798,N_36771);
nand U39057 (N_39057,N_37845,N_36098);
nor U39058 (N_39058,N_36260,N_37929);
and U39059 (N_39059,N_37476,N_37205);
nor U39060 (N_39060,N_37737,N_36158);
and U39061 (N_39061,N_37266,N_37251);
and U39062 (N_39062,N_37455,N_37723);
nand U39063 (N_39063,N_36340,N_37229);
nor U39064 (N_39064,N_37341,N_37527);
xor U39065 (N_39065,N_36794,N_36408);
nand U39066 (N_39066,N_37524,N_37792);
and U39067 (N_39067,N_36892,N_37070);
or U39068 (N_39068,N_37829,N_37731);
xor U39069 (N_39069,N_37600,N_37964);
xor U39070 (N_39070,N_37559,N_37890);
xnor U39071 (N_39071,N_36408,N_36102);
xor U39072 (N_39072,N_37443,N_37184);
nor U39073 (N_39073,N_37193,N_37009);
xnor U39074 (N_39074,N_36410,N_36692);
nand U39075 (N_39075,N_36768,N_37700);
xor U39076 (N_39076,N_37571,N_37624);
nor U39077 (N_39077,N_37814,N_37703);
nand U39078 (N_39078,N_37862,N_36976);
nor U39079 (N_39079,N_36371,N_37680);
nor U39080 (N_39080,N_36853,N_37260);
nor U39081 (N_39081,N_36118,N_36532);
xor U39082 (N_39082,N_36548,N_36750);
xor U39083 (N_39083,N_37223,N_36367);
xor U39084 (N_39084,N_36666,N_37741);
nand U39085 (N_39085,N_37304,N_37680);
nand U39086 (N_39086,N_37297,N_36359);
and U39087 (N_39087,N_36025,N_36109);
xor U39088 (N_39088,N_37356,N_37382);
xor U39089 (N_39089,N_37509,N_36471);
nor U39090 (N_39090,N_36419,N_37856);
nand U39091 (N_39091,N_37213,N_37307);
xor U39092 (N_39092,N_37595,N_37498);
nand U39093 (N_39093,N_36350,N_36112);
xor U39094 (N_39094,N_36878,N_37266);
nor U39095 (N_39095,N_37189,N_36267);
nor U39096 (N_39096,N_36873,N_36179);
nor U39097 (N_39097,N_36630,N_37742);
or U39098 (N_39098,N_36796,N_37971);
nor U39099 (N_39099,N_37914,N_36708);
nor U39100 (N_39100,N_36421,N_37780);
and U39101 (N_39101,N_36215,N_36042);
xor U39102 (N_39102,N_36902,N_37238);
or U39103 (N_39103,N_37173,N_36422);
xnor U39104 (N_39104,N_36729,N_36396);
nand U39105 (N_39105,N_37956,N_36055);
nand U39106 (N_39106,N_37098,N_37420);
nor U39107 (N_39107,N_37833,N_37387);
or U39108 (N_39108,N_36878,N_36798);
xnor U39109 (N_39109,N_36787,N_36478);
nor U39110 (N_39110,N_37226,N_36020);
and U39111 (N_39111,N_36230,N_37289);
or U39112 (N_39112,N_37373,N_36743);
nor U39113 (N_39113,N_36974,N_36953);
or U39114 (N_39114,N_37431,N_36125);
and U39115 (N_39115,N_37934,N_36606);
nor U39116 (N_39116,N_36025,N_37650);
xnor U39117 (N_39117,N_37135,N_37067);
nand U39118 (N_39118,N_36434,N_36814);
or U39119 (N_39119,N_37101,N_37944);
nor U39120 (N_39120,N_36692,N_37279);
nor U39121 (N_39121,N_36835,N_36383);
nor U39122 (N_39122,N_36564,N_37454);
xnor U39123 (N_39123,N_36634,N_36424);
xor U39124 (N_39124,N_36726,N_36389);
nor U39125 (N_39125,N_37316,N_37230);
and U39126 (N_39126,N_36935,N_37765);
xnor U39127 (N_39127,N_36178,N_37018);
and U39128 (N_39128,N_36891,N_36493);
nand U39129 (N_39129,N_36089,N_37229);
and U39130 (N_39130,N_37673,N_36705);
xor U39131 (N_39131,N_37279,N_37282);
xor U39132 (N_39132,N_36285,N_37495);
and U39133 (N_39133,N_36183,N_37654);
or U39134 (N_39134,N_37268,N_36341);
nor U39135 (N_39135,N_36447,N_36910);
and U39136 (N_39136,N_36247,N_37245);
and U39137 (N_39137,N_37995,N_37648);
or U39138 (N_39138,N_36948,N_36904);
nor U39139 (N_39139,N_36779,N_37424);
or U39140 (N_39140,N_37184,N_37714);
xnor U39141 (N_39141,N_36840,N_37656);
and U39142 (N_39142,N_37050,N_36397);
xnor U39143 (N_39143,N_36336,N_37357);
nand U39144 (N_39144,N_37639,N_36387);
and U39145 (N_39145,N_36752,N_36664);
or U39146 (N_39146,N_37904,N_36904);
nand U39147 (N_39147,N_37104,N_36206);
xor U39148 (N_39148,N_37476,N_37799);
or U39149 (N_39149,N_37511,N_37187);
nand U39150 (N_39150,N_36041,N_36564);
nand U39151 (N_39151,N_37911,N_37894);
nand U39152 (N_39152,N_36616,N_37287);
nor U39153 (N_39153,N_36730,N_36749);
xnor U39154 (N_39154,N_37954,N_37338);
or U39155 (N_39155,N_36101,N_36806);
nor U39156 (N_39156,N_37082,N_37337);
xnor U39157 (N_39157,N_37776,N_36406);
nand U39158 (N_39158,N_37953,N_36648);
xnor U39159 (N_39159,N_36098,N_37686);
nor U39160 (N_39160,N_36909,N_37833);
nor U39161 (N_39161,N_37251,N_36537);
and U39162 (N_39162,N_36797,N_36927);
nor U39163 (N_39163,N_37460,N_36593);
nor U39164 (N_39164,N_37774,N_37622);
nand U39165 (N_39165,N_37439,N_37306);
nand U39166 (N_39166,N_37516,N_37811);
nand U39167 (N_39167,N_37415,N_37010);
or U39168 (N_39168,N_36039,N_36244);
nor U39169 (N_39169,N_36621,N_37134);
nand U39170 (N_39170,N_36549,N_37594);
or U39171 (N_39171,N_36366,N_36246);
and U39172 (N_39172,N_37029,N_37445);
xnor U39173 (N_39173,N_36930,N_36061);
and U39174 (N_39174,N_36380,N_37630);
or U39175 (N_39175,N_37787,N_36256);
nand U39176 (N_39176,N_37663,N_36093);
xnor U39177 (N_39177,N_36181,N_37830);
or U39178 (N_39178,N_37579,N_37889);
nor U39179 (N_39179,N_36456,N_36291);
nor U39180 (N_39180,N_37367,N_37630);
nand U39181 (N_39181,N_36829,N_36462);
or U39182 (N_39182,N_36244,N_36486);
xnor U39183 (N_39183,N_36834,N_36701);
xor U39184 (N_39184,N_36769,N_36027);
or U39185 (N_39185,N_36675,N_36080);
nand U39186 (N_39186,N_36620,N_37721);
nand U39187 (N_39187,N_36473,N_36175);
and U39188 (N_39188,N_37033,N_36126);
xnor U39189 (N_39189,N_36851,N_36950);
and U39190 (N_39190,N_36345,N_37684);
or U39191 (N_39191,N_36527,N_36220);
and U39192 (N_39192,N_36716,N_37391);
and U39193 (N_39193,N_37805,N_37932);
nand U39194 (N_39194,N_36993,N_37383);
nor U39195 (N_39195,N_36836,N_37783);
xor U39196 (N_39196,N_36931,N_37382);
or U39197 (N_39197,N_36841,N_36047);
nor U39198 (N_39198,N_36409,N_37205);
and U39199 (N_39199,N_37860,N_36796);
nor U39200 (N_39200,N_36282,N_36804);
or U39201 (N_39201,N_37201,N_37069);
or U39202 (N_39202,N_36735,N_37954);
and U39203 (N_39203,N_36082,N_36287);
and U39204 (N_39204,N_36475,N_36193);
or U39205 (N_39205,N_36180,N_36991);
or U39206 (N_39206,N_37462,N_36376);
or U39207 (N_39207,N_36153,N_36118);
and U39208 (N_39208,N_36880,N_37936);
nor U39209 (N_39209,N_36583,N_37776);
nand U39210 (N_39210,N_37237,N_36116);
nor U39211 (N_39211,N_36196,N_36812);
nor U39212 (N_39212,N_36988,N_37164);
xor U39213 (N_39213,N_36300,N_36977);
nor U39214 (N_39214,N_36775,N_37967);
nand U39215 (N_39215,N_37147,N_37686);
and U39216 (N_39216,N_37972,N_37874);
or U39217 (N_39217,N_37250,N_37914);
xor U39218 (N_39218,N_37507,N_37896);
nand U39219 (N_39219,N_37729,N_37090);
and U39220 (N_39220,N_36251,N_36874);
xnor U39221 (N_39221,N_36479,N_36223);
xnor U39222 (N_39222,N_36908,N_37570);
or U39223 (N_39223,N_37418,N_36828);
and U39224 (N_39224,N_36288,N_37895);
nand U39225 (N_39225,N_37344,N_36526);
nand U39226 (N_39226,N_37245,N_36458);
or U39227 (N_39227,N_36474,N_36150);
xnor U39228 (N_39228,N_36247,N_37559);
xnor U39229 (N_39229,N_37658,N_37218);
nor U39230 (N_39230,N_37352,N_36445);
nor U39231 (N_39231,N_37863,N_36231);
nor U39232 (N_39232,N_36146,N_36029);
xor U39233 (N_39233,N_37597,N_36833);
or U39234 (N_39234,N_36588,N_36091);
nor U39235 (N_39235,N_37383,N_37895);
nor U39236 (N_39236,N_37617,N_36684);
and U39237 (N_39237,N_37172,N_36067);
or U39238 (N_39238,N_36612,N_36033);
nand U39239 (N_39239,N_36732,N_37080);
nor U39240 (N_39240,N_36426,N_37317);
xnor U39241 (N_39241,N_36606,N_36013);
and U39242 (N_39242,N_37722,N_36666);
or U39243 (N_39243,N_37969,N_36849);
and U39244 (N_39244,N_37380,N_36725);
nand U39245 (N_39245,N_37140,N_36342);
and U39246 (N_39246,N_37446,N_37632);
and U39247 (N_39247,N_36578,N_37270);
or U39248 (N_39248,N_37843,N_36386);
and U39249 (N_39249,N_36112,N_36544);
nand U39250 (N_39250,N_36125,N_36188);
or U39251 (N_39251,N_36154,N_36319);
nor U39252 (N_39252,N_36458,N_37701);
xnor U39253 (N_39253,N_37419,N_36669);
xor U39254 (N_39254,N_37078,N_36095);
and U39255 (N_39255,N_36483,N_37735);
nor U39256 (N_39256,N_36319,N_37737);
nand U39257 (N_39257,N_36742,N_37270);
xor U39258 (N_39258,N_36676,N_37556);
xor U39259 (N_39259,N_36933,N_36360);
xor U39260 (N_39260,N_37478,N_36103);
nand U39261 (N_39261,N_37178,N_36969);
nor U39262 (N_39262,N_36732,N_36084);
nor U39263 (N_39263,N_36087,N_37881);
or U39264 (N_39264,N_36043,N_36372);
nor U39265 (N_39265,N_37338,N_37673);
nand U39266 (N_39266,N_37682,N_37302);
and U39267 (N_39267,N_37577,N_37115);
nor U39268 (N_39268,N_37988,N_36656);
nor U39269 (N_39269,N_36208,N_37342);
xnor U39270 (N_39270,N_37908,N_37451);
or U39271 (N_39271,N_37953,N_36382);
and U39272 (N_39272,N_36342,N_36984);
xnor U39273 (N_39273,N_37433,N_37670);
and U39274 (N_39274,N_37894,N_36460);
xnor U39275 (N_39275,N_36012,N_36554);
xnor U39276 (N_39276,N_37734,N_36490);
nor U39277 (N_39277,N_37209,N_36544);
xnor U39278 (N_39278,N_36976,N_36882);
or U39279 (N_39279,N_36059,N_36533);
xor U39280 (N_39280,N_37256,N_37083);
nand U39281 (N_39281,N_37221,N_37622);
or U39282 (N_39282,N_36266,N_37261);
and U39283 (N_39283,N_36214,N_37115);
and U39284 (N_39284,N_36965,N_37602);
or U39285 (N_39285,N_37157,N_36095);
and U39286 (N_39286,N_36368,N_37324);
nand U39287 (N_39287,N_36398,N_36032);
or U39288 (N_39288,N_37195,N_36636);
nor U39289 (N_39289,N_37150,N_37771);
xor U39290 (N_39290,N_36090,N_36462);
and U39291 (N_39291,N_37006,N_37946);
or U39292 (N_39292,N_37144,N_36103);
xor U39293 (N_39293,N_36565,N_37396);
xor U39294 (N_39294,N_37188,N_36212);
nor U39295 (N_39295,N_36394,N_36354);
nor U39296 (N_39296,N_37572,N_37190);
and U39297 (N_39297,N_37486,N_37558);
and U39298 (N_39298,N_36581,N_36519);
nand U39299 (N_39299,N_36552,N_37612);
nand U39300 (N_39300,N_37759,N_37270);
xor U39301 (N_39301,N_36563,N_36100);
and U39302 (N_39302,N_37458,N_37561);
nor U39303 (N_39303,N_36318,N_36384);
nand U39304 (N_39304,N_37529,N_37032);
nand U39305 (N_39305,N_37277,N_37822);
nor U39306 (N_39306,N_36950,N_37598);
nand U39307 (N_39307,N_37671,N_37126);
or U39308 (N_39308,N_37565,N_36016);
and U39309 (N_39309,N_37840,N_37357);
and U39310 (N_39310,N_37503,N_36867);
xor U39311 (N_39311,N_37544,N_37255);
nand U39312 (N_39312,N_37966,N_37555);
nand U39313 (N_39313,N_36578,N_37479);
and U39314 (N_39314,N_36060,N_36091);
nand U39315 (N_39315,N_37221,N_36765);
xor U39316 (N_39316,N_37979,N_37398);
xor U39317 (N_39317,N_37026,N_37447);
nand U39318 (N_39318,N_36411,N_36900);
nand U39319 (N_39319,N_37286,N_37811);
xnor U39320 (N_39320,N_37272,N_36607);
nor U39321 (N_39321,N_37089,N_36818);
and U39322 (N_39322,N_37294,N_37068);
xor U39323 (N_39323,N_36182,N_36810);
or U39324 (N_39324,N_36273,N_36140);
nor U39325 (N_39325,N_36172,N_36382);
or U39326 (N_39326,N_36672,N_36595);
xor U39327 (N_39327,N_36330,N_37198);
or U39328 (N_39328,N_37163,N_37451);
xnor U39329 (N_39329,N_37278,N_37251);
and U39330 (N_39330,N_37106,N_36327);
xor U39331 (N_39331,N_37718,N_37301);
nand U39332 (N_39332,N_36459,N_37668);
and U39333 (N_39333,N_37481,N_37360);
and U39334 (N_39334,N_37956,N_36392);
and U39335 (N_39335,N_36977,N_37988);
and U39336 (N_39336,N_36964,N_36512);
nand U39337 (N_39337,N_37357,N_36215);
nor U39338 (N_39338,N_36878,N_36747);
and U39339 (N_39339,N_37501,N_36001);
or U39340 (N_39340,N_37303,N_36133);
nor U39341 (N_39341,N_36774,N_36222);
xor U39342 (N_39342,N_37218,N_36231);
nand U39343 (N_39343,N_36206,N_36521);
and U39344 (N_39344,N_37641,N_36298);
nand U39345 (N_39345,N_37546,N_37661);
or U39346 (N_39346,N_36934,N_36704);
xnor U39347 (N_39347,N_37919,N_36278);
and U39348 (N_39348,N_37447,N_36112);
nor U39349 (N_39349,N_37502,N_37981);
or U39350 (N_39350,N_36668,N_37693);
or U39351 (N_39351,N_37436,N_36469);
nor U39352 (N_39352,N_37773,N_37634);
and U39353 (N_39353,N_37704,N_37111);
nand U39354 (N_39354,N_37727,N_37288);
nor U39355 (N_39355,N_37962,N_37919);
and U39356 (N_39356,N_36448,N_37343);
and U39357 (N_39357,N_36594,N_36286);
or U39358 (N_39358,N_37434,N_37043);
nor U39359 (N_39359,N_37496,N_37489);
nand U39360 (N_39360,N_37651,N_36226);
nand U39361 (N_39361,N_37336,N_36469);
nor U39362 (N_39362,N_37838,N_36209);
xor U39363 (N_39363,N_37728,N_36304);
xnor U39364 (N_39364,N_37900,N_36831);
or U39365 (N_39365,N_37962,N_36964);
nor U39366 (N_39366,N_37943,N_37627);
or U39367 (N_39367,N_36402,N_36752);
and U39368 (N_39368,N_37059,N_37193);
nor U39369 (N_39369,N_37537,N_36548);
nor U39370 (N_39370,N_37960,N_37519);
nor U39371 (N_39371,N_36891,N_37208);
and U39372 (N_39372,N_37128,N_37465);
or U39373 (N_39373,N_36326,N_36559);
xnor U39374 (N_39374,N_37732,N_36739);
nor U39375 (N_39375,N_36387,N_36381);
nand U39376 (N_39376,N_36619,N_37738);
and U39377 (N_39377,N_36571,N_36242);
nor U39378 (N_39378,N_37313,N_36894);
nor U39379 (N_39379,N_37418,N_37477);
nor U39380 (N_39380,N_36914,N_36051);
nor U39381 (N_39381,N_36881,N_37934);
or U39382 (N_39382,N_37922,N_37380);
and U39383 (N_39383,N_36593,N_37552);
and U39384 (N_39384,N_37813,N_37668);
and U39385 (N_39385,N_37999,N_36428);
xnor U39386 (N_39386,N_36506,N_36500);
nand U39387 (N_39387,N_36476,N_37939);
and U39388 (N_39388,N_36117,N_36514);
xnor U39389 (N_39389,N_36612,N_36725);
xor U39390 (N_39390,N_36373,N_36038);
nor U39391 (N_39391,N_37153,N_36330);
nand U39392 (N_39392,N_36507,N_36742);
nand U39393 (N_39393,N_36343,N_37909);
or U39394 (N_39394,N_36412,N_37253);
xnor U39395 (N_39395,N_37642,N_37573);
nor U39396 (N_39396,N_37118,N_37240);
or U39397 (N_39397,N_37897,N_37310);
or U39398 (N_39398,N_36652,N_36603);
or U39399 (N_39399,N_36891,N_37396);
xnor U39400 (N_39400,N_36555,N_37565);
xnor U39401 (N_39401,N_36770,N_36408);
nor U39402 (N_39402,N_37745,N_36697);
xor U39403 (N_39403,N_37114,N_36772);
and U39404 (N_39404,N_36256,N_36717);
nor U39405 (N_39405,N_36541,N_37119);
and U39406 (N_39406,N_36248,N_36568);
or U39407 (N_39407,N_37968,N_37206);
xor U39408 (N_39408,N_37080,N_36771);
nor U39409 (N_39409,N_37788,N_36279);
or U39410 (N_39410,N_37117,N_36432);
xor U39411 (N_39411,N_37819,N_36029);
or U39412 (N_39412,N_36699,N_37479);
xnor U39413 (N_39413,N_37062,N_37546);
xnor U39414 (N_39414,N_36056,N_36093);
nor U39415 (N_39415,N_36617,N_36379);
xor U39416 (N_39416,N_37262,N_37903);
nand U39417 (N_39417,N_37955,N_37800);
and U39418 (N_39418,N_37404,N_36626);
xor U39419 (N_39419,N_37457,N_37592);
or U39420 (N_39420,N_37372,N_37423);
nand U39421 (N_39421,N_36315,N_37675);
nand U39422 (N_39422,N_37548,N_37317);
nand U39423 (N_39423,N_36505,N_37555);
or U39424 (N_39424,N_37368,N_36577);
nand U39425 (N_39425,N_37162,N_36764);
nand U39426 (N_39426,N_36904,N_36590);
nand U39427 (N_39427,N_36261,N_37858);
nand U39428 (N_39428,N_36819,N_36206);
and U39429 (N_39429,N_37647,N_37169);
xnor U39430 (N_39430,N_36369,N_37223);
nor U39431 (N_39431,N_36144,N_36495);
nor U39432 (N_39432,N_36992,N_36295);
or U39433 (N_39433,N_37153,N_36463);
or U39434 (N_39434,N_37064,N_36142);
nor U39435 (N_39435,N_36590,N_37144);
and U39436 (N_39436,N_36879,N_36707);
nand U39437 (N_39437,N_36160,N_37061);
nor U39438 (N_39438,N_36580,N_36756);
and U39439 (N_39439,N_36348,N_37200);
nand U39440 (N_39440,N_37664,N_37728);
xor U39441 (N_39441,N_36625,N_37476);
xor U39442 (N_39442,N_37785,N_37673);
and U39443 (N_39443,N_36315,N_36172);
and U39444 (N_39444,N_37519,N_36666);
nor U39445 (N_39445,N_36454,N_36038);
and U39446 (N_39446,N_37016,N_37870);
or U39447 (N_39447,N_36559,N_37902);
and U39448 (N_39448,N_37771,N_37274);
and U39449 (N_39449,N_36954,N_36329);
xor U39450 (N_39450,N_36367,N_36914);
xor U39451 (N_39451,N_36211,N_37099);
nor U39452 (N_39452,N_36793,N_36513);
xor U39453 (N_39453,N_37468,N_36917);
or U39454 (N_39454,N_37599,N_37545);
nand U39455 (N_39455,N_36776,N_36116);
or U39456 (N_39456,N_37931,N_37367);
xor U39457 (N_39457,N_36361,N_36405);
xnor U39458 (N_39458,N_36188,N_36542);
nand U39459 (N_39459,N_36761,N_37886);
nand U39460 (N_39460,N_37891,N_37509);
or U39461 (N_39461,N_37543,N_37718);
nor U39462 (N_39462,N_36678,N_37482);
nor U39463 (N_39463,N_37121,N_37046);
xor U39464 (N_39464,N_36844,N_37875);
nand U39465 (N_39465,N_36304,N_36853);
and U39466 (N_39466,N_37214,N_37571);
xor U39467 (N_39467,N_37266,N_37923);
nor U39468 (N_39468,N_36268,N_36519);
xnor U39469 (N_39469,N_37960,N_36455);
xor U39470 (N_39470,N_37459,N_37779);
nand U39471 (N_39471,N_37221,N_36728);
or U39472 (N_39472,N_36930,N_37357);
xor U39473 (N_39473,N_36387,N_36904);
and U39474 (N_39474,N_37452,N_37865);
or U39475 (N_39475,N_37304,N_37593);
or U39476 (N_39476,N_36330,N_37259);
and U39477 (N_39477,N_36094,N_37091);
xor U39478 (N_39478,N_36033,N_36834);
and U39479 (N_39479,N_36592,N_37685);
nand U39480 (N_39480,N_37985,N_36732);
nor U39481 (N_39481,N_37732,N_37909);
nand U39482 (N_39482,N_36643,N_37857);
or U39483 (N_39483,N_36635,N_36259);
or U39484 (N_39484,N_37892,N_37404);
nor U39485 (N_39485,N_36944,N_37376);
nand U39486 (N_39486,N_37695,N_37170);
and U39487 (N_39487,N_36506,N_36683);
nor U39488 (N_39488,N_36130,N_37460);
and U39489 (N_39489,N_37254,N_37000);
nor U39490 (N_39490,N_37813,N_37353);
xnor U39491 (N_39491,N_36740,N_37003);
and U39492 (N_39492,N_37059,N_37827);
nand U39493 (N_39493,N_36705,N_36727);
xor U39494 (N_39494,N_37065,N_36383);
or U39495 (N_39495,N_37328,N_36611);
nor U39496 (N_39496,N_37496,N_37851);
and U39497 (N_39497,N_36643,N_37776);
nor U39498 (N_39498,N_37473,N_36920);
nor U39499 (N_39499,N_37266,N_37730);
nand U39500 (N_39500,N_37660,N_37753);
xnor U39501 (N_39501,N_37099,N_36698);
xnor U39502 (N_39502,N_36711,N_37767);
and U39503 (N_39503,N_36886,N_37466);
or U39504 (N_39504,N_37825,N_37728);
nor U39505 (N_39505,N_36338,N_36181);
xor U39506 (N_39506,N_37811,N_37605);
nor U39507 (N_39507,N_36257,N_36012);
xor U39508 (N_39508,N_37816,N_37755);
nand U39509 (N_39509,N_36292,N_36891);
or U39510 (N_39510,N_36250,N_36162);
nand U39511 (N_39511,N_36959,N_37532);
nor U39512 (N_39512,N_37333,N_36144);
nor U39513 (N_39513,N_36567,N_37972);
nor U39514 (N_39514,N_37026,N_36460);
xor U39515 (N_39515,N_36405,N_36110);
xnor U39516 (N_39516,N_36845,N_36112);
nor U39517 (N_39517,N_37266,N_36849);
xnor U39518 (N_39518,N_37858,N_36422);
or U39519 (N_39519,N_36900,N_37641);
and U39520 (N_39520,N_36887,N_36970);
xnor U39521 (N_39521,N_36098,N_37763);
nor U39522 (N_39522,N_36522,N_36305);
xnor U39523 (N_39523,N_36633,N_37402);
and U39524 (N_39524,N_36401,N_36083);
and U39525 (N_39525,N_37326,N_37800);
xor U39526 (N_39526,N_37242,N_37968);
nand U39527 (N_39527,N_37372,N_37577);
nand U39528 (N_39528,N_37659,N_37296);
nand U39529 (N_39529,N_36245,N_36069);
or U39530 (N_39530,N_36835,N_36644);
and U39531 (N_39531,N_37443,N_37746);
nor U39532 (N_39532,N_36208,N_36906);
xor U39533 (N_39533,N_37037,N_36316);
or U39534 (N_39534,N_36921,N_37882);
or U39535 (N_39535,N_37202,N_36807);
or U39536 (N_39536,N_36317,N_36361);
nor U39537 (N_39537,N_36443,N_36794);
nand U39538 (N_39538,N_36067,N_36295);
xor U39539 (N_39539,N_36644,N_36739);
nor U39540 (N_39540,N_37309,N_37392);
nand U39541 (N_39541,N_37356,N_36442);
and U39542 (N_39542,N_36770,N_37443);
or U39543 (N_39543,N_36077,N_36793);
or U39544 (N_39544,N_36092,N_36695);
xor U39545 (N_39545,N_37915,N_37849);
nand U39546 (N_39546,N_37085,N_36137);
xor U39547 (N_39547,N_36637,N_37789);
and U39548 (N_39548,N_37540,N_36684);
nand U39549 (N_39549,N_37865,N_36084);
nor U39550 (N_39550,N_37783,N_36317);
xnor U39551 (N_39551,N_37913,N_36238);
nand U39552 (N_39552,N_37748,N_37535);
and U39553 (N_39553,N_36162,N_36466);
or U39554 (N_39554,N_36763,N_36310);
xnor U39555 (N_39555,N_37812,N_37369);
xor U39556 (N_39556,N_37808,N_36034);
and U39557 (N_39557,N_37600,N_37372);
nand U39558 (N_39558,N_37772,N_37713);
nor U39559 (N_39559,N_37368,N_37504);
xnor U39560 (N_39560,N_37807,N_36136);
xnor U39561 (N_39561,N_37014,N_36389);
xor U39562 (N_39562,N_36618,N_37347);
and U39563 (N_39563,N_37057,N_36061);
nor U39564 (N_39564,N_36607,N_36797);
nor U39565 (N_39565,N_37892,N_37726);
nand U39566 (N_39566,N_37568,N_37011);
nand U39567 (N_39567,N_36777,N_37524);
nand U39568 (N_39568,N_36531,N_37579);
xnor U39569 (N_39569,N_36410,N_37341);
xnor U39570 (N_39570,N_36163,N_37814);
or U39571 (N_39571,N_37933,N_37508);
nand U39572 (N_39572,N_36809,N_36569);
or U39573 (N_39573,N_37751,N_37938);
and U39574 (N_39574,N_36834,N_37694);
xor U39575 (N_39575,N_36109,N_36092);
or U39576 (N_39576,N_36904,N_36458);
nand U39577 (N_39577,N_36466,N_36546);
xor U39578 (N_39578,N_36681,N_36323);
and U39579 (N_39579,N_36581,N_36105);
xor U39580 (N_39580,N_36389,N_37009);
nand U39581 (N_39581,N_36037,N_37330);
and U39582 (N_39582,N_36684,N_37823);
xor U39583 (N_39583,N_36046,N_37685);
xnor U39584 (N_39584,N_37747,N_37059);
xor U39585 (N_39585,N_36252,N_37288);
and U39586 (N_39586,N_37180,N_36001);
or U39587 (N_39587,N_36064,N_37767);
nor U39588 (N_39588,N_37654,N_37971);
or U39589 (N_39589,N_36582,N_37388);
nand U39590 (N_39590,N_36484,N_37122);
nor U39591 (N_39591,N_37712,N_37821);
xnor U39592 (N_39592,N_37618,N_36701);
xor U39593 (N_39593,N_37574,N_37431);
xnor U39594 (N_39594,N_36753,N_36151);
or U39595 (N_39595,N_37481,N_36901);
nand U39596 (N_39596,N_36807,N_36081);
or U39597 (N_39597,N_37049,N_36618);
or U39598 (N_39598,N_37824,N_37884);
xor U39599 (N_39599,N_37485,N_37649);
xnor U39600 (N_39600,N_36551,N_36088);
or U39601 (N_39601,N_36238,N_37764);
and U39602 (N_39602,N_37965,N_37086);
and U39603 (N_39603,N_36444,N_37393);
xnor U39604 (N_39604,N_37125,N_37154);
nand U39605 (N_39605,N_36223,N_36004);
and U39606 (N_39606,N_36588,N_36206);
or U39607 (N_39607,N_36322,N_36353);
nor U39608 (N_39608,N_37127,N_36557);
nand U39609 (N_39609,N_37848,N_37864);
nand U39610 (N_39610,N_36150,N_37146);
xor U39611 (N_39611,N_37548,N_37291);
nand U39612 (N_39612,N_37937,N_37311);
nor U39613 (N_39613,N_36315,N_37102);
xnor U39614 (N_39614,N_37145,N_37199);
or U39615 (N_39615,N_37174,N_37987);
or U39616 (N_39616,N_37901,N_36047);
and U39617 (N_39617,N_36554,N_36694);
nand U39618 (N_39618,N_36125,N_37612);
xnor U39619 (N_39619,N_37884,N_37210);
nor U39620 (N_39620,N_37299,N_36202);
and U39621 (N_39621,N_36759,N_36686);
and U39622 (N_39622,N_36197,N_37536);
nand U39623 (N_39623,N_36350,N_36211);
nor U39624 (N_39624,N_36379,N_36434);
and U39625 (N_39625,N_37845,N_36682);
nand U39626 (N_39626,N_37823,N_36203);
nand U39627 (N_39627,N_37329,N_36269);
or U39628 (N_39628,N_36972,N_37726);
xor U39629 (N_39629,N_36285,N_36557);
and U39630 (N_39630,N_36725,N_37242);
xor U39631 (N_39631,N_37600,N_37611);
and U39632 (N_39632,N_37909,N_37166);
nor U39633 (N_39633,N_36925,N_36804);
and U39634 (N_39634,N_36573,N_36183);
xor U39635 (N_39635,N_37722,N_37944);
nor U39636 (N_39636,N_36860,N_36836);
nand U39637 (N_39637,N_37042,N_36197);
xnor U39638 (N_39638,N_37932,N_36207);
and U39639 (N_39639,N_36307,N_36270);
nand U39640 (N_39640,N_37728,N_36105);
nand U39641 (N_39641,N_36333,N_36348);
nor U39642 (N_39642,N_36558,N_37349);
and U39643 (N_39643,N_36291,N_37686);
nand U39644 (N_39644,N_36970,N_37209);
or U39645 (N_39645,N_36214,N_36361);
and U39646 (N_39646,N_37344,N_36188);
xor U39647 (N_39647,N_37070,N_37282);
and U39648 (N_39648,N_36233,N_37113);
nand U39649 (N_39649,N_37828,N_37216);
and U39650 (N_39650,N_37037,N_37013);
and U39651 (N_39651,N_36739,N_36303);
and U39652 (N_39652,N_37066,N_36738);
or U39653 (N_39653,N_37260,N_37390);
xnor U39654 (N_39654,N_37405,N_36094);
xnor U39655 (N_39655,N_37649,N_36194);
xnor U39656 (N_39656,N_36766,N_36353);
xnor U39657 (N_39657,N_37371,N_37244);
nor U39658 (N_39658,N_36351,N_37005);
xnor U39659 (N_39659,N_37220,N_37863);
xor U39660 (N_39660,N_37914,N_37993);
and U39661 (N_39661,N_36044,N_37777);
or U39662 (N_39662,N_36581,N_37688);
and U39663 (N_39663,N_37067,N_37004);
nand U39664 (N_39664,N_37843,N_36099);
and U39665 (N_39665,N_37337,N_37580);
nor U39666 (N_39666,N_37652,N_37756);
nor U39667 (N_39667,N_36763,N_36301);
xnor U39668 (N_39668,N_36517,N_36081);
or U39669 (N_39669,N_37176,N_36747);
nor U39670 (N_39670,N_37558,N_37901);
and U39671 (N_39671,N_36907,N_36078);
and U39672 (N_39672,N_37119,N_36757);
and U39673 (N_39673,N_36309,N_36294);
and U39674 (N_39674,N_37992,N_37748);
or U39675 (N_39675,N_37267,N_37886);
xor U39676 (N_39676,N_37369,N_36436);
and U39677 (N_39677,N_36490,N_37221);
nand U39678 (N_39678,N_37156,N_36471);
nand U39679 (N_39679,N_37286,N_36154);
and U39680 (N_39680,N_36575,N_37799);
nand U39681 (N_39681,N_37377,N_37953);
xnor U39682 (N_39682,N_36179,N_36929);
nor U39683 (N_39683,N_37500,N_36744);
nand U39684 (N_39684,N_37404,N_37549);
nor U39685 (N_39685,N_37065,N_36597);
or U39686 (N_39686,N_36181,N_37272);
xor U39687 (N_39687,N_36830,N_37717);
and U39688 (N_39688,N_37893,N_37101);
or U39689 (N_39689,N_36614,N_36448);
xnor U39690 (N_39690,N_37912,N_36922);
xnor U39691 (N_39691,N_37941,N_37913);
or U39692 (N_39692,N_36076,N_36551);
nor U39693 (N_39693,N_36972,N_36132);
nor U39694 (N_39694,N_36135,N_36795);
xnor U39695 (N_39695,N_37736,N_37823);
or U39696 (N_39696,N_37650,N_36997);
and U39697 (N_39697,N_36372,N_37485);
and U39698 (N_39698,N_37050,N_36037);
or U39699 (N_39699,N_36927,N_37647);
nor U39700 (N_39700,N_37434,N_37517);
nor U39701 (N_39701,N_36262,N_37990);
or U39702 (N_39702,N_36573,N_36272);
nor U39703 (N_39703,N_37628,N_36924);
nand U39704 (N_39704,N_37648,N_36809);
nand U39705 (N_39705,N_37798,N_36443);
nand U39706 (N_39706,N_36919,N_37177);
xor U39707 (N_39707,N_37848,N_36310);
nor U39708 (N_39708,N_36634,N_36905);
nand U39709 (N_39709,N_36581,N_37517);
or U39710 (N_39710,N_37589,N_36054);
and U39711 (N_39711,N_36358,N_37078);
nand U39712 (N_39712,N_37709,N_37637);
and U39713 (N_39713,N_37104,N_37647);
nand U39714 (N_39714,N_36071,N_37612);
xnor U39715 (N_39715,N_36689,N_37813);
xnor U39716 (N_39716,N_36842,N_36616);
nand U39717 (N_39717,N_36921,N_37378);
xor U39718 (N_39718,N_37745,N_36161);
nor U39719 (N_39719,N_37483,N_36375);
xor U39720 (N_39720,N_36767,N_36233);
or U39721 (N_39721,N_37722,N_36995);
or U39722 (N_39722,N_36629,N_37239);
xnor U39723 (N_39723,N_36612,N_37334);
nor U39724 (N_39724,N_37862,N_37589);
or U39725 (N_39725,N_37946,N_36789);
or U39726 (N_39726,N_37359,N_36369);
xor U39727 (N_39727,N_36936,N_36960);
or U39728 (N_39728,N_37651,N_36458);
nor U39729 (N_39729,N_37073,N_37897);
or U39730 (N_39730,N_37657,N_37941);
nand U39731 (N_39731,N_36780,N_37158);
or U39732 (N_39732,N_37951,N_36956);
xnor U39733 (N_39733,N_37112,N_36373);
nand U39734 (N_39734,N_36717,N_37211);
or U39735 (N_39735,N_36658,N_36145);
xnor U39736 (N_39736,N_36890,N_37780);
or U39737 (N_39737,N_37089,N_36300);
or U39738 (N_39738,N_37581,N_37535);
nand U39739 (N_39739,N_36406,N_37352);
and U39740 (N_39740,N_36982,N_37075);
xnor U39741 (N_39741,N_36415,N_37207);
nand U39742 (N_39742,N_36726,N_37090);
or U39743 (N_39743,N_36135,N_36908);
and U39744 (N_39744,N_36913,N_36765);
and U39745 (N_39745,N_37156,N_36278);
nor U39746 (N_39746,N_37892,N_36900);
nor U39747 (N_39747,N_36545,N_36950);
or U39748 (N_39748,N_36721,N_36799);
and U39749 (N_39749,N_37528,N_36448);
nor U39750 (N_39750,N_37726,N_37180);
xnor U39751 (N_39751,N_37716,N_37772);
nor U39752 (N_39752,N_36124,N_36369);
nand U39753 (N_39753,N_36715,N_36265);
xor U39754 (N_39754,N_36943,N_37096);
nor U39755 (N_39755,N_37537,N_36448);
nand U39756 (N_39756,N_37130,N_37630);
nor U39757 (N_39757,N_37415,N_36340);
or U39758 (N_39758,N_37702,N_37772);
and U39759 (N_39759,N_37558,N_36009);
nand U39760 (N_39760,N_36804,N_37905);
nor U39761 (N_39761,N_36086,N_36346);
nand U39762 (N_39762,N_36389,N_37646);
nand U39763 (N_39763,N_37347,N_37450);
and U39764 (N_39764,N_37647,N_37417);
nor U39765 (N_39765,N_36857,N_36294);
and U39766 (N_39766,N_36385,N_36065);
or U39767 (N_39767,N_36742,N_36562);
xor U39768 (N_39768,N_37124,N_37545);
nor U39769 (N_39769,N_37491,N_36544);
and U39770 (N_39770,N_36087,N_36143);
or U39771 (N_39771,N_36687,N_36878);
nor U39772 (N_39772,N_36443,N_36357);
and U39773 (N_39773,N_36206,N_36478);
nor U39774 (N_39774,N_37575,N_37787);
nor U39775 (N_39775,N_36299,N_36256);
nand U39776 (N_39776,N_36497,N_36872);
nor U39777 (N_39777,N_37001,N_37918);
xnor U39778 (N_39778,N_37048,N_37515);
nand U39779 (N_39779,N_36591,N_37886);
or U39780 (N_39780,N_37758,N_37501);
nand U39781 (N_39781,N_37800,N_37143);
and U39782 (N_39782,N_36887,N_36118);
or U39783 (N_39783,N_37229,N_37661);
nand U39784 (N_39784,N_37932,N_36363);
or U39785 (N_39785,N_36479,N_36183);
nand U39786 (N_39786,N_37510,N_37407);
and U39787 (N_39787,N_37840,N_37107);
and U39788 (N_39788,N_36992,N_37434);
xnor U39789 (N_39789,N_36197,N_36579);
nand U39790 (N_39790,N_36582,N_36527);
nand U39791 (N_39791,N_36391,N_36701);
nand U39792 (N_39792,N_36281,N_37461);
xnor U39793 (N_39793,N_36365,N_36341);
or U39794 (N_39794,N_36296,N_37833);
or U39795 (N_39795,N_36063,N_36955);
nor U39796 (N_39796,N_37369,N_37989);
nor U39797 (N_39797,N_36119,N_36005);
xnor U39798 (N_39798,N_36600,N_36222);
nor U39799 (N_39799,N_37840,N_37019);
nor U39800 (N_39800,N_37318,N_37456);
and U39801 (N_39801,N_37152,N_37347);
xnor U39802 (N_39802,N_36673,N_36765);
or U39803 (N_39803,N_37894,N_37452);
xnor U39804 (N_39804,N_36118,N_37554);
nor U39805 (N_39805,N_36992,N_36086);
xnor U39806 (N_39806,N_37281,N_36382);
xor U39807 (N_39807,N_36009,N_36011);
and U39808 (N_39808,N_37601,N_36023);
nor U39809 (N_39809,N_36652,N_37873);
xor U39810 (N_39810,N_36653,N_36025);
or U39811 (N_39811,N_37297,N_37985);
or U39812 (N_39812,N_37080,N_36042);
and U39813 (N_39813,N_37172,N_37317);
xnor U39814 (N_39814,N_37940,N_36237);
nor U39815 (N_39815,N_37714,N_37740);
xnor U39816 (N_39816,N_36681,N_37714);
xnor U39817 (N_39817,N_36904,N_36607);
nand U39818 (N_39818,N_37854,N_37694);
nor U39819 (N_39819,N_37378,N_37429);
xnor U39820 (N_39820,N_36147,N_37704);
nor U39821 (N_39821,N_37431,N_37003);
xnor U39822 (N_39822,N_36025,N_36508);
nand U39823 (N_39823,N_37614,N_37126);
or U39824 (N_39824,N_37279,N_36311);
nor U39825 (N_39825,N_37757,N_37244);
and U39826 (N_39826,N_36885,N_36013);
xor U39827 (N_39827,N_37548,N_37478);
and U39828 (N_39828,N_37366,N_37745);
or U39829 (N_39829,N_37041,N_36628);
or U39830 (N_39830,N_37663,N_37502);
or U39831 (N_39831,N_37447,N_37376);
and U39832 (N_39832,N_36451,N_37236);
nand U39833 (N_39833,N_36335,N_37347);
nand U39834 (N_39834,N_36244,N_36695);
nor U39835 (N_39835,N_37727,N_37503);
and U39836 (N_39836,N_36999,N_36744);
or U39837 (N_39837,N_36105,N_36766);
or U39838 (N_39838,N_37703,N_37439);
nor U39839 (N_39839,N_37016,N_36318);
and U39840 (N_39840,N_37713,N_37286);
xnor U39841 (N_39841,N_36094,N_36861);
nor U39842 (N_39842,N_37434,N_37307);
nand U39843 (N_39843,N_37026,N_36428);
or U39844 (N_39844,N_37135,N_37665);
nor U39845 (N_39845,N_36184,N_37072);
and U39846 (N_39846,N_37924,N_37465);
nand U39847 (N_39847,N_37336,N_37202);
xor U39848 (N_39848,N_37403,N_37767);
and U39849 (N_39849,N_37000,N_37790);
or U39850 (N_39850,N_37571,N_36001);
xor U39851 (N_39851,N_36213,N_37881);
nor U39852 (N_39852,N_37301,N_36389);
or U39853 (N_39853,N_36243,N_37067);
and U39854 (N_39854,N_36943,N_37454);
xor U39855 (N_39855,N_37181,N_36123);
xnor U39856 (N_39856,N_36507,N_36103);
and U39857 (N_39857,N_36733,N_36555);
nor U39858 (N_39858,N_36724,N_36834);
nand U39859 (N_39859,N_37181,N_36488);
nor U39860 (N_39860,N_37125,N_36686);
nand U39861 (N_39861,N_36971,N_37127);
nand U39862 (N_39862,N_36930,N_36158);
xor U39863 (N_39863,N_37307,N_36735);
nand U39864 (N_39864,N_37941,N_37915);
xnor U39865 (N_39865,N_36644,N_37981);
nand U39866 (N_39866,N_36184,N_36028);
nand U39867 (N_39867,N_37979,N_36080);
or U39868 (N_39868,N_37304,N_36313);
nor U39869 (N_39869,N_37621,N_37288);
nor U39870 (N_39870,N_36211,N_36638);
nor U39871 (N_39871,N_37542,N_36043);
nor U39872 (N_39872,N_37520,N_37547);
and U39873 (N_39873,N_36981,N_36998);
or U39874 (N_39874,N_36959,N_37050);
nor U39875 (N_39875,N_36503,N_37269);
nor U39876 (N_39876,N_36666,N_37227);
nand U39877 (N_39877,N_36830,N_36358);
xor U39878 (N_39878,N_37715,N_37435);
xor U39879 (N_39879,N_36822,N_36720);
or U39880 (N_39880,N_36605,N_37323);
nor U39881 (N_39881,N_36007,N_36821);
nor U39882 (N_39882,N_37311,N_37290);
nand U39883 (N_39883,N_37276,N_37113);
xor U39884 (N_39884,N_37208,N_37517);
nor U39885 (N_39885,N_37892,N_36293);
xor U39886 (N_39886,N_36828,N_36364);
xor U39887 (N_39887,N_36809,N_37483);
nor U39888 (N_39888,N_37010,N_37434);
and U39889 (N_39889,N_36644,N_37798);
or U39890 (N_39890,N_36411,N_36136);
xnor U39891 (N_39891,N_37750,N_37758);
xor U39892 (N_39892,N_36455,N_36593);
and U39893 (N_39893,N_36395,N_36176);
or U39894 (N_39894,N_37787,N_37824);
and U39895 (N_39895,N_36399,N_37405);
and U39896 (N_39896,N_36819,N_37286);
nor U39897 (N_39897,N_36252,N_36214);
nand U39898 (N_39898,N_37162,N_37056);
and U39899 (N_39899,N_36959,N_36771);
or U39900 (N_39900,N_37459,N_37486);
xor U39901 (N_39901,N_36315,N_37103);
or U39902 (N_39902,N_37220,N_36889);
and U39903 (N_39903,N_37306,N_37601);
and U39904 (N_39904,N_37374,N_36508);
or U39905 (N_39905,N_37916,N_37392);
or U39906 (N_39906,N_37086,N_36136);
xor U39907 (N_39907,N_36302,N_36096);
and U39908 (N_39908,N_36347,N_37348);
nand U39909 (N_39909,N_36589,N_37761);
or U39910 (N_39910,N_36745,N_37872);
xnor U39911 (N_39911,N_37105,N_37611);
nand U39912 (N_39912,N_36810,N_37345);
nor U39913 (N_39913,N_37382,N_36662);
xor U39914 (N_39914,N_37516,N_36567);
nor U39915 (N_39915,N_36078,N_36069);
and U39916 (N_39916,N_37765,N_37926);
and U39917 (N_39917,N_37920,N_36550);
or U39918 (N_39918,N_36481,N_36492);
nand U39919 (N_39919,N_36036,N_37975);
or U39920 (N_39920,N_37727,N_37980);
or U39921 (N_39921,N_37738,N_36907);
xor U39922 (N_39922,N_37790,N_37432);
nand U39923 (N_39923,N_37932,N_36107);
xnor U39924 (N_39924,N_36308,N_37425);
nand U39925 (N_39925,N_37329,N_36420);
nand U39926 (N_39926,N_37833,N_36970);
or U39927 (N_39927,N_36341,N_36718);
or U39928 (N_39928,N_37913,N_36437);
or U39929 (N_39929,N_37172,N_36428);
nand U39930 (N_39930,N_37085,N_37318);
nand U39931 (N_39931,N_36402,N_36539);
nand U39932 (N_39932,N_37000,N_36300);
or U39933 (N_39933,N_37334,N_36165);
nand U39934 (N_39934,N_36794,N_36665);
or U39935 (N_39935,N_36245,N_37497);
nand U39936 (N_39936,N_36655,N_36277);
and U39937 (N_39937,N_36512,N_36788);
nand U39938 (N_39938,N_37735,N_37034);
and U39939 (N_39939,N_37887,N_37524);
or U39940 (N_39940,N_37727,N_36336);
or U39941 (N_39941,N_36121,N_36076);
nor U39942 (N_39942,N_36597,N_36295);
and U39943 (N_39943,N_37455,N_36471);
and U39944 (N_39944,N_37916,N_37566);
nand U39945 (N_39945,N_36510,N_36020);
nor U39946 (N_39946,N_37314,N_37440);
xor U39947 (N_39947,N_36821,N_37168);
xor U39948 (N_39948,N_36467,N_37544);
and U39949 (N_39949,N_37790,N_36751);
nor U39950 (N_39950,N_36677,N_36332);
and U39951 (N_39951,N_37355,N_37594);
nor U39952 (N_39952,N_36218,N_36306);
and U39953 (N_39953,N_36087,N_37697);
nor U39954 (N_39954,N_36089,N_36249);
or U39955 (N_39955,N_37095,N_37306);
or U39956 (N_39956,N_36354,N_37788);
xor U39957 (N_39957,N_36275,N_36058);
and U39958 (N_39958,N_36388,N_36238);
and U39959 (N_39959,N_37693,N_37536);
or U39960 (N_39960,N_37870,N_37678);
nand U39961 (N_39961,N_36613,N_36667);
or U39962 (N_39962,N_36670,N_37554);
or U39963 (N_39963,N_36878,N_37834);
nor U39964 (N_39964,N_37323,N_37600);
and U39965 (N_39965,N_36240,N_36491);
nand U39966 (N_39966,N_36881,N_36797);
nand U39967 (N_39967,N_37673,N_36811);
xor U39968 (N_39968,N_37170,N_37117);
or U39969 (N_39969,N_37272,N_37168);
or U39970 (N_39970,N_37987,N_36286);
nor U39971 (N_39971,N_36490,N_36887);
xnor U39972 (N_39972,N_36240,N_37833);
nor U39973 (N_39973,N_37966,N_37323);
or U39974 (N_39974,N_36052,N_37528);
xor U39975 (N_39975,N_37702,N_36328);
xnor U39976 (N_39976,N_36215,N_36193);
nand U39977 (N_39977,N_37201,N_36461);
nand U39978 (N_39978,N_37390,N_37228);
xor U39979 (N_39979,N_36751,N_36738);
nand U39980 (N_39980,N_36693,N_37378);
nand U39981 (N_39981,N_37346,N_36462);
and U39982 (N_39982,N_36752,N_37326);
xnor U39983 (N_39983,N_37073,N_36670);
xnor U39984 (N_39984,N_37581,N_36119);
nor U39985 (N_39985,N_37857,N_37739);
nand U39986 (N_39986,N_37429,N_37491);
nand U39987 (N_39987,N_37279,N_36982);
nand U39988 (N_39988,N_37774,N_37979);
xnor U39989 (N_39989,N_36900,N_37175);
nand U39990 (N_39990,N_36728,N_36481);
or U39991 (N_39991,N_37986,N_36647);
nor U39992 (N_39992,N_36576,N_37473);
xnor U39993 (N_39993,N_36380,N_37036);
xor U39994 (N_39994,N_36855,N_37182);
and U39995 (N_39995,N_37717,N_37241);
nor U39996 (N_39996,N_36280,N_37983);
or U39997 (N_39997,N_37788,N_37722);
nand U39998 (N_39998,N_36367,N_36706);
nor U39999 (N_39999,N_37650,N_37841);
nand U40000 (N_40000,N_38055,N_38062);
nor U40001 (N_40001,N_38398,N_38788);
and U40002 (N_40002,N_38854,N_39090);
and U40003 (N_40003,N_38798,N_38686);
nand U40004 (N_40004,N_38615,N_39048);
and U40005 (N_40005,N_39647,N_39585);
or U40006 (N_40006,N_39083,N_39021);
xnor U40007 (N_40007,N_38784,N_38372);
xor U40008 (N_40008,N_39349,N_38144);
nand U40009 (N_40009,N_39161,N_39502);
xor U40010 (N_40010,N_39543,N_39322);
nand U40011 (N_40011,N_39866,N_39217);
and U40012 (N_40012,N_39186,N_38648);
xnor U40013 (N_40013,N_39886,N_39984);
nor U40014 (N_40014,N_38452,N_39261);
nor U40015 (N_40015,N_39494,N_39417);
xnor U40016 (N_40016,N_38729,N_39882);
xnor U40017 (N_40017,N_39373,N_39997);
nor U40018 (N_40018,N_39939,N_38429);
nand U40019 (N_40019,N_38698,N_38426);
and U40020 (N_40020,N_38265,N_39781);
or U40021 (N_40021,N_39482,N_39857);
nor U40022 (N_40022,N_39497,N_38043);
or U40023 (N_40023,N_39218,N_38186);
and U40024 (N_40024,N_38827,N_39243);
and U40025 (N_40025,N_39589,N_38324);
and U40026 (N_40026,N_39446,N_38194);
and U40027 (N_40027,N_38039,N_38303);
nand U40028 (N_40028,N_39131,N_39343);
or U40029 (N_40029,N_39526,N_39138);
or U40030 (N_40030,N_39480,N_39535);
nor U40031 (N_40031,N_39075,N_38430);
nor U40032 (N_40032,N_39118,N_38734);
nor U40033 (N_40033,N_39979,N_39838);
xor U40034 (N_40034,N_39178,N_38713);
or U40035 (N_40035,N_38354,N_39995);
xnor U40036 (N_40036,N_39077,N_39358);
nor U40037 (N_40037,N_39677,N_39806);
xor U40038 (N_40038,N_38147,N_38860);
nor U40039 (N_40039,N_38486,N_39227);
xnor U40040 (N_40040,N_38374,N_39208);
nand U40041 (N_40041,N_39050,N_39938);
nor U40042 (N_40042,N_38720,N_38752);
or U40043 (N_40043,N_39923,N_38738);
nand U40044 (N_40044,N_38740,N_39928);
xnor U40045 (N_40045,N_38812,N_39903);
and U40046 (N_40046,N_39709,N_38819);
xor U40047 (N_40047,N_39418,N_39689);
nor U40048 (N_40048,N_38905,N_39952);
xnor U40049 (N_40049,N_38549,N_39286);
nand U40050 (N_40050,N_39609,N_38356);
xnor U40051 (N_40051,N_39421,N_39123);
and U40052 (N_40052,N_38278,N_39154);
or U40053 (N_40053,N_38657,N_38973);
and U40054 (N_40054,N_39725,N_38660);
and U40055 (N_40055,N_39405,N_39086);
xor U40056 (N_40056,N_39622,N_39630);
nand U40057 (N_40057,N_38034,N_39910);
and U40058 (N_40058,N_38557,N_38795);
nor U40059 (N_40059,N_38191,N_39026);
nor U40060 (N_40060,N_38273,N_38439);
xor U40061 (N_40061,N_38754,N_39691);
or U40062 (N_40062,N_39255,N_38029);
and U40063 (N_40063,N_39345,N_38662);
or U40064 (N_40064,N_38443,N_38682);
xnor U40065 (N_40065,N_39614,N_38182);
or U40066 (N_40066,N_39173,N_38096);
nand U40067 (N_40067,N_39750,N_39909);
xnor U40068 (N_40068,N_39003,N_38117);
xnor U40069 (N_40069,N_38652,N_39862);
and U40070 (N_40070,N_38427,N_39445);
nor U40071 (N_40071,N_38759,N_38536);
nand U40072 (N_40072,N_39382,N_39391);
or U40073 (N_40073,N_38506,N_38098);
or U40074 (N_40074,N_38309,N_38166);
or U40075 (N_40075,N_38688,N_39238);
or U40076 (N_40076,N_38793,N_38073);
or U40077 (N_40077,N_39976,N_39377);
xnor U40078 (N_40078,N_39333,N_38215);
or U40079 (N_40079,N_38010,N_39430);
xor U40080 (N_40080,N_39011,N_38663);
or U40081 (N_40081,N_39561,N_38004);
or U40082 (N_40082,N_38808,N_38512);
and U40083 (N_40083,N_38944,N_38751);
or U40084 (N_40084,N_39608,N_38640);
and U40085 (N_40085,N_38375,N_39245);
or U40086 (N_40086,N_39853,N_39848);
and U40087 (N_40087,N_38026,N_38507);
and U40088 (N_40088,N_39594,N_39168);
xor U40089 (N_40089,N_38395,N_38529);
or U40090 (N_40090,N_39125,N_38225);
nand U40091 (N_40091,N_38570,N_39996);
xnor U40092 (N_40092,N_38041,N_39571);
xor U40093 (N_40093,N_38597,N_39287);
or U40094 (N_40094,N_39890,N_39635);
or U40095 (N_40095,N_38792,N_38164);
xor U40096 (N_40096,N_39302,N_39401);
xnor U40097 (N_40097,N_39751,N_38092);
or U40098 (N_40098,N_38327,N_38765);
nand U40099 (N_40099,N_38176,N_38878);
or U40100 (N_40100,N_38775,N_38442);
xor U40101 (N_40101,N_39189,N_39694);
xor U40102 (N_40102,N_38080,N_39303);
nand U40103 (N_40103,N_39711,N_38932);
xnor U40104 (N_40104,N_39926,N_39463);
xnor U40105 (N_40105,N_38755,N_39214);
nand U40106 (N_40106,N_38379,N_39182);
nand U40107 (N_40107,N_38789,N_38076);
and U40108 (N_40108,N_39896,N_38619);
and U40109 (N_40109,N_38220,N_39251);
xor U40110 (N_40110,N_38779,N_38000);
or U40111 (N_40111,N_38226,N_38006);
nor U40112 (N_40112,N_39328,N_39868);
nor U40113 (N_40113,N_38193,N_39241);
nor U40114 (N_40114,N_38678,N_39768);
nor U40115 (N_40115,N_39789,N_38484);
and U40116 (N_40116,N_38264,N_38032);
and U40117 (N_40117,N_39422,N_39198);
nand U40118 (N_40118,N_38742,N_39252);
xor U40119 (N_40119,N_39546,N_39234);
nor U40120 (N_40120,N_39568,N_39216);
xnor U40121 (N_40121,N_39793,N_39701);
xnor U40122 (N_40122,N_38773,N_38883);
xor U40123 (N_40123,N_38391,N_39784);
nand U40124 (N_40124,N_38940,N_38873);
nor U40125 (N_40125,N_38587,N_38192);
nor U40126 (N_40126,N_38360,N_38780);
or U40127 (N_40127,N_39437,N_39796);
nor U40128 (N_40128,N_39628,N_38224);
and U40129 (N_40129,N_38051,N_39072);
nor U40130 (N_40130,N_39335,N_39912);
and U40131 (N_40131,N_38605,N_39905);
or U40132 (N_40132,N_38556,N_38376);
or U40133 (N_40133,N_38377,N_39069);
or U40134 (N_40134,N_38511,N_39961);
and U40135 (N_40135,N_39672,N_38976);
xor U40136 (N_40136,N_39079,N_38340);
nor U40137 (N_40137,N_38135,N_38210);
xnor U40138 (N_40138,N_39670,N_38977);
nor U40139 (N_40139,N_39371,N_38960);
xor U40140 (N_40140,N_39901,N_38544);
or U40141 (N_40141,N_39106,N_38269);
nor U40142 (N_40142,N_39393,N_39586);
nand U40143 (N_40143,N_38563,N_39511);
and U40144 (N_40144,N_39441,N_39885);
nor U40145 (N_40145,N_38542,N_39311);
nand U40146 (N_40146,N_39347,N_38679);
xor U40147 (N_40147,N_39936,N_39974);
xor U40148 (N_40148,N_39877,N_39193);
nor U40149 (N_40149,N_39855,N_38343);
xnor U40150 (N_40150,N_39743,N_39498);
xnor U40151 (N_40151,N_38986,N_38124);
nand U40152 (N_40152,N_38867,N_38611);
xnor U40153 (N_40153,N_39529,N_38888);
or U40154 (N_40154,N_38332,N_39596);
xnor U40155 (N_40155,N_38084,N_39712);
xor U40156 (N_40156,N_38150,N_38001);
or U40157 (N_40157,N_39752,N_38071);
xor U40158 (N_40158,N_38562,N_39331);
nor U40159 (N_40159,N_39068,N_39368);
or U40160 (N_40160,N_39676,N_39863);
and U40161 (N_40161,N_38585,N_39757);
or U40162 (N_40162,N_38958,N_39969);
or U40163 (N_40163,N_39142,N_38548);
xor U40164 (N_40164,N_39872,N_39816);
nor U40165 (N_40165,N_38524,N_39459);
or U40166 (N_40166,N_39272,N_38475);
and U40167 (N_40167,N_38467,N_39305);
xor U40168 (N_40168,N_39550,N_39388);
xor U40169 (N_40169,N_39284,N_38820);
or U40170 (N_40170,N_38290,N_39247);
nand U40171 (N_40171,N_39668,N_38276);
xor U40172 (N_40172,N_39966,N_39661);
nor U40173 (N_40173,N_38982,N_38105);
nand U40174 (N_40174,N_39637,N_38380);
xor U40175 (N_40175,N_38338,N_38440);
or U40176 (N_40176,N_39508,N_39600);
nand U40177 (N_40177,N_39492,N_39491);
xnor U40178 (N_40178,N_39562,N_38271);
nor U40179 (N_40179,N_38540,N_38127);
or U40180 (N_40180,N_39879,N_38400);
nand U40181 (N_40181,N_38983,N_39950);
and U40182 (N_40182,N_38647,N_39899);
nor U40183 (N_40183,N_38911,N_39120);
and U40184 (N_40184,N_39232,N_38152);
xnor U40185 (N_40185,N_39636,N_38764);
xnor U40186 (N_40186,N_38632,N_39144);
or U40187 (N_40187,N_39854,N_38670);
nor U40188 (N_40188,N_39051,N_38618);
xnor U40189 (N_40189,N_38950,N_39192);
nor U40190 (N_40190,N_38884,N_39755);
xor U40191 (N_40191,N_39802,N_38805);
nand U40192 (N_40192,N_38591,N_39046);
and U40193 (N_40193,N_39031,N_39867);
nor U40194 (N_40194,N_39704,N_38684);
xnor U40195 (N_40195,N_38658,N_38261);
nor U40196 (N_40196,N_39549,N_38716);
and U40197 (N_40197,N_38997,N_39840);
nand U40198 (N_40198,N_38833,N_39460);
nor U40199 (N_40199,N_39185,N_38140);
xnor U40200 (N_40200,N_38125,N_38546);
or U40201 (N_40201,N_38769,N_39429);
xor U40202 (N_40202,N_39572,N_38661);
xnor U40203 (N_40203,N_39257,N_38211);
xnor U40204 (N_40204,N_38862,N_39276);
nor U40205 (N_40205,N_39524,N_39728);
nand U40206 (N_40206,N_39036,N_38250);
and U40207 (N_40207,N_39773,N_39239);
nand U40208 (N_40208,N_39532,N_38412);
xor U40209 (N_40209,N_39457,N_39865);
xor U40210 (N_40210,N_39058,N_38757);
or U40211 (N_40211,N_38199,N_39558);
and U40212 (N_40212,N_38596,N_39327);
nand U40213 (N_40213,N_39620,N_39501);
nand U40214 (N_40214,N_38943,N_39645);
and U40215 (N_40215,N_39012,N_38623);
nor U40216 (N_40216,N_39891,N_39392);
xor U40217 (N_40217,N_38057,N_39930);
nor U40218 (N_40218,N_39692,N_38020);
or U40219 (N_40219,N_39530,N_39248);
or U40220 (N_40220,N_38525,N_38846);
and U40221 (N_40221,N_38279,N_38257);
or U40222 (N_40222,N_39250,N_39597);
xor U40223 (N_40223,N_38009,N_38107);
xor U40224 (N_40224,N_38803,N_38709);
and U40225 (N_40225,N_38247,N_39619);
nand U40226 (N_40226,N_39512,N_39657);
xor U40227 (N_40227,N_39367,N_38415);
or U40228 (N_40228,N_38835,N_38069);
nor U40229 (N_40229,N_38244,N_39481);
and U40230 (N_40230,N_39499,N_39813);
xnor U40231 (N_40231,N_38879,N_39658);
nand U40232 (N_40232,N_39778,N_39700);
xnor U40233 (N_40233,N_38558,N_39389);
nand U40234 (N_40234,N_39766,N_39883);
nor U40235 (N_40235,N_38896,N_38025);
or U40236 (N_40236,N_38059,N_39528);
xor U40237 (N_40237,N_39861,N_39605);
xor U40238 (N_40238,N_38504,N_39588);
nor U40239 (N_40239,N_39834,N_38749);
xor U40240 (N_40240,N_39108,N_39917);
and U40241 (N_40241,N_39277,N_38876);
nand U40242 (N_40242,N_39111,N_38527);
or U40243 (N_40243,N_38482,N_39856);
nand U40244 (N_40244,N_39795,N_39733);
xor U40245 (N_40245,N_38785,N_39330);
or U40246 (N_40246,N_38696,N_39159);
or U40247 (N_40247,N_38077,N_39196);
xnor U40248 (N_40248,N_38385,N_38207);
nor U40249 (N_40249,N_38807,N_38665);
and U40250 (N_40250,N_38566,N_38310);
xnor U40251 (N_40251,N_38460,N_39082);
nand U40252 (N_40252,N_39522,N_38510);
and U40253 (N_40253,N_39506,N_39209);
nor U40254 (N_40254,N_39279,N_38913);
nand U40255 (N_40255,N_38607,N_38367);
nor U40256 (N_40256,N_39607,N_38937);
and U40257 (N_40257,N_39307,N_39019);
and U40258 (N_40258,N_39285,N_39032);
xor U40259 (N_40259,N_39925,N_38704);
nand U40260 (N_40260,N_39317,N_39361);
nand U40261 (N_40261,N_38768,N_38142);
xor U40262 (N_40262,N_39881,N_39246);
and U40263 (N_40263,N_38438,N_38169);
or U40264 (N_40264,N_38708,N_39764);
or U40265 (N_40265,N_38617,N_39436);
xor U40266 (N_40266,N_39315,N_39800);
nand U40267 (N_40267,N_39387,N_38520);
and U40268 (N_40268,N_39166,N_39828);
or U40269 (N_40269,N_39739,N_38177);
nand U40270 (N_40270,N_39306,N_39987);
xnor U40271 (N_40271,N_38772,N_39413);
nand U40272 (N_40272,N_38168,N_38299);
nand U40273 (N_40273,N_38840,N_38894);
nand U40274 (N_40274,N_39225,N_39310);
and U40275 (N_40275,N_38907,N_39814);
nor U40276 (N_40276,N_39578,N_39129);
or U40277 (N_40277,N_39841,N_38202);
nor U40278 (N_40278,N_38848,N_38394);
nor U40279 (N_40279,N_38167,N_38518);
or U40280 (N_40280,N_38501,N_39598);
and U40281 (N_40281,N_39992,N_38047);
xnor U40282 (N_40282,N_39559,N_38578);
or U40283 (N_40283,N_38655,N_39282);
xnor U40284 (N_40284,N_38996,N_39153);
nand U40285 (N_40285,N_38629,N_38471);
and U40286 (N_40286,N_39473,N_39080);
or U40287 (N_40287,N_39695,N_38703);
nor U40288 (N_40288,N_38783,N_39456);
nand U40289 (N_40289,N_39716,N_39355);
xor U40290 (N_40290,N_38650,N_39434);
and U40291 (N_40291,N_38317,N_39043);
nor U40292 (N_40292,N_39544,N_38106);
or U40293 (N_40293,N_38005,N_38728);
and U40294 (N_40294,N_38750,N_39407);
and U40295 (N_40295,N_38252,N_38260);
or U40296 (N_40296,N_38786,N_39797);
nand U40297 (N_40297,N_38571,N_39150);
or U40298 (N_40298,N_39443,N_38042);
or U40299 (N_40299,N_38450,N_39337);
xor U40300 (N_40300,N_39729,N_38551);
nand U40301 (N_40301,N_38736,N_39644);
nand U40302 (N_40302,N_38651,N_39496);
or U40303 (N_40303,N_38108,N_39455);
and U40304 (N_40304,N_38344,N_39531);
xor U40305 (N_40305,N_39479,N_38402);
and U40306 (N_40306,N_38267,N_39348);
and U40307 (N_40307,N_39638,N_38702);
nor U40308 (N_40308,N_38075,N_39915);
nand U40309 (N_40309,N_39954,N_38404);
and U40310 (N_40310,N_38885,N_38614);
nor U40311 (N_40311,N_39230,N_38936);
or U40312 (N_40312,N_39290,N_39624);
xor U40313 (N_40313,N_39612,N_38601);
nor U40314 (N_40314,N_39794,N_39761);
nand U40315 (N_40315,N_38850,N_38526);
xor U40316 (N_40316,N_39146,N_39871);
and U40317 (N_40317,N_39516,N_38435);
or U40318 (N_40318,N_39267,N_39163);
nor U40319 (N_40319,N_39213,N_39601);
or U40320 (N_40320,N_39567,N_39289);
nand U40321 (N_40321,N_39061,N_39533);
and U40322 (N_40322,N_39742,N_38018);
nand U40323 (N_40323,N_39321,N_38090);
nand U40324 (N_40324,N_39047,N_38281);
nor U40325 (N_40325,N_38628,N_38351);
nand U40326 (N_40326,N_38538,N_39030);
xnor U40327 (N_40327,N_38710,N_39651);
xnor U40328 (N_40328,N_39523,N_39648);
xor U40329 (N_40329,N_38992,N_39249);
and U40330 (N_40330,N_39420,N_38534);
nand U40331 (N_40331,N_38744,N_38256);
nand U40332 (N_40332,N_39563,N_39374);
xnor U40333 (N_40333,N_39682,N_38500);
xor U40334 (N_40334,N_39200,N_38831);
nor U40335 (N_40335,N_38401,N_39897);
nor U40336 (N_40336,N_39775,N_38929);
or U40337 (N_40337,N_39167,N_38243);
nor U40338 (N_40338,N_39099,N_39313);
and U40339 (N_40339,N_38102,N_38590);
or U40340 (N_40340,N_39965,N_38564);
or U40341 (N_40341,N_39464,N_39101);
and U40342 (N_40342,N_38245,N_39020);
xnor U40343 (N_40343,N_38300,N_38131);
nor U40344 (N_40344,N_39112,N_38675);
xor U40345 (N_40345,N_38414,N_39835);
or U40346 (N_40346,N_39844,N_38778);
nand U40347 (N_40347,N_39450,N_39300);
or U40348 (N_40348,N_39874,N_38040);
and U40349 (N_40349,N_39518,N_38689);
xor U40350 (N_40350,N_39958,N_38012);
and U40351 (N_40351,N_39339,N_38494);
and U40352 (N_40352,N_39957,N_38492);
xor U40353 (N_40353,N_39109,N_38120);
and U40354 (N_40354,N_38236,N_39115);
nor U40355 (N_40355,N_39096,N_39016);
or U40356 (N_40356,N_39918,N_39215);
nand U40357 (N_40357,N_39475,N_39162);
and U40358 (N_40358,N_39470,N_39363);
or U40359 (N_40359,N_38639,N_39852);
and U40360 (N_40360,N_39888,N_38061);
and U40361 (N_40361,N_39147,N_38346);
or U40362 (N_40362,N_38070,N_39024);
nor U40363 (N_40363,N_38325,N_38606);
or U40364 (N_40364,N_38531,N_38493);
xor U40365 (N_40365,N_39500,N_39357);
or U40366 (N_40366,N_39476,N_39157);
xnor U40367 (N_40367,N_38770,N_38221);
nor U40368 (N_40368,N_39876,N_39254);
and U40369 (N_40369,N_38088,N_38464);
nand U40370 (N_40370,N_38368,N_39604);
or U40371 (N_40371,N_38459,N_39107);
nand U40372 (N_40372,N_39639,N_38762);
nor U40373 (N_40373,N_38503,N_39573);
and U40374 (N_40374,N_38463,N_38923);
nor U40375 (N_40375,N_39960,N_38809);
and U40376 (N_40376,N_38110,N_38263);
and U40377 (N_40377,N_38248,N_38565);
or U40378 (N_40378,N_38007,N_39929);
and U40379 (N_40379,N_38083,N_39833);
and U40380 (N_40380,N_38863,N_39595);
or U40381 (N_40381,N_39849,N_39462);
nor U40382 (N_40382,N_39486,N_38593);
or U40383 (N_40383,N_39937,N_38654);
or U40384 (N_40384,N_39171,N_39314);
and U40385 (N_40385,N_39934,N_39360);
nor U40386 (N_40386,N_38800,N_38295);
or U40387 (N_40387,N_38700,N_39121);
nand U40388 (N_40388,N_38002,N_38592);
nand U40389 (N_40389,N_39825,N_38289);
xnor U40390 (N_40390,N_38031,N_38465);
nor U40391 (N_40391,N_39205,N_38610);
nand U40392 (N_40392,N_39296,N_38706);
nor U40393 (N_40393,N_38516,N_38392);
or U40394 (N_40394,N_38297,N_39606);
xnor U40395 (N_40395,N_38946,N_38361);
xor U40396 (N_40396,N_39968,N_38447);
or U40397 (N_40397,N_38683,N_39893);
nor U40398 (N_40398,N_38927,N_39483);
and U40399 (N_40399,N_38370,N_39801);
nor U40400 (N_40400,N_38561,N_38119);
nand U40401 (N_40401,N_39381,N_39375);
nand U40402 (N_40402,N_39820,N_39579);
xor U40403 (N_40403,N_39116,N_38645);
or U40404 (N_40404,N_38046,N_39057);
nor U40405 (N_40405,N_39466,N_38909);
xor U40406 (N_40406,N_39372,N_38373);
nand U40407 (N_40407,N_38624,N_38916);
nand U40408 (N_40408,N_39665,N_39574);
nand U40409 (N_40409,N_38235,N_39566);
nand U40410 (N_40410,N_39233,N_39334);
xor U40411 (N_40411,N_39014,N_39100);
nor U40412 (N_40412,N_38910,N_38126);
and U40413 (N_40413,N_39660,N_39913);
or U40414 (N_40414,N_39089,N_39452);
or U40415 (N_40415,N_39542,N_38335);
nand U40416 (N_40416,N_39053,N_38583);
nand U40417 (N_40417,N_39428,N_38719);
and U40418 (N_40418,N_39133,N_38353);
nor U40419 (N_40419,N_38348,N_39626);
nand U40420 (N_40420,N_39478,N_39256);
or U40421 (N_40421,N_38214,N_38781);
xnor U40422 (N_40422,N_38477,N_39774);
xnor U40423 (N_40423,N_39224,N_39830);
nor U40424 (N_40424,N_39149,N_39786);
nor U40425 (N_40425,N_38918,N_39599);
or U40426 (N_40426,N_39845,N_38315);
xnor U40427 (N_40427,N_39654,N_38422);
nand U40428 (N_40428,N_39610,N_38919);
and U40429 (N_40429,N_39693,N_38741);
nand U40430 (N_40430,N_39850,N_38444);
xnor U40431 (N_40431,N_39932,N_39134);
nor U40432 (N_40432,N_38406,N_38457);
xnor U40433 (N_40433,N_39760,N_38200);
nand U40434 (N_40434,N_38160,N_38359);
or U40435 (N_40435,N_38664,N_38331);
nand U40436 (N_40436,N_38013,N_38817);
xnor U40437 (N_40437,N_38816,N_38172);
and U40438 (N_40438,N_39587,N_39195);
nor U40439 (N_40439,N_38292,N_38727);
nor U40440 (N_40440,N_39414,N_38532);
or U40441 (N_40441,N_39160,N_39105);
xnor U40442 (N_40442,N_39527,N_38287);
xnor U40443 (N_40443,N_38478,N_38753);
and U40444 (N_40444,N_38307,N_38174);
nand U40445 (N_40445,N_38815,N_38205);
xnor U40446 (N_40446,N_39633,N_39539);
and U40447 (N_40447,N_38636,N_39010);
nand U40448 (N_40448,N_39265,N_39076);
and U40449 (N_40449,N_39004,N_38397);
nor U40450 (N_40450,N_38712,N_39324);
xor U40451 (N_40451,N_39967,N_39035);
and U40452 (N_40452,N_38978,N_38724);
xor U40453 (N_40453,N_39447,N_38533);
or U40454 (N_40454,N_38165,N_39091);
nor U40455 (N_40455,N_39583,N_38431);
xnor U40456 (N_40456,N_39551,N_39590);
and U40457 (N_40457,N_39749,N_38818);
or U40458 (N_40458,N_38642,N_38044);
nor U40459 (N_40459,N_38355,N_39180);
xnor U40460 (N_40460,N_39504,N_38425);
xnor U40461 (N_40461,N_39380,N_39045);
xnor U40462 (N_40462,N_39085,N_39517);
or U40463 (N_40463,N_39124,N_38113);
and U40464 (N_40464,N_38588,N_38458);
nand U40465 (N_40465,N_38198,N_38694);
or U40466 (N_40466,N_38861,N_38421);
nand U40467 (N_40467,N_39094,N_38237);
xor U40468 (N_40468,N_38972,N_38541);
nor U40469 (N_40469,N_38382,N_39439);
nand U40470 (N_40470,N_38731,N_38739);
nand U40471 (N_40471,N_38231,N_39395);
xor U40472 (N_40472,N_38449,N_38917);
nor U40473 (N_40473,N_38175,N_39400);
xor U40474 (N_40474,N_39364,N_39956);
and U40475 (N_40475,N_39565,N_38569);
xnor U40476 (N_40476,N_38802,N_39351);
nand U40477 (N_40477,N_39275,N_39454);
xor U40478 (N_40478,N_38383,N_38399);
nor U40479 (N_40479,N_39093,N_39329);
xor U40480 (N_40480,N_38304,N_39495);
or U40481 (N_40481,N_38015,N_39262);
nor U40482 (N_40482,N_39719,N_38058);
xor U40483 (N_40483,N_39706,N_39911);
xor U40484 (N_40484,N_39365,N_38212);
or U40485 (N_40485,N_38389,N_38613);
xnor U40486 (N_40486,N_38242,N_38743);
or U40487 (N_40487,N_38934,N_39727);
xor U40488 (N_40488,N_39687,N_39895);
xnor U40489 (N_40489,N_39044,N_38900);
xnor U40490 (N_40490,N_39705,N_38037);
nand U40491 (N_40491,N_39005,N_39366);
nor U40492 (N_40492,N_39070,N_39319);
nor U40493 (N_40493,N_39155,N_38513);
nor U40494 (N_40494,N_38574,N_39908);
and U40495 (N_40495,N_39402,N_39458);
nand U40496 (N_40496,N_38790,N_38259);
xnor U40497 (N_40497,N_39323,N_38767);
nor U40498 (N_40498,N_38858,N_39634);
nor U40499 (N_40499,N_38143,N_38521);
nand U40500 (N_40500,N_39702,N_39181);
xnor U40501 (N_40501,N_38998,N_39415);
and U40502 (N_40502,N_39425,N_38312);
nor U40503 (N_40503,N_38216,N_38311);
nand U40504 (N_40504,N_38011,N_38514);
and U40505 (N_40505,N_39582,N_38991);
and U40506 (N_40506,N_38386,N_39972);
nand U40507 (N_40507,N_38436,N_38875);
xnor U40508 (N_40508,N_39873,N_38953);
nor U40509 (N_40509,N_38987,N_39944);
xor U40510 (N_40510,N_39191,N_38417);
nor U40511 (N_40511,N_38320,N_39993);
or U40512 (N_40512,N_39103,N_38705);
xnor U40513 (N_40513,N_39907,N_39266);
xor U40514 (N_40514,N_39678,N_38616);
nand U40515 (N_40515,N_38522,N_39617);
xor U40516 (N_40516,N_39312,N_38568);
or U40517 (N_40517,N_38886,N_38104);
and U40518 (N_40518,N_39240,N_39145);
and U40519 (N_40519,N_39514,N_38329);
nand U40520 (N_40520,N_39744,N_39722);
nand U40521 (N_40521,N_38515,N_38163);
nor U40522 (N_40522,N_38956,N_38366);
xnor U40523 (N_40523,N_39949,N_39540);
nand U40524 (N_40524,N_39832,N_39730);
nand U40525 (N_40525,N_38887,N_39602);
nand U40526 (N_40526,N_39667,N_39386);
nor U40527 (N_40527,N_38272,N_39931);
and U40528 (N_40528,N_39674,N_38864);
and U40529 (N_40529,N_39488,N_39431);
or U40530 (N_40530,N_38218,N_39538);
and U40531 (N_40531,N_38673,N_39221);
or U40532 (N_40532,N_38302,N_39183);
nand U40533 (N_40533,N_39826,N_39097);
and U40534 (N_40534,N_39244,N_38687);
and U40535 (N_40535,N_38859,N_39962);
nand U40536 (N_40536,N_38804,N_38951);
xnor U40537 (N_40537,N_38085,N_39941);
nor U40538 (N_40538,N_38238,N_38045);
and U40539 (N_40539,N_39114,N_38298);
nor U40540 (N_40540,N_38137,N_39229);
nand U40541 (N_40541,N_39461,N_38232);
nor U40542 (N_40542,N_39137,N_39788);
nand U40543 (N_40543,N_39717,N_39318);
nand U40544 (N_40544,N_39738,N_38847);
or U40545 (N_40545,N_39188,N_38187);
nor U40546 (N_40546,N_39013,N_38074);
nand U40547 (N_40547,N_38068,N_39273);
and U40548 (N_40548,N_38054,N_38189);
and U40549 (N_40549,N_38920,N_38667);
or U40550 (N_40550,N_38509,N_39734);
and U40551 (N_40551,N_38358,N_39762);
xor U40552 (N_40552,N_38363,N_38908);
xnor U40553 (N_40553,N_39545,N_39552);
xor U40554 (N_40554,N_38322,N_39304);
nor U40555 (N_40555,N_39293,N_38369);
xnor U40556 (N_40556,N_38239,N_39127);
nand U40557 (N_40557,N_38153,N_39332);
nand U40558 (N_40558,N_38902,N_38584);
xor U40559 (N_40559,N_39681,N_39060);
nor U40560 (N_40560,N_38112,N_38453);
or U40561 (N_40561,N_38326,N_38756);
or U40562 (N_40562,N_39135,N_39536);
nor U40563 (N_40563,N_38387,N_39721);
and U40564 (N_40564,N_38576,N_38969);
xor U40565 (N_40565,N_39655,N_39819);
nand U40566 (N_40566,N_39268,N_38249);
nand U40567 (N_40567,N_39356,N_38283);
or U40568 (N_40568,N_38188,N_38897);
and U40569 (N_40569,N_39172,N_39715);
nand U40570 (N_40570,N_39067,N_38284);
xor U40571 (N_40571,N_38722,N_39827);
nor U40572 (N_40572,N_39477,N_38121);
or U40573 (N_40573,N_39298,N_38388);
and U40574 (N_40574,N_38446,N_38294);
or U40575 (N_40575,N_39869,N_38843);
nor U40576 (N_40576,N_38553,N_39643);
or U40577 (N_40577,N_39656,N_39880);
nor U40578 (N_40578,N_38766,N_39821);
nand U40579 (N_40579,N_38674,N_39404);
xnor U40580 (N_40580,N_39338,N_38423);
nor U40581 (N_40581,N_39570,N_39892);
nand U40582 (N_40582,N_38620,N_38844);
xnor U40583 (N_40583,N_39785,N_39791);
nand U40584 (N_40584,N_39170,N_39291);
nor U40585 (N_40585,N_38924,N_39983);
or U40586 (N_40586,N_39056,N_39971);
nand U40587 (N_40587,N_38139,N_39703);
and U40588 (N_40588,N_39697,N_39226);
and U40589 (N_40589,N_38266,N_39688);
xnor U40590 (N_40590,N_38649,N_39509);
nor U40591 (N_40591,N_38081,N_39714);
nand U40592 (N_40592,N_39263,N_39350);
and U40593 (N_40593,N_38837,N_39440);
xnor U40594 (N_40594,N_38697,N_38038);
xnor U40595 (N_40595,N_38173,N_38171);
nand U40596 (N_40596,N_38747,N_39342);
and U40597 (N_40597,N_38251,N_39088);
nand U40598 (N_40598,N_39669,N_38485);
nand U40599 (N_40599,N_38407,N_38988);
xor U40600 (N_40600,N_39988,N_38103);
or U40601 (N_40601,N_38123,N_39449);
and U40602 (N_40602,N_38646,N_38487);
or U40603 (N_40603,N_38162,N_38087);
nor U40604 (N_40604,N_39884,N_38470);
nor U40605 (N_40605,N_39320,N_38197);
and U40606 (N_40606,N_38994,N_38832);
nor U40607 (N_40607,N_39165,N_39748);
xnor U40608 (N_40608,N_38262,N_39822);
nor U40609 (N_40609,N_39887,N_38296);
and U40610 (N_40610,N_39027,N_39746);
xor U40611 (N_40611,N_38644,N_39878);
nand U40612 (N_40612,N_39927,N_38723);
or U40613 (N_40613,N_39484,N_38180);
nand U40614 (N_40614,N_38550,N_38641);
nor U40615 (N_40615,N_39442,N_39117);
or U40616 (N_40616,N_39237,N_39591);
nor U40617 (N_40617,N_39641,N_39554);
and U40618 (N_40618,N_38828,N_39253);
and U40619 (N_40619,N_38357,N_38699);
or U40620 (N_40620,N_39487,N_39354);
and U40621 (N_40621,N_39900,N_38797);
xor U40622 (N_40622,N_38508,N_38880);
and U40623 (N_40623,N_38483,N_39817);
or U40624 (N_40624,N_39033,N_38637);
nand U40625 (N_40625,N_39779,N_38865);
xor U40626 (N_40626,N_39411,N_39264);
or U40627 (N_40627,N_38016,N_38008);
or U40628 (N_40628,N_38445,N_38995);
xor U40629 (N_40629,N_38362,N_39846);
or U40630 (N_40630,N_38547,N_39468);
and U40631 (N_40631,N_39054,N_38949);
and U40632 (N_40632,N_38408,N_39152);
or U40633 (N_40633,N_39611,N_38672);
nand U40634 (N_40634,N_39653,N_38554);
and U40635 (N_40635,N_38733,N_39803);
xnor U40636 (N_40636,N_38134,N_38849);
nand U40637 (N_40637,N_38128,N_39283);
and U40638 (N_40638,N_38676,N_39141);
xor U40639 (N_40639,N_39875,N_39771);
nand U40640 (N_40640,N_38282,N_38801);
and U40641 (N_40641,N_39964,N_38925);
nor U40642 (N_40642,N_39560,N_38609);
nor U40643 (N_40643,N_38922,N_38715);
and U40644 (N_40644,N_39613,N_39942);
xnor U40645 (N_40645,N_38491,N_38378);
or U40646 (N_40646,N_39556,N_38079);
and U40647 (N_40647,N_39690,N_39919);
nand U40648 (N_40648,N_38314,N_39754);
nor U40649 (N_40649,N_38203,N_38967);
nor U40650 (N_40650,N_39346,N_39933);
and U40651 (N_40651,N_38656,N_39662);
xor U40652 (N_40652,N_39977,N_39489);
and U40653 (N_40653,N_39490,N_39696);
nand U40654 (N_40654,N_38573,N_39219);
or U40655 (N_40655,N_39071,N_39999);
or U40656 (N_40656,N_39889,N_38813);
nand U40657 (N_40657,N_39023,N_39438);
nor U40658 (N_40658,N_38653,N_38877);
nor U40659 (N_40659,N_38681,N_38122);
or U40660 (N_40660,N_38050,N_39242);
and U40661 (N_40661,N_39001,N_38286);
or U40662 (N_40662,N_39408,N_38869);
and U40663 (N_40663,N_38567,N_38321);
or U40664 (N_40664,N_38063,N_38116);
or U40665 (N_40665,N_39741,N_38035);
nor U40666 (N_40666,N_39008,N_39548);
and U40667 (N_40667,N_38086,N_39629);
nand U40668 (N_40668,N_38490,N_38274);
nand U40669 (N_40669,N_39615,N_38669);
nand U40670 (N_40670,N_38961,N_39914);
and U40671 (N_40671,N_38851,N_38707);
nand U40672 (N_40672,N_38060,N_39507);
nand U40673 (N_40673,N_38901,N_38622);
nand U40674 (N_40674,N_39809,N_39745);
nor U40675 (N_40675,N_38141,N_38030);
nand U40676 (N_40676,N_39953,N_39994);
or U40677 (N_40677,N_39410,N_39663);
nor U40678 (N_40678,N_39148,N_39406);
nor U40679 (N_40679,N_38732,N_38939);
or U40680 (N_40680,N_39906,N_38761);
xor U40681 (N_40681,N_38730,N_39151);
nor U40682 (N_40682,N_38777,N_38240);
nand U40683 (N_40683,N_39308,N_38630);
or U40684 (N_40684,N_38489,N_39823);
nand U40685 (N_40685,N_38330,N_39747);
xor U40686 (N_40686,N_38975,N_38337);
and U40687 (N_40687,N_39359,N_39471);
xor U40688 (N_40688,N_38974,N_38898);
or U40689 (N_40689,N_38158,N_39493);
and U40690 (N_40690,N_38196,N_39081);
xor U40691 (N_40691,N_39963,N_38814);
and U40692 (N_40692,N_38291,N_39126);
nor U40693 (N_40693,N_39902,N_39707);
and U40694 (N_40694,N_38822,N_39753);
nor U40695 (N_40695,N_38468,N_38496);
nor U40696 (N_40696,N_39592,N_38537);
nor U40697 (N_40697,N_38701,N_38912);
and U40698 (N_40698,N_39922,N_38277);
or U40699 (N_40699,N_38268,N_38495);
xor U40700 (N_40700,N_38945,N_38714);
nand U40701 (N_40701,N_38223,N_39158);
or U40702 (N_40702,N_39184,N_38275);
and U40703 (N_40703,N_38935,N_38638);
or U40704 (N_40704,N_38981,N_39783);
nand U40705 (N_40705,N_38019,N_38787);
and U40706 (N_40706,N_39799,N_38365);
xor U40707 (N_40707,N_39007,N_39078);
and U40708 (N_40708,N_38933,N_39175);
and U40709 (N_40709,N_38233,N_38690);
nand U40710 (N_40710,N_39798,N_38179);
or U40711 (N_40711,N_39955,N_38726);
nand U40712 (N_40712,N_39095,N_38842);
xor U40713 (N_40713,N_39623,N_38581);
nor U40714 (N_40714,N_38342,N_39792);
nor U40715 (N_40715,N_38095,N_39426);
nor U40716 (N_40716,N_38145,N_39223);
and U40717 (N_40717,N_38985,N_38717);
and U40718 (N_40718,N_39824,N_39519);
xnor U40719 (N_40719,N_39732,N_38066);
nor U40720 (N_40720,N_39396,N_38448);
nor U40721 (N_40721,N_38746,N_39110);
nand U40722 (N_40722,N_39119,N_39326);
nand U40723 (N_40723,N_39812,N_38474);
or U40724 (N_40724,N_38824,N_39731);
or U40725 (N_40725,N_38666,N_39710);
nand U40726 (N_40726,N_39258,N_38479);
and U40727 (N_40727,N_39385,N_39222);
nor U40728 (N_40728,N_39763,N_38183);
or U40729 (N_40729,N_39190,N_38146);
or U40730 (N_40730,N_39453,N_39353);
or U40731 (N_40731,N_39616,N_38148);
nor U40732 (N_40732,N_39260,N_39837);
or U40733 (N_40733,N_39341,N_39064);
xnor U40734 (N_40734,N_39235,N_38352);
nand U40735 (N_40735,N_38668,N_39916);
and U40736 (N_40736,N_38345,N_39780);
nand U40737 (N_40737,N_39084,N_38659);
nand U40738 (N_40738,N_39006,N_39818);
and U40739 (N_40739,N_38100,N_38586);
nor U40740 (N_40740,N_39278,N_39581);
nand U40741 (N_40741,N_39295,N_38857);
nor U40742 (N_40742,N_38065,N_38539);
and U40743 (N_40743,N_38390,N_39584);
xor U40744 (N_40744,N_39652,N_38301);
xnor U40745 (N_40745,N_39206,N_39336);
nor U40746 (N_40746,N_39720,N_38454);
nand U40747 (N_40747,N_38206,N_38253);
nor U40748 (N_40748,N_38170,N_39646);
nor U40749 (N_40749,N_38130,N_39758);
or U40750 (N_40750,N_39860,N_38826);
nand U40751 (N_40751,N_38293,N_38280);
nor U40752 (N_40752,N_39427,N_38685);
xnor U40753 (N_40753,N_38056,N_39981);
or U40754 (N_40754,N_39843,N_38955);
xnor U40755 (N_40755,N_38627,N_38118);
or U40756 (N_40756,N_38693,N_39569);
and U40757 (N_40757,N_38990,N_38021);
nand U40758 (N_40758,N_38579,N_38904);
nand U40759 (N_40759,N_38254,N_38204);
or U40760 (N_40760,N_39073,N_38381);
nand U40761 (N_40761,N_39423,N_38328);
and U40762 (N_40762,N_39174,N_39042);
xnor U40763 (N_40763,N_38535,N_39894);
nor U40764 (N_40764,N_39292,N_38416);
or U40765 (N_40765,N_38288,N_38316);
or U40766 (N_40766,N_38796,N_38003);
nor U40767 (N_40767,N_39541,N_38711);
and U40768 (N_40768,N_38078,N_38409);
and U40769 (N_40769,N_39537,N_38677);
nor U40770 (N_40770,N_38469,N_39943);
or U40771 (N_40771,N_38577,N_39187);
and U40772 (N_40772,N_38871,N_39759);
and U40773 (N_40773,N_39102,N_38965);
or U40774 (N_40774,N_38109,N_39947);
nand U40775 (N_40775,N_39765,N_39139);
or U40776 (N_40776,N_39140,N_38608);
nand U40777 (N_40777,N_39383,N_39288);
xnor U40778 (N_40778,N_39940,N_38941);
and U40779 (N_40779,N_39419,N_39621);
xnor U40780 (N_40780,N_39946,N_38014);
xor U40781 (N_40781,N_38954,N_39555);
or U40782 (N_40782,N_39433,N_38589);
nand U40783 (N_40783,N_39451,N_38217);
nand U40784 (N_40784,N_39576,N_38963);
or U40785 (N_40785,N_39063,N_38219);
or U40786 (N_40786,N_39970,N_38455);
and U40787 (N_40787,N_39831,N_38089);
nor U40788 (N_40788,N_38270,N_38082);
nand U40789 (N_40789,N_38097,N_39340);
nor U40790 (N_40790,N_38201,N_38451);
nand U40791 (N_40791,N_38151,N_38595);
and U40792 (N_40792,N_38993,N_39113);
nand U40793 (N_40793,N_38499,N_39474);
nor U40794 (N_40794,N_38334,N_39948);
nand U40795 (N_40795,N_39485,N_39397);
nor U40796 (N_40796,N_39384,N_38836);
nand U40797 (N_40797,N_38774,N_39829);
nand U40798 (N_40798,N_38555,N_38845);
nor U40799 (N_40799,N_39924,N_38420);
or U40800 (N_40800,N_39281,N_38895);
or U40801 (N_40801,N_39776,N_38462);
nand U40802 (N_40802,N_39990,N_39087);
nand U40803 (N_40803,N_39737,N_39699);
nand U40804 (N_40804,N_39199,N_38072);
or U40805 (N_40805,N_39580,N_39301);
nand U40806 (N_40806,N_39128,N_38306);
nor U40807 (N_40807,N_39122,N_38227);
nor U40808 (N_40808,N_39679,N_38602);
xnor U40809 (N_40809,N_39210,N_39203);
xor U40810 (N_40810,N_38545,N_39898);
xnor U40811 (N_40811,N_38419,N_39176);
or U40812 (N_40812,N_38979,N_39376);
xor U40813 (N_40813,N_38695,N_38229);
xnor U40814 (N_40814,N_38748,N_39564);
xnor U40815 (N_40815,N_38154,N_39211);
or U40816 (N_40816,N_38052,N_38393);
nor U40817 (N_40817,N_39274,N_38799);
xnor U40818 (N_40818,N_38184,N_38735);
or U40819 (N_40819,N_39625,N_38350);
xnor U40820 (N_40820,N_39398,N_38626);
xnor U40821 (N_40821,N_38418,N_39065);
nand U40822 (N_40822,N_38517,N_38889);
xor U40823 (N_40823,N_39098,N_39231);
xnor U40824 (N_40824,N_38906,N_38926);
nor U40825 (N_40825,N_38133,N_39593);
nor U40826 (N_40826,N_39680,N_38856);
and U40827 (N_40827,N_39577,N_39777);
nor U40828 (N_40828,N_39618,N_38671);
xor U40829 (N_40829,N_38157,N_39207);
nor U40830 (N_40830,N_39815,N_39982);
nand U40831 (N_40831,N_39204,N_38921);
nand U40832 (N_40832,N_39416,N_39018);
xnor U40833 (N_40833,N_38024,N_39390);
xor U40834 (N_40834,N_39448,N_39740);
xor U40835 (N_40835,N_38149,N_38604);
or U40836 (N_40836,N_38466,N_38692);
and U40837 (N_40837,N_38258,N_39513);
and U40838 (N_40838,N_38138,N_38308);
nand U40839 (N_40839,N_38319,N_39038);
nand U40840 (N_40840,N_38903,N_38721);
and U40841 (N_40841,N_39525,N_38036);
nand U40842 (N_40842,N_39603,N_39299);
nor U40843 (N_40843,N_38434,N_38246);
nor U40844 (N_40844,N_38968,N_39378);
nor U40845 (N_40845,N_39698,N_39708);
xnor U40846 (N_40846,N_38855,N_38333);
nor U40847 (N_40847,N_39510,N_38552);
nand U40848 (N_40848,N_39370,N_38405);
or U40849 (N_40849,N_38870,N_39270);
nor U40850 (N_40850,N_39713,N_39029);
nand U40851 (N_40851,N_38760,N_39575);
or U40852 (N_40852,N_38582,N_39664);
or U40853 (N_40853,N_38758,N_39352);
xnor U40854 (N_40854,N_38208,N_39904);
or U40855 (N_40855,N_39980,N_38942);
or U40856 (N_40856,N_38964,N_39309);
xnor U40857 (N_40857,N_38560,N_38213);
or U40858 (N_40858,N_38371,N_38285);
and U40859 (N_40859,N_38841,N_39472);
xnor U40860 (N_40860,N_38480,N_39839);
xnor U40861 (N_40861,N_39627,N_39394);
xnor U40862 (N_40862,N_39985,N_38364);
or U40863 (N_40863,N_39212,N_39683);
or U40864 (N_40864,N_39034,N_39369);
or U40865 (N_40865,N_38099,N_38530);
nand U40866 (N_40866,N_39769,N_39991);
or U40867 (N_40867,N_39808,N_38209);
and U40868 (N_40868,N_38612,N_39666);
nor U40869 (N_40869,N_38437,N_38255);
and U40870 (N_40870,N_38830,N_39684);
nand U40871 (N_40871,N_39521,N_39022);
xor U40872 (N_40872,N_38603,N_38971);
nor U40873 (N_40873,N_38505,N_38519);
and U40874 (N_40874,N_38424,N_39859);
xnor U40875 (N_40875,N_38456,N_38745);
and U40876 (N_40876,N_38323,N_38241);
nor U40877 (N_40877,N_39686,N_39092);
and U40878 (N_40878,N_39040,N_39202);
and U40879 (N_40879,N_39505,N_39650);
and U40880 (N_40880,N_38811,N_38853);
and U40881 (N_40881,N_38053,N_38432);
and U40882 (N_40882,N_38635,N_39659);
or U40883 (N_40883,N_38049,N_38594);
or U40884 (N_40884,N_39810,N_39685);
and U40885 (N_40885,N_39870,N_39553);
xor U40886 (N_40886,N_38159,N_38599);
and U40887 (N_40887,N_38838,N_39362);
nor U40888 (N_40888,N_39228,N_39989);
and U40889 (N_40889,N_38528,N_38989);
or U40890 (N_40890,N_38155,N_38882);
xor U40891 (N_40891,N_38472,N_38782);
nand U40892 (N_40892,N_39220,N_39297);
and U40893 (N_40893,N_38866,N_38829);
xnor U40894 (N_40894,N_38093,N_39017);
xnor U40895 (N_40895,N_38481,N_38339);
nor U40896 (N_40896,N_39959,N_39735);
and U40897 (N_40897,N_39469,N_39136);
or U40898 (N_40898,N_38349,N_38928);
xor U40899 (N_40899,N_39015,N_38132);
xor U40900 (N_40900,N_38341,N_38852);
nor U40901 (N_40901,N_38948,N_39772);
xor U40902 (N_40902,N_39236,N_39435);
or U40903 (N_40903,N_39805,N_39847);
nor U40904 (N_40904,N_38839,N_39049);
nor U40905 (N_40905,N_39059,N_39756);
xor U40906 (N_40906,N_39787,N_38825);
or U40907 (N_40907,N_39432,N_39201);
nor U40908 (N_40908,N_38890,N_38411);
nand U40909 (N_40909,N_38868,N_39770);
nor U40910 (N_40910,N_39409,N_38136);
nor U40911 (N_40911,N_39130,N_39557);
nor U40912 (N_40912,N_39975,N_38957);
or U40913 (N_40913,N_38834,N_38488);
or U40914 (N_40914,N_38580,N_39515);
xor U40915 (N_40915,N_39851,N_38633);
and U40916 (N_40916,N_39921,N_38543);
xnor U40917 (N_40917,N_39673,N_38433);
nand U40918 (N_40918,N_39052,N_38190);
xor U40919 (N_40919,N_39000,N_39039);
nand U40920 (N_40920,N_39842,N_38502);
nor U40921 (N_40921,N_39325,N_39294);
and U40922 (N_40922,N_39945,N_38600);
and U40923 (N_40923,N_38234,N_38625);
or U40924 (N_40924,N_38336,N_38347);
nor U40925 (N_40925,N_39271,N_38461);
nor U40926 (N_40926,N_38892,N_38980);
and U40927 (N_40927,N_39062,N_39156);
nand U40928 (N_40928,N_38129,N_39143);
xor U40929 (N_40929,N_38771,N_38915);
nor U40930 (N_40930,N_38441,N_39782);
or U40931 (N_40931,N_39412,N_38952);
and U40932 (N_40932,N_38984,N_39316);
nand U40933 (N_40933,N_39169,N_39197);
nand U40934 (N_40934,N_38872,N_38572);
nand U40935 (N_40935,N_38794,N_38161);
nand U40936 (N_40936,N_39807,N_38111);
nor U40937 (N_40937,N_38305,N_38017);
xnor U40938 (N_40938,N_39259,N_38023);
nand U40939 (N_40939,N_39104,N_38631);
or U40940 (N_40940,N_39041,N_39864);
and U40941 (N_40941,N_38230,N_39465);
and U40942 (N_40942,N_39344,N_39951);
nand U40943 (N_40943,N_38821,N_39403);
or U40944 (N_40944,N_39002,N_38938);
nor U40945 (N_40945,N_39379,N_39179);
and U40946 (N_40946,N_38899,N_38091);
nand U40947 (N_40947,N_38497,N_38737);
xnor U40948 (N_40948,N_38048,N_38621);
and U40949 (N_40949,N_38033,N_39998);
nand U40950 (N_40950,N_39718,N_39804);
or U40951 (N_40951,N_38156,N_39074);
or U40952 (N_40952,N_38691,N_39028);
and U40953 (N_40953,N_38094,N_38476);
nor U40954 (N_40954,N_39025,N_39920);
xor U40955 (N_40955,N_39790,N_39724);
or U40956 (N_40956,N_38410,N_38523);
xnor U40957 (N_40957,N_39671,N_38718);
xor U40958 (N_40958,N_39811,N_39858);
and U40959 (N_40959,N_38396,N_38680);
xor U40960 (N_40960,N_39177,N_38185);
nand U40961 (N_40961,N_38228,N_39399);
nor U40962 (N_40962,N_38931,N_38725);
or U40963 (N_40963,N_39642,N_38498);
nand U40964 (N_40964,N_39973,N_38930);
xor U40965 (N_40965,N_38575,N_39978);
nor U40966 (N_40966,N_39269,N_38222);
nor U40967 (N_40967,N_38318,N_38823);
xor U40968 (N_40968,N_39164,N_38114);
nand U40969 (N_40969,N_38181,N_38028);
nand U40970 (N_40970,N_38178,N_39723);
nor U40971 (N_40971,N_38959,N_39640);
and U40972 (N_40972,N_38874,N_39037);
nor U40973 (N_40973,N_38559,N_38473);
or U40974 (N_40974,N_38027,N_38776);
nand U40975 (N_40975,N_38966,N_39467);
or U40976 (N_40976,N_39767,N_39444);
and U40977 (N_40977,N_39632,N_39280);
or U40978 (N_40978,N_39055,N_39986);
xor U40979 (N_40979,N_38970,N_38914);
xnor U40980 (N_40980,N_38763,N_38403);
and U40981 (N_40981,N_39547,N_39836);
and U40982 (N_40982,N_39520,N_38806);
or U40983 (N_40983,N_39726,N_39736);
or U40984 (N_40984,N_38022,N_39009);
and U40985 (N_40985,N_38064,N_38891);
xnor U40986 (N_40986,N_38413,N_38067);
xnor U40987 (N_40987,N_39534,N_38893);
and U40988 (N_40988,N_38634,N_39649);
xor U40989 (N_40989,N_39132,N_39066);
and U40990 (N_40990,N_38313,N_38947);
nor U40991 (N_40991,N_38999,N_39424);
or U40992 (N_40992,N_38384,N_38101);
and U40993 (N_40993,N_38643,N_38881);
xor U40994 (N_40994,N_39631,N_39194);
and U40995 (N_40995,N_38195,N_38428);
nand U40996 (N_40996,N_38115,N_39503);
and U40997 (N_40997,N_39675,N_38962);
or U40998 (N_40998,N_38791,N_39935);
and U40999 (N_40999,N_38810,N_38598);
and U41000 (N_41000,N_39863,N_39177);
nor U41001 (N_41001,N_38187,N_38357);
and U41002 (N_41002,N_39782,N_38087);
xnor U41003 (N_41003,N_39954,N_38376);
and U41004 (N_41004,N_39687,N_39713);
xnor U41005 (N_41005,N_38002,N_39750);
and U41006 (N_41006,N_38442,N_38690);
nor U41007 (N_41007,N_39735,N_39548);
or U41008 (N_41008,N_38073,N_38390);
and U41009 (N_41009,N_39847,N_39542);
nand U41010 (N_41010,N_38741,N_38103);
and U41011 (N_41011,N_38715,N_38398);
or U41012 (N_41012,N_39303,N_39342);
and U41013 (N_41013,N_38277,N_39257);
xnor U41014 (N_41014,N_38661,N_39430);
nor U41015 (N_41015,N_39595,N_38106);
and U41016 (N_41016,N_38916,N_38136);
nand U41017 (N_41017,N_38632,N_39747);
or U41018 (N_41018,N_38070,N_38674);
or U41019 (N_41019,N_38355,N_39296);
and U41020 (N_41020,N_38646,N_38479);
xor U41021 (N_41021,N_39116,N_39503);
and U41022 (N_41022,N_38178,N_38220);
or U41023 (N_41023,N_38728,N_39087);
or U41024 (N_41024,N_39987,N_39799);
nor U41025 (N_41025,N_38213,N_39710);
or U41026 (N_41026,N_38523,N_39269);
nor U41027 (N_41027,N_39718,N_39731);
xnor U41028 (N_41028,N_39918,N_38584);
xnor U41029 (N_41029,N_39021,N_39196);
nand U41030 (N_41030,N_39305,N_38751);
nor U41031 (N_41031,N_38354,N_39696);
and U41032 (N_41032,N_39344,N_38355);
xnor U41033 (N_41033,N_39441,N_38923);
nor U41034 (N_41034,N_39536,N_39618);
or U41035 (N_41035,N_39484,N_38459);
or U41036 (N_41036,N_39538,N_39759);
nand U41037 (N_41037,N_39666,N_39182);
nand U41038 (N_41038,N_38498,N_38589);
xnor U41039 (N_41039,N_38653,N_38941);
nand U41040 (N_41040,N_38528,N_38363);
or U41041 (N_41041,N_39822,N_39846);
and U41042 (N_41042,N_39814,N_38419);
or U41043 (N_41043,N_39147,N_39320);
or U41044 (N_41044,N_38453,N_39519);
and U41045 (N_41045,N_38641,N_39624);
xnor U41046 (N_41046,N_39687,N_38522);
or U41047 (N_41047,N_38151,N_39068);
and U41048 (N_41048,N_39761,N_38783);
xnor U41049 (N_41049,N_38528,N_39560);
nand U41050 (N_41050,N_39222,N_39679);
nor U41051 (N_41051,N_39722,N_39914);
and U41052 (N_41052,N_39602,N_38416);
xor U41053 (N_41053,N_39853,N_39872);
xnor U41054 (N_41054,N_39847,N_38875);
nor U41055 (N_41055,N_38092,N_38361);
or U41056 (N_41056,N_39471,N_39267);
nor U41057 (N_41057,N_38176,N_38562);
and U41058 (N_41058,N_38505,N_38149);
and U41059 (N_41059,N_38426,N_39255);
nand U41060 (N_41060,N_38518,N_39216);
xnor U41061 (N_41061,N_38325,N_39867);
and U41062 (N_41062,N_39549,N_38672);
nor U41063 (N_41063,N_38947,N_38850);
xor U41064 (N_41064,N_38006,N_38310);
and U41065 (N_41065,N_39067,N_38813);
or U41066 (N_41066,N_38148,N_39066);
and U41067 (N_41067,N_39322,N_39642);
nor U41068 (N_41068,N_39348,N_39584);
and U41069 (N_41069,N_39140,N_39202);
or U41070 (N_41070,N_39272,N_39584);
nor U41071 (N_41071,N_38561,N_38377);
or U41072 (N_41072,N_39702,N_38408);
or U41073 (N_41073,N_39537,N_38649);
and U41074 (N_41074,N_38581,N_39966);
xnor U41075 (N_41075,N_39667,N_39037);
nand U41076 (N_41076,N_38877,N_39470);
nand U41077 (N_41077,N_39509,N_38499);
xor U41078 (N_41078,N_39411,N_39176);
xor U41079 (N_41079,N_39663,N_39042);
xor U41080 (N_41080,N_39978,N_39247);
nor U41081 (N_41081,N_38128,N_39064);
and U41082 (N_41082,N_39741,N_39276);
xnor U41083 (N_41083,N_39337,N_38283);
or U41084 (N_41084,N_38249,N_38008);
nor U41085 (N_41085,N_39313,N_39927);
nand U41086 (N_41086,N_38798,N_38901);
nor U41087 (N_41087,N_39482,N_39287);
nand U41088 (N_41088,N_38474,N_38975);
or U41089 (N_41089,N_39522,N_38905);
xor U41090 (N_41090,N_39528,N_39359);
nand U41091 (N_41091,N_39678,N_38532);
nand U41092 (N_41092,N_38694,N_38132);
nor U41093 (N_41093,N_38299,N_38074);
nand U41094 (N_41094,N_39227,N_39148);
nor U41095 (N_41095,N_39200,N_39162);
xnor U41096 (N_41096,N_38830,N_38393);
or U41097 (N_41097,N_38448,N_39938);
or U41098 (N_41098,N_38001,N_38209);
nor U41099 (N_41099,N_38863,N_39038);
or U41100 (N_41100,N_38333,N_38011);
nand U41101 (N_41101,N_39665,N_39895);
and U41102 (N_41102,N_38618,N_38296);
nor U41103 (N_41103,N_38698,N_39425);
nand U41104 (N_41104,N_39586,N_39804);
nand U41105 (N_41105,N_39840,N_38373);
nand U41106 (N_41106,N_39924,N_38820);
xor U41107 (N_41107,N_38581,N_39070);
and U41108 (N_41108,N_39043,N_39494);
nor U41109 (N_41109,N_38402,N_39491);
and U41110 (N_41110,N_39127,N_39134);
and U41111 (N_41111,N_38601,N_38847);
nand U41112 (N_41112,N_39840,N_39904);
nor U41113 (N_41113,N_39970,N_38231);
and U41114 (N_41114,N_39709,N_39616);
nand U41115 (N_41115,N_38987,N_38972);
or U41116 (N_41116,N_39182,N_39062);
nor U41117 (N_41117,N_39300,N_39574);
nand U41118 (N_41118,N_38808,N_38572);
and U41119 (N_41119,N_38566,N_39027);
nor U41120 (N_41120,N_38881,N_38871);
xnor U41121 (N_41121,N_38890,N_38550);
and U41122 (N_41122,N_39942,N_38662);
xnor U41123 (N_41123,N_38187,N_38689);
nor U41124 (N_41124,N_38853,N_39367);
and U41125 (N_41125,N_38561,N_38345);
and U41126 (N_41126,N_39186,N_38352);
xor U41127 (N_41127,N_39029,N_39864);
nand U41128 (N_41128,N_39658,N_39422);
nand U41129 (N_41129,N_39070,N_38867);
xor U41130 (N_41130,N_39219,N_38408);
or U41131 (N_41131,N_38722,N_39046);
nand U41132 (N_41132,N_38366,N_38122);
nand U41133 (N_41133,N_39550,N_39291);
xor U41134 (N_41134,N_38573,N_38922);
and U41135 (N_41135,N_39739,N_39033);
nand U41136 (N_41136,N_38573,N_39627);
nand U41137 (N_41137,N_38777,N_39229);
nor U41138 (N_41138,N_38429,N_39362);
nand U41139 (N_41139,N_39013,N_38221);
nand U41140 (N_41140,N_38134,N_39636);
xnor U41141 (N_41141,N_38987,N_39881);
nand U41142 (N_41142,N_38955,N_39563);
nor U41143 (N_41143,N_39836,N_38725);
nand U41144 (N_41144,N_39298,N_39086);
and U41145 (N_41145,N_38693,N_38892);
nand U41146 (N_41146,N_39563,N_39442);
or U41147 (N_41147,N_39019,N_39251);
and U41148 (N_41148,N_39545,N_39847);
and U41149 (N_41149,N_39754,N_39753);
nor U41150 (N_41150,N_38501,N_38348);
or U41151 (N_41151,N_39139,N_39847);
or U41152 (N_41152,N_38283,N_38491);
nor U41153 (N_41153,N_39896,N_38095);
xnor U41154 (N_41154,N_38859,N_39390);
or U41155 (N_41155,N_38424,N_38410);
or U41156 (N_41156,N_38415,N_39284);
nor U41157 (N_41157,N_38881,N_38158);
or U41158 (N_41158,N_38437,N_39441);
nand U41159 (N_41159,N_39336,N_38648);
nand U41160 (N_41160,N_38857,N_38017);
xor U41161 (N_41161,N_38883,N_38033);
or U41162 (N_41162,N_38263,N_39176);
nand U41163 (N_41163,N_38701,N_38254);
or U41164 (N_41164,N_38033,N_38742);
nor U41165 (N_41165,N_39897,N_39334);
and U41166 (N_41166,N_38608,N_38515);
nor U41167 (N_41167,N_39570,N_38569);
xnor U41168 (N_41168,N_39396,N_39766);
nor U41169 (N_41169,N_38734,N_38797);
and U41170 (N_41170,N_38684,N_38385);
and U41171 (N_41171,N_38306,N_38662);
or U41172 (N_41172,N_39151,N_39326);
nor U41173 (N_41173,N_39158,N_38393);
nor U41174 (N_41174,N_39009,N_39895);
or U41175 (N_41175,N_39763,N_38005);
xor U41176 (N_41176,N_39338,N_39012);
and U41177 (N_41177,N_38422,N_39569);
xnor U41178 (N_41178,N_39351,N_39518);
nand U41179 (N_41179,N_39806,N_38375);
or U41180 (N_41180,N_38179,N_38341);
xor U41181 (N_41181,N_39317,N_39252);
nand U41182 (N_41182,N_38001,N_39735);
and U41183 (N_41183,N_38917,N_39032);
nor U41184 (N_41184,N_39261,N_39777);
xor U41185 (N_41185,N_39582,N_38621);
xor U41186 (N_41186,N_39461,N_38642);
nand U41187 (N_41187,N_39141,N_38540);
nor U41188 (N_41188,N_38017,N_39762);
xor U41189 (N_41189,N_38962,N_39780);
and U41190 (N_41190,N_38264,N_39982);
nor U41191 (N_41191,N_38008,N_39045);
or U41192 (N_41192,N_38030,N_38847);
nand U41193 (N_41193,N_38238,N_38222);
and U41194 (N_41194,N_39392,N_39779);
or U41195 (N_41195,N_39501,N_38251);
and U41196 (N_41196,N_38217,N_39925);
nor U41197 (N_41197,N_39329,N_38292);
nor U41198 (N_41198,N_39851,N_38381);
and U41199 (N_41199,N_39607,N_39506);
nand U41200 (N_41200,N_38788,N_38001);
or U41201 (N_41201,N_38411,N_39789);
or U41202 (N_41202,N_38894,N_38069);
and U41203 (N_41203,N_39945,N_39422);
nor U41204 (N_41204,N_39565,N_39764);
xor U41205 (N_41205,N_38475,N_38706);
nor U41206 (N_41206,N_39119,N_39111);
nor U41207 (N_41207,N_39835,N_39584);
and U41208 (N_41208,N_38748,N_38876);
or U41209 (N_41209,N_39404,N_39631);
or U41210 (N_41210,N_38793,N_39293);
nand U41211 (N_41211,N_38616,N_38634);
xnor U41212 (N_41212,N_39284,N_38322);
nor U41213 (N_41213,N_38802,N_38930);
nor U41214 (N_41214,N_38482,N_39151);
and U41215 (N_41215,N_38392,N_39915);
nand U41216 (N_41216,N_39501,N_39088);
xnor U41217 (N_41217,N_38516,N_38174);
or U41218 (N_41218,N_38412,N_39865);
xnor U41219 (N_41219,N_39881,N_38567);
xor U41220 (N_41220,N_38020,N_38220);
and U41221 (N_41221,N_39958,N_39213);
nor U41222 (N_41222,N_39167,N_38129);
or U41223 (N_41223,N_39653,N_39170);
or U41224 (N_41224,N_39214,N_39139);
or U41225 (N_41225,N_38626,N_38377);
nand U41226 (N_41226,N_38356,N_38918);
nor U41227 (N_41227,N_38895,N_39993);
nand U41228 (N_41228,N_38973,N_38623);
nor U41229 (N_41229,N_39519,N_38868);
or U41230 (N_41230,N_38500,N_39756);
nor U41231 (N_41231,N_39268,N_39506);
xnor U41232 (N_41232,N_39561,N_39978);
nand U41233 (N_41233,N_38626,N_38565);
nand U41234 (N_41234,N_38674,N_39104);
or U41235 (N_41235,N_39540,N_38457);
nor U41236 (N_41236,N_39586,N_39253);
xor U41237 (N_41237,N_39348,N_38098);
nor U41238 (N_41238,N_39731,N_38157);
or U41239 (N_41239,N_38116,N_39414);
nand U41240 (N_41240,N_39307,N_39543);
nor U41241 (N_41241,N_38328,N_39584);
nor U41242 (N_41242,N_39553,N_38963);
and U41243 (N_41243,N_39607,N_38841);
nand U41244 (N_41244,N_38504,N_38369);
nand U41245 (N_41245,N_39014,N_39043);
and U41246 (N_41246,N_38503,N_38963);
and U41247 (N_41247,N_38794,N_39018);
nand U41248 (N_41248,N_39041,N_38135);
and U41249 (N_41249,N_39263,N_39580);
nand U41250 (N_41250,N_39210,N_38488);
nand U41251 (N_41251,N_38181,N_38328);
and U41252 (N_41252,N_38127,N_39400);
and U41253 (N_41253,N_38491,N_38840);
and U41254 (N_41254,N_39981,N_38514);
and U41255 (N_41255,N_39239,N_38597);
and U41256 (N_41256,N_38494,N_38885);
and U41257 (N_41257,N_38003,N_38599);
xor U41258 (N_41258,N_39784,N_38631);
nand U41259 (N_41259,N_39244,N_38653);
or U41260 (N_41260,N_38899,N_38559);
and U41261 (N_41261,N_38055,N_38585);
nor U41262 (N_41262,N_39666,N_38102);
nor U41263 (N_41263,N_39728,N_39658);
or U41264 (N_41264,N_38153,N_39186);
or U41265 (N_41265,N_38792,N_39285);
nor U41266 (N_41266,N_39207,N_38063);
nor U41267 (N_41267,N_39922,N_38059);
or U41268 (N_41268,N_39027,N_38937);
and U41269 (N_41269,N_39611,N_39364);
nand U41270 (N_41270,N_38802,N_38359);
or U41271 (N_41271,N_38671,N_39684);
xnor U41272 (N_41272,N_39849,N_38297);
nor U41273 (N_41273,N_39059,N_39513);
or U41274 (N_41274,N_38304,N_39173);
and U41275 (N_41275,N_38655,N_39816);
xor U41276 (N_41276,N_38397,N_38519);
xnor U41277 (N_41277,N_38741,N_38822);
nand U41278 (N_41278,N_38288,N_39977);
and U41279 (N_41279,N_39958,N_38998);
nand U41280 (N_41280,N_39078,N_39275);
and U41281 (N_41281,N_38872,N_38561);
nand U41282 (N_41282,N_39180,N_38767);
or U41283 (N_41283,N_38269,N_38926);
and U41284 (N_41284,N_39685,N_38936);
nand U41285 (N_41285,N_38935,N_39344);
xor U41286 (N_41286,N_39560,N_39501);
nor U41287 (N_41287,N_39460,N_39536);
nand U41288 (N_41288,N_38549,N_39524);
and U41289 (N_41289,N_38517,N_39310);
or U41290 (N_41290,N_39738,N_39381);
xnor U41291 (N_41291,N_39341,N_38681);
nand U41292 (N_41292,N_39683,N_39413);
xor U41293 (N_41293,N_39513,N_38917);
or U41294 (N_41294,N_38468,N_39657);
nand U41295 (N_41295,N_39751,N_38773);
or U41296 (N_41296,N_39028,N_39552);
and U41297 (N_41297,N_39922,N_38563);
nand U41298 (N_41298,N_38974,N_39532);
or U41299 (N_41299,N_39480,N_39420);
xnor U41300 (N_41300,N_39267,N_39122);
nor U41301 (N_41301,N_39015,N_39056);
or U41302 (N_41302,N_39568,N_39330);
nor U41303 (N_41303,N_38963,N_38616);
xor U41304 (N_41304,N_39883,N_38545);
nand U41305 (N_41305,N_38982,N_39451);
and U41306 (N_41306,N_38427,N_39083);
and U41307 (N_41307,N_39558,N_39074);
xnor U41308 (N_41308,N_38697,N_39335);
nor U41309 (N_41309,N_38656,N_39076);
nand U41310 (N_41310,N_39699,N_39616);
xor U41311 (N_41311,N_39760,N_38186);
nand U41312 (N_41312,N_38928,N_39307);
xnor U41313 (N_41313,N_38659,N_39451);
and U41314 (N_41314,N_38256,N_38573);
xnor U41315 (N_41315,N_39020,N_38761);
xor U41316 (N_41316,N_38796,N_38620);
nor U41317 (N_41317,N_39579,N_38627);
xnor U41318 (N_41318,N_38692,N_39655);
or U41319 (N_41319,N_39627,N_38850);
or U41320 (N_41320,N_39740,N_39765);
or U41321 (N_41321,N_38424,N_39881);
and U41322 (N_41322,N_38749,N_39672);
nor U41323 (N_41323,N_39072,N_39504);
or U41324 (N_41324,N_39560,N_38590);
xnor U41325 (N_41325,N_38102,N_38464);
xnor U41326 (N_41326,N_39251,N_39198);
nand U41327 (N_41327,N_38587,N_39282);
and U41328 (N_41328,N_38817,N_38920);
or U41329 (N_41329,N_38166,N_39966);
or U41330 (N_41330,N_39326,N_39871);
and U41331 (N_41331,N_38923,N_38985);
and U41332 (N_41332,N_38912,N_39202);
or U41333 (N_41333,N_39407,N_39563);
xnor U41334 (N_41334,N_39977,N_38535);
or U41335 (N_41335,N_38632,N_38709);
or U41336 (N_41336,N_39512,N_38308);
nor U41337 (N_41337,N_38605,N_38063);
or U41338 (N_41338,N_38603,N_38157);
xnor U41339 (N_41339,N_39388,N_39043);
nand U41340 (N_41340,N_38062,N_38932);
and U41341 (N_41341,N_39491,N_39455);
or U41342 (N_41342,N_39723,N_38871);
nor U41343 (N_41343,N_39761,N_38109);
or U41344 (N_41344,N_38125,N_39012);
and U41345 (N_41345,N_38966,N_39409);
nand U41346 (N_41346,N_39089,N_38697);
nand U41347 (N_41347,N_38943,N_38806);
nand U41348 (N_41348,N_39002,N_39290);
nand U41349 (N_41349,N_39933,N_38354);
or U41350 (N_41350,N_39627,N_39458);
and U41351 (N_41351,N_38708,N_38956);
nor U41352 (N_41352,N_39450,N_38215);
and U41353 (N_41353,N_38818,N_38590);
or U41354 (N_41354,N_38395,N_39532);
and U41355 (N_41355,N_39037,N_38662);
and U41356 (N_41356,N_38087,N_38495);
nor U41357 (N_41357,N_39428,N_39029);
and U41358 (N_41358,N_39758,N_38737);
xnor U41359 (N_41359,N_39153,N_38019);
or U41360 (N_41360,N_38854,N_38470);
xnor U41361 (N_41361,N_39003,N_38402);
nand U41362 (N_41362,N_39806,N_38407);
or U41363 (N_41363,N_39855,N_38158);
xor U41364 (N_41364,N_38277,N_39798);
and U41365 (N_41365,N_38708,N_39120);
xor U41366 (N_41366,N_39884,N_38508);
nand U41367 (N_41367,N_38477,N_39155);
or U41368 (N_41368,N_39355,N_39400);
or U41369 (N_41369,N_38677,N_38682);
or U41370 (N_41370,N_39293,N_38636);
xnor U41371 (N_41371,N_38611,N_39552);
xnor U41372 (N_41372,N_38314,N_39342);
or U41373 (N_41373,N_38174,N_38225);
and U41374 (N_41374,N_39596,N_38965);
and U41375 (N_41375,N_39590,N_39109);
nor U41376 (N_41376,N_39626,N_39918);
or U41377 (N_41377,N_39895,N_38622);
nand U41378 (N_41378,N_39563,N_38219);
and U41379 (N_41379,N_39040,N_39078);
or U41380 (N_41380,N_39947,N_39941);
and U41381 (N_41381,N_39513,N_38486);
and U41382 (N_41382,N_38500,N_39748);
and U41383 (N_41383,N_39502,N_39496);
nor U41384 (N_41384,N_38142,N_39455);
or U41385 (N_41385,N_39941,N_38702);
or U41386 (N_41386,N_38177,N_39701);
nand U41387 (N_41387,N_39874,N_39416);
nor U41388 (N_41388,N_38701,N_39327);
and U41389 (N_41389,N_38465,N_39103);
nand U41390 (N_41390,N_38367,N_38909);
or U41391 (N_41391,N_38889,N_39701);
or U41392 (N_41392,N_38076,N_39197);
or U41393 (N_41393,N_38639,N_39312);
or U41394 (N_41394,N_39831,N_39870);
or U41395 (N_41395,N_38742,N_38147);
nor U41396 (N_41396,N_39746,N_39278);
nand U41397 (N_41397,N_38499,N_39704);
nand U41398 (N_41398,N_38396,N_39384);
nand U41399 (N_41399,N_39297,N_39804);
and U41400 (N_41400,N_39805,N_39003);
nand U41401 (N_41401,N_38705,N_39245);
xor U41402 (N_41402,N_38511,N_38471);
and U41403 (N_41403,N_38069,N_39130);
nand U41404 (N_41404,N_39753,N_38407);
or U41405 (N_41405,N_39946,N_39549);
xnor U41406 (N_41406,N_38537,N_39299);
nand U41407 (N_41407,N_38930,N_39030);
and U41408 (N_41408,N_38259,N_39532);
nand U41409 (N_41409,N_39478,N_39325);
xnor U41410 (N_41410,N_38243,N_38749);
nor U41411 (N_41411,N_39883,N_38304);
nand U41412 (N_41412,N_39375,N_38671);
or U41413 (N_41413,N_38879,N_39460);
nand U41414 (N_41414,N_39079,N_39366);
or U41415 (N_41415,N_38821,N_38742);
and U41416 (N_41416,N_39355,N_39633);
nand U41417 (N_41417,N_38527,N_38349);
xor U41418 (N_41418,N_38266,N_38309);
and U41419 (N_41419,N_39151,N_38073);
xor U41420 (N_41420,N_39961,N_39721);
or U41421 (N_41421,N_38883,N_39272);
or U41422 (N_41422,N_39104,N_39620);
xnor U41423 (N_41423,N_38089,N_38818);
nor U41424 (N_41424,N_38548,N_39622);
nor U41425 (N_41425,N_38948,N_38111);
nand U41426 (N_41426,N_39456,N_38208);
nor U41427 (N_41427,N_39745,N_38393);
nor U41428 (N_41428,N_39923,N_39683);
nor U41429 (N_41429,N_38607,N_38307);
or U41430 (N_41430,N_39177,N_38715);
or U41431 (N_41431,N_39475,N_38432);
or U41432 (N_41432,N_39533,N_39786);
and U41433 (N_41433,N_39998,N_38249);
or U41434 (N_41434,N_38211,N_39674);
and U41435 (N_41435,N_38695,N_39193);
xnor U41436 (N_41436,N_38363,N_39453);
nand U41437 (N_41437,N_39877,N_38360);
nand U41438 (N_41438,N_38739,N_38804);
and U41439 (N_41439,N_39605,N_39552);
nor U41440 (N_41440,N_39481,N_39723);
xnor U41441 (N_41441,N_39979,N_38950);
nor U41442 (N_41442,N_39393,N_39939);
or U41443 (N_41443,N_38641,N_39846);
and U41444 (N_41444,N_39499,N_38222);
nor U41445 (N_41445,N_38418,N_38765);
xor U41446 (N_41446,N_38682,N_39265);
xnor U41447 (N_41447,N_39446,N_39349);
xnor U41448 (N_41448,N_38521,N_38559);
or U41449 (N_41449,N_39781,N_38095);
nand U41450 (N_41450,N_39216,N_38942);
xor U41451 (N_41451,N_39000,N_39163);
and U41452 (N_41452,N_38596,N_39456);
nand U41453 (N_41453,N_38180,N_38237);
nor U41454 (N_41454,N_38864,N_39706);
xnor U41455 (N_41455,N_38199,N_39163);
and U41456 (N_41456,N_38173,N_38072);
xor U41457 (N_41457,N_38228,N_38067);
nor U41458 (N_41458,N_38719,N_38159);
nand U41459 (N_41459,N_38483,N_39374);
xnor U41460 (N_41460,N_38633,N_39707);
nor U41461 (N_41461,N_39748,N_38767);
nand U41462 (N_41462,N_38604,N_38060);
xnor U41463 (N_41463,N_38219,N_38179);
nand U41464 (N_41464,N_38832,N_38253);
xnor U41465 (N_41465,N_39095,N_39431);
nand U41466 (N_41466,N_38782,N_39011);
or U41467 (N_41467,N_39545,N_38259);
xnor U41468 (N_41468,N_39979,N_39727);
nor U41469 (N_41469,N_38271,N_38984);
nand U41470 (N_41470,N_38148,N_38084);
and U41471 (N_41471,N_38247,N_39274);
xor U41472 (N_41472,N_39672,N_39540);
nor U41473 (N_41473,N_38179,N_39000);
and U41474 (N_41474,N_38223,N_39108);
nor U41475 (N_41475,N_39082,N_39778);
or U41476 (N_41476,N_39161,N_39726);
and U41477 (N_41477,N_38716,N_38324);
nand U41478 (N_41478,N_38290,N_38748);
xnor U41479 (N_41479,N_39804,N_39584);
xnor U41480 (N_41480,N_39416,N_38196);
and U41481 (N_41481,N_38343,N_38045);
nand U41482 (N_41482,N_39991,N_38491);
nor U41483 (N_41483,N_38046,N_38617);
nor U41484 (N_41484,N_39524,N_38667);
and U41485 (N_41485,N_39527,N_39847);
or U41486 (N_41486,N_39179,N_38196);
or U41487 (N_41487,N_38677,N_38507);
and U41488 (N_41488,N_38829,N_39141);
and U41489 (N_41489,N_38927,N_39016);
or U41490 (N_41490,N_39526,N_39802);
nor U41491 (N_41491,N_38608,N_38883);
nand U41492 (N_41492,N_39536,N_39970);
or U41493 (N_41493,N_39997,N_39219);
nor U41494 (N_41494,N_38666,N_38673);
and U41495 (N_41495,N_38659,N_39622);
or U41496 (N_41496,N_39360,N_38613);
nand U41497 (N_41497,N_38089,N_39520);
xnor U41498 (N_41498,N_39475,N_39524);
nor U41499 (N_41499,N_39409,N_39498);
or U41500 (N_41500,N_39181,N_39271);
nor U41501 (N_41501,N_38473,N_38008);
and U41502 (N_41502,N_39913,N_38602);
nor U41503 (N_41503,N_39671,N_39326);
nand U41504 (N_41504,N_39241,N_38572);
xnor U41505 (N_41505,N_38124,N_38829);
and U41506 (N_41506,N_39019,N_38010);
or U41507 (N_41507,N_39965,N_39828);
and U41508 (N_41508,N_39032,N_38531);
xnor U41509 (N_41509,N_39320,N_38021);
or U41510 (N_41510,N_39304,N_39047);
and U41511 (N_41511,N_39951,N_39345);
nor U41512 (N_41512,N_38283,N_39334);
or U41513 (N_41513,N_39277,N_39785);
nand U41514 (N_41514,N_38897,N_39551);
nand U41515 (N_41515,N_39784,N_38129);
nor U41516 (N_41516,N_38952,N_39593);
nor U41517 (N_41517,N_39031,N_39931);
or U41518 (N_41518,N_38614,N_38193);
nand U41519 (N_41519,N_39005,N_39717);
or U41520 (N_41520,N_38651,N_38788);
or U41521 (N_41521,N_38493,N_38041);
nand U41522 (N_41522,N_38920,N_39446);
nand U41523 (N_41523,N_38566,N_38027);
and U41524 (N_41524,N_38744,N_39449);
xor U41525 (N_41525,N_38016,N_38973);
and U41526 (N_41526,N_38652,N_38989);
or U41527 (N_41527,N_39094,N_38316);
nand U41528 (N_41528,N_39459,N_38243);
xnor U41529 (N_41529,N_38110,N_39026);
nor U41530 (N_41530,N_38745,N_38633);
nor U41531 (N_41531,N_39638,N_38741);
and U41532 (N_41532,N_38651,N_39810);
or U41533 (N_41533,N_39930,N_39589);
nand U41534 (N_41534,N_38520,N_39002);
or U41535 (N_41535,N_39712,N_39366);
or U41536 (N_41536,N_39851,N_39151);
nor U41537 (N_41537,N_39370,N_38583);
xor U41538 (N_41538,N_38522,N_39842);
xnor U41539 (N_41539,N_38514,N_38603);
or U41540 (N_41540,N_39015,N_38804);
nor U41541 (N_41541,N_39671,N_39436);
nand U41542 (N_41542,N_39051,N_38641);
nand U41543 (N_41543,N_39700,N_38170);
and U41544 (N_41544,N_38300,N_39066);
nor U41545 (N_41545,N_38682,N_38987);
nand U41546 (N_41546,N_38320,N_38060);
nand U41547 (N_41547,N_39564,N_38478);
nor U41548 (N_41548,N_39175,N_38290);
nand U41549 (N_41549,N_38220,N_38442);
xor U41550 (N_41550,N_39303,N_38900);
nand U41551 (N_41551,N_38682,N_39433);
xor U41552 (N_41552,N_39366,N_39078);
nand U41553 (N_41553,N_39663,N_38937);
or U41554 (N_41554,N_38612,N_39571);
and U41555 (N_41555,N_38591,N_39828);
xor U41556 (N_41556,N_38090,N_38885);
nor U41557 (N_41557,N_38176,N_38553);
or U41558 (N_41558,N_39896,N_38448);
nand U41559 (N_41559,N_38750,N_38314);
nor U41560 (N_41560,N_39698,N_38080);
nand U41561 (N_41561,N_39846,N_39015);
or U41562 (N_41562,N_38153,N_39736);
nand U41563 (N_41563,N_38821,N_39433);
xnor U41564 (N_41564,N_39698,N_38304);
or U41565 (N_41565,N_38062,N_38180);
xnor U41566 (N_41566,N_38887,N_38683);
nor U41567 (N_41567,N_39916,N_38410);
and U41568 (N_41568,N_38856,N_39001);
nor U41569 (N_41569,N_38321,N_39757);
nand U41570 (N_41570,N_39542,N_38589);
or U41571 (N_41571,N_39220,N_38514);
or U41572 (N_41572,N_38067,N_39305);
or U41573 (N_41573,N_38716,N_38868);
xor U41574 (N_41574,N_39991,N_38984);
and U41575 (N_41575,N_39520,N_39996);
or U41576 (N_41576,N_39724,N_38411);
nor U41577 (N_41577,N_38639,N_39777);
nand U41578 (N_41578,N_39999,N_38724);
and U41579 (N_41579,N_39917,N_39985);
and U41580 (N_41580,N_39351,N_38140);
and U41581 (N_41581,N_38149,N_38371);
nor U41582 (N_41582,N_38417,N_39469);
and U41583 (N_41583,N_38398,N_38095);
or U41584 (N_41584,N_38491,N_38978);
or U41585 (N_41585,N_39396,N_39095);
xor U41586 (N_41586,N_39097,N_38468);
or U41587 (N_41587,N_38555,N_38782);
or U41588 (N_41588,N_38997,N_39837);
or U41589 (N_41589,N_39457,N_38022);
xor U41590 (N_41590,N_39216,N_38143);
or U41591 (N_41591,N_38003,N_38605);
nand U41592 (N_41592,N_39020,N_38015);
and U41593 (N_41593,N_39558,N_39646);
and U41594 (N_41594,N_39591,N_39036);
nand U41595 (N_41595,N_39393,N_38180);
nand U41596 (N_41596,N_39231,N_39268);
and U41597 (N_41597,N_38745,N_38838);
or U41598 (N_41598,N_39219,N_38017);
or U41599 (N_41599,N_38976,N_38226);
or U41600 (N_41600,N_38850,N_39360);
xnor U41601 (N_41601,N_38217,N_38321);
nand U41602 (N_41602,N_38714,N_39257);
or U41603 (N_41603,N_38013,N_39829);
xnor U41604 (N_41604,N_38839,N_39502);
xor U41605 (N_41605,N_38363,N_38798);
nor U41606 (N_41606,N_38324,N_38339);
nor U41607 (N_41607,N_39535,N_38265);
xnor U41608 (N_41608,N_38067,N_39604);
or U41609 (N_41609,N_38612,N_38645);
nor U41610 (N_41610,N_38327,N_39359);
or U41611 (N_41611,N_39747,N_38105);
or U41612 (N_41612,N_39904,N_39226);
nor U41613 (N_41613,N_39385,N_38111);
nor U41614 (N_41614,N_39944,N_38081);
nand U41615 (N_41615,N_39657,N_39939);
nor U41616 (N_41616,N_38459,N_38817);
and U41617 (N_41617,N_38687,N_38521);
and U41618 (N_41618,N_38685,N_39544);
xnor U41619 (N_41619,N_38696,N_39735);
or U41620 (N_41620,N_38863,N_39895);
nand U41621 (N_41621,N_39373,N_39588);
nor U41622 (N_41622,N_38972,N_38686);
and U41623 (N_41623,N_39820,N_38861);
or U41624 (N_41624,N_39647,N_38099);
xnor U41625 (N_41625,N_38507,N_38131);
or U41626 (N_41626,N_39657,N_39767);
nand U41627 (N_41627,N_38959,N_39491);
or U41628 (N_41628,N_39967,N_39121);
xor U41629 (N_41629,N_39721,N_39464);
and U41630 (N_41630,N_39356,N_38104);
xor U41631 (N_41631,N_38895,N_39316);
xnor U41632 (N_41632,N_39810,N_38275);
xnor U41633 (N_41633,N_38709,N_38457);
xor U41634 (N_41634,N_38997,N_39638);
and U41635 (N_41635,N_38251,N_38780);
or U41636 (N_41636,N_39093,N_38357);
or U41637 (N_41637,N_39192,N_38359);
and U41638 (N_41638,N_39705,N_39831);
nor U41639 (N_41639,N_38399,N_39782);
nand U41640 (N_41640,N_39763,N_38816);
nand U41641 (N_41641,N_38771,N_39262);
or U41642 (N_41642,N_39804,N_38836);
or U41643 (N_41643,N_39757,N_39237);
nor U41644 (N_41644,N_39518,N_39106);
nand U41645 (N_41645,N_38066,N_38716);
or U41646 (N_41646,N_39159,N_38267);
nand U41647 (N_41647,N_38603,N_38812);
xor U41648 (N_41648,N_39994,N_39067);
nand U41649 (N_41649,N_39274,N_39249);
or U41650 (N_41650,N_38543,N_39780);
nor U41651 (N_41651,N_38375,N_39240);
nor U41652 (N_41652,N_38956,N_38044);
xnor U41653 (N_41653,N_38518,N_39369);
nor U41654 (N_41654,N_39151,N_39850);
and U41655 (N_41655,N_39901,N_39454);
or U41656 (N_41656,N_38252,N_39484);
or U41657 (N_41657,N_38314,N_39100);
nor U41658 (N_41658,N_38266,N_39546);
nand U41659 (N_41659,N_39400,N_38958);
nand U41660 (N_41660,N_38226,N_38884);
xor U41661 (N_41661,N_38198,N_39535);
nor U41662 (N_41662,N_39246,N_39434);
nand U41663 (N_41663,N_38571,N_38811);
and U41664 (N_41664,N_39447,N_38162);
and U41665 (N_41665,N_39200,N_38262);
and U41666 (N_41666,N_38238,N_39664);
or U41667 (N_41667,N_38471,N_39320);
or U41668 (N_41668,N_38789,N_38160);
and U41669 (N_41669,N_39522,N_39974);
or U41670 (N_41670,N_39579,N_39370);
nand U41671 (N_41671,N_39545,N_39242);
nor U41672 (N_41672,N_38896,N_38235);
nand U41673 (N_41673,N_39002,N_39123);
nand U41674 (N_41674,N_38035,N_39315);
or U41675 (N_41675,N_39819,N_39520);
xnor U41676 (N_41676,N_39777,N_39642);
or U41677 (N_41677,N_39758,N_39715);
nor U41678 (N_41678,N_39647,N_38174);
nand U41679 (N_41679,N_39395,N_39389);
or U41680 (N_41680,N_39953,N_38107);
nor U41681 (N_41681,N_38838,N_39432);
xnor U41682 (N_41682,N_39243,N_39235);
nand U41683 (N_41683,N_38641,N_39374);
nand U41684 (N_41684,N_38820,N_39148);
xnor U41685 (N_41685,N_38769,N_39321);
or U41686 (N_41686,N_38750,N_39896);
nand U41687 (N_41687,N_38938,N_39059);
nor U41688 (N_41688,N_39525,N_39469);
nor U41689 (N_41689,N_38837,N_38333);
and U41690 (N_41690,N_39184,N_39472);
xnor U41691 (N_41691,N_38115,N_39322);
nor U41692 (N_41692,N_38911,N_39947);
and U41693 (N_41693,N_39084,N_38467);
and U41694 (N_41694,N_39066,N_39418);
nand U41695 (N_41695,N_39720,N_39091);
or U41696 (N_41696,N_38085,N_39516);
nor U41697 (N_41697,N_38703,N_39946);
or U41698 (N_41698,N_38186,N_38162);
nor U41699 (N_41699,N_39188,N_38035);
xnor U41700 (N_41700,N_39525,N_39614);
or U41701 (N_41701,N_38485,N_39075);
nor U41702 (N_41702,N_38383,N_38245);
and U41703 (N_41703,N_39716,N_39807);
and U41704 (N_41704,N_38981,N_39320);
nand U41705 (N_41705,N_39622,N_39300);
or U41706 (N_41706,N_39389,N_38852);
and U41707 (N_41707,N_38517,N_38822);
or U41708 (N_41708,N_39586,N_38007);
and U41709 (N_41709,N_39976,N_39106);
nand U41710 (N_41710,N_39814,N_39483);
xor U41711 (N_41711,N_39276,N_39933);
nor U41712 (N_41712,N_39976,N_38277);
nand U41713 (N_41713,N_38043,N_39323);
and U41714 (N_41714,N_38317,N_39337);
xnor U41715 (N_41715,N_39770,N_38657);
xnor U41716 (N_41716,N_39637,N_39689);
or U41717 (N_41717,N_38762,N_38293);
and U41718 (N_41718,N_38069,N_38919);
and U41719 (N_41719,N_38477,N_38988);
and U41720 (N_41720,N_39899,N_38298);
and U41721 (N_41721,N_39772,N_38868);
and U41722 (N_41722,N_39318,N_39809);
nor U41723 (N_41723,N_39894,N_38234);
nand U41724 (N_41724,N_38883,N_39866);
nor U41725 (N_41725,N_39032,N_39396);
or U41726 (N_41726,N_38902,N_38528);
xnor U41727 (N_41727,N_39484,N_38477);
nor U41728 (N_41728,N_39065,N_38848);
or U41729 (N_41729,N_39453,N_38752);
nor U41730 (N_41730,N_39571,N_39447);
xnor U41731 (N_41731,N_38579,N_39606);
and U41732 (N_41732,N_39985,N_39184);
and U41733 (N_41733,N_38512,N_39679);
or U41734 (N_41734,N_38862,N_39749);
and U41735 (N_41735,N_38237,N_39701);
nand U41736 (N_41736,N_38503,N_39757);
or U41737 (N_41737,N_39706,N_39517);
and U41738 (N_41738,N_39768,N_39346);
or U41739 (N_41739,N_39636,N_39942);
nand U41740 (N_41740,N_38956,N_39841);
xnor U41741 (N_41741,N_38430,N_38666);
and U41742 (N_41742,N_39215,N_39972);
xnor U41743 (N_41743,N_38424,N_39412);
xor U41744 (N_41744,N_39626,N_38257);
or U41745 (N_41745,N_39024,N_39022);
and U41746 (N_41746,N_38767,N_38324);
nand U41747 (N_41747,N_38173,N_39594);
xor U41748 (N_41748,N_39178,N_38094);
nor U41749 (N_41749,N_38057,N_39508);
xor U41750 (N_41750,N_38099,N_39480);
nor U41751 (N_41751,N_39766,N_39325);
nor U41752 (N_41752,N_38165,N_39453);
and U41753 (N_41753,N_38793,N_38014);
xor U41754 (N_41754,N_38589,N_38525);
nor U41755 (N_41755,N_39188,N_38224);
nand U41756 (N_41756,N_39622,N_38665);
or U41757 (N_41757,N_38264,N_38629);
and U41758 (N_41758,N_39413,N_38529);
or U41759 (N_41759,N_39250,N_38397);
and U41760 (N_41760,N_38811,N_39389);
or U41761 (N_41761,N_38437,N_38137);
or U41762 (N_41762,N_39175,N_38962);
xor U41763 (N_41763,N_38990,N_38032);
and U41764 (N_41764,N_38163,N_38436);
nor U41765 (N_41765,N_39947,N_38043);
nor U41766 (N_41766,N_39790,N_38025);
and U41767 (N_41767,N_38436,N_39386);
or U41768 (N_41768,N_38869,N_38794);
nand U41769 (N_41769,N_38429,N_38577);
xor U41770 (N_41770,N_39399,N_39138);
xnor U41771 (N_41771,N_38894,N_39392);
nor U41772 (N_41772,N_38119,N_39711);
xor U41773 (N_41773,N_39199,N_39873);
xor U41774 (N_41774,N_38670,N_38532);
xnor U41775 (N_41775,N_38308,N_38253);
xnor U41776 (N_41776,N_39178,N_39719);
nor U41777 (N_41777,N_39210,N_38713);
or U41778 (N_41778,N_38136,N_39713);
and U41779 (N_41779,N_39756,N_38498);
nor U41780 (N_41780,N_39577,N_38009);
nand U41781 (N_41781,N_38230,N_39864);
or U41782 (N_41782,N_39811,N_38127);
or U41783 (N_41783,N_38668,N_39917);
nor U41784 (N_41784,N_38287,N_38742);
or U41785 (N_41785,N_38187,N_39909);
and U41786 (N_41786,N_39315,N_38463);
nand U41787 (N_41787,N_39582,N_39559);
and U41788 (N_41788,N_39248,N_38798);
xnor U41789 (N_41789,N_38540,N_38748);
nand U41790 (N_41790,N_39845,N_39366);
and U41791 (N_41791,N_38285,N_38544);
or U41792 (N_41792,N_39262,N_38173);
nand U41793 (N_41793,N_39657,N_39571);
nand U41794 (N_41794,N_38018,N_39402);
nand U41795 (N_41795,N_38476,N_39443);
xnor U41796 (N_41796,N_38272,N_39287);
nand U41797 (N_41797,N_39899,N_39100);
or U41798 (N_41798,N_39727,N_39420);
and U41799 (N_41799,N_39524,N_39283);
nor U41800 (N_41800,N_38982,N_39015);
and U41801 (N_41801,N_39738,N_38817);
nand U41802 (N_41802,N_39852,N_38583);
nor U41803 (N_41803,N_39671,N_38057);
and U41804 (N_41804,N_38850,N_38910);
xnor U41805 (N_41805,N_38293,N_38398);
or U41806 (N_41806,N_39543,N_39052);
nor U41807 (N_41807,N_39039,N_39581);
and U41808 (N_41808,N_39991,N_38917);
and U41809 (N_41809,N_38188,N_38054);
nand U41810 (N_41810,N_38764,N_38954);
nor U41811 (N_41811,N_39956,N_39784);
nor U41812 (N_41812,N_39274,N_39245);
xor U41813 (N_41813,N_39411,N_39638);
nor U41814 (N_41814,N_38335,N_38595);
nand U41815 (N_41815,N_38913,N_38311);
xnor U41816 (N_41816,N_39492,N_38365);
nor U41817 (N_41817,N_38348,N_39886);
xor U41818 (N_41818,N_39635,N_39166);
xor U41819 (N_41819,N_38248,N_38937);
or U41820 (N_41820,N_39395,N_38801);
xor U41821 (N_41821,N_38249,N_39869);
nand U41822 (N_41822,N_39404,N_38478);
or U41823 (N_41823,N_39633,N_39613);
xor U41824 (N_41824,N_39353,N_38819);
and U41825 (N_41825,N_38605,N_38178);
and U41826 (N_41826,N_38119,N_39507);
xor U41827 (N_41827,N_39753,N_38349);
nor U41828 (N_41828,N_39030,N_39080);
nand U41829 (N_41829,N_39364,N_38555);
or U41830 (N_41830,N_38699,N_38183);
nor U41831 (N_41831,N_39460,N_39264);
or U41832 (N_41832,N_38258,N_38820);
or U41833 (N_41833,N_39060,N_38770);
nand U41834 (N_41834,N_38352,N_38119);
nor U41835 (N_41835,N_39325,N_38627);
nor U41836 (N_41836,N_39773,N_38759);
or U41837 (N_41837,N_39026,N_38365);
nand U41838 (N_41838,N_39685,N_38442);
nor U41839 (N_41839,N_39777,N_38856);
and U41840 (N_41840,N_39329,N_38957);
and U41841 (N_41841,N_39072,N_39084);
nor U41842 (N_41842,N_38795,N_38804);
nand U41843 (N_41843,N_39829,N_39318);
nor U41844 (N_41844,N_38631,N_38877);
and U41845 (N_41845,N_39675,N_38875);
nor U41846 (N_41846,N_38832,N_39334);
or U41847 (N_41847,N_39345,N_38185);
nand U41848 (N_41848,N_38889,N_38912);
xor U41849 (N_41849,N_39225,N_38085);
nor U41850 (N_41850,N_38229,N_38160);
xor U41851 (N_41851,N_39002,N_39908);
and U41852 (N_41852,N_38519,N_39806);
nand U41853 (N_41853,N_39118,N_39753);
nor U41854 (N_41854,N_38867,N_38691);
and U41855 (N_41855,N_38811,N_38874);
and U41856 (N_41856,N_39176,N_39550);
or U41857 (N_41857,N_39798,N_38683);
or U41858 (N_41858,N_38260,N_38166);
nor U41859 (N_41859,N_39601,N_38159);
nand U41860 (N_41860,N_38991,N_38509);
xnor U41861 (N_41861,N_39741,N_39610);
nand U41862 (N_41862,N_39349,N_39707);
xor U41863 (N_41863,N_38624,N_39817);
and U41864 (N_41864,N_38004,N_39535);
and U41865 (N_41865,N_38287,N_39450);
xnor U41866 (N_41866,N_38722,N_38487);
nor U41867 (N_41867,N_38199,N_38090);
nor U41868 (N_41868,N_38723,N_39647);
or U41869 (N_41869,N_38420,N_38241);
xor U41870 (N_41870,N_39711,N_38855);
xnor U41871 (N_41871,N_39013,N_38505);
and U41872 (N_41872,N_38732,N_39571);
and U41873 (N_41873,N_38434,N_39428);
nand U41874 (N_41874,N_38325,N_38776);
xnor U41875 (N_41875,N_39349,N_39862);
and U41876 (N_41876,N_38640,N_38781);
or U41877 (N_41877,N_39343,N_38327);
xnor U41878 (N_41878,N_38420,N_38702);
nand U41879 (N_41879,N_39717,N_38959);
and U41880 (N_41880,N_39608,N_38284);
xnor U41881 (N_41881,N_39322,N_39885);
xor U41882 (N_41882,N_39827,N_38030);
nand U41883 (N_41883,N_39547,N_39383);
and U41884 (N_41884,N_38327,N_39669);
xnor U41885 (N_41885,N_38134,N_39872);
nor U41886 (N_41886,N_39220,N_38634);
or U41887 (N_41887,N_39461,N_39291);
xnor U41888 (N_41888,N_39177,N_39182);
and U41889 (N_41889,N_39101,N_38484);
xor U41890 (N_41890,N_39400,N_38196);
and U41891 (N_41891,N_39339,N_38621);
nor U41892 (N_41892,N_39098,N_39934);
or U41893 (N_41893,N_38379,N_39854);
xnor U41894 (N_41894,N_38264,N_39383);
xnor U41895 (N_41895,N_39919,N_38290);
nand U41896 (N_41896,N_38017,N_38038);
nor U41897 (N_41897,N_38512,N_38515);
nor U41898 (N_41898,N_38634,N_39672);
xnor U41899 (N_41899,N_39001,N_38293);
nor U41900 (N_41900,N_38543,N_39814);
and U41901 (N_41901,N_38078,N_38030);
nor U41902 (N_41902,N_39677,N_39792);
nand U41903 (N_41903,N_38335,N_39878);
or U41904 (N_41904,N_38997,N_38402);
or U41905 (N_41905,N_38572,N_39602);
and U41906 (N_41906,N_39562,N_39172);
nor U41907 (N_41907,N_39651,N_39776);
and U41908 (N_41908,N_38207,N_39856);
nand U41909 (N_41909,N_39249,N_38604);
xor U41910 (N_41910,N_38103,N_38211);
nand U41911 (N_41911,N_38986,N_38186);
nand U41912 (N_41912,N_39446,N_39026);
nand U41913 (N_41913,N_38554,N_38543);
nand U41914 (N_41914,N_38062,N_39194);
and U41915 (N_41915,N_39843,N_38657);
and U41916 (N_41916,N_38245,N_38277);
nand U41917 (N_41917,N_39830,N_38240);
and U41918 (N_41918,N_39713,N_38679);
or U41919 (N_41919,N_39681,N_38885);
nand U41920 (N_41920,N_39328,N_38726);
and U41921 (N_41921,N_38605,N_38966);
nor U41922 (N_41922,N_39526,N_38483);
or U41923 (N_41923,N_39242,N_38423);
and U41924 (N_41924,N_38500,N_39236);
or U41925 (N_41925,N_39411,N_39501);
or U41926 (N_41926,N_39738,N_39891);
xnor U41927 (N_41927,N_39965,N_39132);
nor U41928 (N_41928,N_38915,N_38255);
and U41929 (N_41929,N_39455,N_38762);
and U41930 (N_41930,N_39121,N_39354);
nand U41931 (N_41931,N_39296,N_39530);
xnor U41932 (N_41932,N_39309,N_38327);
nand U41933 (N_41933,N_39951,N_39178);
and U41934 (N_41934,N_39340,N_39565);
xor U41935 (N_41935,N_38634,N_38747);
xor U41936 (N_41936,N_38009,N_38947);
or U41937 (N_41937,N_39102,N_39932);
nand U41938 (N_41938,N_38811,N_38307);
and U41939 (N_41939,N_38555,N_38063);
nor U41940 (N_41940,N_38069,N_38649);
xor U41941 (N_41941,N_38277,N_39813);
nand U41942 (N_41942,N_39372,N_38513);
or U41943 (N_41943,N_39265,N_39912);
and U41944 (N_41944,N_39809,N_38026);
or U41945 (N_41945,N_39849,N_38783);
and U41946 (N_41946,N_38628,N_39561);
or U41947 (N_41947,N_39635,N_38384);
nand U41948 (N_41948,N_38667,N_39681);
nor U41949 (N_41949,N_39196,N_38666);
and U41950 (N_41950,N_39425,N_39253);
and U41951 (N_41951,N_39691,N_39281);
xnor U41952 (N_41952,N_39425,N_38511);
xnor U41953 (N_41953,N_39481,N_38725);
nor U41954 (N_41954,N_39040,N_38859);
nand U41955 (N_41955,N_39653,N_38350);
and U41956 (N_41956,N_39552,N_39161);
nand U41957 (N_41957,N_39414,N_39915);
or U41958 (N_41958,N_39908,N_39986);
xnor U41959 (N_41959,N_39428,N_39337);
nand U41960 (N_41960,N_39038,N_39152);
nand U41961 (N_41961,N_38733,N_39469);
or U41962 (N_41962,N_39003,N_38907);
xnor U41963 (N_41963,N_39164,N_38946);
and U41964 (N_41964,N_38786,N_39778);
xnor U41965 (N_41965,N_38244,N_39005);
nor U41966 (N_41966,N_38172,N_38286);
nand U41967 (N_41967,N_39682,N_38857);
and U41968 (N_41968,N_39892,N_39536);
xor U41969 (N_41969,N_38523,N_39152);
and U41970 (N_41970,N_38711,N_39752);
and U41971 (N_41971,N_38052,N_38444);
or U41972 (N_41972,N_38555,N_39238);
xor U41973 (N_41973,N_38340,N_39316);
nand U41974 (N_41974,N_39802,N_39390);
and U41975 (N_41975,N_38164,N_38668);
nor U41976 (N_41976,N_38531,N_38951);
nand U41977 (N_41977,N_39175,N_38566);
nor U41978 (N_41978,N_39532,N_39459);
xnor U41979 (N_41979,N_39539,N_39806);
and U41980 (N_41980,N_38350,N_38379);
nor U41981 (N_41981,N_39812,N_39662);
or U41982 (N_41982,N_38430,N_39345);
nand U41983 (N_41983,N_39436,N_38675);
xor U41984 (N_41984,N_39241,N_39057);
xnor U41985 (N_41985,N_38255,N_38618);
and U41986 (N_41986,N_38513,N_38148);
or U41987 (N_41987,N_39337,N_39038);
xor U41988 (N_41988,N_39516,N_38688);
nor U41989 (N_41989,N_39435,N_38004);
nand U41990 (N_41990,N_39798,N_39979);
xor U41991 (N_41991,N_39182,N_38298);
nand U41992 (N_41992,N_38057,N_38664);
nor U41993 (N_41993,N_38876,N_38774);
and U41994 (N_41994,N_38653,N_39765);
and U41995 (N_41995,N_39039,N_38920);
nand U41996 (N_41996,N_38042,N_38276);
and U41997 (N_41997,N_39782,N_39331);
nor U41998 (N_41998,N_38352,N_39252);
xor U41999 (N_41999,N_38876,N_38070);
or U42000 (N_42000,N_41458,N_40692);
and U42001 (N_42001,N_40660,N_41206);
nor U42002 (N_42002,N_40297,N_40547);
and U42003 (N_42003,N_40197,N_40840);
or U42004 (N_42004,N_40039,N_41593);
nand U42005 (N_42005,N_41711,N_41202);
and U42006 (N_42006,N_41392,N_41186);
xnor U42007 (N_42007,N_40009,N_41180);
nor U42008 (N_42008,N_40119,N_40595);
xnor U42009 (N_42009,N_41484,N_40135);
xor U42010 (N_42010,N_41495,N_41883);
xnor U42011 (N_42011,N_40513,N_40596);
or U42012 (N_42012,N_41130,N_40811);
xnor U42013 (N_42013,N_40054,N_41742);
or U42014 (N_42014,N_40201,N_41140);
xnor U42015 (N_42015,N_40299,N_40402);
xor U42016 (N_42016,N_41995,N_41896);
or U42017 (N_42017,N_41113,N_41248);
and U42018 (N_42018,N_41803,N_40233);
or U42019 (N_42019,N_40875,N_40609);
or U42020 (N_42020,N_40000,N_40731);
and U42021 (N_42021,N_41900,N_40842);
nand U42022 (N_42022,N_41482,N_40262);
or U42023 (N_42023,N_41270,N_41025);
xnor U42024 (N_42024,N_40223,N_41088);
nor U42025 (N_42025,N_40824,N_41759);
xor U42026 (N_42026,N_40294,N_41481);
nor U42027 (N_42027,N_40599,N_40554);
and U42028 (N_42028,N_41571,N_41216);
and U42029 (N_42029,N_40548,N_41899);
or U42030 (N_42030,N_40458,N_40486);
and U42031 (N_42031,N_40828,N_40801);
nand U42032 (N_42032,N_41697,N_41542);
and U42033 (N_42033,N_41148,N_40056);
nand U42034 (N_42034,N_41501,N_40709);
or U42035 (N_42035,N_40982,N_40154);
xor U42036 (N_42036,N_40524,N_41859);
or U42037 (N_42037,N_40913,N_41311);
and U42038 (N_42038,N_40863,N_41400);
xnor U42039 (N_42039,N_40807,N_40330);
xor U42040 (N_42040,N_40366,N_40045);
nor U42041 (N_42041,N_41766,N_41987);
xnor U42042 (N_42042,N_40158,N_40254);
xor U42043 (N_42043,N_40416,N_40950);
and U42044 (N_42044,N_41366,N_40217);
xnor U42045 (N_42045,N_41351,N_41373);
nand U42046 (N_42046,N_41097,N_41503);
nand U42047 (N_42047,N_40138,N_40246);
or U42048 (N_42048,N_40674,N_41273);
and U42049 (N_42049,N_41625,N_41595);
and U42050 (N_42050,N_40350,N_41645);
nand U42051 (N_42051,N_40694,N_40080);
nor U42052 (N_42052,N_40258,N_41961);
or U42053 (N_42053,N_40188,N_40150);
xnor U42054 (N_42054,N_40210,N_40467);
nand U42055 (N_42055,N_41889,N_41999);
nor U42056 (N_42056,N_41958,N_40805);
xnor U42057 (N_42057,N_40374,N_40221);
and U42058 (N_42058,N_41205,N_41124);
xnor U42059 (N_42059,N_41081,N_41380);
or U42060 (N_42060,N_40745,N_41396);
nand U42061 (N_42061,N_40979,N_40860);
or U42062 (N_42062,N_41211,N_41388);
nand U42063 (N_42063,N_41015,N_40604);
or U42064 (N_42064,N_40772,N_41941);
xnor U42065 (N_42065,N_41342,N_40174);
or U42066 (N_42066,N_41150,N_41310);
xnor U42067 (N_42067,N_40172,N_41829);
xor U42068 (N_42068,N_41801,N_40491);
xnor U42069 (N_42069,N_41655,N_41257);
xnor U42070 (N_42070,N_40556,N_41779);
nor U42071 (N_42071,N_41071,N_41127);
xor U42072 (N_42072,N_41973,N_40632);
nor U42073 (N_42073,N_41689,N_41720);
xor U42074 (N_42074,N_41797,N_40643);
nor U42075 (N_42075,N_41622,N_41439);
nor U42076 (N_42076,N_41324,N_41437);
xor U42077 (N_42077,N_41804,N_40785);
and U42078 (N_42078,N_41284,N_40409);
xor U42079 (N_42079,N_41173,N_40382);
or U42080 (N_42080,N_41606,N_41201);
nor U42081 (N_42081,N_41767,N_41932);
nand U42082 (N_42082,N_41098,N_40292);
and U42083 (N_42083,N_41823,N_40126);
xnor U42084 (N_42084,N_41534,N_41541);
or U42085 (N_42085,N_40652,N_41674);
and U42086 (N_42086,N_41919,N_40878);
and U42087 (N_42087,N_41347,N_40372);
or U42088 (N_42088,N_40047,N_41134);
and U42089 (N_42089,N_40517,N_40589);
and U42090 (N_42090,N_41557,N_41723);
nor U42091 (N_42091,N_41893,N_41675);
xnor U42092 (N_42092,N_40265,N_40362);
and U42093 (N_42093,N_40144,N_41929);
nor U42094 (N_42094,N_40737,N_40378);
nand U42095 (N_42095,N_40202,N_40853);
xor U42096 (N_42096,N_41972,N_40898);
xor U42097 (N_42097,N_41292,N_41688);
and U42098 (N_42098,N_41868,N_40730);
xor U42099 (N_42099,N_40420,N_40827);
or U42100 (N_42100,N_41844,N_40061);
nand U42101 (N_42101,N_41632,N_40826);
nand U42102 (N_42102,N_40108,N_41189);
nand U42103 (N_42103,N_41294,N_40738);
xor U42104 (N_42104,N_40872,N_40451);
nand U42105 (N_42105,N_41298,N_40269);
nor U42106 (N_42106,N_40778,N_40968);
nor U42107 (N_42107,N_40569,N_41390);
nor U42108 (N_42108,N_41590,N_41906);
nor U42109 (N_42109,N_41821,N_41352);
and U42110 (N_42110,N_40588,N_40487);
or U42111 (N_42111,N_40868,N_41884);
or U42112 (N_42112,N_40706,N_41360);
nor U42113 (N_42113,N_40928,N_41279);
xor U42114 (N_42114,N_41833,N_40525);
nor U42115 (N_42115,N_41671,N_40748);
or U42116 (N_42116,N_40276,N_41525);
nor U42117 (N_42117,N_41576,N_41653);
xor U42118 (N_42118,N_40685,N_40026);
and U42119 (N_42119,N_41315,N_41232);
and U42120 (N_42120,N_41734,N_40033);
xnor U42121 (N_42121,N_41815,N_41087);
xnor U42122 (N_42122,N_41370,N_41049);
nor U42123 (N_42123,N_40152,N_40908);
nand U42124 (N_42124,N_40099,N_41936);
and U42125 (N_42125,N_41020,N_41656);
or U42126 (N_42126,N_40016,N_40170);
and U42127 (N_42127,N_41041,N_41713);
or U42128 (N_42128,N_41267,N_41061);
or U42129 (N_42129,N_40399,N_40184);
nor U42130 (N_42130,N_41916,N_40790);
or U42131 (N_42131,N_41398,N_40696);
and U42132 (N_42132,N_41058,N_40205);
nor U42133 (N_42133,N_40943,N_40405);
nor U42134 (N_42134,N_41582,N_41013);
and U42135 (N_42135,N_41307,N_41253);
nor U42136 (N_42136,N_40847,N_40640);
nor U42137 (N_42137,N_41498,N_40229);
or U42138 (N_42138,N_40862,N_40115);
and U42139 (N_42139,N_41321,N_41696);
nor U42140 (N_42140,N_40920,N_41874);
xor U42141 (N_42141,N_40695,N_41357);
xnor U42142 (N_42142,N_40756,N_41170);
or U42143 (N_42143,N_40106,N_40673);
or U42144 (N_42144,N_40794,N_41668);
and U42145 (N_42145,N_41008,N_40736);
xnor U42146 (N_42146,N_41473,N_40340);
xnor U42147 (N_42147,N_41805,N_40264);
and U42148 (N_42148,N_40581,N_40488);
nor U42149 (N_42149,N_41258,N_40478);
nand U42150 (N_42150,N_41223,N_41902);
nor U42151 (N_42151,N_41107,N_41788);
nand U42152 (N_42152,N_41536,N_40658);
nand U42153 (N_42153,N_41903,N_41132);
xor U42154 (N_42154,N_40257,N_40575);
and U42155 (N_42155,N_40430,N_41581);
or U42156 (N_42156,N_41714,N_41161);
or U42157 (N_42157,N_40481,N_41565);
nor U42158 (N_42158,N_40303,N_40594);
nand U42159 (N_42159,N_41436,N_40354);
and U42160 (N_42160,N_40602,N_41184);
or U42161 (N_42161,N_41092,N_41399);
xnor U42162 (N_42162,N_41783,N_41171);
nor U42163 (N_42163,N_41985,N_40048);
xnor U42164 (N_42164,N_41413,N_41485);
or U42165 (N_42165,N_40230,N_40279);
xnor U42166 (N_42166,N_41955,N_41633);
nor U42167 (N_42167,N_40961,N_41462);
nor U42168 (N_42168,N_41680,N_41453);
nor U42169 (N_42169,N_41247,N_40113);
nor U42170 (N_42170,N_40398,N_40553);
xor U42171 (N_42171,N_41006,N_40975);
nor U42172 (N_42172,N_41265,N_41573);
xnor U42173 (N_42173,N_40784,N_41405);
or U42174 (N_42174,N_40068,N_41984);
nand U42175 (N_42175,N_41569,N_41073);
nand U42176 (N_42176,N_41203,N_41809);
or U42177 (N_42177,N_40882,N_40175);
nor U42178 (N_42178,N_40831,N_40322);
xor U42179 (N_42179,N_41187,N_41052);
xnor U42180 (N_42180,N_40997,N_40911);
and U42181 (N_42181,N_40028,N_40846);
and U42182 (N_42182,N_41262,N_41699);
and U42183 (N_42183,N_40851,N_41724);
and U42184 (N_42184,N_41358,N_41603);
nand U42185 (N_42185,N_41468,N_40460);
xor U42186 (N_42186,N_40022,N_41979);
nor U42187 (N_42187,N_41109,N_40511);
or U42188 (N_42188,N_41012,N_41085);
nor U42189 (N_42189,N_41494,N_40841);
nor U42190 (N_42190,N_40032,N_41287);
and U42191 (N_42191,N_40617,N_41281);
nand U42192 (N_42192,N_40450,N_41617);
nand U42193 (N_42193,N_40683,N_40567);
or U42194 (N_42194,N_40171,N_40570);
and U42195 (N_42195,N_40275,N_41673);
and U42196 (N_42196,N_40479,N_41445);
or U42197 (N_42197,N_40880,N_40742);
or U42198 (N_42198,N_40796,N_40601);
and U42199 (N_42199,N_40238,N_41100);
and U42200 (N_42200,N_41295,N_40788);
and U42201 (N_42201,N_40693,N_41881);
nand U42202 (N_42202,N_41497,N_41639);
and U42203 (N_42203,N_41055,N_41792);
nor U42204 (N_42204,N_40131,N_41858);
nand U42205 (N_42205,N_40884,N_41735);
and U42206 (N_42206,N_40311,N_40003);
and U42207 (N_42207,N_41167,N_41496);
nor U42208 (N_42208,N_40359,N_40100);
nor U42209 (N_42209,N_40485,N_41317);
xnor U42210 (N_42210,N_41239,N_40498);
xor U42211 (N_42211,N_41867,N_40281);
or U42212 (N_42212,N_40370,N_41377);
nor U42213 (N_42213,N_40606,N_41679);
or U42214 (N_42214,N_40072,N_40206);
or U42215 (N_42215,N_41887,N_41146);
or U42216 (N_42216,N_40422,N_40924);
or U42217 (N_42217,N_40984,N_40084);
and U42218 (N_42218,N_40743,N_41784);
and U42219 (N_42219,N_41586,N_41272);
xnor U42220 (N_42220,N_41523,N_40852);
xor U42221 (N_42221,N_41153,N_41374);
and U42222 (N_42222,N_41337,N_40544);
and U42223 (N_42223,N_41610,N_40474);
nor U42224 (N_42224,N_41616,N_40413);
or U42225 (N_42225,N_40055,N_41076);
nor U42226 (N_42226,N_40563,N_41849);
nor U42227 (N_42227,N_40668,N_40365);
or U42228 (N_42228,N_40459,N_40700);
xnor U42229 (N_42229,N_41313,N_40477);
nor U42230 (N_42230,N_41117,N_41597);
and U42231 (N_42231,N_41449,N_40074);
or U42232 (N_42232,N_40196,N_41731);
nand U42233 (N_42233,N_41432,N_41214);
or U42234 (N_42234,N_41886,N_40130);
nor U42235 (N_42235,N_41678,N_41068);
xnor U42236 (N_42236,N_40751,N_40679);
nand U42237 (N_42237,N_40501,N_41718);
nand U42238 (N_42238,N_40319,N_40043);
nor U42239 (N_42239,N_40716,N_41676);
nor U42240 (N_42240,N_41543,N_40819);
and U42241 (N_42241,N_40816,N_41240);
or U42242 (N_42242,N_41021,N_41210);
and U42243 (N_42243,N_41391,N_40240);
nor U42244 (N_42244,N_40779,N_40821);
nor U42245 (N_42245,N_40845,N_41540);
xor U42246 (N_42246,N_40998,N_41561);
xnor U42247 (N_42247,N_40226,N_40042);
nand U42248 (N_42248,N_40906,N_41199);
nand U42249 (N_42249,N_40466,N_41083);
nor U42250 (N_42250,N_41765,N_41064);
xnor U42251 (N_42251,N_40815,N_41040);
xor U42252 (N_42252,N_40665,N_41490);
and U42253 (N_42253,N_40139,N_41997);
nor U42254 (N_42254,N_41553,N_41574);
and U42255 (N_42255,N_40373,N_41957);
nor U42256 (N_42256,N_40381,N_40909);
or U42257 (N_42257,N_40535,N_40403);
and U42258 (N_42258,N_40489,N_41977);
nand U42259 (N_42259,N_40521,N_41280);
nor U42260 (N_42260,N_41641,N_41825);
nand U42261 (N_42261,N_41126,N_40935);
or U42262 (N_42262,N_40313,N_40947);
and U42263 (N_42263,N_40199,N_41728);
and U42264 (N_42264,N_40284,N_41605);
nor U42265 (N_42265,N_40353,N_40082);
or U42266 (N_42266,N_41736,N_40304);
xor U42267 (N_42267,N_40977,N_41612);
nor U42268 (N_42268,N_40015,N_41291);
and U42269 (N_42269,N_40406,N_41269);
nor U42270 (N_42270,N_41131,N_41572);
or U42271 (N_42271,N_41094,N_40160);
nand U42272 (N_42272,N_41465,N_40728);
or U42273 (N_42273,N_40194,N_41178);
nor U42274 (N_42274,N_40295,N_40809);
nand U42275 (N_42275,N_40443,N_40777);
or U42276 (N_42276,N_41548,N_41500);
nand U42277 (N_42277,N_41386,N_40191);
nand U42278 (N_42278,N_41813,N_41431);
xnor U42279 (N_42279,N_40081,N_40427);
nor U42280 (N_42280,N_41221,N_41948);
and U42281 (N_42281,N_40830,N_40659);
and U42282 (N_42282,N_40985,N_40331);
nand U42283 (N_42283,N_40509,N_41296);
nor U42284 (N_42284,N_40177,N_41387);
nor U42285 (N_42285,N_41537,N_40356);
nand U42286 (N_42286,N_40289,N_40934);
nand U42287 (N_42287,N_41556,N_41301);
or U42288 (N_42288,N_41819,N_40253);
or U42289 (N_42289,N_40957,N_40507);
and U42290 (N_42290,N_40343,N_40309);
or U42291 (N_42291,N_40165,N_41330);
nand U42292 (N_42292,N_41782,N_41433);
or U42293 (N_42293,N_40070,N_41264);
or U42294 (N_42294,N_41125,N_41506);
nand U42295 (N_42295,N_40314,N_41022);
nor U42296 (N_42296,N_41507,N_41527);
xor U42297 (N_42297,N_40927,N_40183);
nor U42298 (N_42298,N_41260,N_40060);
and U42299 (N_42299,N_41185,N_40121);
and U42300 (N_42300,N_41528,N_41212);
nor U42301 (N_42301,N_41225,N_40502);
nor U42302 (N_42302,N_41024,N_40316);
and U42303 (N_42303,N_40442,N_41290);
or U42304 (N_42304,N_41469,N_40133);
or U42305 (N_42305,N_41152,N_40005);
and U42306 (N_42306,N_41192,N_40883);
xor U42307 (N_42307,N_40225,N_41602);
nand U42308 (N_42308,N_40143,N_41082);
xnor U42309 (N_42309,N_40954,N_41004);
nand U42310 (N_42310,N_40902,N_40699);
and U42311 (N_42311,N_41194,N_40886);
and U42312 (N_42312,N_41851,N_41873);
xnor U42313 (N_42313,N_40159,N_41865);
nor U42314 (N_42314,N_41238,N_40505);
nor U42315 (N_42315,N_40008,N_40173);
nand U42316 (N_42316,N_40799,N_41560);
xnor U42317 (N_42317,N_41798,N_41050);
nand U42318 (N_42318,N_41908,N_40671);
nand U42319 (N_42319,N_40965,N_41613);
nand U42320 (N_42320,N_40578,N_40376);
and U42321 (N_42321,N_40648,N_40732);
nand U42322 (N_42322,N_41364,N_41406);
or U42323 (N_42323,N_40465,N_40369);
and U42324 (N_42324,N_41562,N_41164);
or U42325 (N_42325,N_40750,N_40027);
nor U42326 (N_42326,N_40823,N_41143);
nor U42327 (N_42327,N_41924,N_41880);
xor U42328 (N_42328,N_41634,N_40439);
xnor U42329 (N_42329,N_40893,N_40181);
xor U42330 (N_42330,N_41425,N_40426);
and U42331 (N_42331,N_40224,N_41455);
xor U42332 (N_42332,N_41103,N_41035);
nor U42333 (N_42333,N_41007,N_40052);
xor U42334 (N_42334,N_41925,N_41354);
xnor U42335 (N_42335,N_41156,N_41348);
nor U42336 (N_42336,N_40948,N_41208);
xor U42337 (N_42337,N_40494,N_41246);
nor U42338 (N_42338,N_41895,N_41619);
xnor U42339 (N_42339,N_41722,N_41244);
nor U42340 (N_42340,N_40468,N_41420);
nor U42341 (N_42341,N_40435,N_40760);
nand U42342 (N_42342,N_40991,N_40773);
and U42343 (N_42343,N_40444,N_41920);
nand U42344 (N_42344,N_41285,N_40140);
or U42345 (N_42345,N_41236,N_40755);
xnor U42346 (N_42346,N_41371,N_40988);
or U42347 (N_42347,N_40338,N_40921);
or U42348 (N_42348,N_41204,N_41694);
xor U42349 (N_42349,N_41717,N_40007);
and U42350 (N_42350,N_40250,N_41359);
nand U42351 (N_42351,N_41636,N_40452);
or U42352 (N_42352,N_40711,N_41875);
xnor U42353 (N_42353,N_41027,N_40004);
nand U42354 (N_42354,N_41276,N_40029);
nor U42355 (N_42355,N_40727,N_41624);
and U42356 (N_42356,N_41785,N_40393);
xor U42357 (N_42357,N_41853,N_41685);
nor U42358 (N_42358,N_41145,N_41786);
and U42359 (N_42359,N_41193,N_40388);
nand U42360 (N_42360,N_40187,N_41181);
nand U42361 (N_42361,N_40286,N_41752);
or U42362 (N_42362,N_40800,N_40169);
nor U42363 (N_42363,N_41057,N_41471);
nor U42364 (N_42364,N_40277,N_40243);
xnor U42365 (N_42365,N_40929,N_40075);
nand U42366 (N_42366,N_41213,N_41644);
and U42367 (N_42367,N_41128,N_40344);
xor U42368 (N_42368,N_41693,N_41029);
nand U42369 (N_42369,N_40326,N_41891);
xnor U42370 (N_42370,N_41862,N_40822);
nor U42371 (N_42371,N_40871,N_41807);
xor U42372 (N_42372,N_40753,N_41234);
nor U42373 (N_42373,N_41716,N_40881);
nor U42374 (N_42374,N_41060,N_41907);
and U42375 (N_42375,N_40059,N_41428);
xor U42376 (N_42376,N_41438,N_40707);
or U42377 (N_42377,N_40995,N_41705);
xor U42378 (N_42378,N_40608,N_41063);
or U42379 (N_42379,N_40834,N_40654);
or U42380 (N_42380,N_41422,N_41476);
xor U42381 (N_42381,N_41847,N_40835);
or U42382 (N_42382,N_41028,N_40768);
and U42383 (N_42383,N_40456,N_40677);
or U42384 (N_42384,N_40646,N_41065);
nor U42385 (N_42385,N_40955,N_40704);
nor U42386 (N_42386,N_40527,N_40129);
and U42387 (N_42387,N_41719,N_41039);
xor U42388 (N_42388,N_40318,N_40974);
nand U42389 (N_42389,N_41376,N_40766);
xor U42390 (N_42390,N_40496,N_40186);
nand U42391 (N_42391,N_41700,N_41250);
nor U42392 (N_42392,N_40508,N_40874);
nand U42393 (N_42393,N_41601,N_40649);
and U42394 (N_42394,N_40142,N_40035);
or U42395 (N_42395,N_40010,N_41524);
nand U42396 (N_42396,N_41615,N_40550);
or U42397 (N_42397,N_40682,N_41839);
nor U42398 (N_42398,N_40280,N_41830);
xnor U42399 (N_42399,N_41756,N_40270);
nand U42400 (N_42400,N_41753,N_40600);
or U42401 (N_42401,N_40215,N_40910);
or U42402 (N_42402,N_41466,N_40904);
or U42403 (N_42403,N_41927,N_41177);
or U42404 (N_42404,N_41799,N_41757);
nor U42405 (N_42405,N_40552,N_40397);
nand U42406 (N_42406,N_40689,N_40441);
xnor U42407 (N_42407,N_41744,N_41174);
nor U42408 (N_42408,N_41460,N_40616);
xor U42409 (N_42409,N_41994,N_41090);
nand U42410 (N_42410,N_40274,N_41811);
or U42411 (N_42411,N_41464,N_40447);
and U42412 (N_42412,N_41532,N_40057);
nand U42413 (N_42413,N_40971,N_41978);
and U42414 (N_42414,N_41959,N_40445);
nand U42415 (N_42415,N_41509,N_40675);
or U42416 (N_42416,N_40421,N_41278);
xor U42417 (N_42417,N_40395,N_41998);
nand U42418 (N_42418,N_40897,N_41489);
nor U42419 (N_42419,N_40661,N_40156);
or U42420 (N_42420,N_40752,N_40708);
or U42421 (N_42421,N_41768,N_40724);
and U42422 (N_42422,N_40938,N_41446);
and U42423 (N_42423,N_40351,N_41487);
nor U42424 (N_42424,N_41754,N_41817);
nand U42425 (N_42425,N_41879,N_41566);
or U42426 (N_42426,N_41772,N_41940);
or U42427 (N_42427,N_41023,N_40078);
nand U42428 (N_42428,N_40622,N_40412);
xnor U42429 (N_42429,N_40355,N_40389);
and U42430 (N_42430,N_40598,N_40166);
xor U42431 (N_42431,N_41318,N_40067);
nor U42432 (N_42432,N_40925,N_40030);
and U42433 (N_42433,N_41443,N_41914);
or U42434 (N_42434,N_40642,N_41365);
nor U42435 (N_42435,N_41794,N_40324);
nand U42436 (N_42436,N_41508,N_41099);
and U42437 (N_42437,N_41677,N_40089);
nand U42438 (N_42438,N_41789,N_41286);
xnor U42439 (N_42439,N_40025,N_40629);
nand U42440 (N_42440,N_41220,N_41312);
nand U42441 (N_42441,N_40305,N_41861);
or U42442 (N_42442,N_40620,N_41578);
nand U42443 (N_42443,N_41596,N_40534);
nand U42444 (N_42444,N_40676,N_40252);
or U42445 (N_42445,N_41254,N_41514);
xnor U42446 (N_42446,N_40619,N_41368);
or U42447 (N_42447,N_40539,N_40687);
and U42448 (N_42448,N_41956,N_40127);
and U42449 (N_42449,N_41993,N_40111);
or U42450 (N_42450,N_41892,N_40408);
and U42451 (N_42451,N_40923,N_41182);
and U42452 (N_42452,N_41059,N_40765);
xor U42453 (N_42453,N_40209,N_40371);
xor U42454 (N_42454,N_40624,N_40580);
and U42455 (N_42455,N_40380,N_41965);
xor U42456 (N_42456,N_41404,N_41224);
nand U42457 (N_42457,N_40446,N_40797);
or U42458 (N_42458,N_40500,N_40256);
nand U42459 (N_42459,N_41982,N_40227);
xor U42460 (N_42460,N_41385,N_40220);
xor U42461 (N_42461,N_40073,N_41827);
and U42462 (N_42462,N_41000,N_41604);
and U42463 (N_42463,N_41300,N_40218);
nor U42464 (N_42464,N_40999,N_40577);
nor U42465 (N_42465,N_40621,N_41255);
or U42466 (N_42466,N_41467,N_40758);
nand U42467 (N_42467,N_40425,N_40896);
or U42468 (N_42468,N_40437,N_41850);
nand U42469 (N_42469,N_41775,N_41795);
xor U42470 (N_42470,N_41609,N_40088);
nand U42471 (N_42471,N_40561,N_40377);
xor U42472 (N_42472,N_40475,N_40390);
nor U42473 (N_42473,N_41589,N_41793);
and U42474 (N_42474,N_40586,N_40278);
xnor U42475 (N_42475,N_41781,N_40385);
xor U42476 (N_42476,N_40232,N_41854);
and U42477 (N_42477,N_41787,N_40321);
or U42478 (N_42478,N_41760,N_41690);
nor U42479 (N_42479,N_40684,N_40203);
nor U42480 (N_42480,N_40944,N_41937);
nand U42481 (N_42481,N_41176,N_41518);
nor U42482 (N_42482,N_41046,N_41245);
xnor U42483 (N_42483,N_40900,N_40597);
nand U42484 (N_42484,N_40951,N_40952);
or U42485 (N_42485,N_40922,N_40669);
or U42486 (N_42486,N_41577,N_41115);
nand U42487 (N_42487,N_40560,N_40866);
and U42488 (N_42488,N_41539,N_40044);
nor U42489 (N_42489,N_41002,N_40087);
nand U42490 (N_42490,N_40564,N_41692);
or U42491 (N_42491,N_41513,N_40583);
xnor U42492 (N_42492,N_40178,N_41031);
and U42493 (N_42493,N_40764,N_41241);
or U42494 (N_42494,N_41303,N_41630);
and U42495 (N_42495,N_41911,N_41974);
and U42496 (N_42496,N_41096,N_40919);
xor U42497 (N_42497,N_40528,N_41309);
or U42498 (N_42498,N_40339,N_41138);
and U42499 (N_42499,N_41499,N_41014);
xnor U42500 (N_42500,N_40763,N_40879);
and U42501 (N_42501,N_40476,N_40960);
and U42502 (N_42502,N_41568,N_41838);
nand U42503 (N_42503,N_41730,N_41806);
or U42504 (N_42504,N_40541,N_41681);
nand U42505 (N_42505,N_40713,N_41336);
xnor U42506 (N_42506,N_40918,N_41910);
xor U42507 (N_42507,N_41663,N_40714);
nand U42508 (N_42508,N_40455,N_40915);
nand U42509 (N_42509,N_41297,N_41598);
and U42510 (N_42510,N_40429,N_40182);
or U42511 (N_42511,N_40231,N_40136);
xor U42512 (N_42512,N_41119,N_40888);
nor U42513 (N_42513,N_41069,N_41256);
or U42514 (N_42514,N_41011,N_40364);
nand U42515 (N_42515,N_40125,N_41163);
nor U42516 (N_42516,N_41950,N_41512);
nor U42517 (N_42517,N_40273,N_41197);
nand U42518 (N_42518,N_41450,N_40293);
nor U42519 (N_42519,N_41791,N_41812);
xor U42520 (N_42520,N_41381,N_41382);
nor U42521 (N_42521,N_40626,N_41456);
nand U42522 (N_42522,N_41480,N_40490);
or U42523 (N_42523,N_40591,N_41361);
or U42524 (N_42524,N_40424,N_40418);
nor U42525 (N_42525,N_40235,N_40431);
or U42526 (N_42526,N_41479,N_41659);
nand U42527 (N_42527,N_41403,N_40098);
or U42528 (N_42528,N_40978,N_40337);
nor U42529 (N_42529,N_41551,N_40516);
nand U42530 (N_42530,N_40631,N_40428);
xnor U42531 (N_42531,N_41748,N_40855);
or U42532 (N_42532,N_41409,N_41802);
and U42533 (N_42533,N_41271,N_41968);
and U42534 (N_42534,N_41415,N_41389);
nand U42535 (N_42535,N_40307,N_41658);
or U42536 (N_42536,N_40833,N_41860);
xnor U42537 (N_42537,N_41416,N_40041);
or U42538 (N_42538,N_40272,N_40046);
and U42539 (N_42539,N_41274,N_41669);
nor U42540 (N_42540,N_40932,N_41062);
nor U42541 (N_42541,N_40124,N_41261);
xnor U42542 (N_42542,N_41139,N_41319);
or U42543 (N_42543,N_41043,N_41314);
nor U42544 (N_42544,N_40655,N_41121);
or U42545 (N_42545,N_41857,N_41703);
nor U42546 (N_42546,N_41047,N_41470);
or U42547 (N_42547,N_40889,N_41643);
nand U42548 (N_42548,N_40638,N_41683);
and U42549 (N_42549,N_41188,N_40829);
nand U42550 (N_42550,N_41661,N_41750);
and U42551 (N_42551,N_40603,N_40503);
nand U42552 (N_42552,N_40050,N_40069);
nor U42553 (N_42553,N_40953,N_40198);
and U42554 (N_42554,N_41461,N_40526);
and U42555 (N_42555,N_40017,N_41747);
nor U42556 (N_42556,N_41888,N_41837);
or U42557 (N_42557,N_40762,N_40532);
xnor U42558 (N_42558,N_41162,N_41898);
nor U42559 (N_42559,N_40894,N_41441);
xor U42560 (N_42560,N_41165,N_41038);
or U42561 (N_42561,N_41990,N_41078);
nor U42562 (N_42562,N_40019,N_41017);
xor U42563 (N_42563,N_40837,N_40283);
xnor U42564 (N_42564,N_41846,N_41623);
or U42565 (N_42565,N_40383,N_41151);
xor U42566 (N_42566,N_40285,N_40949);
xnor U42567 (N_42567,N_41423,N_41822);
nand U42568 (N_42568,N_40973,N_40034);
or U42569 (N_42569,N_41664,N_41922);
nor U42570 (N_42570,N_41943,N_40367);
or U42571 (N_42571,N_41308,N_41621);
and U42572 (N_42572,N_41960,N_41531);
or U42573 (N_42573,N_41379,N_40401);
nor U42574 (N_42574,N_41550,N_40216);
nor U42575 (N_42575,N_41535,N_40291);
xor U42576 (N_42576,N_41538,N_41918);
or U42577 (N_42577,N_40471,N_40207);
nor U42578 (N_42578,N_41777,N_41072);
or U42579 (N_42579,N_40972,N_40566);
and U42580 (N_42580,N_41642,N_41339);
or U42581 (N_42581,N_41492,N_40959);
or U42582 (N_42582,N_41953,N_40247);
nand U42583 (N_42583,N_40681,N_41894);
nor U42584 (N_42584,N_40146,N_41414);
xnor U42585 (N_42585,N_41770,N_40168);
or U42586 (N_42586,N_40176,N_41575);
nor U42587 (N_42587,N_41116,N_40261);
and U42588 (N_42588,N_41305,N_41394);
or U42589 (N_42589,N_40147,N_41169);
nor U42590 (N_42590,N_41939,N_41475);
xor U42591 (N_42591,N_40533,N_41229);
xor U42592 (N_42592,N_41749,N_40522);
xor U42593 (N_42593,N_41981,N_41660);
or U42594 (N_42594,N_41901,N_40697);
nand U42595 (N_42595,N_40636,N_40754);
xnor U42596 (N_42596,N_41832,N_40260);
xnor U42597 (N_42597,N_40332,N_41652);
and U42598 (N_42598,N_40776,N_41369);
or U42599 (N_42599,N_41963,N_41564);
xnor U42600 (N_42600,N_41034,N_41931);
nor U42601 (N_42601,N_40802,N_40793);
and U42602 (N_42602,N_41712,N_41110);
xor U42603 (N_42603,N_40720,N_41463);
and U42604 (N_42604,N_41546,N_41328);
nand U42605 (N_42605,N_41005,N_40551);
nor U42606 (N_42606,N_40086,N_40244);
nor U42607 (N_42607,N_41504,N_40810);
nor U42608 (N_42608,N_40512,N_40634);
and U42609 (N_42609,N_41030,N_40549);
and U42610 (N_42610,N_40686,N_40719);
and U42611 (N_42611,N_40892,N_40110);
xnor U42612 (N_42612,N_41522,N_40219);
nor U42613 (N_42613,N_40901,N_40391);
nand U42614 (N_42614,N_40315,N_41144);
xor U42615 (N_42615,N_40287,N_40464);
nor U42616 (N_42616,N_41684,N_40688);
and U42617 (N_42617,N_41588,N_40386);
or U42618 (N_42618,N_40936,N_40132);
and U42619 (N_42619,N_41042,N_40001);
nand U42620 (N_42620,N_40939,N_41408);
nor U42621 (N_42621,N_41421,N_40128);
or U42622 (N_42622,N_41758,N_41045);
xor U42623 (N_42623,N_40703,N_40798);
nor U42624 (N_42624,N_41349,N_40066);
or U42625 (N_42625,N_40290,N_40786);
xor U42626 (N_42626,N_40328,N_40095);
and U42627 (N_42627,N_40926,N_41283);
xnor U42628 (N_42628,N_40817,N_41102);
and U42629 (N_42629,N_40407,N_40813);
nand U42630 (N_42630,N_41447,N_40849);
and U42631 (N_42631,N_40870,N_40375);
nor U42632 (N_42632,N_41010,N_40590);
xnor U42633 (N_42633,N_40733,N_41160);
or U42634 (N_42634,N_40484,N_40259);
nor U42635 (N_42635,N_41218,N_40791);
nor U42636 (N_42636,N_41019,N_41727);
nand U42637 (N_42637,N_40092,N_41054);
xor U42638 (N_42638,N_40114,N_41627);
nand U42639 (N_42639,N_40449,N_40637);
nor U42640 (N_42640,N_41219,N_40268);
or U42641 (N_42641,N_41738,N_40345);
nor U42642 (N_42642,N_41667,N_40392);
and U42643 (N_42643,N_41093,N_40077);
nor U42644 (N_42644,N_41488,N_41268);
or U42645 (N_42645,N_41356,N_40645);
and U42646 (N_42646,N_40651,N_40400);
nand U42647 (N_42647,N_41618,N_41835);
xor U42648 (N_42648,N_41587,N_40931);
or U42649 (N_42649,N_41095,N_40335);
nor U42650 (N_42650,N_40615,N_41761);
or U42651 (N_42651,N_41526,N_40722);
and U42652 (N_42652,N_41967,N_41962);
and U42653 (N_42653,N_40482,N_41217);
nor U42654 (N_42654,N_41491,N_41483);
xor U42655 (N_42655,N_41316,N_41118);
xor U42656 (N_42656,N_40134,N_40780);
or U42657 (N_42657,N_40239,N_40582);
or U42658 (N_42658,N_41183,N_41338);
nand U42659 (N_42659,N_40079,N_41175);
nor U42660 (N_42660,N_40037,N_40543);
nand U42661 (N_42661,N_41746,N_40734);
and U42662 (N_42662,N_40499,N_40986);
nand U42663 (N_42663,N_41231,N_40559);
and U42664 (N_42664,N_41944,N_40320);
nand U42665 (N_42665,N_41947,N_41411);
nand U42666 (N_42666,N_40825,N_41427);
xor U42667 (N_42667,N_41448,N_40323);
nor U42668 (N_42668,N_41111,N_40112);
nand U42669 (N_42669,N_41515,N_40091);
or U42670 (N_42670,N_40739,N_40266);
xor U42671 (N_42671,N_40558,N_40940);
xor U42672 (N_42672,N_40747,N_41808);
nor U42673 (N_42673,N_41263,N_40804);
or U42674 (N_42674,N_41033,N_41654);
or U42675 (N_42675,N_40436,N_40248);
nand U42676 (N_42676,N_41790,N_40523);
nand U42677 (N_42677,N_41478,N_41584);
nand U42678 (N_42678,N_41105,N_40434);
nand U42679 (N_42679,N_40605,N_40148);
and U42680 (N_42680,N_40317,N_40506);
nor U42681 (N_42681,N_41824,N_40832);
nor U42682 (N_42682,N_41848,N_40593);
or U42683 (N_42683,N_41558,N_41774);
or U42684 (N_42684,N_40680,N_41429);
nor U42685 (N_42685,N_40877,N_40312);
nand U42686 (N_42686,N_41155,N_41521);
xor U42687 (N_42687,N_41607,N_40789);
nor U42688 (N_42688,N_41649,N_41136);
nor U42689 (N_42689,N_41340,N_40820);
and U42690 (N_42690,N_41190,N_41552);
and U42691 (N_42691,N_41769,N_41764);
or U42692 (N_42692,N_40249,N_41628);
or U42693 (N_42693,N_40020,N_40639);
xor U42694 (N_42694,N_41334,N_40519);
and U42695 (N_42695,N_41114,N_40510);
nand U42696 (N_42696,N_40876,N_40329);
or U42697 (N_42697,N_41904,N_40222);
and U42698 (N_42698,N_40469,N_40865);
nand U42699 (N_42699,N_40610,N_40193);
and U42700 (N_42700,N_40463,N_40301);
and U42701 (N_42701,N_41650,N_40990);
xnor U42702 (N_42702,N_41122,N_41195);
nor U42703 (N_42703,N_41662,N_41003);
nor U42704 (N_42704,N_40438,N_41242);
xor U42705 (N_42705,N_40650,N_41323);
nor U42706 (N_42706,N_41166,N_40123);
and U42707 (N_42707,N_41149,N_40347);
nand U42708 (N_42708,N_40964,N_41529);
nor U42709 (N_42709,N_40630,N_41344);
nor U42710 (N_42710,N_40917,N_41179);
nor U42711 (N_42711,N_41329,N_40103);
and U42712 (N_42712,N_40085,N_41698);
or U42713 (N_42713,N_40018,N_41691);
and U42714 (N_42714,N_40208,N_41048);
or U42715 (N_42715,N_40036,N_41695);
xnor U42716 (N_42716,N_41547,N_41852);
or U42717 (N_42717,N_40657,N_40164);
nand U42718 (N_42718,N_41951,N_40962);
and U42719 (N_42719,N_40483,N_41814);
nor U42720 (N_42720,N_41454,N_41157);
xor U42721 (N_42721,N_41106,N_41112);
or U42722 (N_42722,N_41966,N_41986);
nand U42723 (N_42723,N_40363,N_41594);
nor U42724 (N_42724,N_41743,N_40228);
and U42725 (N_42725,N_41882,N_40945);
nor U42726 (N_42726,N_41333,N_40814);
and U42727 (N_42727,N_41773,N_40234);
and U42728 (N_42728,N_40769,N_40691);
and U42729 (N_42729,N_40710,N_40163);
and U42730 (N_42730,N_40783,N_41493);
and U42731 (N_42731,N_41089,N_40414);
nor U42732 (N_42732,N_41969,N_41980);
xnor U42733 (N_42733,N_40013,N_41519);
or U42734 (N_42734,N_40994,N_40848);
nor U42735 (N_42735,N_41402,N_41555);
and U42736 (N_42736,N_41629,N_40192);
xnor U42737 (N_42737,N_41580,N_41614);
xor U42738 (N_42738,N_41410,N_40096);
or U42739 (N_42739,N_41935,N_40415);
xnor U42740 (N_42740,N_40093,N_40867);
or U42741 (N_42741,N_40090,N_41810);
nor U42742 (N_42742,N_40053,N_41826);
nand U42743 (N_42743,N_41407,N_40613);
xnor U42744 (N_42744,N_40242,N_40993);
nand U42745 (N_42745,N_41870,N_40656);
nand U42746 (N_42746,N_41036,N_40930);
nand U42747 (N_42747,N_41141,N_41018);
xnor U42748 (N_42748,N_41320,N_40298);
xor U42749 (N_42749,N_41215,N_41230);
and U42750 (N_42750,N_40157,N_41074);
nor U42751 (N_42751,N_40063,N_41708);
and U42752 (N_42752,N_41954,N_41530);
nand U42753 (N_42753,N_40520,N_40647);
xnor U42754 (N_42754,N_41834,N_41520);
or U42755 (N_42755,N_40122,N_41745);
and U42756 (N_42756,N_40213,N_40767);
or U42757 (N_42757,N_41159,N_40155);
nor U42758 (N_42758,N_41293,N_40903);
or U42759 (N_42759,N_40120,N_41345);
or U42760 (N_42760,N_41554,N_40263);
xor U42761 (N_42761,N_40774,N_41158);
nor U42762 (N_42762,N_40854,N_40690);
or U42763 (N_42763,N_40470,N_40379);
or U42764 (N_42764,N_41776,N_40803);
xor U42765 (N_42765,N_40698,N_41383);
or U42766 (N_42766,N_40384,N_41266);
nor U42767 (N_42767,N_41077,N_40987);
nand U42768 (N_42768,N_41942,N_40040);
or U42769 (N_42769,N_40933,N_40497);
nand U42770 (N_42770,N_41666,N_41299);
nand U42771 (N_42771,N_41282,N_40109);
nand U42772 (N_42772,N_41457,N_40083);
or U42773 (N_42773,N_41591,N_40387);
xor U42774 (N_42774,N_41372,N_40633);
and U42775 (N_42775,N_41992,N_40141);
xnor U42776 (N_42776,N_41945,N_41451);
nor U42777 (N_42777,N_40678,N_41362);
and U42778 (N_42778,N_40942,N_41237);
xnor U42779 (N_42779,N_40480,N_40856);
xnor U42780 (N_42780,N_41142,N_41905);
and U42781 (N_42781,N_41251,N_40757);
or U42782 (N_42782,N_41209,N_41395);
nor U42783 (N_42783,N_40749,N_40614);
xnor U42784 (N_42784,N_40368,N_41665);
or U42785 (N_42785,N_41740,N_41640);
and U42786 (N_42786,N_40530,N_40555);
nand U42787 (N_42787,N_40417,N_40861);
nand U42788 (N_42788,N_41646,N_41544);
nand U42789 (N_42789,N_40542,N_40267);
or U42790 (N_42790,N_41545,N_41913);
or U42791 (N_42791,N_41335,N_40190);
nand U42792 (N_42792,N_41739,N_40179);
nor U42793 (N_42793,N_40195,N_40565);
nor U42794 (N_42794,N_40302,N_40394);
nand U42795 (N_42795,N_41133,N_41648);
nand U42796 (N_42796,N_41129,N_40741);
or U42797 (N_42797,N_41983,N_41579);
nor U42798 (N_42798,N_40352,N_41472);
and U42799 (N_42799,N_40334,N_40670);
nand U42800 (N_42800,N_40006,N_40573);
nor U42801 (N_42801,N_40557,N_41288);
xnor U42802 (N_42802,N_41921,N_40325);
and U42803 (N_42803,N_40101,N_41933);
or U42804 (N_42804,N_40571,N_41331);
nand U42805 (N_42805,N_41706,N_40031);
xnor U42806 (N_42806,N_40980,N_40761);
xor U42807 (N_42807,N_41434,N_40461);
xnor U42808 (N_42808,N_41855,N_40255);
and U42809 (N_42809,N_41243,N_41592);
nor U42810 (N_42810,N_41108,N_40587);
nand U42811 (N_42811,N_41353,N_40653);
nand U42812 (N_42812,N_40912,N_41393);
xor U42813 (N_42813,N_41346,N_41341);
or U42814 (N_42814,N_40038,N_41721);
nor U42815 (N_42815,N_41016,N_40664);
xnor U42816 (N_42816,N_41367,N_41249);
xnor U42817 (N_42817,N_40473,N_41631);
or U42818 (N_42818,N_40970,N_40718);
or U42819 (N_42819,N_40891,N_40357);
nor U42820 (N_42820,N_40844,N_40989);
and U42821 (N_42821,N_41816,N_41401);
or U42822 (N_42822,N_41946,N_40976);
and U42823 (N_42823,N_41001,N_40021);
or U42824 (N_42824,N_40336,N_40946);
xnor U42825 (N_42825,N_40585,N_41228);
nor U42826 (N_42826,N_40518,N_40251);
or U42827 (N_42827,N_41608,N_40342);
nand U42828 (N_42828,N_41732,N_41583);
xnor U42829 (N_42829,N_41056,N_41687);
nor U42830 (N_42830,N_40836,N_40937);
nand U42831 (N_42831,N_41635,N_40723);
xnor U42832 (N_42832,N_41701,N_40204);
xor U42833 (N_42833,N_40094,N_40969);
nand U42834 (N_42834,N_40162,N_40423);
and U42835 (N_42835,N_41988,N_40145);
xor U42836 (N_42836,N_41440,N_41704);
nor U42837 (N_42837,N_40361,N_41976);
xnor U42838 (N_42838,N_41996,N_40457);
nand U42839 (N_42839,N_40996,N_41517);
nand U42840 (N_42840,N_41709,N_41430);
nand U42841 (N_42841,N_40725,N_41725);
or U42842 (N_42842,N_41289,N_40440);
and U42843 (N_42843,N_41477,N_41600);
nand U42844 (N_42844,N_40271,N_40759);
nor U42845 (N_42845,N_41871,N_40956);
nor U42846 (N_42846,N_41200,N_41866);
and U42847 (N_42847,N_41384,N_41009);
or U42848 (N_42848,N_40981,N_40705);
and U42849 (N_42849,N_40538,N_40858);
or U42850 (N_42850,N_40076,N_40282);
and U42851 (N_42851,N_40721,N_40712);
nand U42852 (N_42852,N_41686,N_40358);
or U42853 (N_42853,N_40346,N_40992);
or U42854 (N_42854,N_40576,N_41975);
or U42855 (N_42855,N_40180,N_40672);
or U42856 (N_42856,N_41412,N_40495);
nand U42857 (N_42857,N_40746,N_40396);
and U42858 (N_42858,N_40536,N_41778);
nor U42859 (N_42859,N_40850,N_41930);
and U42860 (N_42860,N_40740,N_41191);
and U42861 (N_42861,N_41828,N_41032);
or U42862 (N_42862,N_40812,N_40167);
and U42863 (N_42863,N_41306,N_40117);
xor U42864 (N_42864,N_40102,N_41585);
or U42865 (N_42865,N_40065,N_41567);
or U42866 (N_42866,N_40062,N_40966);
and U42867 (N_42867,N_41836,N_41363);
or U42868 (N_42868,N_41207,N_40327);
and U42869 (N_42869,N_41928,N_41442);
nor U42870 (N_42870,N_41733,N_40404);
and U42871 (N_42871,N_41970,N_41120);
xnor U42872 (N_42872,N_41026,N_41820);
or U42873 (N_42873,N_40726,N_40958);
nor U42874 (N_42874,N_40635,N_40781);
nor U42875 (N_42875,N_41559,N_41952);
nor U42876 (N_42876,N_40771,N_40151);
nor U42877 (N_42877,N_41863,N_41964);
xnor U42878 (N_42878,N_40735,N_41570);
nor U42879 (N_42879,N_40702,N_40448);
nor U42880 (N_42880,N_41135,N_40237);
or U42881 (N_42881,N_41877,N_41419);
and U42882 (N_42882,N_41226,N_41780);
and U42883 (N_42883,N_40572,N_41710);
xor U42884 (N_42884,N_41737,N_41343);
nand U42885 (N_42885,N_40562,N_41452);
nand U42886 (N_42886,N_40288,N_41397);
and U42887 (N_42887,N_40843,N_40838);
xnor U42888 (N_42888,N_41926,N_40104);
nor U42889 (N_42889,N_41751,N_40012);
nor U42890 (N_42890,N_40051,N_41549);
nand U42891 (N_42891,N_40308,N_40023);
nand U42892 (N_42892,N_41626,N_41620);
or U42893 (N_42893,N_40545,N_41304);
nor U42894 (N_42894,N_41222,N_40245);
and U42895 (N_42895,N_41459,N_41322);
xor U42896 (N_42896,N_41670,N_40701);
nand U42897 (N_42897,N_40983,N_41067);
and U42898 (N_42898,N_41486,N_40118);
nor U42899 (N_42899,N_40107,N_40895);
nand U42900 (N_42900,N_41771,N_41949);
xnor U42901 (N_42901,N_40568,N_41505);
or U42902 (N_42902,N_41051,N_41638);
or U42903 (N_42903,N_40963,N_40899);
xnor U42904 (N_42904,N_41934,N_41326);
or U42905 (N_42905,N_40662,N_40472);
xor U42906 (N_42906,N_40493,N_41375);
nand U42907 (N_42907,N_40729,N_41091);
nor U42908 (N_42908,N_41474,N_40540);
xor U42909 (N_42909,N_40531,N_41172);
or U42910 (N_42910,N_41444,N_41502);
or U42911 (N_42911,N_40161,N_40775);
and U42912 (N_42912,N_40515,N_41637);
xor U42913 (N_42913,N_40200,N_40839);
xor U42914 (N_42914,N_41510,N_40300);
and U42915 (N_42915,N_41599,N_40574);
nor U42916 (N_42916,N_41075,N_40806);
xor U42917 (N_42917,N_41818,N_41227);
xnor U42918 (N_42918,N_41137,N_40211);
nor U42919 (N_42919,N_40002,N_41426);
or U42920 (N_42920,N_40241,N_40411);
or U42921 (N_42921,N_40348,N_41864);
nand U42922 (N_42922,N_40153,N_40492);
nor U42923 (N_42923,N_40537,N_40859);
nand U42924 (N_42924,N_41800,N_40623);
nand U42925 (N_42925,N_40214,N_41923);
xor U42926 (N_42926,N_40625,N_41672);
nor U42927 (N_42927,N_41726,N_41168);
and U42928 (N_42928,N_40432,N_40360);
and U42929 (N_42929,N_41378,N_41424);
or U42930 (N_42930,N_40236,N_41080);
nor U42931 (N_42931,N_41233,N_40049);
and U42932 (N_42932,N_40453,N_40454);
nor U42933 (N_42933,N_41909,N_41327);
nand U42934 (N_42934,N_40349,N_41275);
xnor U42935 (N_42935,N_40546,N_40885);
or U42936 (N_42936,N_40529,N_40097);
nor U42937 (N_42937,N_41302,N_41196);
xnor U42938 (N_42938,N_41702,N_41845);
nand U42939 (N_42939,N_40189,N_41843);
nand U42940 (N_42940,N_40618,N_40627);
nand U42941 (N_42941,N_40592,N_40310);
or U42942 (N_42942,N_41418,N_41831);
or U42943 (N_42943,N_40612,N_40641);
nor U42944 (N_42944,N_41657,N_41856);
nand U42945 (N_42945,N_41355,N_41729);
nand U42946 (N_42946,N_41198,N_40808);
and U42947 (N_42947,N_41053,N_41682);
xnor U42948 (N_42948,N_40137,N_41841);
or U42949 (N_42949,N_40795,N_40410);
and U42950 (N_42950,N_41878,N_41842);
nand U42951 (N_42951,N_41044,N_41796);
nand U42952 (N_42952,N_40462,N_40770);
and U42953 (N_42953,N_40433,N_40890);
or U42954 (N_42954,N_41989,N_40514);
nor U42955 (N_42955,N_40011,N_40715);
and U42956 (N_42956,N_41563,N_40869);
nand U42957 (N_42957,N_40333,N_40787);
and U42958 (N_42958,N_41707,N_40116);
xor U42959 (N_42959,N_41101,N_41325);
and U42960 (N_42960,N_40914,N_40058);
nand U42961 (N_42961,N_41991,N_41070);
or U42962 (N_42962,N_40341,N_40818);
xnor U42963 (N_42963,N_41840,N_40905);
nor U42964 (N_42964,N_40873,N_41086);
nor U42965 (N_42965,N_40663,N_41435);
or U42966 (N_42966,N_41037,N_41277);
nor U42967 (N_42967,N_40024,N_40628);
or U42968 (N_42968,N_40296,N_41872);
nor U42969 (N_42969,N_41516,N_40611);
nor U42970 (N_42970,N_41763,N_40584);
or U42971 (N_42971,N_41066,N_40941);
xor U42972 (N_42972,N_41938,N_41104);
and U42973 (N_42973,N_40744,N_40782);
and U42974 (N_42974,N_41252,N_41885);
or U42975 (N_42975,N_40607,N_40666);
and U42976 (N_42976,N_41533,N_40887);
or U42977 (N_42977,N_40306,N_40212);
nor U42978 (N_42978,N_41755,N_40419);
nor U42979 (N_42979,N_41876,N_40105);
or U42980 (N_42980,N_40504,N_41350);
xor U42981 (N_42981,N_41332,N_41715);
or U42982 (N_42982,N_41235,N_40185);
xor U42983 (N_42983,N_41511,N_41869);
xnor U42984 (N_42984,N_41890,N_40864);
nand U42985 (N_42985,N_41123,N_41917);
or U42986 (N_42986,N_40916,N_40014);
and U42987 (N_42987,N_40667,N_41915);
xnor U42988 (N_42988,N_40792,N_41741);
nand U42989 (N_42989,N_40967,N_40071);
nand U42990 (N_42990,N_40064,N_40717);
nand U42991 (N_42991,N_40149,N_41651);
nor U42992 (N_42992,N_41647,N_41971);
xnor U42993 (N_42993,N_41912,N_40579);
or U42994 (N_42994,N_41147,N_41897);
nand U42995 (N_42995,N_40857,N_41762);
nor U42996 (N_42996,N_41611,N_41079);
and U42997 (N_42997,N_41084,N_40907);
nor U42998 (N_42998,N_41417,N_41259);
xnor U42999 (N_42999,N_41154,N_40644);
and U43000 (N_43000,N_41578,N_40754);
nand U43001 (N_43001,N_40322,N_40250);
xnor U43002 (N_43002,N_41835,N_41350);
and U43003 (N_43003,N_40190,N_41843);
nand U43004 (N_43004,N_41545,N_41580);
xnor U43005 (N_43005,N_40972,N_40100);
and U43006 (N_43006,N_40029,N_40514);
nor U43007 (N_43007,N_40930,N_40034);
nand U43008 (N_43008,N_40986,N_40232);
nor U43009 (N_43009,N_41545,N_41630);
nor U43010 (N_43010,N_41034,N_40363);
or U43011 (N_43011,N_40919,N_41474);
nand U43012 (N_43012,N_40689,N_41671);
and U43013 (N_43013,N_41142,N_41831);
or U43014 (N_43014,N_41384,N_40035);
xnor U43015 (N_43015,N_41181,N_40273);
xnor U43016 (N_43016,N_40008,N_40193);
or U43017 (N_43017,N_40883,N_41732);
or U43018 (N_43018,N_40205,N_41382);
or U43019 (N_43019,N_41907,N_41537);
and U43020 (N_43020,N_41091,N_40302);
or U43021 (N_43021,N_40040,N_40487);
nand U43022 (N_43022,N_40356,N_41487);
nand U43023 (N_43023,N_40640,N_41672);
xor U43024 (N_43024,N_41837,N_40773);
or U43025 (N_43025,N_40763,N_41077);
nand U43026 (N_43026,N_41132,N_40299);
or U43027 (N_43027,N_41993,N_41858);
or U43028 (N_43028,N_40884,N_41587);
nor U43029 (N_43029,N_40022,N_41097);
nor U43030 (N_43030,N_40569,N_41555);
nand U43031 (N_43031,N_40153,N_41976);
xor U43032 (N_43032,N_40389,N_41468);
nand U43033 (N_43033,N_41851,N_40073);
nand U43034 (N_43034,N_41066,N_40843);
nand U43035 (N_43035,N_41145,N_41031);
nand U43036 (N_43036,N_41736,N_40862);
nor U43037 (N_43037,N_41262,N_40905);
nand U43038 (N_43038,N_41291,N_41464);
nand U43039 (N_43039,N_40293,N_40266);
or U43040 (N_43040,N_40985,N_41616);
nand U43041 (N_43041,N_40010,N_41617);
and U43042 (N_43042,N_40545,N_40233);
or U43043 (N_43043,N_41225,N_41478);
or U43044 (N_43044,N_40764,N_41049);
nor U43045 (N_43045,N_40220,N_40629);
or U43046 (N_43046,N_41615,N_40332);
and U43047 (N_43047,N_41044,N_40164);
and U43048 (N_43048,N_41177,N_40451);
and U43049 (N_43049,N_41896,N_40830);
or U43050 (N_43050,N_41781,N_40005);
or U43051 (N_43051,N_41744,N_40265);
nand U43052 (N_43052,N_40248,N_41612);
nand U43053 (N_43053,N_40649,N_40003);
and U43054 (N_43054,N_40061,N_41558);
nor U43055 (N_43055,N_40634,N_41400);
nand U43056 (N_43056,N_41097,N_41514);
and U43057 (N_43057,N_40477,N_41366);
xor U43058 (N_43058,N_41050,N_41947);
and U43059 (N_43059,N_40024,N_41374);
and U43060 (N_43060,N_40566,N_41139);
or U43061 (N_43061,N_40654,N_41408);
nand U43062 (N_43062,N_40721,N_41036);
nor U43063 (N_43063,N_41790,N_41797);
or U43064 (N_43064,N_40342,N_40512);
nand U43065 (N_43065,N_41106,N_41834);
nor U43066 (N_43066,N_40955,N_40548);
nand U43067 (N_43067,N_41616,N_41150);
nor U43068 (N_43068,N_40388,N_41204);
or U43069 (N_43069,N_40070,N_40137);
nand U43070 (N_43070,N_40270,N_41901);
nor U43071 (N_43071,N_41201,N_41782);
and U43072 (N_43072,N_40001,N_40809);
nor U43073 (N_43073,N_40811,N_41267);
nand U43074 (N_43074,N_40693,N_40904);
and U43075 (N_43075,N_41487,N_40096);
nand U43076 (N_43076,N_41479,N_40067);
xnor U43077 (N_43077,N_40655,N_40825);
or U43078 (N_43078,N_41623,N_41289);
nand U43079 (N_43079,N_41936,N_40475);
nand U43080 (N_43080,N_40208,N_41621);
and U43081 (N_43081,N_40486,N_40435);
or U43082 (N_43082,N_41465,N_40328);
nor U43083 (N_43083,N_41497,N_41993);
nor U43084 (N_43084,N_41500,N_40862);
nand U43085 (N_43085,N_41814,N_40284);
or U43086 (N_43086,N_41453,N_41475);
and U43087 (N_43087,N_41392,N_40113);
or U43088 (N_43088,N_41763,N_40092);
nor U43089 (N_43089,N_40834,N_41293);
nand U43090 (N_43090,N_40745,N_41958);
nand U43091 (N_43091,N_41006,N_40073);
nand U43092 (N_43092,N_40747,N_40033);
nand U43093 (N_43093,N_41018,N_40696);
or U43094 (N_43094,N_40630,N_40661);
or U43095 (N_43095,N_41492,N_40368);
xnor U43096 (N_43096,N_41350,N_41408);
or U43097 (N_43097,N_40377,N_40245);
xnor U43098 (N_43098,N_41932,N_40386);
or U43099 (N_43099,N_41125,N_40184);
xor U43100 (N_43100,N_41612,N_41173);
and U43101 (N_43101,N_40516,N_40521);
xor U43102 (N_43102,N_40860,N_40329);
or U43103 (N_43103,N_40997,N_41194);
or U43104 (N_43104,N_40751,N_40040);
or U43105 (N_43105,N_40826,N_41661);
xnor U43106 (N_43106,N_40298,N_40796);
nand U43107 (N_43107,N_40507,N_40009);
or U43108 (N_43108,N_40449,N_41376);
nand U43109 (N_43109,N_41867,N_40196);
and U43110 (N_43110,N_40543,N_41547);
nor U43111 (N_43111,N_40548,N_40809);
nand U43112 (N_43112,N_41872,N_41481);
and U43113 (N_43113,N_41136,N_40729);
and U43114 (N_43114,N_41927,N_40071);
or U43115 (N_43115,N_41081,N_41770);
nor U43116 (N_43116,N_40235,N_41937);
nor U43117 (N_43117,N_41003,N_40244);
nor U43118 (N_43118,N_41240,N_41442);
nor U43119 (N_43119,N_40570,N_41547);
nor U43120 (N_43120,N_40626,N_40812);
and U43121 (N_43121,N_41529,N_41796);
and U43122 (N_43122,N_40894,N_41335);
xnor U43123 (N_43123,N_41510,N_41418);
xnor U43124 (N_43124,N_41285,N_41350);
nand U43125 (N_43125,N_41509,N_40436);
nor U43126 (N_43126,N_41146,N_40633);
nand U43127 (N_43127,N_40802,N_40103);
and U43128 (N_43128,N_40861,N_41651);
nand U43129 (N_43129,N_41642,N_40635);
or U43130 (N_43130,N_40111,N_41032);
and U43131 (N_43131,N_41589,N_41567);
xnor U43132 (N_43132,N_41790,N_41019);
nand U43133 (N_43133,N_41040,N_40823);
nor U43134 (N_43134,N_41870,N_40715);
or U43135 (N_43135,N_41785,N_40018);
nor U43136 (N_43136,N_41414,N_41022);
and U43137 (N_43137,N_40383,N_41495);
xor U43138 (N_43138,N_40002,N_41251);
nor U43139 (N_43139,N_40157,N_41541);
nor U43140 (N_43140,N_41171,N_41168);
nor U43141 (N_43141,N_40946,N_40131);
xor U43142 (N_43142,N_41704,N_41957);
nand U43143 (N_43143,N_40682,N_40611);
or U43144 (N_43144,N_40122,N_40286);
nand U43145 (N_43145,N_41096,N_40983);
and U43146 (N_43146,N_40683,N_41923);
or U43147 (N_43147,N_41386,N_41239);
and U43148 (N_43148,N_40326,N_40368);
or U43149 (N_43149,N_40081,N_41306);
and U43150 (N_43150,N_41624,N_40800);
nor U43151 (N_43151,N_41110,N_41632);
or U43152 (N_43152,N_40890,N_41748);
and U43153 (N_43153,N_41010,N_41152);
nor U43154 (N_43154,N_41863,N_41752);
nand U43155 (N_43155,N_41268,N_41609);
nor U43156 (N_43156,N_40981,N_41062);
xnor U43157 (N_43157,N_41326,N_41132);
xor U43158 (N_43158,N_40274,N_40589);
nand U43159 (N_43159,N_40244,N_41815);
and U43160 (N_43160,N_40846,N_41384);
and U43161 (N_43161,N_40651,N_41425);
or U43162 (N_43162,N_40359,N_41453);
and U43163 (N_43163,N_40225,N_41017);
nand U43164 (N_43164,N_40595,N_40766);
or U43165 (N_43165,N_41398,N_40318);
or U43166 (N_43166,N_41365,N_40000);
or U43167 (N_43167,N_40961,N_41742);
nand U43168 (N_43168,N_41964,N_41288);
and U43169 (N_43169,N_40292,N_40742);
or U43170 (N_43170,N_41397,N_40937);
nand U43171 (N_43171,N_41510,N_40485);
or U43172 (N_43172,N_40085,N_40376);
and U43173 (N_43173,N_40502,N_40362);
nor U43174 (N_43174,N_41918,N_40491);
and U43175 (N_43175,N_40424,N_41592);
or U43176 (N_43176,N_40575,N_41406);
nand U43177 (N_43177,N_41785,N_40055);
nand U43178 (N_43178,N_40467,N_40521);
and U43179 (N_43179,N_41354,N_40413);
xnor U43180 (N_43180,N_40011,N_41986);
and U43181 (N_43181,N_40046,N_40694);
xor U43182 (N_43182,N_40777,N_41783);
nand U43183 (N_43183,N_40164,N_40079);
and U43184 (N_43184,N_41435,N_40176);
nand U43185 (N_43185,N_40976,N_41483);
nor U43186 (N_43186,N_40245,N_40980);
or U43187 (N_43187,N_40509,N_41167);
and U43188 (N_43188,N_40043,N_40805);
or U43189 (N_43189,N_40397,N_40950);
and U43190 (N_43190,N_41619,N_40983);
xor U43191 (N_43191,N_40980,N_41917);
xor U43192 (N_43192,N_40958,N_40113);
nor U43193 (N_43193,N_40304,N_40674);
nand U43194 (N_43194,N_41227,N_40049);
or U43195 (N_43195,N_40232,N_40450);
or U43196 (N_43196,N_41677,N_41813);
or U43197 (N_43197,N_40990,N_40522);
or U43198 (N_43198,N_40885,N_41244);
or U43199 (N_43199,N_41633,N_41124);
or U43200 (N_43200,N_41427,N_41591);
nand U43201 (N_43201,N_41643,N_40485);
nor U43202 (N_43202,N_41151,N_41588);
nand U43203 (N_43203,N_41898,N_41830);
and U43204 (N_43204,N_41478,N_41257);
and U43205 (N_43205,N_41482,N_41532);
nor U43206 (N_43206,N_40729,N_41581);
or U43207 (N_43207,N_40772,N_40860);
nand U43208 (N_43208,N_40758,N_41647);
and U43209 (N_43209,N_41676,N_41246);
nor U43210 (N_43210,N_41355,N_40824);
xnor U43211 (N_43211,N_41083,N_40157);
xor U43212 (N_43212,N_40423,N_40295);
nand U43213 (N_43213,N_40519,N_41716);
nand U43214 (N_43214,N_40182,N_40998);
nor U43215 (N_43215,N_40658,N_41109);
xor U43216 (N_43216,N_41740,N_41911);
nand U43217 (N_43217,N_41539,N_41290);
or U43218 (N_43218,N_41582,N_40479);
nor U43219 (N_43219,N_40299,N_41254);
nor U43220 (N_43220,N_41069,N_41923);
and U43221 (N_43221,N_41569,N_40616);
and U43222 (N_43222,N_40012,N_41933);
nor U43223 (N_43223,N_40572,N_41709);
nand U43224 (N_43224,N_40726,N_41758);
nand U43225 (N_43225,N_41076,N_41648);
xnor U43226 (N_43226,N_40763,N_40217);
xnor U43227 (N_43227,N_40310,N_41188);
nand U43228 (N_43228,N_41564,N_41998);
and U43229 (N_43229,N_40731,N_41599);
xnor U43230 (N_43230,N_41688,N_40471);
or U43231 (N_43231,N_40097,N_40317);
nor U43232 (N_43232,N_40947,N_40194);
or U43233 (N_43233,N_40674,N_40651);
and U43234 (N_43234,N_41031,N_41100);
and U43235 (N_43235,N_40687,N_41823);
nand U43236 (N_43236,N_40206,N_40942);
xnor U43237 (N_43237,N_40325,N_40344);
or U43238 (N_43238,N_41617,N_41861);
xnor U43239 (N_43239,N_40719,N_41760);
nand U43240 (N_43240,N_40667,N_41437);
or U43241 (N_43241,N_41217,N_40607);
nand U43242 (N_43242,N_41276,N_41176);
nand U43243 (N_43243,N_41147,N_41051);
nor U43244 (N_43244,N_40416,N_40189);
and U43245 (N_43245,N_40313,N_40043);
xnor U43246 (N_43246,N_40297,N_41229);
nor U43247 (N_43247,N_41523,N_40850);
and U43248 (N_43248,N_41981,N_40387);
and U43249 (N_43249,N_41416,N_40744);
or U43250 (N_43250,N_40415,N_41739);
nand U43251 (N_43251,N_40905,N_41692);
nor U43252 (N_43252,N_40800,N_40468);
nor U43253 (N_43253,N_41657,N_41948);
xnor U43254 (N_43254,N_41446,N_40066);
nand U43255 (N_43255,N_41182,N_40429);
nor U43256 (N_43256,N_40142,N_41436);
and U43257 (N_43257,N_41947,N_40629);
nor U43258 (N_43258,N_41477,N_40672);
nor U43259 (N_43259,N_40844,N_41034);
xnor U43260 (N_43260,N_41057,N_41987);
xnor U43261 (N_43261,N_41443,N_41536);
or U43262 (N_43262,N_41408,N_40767);
or U43263 (N_43263,N_41857,N_41825);
nor U43264 (N_43264,N_40139,N_41563);
nand U43265 (N_43265,N_41589,N_40538);
or U43266 (N_43266,N_41333,N_40428);
nand U43267 (N_43267,N_41081,N_41266);
or U43268 (N_43268,N_41281,N_40769);
nor U43269 (N_43269,N_40982,N_40269);
or U43270 (N_43270,N_40400,N_40298);
xor U43271 (N_43271,N_40721,N_41342);
xor U43272 (N_43272,N_40556,N_41463);
nand U43273 (N_43273,N_40368,N_41745);
xnor U43274 (N_43274,N_41341,N_41939);
nand U43275 (N_43275,N_40275,N_40870);
or U43276 (N_43276,N_40418,N_41108);
and U43277 (N_43277,N_40034,N_41622);
nand U43278 (N_43278,N_41830,N_40357);
nand U43279 (N_43279,N_40995,N_40218);
or U43280 (N_43280,N_41530,N_40832);
or U43281 (N_43281,N_41911,N_40016);
nand U43282 (N_43282,N_40903,N_40113);
and U43283 (N_43283,N_40791,N_41030);
nand U43284 (N_43284,N_40698,N_40889);
or U43285 (N_43285,N_40523,N_40865);
nand U43286 (N_43286,N_41229,N_41608);
xnor U43287 (N_43287,N_41863,N_40781);
nor U43288 (N_43288,N_40306,N_41452);
nor U43289 (N_43289,N_40611,N_41903);
and U43290 (N_43290,N_40258,N_41734);
xnor U43291 (N_43291,N_41148,N_41446);
nor U43292 (N_43292,N_41168,N_40827);
and U43293 (N_43293,N_40121,N_40977);
nor U43294 (N_43294,N_41418,N_40369);
xnor U43295 (N_43295,N_41880,N_40226);
or U43296 (N_43296,N_41601,N_40462);
or U43297 (N_43297,N_40478,N_40409);
xor U43298 (N_43298,N_40506,N_41136);
xnor U43299 (N_43299,N_41171,N_40261);
xor U43300 (N_43300,N_41736,N_41898);
or U43301 (N_43301,N_40715,N_41007);
xor U43302 (N_43302,N_40303,N_41838);
xor U43303 (N_43303,N_41712,N_40881);
nand U43304 (N_43304,N_41434,N_41500);
and U43305 (N_43305,N_41464,N_40861);
nand U43306 (N_43306,N_40435,N_41711);
or U43307 (N_43307,N_40520,N_40657);
nand U43308 (N_43308,N_40335,N_41955);
nand U43309 (N_43309,N_40673,N_41749);
or U43310 (N_43310,N_41362,N_40987);
or U43311 (N_43311,N_40197,N_40124);
nand U43312 (N_43312,N_40903,N_41456);
or U43313 (N_43313,N_41704,N_41695);
or U43314 (N_43314,N_41499,N_40645);
and U43315 (N_43315,N_41219,N_40656);
and U43316 (N_43316,N_41696,N_41539);
or U43317 (N_43317,N_41328,N_41083);
or U43318 (N_43318,N_41328,N_40680);
xor U43319 (N_43319,N_40633,N_40687);
nand U43320 (N_43320,N_41191,N_41020);
or U43321 (N_43321,N_41656,N_40204);
nand U43322 (N_43322,N_40657,N_40479);
or U43323 (N_43323,N_40665,N_40041);
nor U43324 (N_43324,N_41354,N_40729);
xor U43325 (N_43325,N_41057,N_41555);
and U43326 (N_43326,N_41435,N_41698);
or U43327 (N_43327,N_40802,N_41241);
and U43328 (N_43328,N_41076,N_40939);
nor U43329 (N_43329,N_41887,N_40343);
nor U43330 (N_43330,N_41937,N_41321);
nor U43331 (N_43331,N_41322,N_41354);
or U43332 (N_43332,N_40875,N_40185);
or U43333 (N_43333,N_41235,N_40123);
or U43334 (N_43334,N_41389,N_41711);
xor U43335 (N_43335,N_40723,N_41379);
or U43336 (N_43336,N_40495,N_41312);
xor U43337 (N_43337,N_41274,N_40737);
or U43338 (N_43338,N_41904,N_41378);
nor U43339 (N_43339,N_40526,N_40191);
and U43340 (N_43340,N_41600,N_40939);
or U43341 (N_43341,N_40765,N_41123);
nand U43342 (N_43342,N_41406,N_40485);
nor U43343 (N_43343,N_40472,N_40655);
nor U43344 (N_43344,N_40102,N_40085);
or U43345 (N_43345,N_40711,N_40476);
xnor U43346 (N_43346,N_40937,N_40386);
xnor U43347 (N_43347,N_41789,N_41540);
nor U43348 (N_43348,N_40108,N_41051);
and U43349 (N_43349,N_41207,N_40869);
and U43350 (N_43350,N_40032,N_40610);
nor U43351 (N_43351,N_40092,N_40875);
nor U43352 (N_43352,N_40556,N_40308);
or U43353 (N_43353,N_41143,N_40721);
nor U43354 (N_43354,N_40812,N_41196);
xor U43355 (N_43355,N_40727,N_41857);
nor U43356 (N_43356,N_41361,N_41722);
nor U43357 (N_43357,N_40408,N_40869);
or U43358 (N_43358,N_40296,N_41307);
and U43359 (N_43359,N_41768,N_41731);
nand U43360 (N_43360,N_40408,N_40235);
or U43361 (N_43361,N_41120,N_40144);
xor U43362 (N_43362,N_40214,N_41743);
and U43363 (N_43363,N_40593,N_41695);
and U43364 (N_43364,N_40342,N_40667);
nor U43365 (N_43365,N_41171,N_40540);
and U43366 (N_43366,N_40706,N_41959);
or U43367 (N_43367,N_41914,N_41786);
xnor U43368 (N_43368,N_40828,N_40703);
xnor U43369 (N_43369,N_41563,N_40618);
and U43370 (N_43370,N_41527,N_41929);
nand U43371 (N_43371,N_41325,N_41959);
nand U43372 (N_43372,N_40720,N_40677);
nor U43373 (N_43373,N_41232,N_40079);
or U43374 (N_43374,N_41747,N_41167);
nor U43375 (N_43375,N_40867,N_40746);
nand U43376 (N_43376,N_41388,N_40610);
nand U43377 (N_43377,N_41996,N_40340);
or U43378 (N_43378,N_41111,N_40900);
nor U43379 (N_43379,N_41971,N_41584);
and U43380 (N_43380,N_41357,N_41178);
nor U43381 (N_43381,N_40439,N_40631);
or U43382 (N_43382,N_41113,N_41961);
and U43383 (N_43383,N_41773,N_41240);
nor U43384 (N_43384,N_41316,N_40091);
nor U43385 (N_43385,N_40679,N_41233);
and U43386 (N_43386,N_41471,N_40438);
or U43387 (N_43387,N_40981,N_41101);
xnor U43388 (N_43388,N_40407,N_40675);
or U43389 (N_43389,N_40763,N_41346);
xor U43390 (N_43390,N_41773,N_41274);
and U43391 (N_43391,N_41630,N_40218);
or U43392 (N_43392,N_41093,N_41462);
nor U43393 (N_43393,N_40349,N_40207);
nor U43394 (N_43394,N_41779,N_40080);
nor U43395 (N_43395,N_40172,N_40981);
nor U43396 (N_43396,N_41928,N_41902);
xor U43397 (N_43397,N_40142,N_40700);
nand U43398 (N_43398,N_41190,N_41862);
nor U43399 (N_43399,N_40299,N_40615);
nor U43400 (N_43400,N_40596,N_40025);
nor U43401 (N_43401,N_41905,N_41068);
and U43402 (N_43402,N_40011,N_40497);
xor U43403 (N_43403,N_40222,N_40184);
or U43404 (N_43404,N_41851,N_40434);
and U43405 (N_43405,N_40463,N_41526);
xnor U43406 (N_43406,N_41987,N_41185);
or U43407 (N_43407,N_41956,N_41320);
xor U43408 (N_43408,N_40317,N_40253);
xnor U43409 (N_43409,N_40703,N_40290);
xor U43410 (N_43410,N_41903,N_41614);
nor U43411 (N_43411,N_41993,N_41438);
nand U43412 (N_43412,N_41808,N_40417);
and U43413 (N_43413,N_40230,N_41767);
nor U43414 (N_43414,N_41216,N_40335);
nand U43415 (N_43415,N_41893,N_40746);
nand U43416 (N_43416,N_41276,N_41907);
and U43417 (N_43417,N_40467,N_40089);
or U43418 (N_43418,N_41135,N_40249);
xnor U43419 (N_43419,N_41957,N_41172);
nand U43420 (N_43420,N_41924,N_41989);
or U43421 (N_43421,N_40447,N_40351);
or U43422 (N_43422,N_41007,N_40459);
or U43423 (N_43423,N_40156,N_40827);
xor U43424 (N_43424,N_41948,N_40840);
or U43425 (N_43425,N_41659,N_40697);
nand U43426 (N_43426,N_41507,N_40209);
xor U43427 (N_43427,N_40121,N_41257);
nand U43428 (N_43428,N_40123,N_41241);
xnor U43429 (N_43429,N_41153,N_40133);
or U43430 (N_43430,N_41369,N_40427);
nand U43431 (N_43431,N_40153,N_41670);
xnor U43432 (N_43432,N_41190,N_41635);
or U43433 (N_43433,N_40667,N_41374);
nand U43434 (N_43434,N_40205,N_40367);
and U43435 (N_43435,N_40457,N_40693);
or U43436 (N_43436,N_40961,N_40278);
nor U43437 (N_43437,N_40206,N_40669);
and U43438 (N_43438,N_40291,N_41445);
nor U43439 (N_43439,N_41356,N_40946);
xnor U43440 (N_43440,N_40988,N_40233);
xor U43441 (N_43441,N_41901,N_41392);
or U43442 (N_43442,N_40302,N_41832);
nand U43443 (N_43443,N_41303,N_40514);
or U43444 (N_43444,N_41823,N_41391);
nand U43445 (N_43445,N_40309,N_40996);
xnor U43446 (N_43446,N_41132,N_40290);
or U43447 (N_43447,N_40176,N_41090);
xnor U43448 (N_43448,N_40372,N_41858);
xor U43449 (N_43449,N_41971,N_40528);
xnor U43450 (N_43450,N_41755,N_40443);
or U43451 (N_43451,N_40321,N_40484);
or U43452 (N_43452,N_41421,N_41511);
nand U43453 (N_43453,N_41762,N_40166);
or U43454 (N_43454,N_40276,N_40798);
and U43455 (N_43455,N_41321,N_41494);
nor U43456 (N_43456,N_41521,N_40578);
xor U43457 (N_43457,N_41361,N_40764);
nand U43458 (N_43458,N_40723,N_40110);
and U43459 (N_43459,N_41943,N_40242);
and U43460 (N_43460,N_41717,N_40304);
and U43461 (N_43461,N_41417,N_40749);
or U43462 (N_43462,N_41522,N_40576);
xnor U43463 (N_43463,N_40226,N_41344);
and U43464 (N_43464,N_41985,N_40239);
nand U43465 (N_43465,N_41214,N_40432);
xnor U43466 (N_43466,N_40256,N_41894);
xnor U43467 (N_43467,N_41543,N_41509);
xnor U43468 (N_43468,N_40830,N_41472);
and U43469 (N_43469,N_40833,N_40264);
or U43470 (N_43470,N_41300,N_40881);
or U43471 (N_43471,N_41789,N_40126);
nor U43472 (N_43472,N_41381,N_41360);
or U43473 (N_43473,N_41320,N_40518);
xor U43474 (N_43474,N_41460,N_41899);
or U43475 (N_43475,N_40152,N_40750);
or U43476 (N_43476,N_41478,N_40120);
and U43477 (N_43477,N_40454,N_40760);
nand U43478 (N_43478,N_40915,N_41373);
nor U43479 (N_43479,N_40640,N_41695);
nor U43480 (N_43480,N_41653,N_41890);
nor U43481 (N_43481,N_40359,N_41515);
xnor U43482 (N_43482,N_41387,N_41322);
nand U43483 (N_43483,N_41410,N_41093);
or U43484 (N_43484,N_41836,N_41547);
nor U43485 (N_43485,N_41489,N_40605);
or U43486 (N_43486,N_41305,N_41015);
or U43487 (N_43487,N_40339,N_41202);
and U43488 (N_43488,N_40826,N_41805);
nand U43489 (N_43489,N_40651,N_41200);
and U43490 (N_43490,N_41801,N_41907);
nand U43491 (N_43491,N_41896,N_40963);
and U43492 (N_43492,N_40416,N_41179);
and U43493 (N_43493,N_40219,N_40741);
nand U43494 (N_43494,N_41527,N_40880);
xor U43495 (N_43495,N_41072,N_40072);
nor U43496 (N_43496,N_41132,N_41200);
xnor U43497 (N_43497,N_40607,N_41244);
and U43498 (N_43498,N_40823,N_40822);
xnor U43499 (N_43499,N_41692,N_41491);
and U43500 (N_43500,N_40964,N_40609);
nor U43501 (N_43501,N_40621,N_41170);
and U43502 (N_43502,N_41774,N_41253);
and U43503 (N_43503,N_40604,N_41998);
nand U43504 (N_43504,N_40139,N_40082);
nand U43505 (N_43505,N_40084,N_41402);
or U43506 (N_43506,N_40497,N_41461);
and U43507 (N_43507,N_41639,N_41179);
nor U43508 (N_43508,N_41714,N_40570);
xnor U43509 (N_43509,N_40680,N_41438);
nand U43510 (N_43510,N_40391,N_40783);
and U43511 (N_43511,N_41124,N_41900);
or U43512 (N_43512,N_40093,N_40957);
nand U43513 (N_43513,N_40885,N_40688);
xnor U43514 (N_43514,N_40652,N_41939);
nand U43515 (N_43515,N_40244,N_41029);
nand U43516 (N_43516,N_40370,N_40388);
nor U43517 (N_43517,N_40464,N_40353);
or U43518 (N_43518,N_40403,N_40646);
nor U43519 (N_43519,N_41512,N_41630);
xnor U43520 (N_43520,N_40482,N_40004);
nand U43521 (N_43521,N_41309,N_40561);
nand U43522 (N_43522,N_41143,N_40633);
xor U43523 (N_43523,N_41627,N_40415);
nor U43524 (N_43524,N_41284,N_41526);
xor U43525 (N_43525,N_40930,N_40840);
nand U43526 (N_43526,N_41991,N_41284);
nand U43527 (N_43527,N_40926,N_40904);
or U43528 (N_43528,N_41576,N_41951);
nor U43529 (N_43529,N_40852,N_41019);
xnor U43530 (N_43530,N_40748,N_41962);
nand U43531 (N_43531,N_40590,N_41166);
nor U43532 (N_43532,N_41466,N_40982);
nand U43533 (N_43533,N_41966,N_41019);
nand U43534 (N_43534,N_41933,N_40265);
or U43535 (N_43535,N_40018,N_41653);
and U43536 (N_43536,N_40908,N_40069);
xnor U43537 (N_43537,N_40561,N_41850);
nand U43538 (N_43538,N_40337,N_41213);
and U43539 (N_43539,N_41930,N_41889);
nor U43540 (N_43540,N_40221,N_41642);
or U43541 (N_43541,N_41923,N_40431);
nor U43542 (N_43542,N_41091,N_40048);
and U43543 (N_43543,N_40330,N_40918);
xnor U43544 (N_43544,N_40337,N_41641);
or U43545 (N_43545,N_40623,N_41558);
nand U43546 (N_43546,N_41363,N_40265);
xor U43547 (N_43547,N_41125,N_41572);
or U43548 (N_43548,N_40765,N_40803);
and U43549 (N_43549,N_40900,N_41059);
and U43550 (N_43550,N_40061,N_41683);
nand U43551 (N_43551,N_40800,N_40143);
xor U43552 (N_43552,N_40712,N_41727);
nand U43553 (N_43553,N_41386,N_41137);
nand U43554 (N_43554,N_41059,N_40472);
nand U43555 (N_43555,N_41934,N_40135);
nand U43556 (N_43556,N_41713,N_41079);
and U43557 (N_43557,N_40684,N_40971);
xnor U43558 (N_43558,N_40629,N_41992);
xor U43559 (N_43559,N_40701,N_40784);
nand U43560 (N_43560,N_41630,N_40017);
and U43561 (N_43561,N_40498,N_41054);
nor U43562 (N_43562,N_40968,N_41884);
nand U43563 (N_43563,N_40471,N_41796);
and U43564 (N_43564,N_41506,N_41575);
or U43565 (N_43565,N_41033,N_40463);
nand U43566 (N_43566,N_40222,N_40424);
nor U43567 (N_43567,N_41160,N_41847);
xnor U43568 (N_43568,N_40817,N_41323);
xnor U43569 (N_43569,N_40166,N_41335);
and U43570 (N_43570,N_41558,N_40900);
nor U43571 (N_43571,N_41869,N_40411);
or U43572 (N_43572,N_40465,N_41535);
nor U43573 (N_43573,N_41697,N_41336);
or U43574 (N_43574,N_40082,N_40391);
nand U43575 (N_43575,N_40442,N_41264);
and U43576 (N_43576,N_40654,N_40325);
xnor U43577 (N_43577,N_41671,N_40562);
nor U43578 (N_43578,N_40669,N_40452);
or U43579 (N_43579,N_41088,N_41643);
or U43580 (N_43580,N_40699,N_40604);
and U43581 (N_43581,N_41712,N_41653);
nor U43582 (N_43582,N_40422,N_41371);
and U43583 (N_43583,N_41713,N_40855);
nand U43584 (N_43584,N_40153,N_40025);
or U43585 (N_43585,N_41662,N_41550);
and U43586 (N_43586,N_40778,N_40825);
or U43587 (N_43587,N_41465,N_41278);
xnor U43588 (N_43588,N_40234,N_40845);
nand U43589 (N_43589,N_40811,N_41497);
nand U43590 (N_43590,N_41722,N_41221);
and U43591 (N_43591,N_40719,N_40276);
xnor U43592 (N_43592,N_40466,N_40123);
xor U43593 (N_43593,N_41682,N_41219);
and U43594 (N_43594,N_41451,N_41111);
nor U43595 (N_43595,N_41572,N_41197);
xnor U43596 (N_43596,N_41995,N_41303);
nand U43597 (N_43597,N_41613,N_40513);
or U43598 (N_43598,N_40209,N_40691);
xnor U43599 (N_43599,N_41200,N_41609);
xor U43600 (N_43600,N_41766,N_41544);
nand U43601 (N_43601,N_40220,N_40326);
nand U43602 (N_43602,N_40971,N_40911);
nand U43603 (N_43603,N_40909,N_40729);
nor U43604 (N_43604,N_40253,N_41873);
or U43605 (N_43605,N_41951,N_41072);
nor U43606 (N_43606,N_40153,N_41058);
or U43607 (N_43607,N_41987,N_41082);
nand U43608 (N_43608,N_40427,N_40304);
nand U43609 (N_43609,N_40601,N_40805);
nand U43610 (N_43610,N_40582,N_41393);
or U43611 (N_43611,N_41004,N_41810);
xnor U43612 (N_43612,N_41748,N_40430);
and U43613 (N_43613,N_40480,N_40332);
and U43614 (N_43614,N_40621,N_41495);
xor U43615 (N_43615,N_40817,N_40848);
nand U43616 (N_43616,N_40119,N_40848);
and U43617 (N_43617,N_40499,N_41284);
nand U43618 (N_43618,N_41570,N_40571);
or U43619 (N_43619,N_40407,N_40102);
and U43620 (N_43620,N_40160,N_40999);
xor U43621 (N_43621,N_40531,N_40311);
or U43622 (N_43622,N_40808,N_40415);
or U43623 (N_43623,N_41446,N_41565);
nor U43624 (N_43624,N_40534,N_41078);
xor U43625 (N_43625,N_41185,N_41658);
or U43626 (N_43626,N_40502,N_40680);
nand U43627 (N_43627,N_40357,N_41827);
xor U43628 (N_43628,N_41971,N_41574);
xor U43629 (N_43629,N_41153,N_40611);
or U43630 (N_43630,N_40757,N_41577);
and U43631 (N_43631,N_41917,N_40133);
nand U43632 (N_43632,N_41722,N_40508);
and U43633 (N_43633,N_40756,N_40153);
or U43634 (N_43634,N_40901,N_40743);
xor U43635 (N_43635,N_41286,N_40615);
nor U43636 (N_43636,N_41162,N_40301);
nand U43637 (N_43637,N_41956,N_40243);
xnor U43638 (N_43638,N_41434,N_40315);
or U43639 (N_43639,N_41544,N_41035);
nand U43640 (N_43640,N_40530,N_40256);
nand U43641 (N_43641,N_41460,N_41820);
nor U43642 (N_43642,N_41682,N_40211);
xnor U43643 (N_43643,N_40787,N_41926);
or U43644 (N_43644,N_41427,N_40736);
or U43645 (N_43645,N_40828,N_41397);
nor U43646 (N_43646,N_40224,N_41989);
nand U43647 (N_43647,N_41651,N_41711);
xor U43648 (N_43648,N_40016,N_41633);
nor U43649 (N_43649,N_40345,N_40121);
xnor U43650 (N_43650,N_40520,N_40154);
nor U43651 (N_43651,N_40520,N_40930);
or U43652 (N_43652,N_41527,N_40716);
nand U43653 (N_43653,N_40104,N_41177);
nor U43654 (N_43654,N_41140,N_40217);
and U43655 (N_43655,N_41185,N_40200);
and U43656 (N_43656,N_41375,N_41736);
or U43657 (N_43657,N_40425,N_40063);
xnor U43658 (N_43658,N_41283,N_41922);
and U43659 (N_43659,N_40294,N_40403);
or U43660 (N_43660,N_41154,N_40225);
and U43661 (N_43661,N_41202,N_41987);
xnor U43662 (N_43662,N_41687,N_41998);
nor U43663 (N_43663,N_40581,N_40774);
and U43664 (N_43664,N_41100,N_41430);
xnor U43665 (N_43665,N_40079,N_40920);
or U43666 (N_43666,N_40965,N_40980);
nor U43667 (N_43667,N_40277,N_40115);
and U43668 (N_43668,N_41359,N_41172);
and U43669 (N_43669,N_41344,N_41701);
and U43670 (N_43670,N_40724,N_41415);
and U43671 (N_43671,N_41768,N_40669);
and U43672 (N_43672,N_40159,N_41731);
nor U43673 (N_43673,N_41838,N_41097);
and U43674 (N_43674,N_41968,N_40125);
or U43675 (N_43675,N_41131,N_41946);
nor U43676 (N_43676,N_41719,N_41303);
nor U43677 (N_43677,N_41719,N_41015);
or U43678 (N_43678,N_41112,N_40183);
nor U43679 (N_43679,N_41869,N_40959);
nand U43680 (N_43680,N_41588,N_40165);
or U43681 (N_43681,N_40788,N_41728);
nor U43682 (N_43682,N_40191,N_41625);
or U43683 (N_43683,N_40395,N_40305);
and U43684 (N_43684,N_40802,N_41195);
nor U43685 (N_43685,N_40130,N_41121);
nand U43686 (N_43686,N_41033,N_40430);
or U43687 (N_43687,N_41790,N_40087);
xnor U43688 (N_43688,N_41925,N_41968);
nand U43689 (N_43689,N_40390,N_41675);
or U43690 (N_43690,N_40608,N_40820);
nand U43691 (N_43691,N_41683,N_41213);
nand U43692 (N_43692,N_40817,N_41697);
or U43693 (N_43693,N_40715,N_40568);
nand U43694 (N_43694,N_40176,N_41767);
and U43695 (N_43695,N_40148,N_40726);
and U43696 (N_43696,N_41168,N_40313);
nor U43697 (N_43697,N_40159,N_40300);
or U43698 (N_43698,N_40710,N_40737);
and U43699 (N_43699,N_41263,N_41287);
nand U43700 (N_43700,N_41789,N_41874);
xnor U43701 (N_43701,N_40168,N_41605);
or U43702 (N_43702,N_40333,N_41405);
xnor U43703 (N_43703,N_41490,N_41148);
and U43704 (N_43704,N_41330,N_41195);
xor U43705 (N_43705,N_40904,N_40185);
or U43706 (N_43706,N_41459,N_41489);
nand U43707 (N_43707,N_40911,N_41597);
or U43708 (N_43708,N_40462,N_41440);
or U43709 (N_43709,N_40709,N_41828);
or U43710 (N_43710,N_40298,N_41111);
nand U43711 (N_43711,N_40829,N_41494);
nand U43712 (N_43712,N_41892,N_41894);
xnor U43713 (N_43713,N_40911,N_41499);
nand U43714 (N_43714,N_41436,N_41726);
and U43715 (N_43715,N_41092,N_40186);
xnor U43716 (N_43716,N_41290,N_41100);
xnor U43717 (N_43717,N_41235,N_40205);
or U43718 (N_43718,N_40421,N_41723);
nor U43719 (N_43719,N_40452,N_40591);
nor U43720 (N_43720,N_40433,N_40603);
and U43721 (N_43721,N_41487,N_41318);
nand U43722 (N_43722,N_40568,N_41126);
nor U43723 (N_43723,N_40866,N_41319);
xor U43724 (N_43724,N_41124,N_40366);
and U43725 (N_43725,N_40939,N_41589);
nor U43726 (N_43726,N_40708,N_40763);
or U43727 (N_43727,N_41981,N_40550);
nand U43728 (N_43728,N_40899,N_41118);
and U43729 (N_43729,N_41781,N_41847);
and U43730 (N_43730,N_40417,N_41573);
nor U43731 (N_43731,N_41308,N_41604);
and U43732 (N_43732,N_40911,N_40312);
or U43733 (N_43733,N_40895,N_40673);
nor U43734 (N_43734,N_40947,N_41834);
nor U43735 (N_43735,N_41437,N_40991);
nor U43736 (N_43736,N_41116,N_41248);
nor U43737 (N_43737,N_40002,N_41773);
nor U43738 (N_43738,N_41672,N_41639);
xnor U43739 (N_43739,N_40023,N_40737);
nor U43740 (N_43740,N_40439,N_41361);
nand U43741 (N_43741,N_40108,N_40064);
nor U43742 (N_43742,N_41964,N_40146);
xor U43743 (N_43743,N_41456,N_40721);
or U43744 (N_43744,N_41877,N_40665);
or U43745 (N_43745,N_40359,N_40065);
xor U43746 (N_43746,N_41034,N_41163);
xnor U43747 (N_43747,N_41082,N_41580);
xnor U43748 (N_43748,N_40695,N_41051);
or U43749 (N_43749,N_40635,N_40913);
nand U43750 (N_43750,N_41568,N_40251);
or U43751 (N_43751,N_40815,N_41066);
and U43752 (N_43752,N_41704,N_41751);
nor U43753 (N_43753,N_41549,N_41236);
nor U43754 (N_43754,N_40898,N_40824);
nand U43755 (N_43755,N_40565,N_40252);
and U43756 (N_43756,N_40663,N_40283);
nand U43757 (N_43757,N_40596,N_40394);
xor U43758 (N_43758,N_40664,N_41455);
xor U43759 (N_43759,N_40823,N_40650);
or U43760 (N_43760,N_41191,N_41846);
and U43761 (N_43761,N_40323,N_41737);
or U43762 (N_43762,N_40185,N_40544);
nor U43763 (N_43763,N_40011,N_40247);
nand U43764 (N_43764,N_40521,N_40064);
xor U43765 (N_43765,N_40335,N_41618);
xor U43766 (N_43766,N_41265,N_41323);
nor U43767 (N_43767,N_41383,N_41173);
or U43768 (N_43768,N_40742,N_41062);
nor U43769 (N_43769,N_41379,N_40631);
nand U43770 (N_43770,N_40542,N_40710);
nand U43771 (N_43771,N_40743,N_41075);
xnor U43772 (N_43772,N_41828,N_40364);
and U43773 (N_43773,N_40806,N_41131);
xor U43774 (N_43774,N_40521,N_41682);
nand U43775 (N_43775,N_40270,N_40156);
and U43776 (N_43776,N_41177,N_41223);
xnor U43777 (N_43777,N_40411,N_41369);
and U43778 (N_43778,N_40380,N_41182);
and U43779 (N_43779,N_40049,N_41360);
xnor U43780 (N_43780,N_41418,N_41864);
nor U43781 (N_43781,N_40892,N_40239);
nor U43782 (N_43782,N_40722,N_41016);
and U43783 (N_43783,N_41222,N_41104);
and U43784 (N_43784,N_41359,N_40046);
nor U43785 (N_43785,N_41588,N_40491);
or U43786 (N_43786,N_40034,N_40302);
or U43787 (N_43787,N_40790,N_41761);
xnor U43788 (N_43788,N_41928,N_41392);
nor U43789 (N_43789,N_41017,N_40030);
nand U43790 (N_43790,N_40524,N_41312);
or U43791 (N_43791,N_41542,N_40872);
or U43792 (N_43792,N_40694,N_40033);
nor U43793 (N_43793,N_41398,N_41737);
nor U43794 (N_43794,N_41282,N_41400);
and U43795 (N_43795,N_40880,N_41862);
and U43796 (N_43796,N_40000,N_40929);
and U43797 (N_43797,N_40179,N_40197);
xor U43798 (N_43798,N_41688,N_41660);
xor U43799 (N_43799,N_40430,N_41631);
nand U43800 (N_43800,N_40929,N_41445);
nor U43801 (N_43801,N_41776,N_41771);
nor U43802 (N_43802,N_40641,N_40929);
nand U43803 (N_43803,N_40867,N_41018);
nor U43804 (N_43804,N_40936,N_41416);
nor U43805 (N_43805,N_41128,N_40368);
nand U43806 (N_43806,N_40731,N_40298);
nor U43807 (N_43807,N_41893,N_41604);
and U43808 (N_43808,N_40474,N_40187);
nor U43809 (N_43809,N_41702,N_40644);
xnor U43810 (N_43810,N_41525,N_40785);
nor U43811 (N_43811,N_40759,N_41967);
nor U43812 (N_43812,N_41542,N_41536);
xor U43813 (N_43813,N_40319,N_41631);
xnor U43814 (N_43814,N_41652,N_40851);
and U43815 (N_43815,N_41129,N_41418);
xnor U43816 (N_43816,N_41583,N_40867);
nor U43817 (N_43817,N_41373,N_41005);
nand U43818 (N_43818,N_40591,N_41383);
or U43819 (N_43819,N_40610,N_41490);
xor U43820 (N_43820,N_41728,N_41256);
or U43821 (N_43821,N_40233,N_41335);
and U43822 (N_43822,N_40010,N_40326);
nor U43823 (N_43823,N_41317,N_41281);
xor U43824 (N_43824,N_40216,N_41507);
nand U43825 (N_43825,N_41006,N_41038);
nor U43826 (N_43826,N_41716,N_41537);
nand U43827 (N_43827,N_41172,N_41808);
nand U43828 (N_43828,N_40344,N_41917);
and U43829 (N_43829,N_40088,N_40098);
or U43830 (N_43830,N_40174,N_40217);
nand U43831 (N_43831,N_41798,N_40309);
and U43832 (N_43832,N_41902,N_40305);
nand U43833 (N_43833,N_40663,N_40710);
xnor U43834 (N_43834,N_40472,N_40495);
nand U43835 (N_43835,N_40489,N_40110);
or U43836 (N_43836,N_41313,N_40480);
and U43837 (N_43837,N_41837,N_40456);
or U43838 (N_43838,N_41637,N_41830);
nand U43839 (N_43839,N_40551,N_41943);
xor U43840 (N_43840,N_40737,N_40563);
xnor U43841 (N_43841,N_41171,N_41905);
xnor U43842 (N_43842,N_41092,N_40273);
nor U43843 (N_43843,N_41388,N_41765);
nand U43844 (N_43844,N_41037,N_41305);
nor U43845 (N_43845,N_40544,N_41830);
xnor U43846 (N_43846,N_41244,N_40154);
or U43847 (N_43847,N_41754,N_41393);
nand U43848 (N_43848,N_40707,N_40312);
nor U43849 (N_43849,N_40981,N_41629);
xor U43850 (N_43850,N_41003,N_41363);
nand U43851 (N_43851,N_41496,N_41699);
xnor U43852 (N_43852,N_41242,N_41370);
or U43853 (N_43853,N_40538,N_41973);
nand U43854 (N_43854,N_41259,N_41984);
xnor U43855 (N_43855,N_41240,N_40706);
nand U43856 (N_43856,N_40861,N_41522);
or U43857 (N_43857,N_41407,N_40958);
nor U43858 (N_43858,N_40818,N_40883);
or U43859 (N_43859,N_40892,N_40175);
xor U43860 (N_43860,N_40887,N_40863);
xor U43861 (N_43861,N_41307,N_41144);
and U43862 (N_43862,N_41010,N_40610);
nand U43863 (N_43863,N_41465,N_40785);
xor U43864 (N_43864,N_41565,N_40230);
nand U43865 (N_43865,N_40035,N_40676);
nor U43866 (N_43866,N_40750,N_40699);
or U43867 (N_43867,N_41729,N_40572);
and U43868 (N_43868,N_41119,N_40049);
nand U43869 (N_43869,N_40087,N_41509);
xor U43870 (N_43870,N_41579,N_41966);
nor U43871 (N_43871,N_40985,N_41573);
and U43872 (N_43872,N_40735,N_40764);
nand U43873 (N_43873,N_40815,N_41064);
xnor U43874 (N_43874,N_41870,N_41439);
nor U43875 (N_43875,N_41940,N_41546);
nor U43876 (N_43876,N_41758,N_40480);
or U43877 (N_43877,N_41650,N_40179);
nand U43878 (N_43878,N_41360,N_41250);
or U43879 (N_43879,N_40184,N_41147);
nand U43880 (N_43880,N_40246,N_40601);
or U43881 (N_43881,N_40546,N_40492);
or U43882 (N_43882,N_41756,N_40454);
nor U43883 (N_43883,N_41996,N_40225);
and U43884 (N_43884,N_41545,N_41720);
nor U43885 (N_43885,N_40766,N_41100);
and U43886 (N_43886,N_41791,N_40768);
and U43887 (N_43887,N_40542,N_41369);
and U43888 (N_43888,N_41624,N_41916);
or U43889 (N_43889,N_40474,N_41244);
or U43890 (N_43890,N_41902,N_40074);
and U43891 (N_43891,N_41573,N_40076);
nor U43892 (N_43892,N_41063,N_40092);
nand U43893 (N_43893,N_41535,N_41517);
and U43894 (N_43894,N_40761,N_41247);
nand U43895 (N_43895,N_41973,N_40008);
and U43896 (N_43896,N_40308,N_41024);
and U43897 (N_43897,N_40808,N_41946);
or U43898 (N_43898,N_40877,N_40032);
nand U43899 (N_43899,N_40499,N_41947);
or U43900 (N_43900,N_41728,N_40546);
nor U43901 (N_43901,N_41385,N_40926);
nor U43902 (N_43902,N_40402,N_40938);
or U43903 (N_43903,N_40238,N_41524);
or U43904 (N_43904,N_41389,N_41429);
nand U43905 (N_43905,N_40899,N_41413);
xor U43906 (N_43906,N_41491,N_41575);
or U43907 (N_43907,N_41461,N_40520);
nand U43908 (N_43908,N_40322,N_40567);
nor U43909 (N_43909,N_41233,N_40712);
or U43910 (N_43910,N_40896,N_41936);
or U43911 (N_43911,N_41615,N_40357);
or U43912 (N_43912,N_41777,N_41923);
xor U43913 (N_43913,N_40054,N_41748);
nand U43914 (N_43914,N_41066,N_40779);
nor U43915 (N_43915,N_40710,N_40525);
xor U43916 (N_43916,N_40900,N_41373);
nand U43917 (N_43917,N_40875,N_41091);
nor U43918 (N_43918,N_40180,N_41705);
or U43919 (N_43919,N_40472,N_40019);
or U43920 (N_43920,N_41849,N_40746);
xor U43921 (N_43921,N_40608,N_40804);
nor U43922 (N_43922,N_40874,N_40179);
or U43923 (N_43923,N_41111,N_40921);
or U43924 (N_43924,N_40560,N_40490);
and U43925 (N_43925,N_41748,N_40730);
or U43926 (N_43926,N_40019,N_41675);
xnor U43927 (N_43927,N_41415,N_41673);
nor U43928 (N_43928,N_40244,N_41642);
xnor U43929 (N_43929,N_40934,N_40116);
xor U43930 (N_43930,N_41240,N_41879);
and U43931 (N_43931,N_41451,N_40109);
nor U43932 (N_43932,N_40319,N_41700);
xnor U43933 (N_43933,N_41179,N_40100);
nor U43934 (N_43934,N_41508,N_41017);
xnor U43935 (N_43935,N_40340,N_40008);
nor U43936 (N_43936,N_40960,N_41178);
nand U43937 (N_43937,N_41597,N_40336);
or U43938 (N_43938,N_41721,N_40278);
and U43939 (N_43939,N_41461,N_41803);
xor U43940 (N_43940,N_41056,N_41180);
and U43941 (N_43941,N_41741,N_40762);
and U43942 (N_43942,N_40649,N_41823);
nand U43943 (N_43943,N_40960,N_41264);
or U43944 (N_43944,N_40530,N_40646);
or U43945 (N_43945,N_41231,N_41945);
xor U43946 (N_43946,N_41271,N_40850);
xnor U43947 (N_43947,N_40622,N_40072);
or U43948 (N_43948,N_40546,N_41365);
or U43949 (N_43949,N_40486,N_41349);
nor U43950 (N_43950,N_41989,N_41970);
nand U43951 (N_43951,N_41665,N_41723);
xor U43952 (N_43952,N_41193,N_40638);
and U43953 (N_43953,N_40272,N_40654);
xor U43954 (N_43954,N_41025,N_40628);
and U43955 (N_43955,N_40608,N_40254);
nor U43956 (N_43956,N_40807,N_40875);
and U43957 (N_43957,N_41863,N_40658);
xor U43958 (N_43958,N_40392,N_41660);
xor U43959 (N_43959,N_40578,N_40848);
or U43960 (N_43960,N_41465,N_41039);
or U43961 (N_43961,N_41364,N_40145);
xor U43962 (N_43962,N_41142,N_41925);
nor U43963 (N_43963,N_40199,N_41612);
xnor U43964 (N_43964,N_41076,N_40606);
and U43965 (N_43965,N_41061,N_41418);
or U43966 (N_43966,N_41819,N_40883);
nand U43967 (N_43967,N_41500,N_40997);
nand U43968 (N_43968,N_40158,N_40925);
xor U43969 (N_43969,N_41110,N_40417);
xor U43970 (N_43970,N_41676,N_40575);
nor U43971 (N_43971,N_40622,N_40287);
and U43972 (N_43972,N_40754,N_40447);
or U43973 (N_43973,N_40360,N_40442);
or U43974 (N_43974,N_40701,N_40406);
and U43975 (N_43975,N_41042,N_40015);
xor U43976 (N_43976,N_41926,N_40912);
and U43977 (N_43977,N_40818,N_41980);
and U43978 (N_43978,N_41808,N_41771);
or U43979 (N_43979,N_40659,N_40585);
and U43980 (N_43980,N_40020,N_41256);
and U43981 (N_43981,N_40087,N_41096);
or U43982 (N_43982,N_41150,N_41322);
xor U43983 (N_43983,N_40426,N_40060);
or U43984 (N_43984,N_40148,N_41390);
xor U43985 (N_43985,N_41099,N_40973);
or U43986 (N_43986,N_40629,N_40930);
and U43987 (N_43987,N_40688,N_40039);
nand U43988 (N_43988,N_41065,N_40245);
or U43989 (N_43989,N_40400,N_40973);
xnor U43990 (N_43990,N_41457,N_41097);
nand U43991 (N_43991,N_40189,N_41733);
or U43992 (N_43992,N_40623,N_41442);
xnor U43993 (N_43993,N_41799,N_40542);
and U43994 (N_43994,N_41404,N_40755);
nand U43995 (N_43995,N_40412,N_41147);
nand U43996 (N_43996,N_41705,N_41314);
xor U43997 (N_43997,N_41843,N_41135);
nand U43998 (N_43998,N_41588,N_41762);
or U43999 (N_43999,N_41111,N_41266);
and U44000 (N_44000,N_43467,N_42227);
or U44001 (N_44001,N_43295,N_43749);
or U44002 (N_44002,N_42016,N_43704);
nand U44003 (N_44003,N_42176,N_43552);
xor U44004 (N_44004,N_43586,N_43409);
nor U44005 (N_44005,N_43419,N_43659);
nor U44006 (N_44006,N_42054,N_43224);
nor U44007 (N_44007,N_42421,N_43183);
and U44008 (N_44008,N_43046,N_42984);
xnor U44009 (N_44009,N_43605,N_42246);
or U44010 (N_44010,N_43466,N_42501);
xnor U44011 (N_44011,N_43114,N_43455);
xor U44012 (N_44012,N_42602,N_43314);
or U44013 (N_44013,N_43221,N_43100);
xnor U44014 (N_44014,N_42353,N_42218);
nor U44015 (N_44015,N_42035,N_42747);
xnor U44016 (N_44016,N_42783,N_42005);
xnor U44017 (N_44017,N_43672,N_43345);
or U44018 (N_44018,N_43778,N_43824);
or U44019 (N_44019,N_43177,N_43410);
and U44020 (N_44020,N_42997,N_42053);
xnor U44021 (N_44021,N_42132,N_42752);
nand U44022 (N_44022,N_43272,N_43601);
or U44023 (N_44023,N_43059,N_43000);
xnor U44024 (N_44024,N_42994,N_43976);
and U44025 (N_44025,N_42812,N_43544);
and U44026 (N_44026,N_43781,N_42210);
xnor U44027 (N_44027,N_42037,N_43225);
and U44028 (N_44028,N_43716,N_43539);
or U44029 (N_44029,N_43408,N_42743);
xnor U44030 (N_44030,N_43149,N_43031);
nand U44031 (N_44031,N_43835,N_43473);
or U44032 (N_44032,N_42120,N_42420);
nor U44033 (N_44033,N_43840,N_43442);
and U44034 (N_44034,N_43500,N_42799);
xor U44035 (N_44035,N_42043,N_42418);
xor U44036 (N_44036,N_42378,N_43958);
and U44037 (N_44037,N_43512,N_42635);
xnor U44038 (N_44038,N_42536,N_42958);
or U44039 (N_44039,N_43872,N_43548);
xor U44040 (N_44040,N_42284,N_42440);
and U44041 (N_44041,N_43596,N_43988);
or U44042 (N_44042,N_42446,N_42433);
and U44043 (N_44043,N_42560,N_42822);
nand U44044 (N_44044,N_43766,N_42065);
nand U44045 (N_44045,N_43517,N_43187);
and U44046 (N_44046,N_42249,N_42983);
nor U44047 (N_44047,N_43330,N_42028);
nand U44048 (N_44048,N_43759,N_42715);
xnor U44049 (N_44049,N_43549,N_43399);
nand U44050 (N_44050,N_42578,N_42322);
or U44051 (N_44051,N_42214,N_43068);
or U44052 (N_44052,N_42186,N_43588);
or U44053 (N_44053,N_42612,N_42962);
nand U44054 (N_44054,N_42463,N_43757);
nor U44055 (N_44055,N_43634,N_43179);
or U44056 (N_44056,N_43867,N_43392);
nor U44057 (N_44057,N_43579,N_43497);
and U44058 (N_44058,N_43746,N_42671);
nand U44059 (N_44059,N_42466,N_43487);
or U44060 (N_44060,N_43034,N_43266);
nand U44061 (N_44061,N_42432,N_43947);
nor U44062 (N_44062,N_42202,N_43087);
nand U44063 (N_44063,N_43133,N_43412);
nand U44064 (N_44064,N_43141,N_42948);
and U44065 (N_44065,N_42335,N_43411);
nand U44066 (N_44066,N_43439,N_43057);
nand U44067 (N_44067,N_42328,N_43858);
and U44068 (N_44068,N_42540,N_43656);
and U44069 (N_44069,N_43420,N_43082);
and U44070 (N_44070,N_43815,N_42113);
or U44071 (N_44071,N_42185,N_42661);
nor U44072 (N_44072,N_42516,N_43361);
xor U44073 (N_44073,N_43931,N_43318);
xor U44074 (N_44074,N_42472,N_43564);
nor U44075 (N_44075,N_42724,N_42911);
nand U44076 (N_44076,N_43001,N_43673);
xor U44077 (N_44077,N_42490,N_43014);
or U44078 (N_44078,N_43274,N_43735);
nand U44079 (N_44079,N_42075,N_43845);
nand U44080 (N_44080,N_42541,N_42175);
xor U44081 (N_44081,N_43256,N_43465);
nor U44082 (N_44082,N_42254,N_43366);
or U44083 (N_44083,N_43677,N_43485);
nor U44084 (N_44084,N_42144,N_42801);
nor U44085 (N_44085,N_42641,N_43075);
or U44086 (N_44086,N_43647,N_42637);
or U44087 (N_44087,N_43774,N_43829);
xnor U44088 (N_44088,N_42355,N_42127);
xnor U44089 (N_44089,N_43414,N_42826);
nand U44090 (N_44090,N_42792,N_42359);
and U44091 (N_44091,N_43237,N_42723);
xnor U44092 (N_44092,N_42347,N_43120);
nand U44093 (N_44093,N_42033,N_42609);
nor U44094 (N_44094,N_43316,N_42905);
xor U44095 (N_44095,N_42384,N_43956);
and U44096 (N_44096,N_42673,N_42924);
or U44097 (N_44097,N_42036,N_43250);
nand U44098 (N_44098,N_42481,N_42684);
xor U44099 (N_44099,N_43033,N_42205);
or U44100 (N_44100,N_43503,N_42230);
and U44101 (N_44101,N_43226,N_43271);
xor U44102 (N_44102,N_42183,N_43418);
and U44103 (N_44103,N_42416,N_43032);
or U44104 (N_44104,N_43709,N_42913);
nand U44105 (N_44105,N_43162,N_42872);
xnor U44106 (N_44106,N_43425,N_43532);
nor U44107 (N_44107,N_43721,N_43923);
xnor U44108 (N_44108,N_43373,N_42790);
nor U44109 (N_44109,N_42173,N_42662);
xor U44110 (N_44110,N_42296,N_42226);
nand U44111 (N_44111,N_42094,N_43152);
and U44112 (N_44112,N_43488,N_42059);
nor U44113 (N_44113,N_42004,N_43665);
nor U44114 (N_44114,N_43343,N_42425);
and U44115 (N_44115,N_42130,N_42804);
nor U44116 (N_44116,N_43834,N_42553);
and U44117 (N_44117,N_42999,N_42566);
nor U44118 (N_44118,N_43195,N_43435);
xor U44119 (N_44119,N_42055,N_42643);
xor U44120 (N_44120,N_42060,N_43383);
and U44121 (N_44121,N_43168,N_43572);
xnor U44122 (N_44122,N_43388,N_43763);
nand U44123 (N_44123,N_43519,N_43798);
nor U44124 (N_44124,N_42403,N_42846);
nor U44125 (N_44125,N_42166,N_43949);
xnor U44126 (N_44126,N_42182,N_42753);
xor U44127 (N_44127,N_43110,N_43955);
and U44128 (N_44128,N_42502,N_42413);
xnor U44129 (N_44129,N_42039,N_42896);
and U44130 (N_44130,N_43328,N_43851);
nor U44131 (N_44131,N_42165,N_43844);
xor U44132 (N_44132,N_43338,N_43401);
nand U44133 (N_44133,N_42557,N_42112);
xnor U44134 (N_44134,N_43627,N_43422);
xnor U44135 (N_44135,N_42306,N_42442);
nand U44136 (N_44136,N_43275,N_42672);
xor U44137 (N_44137,N_43102,N_42504);
and U44138 (N_44138,N_43458,N_43535);
xor U44139 (N_44139,N_42239,N_43148);
nor U44140 (N_44140,N_43406,N_42996);
and U44141 (N_44141,N_42253,N_42260);
nand U44142 (N_44142,N_42800,N_43067);
xnor U44143 (N_44143,N_42122,N_43350);
xor U44144 (N_44144,N_42711,N_43946);
or U44145 (N_44145,N_42492,N_42595);
nand U44146 (N_44146,N_43784,N_42029);
or U44147 (N_44147,N_42302,N_42926);
xor U44148 (N_44148,N_43352,N_42273);
nor U44149 (N_44149,N_42966,N_43918);
or U44150 (N_44150,N_43702,N_43642);
and U44151 (N_44151,N_43699,N_42589);
or U44152 (N_44152,N_43003,N_42052);
nand U44153 (N_44153,N_43807,N_42380);
nand U44154 (N_44154,N_43636,N_42277);
or U44155 (N_44155,N_43813,N_43556);
or U44156 (N_44156,N_43289,N_42939);
or U44157 (N_44157,N_43600,N_42476);
and U44158 (N_44158,N_43966,N_43922);
and U44159 (N_44159,N_42096,N_42545);
or U44160 (N_44160,N_43996,N_43842);
or U44161 (N_44161,N_43850,N_43079);
and U44162 (N_44162,N_43028,N_43896);
xor U44163 (N_44163,N_43492,N_43066);
nor U44164 (N_44164,N_42168,N_42579);
nor U44165 (N_44165,N_43712,N_43360);
or U44166 (N_44166,N_42320,N_42487);
nand U44167 (N_44167,N_42204,N_43443);
and U44168 (N_44168,N_42430,N_43002);
nor U44169 (N_44169,N_42586,N_43142);
and U44170 (N_44170,N_43528,N_43459);
nand U44171 (N_44171,N_43899,N_42402);
nand U44172 (N_44172,N_42041,N_42484);
nor U44173 (N_44173,N_42934,N_43260);
nor U44174 (N_44174,N_42843,N_42827);
nand U44175 (N_44175,N_42217,N_43501);
nor U44176 (N_44176,N_42660,N_43597);
nor U44177 (N_44177,N_42293,N_42895);
nand U44178 (N_44178,N_43264,N_42678);
nor U44179 (N_44179,N_42953,N_43733);
and U44180 (N_44180,N_42746,N_43630);
nand U44181 (N_44181,N_42759,N_43523);
or U44182 (N_44182,N_42577,N_42704);
and U44183 (N_44183,N_43104,N_42462);
and U44184 (N_44184,N_42606,N_42977);
and U44185 (N_44185,N_42073,N_42960);
xor U44186 (N_44186,N_42232,N_43232);
and U44187 (N_44187,N_43444,N_42633);
nor U44188 (N_44188,N_42990,N_43341);
xnor U44189 (N_44189,N_42344,N_43827);
xor U44190 (N_44190,N_42103,N_43276);
xor U44191 (N_44191,N_43995,N_43773);
and U44192 (N_44192,N_43667,N_43510);
nand U44193 (N_44193,N_42884,N_43038);
or U44194 (N_44194,N_42118,N_43215);
nand U44195 (N_44195,N_43959,N_42568);
or U44196 (N_44196,N_42923,N_43036);
nor U44197 (N_44197,N_42066,N_43337);
nand U44198 (N_44198,N_43287,N_42729);
nor U44199 (N_44199,N_42315,N_42495);
and U44200 (N_44200,N_42388,N_43629);
or U44201 (N_44201,N_42508,N_42365);
nand U44202 (N_44202,N_42791,N_43894);
nor U44203 (N_44203,N_42313,N_43595);
xnor U44204 (N_44204,N_43270,N_43646);
nand U44205 (N_44205,N_43843,N_42238);
xnor U44206 (N_44206,N_42292,N_43201);
nor U44207 (N_44207,N_42959,N_42093);
and U44208 (N_44208,N_43008,N_42698);
or U44209 (N_44209,N_42841,N_43365);
nand U44210 (N_44210,N_42377,N_43904);
nor U44211 (N_44211,N_43675,N_42649);
nor U44212 (N_44212,N_43053,N_43967);
xnor U44213 (N_44213,N_42610,N_43219);
or U44214 (N_44214,N_43056,N_43372);
nand U44215 (N_44215,N_42592,N_43864);
xnor U44216 (N_44216,N_43099,N_42778);
or U44217 (N_44217,N_43805,N_42625);
nand U44218 (N_44218,N_43891,N_42019);
nor U44219 (N_44219,N_43080,N_43371);
nand U44220 (N_44220,N_43151,N_42584);
nand U44221 (N_44221,N_42162,N_42447);
and U44222 (N_44222,N_43358,N_43578);
nand U44223 (N_44223,N_42471,N_43426);
and U44224 (N_44224,N_42648,N_43189);
nor U44225 (N_44225,N_42349,N_43892);
nand U44226 (N_44226,N_42235,N_43823);
xor U44227 (N_44227,N_43332,N_43755);
xor U44228 (N_44228,N_42668,N_42814);
or U44229 (N_44229,N_43668,N_43283);
xnor U44230 (N_44230,N_43878,N_43292);
xor U44231 (N_44231,N_42617,N_42098);
or U44232 (N_44232,N_43153,N_42395);
nor U44233 (N_44233,N_42844,N_42564);
or U44234 (N_44234,N_42786,N_43602);
or U44235 (N_44235,N_42255,N_42770);
and U44236 (N_44236,N_42963,N_43170);
nand U44237 (N_44237,N_43980,N_43527);
or U44238 (N_44238,N_42299,N_42308);
nand U44239 (N_44239,N_42158,N_42642);
or U44240 (N_44240,N_42247,N_42138);
or U44241 (N_44241,N_43689,N_42242);
nor U44242 (N_44242,N_42782,N_43690);
xnor U44243 (N_44243,N_43395,N_42156);
or U44244 (N_44244,N_42892,N_43553);
nor U44245 (N_44245,N_43971,N_43954);
and U44246 (N_44246,N_42062,N_42412);
nor U44247 (N_44247,N_43562,N_42265);
or U44248 (N_44248,N_42636,N_42494);
or U44249 (N_44249,N_42269,N_42017);
or U44250 (N_44250,N_42032,N_43883);
nor U44251 (N_44251,N_42988,N_42219);
and U44252 (N_44252,N_42531,N_42789);
or U44253 (N_44253,N_42864,N_43180);
xnor U44254 (N_44254,N_43960,N_42979);
nor U44255 (N_44255,N_42554,N_42739);
xor U44256 (N_44256,N_42220,N_43545);
nand U44257 (N_44257,N_42187,N_43163);
nand U44258 (N_44258,N_42954,N_43612);
or U44259 (N_44259,N_42942,N_42058);
or U44260 (N_44260,N_42616,N_42525);
and U44261 (N_44261,N_43417,N_43574);
and U44262 (N_44262,N_42414,N_43818);
and U44263 (N_44263,N_42693,N_43020);
xnor U44264 (N_44264,N_43836,N_42200);
xnor U44265 (N_44265,N_43786,N_42726);
xnor U44266 (N_44266,N_43802,N_42904);
nor U44267 (N_44267,N_43012,N_43688);
xor U44268 (N_44268,N_43587,N_43136);
nor U44269 (N_44269,N_43308,N_42184);
or U44270 (N_44270,N_43261,N_42917);
xnor U44271 (N_44271,N_42470,N_42945);
nor U44272 (N_44272,N_42888,N_42580);
nand U44273 (N_44273,N_42074,N_43606);
and U44274 (N_44274,N_42458,N_43622);
or U44275 (N_44275,N_42670,N_43022);
nand U44276 (N_44276,N_42061,N_43450);
xor U44277 (N_44277,N_43491,N_42601);
and U44278 (N_44278,N_42719,N_42679);
and U44279 (N_44279,N_43977,N_43357);
nor U44280 (N_44280,N_43464,N_43771);
nor U44281 (N_44281,N_43514,N_43278);
xor U44282 (N_44282,N_43205,N_43936);
xnor U44283 (N_44283,N_43496,N_43310);
or U44284 (N_44284,N_43961,N_43397);
and U44285 (N_44285,N_43507,N_43860);
nand U44286 (N_44286,N_42126,N_43017);
and U44287 (N_44287,N_43653,N_43915);
xnor U44288 (N_44288,N_42408,N_43989);
or U44289 (N_44289,N_43213,N_43811);
or U44290 (N_44290,N_42027,N_42142);
or U44291 (N_44291,N_43719,N_43710);
and U44292 (N_44292,N_43633,N_42282);
xor U44293 (N_44293,N_42370,N_43926);
nor U44294 (N_44294,N_42329,N_42985);
or U44295 (N_44295,N_43516,N_43304);
nand U44296 (N_44296,N_42600,N_43782);
nor U44297 (N_44297,N_43228,N_42718);
or U44298 (N_44298,N_42821,N_43502);
or U44299 (N_44299,N_42652,N_43683);
xor U44300 (N_44300,N_43290,N_42833);
or U44301 (N_44301,N_43489,N_42351);
or U44302 (N_44302,N_42526,N_43463);
nor U44303 (N_44303,N_42473,N_43529);
nor U44304 (N_44304,N_42250,N_43713);
or U44305 (N_44305,N_43174,N_42312);
or U44306 (N_44306,N_43255,N_42509);
nand U44307 (N_44307,N_43865,N_42928);
and U44308 (N_44308,N_42100,N_43631);
and U44309 (N_44309,N_42936,N_43592);
xnor U44310 (N_44310,N_43288,N_43819);
xnor U44311 (N_44311,N_43866,N_42793);
xor U44312 (N_44312,N_42129,N_43374);
xor U44313 (N_44313,N_42266,N_42342);
nand U44314 (N_44314,N_43962,N_42276);
nand U44315 (N_44315,N_42528,N_43073);
nand U44316 (N_44316,N_42860,N_42179);
and U44317 (N_44317,N_42089,N_43217);
or U44318 (N_44318,N_43969,N_43795);
and U44319 (N_44319,N_42288,N_42434);
nand U44320 (N_44320,N_42640,N_42518);
or U44321 (N_44321,N_43349,N_42912);
nand U44322 (N_44322,N_42309,N_43339);
nand U44323 (N_44323,N_42608,N_42261);
nor U44324 (N_44324,N_43809,N_43265);
xor U44325 (N_44325,N_42961,N_43794);
and U44326 (N_44326,N_42976,N_43761);
nand U44327 (N_44327,N_43251,N_43585);
or U44328 (N_44328,N_43476,N_43311);
nor U44329 (N_44329,N_43301,N_42215);
xor U44330 (N_44330,N_43820,N_42154);
or U44331 (N_44331,N_42387,N_42597);
nand U44332 (N_44332,N_43812,N_43209);
nand U44333 (N_44333,N_43789,N_43286);
nor U44334 (N_44334,N_42360,N_43772);
xnor U44335 (N_44335,N_43048,N_42588);
or U44336 (N_44336,N_42972,N_42444);
xnor U44337 (N_44337,N_42677,N_42570);
and U44338 (N_44338,N_42088,N_43103);
nand U44339 (N_44339,N_42879,N_43831);
nor U44340 (N_44340,N_42286,N_43015);
nand U44341 (N_44341,N_43856,N_42157);
xor U44342 (N_44342,N_43167,N_43281);
and U44343 (N_44343,N_42141,N_43307);
and U44344 (N_44344,N_43857,N_43568);
nor U44345 (N_44345,N_43398,N_43779);
xnor U44346 (N_44346,N_42406,N_42569);
nand U44347 (N_44347,N_42803,N_42951);
or U44348 (N_44348,N_42427,N_42909);
xnor U44349 (N_44349,N_43729,N_42398);
nor U44350 (N_44350,N_42757,N_42042);
nor U44351 (N_44351,N_43849,N_43747);
nor U44352 (N_44352,N_43609,N_42875);
nand U44353 (N_44353,N_42931,N_43460);
nand U44354 (N_44354,N_43436,N_42764);
nand U44355 (N_44355,N_43333,N_43957);
or U44356 (N_44356,N_42663,N_42417);
nand U44357 (N_44357,N_43921,N_42517);
xor U44358 (N_44358,N_42974,N_43979);
xor U44359 (N_44359,N_43092,N_43113);
and U44360 (N_44360,N_43192,N_43885);
nand U44361 (N_44361,N_42030,N_42787);
nand U44362 (N_44362,N_42675,N_42705);
and U44363 (N_44363,N_43269,N_42524);
xor U44364 (N_44364,N_42949,N_42171);
and U44365 (N_44365,N_42534,N_42263);
or U44366 (N_44366,N_43116,N_42295);
nor U44367 (N_44367,N_43821,N_42883);
or U44368 (N_44368,N_42703,N_42085);
xor U44369 (N_44369,N_42762,N_43663);
or U44370 (N_44370,N_43662,N_43137);
and U44371 (N_44371,N_43078,N_43504);
nand U44372 (N_44372,N_42251,N_42319);
nand U44373 (N_44373,N_43475,N_43906);
and U44374 (N_44374,N_43970,N_42590);
xor U44375 (N_44375,N_42223,N_43223);
and U44376 (N_44376,N_42858,N_42245);
nand U44377 (N_44377,N_42267,N_42482);
and U44378 (N_44378,N_42136,N_43680);
xnor U44379 (N_44379,N_43244,N_43783);
or U44380 (N_44380,N_42910,N_42003);
or U44381 (N_44381,N_42669,N_43981);
xor U44382 (N_44382,N_42535,N_43128);
nand U44383 (N_44383,N_43050,N_42725);
xnor U44384 (N_44384,N_43071,N_43211);
xnor U44385 (N_44385,N_42734,N_42667);
or U44386 (N_44386,N_42823,N_43147);
or U44387 (N_44387,N_43893,N_43615);
nor U44388 (N_44388,N_42092,N_42348);
or U44389 (N_44389,N_43441,N_42451);
and U44390 (N_44390,N_43108,N_43472);
and U44391 (N_44391,N_43847,N_42109);
or U44392 (N_44392,N_42190,N_42523);
xnor U44393 (N_44393,N_42537,N_43355);
and U44394 (N_44394,N_42995,N_43069);
nor U44395 (N_44395,N_42964,N_42201);
nor U44396 (N_44396,N_43524,N_43508);
xor U44397 (N_44397,N_43203,N_43920);
or U44398 (N_44398,N_42975,N_43715);
nand U44399 (N_44399,N_42376,N_42708);
nor U44400 (N_44400,N_42091,N_43939);
nor U44401 (N_44401,N_43691,N_42824);
nor U44402 (N_44402,N_42225,N_42483);
xnor U44403 (N_44403,N_43933,N_42614);
nor U44404 (N_44404,N_42479,N_43446);
nor U44405 (N_44405,N_42565,N_43098);
nand U44406 (N_44406,N_42889,N_42262);
or U44407 (N_44407,N_42856,N_43953);
nor U44408 (N_44408,N_42257,N_43799);
xor U44409 (N_44409,N_42611,N_43983);
or U44410 (N_44410,N_42765,N_42933);
xor U44411 (N_44411,N_42522,N_42515);
nor U44412 (N_44412,N_43364,N_42099);
or U44413 (N_44413,N_43706,N_43238);
nor U44414 (N_44414,N_43023,N_42072);
nand U44415 (N_44415,N_42874,N_43387);
and U44416 (N_44416,N_42015,N_42820);
nor U44417 (N_44417,N_43164,N_42702);
and U44418 (N_44418,N_42932,N_43598);
xor U44419 (N_44419,N_43537,N_43610);
xnor U44420 (N_44420,N_43732,N_42773);
xor U44421 (N_44421,N_42116,N_42002);
xnor U44422 (N_44422,N_43369,N_42305);
nor U44423 (N_44423,N_42682,N_42758);
and U44424 (N_44424,N_43186,N_43438);
xor U44425 (N_44425,N_42125,N_43871);
or U44426 (N_44426,N_43384,N_42631);
nor U44427 (N_44427,N_42596,N_42343);
nor U44428 (N_44428,N_43551,N_43005);
and U44429 (N_44429,N_42837,N_42083);
or U44430 (N_44430,N_43984,N_42374);
nor U44431 (N_44431,N_42285,N_42546);
nor U44432 (N_44432,N_43185,N_43089);
or U44433 (N_44433,N_43723,N_43862);
and U44434 (N_44434,N_43039,N_43934);
xnor U44435 (N_44435,N_43375,N_42688);
or U44436 (N_44436,N_42203,N_42903);
nand U44437 (N_44437,N_43344,N_43254);
or U44438 (N_44438,N_42195,N_43396);
and U44439 (N_44439,N_42808,N_42922);
xor U44440 (N_44440,N_42271,N_43166);
nand U44441 (N_44441,N_43267,N_43144);
nand U44442 (N_44442,N_43335,N_43509);
nor U44443 (N_44443,N_42768,N_42727);
and U44444 (N_44444,N_42957,N_43908);
nor U44445 (N_44445,N_42323,N_43705);
xnor U44446 (N_44446,N_42071,N_43695);
or U44447 (N_44447,N_42045,N_42605);
xnor U44448 (N_44448,N_42356,N_43560);
or U44449 (N_44449,N_43196,N_42064);
nand U44450 (N_44450,N_43479,N_43282);
xor U44451 (N_44451,N_42234,N_43070);
or U44452 (N_44452,N_43513,N_42164);
and U44453 (N_44453,N_42873,N_42256);
nor U44454 (N_44454,N_42973,N_43521);
and U44455 (N_44455,N_42172,N_43682);
xor U44456 (N_44456,N_43990,N_42151);
nor U44457 (N_44457,N_42587,N_42209);
or U44458 (N_44458,N_43714,N_42352);
or U44459 (N_44459,N_42298,N_42863);
or U44460 (N_44460,N_43846,N_43105);
or U44461 (N_44461,N_42815,N_42701);
nand U44462 (N_44462,N_43007,N_42330);
xor U44463 (N_44463,N_42221,N_42969);
or U44464 (N_44464,N_43814,N_43728);
and U44465 (N_44465,N_43101,N_42681);
xnor U44466 (N_44466,N_43382,N_43139);
xor U44467 (N_44467,N_42057,N_43796);
and U44468 (N_44468,N_42010,N_42385);
nor U44469 (N_44469,N_42628,N_43480);
nor U44470 (N_44470,N_42771,N_42728);
nand U44471 (N_44471,N_43770,N_42084);
nand U44472 (N_44472,N_43888,N_43877);
xnor U44473 (N_44473,N_42935,N_43526);
nand U44474 (N_44474,N_42834,N_43077);
nand U44475 (N_44475,N_42593,N_43145);
nand U44476 (N_44476,N_43016,N_43154);
or U44477 (N_44477,N_42538,N_42645);
nand U44478 (N_44478,N_43233,N_43115);
or U44479 (N_44479,N_42333,N_42252);
xor U44480 (N_44480,N_43804,N_42798);
xor U44481 (N_44481,N_42676,N_42629);
nor U44482 (N_44482,N_43905,N_42599);
xnor U44483 (N_44483,N_43277,N_42613);
xor U44484 (N_44484,N_42871,N_42880);
nand U44485 (N_44485,N_43754,N_43321);
nand U44486 (N_44486,N_43416,N_42435);
xor U44487 (N_44487,N_42916,N_42742);
and U44488 (N_44488,N_43869,N_43756);
xnor U44489 (N_44489,N_43536,N_42455);
and U44490 (N_44490,N_42542,N_43900);
xor U44491 (N_44491,N_42244,N_43035);
nor U44492 (N_44492,N_42733,N_43402);
and U44493 (N_44493,N_43096,N_42735);
nor U44494 (N_44494,N_42108,N_43368);
nand U44495 (N_44495,N_43701,N_42051);
xor U44496 (N_44496,N_43546,N_43268);
nor U44497 (N_44497,N_43639,N_42169);
or U44498 (N_44498,N_42111,N_42174);
or U44499 (N_44499,N_43135,N_42946);
xnor U44500 (N_44500,N_43379,N_42008);
or U44501 (N_44501,N_42110,N_43808);
nor U44502 (N_44502,N_43863,N_43661);
or U44503 (N_44503,N_43161,N_43566);
xnor U44504 (N_44504,N_42485,N_43944);
and U44505 (N_44505,N_43220,N_42192);
nor U44506 (N_44506,N_43429,N_43243);
or U44507 (N_44507,N_43725,N_42744);
xor U44508 (N_44508,N_42213,N_42887);
or U44509 (N_44509,N_43126,N_42797);
nor U44510 (N_44510,N_42324,N_42776);
nand U44511 (N_44511,N_43743,N_43676);
xor U44512 (N_44512,N_43279,N_43950);
nor U44513 (N_44513,N_43839,N_43447);
nand U44514 (N_44514,N_43470,N_42382);
nor U44515 (N_44515,N_43987,N_42749);
nor U44516 (N_44516,N_42573,N_42332);
and U44517 (N_44517,N_42178,N_42297);
xor U44518 (N_44518,N_43583,N_42707);
nor U44519 (N_44519,N_42687,N_42775);
or U44520 (N_44520,N_43451,N_42607);
nor U44521 (N_44521,N_42231,N_42357);
xnor U44522 (N_44522,N_43297,N_43938);
nor U44523 (N_44523,N_43356,N_43009);
nor U44524 (N_44524,N_43671,N_42987);
or U44525 (N_44525,N_43280,N_43452);
nand U44526 (N_44526,N_42379,N_43870);
xnor U44527 (N_44527,N_43543,N_42943);
nand U44528 (N_44528,N_43090,N_42713);
xor U44529 (N_44529,N_42119,N_43717);
or U44530 (N_44530,N_43775,N_42626);
and U44531 (N_44531,N_42639,N_43591);
or U44532 (N_44532,N_43964,N_43171);
and U44533 (N_44533,N_42893,N_42530);
xnor U44534 (N_44534,N_42894,N_42448);
xor U44535 (N_44535,N_43780,N_42369);
xnor U44536 (N_44536,N_43614,N_42291);
nand U44537 (N_44537,N_43525,N_42604);
nor U44538 (N_44538,N_42489,N_42167);
nand U44539 (N_44539,N_42086,N_42488);
or U44540 (N_44540,N_43004,N_42411);
xnor U44541 (N_44541,N_43222,N_42919);
or U44542 (N_44542,N_42270,N_42177);
or U44543 (N_44543,N_43534,N_43972);
or U44544 (N_44544,N_42303,N_42849);
or U44545 (N_44545,N_43117,N_42627);
nor U44546 (N_44546,N_42337,N_43478);
nor U44547 (N_44547,N_42576,N_43389);
or U44548 (N_44548,N_43928,N_42046);
xnor U44549 (N_44549,N_42623,N_42760);
nor U44550 (N_44550,N_42690,N_43291);
nand U44551 (N_44551,N_43937,N_43868);
and U44552 (N_44552,N_42133,N_43351);
or U44553 (N_44553,N_43386,N_42137);
and U44554 (N_44554,N_42547,N_42877);
nor U44555 (N_44555,N_42781,N_43816);
xor U44556 (N_44556,N_42044,N_43570);
nor U44557 (N_44557,N_42851,N_43182);
and U44558 (N_44558,N_42721,N_43194);
and U44559 (N_44559,N_42140,N_43236);
nand U44560 (N_44560,N_43686,N_42965);
xnor U44561 (N_44561,N_42067,N_42620);
xnor U44562 (N_44562,N_43259,N_43837);
xnor U44563 (N_44563,N_43160,N_43319);
nor U44564 (N_44564,N_43049,N_43577);
nor U44565 (N_44565,N_42556,N_42659);
nor U44566 (N_44566,N_43041,N_42272);
xor U44567 (N_44567,N_43094,N_43058);
and U44568 (N_44568,N_43952,N_43889);
nand U44569 (N_44569,N_42991,N_43657);
or U44570 (N_44570,N_42867,N_43156);
and U44571 (N_44571,N_42658,N_42321);
xor U44572 (N_44572,N_43481,N_43736);
nand U44573 (N_44573,N_43764,N_42241);
nand U44574 (N_44574,N_43258,N_42281);
or U44575 (N_44575,N_42906,N_42069);
nor U44576 (N_44576,N_43346,N_43134);
or U44577 (N_44577,N_42011,N_43084);
and U44578 (N_44578,N_42898,N_42710);
xnor U44579 (N_44579,N_43390,N_42498);
nor U44580 (N_44580,N_43626,N_42034);
and U44581 (N_44581,N_43212,N_42730);
nand U44582 (N_44582,N_42853,N_43231);
and U44583 (N_44583,N_43257,N_42716);
and U44584 (N_44584,N_42754,N_42929);
and U44585 (N_44585,N_42310,N_43722);
or U44586 (N_44586,N_42236,N_42212);
nor U44587 (N_44587,N_42339,N_42712);
and U44588 (N_44588,N_42740,N_42574);
and U44589 (N_44589,N_43284,N_43127);
or U44590 (N_44590,N_43940,N_42756);
nor U44591 (N_44591,N_42886,N_43571);
nand U44592 (N_44592,N_42717,N_42558);
nor U44593 (N_44593,N_42750,N_42373);
nor U44594 (N_44594,N_43632,N_43506);
and U44595 (N_44595,N_43711,N_43617);
and U44596 (N_44596,N_42520,N_42026);
or U44597 (N_44597,N_43707,N_42428);
nand U44598 (N_44598,N_43065,N_43454);
xor U44599 (N_44599,N_42647,N_42706);
nor U44600 (N_44600,N_42104,N_43623);
nor U44601 (N_44601,N_43037,N_42304);
nor U44602 (N_44602,N_42567,N_43299);
nand U44603 (N_44603,N_42048,N_43190);
nor U44604 (N_44604,N_43252,N_42869);
and U44605 (N_44605,N_42774,N_43051);
or U44606 (N_44606,N_43354,N_42855);
and U44607 (N_44607,N_43143,N_42474);
or U44608 (N_44608,N_42307,N_42393);
xor U44609 (N_44609,N_42038,N_42422);
or U44610 (N_44610,N_42114,N_43391);
nand U44611 (N_44611,N_42346,N_42147);
nand U44612 (N_44612,N_42615,N_43580);
nor U44613 (N_44613,N_42087,N_43178);
nand U44614 (N_44614,N_43731,N_43482);
xnor U44615 (N_44615,N_42022,N_42674);
or U44616 (N_44616,N_43428,N_43927);
nand U44617 (N_44617,N_42861,N_43013);
or U44618 (N_44618,N_42143,N_42908);
nor U44619 (N_44619,N_43776,N_43019);
nand U44620 (N_44620,N_42850,N_42624);
nand U44621 (N_44621,N_42603,N_43604);
xor U44622 (N_44622,N_42978,N_42311);
and U44623 (N_44623,N_43474,N_42134);
and U44624 (N_44624,N_42409,N_43649);
nand U44625 (N_44625,N_43146,N_42780);
nor U44626 (N_44626,N_43229,N_42848);
nor U44627 (N_44627,N_43363,N_42769);
nand U44628 (N_44628,N_43745,N_42155);
or U44629 (N_44629,N_42274,N_43403);
or U44630 (N_44630,N_43685,N_42539);
or U44631 (N_44631,N_42181,N_42170);
nor U44632 (N_44632,N_43531,N_43911);
nand U44633 (N_44633,N_42090,N_43569);
nor U44634 (N_44634,N_43262,N_43320);
and U44635 (N_44635,N_42076,N_42594);
nand U44636 (N_44636,N_42287,N_43184);
or U44637 (N_44637,N_42441,N_43787);
or U44638 (N_44638,N_43674,N_43624);
and U44639 (N_44639,N_42656,N_42868);
xnor U44640 (N_44640,N_43030,N_42362);
nor U44641 (N_44641,N_43925,N_42243);
nand U44642 (N_44642,N_42439,N_42510);
or U44643 (N_44643,N_43724,N_43554);
or U44644 (N_44644,N_42581,N_43206);
nor U44645 (N_44645,N_42731,N_42437);
nand U44646 (N_44646,N_42081,N_42993);
xnor U44647 (N_44647,N_43678,N_43765);
xor U44648 (N_44648,N_42228,N_42828);
or U44649 (N_44649,N_42000,N_42189);
nand U44650 (N_44650,N_42819,N_43744);
and U44651 (N_44651,N_42618,N_43887);
nor U44652 (N_44652,N_42882,N_42070);
and U44653 (N_44653,N_42665,N_43826);
nor U44654 (N_44654,N_42582,N_43449);
nand U44655 (N_44655,N_43493,N_43106);
nand U44656 (N_44656,N_43091,N_43898);
xnor U44657 (N_44657,N_42024,N_43565);
and U44658 (N_44658,N_42237,N_42766);
xor U44659 (N_44659,N_43313,N_42810);
or U44660 (N_44660,N_42902,N_42680);
and U44661 (N_44661,N_42115,N_42561);
or U44662 (N_44662,N_43107,N_43159);
or U44663 (N_44663,N_42180,N_42275);
nand U44664 (N_44664,N_42938,N_42334);
or U44665 (N_44665,N_42859,N_42638);
and U44666 (N_44666,N_42410,N_43248);
nand U44667 (N_44667,N_42336,N_42404);
and U44668 (N_44668,N_42082,N_42842);
nand U44669 (N_44669,N_42646,N_42499);
nor U44670 (N_44670,N_42549,N_42533);
and U44671 (N_44671,N_42796,N_42469);
and U44672 (N_44672,N_43999,N_42248);
or U44673 (N_44673,N_42852,N_42198);
nor U44674 (N_44674,N_42159,N_43693);
and U44675 (N_44675,N_42461,N_43948);
xnor U44676 (N_44676,N_42364,N_42967);
nor U44677 (N_44677,N_42023,N_42583);
nor U44678 (N_44678,N_42619,N_42527);
nand U44679 (N_44679,N_42424,N_43325);
nor U44680 (N_44680,N_43242,N_42552);
nor U44681 (N_44681,N_42575,N_43024);
or U44682 (N_44682,N_42367,N_42865);
or U44683 (N_44683,N_43942,N_42318);
nor U44684 (N_44684,N_43247,N_42009);
nand U44685 (N_44685,N_43300,N_42920);
xnor U44686 (N_44686,N_43573,N_42788);
xor U44687 (N_44687,N_42194,N_42921);
nand U44688 (N_44688,N_43750,N_42486);
and U44689 (N_44689,N_43912,N_43825);
xor U44690 (N_44690,N_43625,N_43611);
nand U44691 (N_44691,N_43302,N_43235);
nor U44692 (N_44692,N_42840,N_43239);
nor U44693 (N_44693,N_43991,N_43405);
or U44694 (N_44694,N_43584,N_43312);
xnor U44695 (N_44695,N_43010,N_43427);
or U44696 (N_44696,N_43806,N_43006);
and U44697 (N_44697,N_43317,N_43326);
nor U44698 (N_44698,N_42278,N_42101);
nand U44699 (N_44699,N_42651,N_43040);
xor U44700 (N_44700,N_42732,N_43055);
and U44701 (N_44701,N_43681,N_43853);
or U44702 (N_44702,N_43130,N_43468);
xnor U44703 (N_44703,N_42006,N_43738);
nor U44704 (N_44704,N_43618,N_43575);
or U44705 (N_44705,N_42222,N_43150);
nand U44706 (N_44706,N_42511,N_43520);
xor U44707 (N_44707,N_43124,N_43640);
xnor U44708 (N_44708,N_42519,N_43498);
nand U44709 (N_44709,N_42654,N_42153);
nand U44710 (N_44710,N_43246,N_43752);
nand U44711 (N_44711,N_43294,N_43801);
nor U44712 (N_44712,N_43423,N_42454);
or U44713 (N_44713,N_43413,N_43457);
or U44714 (N_44714,N_43666,N_43643);
and U44715 (N_44715,N_42372,N_42761);
and U44716 (N_44716,N_43767,N_43285);
nand U44717 (N_44717,N_43982,N_43793);
nand U44718 (N_44718,N_43861,N_43902);
xor U44719 (N_44719,N_43791,N_42741);
xnor U44720 (N_44720,N_43359,N_43559);
xor U44721 (N_44721,N_42331,N_43433);
xnor U44722 (N_44722,N_43093,N_42007);
nor U44723 (N_44723,N_42885,N_42396);
or U44724 (N_44724,N_42106,N_43172);
nand U44725 (N_44725,N_43828,N_42653);
nand U44726 (N_44726,N_42224,N_42438);
xor U44727 (N_44727,N_42857,N_43916);
or U44728 (N_44728,N_42998,N_43930);
and U44729 (N_44729,N_42683,N_42426);
nor U44730 (N_44730,N_42700,N_42366);
and U44731 (N_44731,N_42947,N_43973);
nor U44732 (N_44732,N_42415,N_43810);
and U44733 (N_44733,N_42878,N_43679);
nand U44734 (N_44734,N_42532,N_42876);
xor U44735 (N_44735,N_42839,N_43230);
nor U44736 (N_44736,N_43726,N_43997);
or U44737 (N_44737,N_42145,N_43329);
or U44738 (N_44738,N_43558,N_42419);
xnor U44739 (N_44739,N_42992,N_43522);
xor U44740 (N_44740,N_42361,N_43785);
nor U44741 (N_44741,N_42279,N_43748);
nand U44742 (N_44742,N_43216,N_42445);
or U44743 (N_44743,N_43788,N_42952);
nor U44744 (N_44744,N_43140,N_43720);
nand U44745 (N_44745,N_42918,N_43567);
nand U44746 (N_44746,N_42105,N_42326);
nand U44747 (N_44747,N_42102,N_42453);
xor U44748 (N_44748,N_42572,N_42350);
nand U44749 (N_44749,N_43191,N_43648);
nor U44750 (N_44750,N_43309,N_42316);
nand U44751 (N_44751,N_43645,N_42513);
and U44752 (N_44752,N_42829,N_43859);
and U44753 (N_44753,N_42040,N_43381);
and U44754 (N_44754,N_42429,N_42063);
nand U44755 (N_44755,N_42930,N_43111);
xor U44756 (N_44756,N_43060,N_42802);
or U44757 (N_44757,N_42686,N_43305);
nor U44758 (N_44758,N_42811,N_42436);
nand U44759 (N_44759,N_42399,N_43064);
nor U44760 (N_44760,N_42818,N_43768);
nor U44761 (N_44761,N_43739,N_43169);
and U44762 (N_44762,N_43533,N_43173);
nand U44763 (N_44763,N_43541,N_43613);
xor U44764 (N_44764,N_43083,N_42751);
and U44765 (N_44765,N_42650,N_42763);
nand U44766 (N_44766,N_43044,N_43207);
or U44767 (N_44767,N_43530,N_42131);
and U44768 (N_44768,N_43085,N_42950);
and U44769 (N_44769,N_43664,N_42736);
and U44770 (N_44770,N_43505,N_42401);
xnor U44771 (N_44771,N_42685,N_43112);
and U44772 (N_44772,N_43331,N_43576);
nand U44773 (N_44773,N_43322,N_42341);
and U44774 (N_44774,N_43603,N_43393);
and U44775 (N_44775,N_43018,N_43241);
nor U44776 (N_44776,N_42585,N_43841);
nor U44777 (N_44777,N_43994,N_43380);
xor U44778 (N_44778,N_43204,N_42123);
xnor U44779 (N_44779,N_42512,N_42407);
and U44780 (N_44780,N_43518,N_43641);
nor U44781 (N_44781,N_42397,N_42191);
nor U44782 (N_44782,N_42817,N_43660);
xor U44783 (N_44783,N_42188,N_42468);
nand U44784 (N_44784,N_42899,N_43097);
or U44785 (N_44785,N_42240,N_43910);
xor U44786 (N_44786,N_43327,N_43121);
nand U44787 (N_44787,N_42836,N_42914);
xor U44788 (N_44788,N_42161,N_42505);
nand U44789 (N_44789,N_43245,N_42078);
and U44790 (N_44790,N_42956,N_42891);
xnor U44791 (N_44791,N_42866,N_43086);
xor U44792 (N_44792,N_42644,N_42907);
or U44793 (N_44793,N_42358,N_43131);
or U44794 (N_44794,N_42544,N_42475);
or U44795 (N_44795,N_42968,N_42621);
and U44796 (N_44796,N_43875,N_43045);
nor U44797 (N_44797,N_43434,N_42135);
nor U44798 (N_44798,N_43907,N_42496);
nand U44799 (N_44799,N_43879,N_42825);
nor U44800 (N_44800,N_43047,N_43833);
and U44801 (N_44801,N_43188,N_43385);
xor U44802 (N_44802,N_43538,N_43376);
nand U44803 (N_44803,N_42300,N_43740);
or U44804 (N_44804,N_43063,N_42363);
xor U44805 (N_44805,N_42862,N_43477);
xor U44806 (N_44806,N_42283,N_42529);
and U44807 (N_44807,N_43430,N_43494);
or U44808 (N_44808,N_42107,N_42630);
nor U44809 (N_44809,N_43323,N_42785);
and U44810 (N_44810,N_42456,N_42149);
or U44811 (N_44811,N_43336,N_42692);
and U44812 (N_44812,N_42477,N_43234);
nand U44813 (N_44813,N_43769,N_42031);
nand U44814 (N_44814,N_42389,N_42809);
nor U44815 (N_44815,N_42289,N_43122);
nand U44816 (N_44816,N_43593,N_43273);
and U44817 (N_44817,N_43751,N_43461);
nand U44818 (N_44818,N_43708,N_42598);
nor U44819 (N_44819,N_43968,N_42691);
xnor U44820 (N_44820,N_43486,N_43790);
nand U44821 (N_44821,N_43118,N_42405);
and U44822 (N_44822,N_43965,N_42507);
or U44823 (N_44823,N_42854,N_42014);
nor U44824 (N_44824,N_42986,N_43471);
or U44825 (N_44825,N_43367,N_43637);
nand U44826 (N_44826,N_42925,N_43890);
or U44827 (N_44827,N_42148,N_42163);
and U44828 (N_44828,N_42460,N_42381);
or U44829 (N_44829,N_43817,N_43998);
and U44830 (N_44830,N_42457,N_43296);
and U44831 (N_44831,N_42980,N_42452);
nand U44832 (N_44832,N_43696,N_42870);
nand U44833 (N_44833,N_42830,N_43882);
nand U44834 (N_44834,N_43158,N_43240);
nand U44835 (N_44835,N_43607,N_42394);
and U44836 (N_44836,N_42591,N_43421);
nand U44837 (N_44837,N_43895,N_43445);
xnor U44838 (N_44838,N_42551,N_43692);
and U44839 (N_44839,N_43986,N_42392);
nand U44840 (N_44840,N_43855,N_43654);
or U44841 (N_44841,N_42699,N_43919);
xnor U44842 (N_44842,N_42193,N_43628);
and U44843 (N_44843,N_43650,N_43088);
nand U44844 (N_44844,N_43072,N_43484);
xnor U44845 (N_44845,N_43909,N_43208);
and U44846 (N_44846,N_43540,N_43431);
xnor U44847 (N_44847,N_43515,N_43555);
nor U44848 (N_44848,N_42443,N_43298);
nor U44849 (N_44849,N_43703,N_43042);
nand U44850 (N_44850,N_42050,N_43700);
nand U44851 (N_44851,N_42937,N_43109);
or U44852 (N_44852,N_42294,N_42121);
and U44853 (N_44853,N_42832,N_42301);
nor U44854 (N_44854,N_43021,N_42386);
or U44855 (N_44855,N_42722,N_42233);
nand U44856 (N_44856,N_42080,N_42216);
or U44857 (N_44857,N_42940,N_43542);
xnor U44858 (N_44858,N_42714,N_42338);
nor U44859 (N_44859,N_42514,N_42464);
xnor U44860 (N_44860,N_42199,N_43125);
and U44861 (N_44861,N_43052,N_42229);
or U44862 (N_44862,N_43616,N_43873);
xnor U44863 (N_44863,N_43176,N_42207);
nand U44864 (N_44864,N_42845,N_43924);
or U44865 (N_44865,N_43218,N_42390);
xor U44866 (N_44866,N_42314,N_42890);
xor U44867 (N_44867,N_42079,N_43658);
and U44868 (N_44868,N_42258,N_42459);
nand U44869 (N_44869,N_43054,N_42559);
nand U44870 (N_44870,N_42097,N_42915);
xor U44871 (N_44871,N_43200,N_42497);
nor U44872 (N_44872,N_43621,N_42971);
nor U44873 (N_44873,N_42368,N_42897);
nor U44874 (N_44874,N_43193,N_42280);
and U44875 (N_44875,N_43437,N_42970);
and U44876 (N_44876,N_43792,N_43483);
nor U44877 (N_44877,N_43822,N_43210);
nand U44878 (N_44878,N_42077,N_43730);
xnor U44879 (N_44879,N_43975,N_43415);
and U44880 (N_44880,N_42622,N_43897);
nor U44881 (N_44881,N_43025,N_42467);
or U44882 (N_44882,N_42927,N_43741);
and U44883 (N_44883,N_42777,N_42146);
nand U44884 (N_44884,N_43227,N_42400);
and U44885 (N_44885,N_42208,N_43456);
or U44886 (N_44886,N_42431,N_42772);
nor U44887 (N_44887,N_43932,N_43306);
and U44888 (N_44888,N_42563,N_43800);
and U44889 (N_44889,N_42197,N_42695);
or U44890 (N_44890,N_42150,N_43499);
xnor U44891 (N_44891,N_43848,N_42941);
or U44892 (N_44892,N_43581,N_42391);
nand U44893 (N_44893,N_42152,N_43495);
or U44894 (N_44894,N_43803,N_42056);
nor U44895 (N_44895,N_43718,N_42449);
nand U44896 (N_44896,N_43651,N_42478);
nand U44897 (N_44897,N_43043,N_43340);
xnor U44898 (N_44898,N_43880,N_43293);
nand U44899 (N_44899,N_42012,N_42555);
xor U44900 (N_44900,N_42794,N_42755);
nor U44901 (N_44901,N_43197,N_42806);
and U44902 (N_44902,N_43945,N_43469);
xor U44903 (N_44903,N_42345,N_43448);
nand U44904 (N_44904,N_42521,N_42139);
and U44905 (N_44905,N_43694,N_43362);
or U44906 (N_44906,N_43737,N_42550);
nand U44907 (N_44907,N_42632,N_42095);
and U44908 (N_44908,N_43832,N_43353);
xnor U44909 (N_44909,N_42634,N_43377);
and U44910 (N_44910,N_43011,N_43742);
xor U44911 (N_44911,N_43440,N_42020);
nor U44912 (N_44912,N_42196,N_42049);
and U44913 (N_44913,N_42709,N_43797);
nand U44914 (N_44914,N_42664,N_43181);
xor U44915 (N_44915,N_43619,N_42264);
nand U44916 (N_44916,N_43138,N_43684);
xnor U44917 (N_44917,N_43914,N_43874);
nand U44918 (N_44918,N_42450,N_42383);
xnor U44919 (N_44919,N_42738,N_42543);
and U44920 (N_44920,N_42340,N_42900);
nor U44921 (N_44921,N_43838,N_43202);
nand U44922 (N_44922,N_42881,N_43563);
nand U44923 (N_44923,N_42548,N_43424);
nand U44924 (N_44924,N_43029,N_42901);
or U44925 (N_44925,N_42423,N_42325);
nand U44926 (N_44926,N_42371,N_43734);
nor U44927 (N_44927,N_43635,N_43978);
or U44928 (N_44928,N_43993,N_43620);
nand U44929 (N_44929,N_43157,N_42784);
nor U44930 (N_44930,N_43876,N_43334);
nor U44931 (N_44931,N_42259,N_43378);
or U44932 (N_44932,N_43453,N_42813);
or U44933 (N_44933,N_42206,N_43490);
nand U44934 (N_44934,N_42944,N_43917);
or U44935 (N_44935,N_42493,N_42506);
xor U44936 (N_44936,N_42767,N_43652);
nand U44937 (N_44937,N_42697,N_43214);
nor U44938 (N_44938,N_43941,N_43698);
nand U44939 (N_44939,N_42021,N_43342);
nor U44940 (N_44940,N_43155,N_43263);
nor U44941 (N_44941,N_42655,N_43903);
or U44942 (N_44942,N_42835,N_43561);
nand U44943 (N_44943,N_43550,N_42124);
or U44944 (N_44944,N_42795,N_42779);
and U44945 (N_44945,N_43963,N_43432);
or U44946 (N_44946,N_42013,N_43249);
and U44947 (N_44947,N_43884,N_43929);
xnor U44948 (N_44948,N_43076,N_43081);
or U44949 (N_44949,N_43886,N_43253);
and U44950 (N_44950,N_42981,N_43974);
and U44951 (N_44951,N_42737,N_42748);
nor U44952 (N_44952,N_42816,N_43074);
xnor U44953 (N_44953,N_42480,N_43985);
or U44954 (N_44954,N_42354,N_42689);
nand U44955 (N_44955,N_42982,N_43129);
nor U44956 (N_44956,N_43992,N_42117);
and U44957 (N_44957,N_43315,N_43061);
and U44958 (N_44958,N_43758,N_42503);
and U44959 (N_44959,N_43655,N_43901);
xor U44960 (N_44960,N_42807,N_43347);
and U44961 (N_44961,N_43599,N_43777);
nand U44962 (N_44962,N_42805,N_43026);
or U44963 (N_44963,N_42128,N_43062);
and U44964 (N_44964,N_43404,N_43670);
nand U44965 (N_44965,N_43123,N_42327);
and U44966 (N_44966,N_42720,N_43913);
and U44967 (N_44967,N_43638,N_43644);
nor U44968 (N_44968,N_42068,N_42745);
xor U44969 (N_44969,N_43669,N_43324);
and U44970 (N_44970,N_43830,N_43400);
and U44971 (N_44971,N_43557,N_42018);
and U44972 (N_44972,N_42290,N_43407);
nand U44973 (N_44973,N_43762,N_42562);
xor U44974 (N_44974,N_43854,N_43198);
xor U44975 (N_44975,N_43175,N_42465);
nor U44976 (N_44976,N_43303,N_43511);
and U44977 (N_44977,N_42571,N_42657);
nor U44978 (N_44978,N_42375,N_43760);
nor U44979 (N_44979,N_43881,N_42317);
or U44980 (N_44980,N_43935,N_42989);
nand U44981 (N_44981,N_43951,N_42160);
or U44982 (N_44982,N_42500,N_43582);
nand U44983 (N_44983,N_43590,N_42955);
nor U44984 (N_44984,N_43608,N_42268);
or U44985 (N_44985,N_43462,N_42001);
nor U44986 (N_44986,N_43547,N_42047);
nand U44987 (N_44987,N_43943,N_42847);
nor U44988 (N_44988,N_43753,N_43119);
xnor U44989 (N_44989,N_43348,N_42838);
nor U44990 (N_44990,N_43095,N_42211);
and U44991 (N_44991,N_42025,N_43594);
nor U44992 (N_44992,N_43589,N_43687);
nand U44993 (N_44993,N_43165,N_43394);
nand U44994 (N_44994,N_43852,N_43697);
or U44995 (N_44995,N_42491,N_43027);
nand U44996 (N_44996,N_42696,N_43370);
nand U44997 (N_44997,N_42666,N_43199);
or U44998 (N_44998,N_43727,N_42831);
nand U44999 (N_44999,N_43132,N_42694);
nand U45000 (N_45000,N_43368,N_43119);
or U45001 (N_45001,N_43438,N_43931);
xor U45002 (N_45002,N_43920,N_43100);
nor U45003 (N_45003,N_42279,N_42106);
or U45004 (N_45004,N_42415,N_43489);
nor U45005 (N_45005,N_43425,N_43612);
nand U45006 (N_45006,N_43037,N_42886);
nand U45007 (N_45007,N_42930,N_42470);
and U45008 (N_45008,N_42474,N_42743);
or U45009 (N_45009,N_42880,N_43998);
nor U45010 (N_45010,N_43973,N_43412);
and U45011 (N_45011,N_42822,N_42029);
and U45012 (N_45012,N_43514,N_42750);
nor U45013 (N_45013,N_43513,N_43140);
nor U45014 (N_45014,N_42718,N_42164);
and U45015 (N_45015,N_42091,N_43879);
or U45016 (N_45016,N_43158,N_43057);
or U45017 (N_45017,N_42525,N_43714);
nand U45018 (N_45018,N_43391,N_42368);
nor U45019 (N_45019,N_42340,N_42496);
or U45020 (N_45020,N_42409,N_43962);
and U45021 (N_45021,N_43500,N_43816);
nand U45022 (N_45022,N_43978,N_43995);
xor U45023 (N_45023,N_43567,N_42791);
nor U45024 (N_45024,N_43760,N_43828);
or U45025 (N_45025,N_42823,N_43674);
and U45026 (N_45026,N_43411,N_43726);
nor U45027 (N_45027,N_43054,N_43350);
xnor U45028 (N_45028,N_42846,N_43016);
nor U45029 (N_45029,N_42676,N_43974);
or U45030 (N_45030,N_42243,N_43920);
nor U45031 (N_45031,N_42798,N_43576);
xnor U45032 (N_45032,N_42629,N_43594);
nand U45033 (N_45033,N_43768,N_43779);
nand U45034 (N_45034,N_42547,N_42637);
or U45035 (N_45035,N_42900,N_43800);
xor U45036 (N_45036,N_42375,N_42966);
xor U45037 (N_45037,N_42441,N_42159);
nor U45038 (N_45038,N_42020,N_42181);
xor U45039 (N_45039,N_43804,N_42628);
xnor U45040 (N_45040,N_43862,N_43142);
and U45041 (N_45041,N_42212,N_42016);
and U45042 (N_45042,N_42758,N_42422);
or U45043 (N_45043,N_42078,N_42071);
and U45044 (N_45044,N_43505,N_43136);
nor U45045 (N_45045,N_42009,N_43452);
and U45046 (N_45046,N_42555,N_42232);
or U45047 (N_45047,N_43900,N_43015);
nand U45048 (N_45048,N_42329,N_42321);
nor U45049 (N_45049,N_43923,N_42761);
nand U45050 (N_45050,N_43718,N_43584);
nor U45051 (N_45051,N_43705,N_42859);
and U45052 (N_45052,N_42069,N_42454);
nand U45053 (N_45053,N_43373,N_43155);
xnor U45054 (N_45054,N_43189,N_43197);
xor U45055 (N_45055,N_42455,N_42170);
xnor U45056 (N_45056,N_42384,N_42492);
xor U45057 (N_45057,N_43282,N_43076);
xor U45058 (N_45058,N_43691,N_43444);
nand U45059 (N_45059,N_43142,N_43147);
or U45060 (N_45060,N_42522,N_42520);
and U45061 (N_45061,N_42210,N_42852);
nor U45062 (N_45062,N_43384,N_42371);
or U45063 (N_45063,N_43222,N_42321);
nand U45064 (N_45064,N_43571,N_43297);
xnor U45065 (N_45065,N_42082,N_42273);
nand U45066 (N_45066,N_43161,N_43864);
xor U45067 (N_45067,N_42222,N_42188);
nor U45068 (N_45068,N_43830,N_43540);
nand U45069 (N_45069,N_42459,N_43226);
nand U45070 (N_45070,N_42814,N_42871);
and U45071 (N_45071,N_43713,N_42200);
and U45072 (N_45072,N_42800,N_42207);
xnor U45073 (N_45073,N_43117,N_42847);
or U45074 (N_45074,N_43626,N_42745);
xnor U45075 (N_45075,N_42808,N_42407);
or U45076 (N_45076,N_42358,N_43049);
nand U45077 (N_45077,N_43607,N_43682);
nor U45078 (N_45078,N_43756,N_42963);
and U45079 (N_45079,N_43410,N_42751);
nor U45080 (N_45080,N_43760,N_43349);
and U45081 (N_45081,N_43737,N_42743);
nor U45082 (N_45082,N_43710,N_43264);
xor U45083 (N_45083,N_42271,N_43438);
nor U45084 (N_45084,N_42803,N_42350);
xnor U45085 (N_45085,N_43463,N_42403);
nand U45086 (N_45086,N_42093,N_42143);
nand U45087 (N_45087,N_43392,N_42759);
nand U45088 (N_45088,N_42299,N_43878);
and U45089 (N_45089,N_42331,N_42908);
xor U45090 (N_45090,N_43491,N_43060);
xor U45091 (N_45091,N_43779,N_43014);
and U45092 (N_45092,N_43108,N_43446);
nor U45093 (N_45093,N_43506,N_42639);
nor U45094 (N_45094,N_42934,N_42078);
nor U45095 (N_45095,N_43034,N_43727);
xor U45096 (N_45096,N_43063,N_43205);
nand U45097 (N_45097,N_42423,N_42947);
or U45098 (N_45098,N_43098,N_43439);
or U45099 (N_45099,N_42048,N_43715);
nand U45100 (N_45100,N_43701,N_43039);
nand U45101 (N_45101,N_42201,N_42253);
nand U45102 (N_45102,N_43453,N_42743);
nand U45103 (N_45103,N_43018,N_42643);
or U45104 (N_45104,N_43336,N_43111);
or U45105 (N_45105,N_42371,N_42512);
nand U45106 (N_45106,N_42315,N_42271);
nand U45107 (N_45107,N_42767,N_42916);
and U45108 (N_45108,N_43516,N_43604);
or U45109 (N_45109,N_43202,N_42413);
xnor U45110 (N_45110,N_42512,N_43865);
xor U45111 (N_45111,N_43787,N_43874);
or U45112 (N_45112,N_42362,N_42232);
nor U45113 (N_45113,N_42355,N_42972);
and U45114 (N_45114,N_43278,N_43026);
and U45115 (N_45115,N_43948,N_42204);
and U45116 (N_45116,N_43502,N_43699);
or U45117 (N_45117,N_43608,N_43845);
or U45118 (N_45118,N_42218,N_42049);
and U45119 (N_45119,N_43667,N_42308);
and U45120 (N_45120,N_43138,N_43041);
xor U45121 (N_45121,N_43311,N_43307);
xnor U45122 (N_45122,N_43986,N_42665);
xor U45123 (N_45123,N_42197,N_42967);
or U45124 (N_45124,N_42288,N_43441);
or U45125 (N_45125,N_42568,N_43798);
or U45126 (N_45126,N_42494,N_43624);
nand U45127 (N_45127,N_43331,N_42797);
or U45128 (N_45128,N_43541,N_43868);
nor U45129 (N_45129,N_42535,N_43624);
and U45130 (N_45130,N_43127,N_42826);
or U45131 (N_45131,N_42320,N_43239);
nor U45132 (N_45132,N_42184,N_42045);
nand U45133 (N_45133,N_42710,N_42299);
and U45134 (N_45134,N_42794,N_42533);
nand U45135 (N_45135,N_43138,N_43393);
and U45136 (N_45136,N_43681,N_43803);
nor U45137 (N_45137,N_42209,N_42846);
or U45138 (N_45138,N_43454,N_43900);
and U45139 (N_45139,N_42824,N_43972);
nor U45140 (N_45140,N_42487,N_42844);
nand U45141 (N_45141,N_42436,N_42665);
xor U45142 (N_45142,N_42405,N_42940);
nand U45143 (N_45143,N_42550,N_42402);
nand U45144 (N_45144,N_42995,N_43262);
or U45145 (N_45145,N_42269,N_42038);
and U45146 (N_45146,N_42994,N_42113);
xnor U45147 (N_45147,N_42179,N_43247);
nand U45148 (N_45148,N_42269,N_43435);
and U45149 (N_45149,N_42706,N_42443);
nand U45150 (N_45150,N_43319,N_42489);
and U45151 (N_45151,N_42784,N_42787);
xor U45152 (N_45152,N_42049,N_42896);
and U45153 (N_45153,N_42247,N_43058);
and U45154 (N_45154,N_42535,N_43351);
nand U45155 (N_45155,N_42145,N_43383);
xnor U45156 (N_45156,N_42896,N_42148);
nand U45157 (N_45157,N_42144,N_43523);
or U45158 (N_45158,N_43844,N_43438);
or U45159 (N_45159,N_43042,N_43904);
nor U45160 (N_45160,N_43045,N_43402);
xnor U45161 (N_45161,N_42751,N_42548);
or U45162 (N_45162,N_43482,N_42448);
and U45163 (N_45163,N_42550,N_43663);
nand U45164 (N_45164,N_42481,N_42143);
or U45165 (N_45165,N_43235,N_43190);
and U45166 (N_45166,N_43197,N_42857);
or U45167 (N_45167,N_42941,N_43073);
nand U45168 (N_45168,N_43501,N_43163);
and U45169 (N_45169,N_42962,N_43137);
xor U45170 (N_45170,N_43376,N_42563);
nand U45171 (N_45171,N_43533,N_43774);
nor U45172 (N_45172,N_42034,N_43973);
nor U45173 (N_45173,N_43833,N_42896);
and U45174 (N_45174,N_42031,N_43079);
nor U45175 (N_45175,N_43856,N_42291);
nand U45176 (N_45176,N_42107,N_42066);
nand U45177 (N_45177,N_42011,N_42870);
nor U45178 (N_45178,N_43423,N_42733);
nand U45179 (N_45179,N_43216,N_43625);
xor U45180 (N_45180,N_42232,N_42289);
nor U45181 (N_45181,N_43625,N_42882);
or U45182 (N_45182,N_43253,N_43056);
or U45183 (N_45183,N_43945,N_43198);
xnor U45184 (N_45184,N_43138,N_42175);
and U45185 (N_45185,N_42805,N_42744);
and U45186 (N_45186,N_43846,N_43317);
nand U45187 (N_45187,N_42142,N_43242);
nor U45188 (N_45188,N_43244,N_43471);
nor U45189 (N_45189,N_42412,N_43321);
nand U45190 (N_45190,N_43330,N_42628);
xor U45191 (N_45191,N_42861,N_43666);
nand U45192 (N_45192,N_42272,N_42769);
nor U45193 (N_45193,N_43177,N_43937);
or U45194 (N_45194,N_42672,N_42631);
nand U45195 (N_45195,N_43922,N_43779);
nor U45196 (N_45196,N_43609,N_42647);
nand U45197 (N_45197,N_43446,N_43760);
xor U45198 (N_45198,N_43334,N_42655);
or U45199 (N_45199,N_43297,N_42493);
nand U45200 (N_45200,N_43272,N_42770);
and U45201 (N_45201,N_42880,N_43628);
or U45202 (N_45202,N_42899,N_43033);
and U45203 (N_45203,N_42099,N_42558);
and U45204 (N_45204,N_43080,N_42521);
or U45205 (N_45205,N_42481,N_42885);
and U45206 (N_45206,N_43392,N_42288);
xor U45207 (N_45207,N_43905,N_42768);
and U45208 (N_45208,N_43278,N_43391);
xor U45209 (N_45209,N_43439,N_43102);
and U45210 (N_45210,N_43593,N_43901);
or U45211 (N_45211,N_42544,N_43492);
or U45212 (N_45212,N_43849,N_43429);
xor U45213 (N_45213,N_43593,N_42703);
xnor U45214 (N_45214,N_43790,N_42756);
nand U45215 (N_45215,N_42603,N_43889);
and U45216 (N_45216,N_42916,N_43580);
nor U45217 (N_45217,N_42265,N_43045);
xnor U45218 (N_45218,N_42224,N_43352);
and U45219 (N_45219,N_42422,N_43323);
nand U45220 (N_45220,N_42572,N_42749);
or U45221 (N_45221,N_42475,N_43323);
xnor U45222 (N_45222,N_43278,N_43500);
and U45223 (N_45223,N_42335,N_42135);
xnor U45224 (N_45224,N_43120,N_42090);
or U45225 (N_45225,N_43134,N_42012);
nand U45226 (N_45226,N_42346,N_42342);
nand U45227 (N_45227,N_42019,N_42832);
and U45228 (N_45228,N_42317,N_43892);
nand U45229 (N_45229,N_42144,N_43820);
or U45230 (N_45230,N_43951,N_43859);
and U45231 (N_45231,N_42371,N_43201);
or U45232 (N_45232,N_43590,N_42593);
nand U45233 (N_45233,N_43723,N_42798);
nand U45234 (N_45234,N_43075,N_43168);
and U45235 (N_45235,N_43709,N_42919);
and U45236 (N_45236,N_43144,N_42232);
and U45237 (N_45237,N_43624,N_42721);
xnor U45238 (N_45238,N_42364,N_43990);
nor U45239 (N_45239,N_43711,N_43805);
and U45240 (N_45240,N_42433,N_42371);
nand U45241 (N_45241,N_43455,N_42836);
or U45242 (N_45242,N_42059,N_42003);
or U45243 (N_45243,N_43498,N_43888);
xor U45244 (N_45244,N_42151,N_43559);
or U45245 (N_45245,N_43512,N_42884);
nand U45246 (N_45246,N_42149,N_42884);
or U45247 (N_45247,N_43763,N_42767);
or U45248 (N_45248,N_42659,N_43860);
xor U45249 (N_45249,N_43649,N_43339);
xnor U45250 (N_45250,N_43449,N_42464);
or U45251 (N_45251,N_42944,N_42179);
or U45252 (N_45252,N_42378,N_43012);
and U45253 (N_45253,N_42011,N_43597);
xor U45254 (N_45254,N_43251,N_43656);
nor U45255 (N_45255,N_43559,N_42169);
nor U45256 (N_45256,N_43663,N_42997);
or U45257 (N_45257,N_43708,N_43231);
xor U45258 (N_45258,N_43996,N_43166);
and U45259 (N_45259,N_42581,N_43648);
nor U45260 (N_45260,N_42073,N_42432);
xnor U45261 (N_45261,N_43689,N_42279);
nor U45262 (N_45262,N_43318,N_42830);
and U45263 (N_45263,N_43369,N_43273);
xor U45264 (N_45264,N_43115,N_42680);
or U45265 (N_45265,N_43991,N_42132);
xnor U45266 (N_45266,N_42392,N_43576);
or U45267 (N_45267,N_42966,N_42557);
and U45268 (N_45268,N_42616,N_42235);
nor U45269 (N_45269,N_43661,N_43035);
nor U45270 (N_45270,N_42215,N_43662);
nor U45271 (N_45271,N_42800,N_42929);
nor U45272 (N_45272,N_43916,N_43785);
nand U45273 (N_45273,N_42420,N_42625);
xor U45274 (N_45274,N_42690,N_42063);
or U45275 (N_45275,N_42843,N_43210);
and U45276 (N_45276,N_42344,N_43140);
nor U45277 (N_45277,N_43176,N_43136);
xnor U45278 (N_45278,N_42052,N_43449);
xor U45279 (N_45279,N_42072,N_42218);
or U45280 (N_45280,N_43817,N_43041);
nand U45281 (N_45281,N_42939,N_43909);
and U45282 (N_45282,N_42530,N_43935);
nand U45283 (N_45283,N_42280,N_43312);
and U45284 (N_45284,N_42369,N_42994);
xnor U45285 (N_45285,N_43191,N_42462);
nand U45286 (N_45286,N_43963,N_43303);
nand U45287 (N_45287,N_43508,N_43046);
or U45288 (N_45288,N_43699,N_42962);
nand U45289 (N_45289,N_42762,N_43167);
nor U45290 (N_45290,N_43040,N_42553);
and U45291 (N_45291,N_43031,N_43972);
nand U45292 (N_45292,N_42471,N_42223);
xnor U45293 (N_45293,N_42809,N_43311);
or U45294 (N_45294,N_43032,N_42613);
xor U45295 (N_45295,N_43563,N_43974);
nor U45296 (N_45296,N_42854,N_43158);
nor U45297 (N_45297,N_42910,N_43580);
and U45298 (N_45298,N_42184,N_42989);
nand U45299 (N_45299,N_43528,N_42532);
nor U45300 (N_45300,N_43459,N_43680);
xor U45301 (N_45301,N_43709,N_43642);
or U45302 (N_45302,N_42726,N_42197);
or U45303 (N_45303,N_42630,N_42200);
nor U45304 (N_45304,N_42373,N_42928);
nor U45305 (N_45305,N_43963,N_43811);
and U45306 (N_45306,N_43226,N_43711);
nor U45307 (N_45307,N_42100,N_42039);
nand U45308 (N_45308,N_43412,N_43943);
and U45309 (N_45309,N_42809,N_42663);
or U45310 (N_45310,N_42452,N_43941);
nand U45311 (N_45311,N_42867,N_42946);
and U45312 (N_45312,N_43991,N_43973);
nand U45313 (N_45313,N_43558,N_43178);
xnor U45314 (N_45314,N_42372,N_42752);
nor U45315 (N_45315,N_43953,N_43009);
or U45316 (N_45316,N_43796,N_43507);
and U45317 (N_45317,N_42867,N_42026);
nand U45318 (N_45318,N_42817,N_42310);
nand U45319 (N_45319,N_43206,N_43747);
nand U45320 (N_45320,N_43633,N_43442);
nand U45321 (N_45321,N_43364,N_42482);
and U45322 (N_45322,N_43781,N_42681);
xnor U45323 (N_45323,N_43986,N_42767);
and U45324 (N_45324,N_43876,N_42104);
or U45325 (N_45325,N_43596,N_43783);
nand U45326 (N_45326,N_43988,N_42586);
or U45327 (N_45327,N_42360,N_43387);
xor U45328 (N_45328,N_43657,N_43337);
xnor U45329 (N_45329,N_43549,N_43010);
nor U45330 (N_45330,N_42492,N_43551);
or U45331 (N_45331,N_42493,N_42890);
nor U45332 (N_45332,N_43563,N_43310);
nand U45333 (N_45333,N_42841,N_43860);
nor U45334 (N_45334,N_42580,N_42163);
and U45335 (N_45335,N_43094,N_42145);
xnor U45336 (N_45336,N_42160,N_42766);
nand U45337 (N_45337,N_43910,N_42171);
xnor U45338 (N_45338,N_43646,N_43002);
and U45339 (N_45339,N_42313,N_43949);
nor U45340 (N_45340,N_43377,N_42460);
or U45341 (N_45341,N_42471,N_42142);
or U45342 (N_45342,N_42274,N_43546);
xor U45343 (N_45343,N_42432,N_42043);
nand U45344 (N_45344,N_43411,N_42361);
xnor U45345 (N_45345,N_43899,N_42563);
xnor U45346 (N_45346,N_42502,N_43302);
and U45347 (N_45347,N_42076,N_42066);
or U45348 (N_45348,N_43743,N_43784);
nor U45349 (N_45349,N_42291,N_42546);
or U45350 (N_45350,N_43053,N_43976);
and U45351 (N_45351,N_42536,N_43728);
or U45352 (N_45352,N_43172,N_42544);
xnor U45353 (N_45353,N_42695,N_42032);
nand U45354 (N_45354,N_43666,N_43609);
or U45355 (N_45355,N_42191,N_43674);
or U45356 (N_45356,N_42315,N_42455);
and U45357 (N_45357,N_42305,N_43598);
nand U45358 (N_45358,N_43274,N_42630);
or U45359 (N_45359,N_42674,N_43464);
and U45360 (N_45360,N_42937,N_43463);
or U45361 (N_45361,N_42815,N_42058);
and U45362 (N_45362,N_43957,N_43293);
nor U45363 (N_45363,N_42790,N_42828);
xor U45364 (N_45364,N_42577,N_43250);
nand U45365 (N_45365,N_43119,N_42528);
nor U45366 (N_45366,N_43511,N_42853);
xor U45367 (N_45367,N_42083,N_43848);
or U45368 (N_45368,N_42400,N_43901);
xor U45369 (N_45369,N_42641,N_43239);
nand U45370 (N_45370,N_43321,N_43656);
xnor U45371 (N_45371,N_42571,N_43579);
and U45372 (N_45372,N_43202,N_43834);
nand U45373 (N_45373,N_43157,N_42297);
and U45374 (N_45374,N_42123,N_43044);
or U45375 (N_45375,N_43862,N_43988);
or U45376 (N_45376,N_42744,N_42594);
nand U45377 (N_45377,N_42288,N_42076);
nor U45378 (N_45378,N_43216,N_42693);
and U45379 (N_45379,N_42362,N_42847);
nor U45380 (N_45380,N_43646,N_42790);
nand U45381 (N_45381,N_43874,N_43166);
xor U45382 (N_45382,N_43022,N_43384);
or U45383 (N_45383,N_42119,N_42543);
nand U45384 (N_45384,N_42787,N_42058);
nor U45385 (N_45385,N_42223,N_43780);
xor U45386 (N_45386,N_42335,N_42197);
or U45387 (N_45387,N_43391,N_43357);
or U45388 (N_45388,N_43820,N_43059);
xnor U45389 (N_45389,N_43805,N_43936);
nand U45390 (N_45390,N_43547,N_42150);
or U45391 (N_45391,N_43483,N_43855);
and U45392 (N_45392,N_43670,N_43277);
and U45393 (N_45393,N_43298,N_42670);
xnor U45394 (N_45394,N_43816,N_42332);
xnor U45395 (N_45395,N_43807,N_42508);
nor U45396 (N_45396,N_42521,N_43841);
nor U45397 (N_45397,N_43601,N_42789);
xnor U45398 (N_45398,N_43272,N_42765);
and U45399 (N_45399,N_43565,N_43938);
or U45400 (N_45400,N_42342,N_43192);
xor U45401 (N_45401,N_42868,N_43950);
nor U45402 (N_45402,N_43300,N_42116);
nor U45403 (N_45403,N_43595,N_42769);
xor U45404 (N_45404,N_42364,N_42085);
nor U45405 (N_45405,N_42513,N_43345);
or U45406 (N_45406,N_43698,N_43344);
nor U45407 (N_45407,N_42750,N_43047);
nand U45408 (N_45408,N_43870,N_43214);
or U45409 (N_45409,N_43940,N_42759);
nand U45410 (N_45410,N_43111,N_42360);
xor U45411 (N_45411,N_42990,N_42603);
xor U45412 (N_45412,N_43809,N_43303);
nand U45413 (N_45413,N_42141,N_43973);
nor U45414 (N_45414,N_43092,N_43829);
nand U45415 (N_45415,N_42481,N_43873);
and U45416 (N_45416,N_42305,N_43866);
nand U45417 (N_45417,N_43980,N_43153);
and U45418 (N_45418,N_42332,N_42302);
nor U45419 (N_45419,N_43788,N_42153);
or U45420 (N_45420,N_43859,N_42939);
nand U45421 (N_45421,N_42602,N_43292);
nand U45422 (N_45422,N_43028,N_42275);
nor U45423 (N_45423,N_43318,N_42633);
nand U45424 (N_45424,N_42224,N_42346);
nand U45425 (N_45425,N_42924,N_42260);
nand U45426 (N_45426,N_43269,N_43238);
and U45427 (N_45427,N_43137,N_42975);
or U45428 (N_45428,N_42138,N_42797);
or U45429 (N_45429,N_42937,N_42335);
or U45430 (N_45430,N_43668,N_42781);
or U45431 (N_45431,N_43212,N_42620);
and U45432 (N_45432,N_42404,N_43206);
nand U45433 (N_45433,N_43714,N_42385);
xor U45434 (N_45434,N_43395,N_43350);
or U45435 (N_45435,N_43747,N_43823);
xor U45436 (N_45436,N_42264,N_43134);
nor U45437 (N_45437,N_43260,N_42747);
and U45438 (N_45438,N_43332,N_42521);
or U45439 (N_45439,N_43046,N_42970);
or U45440 (N_45440,N_42287,N_42414);
xor U45441 (N_45441,N_42708,N_42433);
and U45442 (N_45442,N_42016,N_43563);
xnor U45443 (N_45443,N_42306,N_43867);
nand U45444 (N_45444,N_43085,N_43651);
or U45445 (N_45445,N_43824,N_42256);
nor U45446 (N_45446,N_43509,N_43273);
nand U45447 (N_45447,N_42203,N_43136);
nor U45448 (N_45448,N_42326,N_43289);
and U45449 (N_45449,N_42898,N_43593);
nor U45450 (N_45450,N_42648,N_42953);
nor U45451 (N_45451,N_43874,N_42408);
xnor U45452 (N_45452,N_43645,N_43634);
nand U45453 (N_45453,N_42608,N_42404);
xnor U45454 (N_45454,N_43178,N_43218);
or U45455 (N_45455,N_42446,N_42270);
or U45456 (N_45456,N_42713,N_42046);
nand U45457 (N_45457,N_42775,N_43794);
and U45458 (N_45458,N_43863,N_42742);
and U45459 (N_45459,N_43489,N_42273);
and U45460 (N_45460,N_42142,N_42877);
or U45461 (N_45461,N_42596,N_43859);
xor U45462 (N_45462,N_42288,N_43018);
nor U45463 (N_45463,N_43360,N_42786);
and U45464 (N_45464,N_43949,N_43545);
xor U45465 (N_45465,N_43491,N_42872);
nand U45466 (N_45466,N_43856,N_42378);
and U45467 (N_45467,N_42546,N_42852);
nor U45468 (N_45468,N_43589,N_43430);
nor U45469 (N_45469,N_42920,N_42897);
nand U45470 (N_45470,N_42733,N_43100);
xnor U45471 (N_45471,N_42982,N_43220);
xor U45472 (N_45472,N_42630,N_42977);
nand U45473 (N_45473,N_42337,N_42425);
nor U45474 (N_45474,N_42012,N_43604);
nand U45475 (N_45475,N_42984,N_43366);
xor U45476 (N_45476,N_43587,N_43339);
xor U45477 (N_45477,N_43246,N_43361);
or U45478 (N_45478,N_42323,N_43762);
nand U45479 (N_45479,N_43837,N_43649);
xnor U45480 (N_45480,N_43655,N_43098);
xnor U45481 (N_45481,N_42426,N_42960);
and U45482 (N_45482,N_43070,N_43725);
nand U45483 (N_45483,N_43345,N_43513);
nor U45484 (N_45484,N_42758,N_43106);
or U45485 (N_45485,N_43528,N_42345);
and U45486 (N_45486,N_43961,N_42326);
nor U45487 (N_45487,N_43191,N_43343);
xor U45488 (N_45488,N_43875,N_42766);
and U45489 (N_45489,N_42881,N_42420);
and U45490 (N_45490,N_42128,N_42130);
nand U45491 (N_45491,N_42332,N_42043);
or U45492 (N_45492,N_43019,N_42925);
nor U45493 (N_45493,N_42029,N_43281);
and U45494 (N_45494,N_43679,N_43246);
nor U45495 (N_45495,N_43629,N_42701);
xnor U45496 (N_45496,N_42470,N_43827);
xnor U45497 (N_45497,N_42342,N_42696);
nand U45498 (N_45498,N_42858,N_43242);
or U45499 (N_45499,N_43998,N_42603);
and U45500 (N_45500,N_43017,N_42755);
nand U45501 (N_45501,N_42951,N_43745);
xor U45502 (N_45502,N_42614,N_43939);
and U45503 (N_45503,N_42415,N_42625);
and U45504 (N_45504,N_42274,N_43673);
nor U45505 (N_45505,N_43083,N_42998);
nand U45506 (N_45506,N_43537,N_43701);
or U45507 (N_45507,N_42307,N_43353);
and U45508 (N_45508,N_42261,N_43094);
nand U45509 (N_45509,N_42900,N_43690);
nor U45510 (N_45510,N_43695,N_43469);
or U45511 (N_45511,N_42675,N_42139);
nor U45512 (N_45512,N_43530,N_42094);
xor U45513 (N_45513,N_42298,N_43653);
xnor U45514 (N_45514,N_43024,N_43834);
xnor U45515 (N_45515,N_43167,N_43227);
xor U45516 (N_45516,N_43125,N_42311);
nand U45517 (N_45517,N_43424,N_42951);
nand U45518 (N_45518,N_43014,N_43035);
xor U45519 (N_45519,N_42821,N_42225);
nand U45520 (N_45520,N_42000,N_42323);
nor U45521 (N_45521,N_43503,N_42662);
nand U45522 (N_45522,N_42412,N_43180);
and U45523 (N_45523,N_43169,N_43656);
or U45524 (N_45524,N_42924,N_43734);
nand U45525 (N_45525,N_43486,N_43791);
xor U45526 (N_45526,N_42257,N_43401);
nand U45527 (N_45527,N_43861,N_43260);
and U45528 (N_45528,N_43645,N_42254);
nor U45529 (N_45529,N_43102,N_43053);
nand U45530 (N_45530,N_42133,N_43856);
nor U45531 (N_45531,N_42999,N_42950);
nor U45532 (N_45532,N_43346,N_43324);
and U45533 (N_45533,N_43843,N_43784);
or U45534 (N_45534,N_42359,N_43800);
nand U45535 (N_45535,N_43089,N_43926);
or U45536 (N_45536,N_42666,N_43237);
nand U45537 (N_45537,N_42321,N_42704);
nor U45538 (N_45538,N_42171,N_43023);
or U45539 (N_45539,N_43917,N_43605);
and U45540 (N_45540,N_43672,N_43678);
and U45541 (N_45541,N_43024,N_42152);
and U45542 (N_45542,N_43145,N_42735);
nand U45543 (N_45543,N_42228,N_42725);
or U45544 (N_45544,N_43801,N_43814);
and U45545 (N_45545,N_43629,N_42689);
and U45546 (N_45546,N_43265,N_42556);
nor U45547 (N_45547,N_43131,N_43926);
and U45548 (N_45548,N_43899,N_43430);
nor U45549 (N_45549,N_42370,N_43509);
nor U45550 (N_45550,N_42237,N_43924);
or U45551 (N_45551,N_43422,N_42990);
nand U45552 (N_45552,N_43816,N_43037);
xnor U45553 (N_45553,N_43822,N_43294);
nor U45554 (N_45554,N_42662,N_43923);
xnor U45555 (N_45555,N_42832,N_42742);
xor U45556 (N_45556,N_42124,N_42260);
nand U45557 (N_45557,N_43125,N_43544);
or U45558 (N_45558,N_42065,N_42719);
and U45559 (N_45559,N_43172,N_43741);
nand U45560 (N_45560,N_43062,N_42911);
nor U45561 (N_45561,N_42521,N_43285);
and U45562 (N_45562,N_43518,N_42094);
nand U45563 (N_45563,N_42297,N_42800);
and U45564 (N_45564,N_43516,N_42367);
xnor U45565 (N_45565,N_43235,N_42595);
and U45566 (N_45566,N_42453,N_42914);
xor U45567 (N_45567,N_42501,N_43128);
or U45568 (N_45568,N_43773,N_42445);
nand U45569 (N_45569,N_43420,N_42646);
nor U45570 (N_45570,N_43346,N_42952);
nand U45571 (N_45571,N_43055,N_42737);
xnor U45572 (N_45572,N_43273,N_43484);
and U45573 (N_45573,N_42309,N_42042);
nand U45574 (N_45574,N_42100,N_42853);
and U45575 (N_45575,N_42966,N_43927);
nand U45576 (N_45576,N_42399,N_42051);
and U45577 (N_45577,N_43599,N_43809);
xor U45578 (N_45578,N_42231,N_43550);
and U45579 (N_45579,N_42407,N_43524);
xnor U45580 (N_45580,N_42949,N_43994);
nor U45581 (N_45581,N_43516,N_42495);
nor U45582 (N_45582,N_42054,N_42649);
and U45583 (N_45583,N_43815,N_42699);
and U45584 (N_45584,N_42855,N_42823);
nand U45585 (N_45585,N_43331,N_43302);
xor U45586 (N_45586,N_42117,N_42382);
xnor U45587 (N_45587,N_43860,N_43717);
or U45588 (N_45588,N_42317,N_42681);
nand U45589 (N_45589,N_43326,N_42417);
xor U45590 (N_45590,N_43523,N_43622);
nor U45591 (N_45591,N_43194,N_43204);
xnor U45592 (N_45592,N_43557,N_42502);
and U45593 (N_45593,N_43843,N_43352);
nor U45594 (N_45594,N_43442,N_42743);
or U45595 (N_45595,N_43820,N_43805);
or U45596 (N_45596,N_43502,N_42083);
and U45597 (N_45597,N_42060,N_42805);
nor U45598 (N_45598,N_43362,N_43425);
nor U45599 (N_45599,N_43551,N_42583);
nor U45600 (N_45600,N_42964,N_42199);
nor U45601 (N_45601,N_42754,N_42132);
or U45602 (N_45602,N_42572,N_42443);
and U45603 (N_45603,N_43715,N_43481);
xor U45604 (N_45604,N_42608,N_42408);
xnor U45605 (N_45605,N_42435,N_43657);
and U45606 (N_45606,N_43171,N_43835);
or U45607 (N_45607,N_42454,N_42007);
xor U45608 (N_45608,N_42869,N_42879);
nand U45609 (N_45609,N_43783,N_43051);
and U45610 (N_45610,N_42434,N_42005);
xnor U45611 (N_45611,N_43585,N_42756);
xor U45612 (N_45612,N_42061,N_43249);
xnor U45613 (N_45613,N_42099,N_43490);
or U45614 (N_45614,N_43530,N_42943);
nand U45615 (N_45615,N_42108,N_43651);
nor U45616 (N_45616,N_42448,N_43177);
nor U45617 (N_45617,N_43938,N_42793);
xnor U45618 (N_45618,N_43691,N_42244);
or U45619 (N_45619,N_43302,N_42251);
nor U45620 (N_45620,N_42564,N_43049);
and U45621 (N_45621,N_42393,N_43854);
nand U45622 (N_45622,N_43577,N_42549);
and U45623 (N_45623,N_42540,N_42894);
nand U45624 (N_45624,N_42195,N_43516);
and U45625 (N_45625,N_43964,N_43686);
xnor U45626 (N_45626,N_43338,N_43902);
nand U45627 (N_45627,N_42549,N_42241);
nor U45628 (N_45628,N_42962,N_42508);
or U45629 (N_45629,N_43074,N_43554);
or U45630 (N_45630,N_43111,N_42927);
xor U45631 (N_45631,N_42981,N_42456);
or U45632 (N_45632,N_42271,N_42122);
or U45633 (N_45633,N_42886,N_43521);
xor U45634 (N_45634,N_42502,N_43928);
and U45635 (N_45635,N_42990,N_43274);
nand U45636 (N_45636,N_43379,N_42692);
or U45637 (N_45637,N_43538,N_43588);
and U45638 (N_45638,N_42596,N_43268);
nor U45639 (N_45639,N_43464,N_42110);
xor U45640 (N_45640,N_43458,N_42003);
and U45641 (N_45641,N_43560,N_43134);
and U45642 (N_45642,N_43934,N_42815);
or U45643 (N_45643,N_42640,N_42878);
xor U45644 (N_45644,N_43693,N_43330);
or U45645 (N_45645,N_43559,N_43333);
and U45646 (N_45646,N_43283,N_42582);
xor U45647 (N_45647,N_43209,N_42705);
and U45648 (N_45648,N_42880,N_43136);
nor U45649 (N_45649,N_43520,N_42910);
xnor U45650 (N_45650,N_42131,N_42615);
or U45651 (N_45651,N_43316,N_42104);
and U45652 (N_45652,N_42979,N_42932);
and U45653 (N_45653,N_42969,N_42224);
or U45654 (N_45654,N_42068,N_43616);
nand U45655 (N_45655,N_42083,N_42056);
nand U45656 (N_45656,N_43698,N_43251);
and U45657 (N_45657,N_43796,N_43536);
nand U45658 (N_45658,N_42435,N_43505);
nor U45659 (N_45659,N_42188,N_42739);
nor U45660 (N_45660,N_43067,N_42933);
and U45661 (N_45661,N_42053,N_42871);
xnor U45662 (N_45662,N_42675,N_42126);
nand U45663 (N_45663,N_43369,N_43788);
nor U45664 (N_45664,N_42113,N_43465);
and U45665 (N_45665,N_43412,N_43364);
nand U45666 (N_45666,N_43743,N_43239);
and U45667 (N_45667,N_42831,N_43576);
nor U45668 (N_45668,N_43701,N_42850);
and U45669 (N_45669,N_43575,N_43332);
nor U45670 (N_45670,N_43364,N_43172);
or U45671 (N_45671,N_42010,N_42651);
nor U45672 (N_45672,N_43128,N_42914);
and U45673 (N_45673,N_43555,N_43274);
nor U45674 (N_45674,N_42502,N_42837);
nand U45675 (N_45675,N_42313,N_42406);
xnor U45676 (N_45676,N_42500,N_43057);
xor U45677 (N_45677,N_43247,N_43478);
xnor U45678 (N_45678,N_42141,N_42056);
or U45679 (N_45679,N_43502,N_42338);
and U45680 (N_45680,N_42087,N_43751);
xnor U45681 (N_45681,N_42258,N_42503);
xnor U45682 (N_45682,N_43441,N_42045);
xor U45683 (N_45683,N_43254,N_42905);
xnor U45684 (N_45684,N_43843,N_42414);
nor U45685 (N_45685,N_43138,N_43444);
or U45686 (N_45686,N_42903,N_43100);
nor U45687 (N_45687,N_43298,N_43661);
nand U45688 (N_45688,N_43950,N_43581);
or U45689 (N_45689,N_43235,N_43613);
nor U45690 (N_45690,N_43634,N_42084);
nand U45691 (N_45691,N_43661,N_42200);
and U45692 (N_45692,N_42471,N_43823);
and U45693 (N_45693,N_43903,N_42654);
nand U45694 (N_45694,N_42955,N_43306);
nand U45695 (N_45695,N_43899,N_43768);
and U45696 (N_45696,N_42580,N_42332);
xor U45697 (N_45697,N_42408,N_43723);
nand U45698 (N_45698,N_42157,N_43280);
or U45699 (N_45699,N_43182,N_42856);
and U45700 (N_45700,N_43359,N_42592);
nand U45701 (N_45701,N_42387,N_43244);
and U45702 (N_45702,N_43639,N_42916);
nor U45703 (N_45703,N_42941,N_43195);
or U45704 (N_45704,N_42430,N_43688);
or U45705 (N_45705,N_43937,N_42153);
nor U45706 (N_45706,N_43559,N_43767);
xnor U45707 (N_45707,N_43040,N_42739);
or U45708 (N_45708,N_42142,N_42990);
nand U45709 (N_45709,N_43688,N_42731);
or U45710 (N_45710,N_43276,N_42207);
or U45711 (N_45711,N_42210,N_42859);
or U45712 (N_45712,N_42890,N_43386);
xor U45713 (N_45713,N_42905,N_43541);
nand U45714 (N_45714,N_43513,N_42897);
nor U45715 (N_45715,N_42124,N_43695);
and U45716 (N_45716,N_42022,N_42499);
nand U45717 (N_45717,N_42820,N_43272);
and U45718 (N_45718,N_43298,N_43012);
nor U45719 (N_45719,N_42597,N_42484);
nor U45720 (N_45720,N_42320,N_42019);
or U45721 (N_45721,N_42570,N_42839);
and U45722 (N_45722,N_42070,N_43645);
or U45723 (N_45723,N_42349,N_43839);
nor U45724 (N_45724,N_43472,N_43239);
and U45725 (N_45725,N_42912,N_43744);
nand U45726 (N_45726,N_43634,N_42735);
xor U45727 (N_45727,N_43380,N_43354);
or U45728 (N_45728,N_42325,N_42238);
nand U45729 (N_45729,N_43958,N_42189);
nor U45730 (N_45730,N_42030,N_43037);
or U45731 (N_45731,N_42009,N_42404);
or U45732 (N_45732,N_43800,N_42101);
nor U45733 (N_45733,N_42816,N_43308);
nand U45734 (N_45734,N_43852,N_43687);
nor U45735 (N_45735,N_43480,N_42062);
and U45736 (N_45736,N_43317,N_43577);
nand U45737 (N_45737,N_42014,N_42346);
xor U45738 (N_45738,N_43207,N_43208);
or U45739 (N_45739,N_43450,N_43798);
nand U45740 (N_45740,N_43376,N_42512);
nor U45741 (N_45741,N_43938,N_43242);
nand U45742 (N_45742,N_42709,N_42980);
and U45743 (N_45743,N_43237,N_43705);
nor U45744 (N_45744,N_43744,N_43134);
or U45745 (N_45745,N_43787,N_43465);
or U45746 (N_45746,N_43145,N_42578);
nand U45747 (N_45747,N_43730,N_42017);
xor U45748 (N_45748,N_43244,N_43344);
xor U45749 (N_45749,N_43110,N_42483);
nand U45750 (N_45750,N_43314,N_43079);
or U45751 (N_45751,N_42102,N_42720);
nand U45752 (N_45752,N_43968,N_42719);
or U45753 (N_45753,N_43948,N_43552);
and U45754 (N_45754,N_42099,N_43520);
xor U45755 (N_45755,N_42931,N_43427);
nand U45756 (N_45756,N_42052,N_42427);
or U45757 (N_45757,N_43936,N_42960);
xnor U45758 (N_45758,N_42732,N_43231);
nand U45759 (N_45759,N_42430,N_43398);
xor U45760 (N_45760,N_43479,N_42562);
xor U45761 (N_45761,N_43957,N_43560);
nand U45762 (N_45762,N_42792,N_42921);
or U45763 (N_45763,N_42780,N_42934);
xor U45764 (N_45764,N_42369,N_42905);
nand U45765 (N_45765,N_42894,N_43658);
nor U45766 (N_45766,N_43597,N_42546);
nand U45767 (N_45767,N_42449,N_42035);
and U45768 (N_45768,N_42303,N_43356);
nor U45769 (N_45769,N_43505,N_43554);
and U45770 (N_45770,N_42826,N_43455);
and U45771 (N_45771,N_42503,N_43986);
nor U45772 (N_45772,N_42407,N_42297);
nand U45773 (N_45773,N_43478,N_43948);
and U45774 (N_45774,N_43500,N_43496);
and U45775 (N_45775,N_43364,N_42255);
nand U45776 (N_45776,N_42149,N_43970);
xor U45777 (N_45777,N_43321,N_43998);
nand U45778 (N_45778,N_43542,N_42675);
xnor U45779 (N_45779,N_43422,N_43986);
nor U45780 (N_45780,N_42354,N_43355);
or U45781 (N_45781,N_42928,N_42407);
nand U45782 (N_45782,N_42969,N_42787);
and U45783 (N_45783,N_43103,N_43497);
or U45784 (N_45784,N_43531,N_42416);
or U45785 (N_45785,N_42461,N_43197);
nor U45786 (N_45786,N_42274,N_42822);
nor U45787 (N_45787,N_43601,N_42613);
and U45788 (N_45788,N_43646,N_43000);
xnor U45789 (N_45789,N_42408,N_42994);
or U45790 (N_45790,N_42918,N_43937);
nand U45791 (N_45791,N_43063,N_43231);
nand U45792 (N_45792,N_43199,N_43083);
xor U45793 (N_45793,N_42457,N_42003);
xnor U45794 (N_45794,N_43063,N_42641);
xor U45795 (N_45795,N_42615,N_42099);
and U45796 (N_45796,N_42302,N_43949);
or U45797 (N_45797,N_42126,N_43898);
nor U45798 (N_45798,N_43726,N_42728);
or U45799 (N_45799,N_43924,N_42678);
nand U45800 (N_45800,N_43094,N_43056);
nor U45801 (N_45801,N_42342,N_43638);
nor U45802 (N_45802,N_42746,N_42616);
and U45803 (N_45803,N_43706,N_43113);
nand U45804 (N_45804,N_42796,N_43884);
nor U45805 (N_45805,N_42710,N_43769);
or U45806 (N_45806,N_43559,N_42148);
nor U45807 (N_45807,N_42531,N_43549);
nor U45808 (N_45808,N_42878,N_43682);
xor U45809 (N_45809,N_42151,N_43029);
and U45810 (N_45810,N_43192,N_43010);
xor U45811 (N_45811,N_42532,N_42189);
xor U45812 (N_45812,N_43700,N_42851);
nor U45813 (N_45813,N_42958,N_42467);
nor U45814 (N_45814,N_43241,N_43310);
and U45815 (N_45815,N_43451,N_42928);
nand U45816 (N_45816,N_42503,N_43416);
xnor U45817 (N_45817,N_42534,N_43475);
nand U45818 (N_45818,N_42129,N_43380);
nor U45819 (N_45819,N_43264,N_42502);
xnor U45820 (N_45820,N_43566,N_42356);
xor U45821 (N_45821,N_43555,N_42502);
nand U45822 (N_45822,N_43839,N_42383);
xor U45823 (N_45823,N_43325,N_43549);
xor U45824 (N_45824,N_43115,N_42463);
and U45825 (N_45825,N_42671,N_42960);
xor U45826 (N_45826,N_42592,N_42128);
nand U45827 (N_45827,N_42773,N_43993);
and U45828 (N_45828,N_43479,N_42766);
xnor U45829 (N_45829,N_42175,N_42101);
xor U45830 (N_45830,N_42097,N_42932);
xnor U45831 (N_45831,N_43945,N_42393);
nor U45832 (N_45832,N_43018,N_43867);
nand U45833 (N_45833,N_42228,N_43409);
nor U45834 (N_45834,N_43684,N_43626);
and U45835 (N_45835,N_42416,N_42484);
nor U45836 (N_45836,N_43782,N_42319);
and U45837 (N_45837,N_42478,N_43680);
nor U45838 (N_45838,N_42214,N_42188);
or U45839 (N_45839,N_42158,N_42948);
nand U45840 (N_45840,N_42617,N_42946);
and U45841 (N_45841,N_42840,N_43345);
and U45842 (N_45842,N_42179,N_43478);
or U45843 (N_45843,N_42198,N_43177);
and U45844 (N_45844,N_42822,N_43971);
or U45845 (N_45845,N_42343,N_43199);
nand U45846 (N_45846,N_43714,N_42235);
xnor U45847 (N_45847,N_42623,N_42697);
and U45848 (N_45848,N_42847,N_43132);
and U45849 (N_45849,N_43915,N_43893);
xnor U45850 (N_45850,N_42373,N_43949);
or U45851 (N_45851,N_43025,N_42380);
or U45852 (N_45852,N_43904,N_42224);
or U45853 (N_45853,N_42618,N_42271);
nand U45854 (N_45854,N_43615,N_42165);
and U45855 (N_45855,N_42805,N_43446);
and U45856 (N_45856,N_42059,N_42656);
and U45857 (N_45857,N_43619,N_43049);
nand U45858 (N_45858,N_42762,N_42359);
nor U45859 (N_45859,N_42700,N_43054);
or U45860 (N_45860,N_43569,N_42597);
nor U45861 (N_45861,N_43666,N_43060);
xor U45862 (N_45862,N_43042,N_43613);
nand U45863 (N_45863,N_42766,N_42344);
or U45864 (N_45864,N_43760,N_43722);
nand U45865 (N_45865,N_43463,N_43752);
and U45866 (N_45866,N_42138,N_43370);
nand U45867 (N_45867,N_42834,N_42148);
nand U45868 (N_45868,N_43062,N_42041);
or U45869 (N_45869,N_42629,N_43687);
and U45870 (N_45870,N_42939,N_42973);
nand U45871 (N_45871,N_42051,N_42038);
and U45872 (N_45872,N_42887,N_42567);
or U45873 (N_45873,N_43569,N_42870);
nand U45874 (N_45874,N_43054,N_42024);
and U45875 (N_45875,N_42290,N_43181);
nand U45876 (N_45876,N_43296,N_43170);
nand U45877 (N_45877,N_42448,N_43428);
nand U45878 (N_45878,N_43019,N_42802);
nor U45879 (N_45879,N_42402,N_42628);
xor U45880 (N_45880,N_42612,N_42274);
nand U45881 (N_45881,N_42649,N_43035);
or U45882 (N_45882,N_42123,N_43808);
nor U45883 (N_45883,N_43631,N_42283);
xnor U45884 (N_45884,N_43696,N_43721);
nand U45885 (N_45885,N_42555,N_43626);
xnor U45886 (N_45886,N_43747,N_43670);
xor U45887 (N_45887,N_42215,N_43183);
xor U45888 (N_45888,N_42289,N_42526);
nand U45889 (N_45889,N_42777,N_42883);
nand U45890 (N_45890,N_42989,N_42176);
nor U45891 (N_45891,N_43202,N_42071);
or U45892 (N_45892,N_42331,N_43704);
or U45893 (N_45893,N_43994,N_42087);
nand U45894 (N_45894,N_43930,N_43489);
and U45895 (N_45895,N_42373,N_42757);
xor U45896 (N_45896,N_43633,N_42227);
xor U45897 (N_45897,N_42926,N_43015);
nor U45898 (N_45898,N_42221,N_43129);
xor U45899 (N_45899,N_43960,N_42184);
nand U45900 (N_45900,N_42459,N_42794);
nand U45901 (N_45901,N_43852,N_42160);
and U45902 (N_45902,N_43808,N_42397);
and U45903 (N_45903,N_42057,N_43994);
and U45904 (N_45904,N_43786,N_43754);
or U45905 (N_45905,N_42617,N_43302);
and U45906 (N_45906,N_42896,N_43054);
nand U45907 (N_45907,N_43571,N_43734);
xnor U45908 (N_45908,N_43383,N_42352);
nor U45909 (N_45909,N_43983,N_43507);
xnor U45910 (N_45910,N_43510,N_43978);
xnor U45911 (N_45911,N_43909,N_43724);
or U45912 (N_45912,N_42405,N_43487);
or U45913 (N_45913,N_43568,N_43889);
nand U45914 (N_45914,N_43324,N_42311);
or U45915 (N_45915,N_43140,N_42228);
and U45916 (N_45916,N_43572,N_43717);
nand U45917 (N_45917,N_42338,N_42517);
or U45918 (N_45918,N_42154,N_43139);
xnor U45919 (N_45919,N_42516,N_43204);
and U45920 (N_45920,N_42337,N_42576);
and U45921 (N_45921,N_42756,N_42598);
nor U45922 (N_45922,N_42667,N_43204);
or U45923 (N_45923,N_43102,N_42949);
nor U45924 (N_45924,N_43112,N_43579);
nand U45925 (N_45925,N_42738,N_43204);
or U45926 (N_45926,N_42850,N_43247);
nand U45927 (N_45927,N_43406,N_42655);
nand U45928 (N_45928,N_43535,N_42384);
and U45929 (N_45929,N_43372,N_42686);
nand U45930 (N_45930,N_43876,N_42161);
xor U45931 (N_45931,N_42685,N_42390);
or U45932 (N_45932,N_43980,N_42217);
and U45933 (N_45933,N_42838,N_43143);
or U45934 (N_45934,N_43831,N_42521);
and U45935 (N_45935,N_42505,N_42761);
xnor U45936 (N_45936,N_42574,N_42058);
nor U45937 (N_45937,N_42501,N_42725);
and U45938 (N_45938,N_42154,N_43567);
or U45939 (N_45939,N_43307,N_42262);
and U45940 (N_45940,N_42173,N_43457);
and U45941 (N_45941,N_42973,N_42727);
nand U45942 (N_45942,N_42155,N_42521);
nor U45943 (N_45943,N_43808,N_42485);
and U45944 (N_45944,N_42063,N_42360);
nor U45945 (N_45945,N_43120,N_42045);
and U45946 (N_45946,N_42702,N_43369);
xor U45947 (N_45947,N_42841,N_43492);
and U45948 (N_45948,N_42599,N_42328);
nor U45949 (N_45949,N_43964,N_42632);
nand U45950 (N_45950,N_43138,N_43772);
nand U45951 (N_45951,N_42217,N_42759);
nand U45952 (N_45952,N_42664,N_43413);
or U45953 (N_45953,N_43256,N_43496);
and U45954 (N_45954,N_42550,N_43071);
or U45955 (N_45955,N_42003,N_43323);
and U45956 (N_45956,N_42941,N_43070);
nand U45957 (N_45957,N_43436,N_43362);
nor U45958 (N_45958,N_42807,N_42665);
and U45959 (N_45959,N_42903,N_43735);
nor U45960 (N_45960,N_42752,N_43104);
nand U45961 (N_45961,N_42026,N_43733);
or U45962 (N_45962,N_43834,N_43507);
xor U45963 (N_45963,N_43183,N_43391);
nand U45964 (N_45964,N_43891,N_42389);
nand U45965 (N_45965,N_42094,N_42254);
and U45966 (N_45966,N_42367,N_42877);
nand U45967 (N_45967,N_43237,N_42322);
nor U45968 (N_45968,N_43331,N_43708);
nor U45969 (N_45969,N_42637,N_43405);
nor U45970 (N_45970,N_43804,N_42706);
nor U45971 (N_45971,N_42222,N_43107);
nand U45972 (N_45972,N_42928,N_42845);
or U45973 (N_45973,N_43450,N_42498);
nand U45974 (N_45974,N_42048,N_43816);
or U45975 (N_45975,N_42932,N_42275);
nor U45976 (N_45976,N_42682,N_42613);
and U45977 (N_45977,N_42168,N_43716);
nor U45978 (N_45978,N_43531,N_42014);
nor U45979 (N_45979,N_42004,N_42794);
nor U45980 (N_45980,N_43999,N_43303);
and U45981 (N_45981,N_43465,N_43054);
or U45982 (N_45982,N_42812,N_42257);
xnor U45983 (N_45983,N_43660,N_43129);
and U45984 (N_45984,N_43901,N_43094);
xor U45985 (N_45985,N_42731,N_42284);
nand U45986 (N_45986,N_42501,N_42450);
nor U45987 (N_45987,N_42546,N_43015);
nor U45988 (N_45988,N_42483,N_43772);
and U45989 (N_45989,N_42619,N_42308);
and U45990 (N_45990,N_43434,N_43309);
nand U45991 (N_45991,N_42290,N_43091);
and U45992 (N_45992,N_43536,N_42588);
nor U45993 (N_45993,N_43307,N_43373);
or U45994 (N_45994,N_43382,N_42535);
xor U45995 (N_45995,N_42217,N_43244);
or U45996 (N_45996,N_42934,N_42729);
nor U45997 (N_45997,N_42481,N_43811);
xor U45998 (N_45998,N_43573,N_43997);
nor U45999 (N_45999,N_43387,N_43683);
and U46000 (N_46000,N_45622,N_44068);
nand U46001 (N_46001,N_45416,N_44732);
nand U46002 (N_46002,N_45571,N_45355);
or U46003 (N_46003,N_44558,N_45884);
and U46004 (N_46004,N_44135,N_45332);
and U46005 (N_46005,N_45360,N_45500);
and U46006 (N_46006,N_44997,N_44377);
nand U46007 (N_46007,N_45475,N_44969);
nand U46008 (N_46008,N_45406,N_44594);
xnor U46009 (N_46009,N_45142,N_45287);
nand U46010 (N_46010,N_44866,N_44101);
nor U46011 (N_46011,N_45684,N_44011);
nor U46012 (N_46012,N_45450,N_45894);
nor U46013 (N_46013,N_44102,N_44167);
xor U46014 (N_46014,N_44878,N_45898);
and U46015 (N_46015,N_44643,N_44257);
or U46016 (N_46016,N_44812,N_45328);
or U46017 (N_46017,N_44548,N_44184);
nand U46018 (N_46018,N_44954,N_44958);
nand U46019 (N_46019,N_45384,N_45508);
and U46020 (N_46020,N_45659,N_45742);
xor U46021 (N_46021,N_45945,N_44961);
nand U46022 (N_46022,N_44745,N_44631);
and U46023 (N_46023,N_44985,N_44026);
or U46024 (N_46024,N_44659,N_45130);
nand U46025 (N_46025,N_44714,N_45433);
nand U46026 (N_46026,N_44045,N_45566);
nor U46027 (N_46027,N_45067,N_44429);
nand U46028 (N_46028,N_44630,N_45310);
nand U46029 (N_46029,N_44953,N_45291);
nand U46030 (N_46030,N_45464,N_44589);
or U46031 (N_46031,N_44927,N_44720);
and U46032 (N_46032,N_44615,N_44095);
or U46033 (N_46033,N_45522,N_45486);
nor U46034 (N_46034,N_44517,N_44655);
and U46035 (N_46035,N_44656,N_44502);
nand U46036 (N_46036,N_44319,N_44638);
or U46037 (N_46037,N_44028,N_45444);
nor U46038 (N_46038,N_45770,N_44382);
nand U46039 (N_46039,N_45178,N_44357);
and U46040 (N_46040,N_45577,N_44837);
nand U46041 (N_46041,N_44206,N_44344);
and U46042 (N_46042,N_45735,N_44981);
nor U46043 (N_46043,N_44566,N_44178);
and U46044 (N_46044,N_44957,N_45611);
nand U46045 (N_46045,N_45674,N_45473);
xnor U46046 (N_46046,N_44932,N_45049);
xor U46047 (N_46047,N_45549,N_44763);
and U46048 (N_46048,N_45928,N_44598);
or U46049 (N_46049,N_44113,N_45306);
nand U46050 (N_46050,N_44419,N_45937);
xnor U46051 (N_46051,N_44930,N_45076);
nor U46052 (N_46052,N_45181,N_45524);
xor U46053 (N_46053,N_45075,N_44340);
nand U46054 (N_46054,N_45580,N_45109);
xnor U46055 (N_46055,N_44512,N_45395);
nand U46056 (N_46056,N_45677,N_44918);
nor U46057 (N_46057,N_45279,N_45853);
nor U46058 (N_46058,N_45010,N_45746);
xnor U46059 (N_46059,N_45361,N_45933);
xnor U46060 (N_46060,N_44282,N_44739);
or U46061 (N_46061,N_45218,N_45123);
nand U46062 (N_46062,N_45833,N_45943);
and U46063 (N_46063,N_44366,N_44704);
nor U46064 (N_46064,N_44457,N_44016);
nor U46065 (N_46065,N_44067,N_44899);
nor U46066 (N_46066,N_44728,N_44423);
nor U46067 (N_46067,N_44752,N_45601);
nor U46068 (N_46068,N_45285,N_45965);
or U46069 (N_46069,N_44904,N_45573);
nand U46070 (N_46070,N_44624,N_45160);
nand U46071 (N_46071,N_45861,N_45213);
and U46072 (N_46072,N_44498,N_44325);
or U46073 (N_46073,N_44943,N_45307);
nand U46074 (N_46074,N_44793,N_45531);
and U46075 (N_46075,N_45507,N_44189);
nand U46076 (N_46076,N_44557,N_44259);
nand U46077 (N_46077,N_44926,N_45238);
or U46078 (N_46078,N_44052,N_45958);
or U46079 (N_46079,N_44249,N_45257);
nor U46080 (N_46080,N_44761,N_45461);
and U46081 (N_46081,N_44649,N_45192);
and U46082 (N_46082,N_45679,N_44785);
nor U46083 (N_46083,N_44315,N_44160);
and U46084 (N_46084,N_45025,N_45617);
xnor U46085 (N_46085,N_45276,N_45024);
nand U46086 (N_46086,N_44891,N_44645);
nand U46087 (N_46087,N_44542,N_45998);
or U46088 (N_46088,N_45216,N_45173);
or U46089 (N_46089,N_44768,N_45650);
and U46090 (N_46090,N_45868,N_44617);
nor U46091 (N_46091,N_44980,N_44609);
and U46092 (N_46092,N_45636,N_44717);
or U46093 (N_46093,N_45744,N_45835);
xnor U46094 (N_46094,N_45858,N_45530);
and U46095 (N_46095,N_45505,N_44778);
and U46096 (N_46096,N_45996,N_45825);
or U46097 (N_46097,N_44786,N_44080);
or U46098 (N_46098,N_44652,N_44553);
and U46099 (N_46099,N_44062,N_44706);
xnor U46100 (N_46100,N_44909,N_44292);
xnor U46101 (N_46101,N_44623,N_44529);
or U46102 (N_46102,N_44724,N_44789);
xor U46103 (N_46103,N_44022,N_45603);
nand U46104 (N_46104,N_45250,N_44523);
and U46105 (N_46105,N_44616,N_45260);
xnor U46106 (N_46106,N_45448,N_44476);
xor U46107 (N_46107,N_44222,N_45890);
nand U46108 (N_46108,N_44039,N_44925);
nor U46109 (N_46109,N_44363,N_45502);
and U46110 (N_46110,N_44865,N_44228);
or U46111 (N_46111,N_44477,N_45443);
and U46112 (N_46112,N_45424,N_45956);
nand U46113 (N_46113,N_45938,N_45102);
xnor U46114 (N_46114,N_45813,N_44684);
nor U46115 (N_46115,N_44966,N_44760);
or U46116 (N_46116,N_45392,N_44238);
xnor U46117 (N_46117,N_45380,N_44077);
nor U46118 (N_46118,N_45869,N_44479);
and U46119 (N_46119,N_44870,N_45815);
or U46120 (N_46120,N_44261,N_45117);
nand U46121 (N_46121,N_44337,N_45204);
nor U46122 (N_46122,N_45511,N_44103);
nand U46123 (N_46123,N_44569,N_45994);
or U46124 (N_46124,N_45856,N_45264);
or U46125 (N_46125,N_44318,N_45005);
and U46126 (N_46126,N_44141,N_44467);
or U46127 (N_46127,N_45949,N_45586);
and U46128 (N_46128,N_45757,N_44956);
xnor U46129 (N_46129,N_44443,N_44678);
nand U46130 (N_46130,N_45168,N_45312);
nand U46131 (N_46131,N_45565,N_44412);
nor U46132 (N_46132,N_44910,N_45261);
xor U46133 (N_46133,N_45594,N_44205);
nor U46134 (N_46134,N_45842,N_44465);
nand U46135 (N_46135,N_45170,N_44765);
nor U46136 (N_46136,N_45644,N_44844);
xor U46137 (N_46137,N_44592,N_44014);
and U46138 (N_46138,N_44688,N_44312);
xnor U46139 (N_46139,N_44025,N_44573);
xor U46140 (N_46140,N_45128,N_44440);
nor U46141 (N_46141,N_44499,N_45655);
nand U46142 (N_46142,N_44667,N_45692);
nand U46143 (N_46143,N_44223,N_44164);
nand U46144 (N_46144,N_44612,N_44952);
nor U46145 (N_46145,N_45660,N_44683);
or U46146 (N_46146,N_44845,N_44829);
nand U46147 (N_46147,N_45280,N_44579);
xor U46148 (N_46148,N_44431,N_44801);
nand U46149 (N_46149,N_45161,N_45789);
nor U46150 (N_46150,N_44977,N_45436);
or U46151 (N_46151,N_45955,N_45387);
nor U46152 (N_46152,N_44816,N_45232);
nor U46153 (N_46153,N_45051,N_44076);
nor U46154 (N_46154,N_45935,N_44203);
nor U46155 (N_46155,N_45923,N_45807);
and U46156 (N_46156,N_45990,N_45834);
and U46157 (N_46157,N_45959,N_44386);
nor U46158 (N_46158,N_44730,N_45050);
nand U46159 (N_46159,N_44729,N_44610);
and U46160 (N_46160,N_45985,N_45341);
or U46161 (N_46161,N_44438,N_44533);
or U46162 (N_46162,N_44577,N_44003);
xor U46163 (N_46163,N_45445,N_45184);
and U46164 (N_46164,N_45925,N_44286);
and U46165 (N_46165,N_44663,N_45014);
xor U46166 (N_46166,N_45018,N_45292);
or U46167 (N_46167,N_44453,N_44371);
nand U46168 (N_46168,N_45367,N_45801);
nand U46169 (N_46169,N_45590,N_45403);
and U46170 (N_46170,N_44716,N_45666);
xor U46171 (N_46171,N_45084,N_45780);
nor U46172 (N_46172,N_45402,N_44736);
xnor U46173 (N_46173,N_45163,N_44660);
nand U46174 (N_46174,N_45086,N_45417);
nand U46175 (N_46175,N_44965,N_44284);
nor U46176 (N_46176,N_45969,N_45855);
xnor U46177 (N_46177,N_45215,N_45224);
or U46178 (N_46178,N_45912,N_44177);
or U46179 (N_46179,N_44063,N_44381);
nand U46180 (N_46180,N_44804,N_45895);
nand U46181 (N_46181,N_44890,N_44416);
and U46182 (N_46182,N_44576,N_45887);
nor U46183 (N_46183,N_45645,N_44964);
or U46184 (N_46184,N_45962,N_44470);
and U46185 (N_46185,N_45680,N_45840);
xor U46186 (N_46186,N_45496,N_45251);
xor U46187 (N_46187,N_45122,N_45922);
or U46188 (N_46188,N_45305,N_44023);
or U46189 (N_46189,N_44575,N_45769);
xor U46190 (N_46190,N_45140,N_44169);
and U46191 (N_46191,N_44859,N_44634);
or U46192 (N_46192,N_44586,N_45519);
or U46193 (N_46193,N_45210,N_44931);
nand U46194 (N_46194,N_45262,N_45850);
nor U46195 (N_46195,N_45981,N_45695);
and U46196 (N_46196,N_44600,N_45046);
or U46197 (N_46197,N_44570,N_45235);
nor U46198 (N_46198,N_44959,N_45973);
nand U46199 (N_46199,N_45609,N_45599);
nor U46200 (N_46200,N_45588,N_45429);
nand U46201 (N_46201,N_44506,N_45982);
or U46202 (N_46202,N_45489,N_44774);
nand U46203 (N_46203,N_45768,N_45670);
nand U46204 (N_46204,N_44661,N_44128);
nand U46205 (N_46205,N_45967,N_45564);
nor U46206 (N_46206,N_44005,N_44935);
or U46207 (N_46207,N_45635,N_45782);
nor U46208 (N_46208,N_44908,N_45960);
and U46209 (N_46209,N_45527,N_44524);
xor U46210 (N_46210,N_44807,N_44034);
xor U46211 (N_46211,N_45608,N_44539);
xnor U46212 (N_46212,N_44188,N_45309);
xor U46213 (N_46213,N_44434,N_44481);
xor U46214 (N_46214,N_45696,N_45072);
and U46215 (N_46215,N_44179,N_45910);
and U46216 (N_46216,N_45986,N_44187);
or U46217 (N_46217,N_45227,N_44469);
or U46218 (N_46218,N_45641,N_44691);
xnor U46219 (N_46219,N_44883,N_44496);
or U46220 (N_46220,N_44492,N_45333);
nor U46221 (N_46221,N_44218,N_44708);
xor U46222 (N_46222,N_45542,N_44798);
and U46223 (N_46223,N_45317,N_44547);
and U46224 (N_46224,N_45092,N_44480);
xnor U46225 (N_46225,N_44352,N_45849);
and U46226 (N_46226,N_45787,N_45797);
or U46227 (N_46227,N_45575,N_45353);
nor U46228 (N_46228,N_45777,N_44040);
xor U46229 (N_46229,N_44850,N_45371);
xnor U46230 (N_46230,N_45576,N_45711);
and U46231 (N_46231,N_44430,N_44613);
xor U46232 (N_46232,N_44146,N_44982);
and U46233 (N_46233,N_45195,N_45897);
and U46234 (N_46234,N_44920,N_45002);
and U46235 (N_46235,N_44420,N_45152);
or U46236 (N_46236,N_44990,N_44256);
nand U46237 (N_46237,N_44614,N_45115);
and U46238 (N_46238,N_44605,N_45303);
and U46239 (N_46239,N_45365,N_44647);
nor U46240 (N_46240,N_45906,N_45526);
xnor U46241 (N_46241,N_44162,N_45151);
or U46242 (N_46242,N_44210,N_44513);
nand U46243 (N_46243,N_44450,N_45085);
nor U46244 (N_46244,N_45009,N_45470);
xor U46245 (N_46245,N_45498,N_44889);
or U46246 (N_46246,N_45681,N_44050);
and U46247 (N_46247,N_45036,N_44670);
nand U46248 (N_46248,N_45785,N_45313);
and U46249 (N_46249,N_44822,N_45000);
nor U46250 (N_46250,N_45931,N_44299);
xnor U46251 (N_46251,N_44628,N_45182);
or U46252 (N_46252,N_44393,N_45598);
or U46253 (N_46253,N_45753,N_45438);
xor U46254 (N_46254,N_45093,N_44722);
xor U46255 (N_46255,N_44084,N_44936);
nor U46256 (N_46256,N_45703,N_45383);
or U46257 (N_46257,N_45664,N_45900);
and U46258 (N_46258,N_45625,N_44584);
and U46259 (N_46259,N_45662,N_44507);
and U46260 (N_46260,N_45675,N_45427);
nor U46261 (N_46261,N_45326,N_44175);
xnor U46262 (N_46262,N_45523,N_45037);
or U46263 (N_46263,N_44975,N_45569);
nor U46264 (N_46264,N_44365,N_44792);
xor U46265 (N_46265,N_44456,N_44407);
xor U46266 (N_46266,N_45832,N_44858);
or U46267 (N_46267,N_44929,N_44354);
and U46268 (N_46268,N_45108,N_45632);
xor U46269 (N_46269,N_44285,N_45125);
and U46270 (N_46270,N_44463,N_45039);
nor U46271 (N_46271,N_45841,N_45258);
and U46272 (N_46272,N_45447,N_44192);
and U46273 (N_46273,N_45784,N_44127);
and U46274 (N_46274,N_44995,N_45282);
and U46275 (N_46275,N_44820,N_45648);
and U46276 (N_46276,N_44305,N_44914);
xnor U46277 (N_46277,N_45284,N_45434);
nor U46278 (N_46278,N_44591,N_45691);
nand U46279 (N_46279,N_45754,N_45714);
nand U46280 (N_46280,N_45359,N_45439);
xnor U46281 (N_46281,N_44585,N_45764);
nand U46282 (N_46282,N_45916,N_45805);
nand U46283 (N_46283,N_44152,N_44979);
or U46284 (N_46284,N_45592,N_44255);
nor U46285 (N_46285,N_45765,N_44313);
and U46286 (N_46286,N_45492,N_44830);
nand U46287 (N_46287,N_44750,N_44818);
xor U46288 (N_46288,N_44385,N_44561);
nand U46289 (N_46289,N_44733,N_45175);
nand U46290 (N_46290,N_45449,N_45254);
or U46291 (N_46291,N_45022,N_44242);
and U46292 (N_46292,N_44648,N_45678);
or U46293 (N_46293,N_44008,N_45545);
xnor U46294 (N_46294,N_44881,N_44079);
or U46295 (N_46295,N_45042,N_44984);
nor U46296 (N_46296,N_44159,N_44073);
nor U46297 (N_46297,N_44071,N_45255);
or U46298 (N_46298,N_45126,N_44689);
or U46299 (N_46299,N_44847,N_45003);
xor U46300 (N_46300,N_44355,N_44239);
or U46301 (N_46301,N_45634,N_45288);
nor U46302 (N_46302,N_45487,N_45249);
nor U46303 (N_46303,N_44056,N_45297);
or U46304 (N_46304,N_44070,N_45459);
and U46305 (N_46305,N_45162,N_45624);
and U46306 (N_46306,N_44713,N_44633);
and U46307 (N_46307,N_44676,N_44358);
or U46308 (N_46308,N_44546,N_44986);
nand U46309 (N_46309,N_45325,N_44916);
xnor U46310 (N_46310,N_45363,N_44311);
nor U46311 (N_46311,N_45047,N_44596);
or U46312 (N_46312,N_45339,N_44963);
or U46313 (N_46313,N_45626,N_44049);
xnor U46314 (N_46314,N_45352,N_45147);
xor U46315 (N_46315,N_44642,N_45335);
nand U46316 (N_46316,N_45035,N_44342);
xnor U46317 (N_46317,N_44675,N_44126);
nand U46318 (N_46318,N_44595,N_44756);
nor U46319 (N_46319,N_44038,N_44769);
and U46320 (N_46320,N_44330,N_44424);
nand U46321 (N_46321,N_44452,N_45267);
nand U46322 (N_46322,N_44897,N_44702);
or U46323 (N_46323,N_44134,N_44636);
or U46324 (N_46324,N_44174,N_45389);
nor U46325 (N_46325,N_44270,N_45011);
nor U46326 (N_46326,N_44161,N_45171);
and U46327 (N_46327,N_45902,N_44644);
xor U46328 (N_46328,N_44211,N_45244);
nor U46329 (N_46329,N_44196,N_44738);
nor U46330 (N_46330,N_44226,N_45286);
and U46331 (N_46331,N_44182,N_45040);
nor U46332 (N_46332,N_45538,N_45368);
nor U46333 (N_46333,N_45847,N_45968);
nand U46334 (N_46334,N_44474,N_45242);
nor U46335 (N_46335,N_45587,N_44111);
or U46336 (N_46336,N_45766,N_44978);
nand U46337 (N_46337,N_45966,N_44762);
xnor U46338 (N_46338,N_45440,N_45778);
and U46339 (N_46339,N_44779,N_44306);
nand U46340 (N_46340,N_44216,N_45839);
or U46341 (N_46341,N_44402,N_44351);
or U46342 (N_46342,N_45506,N_44705);
nor U46343 (N_46343,N_45055,N_45773);
and U46344 (N_46344,N_44968,N_45205);
xnor U46345 (N_46345,N_44274,N_44398);
and U46346 (N_46346,N_44747,N_45709);
nand U46347 (N_46347,N_45667,N_44998);
nand U46348 (N_46348,N_45469,N_44940);
and U46349 (N_46349,N_44973,N_45038);
nor U46350 (N_46350,N_44171,N_44399);
nor U46351 (N_46351,N_44827,N_45831);
and U46352 (N_46352,N_45547,N_44905);
nand U46353 (N_46353,N_44537,N_45405);
nand U46354 (N_46354,N_45225,N_44603);
or U46355 (N_46355,N_44240,N_45408);
nor U46356 (N_46356,N_45062,N_44105);
nand U46357 (N_46357,N_44322,N_45026);
nor U46358 (N_46358,N_45426,N_44097);
or U46359 (N_46359,N_45907,N_45838);
or U46360 (N_46360,N_45993,N_45995);
or U46361 (N_46361,N_45030,N_44018);
and U46362 (N_46362,N_45722,N_44796);
nand U46363 (N_46363,N_44976,N_44461);
nor U46364 (N_46364,N_44404,N_44520);
nor U46365 (N_46365,N_44515,N_45957);
nand U46366 (N_46366,N_45324,N_44046);
or U46367 (N_46367,N_44157,N_44298);
nand U46368 (N_46368,N_45669,N_45300);
xnor U46369 (N_46369,N_44180,N_44031);
xnor U46370 (N_46370,N_45546,N_44626);
and U46371 (N_46371,N_44323,N_45658);
and U46372 (N_46372,N_44526,N_44362);
nand U46373 (N_46373,N_44999,N_45915);
xnor U46374 (N_46374,N_45615,N_45817);
xor U46375 (N_46375,N_44967,N_44301);
or U46376 (N_46376,N_44735,N_45442);
xnor U46377 (N_46377,N_44601,N_45478);
nand U46378 (N_46378,N_45087,N_45827);
nand U46379 (N_46379,N_45929,N_45795);
or U46380 (N_46380,N_44173,N_44266);
nand U46381 (N_46381,N_44780,N_44848);
or U46382 (N_46382,N_44597,N_44823);
or U46383 (N_46383,N_44725,N_45471);
or U46384 (N_46384,N_45953,N_45535);
nor U46385 (N_46385,N_45146,N_44484);
or U46386 (N_46386,N_45820,N_45865);
or U46387 (N_46387,N_45020,N_44225);
nand U46388 (N_46388,N_45734,N_44490);
nand U46389 (N_46389,N_45707,N_45863);
xnor U46390 (N_46390,N_45208,N_44587);
and U46391 (N_46391,N_44408,N_45950);
nand U46392 (N_46392,N_45373,N_44378);
or U46393 (N_46393,N_45846,N_44532);
nand U46394 (N_46394,N_44139,N_45023);
or U46395 (N_46395,N_44204,N_45548);
and U46396 (N_46396,N_44445,N_45316);
and U46397 (N_46397,N_44849,N_44941);
and U46398 (N_46398,N_45490,N_44446);
or U46399 (N_46399,N_44861,N_45268);
or U46400 (N_46400,N_45372,N_45344);
nor U46401 (N_46401,N_45630,N_45008);
nor U46402 (N_46402,N_45435,N_45245);
nand U46403 (N_46403,N_45762,N_44811);
nor U46404 (N_46404,N_45911,N_44168);
xor U46405 (N_46405,N_44458,N_45043);
nor U46406 (N_46406,N_45515,N_45089);
and U46407 (N_46407,N_44370,N_45314);
xor U46408 (N_46408,N_44232,N_44640);
nor U46409 (N_46409,N_45240,N_44133);
xor U46410 (N_46410,N_44621,N_45737);
or U46411 (N_46411,N_44074,N_44083);
nor U46412 (N_46412,N_44380,N_44685);
or U46413 (N_46413,N_45829,N_45493);
nor U46414 (N_46414,N_45918,N_45059);
xor U46415 (N_46415,N_44950,N_45885);
and U46416 (N_46416,N_45243,N_45407);
and U46417 (N_46417,N_45256,N_44972);
or U46418 (N_46418,N_44607,N_45338);
xnor U46419 (N_46419,N_45759,N_44078);
or U46420 (N_46420,N_44391,N_45909);
or U46421 (N_46421,N_45673,N_45068);
xnor U46422 (N_46422,N_44740,N_45697);
nor U46423 (N_46423,N_44483,N_45143);
or U46424 (N_46424,N_45551,N_44277);
nand U46425 (N_46425,N_44921,N_44214);
nand U46426 (N_46426,N_45891,N_45396);
or U46427 (N_46427,N_45639,N_44015);
or U46428 (N_46428,N_44686,N_44158);
nor U46429 (N_46429,N_45428,N_45920);
or U46430 (N_46430,N_44749,N_45141);
or U46431 (N_46431,N_44772,N_44123);
xor U46432 (N_46432,N_45378,N_45921);
nand U46433 (N_46433,N_44939,N_44703);
nand U46434 (N_46434,N_45088,N_45961);
nor U46435 (N_46435,N_44806,N_44061);
or U46436 (N_46436,N_45226,N_44665);
and U46437 (N_46437,N_44087,N_45366);
xnor U46438 (N_46438,N_44753,N_44369);
nand U46439 (N_46439,N_44207,N_45032);
nand U46440 (N_46440,N_45377,N_44876);
nor U46441 (N_46441,N_44275,N_44280);
nand U46442 (N_46442,N_44563,N_44448);
nor U46443 (N_46443,N_44013,N_45880);
xnor U46444 (N_46444,N_45804,N_44244);
xor U46445 (N_46445,N_44166,N_44554);
nand U46446 (N_46446,N_45246,N_45044);
and U46447 (N_46447,N_45823,N_44220);
nand U46448 (N_46448,N_44096,N_45977);
nor U46449 (N_46449,N_45200,N_45275);
or U46450 (N_46450,N_45934,N_45618);
or U46451 (N_46451,N_45582,N_45710);
or U46452 (N_46452,N_44521,N_45074);
nand U46453 (N_46453,N_44588,N_45570);
nand U46454 (N_46454,N_44948,N_45421);
and U46455 (N_46455,N_45975,N_44933);
nor U46456 (N_46456,N_44142,N_45239);
nand U46457 (N_46457,N_44383,N_44508);
or U46458 (N_46458,N_44267,N_45437);
nand U46459 (N_46459,N_45631,N_45179);
xnor U46460 (N_46460,N_45733,N_44287);
xor U46461 (N_46461,N_44020,N_44754);
xnor U46462 (N_46462,N_44599,N_45431);
xnor U46463 (N_46463,N_44264,N_44001);
or U46464 (N_46464,N_44938,N_44923);
nor U46465 (N_46465,N_45253,N_45241);
and U46466 (N_46466,N_45661,N_44864);
nor U46467 (N_46467,N_44934,N_45100);
and U46468 (N_46468,N_44217,N_44224);
nor U46469 (N_46469,N_45164,N_44012);
nor U46470 (N_46470,N_45413,N_45460);
nor U46471 (N_46471,N_44898,N_44843);
nor U46472 (N_46472,N_45533,N_44873);
nor U46473 (N_46473,N_44130,N_44880);
xor U46474 (N_46474,N_45984,N_44550);
or U46475 (N_46475,N_44482,N_44696);
or U46476 (N_46476,N_45001,N_44671);
or U46477 (N_46477,N_44574,N_44272);
nand U46478 (N_46478,N_44291,N_45554);
xor U46479 (N_46479,N_45864,N_45583);
nor U46480 (N_46480,N_44110,N_45881);
xnor U46481 (N_46481,N_44304,N_44233);
nor U46482 (N_46482,N_44854,N_44345);
xor U46483 (N_46483,N_44544,N_45796);
and U46484 (N_46484,N_45323,N_45124);
and U46485 (N_46485,N_44571,N_44118);
xor U46486 (N_46486,N_45057,N_45265);
xnor U46487 (N_46487,N_44622,N_44019);
xor U46488 (N_46488,N_44751,N_45504);
nand U46489 (N_46489,N_44121,N_45936);
and U46490 (N_46490,N_45016,N_45061);
xor U46491 (N_46491,N_44900,N_44122);
nor U46492 (N_46492,N_45400,N_45159);
and U46493 (N_46493,N_44698,N_44032);
or U46494 (N_46494,N_45153,N_45792);
nand U46495 (N_46495,N_45474,N_44755);
nand U46496 (N_46496,N_44359,N_44867);
nor U46497 (N_46497,N_45941,N_44758);
nand U46498 (N_46498,N_45563,N_45132);
nor U46499 (N_46499,N_45206,N_44697);
and U46500 (N_46500,N_44401,N_44856);
nor U46501 (N_46501,N_45786,N_44269);
xnor U46502 (N_46502,N_45099,N_45129);
or U46503 (N_46503,N_44006,N_45236);
or U46504 (N_46504,N_44803,N_44875);
and U46505 (N_46505,N_44472,N_44009);
nor U46506 (N_46506,N_45150,N_44568);
or U46507 (N_46507,N_44279,N_44428);
nor U46508 (N_46508,N_45561,N_45248);
and U46509 (N_46509,N_45376,N_45724);
xor U46510 (N_46510,N_45104,N_44403);
nor U46511 (N_46511,N_44872,N_45628);
nand U46512 (N_46512,N_45627,N_45203);
or U46513 (N_46513,N_44992,N_45391);
or U46514 (N_46514,N_45197,N_44788);
xor U46515 (N_46515,N_44148,N_44759);
nor U46516 (N_46516,N_45579,N_45555);
nand U46517 (N_46517,N_45116,N_45472);
xor U46518 (N_46518,N_44149,N_45690);
xnor U46519 (N_46519,N_45019,N_44527);
nor U46520 (N_46520,N_44593,N_45467);
and U46521 (N_46521,N_45451,N_45708);
or U46522 (N_46522,N_45476,N_44770);
nand U46523 (N_46523,N_44879,N_45940);
or U46524 (N_46524,N_44629,N_45081);
xnor U46525 (N_46525,N_44258,N_45514);
nand U46526 (N_46526,N_45388,N_45346);
nor U46527 (N_46527,N_45409,N_45557);
and U46528 (N_46528,N_44417,N_45188);
xnor U46529 (N_46529,N_45272,N_44602);
xnor U46530 (N_46530,N_44468,N_44027);
xor U46531 (N_46531,N_44326,N_44343);
nand U46532 (N_46532,N_44887,N_44518);
and U46533 (N_46533,N_45857,N_44783);
and U46534 (N_46534,N_45157,N_44666);
nor U46535 (N_46535,N_45550,N_45231);
or U46536 (N_46536,N_44246,N_45513);
nor U46537 (N_46537,N_44137,N_44580);
or U46538 (N_46538,N_44766,N_45144);
xor U46539 (N_46539,N_45620,N_45760);
or U46540 (N_46540,N_45390,N_44810);
and U46541 (N_46541,N_45070,N_44396);
or U46542 (N_46542,N_45462,N_44388);
and U46543 (N_46543,N_44449,N_44185);
nor U46544 (N_46544,N_44115,N_45774);
nor U46545 (N_46545,N_44338,N_44372);
or U46546 (N_46546,N_44497,N_44324);
nor U46547 (N_46547,N_44700,N_44278);
or U46548 (N_46548,N_45412,N_45930);
and U46549 (N_46549,N_45336,N_45458);
and U46550 (N_46550,N_45539,N_44119);
nand U46551 (N_46551,N_45277,N_45721);
nor U46552 (N_46552,N_44058,N_44748);
nor U46553 (N_46553,N_45494,N_45029);
or U46554 (N_46554,N_45337,N_45422);
xor U46555 (N_46555,N_44555,N_44088);
or U46556 (N_46556,N_45199,N_45607);
nor U46557 (N_46557,N_45154,N_45781);
or U46558 (N_46558,N_45481,N_44677);
and U46559 (N_46559,N_45657,N_45399);
nor U46560 (N_46560,N_45537,N_44007);
or U46561 (N_46561,N_44197,N_45616);
xor U46562 (N_46562,N_45191,N_45556);
nor U46563 (N_46563,N_44081,N_44066);
nand U46564 (N_46564,N_45614,N_45814);
nor U46565 (N_46565,N_45356,N_45954);
and U46566 (N_46566,N_44535,N_44030);
and U46567 (N_46567,N_44409,N_44290);
xor U46568 (N_46568,N_45113,N_45234);
and U46569 (N_46569,N_45802,N_45649);
and U46570 (N_46570,N_44131,N_45826);
xor U46571 (N_46571,N_44951,N_45198);
nand U46572 (N_46572,N_44243,N_45385);
nand U46573 (N_46573,N_45033,N_45712);
or U46574 (N_46574,N_44072,N_45379);
xnor U46575 (N_46575,N_45758,N_45223);
and U46576 (N_46576,N_44029,N_45135);
nand U46577 (N_46577,N_45193,N_45860);
nand U46578 (N_46578,N_44065,N_44627);
nor U46579 (N_46579,N_45738,N_45386);
xor U46580 (N_46580,N_44971,N_44021);
and U46581 (N_46581,N_45879,N_44726);
or U46582 (N_46582,N_45706,N_44392);
nand U46583 (N_46583,N_45844,N_44254);
and U46584 (N_46584,N_45393,N_45553);
or U46585 (N_46585,N_44799,N_44907);
nand U46586 (N_46586,N_45452,N_44945);
nand U46587 (N_46587,N_45158,N_45619);
or U46588 (N_46588,N_45091,N_45882);
nand U46589 (N_46589,N_44819,N_45134);
xnor U46590 (N_46590,N_44035,N_44501);
and U46591 (N_46591,N_45719,N_44495);
and U46592 (N_46592,N_44509,N_44731);
nor U46593 (N_46593,N_45340,N_45121);
xor U46594 (N_46594,N_44701,N_45988);
nor U46595 (N_46595,N_45873,N_45584);
or U46596 (N_46596,N_44485,N_45512);
xor U46597 (N_46597,N_45394,N_44737);
xor U46598 (N_46598,N_45717,N_45763);
nand U46599 (N_46599,N_45167,N_44106);
xnor U46600 (N_46600,N_45209,N_45034);
xor U46601 (N_46601,N_45843,N_45118);
or U46602 (N_46602,N_45334,N_44112);
xnor U46603 (N_46603,N_45836,N_44790);
and U46604 (N_46604,N_45327,N_45913);
nand U46605 (N_46605,N_45343,N_45252);
nor U46606 (N_46606,N_45596,N_44471);
and U46607 (N_46607,N_44549,N_44813);
nor U46608 (N_46608,N_45640,N_44619);
and U46609 (N_46609,N_44036,N_44252);
xor U46610 (N_46610,N_45228,N_44427);
nor U46611 (N_46611,N_45183,N_44917);
xor U46612 (N_46612,N_44988,N_45120);
nand U46613 (N_46613,N_44390,N_44209);
xor U46614 (N_46614,N_44309,N_44145);
nor U46615 (N_46615,N_44743,N_45687);
or U46616 (N_46616,N_44341,N_44459);
nor U46617 (N_46617,N_44718,N_44672);
nor U46618 (N_46618,N_45318,N_44247);
and U46619 (N_46619,N_45974,N_44505);
or U46620 (N_46620,N_45845,N_45430);
xor U46621 (N_46621,N_44208,N_45411);
nand U46622 (N_46622,N_45516,N_45979);
or U46623 (N_46623,N_44654,N_44650);
nor U46624 (N_46624,N_44831,N_45718);
nand U46625 (N_46625,N_44664,N_44776);
nor U46626 (N_46626,N_45745,N_44771);
nand U46627 (N_46627,N_44974,N_45012);
nor U46628 (N_46628,N_44727,N_44947);
nor U46629 (N_46629,N_44693,N_44153);
nor U46630 (N_46630,N_45971,N_45976);
and U46631 (N_46631,N_45852,N_45441);
and U46632 (N_46632,N_44397,N_45107);
nor U46633 (N_46633,N_44543,N_44384);
and U46634 (N_46634,N_45497,N_44098);
nand U46635 (N_46635,N_45942,N_44832);
nand U46636 (N_46636,N_45875,N_44912);
nor U46637 (N_46637,N_44886,N_44042);
nor U46638 (N_46638,N_44902,N_44635);
nand U46639 (N_46639,N_44987,N_45311);
xnor U46640 (N_46640,N_44389,N_45963);
xnor U46641 (N_46641,N_45063,N_44679);
nand U46642 (N_46642,N_45876,N_44333);
nor U46643 (N_46643,N_45006,N_44519);
xor U46644 (N_46644,N_44289,N_44565);
nand U46645 (N_46645,N_44682,N_44294);
or U46646 (N_46646,N_44415,N_44320);
nand U46647 (N_46647,N_44809,N_45806);
and U46648 (N_46648,N_44395,N_44946);
xor U46649 (N_46649,N_45810,N_45320);
nand U46650 (N_46650,N_45237,N_45767);
nand U46651 (N_46651,N_44332,N_45207);
and U46652 (N_46652,N_44882,N_45138);
nor U46653 (N_46653,N_45056,N_44406);
xnor U46654 (N_46654,N_44156,N_45349);
or U46655 (N_46655,N_45647,N_45382);
or U46656 (N_46656,N_44489,N_44002);
xnor U46657 (N_46657,N_45591,N_44486);
nand U46658 (N_46658,N_44690,N_45716);
and U46659 (N_46659,N_44314,N_44852);
nor U46660 (N_46660,N_44608,N_44347);
xnor U46661 (N_46661,N_44541,N_44410);
and U46662 (N_46662,N_44163,N_45214);
nor U46663 (N_46663,N_44564,N_45221);
and U46664 (N_46664,N_44464,N_45106);
or U46665 (N_46665,N_45488,N_45702);
nor U46666 (N_46666,N_45298,N_44567);
xor U46667 (N_46667,N_45069,N_45779);
xor U46668 (N_46668,N_44960,N_44212);
nor U46669 (N_46669,N_44268,N_44723);
or U46670 (N_46670,N_45790,N_44949);
xor U46671 (N_46671,N_45299,N_45828);
and U46672 (N_46672,N_45651,N_45822);
nand U46673 (N_46673,N_45137,N_45045);
nand U46674 (N_46674,N_45877,N_44488);
nand U46675 (N_46675,N_44841,N_45874);
nand U46676 (N_46676,N_44435,N_44017);
nor U46677 (N_46677,N_45211,N_45740);
nor U46678 (N_46678,N_45948,N_45871);
xnor U46679 (N_46679,N_45604,N_45397);
or U46680 (N_46680,N_44868,N_44924);
nor U46681 (N_46681,N_44316,N_44514);
and U46682 (N_46682,N_45079,N_44353);
or U46683 (N_46683,N_44432,N_45453);
or U46684 (N_46684,N_45800,N_44944);
xor U46685 (N_46685,N_44441,N_44194);
xor U46686 (N_46686,N_44138,N_45090);
or U46687 (N_46687,N_45720,N_44245);
nand U46688 (N_46688,N_45541,N_44114);
nor U46689 (N_46689,N_45987,N_44414);
nand U46690 (N_46690,N_44674,N_45263);
or U46691 (N_46691,N_44530,N_44170);
and U46692 (N_46692,N_45701,N_45525);
xor U46693 (N_46693,N_44504,N_45775);
nor U46694 (N_46694,N_44994,N_44540);
and U46695 (N_46695,N_45111,N_44104);
xor U46696 (N_46696,N_44694,N_44787);
and U46697 (N_46697,N_45133,N_44767);
or U46698 (N_46698,N_45585,N_45007);
or U46699 (N_46699,N_44082,N_44842);
nor U46700 (N_46700,N_45364,N_44895);
or U46701 (N_46701,N_44707,N_45621);
xnor U46702 (N_46702,N_44581,N_45904);
or U46703 (N_46703,N_44863,N_45886);
nand U46704 (N_46704,N_45156,N_45653);
or U46705 (N_46705,N_44795,N_45972);
or U46706 (N_46706,N_45521,N_44374);
and U46707 (N_46707,N_45015,N_45177);
xor U46708 (N_46708,N_44562,N_45713);
xnor U46709 (N_46709,N_45727,N_45892);
xor U46710 (N_46710,N_45686,N_44712);
and U46711 (N_46711,N_44885,N_45914);
xor U46712 (N_46712,N_44805,N_45612);
xor U46713 (N_46713,N_45872,N_44117);
nand U46714 (N_46714,N_45824,N_44651);
and U46715 (N_46715,N_44055,N_44777);
nand U46716 (N_46716,N_44336,N_45362);
or U46717 (N_46717,N_45559,N_45999);
nand U46718 (N_46718,N_44283,N_45301);
and U46719 (N_46719,N_45101,N_45058);
or U46720 (N_46720,N_45665,N_44797);
and U46721 (N_46721,N_45149,N_44375);
or U46722 (N_46722,N_45060,N_45704);
and U46723 (N_46723,N_44276,N_45495);
and U46724 (N_46724,N_45751,N_45819);
xor U46725 (N_46725,N_44181,N_45944);
nand U46726 (N_46726,N_44937,N_45747);
and U46727 (N_46727,N_44308,N_44583);
nor U46728 (N_46728,N_45351,N_45139);
nand U46729 (N_46729,N_45329,N_45041);
or U46730 (N_46730,N_45187,N_44100);
and U46731 (N_46731,N_45919,N_44201);
nor U46732 (N_46732,N_45552,N_45342);
xor U46733 (N_46733,N_45509,N_45520);
nand U46734 (N_46734,N_45233,N_44996);
xnor U46735 (N_46735,N_44687,N_44198);
nand U46736 (N_46736,N_44422,N_45694);
nand U46737 (N_46737,N_45862,N_45110);
nor U46738 (N_46738,N_44692,N_45155);
nand U46739 (N_46739,N_44360,N_44922);
nor U46740 (N_46740,N_45172,N_44411);
nor U46741 (N_46741,N_45321,N_45532);
and U46742 (N_46742,N_45031,N_45811);
nand U46743 (N_46743,N_44227,N_44154);
nor U46744 (N_46744,N_44120,N_44741);
xnor U46745 (N_46745,N_45726,N_44295);
or U46746 (N_46746,N_45283,N_45315);
nand U46747 (N_46747,N_44044,N_44293);
nor U46748 (N_46748,N_44710,N_45048);
nor U46749 (N_46749,N_44099,N_44913);
or U46750 (N_46750,N_44186,N_44089);
nand U46751 (N_46751,N_45004,N_45176);
nand U46752 (N_46752,N_45851,N_44376);
nand U46753 (N_46753,N_44680,N_44400);
and U46754 (N_46754,N_44840,N_44893);
and U46755 (N_46755,N_45883,N_45830);
xor U46756 (N_46756,N_44764,N_44715);
nand U46757 (N_46757,N_44136,N_44413);
or U46758 (N_46758,N_45878,N_45290);
or U46759 (N_46759,N_45053,N_44057);
xor U46760 (N_46760,N_45222,N_45278);
and U46761 (N_46761,N_45201,N_44473);
xor U46762 (N_46762,N_45230,N_45027);
nand U46763 (N_46763,N_44086,N_45078);
or U46764 (N_46764,N_45273,N_44503);
xnor U46765 (N_46765,N_44894,N_44172);
xor U46766 (N_46766,N_44611,N_44578);
or U46767 (N_46767,N_44281,N_45700);
and U46768 (N_46768,N_45748,N_45484);
nor U46769 (N_46769,N_45927,N_45859);
and U46770 (N_46770,N_44511,N_44888);
and U46771 (N_46771,N_44321,N_45866);
xnor U46772 (N_46772,N_44983,N_44637);
xnor U46773 (N_46773,N_45348,N_44200);
nand U46774 (N_46774,N_44229,N_44199);
xnor U46775 (N_46775,N_44625,N_45082);
or U46776 (N_46776,N_44202,N_45415);
or U46777 (N_46777,N_44433,N_45629);
and U46778 (N_46778,N_44455,N_45743);
nand U46779 (N_46779,N_45783,N_45997);
or U46780 (N_46780,N_45483,N_45127);
or U46781 (N_46781,N_45560,N_44781);
xor U46782 (N_46782,N_44884,N_45296);
nand U46783 (N_46783,N_44653,N_44919);
and U46784 (N_46784,N_44835,N_44699);
or U46785 (N_46785,N_45728,N_45350);
nand U46786 (N_46786,N_45593,N_44271);
or U46787 (N_46787,N_45568,N_45419);
nand U46788 (N_46788,N_45503,N_44439);
xnor U46789 (N_46789,N_45304,N_44193);
and U46790 (N_46790,N_44425,N_45098);
xor U46791 (N_46791,N_44426,N_45259);
nor U46792 (N_46792,N_44307,N_45270);
and U46793 (N_46793,N_44231,N_45951);
xor U46794 (N_46794,N_45212,N_45964);
or U46795 (N_46795,N_45656,N_44328);
or U46796 (N_46796,N_45269,N_44668);
nor U46797 (N_46797,N_45572,N_44190);
nand U46798 (N_46798,N_45463,N_44379);
nor U46799 (N_46799,N_45423,N_45404);
nor U46800 (N_46800,N_45903,N_45347);
nor U46801 (N_46801,N_45798,N_44147);
or U46802 (N_46802,N_44075,N_45889);
xnor U46803 (N_46803,N_44059,N_44551);
and U46804 (N_46804,N_44250,N_45723);
and U46805 (N_46805,N_45705,N_44460);
nor U46806 (N_46806,N_44522,N_45169);
nand U46807 (N_46807,N_45491,N_45698);
xnor U46808 (N_46808,N_44641,N_44010);
and U46809 (N_46809,N_44421,N_44033);
nor U46810 (N_46810,N_45073,N_44491);
xor U46811 (N_46811,N_45454,N_45788);
nand U46812 (N_46812,N_44855,N_45374);
nand U46813 (N_46813,N_45637,N_45540);
and U46814 (N_46814,N_44262,N_44744);
nor U46815 (N_46815,N_45741,N_44773);
nand U46816 (N_46816,N_44942,N_44348);
or U46817 (N_46817,N_45021,N_44361);
or U46818 (N_46818,N_45623,N_45054);
nor U46819 (N_46819,N_45932,N_44572);
and U46820 (N_46820,N_45668,N_45893);
nor U46821 (N_46821,N_44037,N_44051);
nor U46822 (N_46822,N_45689,N_45148);
nor U46823 (N_46823,N_44639,N_44838);
xor U46824 (N_46824,N_45185,N_44874);
nor U46825 (N_46825,N_44327,N_45190);
or U46826 (N_46826,N_44815,N_45414);
nor U46827 (N_46827,N_45633,N_44466);
and U46828 (N_46828,N_44437,N_44405);
xnor U46829 (N_46829,N_44297,N_44303);
nand U46830 (N_46830,N_45370,N_45752);
xnor U46831 (N_46831,N_45518,N_44828);
and U46832 (N_46832,N_45605,N_45529);
nor U46833 (N_46833,N_45812,N_44869);
nor U46834 (N_46834,N_44241,N_44263);
xnor U46835 (N_46835,N_45725,N_45544);
or U46836 (N_46836,N_45468,N_44043);
and U46837 (N_46837,N_44176,N_45736);
nand U46838 (N_46838,N_45715,N_44814);
nor U46839 (N_46839,N_45077,N_45685);
nor U46840 (N_46840,N_45870,N_44494);
or U46841 (N_46841,N_45600,N_44183);
xnor U46842 (N_46842,N_44090,N_44364);
or U46843 (N_46843,N_44132,N_44143);
xor U46844 (N_46844,N_45194,N_45799);
xnor U46845 (N_46845,N_44516,N_45457);
or U46846 (N_46846,N_45776,N_44782);
nor U46847 (N_46847,N_45980,N_44195);
nor U46848 (N_46848,N_44093,N_44054);
nand U46849 (N_46849,N_45166,N_45432);
or U46850 (N_46850,N_45064,N_44525);
nor U46851 (N_46851,N_45165,N_45808);
nand U46852 (N_46852,N_44116,N_44373);
or U46853 (N_46853,N_45477,N_45456);
and U46854 (N_46854,N_45096,N_44253);
nand U46855 (N_46855,N_45247,N_45848);
nand U46856 (N_46856,N_45646,N_45501);
or U46857 (N_46857,N_45699,N_45606);
xnor U46858 (N_46858,N_45136,N_45398);
xnor U46859 (N_46859,N_44356,N_45731);
xnor U46860 (N_46860,N_45693,N_44955);
and U46861 (N_46861,N_44124,N_44510);
nand U46862 (N_46862,N_44387,N_45578);
or U46863 (N_46863,N_44791,N_44296);
and U46864 (N_46864,N_44896,N_45947);
nor U46865 (N_46865,N_44534,N_44528);
xnor U46866 (N_46866,N_45103,N_45602);
or U46867 (N_46867,N_45528,N_44493);
xor U46868 (N_46868,N_44709,N_45581);
nor U46869 (N_46869,N_45358,N_44669);
xnor U46870 (N_46870,N_45749,N_44552);
or U46871 (N_46871,N_45671,N_45465);
or U46872 (N_46872,N_44094,N_45446);
nor U46873 (N_46873,N_44234,N_45683);
or U46874 (N_46874,N_45517,N_44346);
nor U46875 (N_46875,N_45418,N_45791);
nor U46876 (N_46876,N_44155,N_44350);
or U46877 (N_46877,N_45017,N_45425);
and U46878 (N_46878,N_44487,N_44331);
nand U46879 (N_46879,N_44004,N_45105);
nand U46880 (N_46880,N_45174,N_44901);
xnor U46881 (N_46881,N_45536,N_45369);
nand U46882 (N_46882,N_45071,N_44418);
nor U46883 (N_46883,N_44911,N_45202);
nor U46884 (N_46884,N_44462,N_44833);
and U46885 (N_46885,N_45375,N_44317);
xnor U46886 (N_46886,N_45319,N_44582);
xnor U46887 (N_46887,N_44604,N_45672);
or U46888 (N_46888,N_44590,N_44235);
nor U46889 (N_46889,N_44144,N_44368);
nand U46890 (N_46890,N_44367,N_44334);
xnor U46891 (N_46891,N_44825,N_45510);
nor U46892 (N_46892,N_45558,N_45066);
nor U46893 (N_46893,N_44024,N_44915);
or U46894 (N_46894,N_45939,N_45732);
or U46895 (N_46895,N_45901,N_44877);
or U46896 (N_46896,N_45485,N_44265);
and U46897 (N_46897,N_45908,N_45574);
xnor U46898 (N_46898,N_45186,N_45357);
xor U46899 (N_46899,N_45345,N_44742);
and U46900 (N_46900,N_45989,N_44681);
nor U46901 (N_46901,N_45331,N_44657);
nor U46902 (N_46902,N_45499,N_45189);
nand U46903 (N_46903,N_45180,N_45643);
and U46904 (N_46904,N_44794,N_45926);
xnor U46905 (N_46905,N_44451,N_44442);
xnor U46906 (N_46906,N_44892,N_45756);
nor U46907 (N_46907,N_45867,N_44129);
and U46908 (N_46908,N_45354,N_44060);
nor U46909 (N_46909,N_45295,N_45455);
xor U46910 (N_46910,N_45816,N_45381);
xnor U46911 (N_46911,N_44288,N_44993);
nand U46912 (N_46912,N_45642,N_45613);
nor U46913 (N_46913,N_45771,N_45854);
xor U46914 (N_46914,N_45401,N_45638);
xor U46915 (N_46915,N_44857,N_44821);
or U46916 (N_46916,N_44335,N_44851);
nor U46917 (N_46917,N_45217,N_44140);
nor U46918 (N_46918,N_44673,N_44302);
nor U46919 (N_46919,N_45730,N_44191);
or U46920 (N_46920,N_45266,N_45543);
or U46921 (N_46921,N_45028,N_44903);
or U46922 (N_46922,N_45610,N_45013);
and U46923 (N_46923,N_44048,N_44757);
or U46924 (N_46924,N_44092,N_45274);
nand U46925 (N_46925,N_45978,N_45970);
and U46926 (N_46926,N_45271,N_44560);
and U46927 (N_46927,N_44047,N_45761);
and U46928 (N_46928,N_44219,N_44800);
xor U46929 (N_46929,N_45739,N_45992);
nand U46930 (N_46930,N_45294,N_44606);
and U46931 (N_46931,N_44646,N_45281);
xor U46932 (N_46932,N_45080,N_45219);
nor U46933 (N_46933,N_44808,N_45905);
xnor U46934 (N_46934,N_44085,N_45595);
nor U46935 (N_46935,N_44041,N_45131);
nor U46936 (N_46936,N_45809,N_44436);
nor U46937 (N_46937,N_45818,N_45793);
nand U46938 (N_46938,N_44784,N_44871);
or U46939 (N_46939,N_45652,N_44478);
or U46940 (N_46940,N_45480,N_45597);
nand U46941 (N_46941,N_44711,N_45688);
nand U46942 (N_46942,N_45750,N_44221);
xnor U46943 (N_46943,N_44853,N_44531);
xor U46944 (N_46944,N_45308,N_45682);
or U46945 (N_46945,N_44826,N_44215);
or U46946 (N_46946,N_45229,N_44928);
nor U46947 (N_46947,N_44775,N_44091);
or U46948 (N_46948,N_44734,N_44836);
nor U46949 (N_46949,N_44444,N_45991);
and U46950 (N_46950,N_44802,N_44620);
xor U46951 (N_46951,N_45420,N_44817);
nand U46952 (N_46952,N_44300,N_44310);
nor U46953 (N_46953,N_44064,N_44053);
nor U46954 (N_46954,N_44069,N_44251);
and U46955 (N_46955,N_44906,N_45479);
xor U46956 (N_46956,N_45896,N_44349);
nor U46957 (N_46957,N_44447,N_45946);
nand U46958 (N_46958,N_45729,N_45466);
and U46959 (N_46959,N_44991,N_44125);
xnor U46960 (N_46960,N_45097,N_44339);
nand U46961 (N_46961,N_44237,N_45330);
xor U46962 (N_46962,N_44662,N_45220);
nor U46963 (N_46963,N_45663,N_45899);
xor U46964 (N_46964,N_45410,N_44108);
or U46965 (N_46965,N_44860,N_45302);
or U46966 (N_46966,N_45983,N_45114);
nand U46967 (N_46967,N_44454,N_45083);
or U46968 (N_46968,N_44862,N_45567);
nand U46969 (N_46969,N_44839,N_44230);
nand U46970 (N_46970,N_44165,N_44536);
nand U46971 (N_46971,N_44475,N_45052);
nor U46972 (N_46972,N_44962,N_44329);
nand U46973 (N_46973,N_45534,N_44834);
and U46974 (N_46974,N_44618,N_44632);
or U46975 (N_46975,N_44695,N_44970);
nand U46976 (N_46976,N_45119,N_44109);
nand U46977 (N_46977,N_45094,N_45095);
or U46978 (N_46978,N_44746,N_45589);
and U46979 (N_46979,N_45482,N_44151);
nand U46980 (N_46980,N_44394,N_45145);
nor U46981 (N_46981,N_44989,N_44658);
or U46982 (N_46982,N_45821,N_44000);
xnor U46983 (N_46983,N_44721,N_45772);
and U46984 (N_46984,N_44538,N_44260);
and U46985 (N_46985,N_44719,N_44213);
or U46986 (N_46986,N_45289,N_44150);
nand U46987 (N_46987,N_45803,N_45917);
nor U46988 (N_46988,N_44559,N_45794);
nor U46989 (N_46989,N_44107,N_45322);
xor U46990 (N_46990,N_45837,N_45888);
nor U46991 (N_46991,N_45676,N_44846);
nand U46992 (N_46992,N_45196,N_44236);
or U46993 (N_46993,N_44248,N_45112);
nand U46994 (N_46994,N_45065,N_44824);
xor U46995 (N_46995,N_45952,N_44545);
nand U46996 (N_46996,N_45654,N_45293);
xnor U46997 (N_46997,N_45755,N_44273);
nor U46998 (N_46998,N_44500,N_45562);
nor U46999 (N_46999,N_45924,N_44556);
or U47000 (N_47000,N_45888,N_44871);
nor U47001 (N_47001,N_45290,N_45916);
xnor U47002 (N_47002,N_44808,N_45605);
xor U47003 (N_47003,N_44836,N_45198);
nand U47004 (N_47004,N_45352,N_44716);
nand U47005 (N_47005,N_44967,N_45080);
nor U47006 (N_47006,N_44600,N_45325);
xor U47007 (N_47007,N_45018,N_44685);
and U47008 (N_47008,N_45717,N_45731);
and U47009 (N_47009,N_44972,N_44772);
xnor U47010 (N_47010,N_45322,N_45821);
xnor U47011 (N_47011,N_45738,N_44972);
or U47012 (N_47012,N_44275,N_45964);
or U47013 (N_47013,N_44748,N_44207);
nor U47014 (N_47014,N_45249,N_45447);
and U47015 (N_47015,N_45272,N_45264);
nor U47016 (N_47016,N_44108,N_45533);
or U47017 (N_47017,N_45790,N_45697);
nor U47018 (N_47018,N_45502,N_45974);
nor U47019 (N_47019,N_44456,N_45927);
nand U47020 (N_47020,N_44594,N_45985);
and U47021 (N_47021,N_45553,N_44263);
nor U47022 (N_47022,N_44419,N_44449);
or U47023 (N_47023,N_45386,N_44625);
xnor U47024 (N_47024,N_44637,N_44914);
or U47025 (N_47025,N_45985,N_45035);
nand U47026 (N_47026,N_45875,N_44413);
and U47027 (N_47027,N_44436,N_44320);
or U47028 (N_47028,N_44311,N_45292);
nand U47029 (N_47029,N_45150,N_45718);
nor U47030 (N_47030,N_45467,N_45078);
and U47031 (N_47031,N_44968,N_45295);
nand U47032 (N_47032,N_45447,N_44242);
and U47033 (N_47033,N_45271,N_45112);
xnor U47034 (N_47034,N_44639,N_45547);
nor U47035 (N_47035,N_45839,N_44580);
xor U47036 (N_47036,N_45418,N_45553);
nor U47037 (N_47037,N_44132,N_44322);
nand U47038 (N_47038,N_44625,N_44114);
nand U47039 (N_47039,N_45334,N_44011);
and U47040 (N_47040,N_45308,N_45649);
nand U47041 (N_47041,N_44374,N_44116);
nor U47042 (N_47042,N_44182,N_44297);
nand U47043 (N_47043,N_44819,N_44613);
and U47044 (N_47044,N_44812,N_44742);
and U47045 (N_47045,N_44235,N_44899);
nand U47046 (N_47046,N_45062,N_45434);
and U47047 (N_47047,N_45907,N_45209);
xnor U47048 (N_47048,N_45677,N_44882);
or U47049 (N_47049,N_44928,N_44090);
nand U47050 (N_47050,N_45575,N_44544);
nand U47051 (N_47051,N_45891,N_45249);
xnor U47052 (N_47052,N_45226,N_45137);
or U47053 (N_47053,N_44588,N_44975);
and U47054 (N_47054,N_44415,N_45247);
nand U47055 (N_47055,N_45752,N_44789);
and U47056 (N_47056,N_45827,N_45161);
nor U47057 (N_47057,N_44091,N_44444);
nand U47058 (N_47058,N_44661,N_45606);
nand U47059 (N_47059,N_44925,N_44432);
nand U47060 (N_47060,N_45851,N_44719);
and U47061 (N_47061,N_45271,N_45967);
nand U47062 (N_47062,N_44215,N_45585);
and U47063 (N_47063,N_45767,N_45953);
xnor U47064 (N_47064,N_44484,N_45942);
and U47065 (N_47065,N_44849,N_45408);
xor U47066 (N_47066,N_45506,N_44429);
nor U47067 (N_47067,N_44502,N_45668);
and U47068 (N_47068,N_45664,N_44052);
nand U47069 (N_47069,N_45959,N_44772);
or U47070 (N_47070,N_45292,N_44782);
or U47071 (N_47071,N_44212,N_44388);
nand U47072 (N_47072,N_45754,N_44013);
nand U47073 (N_47073,N_44734,N_44953);
and U47074 (N_47074,N_45147,N_44122);
or U47075 (N_47075,N_45570,N_44854);
or U47076 (N_47076,N_44630,N_44626);
nand U47077 (N_47077,N_44361,N_44551);
nor U47078 (N_47078,N_45995,N_45879);
nand U47079 (N_47079,N_44446,N_45472);
nor U47080 (N_47080,N_45142,N_45724);
nand U47081 (N_47081,N_45992,N_44401);
nand U47082 (N_47082,N_44972,N_45729);
and U47083 (N_47083,N_44520,N_44168);
xor U47084 (N_47084,N_45034,N_45765);
and U47085 (N_47085,N_44014,N_45354);
nor U47086 (N_47086,N_45154,N_45931);
and U47087 (N_47087,N_45540,N_45714);
nor U47088 (N_47088,N_45706,N_45489);
or U47089 (N_47089,N_45213,N_45346);
nand U47090 (N_47090,N_45483,N_45998);
nor U47091 (N_47091,N_45638,N_44835);
or U47092 (N_47092,N_44851,N_45310);
nand U47093 (N_47093,N_44693,N_45461);
xor U47094 (N_47094,N_45457,N_44541);
xnor U47095 (N_47095,N_45470,N_44418);
nand U47096 (N_47096,N_44873,N_45480);
or U47097 (N_47097,N_45313,N_44088);
or U47098 (N_47098,N_45388,N_45739);
xnor U47099 (N_47099,N_44478,N_45443);
nand U47100 (N_47100,N_45073,N_45461);
xor U47101 (N_47101,N_44373,N_44410);
and U47102 (N_47102,N_45187,N_44492);
or U47103 (N_47103,N_44761,N_45352);
nand U47104 (N_47104,N_45115,N_44097);
or U47105 (N_47105,N_44954,N_44573);
xnor U47106 (N_47106,N_44832,N_45506);
and U47107 (N_47107,N_44266,N_44196);
nor U47108 (N_47108,N_45570,N_44769);
or U47109 (N_47109,N_44087,N_44455);
and U47110 (N_47110,N_44642,N_45926);
nand U47111 (N_47111,N_44186,N_44246);
nand U47112 (N_47112,N_44118,N_44045);
nor U47113 (N_47113,N_45890,N_44323);
and U47114 (N_47114,N_45853,N_44668);
xor U47115 (N_47115,N_44183,N_45042);
xor U47116 (N_47116,N_45284,N_45325);
nor U47117 (N_47117,N_44132,N_45346);
or U47118 (N_47118,N_44825,N_45456);
nand U47119 (N_47119,N_44438,N_45165);
xnor U47120 (N_47120,N_44956,N_44041);
nand U47121 (N_47121,N_44701,N_45137);
nor U47122 (N_47122,N_45824,N_44415);
or U47123 (N_47123,N_44218,N_45075);
and U47124 (N_47124,N_45970,N_44742);
nor U47125 (N_47125,N_45253,N_45184);
nor U47126 (N_47126,N_45265,N_45559);
nand U47127 (N_47127,N_45080,N_44420);
nor U47128 (N_47128,N_44337,N_45014);
and U47129 (N_47129,N_44887,N_45997);
xnor U47130 (N_47130,N_45509,N_45929);
nor U47131 (N_47131,N_44925,N_45242);
nor U47132 (N_47132,N_44951,N_45106);
and U47133 (N_47133,N_45631,N_45415);
nor U47134 (N_47134,N_44597,N_45149);
and U47135 (N_47135,N_44601,N_44715);
xor U47136 (N_47136,N_44692,N_44127);
or U47137 (N_47137,N_45185,N_44361);
and U47138 (N_47138,N_45622,N_45858);
nor U47139 (N_47139,N_45436,N_44220);
and U47140 (N_47140,N_44603,N_44872);
nor U47141 (N_47141,N_45759,N_44089);
xnor U47142 (N_47142,N_44021,N_45636);
nand U47143 (N_47143,N_45893,N_44187);
or U47144 (N_47144,N_45099,N_45916);
or U47145 (N_47145,N_45888,N_44765);
and U47146 (N_47146,N_45571,N_45285);
nor U47147 (N_47147,N_44786,N_45705);
or U47148 (N_47148,N_44341,N_45788);
nor U47149 (N_47149,N_45564,N_45569);
nor U47150 (N_47150,N_45764,N_44126);
xnor U47151 (N_47151,N_45332,N_45162);
nand U47152 (N_47152,N_45569,N_45044);
and U47153 (N_47153,N_45308,N_45814);
xnor U47154 (N_47154,N_45672,N_44599);
nand U47155 (N_47155,N_45969,N_44136);
or U47156 (N_47156,N_44458,N_44183);
and U47157 (N_47157,N_45450,N_44439);
and U47158 (N_47158,N_44628,N_45838);
xnor U47159 (N_47159,N_44001,N_45698);
nand U47160 (N_47160,N_45914,N_44910);
nand U47161 (N_47161,N_44099,N_44478);
nor U47162 (N_47162,N_44369,N_45351);
nand U47163 (N_47163,N_45024,N_44925);
xnor U47164 (N_47164,N_44540,N_44314);
xnor U47165 (N_47165,N_44372,N_45311);
xnor U47166 (N_47166,N_44708,N_44762);
nor U47167 (N_47167,N_45415,N_44845);
and U47168 (N_47168,N_44650,N_45902);
nand U47169 (N_47169,N_45893,N_45843);
nor U47170 (N_47170,N_45094,N_44964);
xnor U47171 (N_47171,N_45930,N_45413);
and U47172 (N_47172,N_45626,N_45545);
nand U47173 (N_47173,N_44497,N_44272);
and U47174 (N_47174,N_45065,N_45337);
nor U47175 (N_47175,N_44697,N_44440);
and U47176 (N_47176,N_44817,N_45444);
xor U47177 (N_47177,N_45254,N_45598);
xor U47178 (N_47178,N_44334,N_44272);
and U47179 (N_47179,N_45348,N_44450);
nand U47180 (N_47180,N_44233,N_44826);
or U47181 (N_47181,N_45141,N_44720);
nand U47182 (N_47182,N_44014,N_45514);
and U47183 (N_47183,N_44613,N_45928);
nor U47184 (N_47184,N_44846,N_44397);
nor U47185 (N_47185,N_45999,N_45807);
nand U47186 (N_47186,N_44743,N_44181);
and U47187 (N_47187,N_45865,N_45065);
or U47188 (N_47188,N_45507,N_44203);
and U47189 (N_47189,N_45433,N_44237);
nand U47190 (N_47190,N_44961,N_45974);
nor U47191 (N_47191,N_44130,N_45508);
and U47192 (N_47192,N_44253,N_45141);
or U47193 (N_47193,N_45164,N_45783);
and U47194 (N_47194,N_44642,N_45529);
nor U47195 (N_47195,N_44385,N_44662);
and U47196 (N_47196,N_44580,N_45084);
xor U47197 (N_47197,N_45347,N_44128);
nand U47198 (N_47198,N_45347,N_45668);
xor U47199 (N_47199,N_45144,N_44632);
and U47200 (N_47200,N_45519,N_44557);
nor U47201 (N_47201,N_44216,N_45616);
or U47202 (N_47202,N_45646,N_45627);
xnor U47203 (N_47203,N_44566,N_44763);
nor U47204 (N_47204,N_45932,N_45206);
or U47205 (N_47205,N_45945,N_44908);
nor U47206 (N_47206,N_45334,N_45432);
nor U47207 (N_47207,N_45101,N_44683);
nand U47208 (N_47208,N_44412,N_44978);
or U47209 (N_47209,N_44765,N_44192);
nor U47210 (N_47210,N_45845,N_45729);
nor U47211 (N_47211,N_44755,N_45484);
xnor U47212 (N_47212,N_45118,N_45593);
and U47213 (N_47213,N_45701,N_45016);
xnor U47214 (N_47214,N_45033,N_44825);
nor U47215 (N_47215,N_44998,N_44235);
and U47216 (N_47216,N_44723,N_44814);
or U47217 (N_47217,N_44062,N_44541);
or U47218 (N_47218,N_45211,N_45981);
or U47219 (N_47219,N_45638,N_44357);
xor U47220 (N_47220,N_44102,N_44335);
or U47221 (N_47221,N_44495,N_44719);
nand U47222 (N_47222,N_44384,N_44885);
nand U47223 (N_47223,N_45776,N_44391);
and U47224 (N_47224,N_44325,N_44726);
xnor U47225 (N_47225,N_44312,N_44932);
or U47226 (N_47226,N_45756,N_45333);
or U47227 (N_47227,N_45019,N_44390);
and U47228 (N_47228,N_44549,N_44866);
nor U47229 (N_47229,N_44007,N_45436);
and U47230 (N_47230,N_45050,N_45703);
nor U47231 (N_47231,N_44832,N_44456);
and U47232 (N_47232,N_45693,N_44529);
nor U47233 (N_47233,N_45743,N_45646);
nand U47234 (N_47234,N_45162,N_44982);
nor U47235 (N_47235,N_44215,N_45590);
nand U47236 (N_47236,N_44940,N_44894);
or U47237 (N_47237,N_45750,N_45049);
nor U47238 (N_47238,N_45993,N_44522);
and U47239 (N_47239,N_44572,N_44594);
nand U47240 (N_47240,N_45024,N_44525);
nand U47241 (N_47241,N_44195,N_44834);
xor U47242 (N_47242,N_44616,N_45235);
or U47243 (N_47243,N_44025,N_45194);
nor U47244 (N_47244,N_45394,N_45563);
or U47245 (N_47245,N_45646,N_44258);
and U47246 (N_47246,N_45983,N_45643);
xnor U47247 (N_47247,N_44736,N_45469);
nand U47248 (N_47248,N_45972,N_44857);
nand U47249 (N_47249,N_44787,N_44092);
and U47250 (N_47250,N_44535,N_45167);
nor U47251 (N_47251,N_45249,N_45484);
nand U47252 (N_47252,N_45008,N_45548);
or U47253 (N_47253,N_44338,N_45298);
nor U47254 (N_47254,N_44910,N_45178);
or U47255 (N_47255,N_44387,N_45155);
xnor U47256 (N_47256,N_44796,N_45665);
and U47257 (N_47257,N_44730,N_45767);
nand U47258 (N_47258,N_44546,N_44978);
and U47259 (N_47259,N_44335,N_45912);
xnor U47260 (N_47260,N_45841,N_44753);
xor U47261 (N_47261,N_45795,N_45813);
xnor U47262 (N_47262,N_44731,N_44153);
nand U47263 (N_47263,N_45944,N_45221);
xnor U47264 (N_47264,N_45937,N_44452);
xor U47265 (N_47265,N_44373,N_44784);
or U47266 (N_47266,N_44079,N_44040);
nor U47267 (N_47267,N_45545,N_45161);
nand U47268 (N_47268,N_44414,N_45833);
and U47269 (N_47269,N_45612,N_45655);
or U47270 (N_47270,N_44598,N_44320);
or U47271 (N_47271,N_44293,N_45441);
or U47272 (N_47272,N_44962,N_44442);
nand U47273 (N_47273,N_45649,N_45192);
nor U47274 (N_47274,N_45232,N_45296);
xor U47275 (N_47275,N_45766,N_44775);
nand U47276 (N_47276,N_45544,N_44241);
and U47277 (N_47277,N_44137,N_44616);
nand U47278 (N_47278,N_45596,N_45100);
nand U47279 (N_47279,N_44740,N_45081);
and U47280 (N_47280,N_44574,N_44706);
or U47281 (N_47281,N_45167,N_44054);
xor U47282 (N_47282,N_44831,N_44162);
and U47283 (N_47283,N_45606,N_44284);
nand U47284 (N_47284,N_44032,N_44105);
nand U47285 (N_47285,N_45698,N_45997);
nand U47286 (N_47286,N_44116,N_44130);
xnor U47287 (N_47287,N_45291,N_44318);
nand U47288 (N_47288,N_45185,N_44902);
nand U47289 (N_47289,N_45040,N_45906);
nand U47290 (N_47290,N_45901,N_45032);
nand U47291 (N_47291,N_45723,N_45869);
nor U47292 (N_47292,N_44403,N_44824);
and U47293 (N_47293,N_45764,N_44845);
or U47294 (N_47294,N_45236,N_44023);
xor U47295 (N_47295,N_45377,N_45447);
xor U47296 (N_47296,N_45352,N_44814);
and U47297 (N_47297,N_45574,N_45382);
and U47298 (N_47298,N_44758,N_44131);
xnor U47299 (N_47299,N_45885,N_44596);
and U47300 (N_47300,N_44871,N_44989);
xnor U47301 (N_47301,N_45370,N_45418);
or U47302 (N_47302,N_44633,N_44144);
nand U47303 (N_47303,N_44759,N_44987);
or U47304 (N_47304,N_45141,N_45765);
and U47305 (N_47305,N_45605,N_45673);
nand U47306 (N_47306,N_44217,N_44685);
and U47307 (N_47307,N_44922,N_44296);
and U47308 (N_47308,N_44020,N_44044);
and U47309 (N_47309,N_45198,N_45854);
xnor U47310 (N_47310,N_44657,N_45577);
nand U47311 (N_47311,N_44231,N_45635);
or U47312 (N_47312,N_45938,N_45788);
nand U47313 (N_47313,N_44079,N_45463);
xnor U47314 (N_47314,N_44581,N_45413);
xor U47315 (N_47315,N_44001,N_44560);
or U47316 (N_47316,N_44001,N_45668);
and U47317 (N_47317,N_44036,N_45739);
or U47318 (N_47318,N_44908,N_45310);
xor U47319 (N_47319,N_44027,N_44036);
nor U47320 (N_47320,N_44432,N_44075);
nand U47321 (N_47321,N_44202,N_45232);
nor U47322 (N_47322,N_44243,N_44164);
xor U47323 (N_47323,N_45194,N_45481);
xor U47324 (N_47324,N_45741,N_45595);
xnor U47325 (N_47325,N_44946,N_44565);
or U47326 (N_47326,N_45097,N_44074);
xnor U47327 (N_47327,N_45279,N_44587);
or U47328 (N_47328,N_44382,N_45219);
or U47329 (N_47329,N_44815,N_45627);
nand U47330 (N_47330,N_45783,N_45565);
nand U47331 (N_47331,N_44622,N_45909);
nor U47332 (N_47332,N_45979,N_44928);
xnor U47333 (N_47333,N_45619,N_45074);
nor U47334 (N_47334,N_45052,N_45444);
nand U47335 (N_47335,N_45012,N_44953);
or U47336 (N_47336,N_45207,N_45027);
nor U47337 (N_47337,N_44872,N_44563);
nor U47338 (N_47338,N_44596,N_45247);
or U47339 (N_47339,N_45443,N_44922);
nor U47340 (N_47340,N_44096,N_44814);
and U47341 (N_47341,N_44150,N_45670);
nor U47342 (N_47342,N_45933,N_44676);
or U47343 (N_47343,N_44693,N_45204);
and U47344 (N_47344,N_44208,N_44407);
nand U47345 (N_47345,N_45833,N_44935);
or U47346 (N_47346,N_45230,N_45900);
or U47347 (N_47347,N_45017,N_44908);
nor U47348 (N_47348,N_45027,N_44732);
or U47349 (N_47349,N_45744,N_44508);
xnor U47350 (N_47350,N_44232,N_44500);
or U47351 (N_47351,N_44464,N_45198);
or U47352 (N_47352,N_45505,N_44817);
nand U47353 (N_47353,N_44831,N_45393);
nor U47354 (N_47354,N_44553,N_44780);
nand U47355 (N_47355,N_45696,N_45387);
and U47356 (N_47356,N_45928,N_45533);
nor U47357 (N_47357,N_44274,N_45850);
and U47358 (N_47358,N_44807,N_45807);
and U47359 (N_47359,N_44760,N_45196);
and U47360 (N_47360,N_44457,N_45582);
and U47361 (N_47361,N_45434,N_44717);
nor U47362 (N_47362,N_44081,N_44940);
nor U47363 (N_47363,N_44998,N_45456);
nand U47364 (N_47364,N_44483,N_45375);
and U47365 (N_47365,N_45506,N_44767);
nand U47366 (N_47366,N_44232,N_44913);
nand U47367 (N_47367,N_44824,N_45588);
nor U47368 (N_47368,N_45755,N_44114);
and U47369 (N_47369,N_45562,N_45787);
xor U47370 (N_47370,N_45466,N_44896);
and U47371 (N_47371,N_45860,N_44632);
or U47372 (N_47372,N_45504,N_45827);
or U47373 (N_47373,N_44430,N_44753);
nand U47374 (N_47374,N_45145,N_45930);
and U47375 (N_47375,N_44168,N_44523);
nor U47376 (N_47376,N_45465,N_44541);
and U47377 (N_47377,N_44860,N_44484);
and U47378 (N_47378,N_44095,N_44157);
nand U47379 (N_47379,N_45288,N_45975);
nand U47380 (N_47380,N_45501,N_44963);
nor U47381 (N_47381,N_45884,N_45490);
xor U47382 (N_47382,N_45903,N_44174);
xor U47383 (N_47383,N_45075,N_45324);
and U47384 (N_47384,N_44073,N_44549);
nor U47385 (N_47385,N_45043,N_45246);
nor U47386 (N_47386,N_44716,N_44724);
and U47387 (N_47387,N_44127,N_44990);
nand U47388 (N_47388,N_45194,N_45253);
nand U47389 (N_47389,N_44282,N_45322);
nor U47390 (N_47390,N_44104,N_45700);
and U47391 (N_47391,N_44467,N_45180);
nand U47392 (N_47392,N_44533,N_44727);
and U47393 (N_47393,N_45030,N_44592);
nand U47394 (N_47394,N_44513,N_44946);
nor U47395 (N_47395,N_44978,N_44257);
nand U47396 (N_47396,N_45865,N_44171);
nand U47397 (N_47397,N_45591,N_45499);
xor U47398 (N_47398,N_45794,N_44939);
nand U47399 (N_47399,N_44204,N_45509);
nand U47400 (N_47400,N_45365,N_44236);
xnor U47401 (N_47401,N_44187,N_44262);
nand U47402 (N_47402,N_44534,N_44485);
and U47403 (N_47403,N_45433,N_44958);
or U47404 (N_47404,N_45605,N_44444);
nor U47405 (N_47405,N_44797,N_45321);
nor U47406 (N_47406,N_44848,N_45631);
and U47407 (N_47407,N_44257,N_45327);
and U47408 (N_47408,N_44193,N_45182);
nor U47409 (N_47409,N_44094,N_44447);
or U47410 (N_47410,N_45035,N_45031);
nor U47411 (N_47411,N_45467,N_45223);
nor U47412 (N_47412,N_44062,N_45528);
nand U47413 (N_47413,N_45309,N_44295);
nor U47414 (N_47414,N_45974,N_45086);
nand U47415 (N_47415,N_45802,N_44575);
xor U47416 (N_47416,N_45182,N_45240);
xor U47417 (N_47417,N_45875,N_44445);
and U47418 (N_47418,N_45792,N_45612);
or U47419 (N_47419,N_45892,N_45035);
nor U47420 (N_47420,N_45253,N_45100);
nand U47421 (N_47421,N_45384,N_45093);
xor U47422 (N_47422,N_44778,N_44930);
or U47423 (N_47423,N_45817,N_44922);
xor U47424 (N_47424,N_44475,N_44358);
nand U47425 (N_47425,N_45140,N_45717);
and U47426 (N_47426,N_44414,N_45048);
nor U47427 (N_47427,N_44679,N_44482);
or U47428 (N_47428,N_44266,N_45356);
and U47429 (N_47429,N_44807,N_44768);
xor U47430 (N_47430,N_44070,N_44614);
xnor U47431 (N_47431,N_45986,N_45522);
or U47432 (N_47432,N_44628,N_45436);
nand U47433 (N_47433,N_44353,N_45878);
nor U47434 (N_47434,N_45876,N_44436);
xnor U47435 (N_47435,N_44643,N_45042);
and U47436 (N_47436,N_44943,N_44096);
nor U47437 (N_47437,N_45168,N_44425);
xor U47438 (N_47438,N_44279,N_44952);
nor U47439 (N_47439,N_45949,N_45964);
xnor U47440 (N_47440,N_44193,N_45895);
xnor U47441 (N_47441,N_44732,N_44001);
nor U47442 (N_47442,N_45829,N_45133);
or U47443 (N_47443,N_45365,N_44933);
nand U47444 (N_47444,N_44340,N_44967);
and U47445 (N_47445,N_44523,N_45590);
nor U47446 (N_47446,N_44699,N_44175);
nand U47447 (N_47447,N_44148,N_45267);
nand U47448 (N_47448,N_44920,N_45989);
xor U47449 (N_47449,N_45710,N_45410);
xor U47450 (N_47450,N_45129,N_44302);
nor U47451 (N_47451,N_45794,N_44482);
nand U47452 (N_47452,N_44501,N_44277);
or U47453 (N_47453,N_44609,N_45366);
nor U47454 (N_47454,N_45045,N_45251);
and U47455 (N_47455,N_45761,N_44505);
xnor U47456 (N_47456,N_44479,N_44548);
nand U47457 (N_47457,N_44178,N_45404);
nor U47458 (N_47458,N_44494,N_44676);
and U47459 (N_47459,N_45765,N_44053);
and U47460 (N_47460,N_45676,N_44977);
nor U47461 (N_47461,N_44898,N_44600);
nand U47462 (N_47462,N_45480,N_45687);
nor U47463 (N_47463,N_45074,N_45043);
and U47464 (N_47464,N_44986,N_45877);
nand U47465 (N_47465,N_44223,N_44820);
xnor U47466 (N_47466,N_45689,N_44580);
nor U47467 (N_47467,N_45558,N_44274);
nor U47468 (N_47468,N_44073,N_45896);
or U47469 (N_47469,N_44123,N_44352);
nand U47470 (N_47470,N_44628,N_44870);
xor U47471 (N_47471,N_45570,N_45663);
and U47472 (N_47472,N_44343,N_45124);
or U47473 (N_47473,N_45406,N_45641);
nand U47474 (N_47474,N_44789,N_45179);
nand U47475 (N_47475,N_44388,N_45688);
or U47476 (N_47476,N_44817,N_45924);
nor U47477 (N_47477,N_45203,N_45098);
and U47478 (N_47478,N_44588,N_45630);
nor U47479 (N_47479,N_45941,N_44908);
nor U47480 (N_47480,N_44020,N_44239);
and U47481 (N_47481,N_44516,N_44118);
xnor U47482 (N_47482,N_44374,N_45175);
xnor U47483 (N_47483,N_44902,N_44155);
or U47484 (N_47484,N_45278,N_44739);
or U47485 (N_47485,N_45981,N_44346);
nor U47486 (N_47486,N_45182,N_45017);
xor U47487 (N_47487,N_45732,N_45415);
or U47488 (N_47488,N_45045,N_45628);
or U47489 (N_47489,N_45283,N_45178);
or U47490 (N_47490,N_45848,N_44264);
or U47491 (N_47491,N_44156,N_44398);
nand U47492 (N_47492,N_45135,N_45131);
or U47493 (N_47493,N_45349,N_45185);
nor U47494 (N_47494,N_45596,N_45297);
xor U47495 (N_47495,N_44735,N_44221);
and U47496 (N_47496,N_44653,N_44405);
or U47497 (N_47497,N_45173,N_44452);
or U47498 (N_47498,N_45643,N_45314);
or U47499 (N_47499,N_44335,N_44040);
and U47500 (N_47500,N_44914,N_45298);
and U47501 (N_47501,N_45684,N_45852);
nor U47502 (N_47502,N_44445,N_44077);
or U47503 (N_47503,N_44826,N_44428);
xnor U47504 (N_47504,N_45432,N_45506);
or U47505 (N_47505,N_44386,N_44623);
and U47506 (N_47506,N_44733,N_44013);
nand U47507 (N_47507,N_45535,N_45494);
and U47508 (N_47508,N_45131,N_44126);
and U47509 (N_47509,N_44485,N_45780);
nor U47510 (N_47510,N_44963,N_44928);
xnor U47511 (N_47511,N_44522,N_45038);
and U47512 (N_47512,N_44402,N_45000);
and U47513 (N_47513,N_45339,N_45571);
xor U47514 (N_47514,N_44340,N_45646);
and U47515 (N_47515,N_44733,N_45305);
or U47516 (N_47516,N_44527,N_44812);
nor U47517 (N_47517,N_45382,N_45204);
nor U47518 (N_47518,N_45312,N_44946);
and U47519 (N_47519,N_44415,N_45883);
xnor U47520 (N_47520,N_44694,N_44399);
and U47521 (N_47521,N_45808,N_44881);
or U47522 (N_47522,N_44444,N_45192);
nand U47523 (N_47523,N_45964,N_45539);
nand U47524 (N_47524,N_44519,N_44513);
or U47525 (N_47525,N_45206,N_45703);
and U47526 (N_47526,N_45802,N_44171);
xor U47527 (N_47527,N_45257,N_45595);
nand U47528 (N_47528,N_44071,N_44124);
or U47529 (N_47529,N_45508,N_45810);
and U47530 (N_47530,N_44051,N_45493);
xnor U47531 (N_47531,N_44871,N_45494);
xnor U47532 (N_47532,N_45578,N_45689);
and U47533 (N_47533,N_45568,N_44775);
nor U47534 (N_47534,N_44944,N_45668);
or U47535 (N_47535,N_45252,N_45987);
nand U47536 (N_47536,N_45853,N_45803);
xnor U47537 (N_47537,N_45057,N_44161);
nor U47538 (N_47538,N_44949,N_45584);
nand U47539 (N_47539,N_45840,N_44630);
xnor U47540 (N_47540,N_44685,N_44409);
and U47541 (N_47541,N_45575,N_45473);
xor U47542 (N_47542,N_45230,N_45431);
xor U47543 (N_47543,N_44029,N_44203);
or U47544 (N_47544,N_45101,N_45423);
or U47545 (N_47545,N_45330,N_45352);
nand U47546 (N_47546,N_44601,N_45551);
xor U47547 (N_47547,N_44331,N_44697);
and U47548 (N_47548,N_44772,N_45909);
xnor U47549 (N_47549,N_44477,N_45440);
nor U47550 (N_47550,N_44097,N_45938);
nand U47551 (N_47551,N_44921,N_44869);
nor U47552 (N_47552,N_45632,N_45444);
nor U47553 (N_47553,N_44795,N_44222);
or U47554 (N_47554,N_45095,N_44102);
nor U47555 (N_47555,N_44406,N_45702);
xor U47556 (N_47556,N_44044,N_44974);
nand U47557 (N_47557,N_44211,N_45067);
nor U47558 (N_47558,N_45373,N_45121);
or U47559 (N_47559,N_45702,N_44280);
or U47560 (N_47560,N_45566,N_44488);
nand U47561 (N_47561,N_44575,N_45455);
xor U47562 (N_47562,N_44436,N_44364);
and U47563 (N_47563,N_45045,N_44035);
xnor U47564 (N_47564,N_45267,N_44196);
and U47565 (N_47565,N_45122,N_44140);
nor U47566 (N_47566,N_45667,N_44828);
nand U47567 (N_47567,N_44913,N_45935);
and U47568 (N_47568,N_44100,N_44619);
nand U47569 (N_47569,N_44655,N_44665);
and U47570 (N_47570,N_45612,N_45920);
and U47571 (N_47571,N_45283,N_45489);
nand U47572 (N_47572,N_45599,N_44646);
nor U47573 (N_47573,N_45430,N_45389);
and U47574 (N_47574,N_45384,N_44108);
xor U47575 (N_47575,N_45371,N_44774);
nand U47576 (N_47576,N_44981,N_45300);
nor U47577 (N_47577,N_45172,N_44428);
nor U47578 (N_47578,N_44800,N_45943);
nor U47579 (N_47579,N_45055,N_44498);
and U47580 (N_47580,N_44109,N_45007);
or U47581 (N_47581,N_44622,N_45618);
nand U47582 (N_47582,N_45231,N_45988);
xor U47583 (N_47583,N_44840,N_45573);
or U47584 (N_47584,N_45488,N_45761);
nor U47585 (N_47585,N_44045,N_45095);
or U47586 (N_47586,N_45294,N_45590);
and U47587 (N_47587,N_45381,N_45476);
nor U47588 (N_47588,N_44363,N_45142);
xnor U47589 (N_47589,N_45042,N_44519);
or U47590 (N_47590,N_45100,N_44145);
and U47591 (N_47591,N_45349,N_44459);
and U47592 (N_47592,N_45033,N_44170);
nand U47593 (N_47593,N_45497,N_44024);
or U47594 (N_47594,N_45290,N_44235);
xnor U47595 (N_47595,N_44491,N_45451);
nand U47596 (N_47596,N_44337,N_44694);
nand U47597 (N_47597,N_45640,N_44033);
xnor U47598 (N_47598,N_44551,N_44115);
or U47599 (N_47599,N_45382,N_44902);
or U47600 (N_47600,N_44340,N_45303);
nor U47601 (N_47601,N_45402,N_44741);
or U47602 (N_47602,N_44409,N_45515);
or U47603 (N_47603,N_45377,N_44744);
nor U47604 (N_47604,N_45917,N_44459);
and U47605 (N_47605,N_44804,N_45977);
xor U47606 (N_47606,N_45449,N_44339);
and U47607 (N_47607,N_45982,N_44500);
nor U47608 (N_47608,N_45339,N_45104);
xor U47609 (N_47609,N_45004,N_45076);
xnor U47610 (N_47610,N_45600,N_45015);
nand U47611 (N_47611,N_44961,N_45634);
and U47612 (N_47612,N_45474,N_44920);
nand U47613 (N_47613,N_45348,N_45349);
xor U47614 (N_47614,N_44924,N_45367);
or U47615 (N_47615,N_45124,N_45585);
and U47616 (N_47616,N_44253,N_44234);
or U47617 (N_47617,N_45472,N_44175);
and U47618 (N_47618,N_44944,N_44345);
nand U47619 (N_47619,N_44002,N_44204);
or U47620 (N_47620,N_44470,N_44698);
or U47621 (N_47621,N_44713,N_45930);
nand U47622 (N_47622,N_44305,N_45262);
and U47623 (N_47623,N_45196,N_45604);
nand U47624 (N_47624,N_45696,N_44764);
nand U47625 (N_47625,N_45290,N_45864);
or U47626 (N_47626,N_44099,N_44335);
and U47627 (N_47627,N_45917,N_45530);
and U47628 (N_47628,N_45546,N_44993);
and U47629 (N_47629,N_45330,N_45647);
and U47630 (N_47630,N_44500,N_45824);
nor U47631 (N_47631,N_44433,N_44578);
nand U47632 (N_47632,N_44748,N_45970);
nor U47633 (N_47633,N_45860,N_45703);
nor U47634 (N_47634,N_44293,N_44509);
nor U47635 (N_47635,N_44193,N_45930);
or U47636 (N_47636,N_44635,N_44132);
xor U47637 (N_47637,N_44126,N_45251);
nor U47638 (N_47638,N_44051,N_44561);
or U47639 (N_47639,N_45993,N_45488);
xnor U47640 (N_47640,N_45145,N_44573);
nor U47641 (N_47641,N_45194,N_44928);
nor U47642 (N_47642,N_44638,N_44230);
xor U47643 (N_47643,N_44166,N_45535);
nor U47644 (N_47644,N_45893,N_44755);
xor U47645 (N_47645,N_45138,N_44981);
nor U47646 (N_47646,N_44340,N_44897);
xnor U47647 (N_47647,N_44008,N_45548);
nor U47648 (N_47648,N_45326,N_45277);
xor U47649 (N_47649,N_44537,N_44264);
xor U47650 (N_47650,N_44410,N_44636);
nor U47651 (N_47651,N_45029,N_44400);
and U47652 (N_47652,N_44753,N_45324);
nand U47653 (N_47653,N_44009,N_44101);
or U47654 (N_47654,N_45678,N_44713);
xnor U47655 (N_47655,N_44663,N_44535);
nand U47656 (N_47656,N_44802,N_44472);
xor U47657 (N_47657,N_45138,N_45241);
or U47658 (N_47658,N_44235,N_45943);
or U47659 (N_47659,N_44497,N_45076);
nor U47660 (N_47660,N_44423,N_45848);
and U47661 (N_47661,N_44270,N_45381);
xnor U47662 (N_47662,N_44253,N_45158);
nor U47663 (N_47663,N_45015,N_44545);
and U47664 (N_47664,N_44258,N_44086);
nand U47665 (N_47665,N_44246,N_44040);
xor U47666 (N_47666,N_44265,N_45019);
or U47667 (N_47667,N_44796,N_45739);
or U47668 (N_47668,N_44290,N_45674);
or U47669 (N_47669,N_44967,N_45369);
nor U47670 (N_47670,N_44783,N_45476);
xnor U47671 (N_47671,N_45551,N_44827);
or U47672 (N_47672,N_45258,N_45652);
nor U47673 (N_47673,N_44939,N_44459);
nor U47674 (N_47674,N_45177,N_45701);
nand U47675 (N_47675,N_45469,N_44357);
or U47676 (N_47676,N_45422,N_44658);
xnor U47677 (N_47677,N_44040,N_45930);
nand U47678 (N_47678,N_44588,N_44090);
nand U47679 (N_47679,N_45310,N_45321);
or U47680 (N_47680,N_45772,N_44705);
nor U47681 (N_47681,N_44194,N_44052);
or U47682 (N_47682,N_44825,N_45874);
xnor U47683 (N_47683,N_44488,N_44990);
and U47684 (N_47684,N_45072,N_44737);
nor U47685 (N_47685,N_44816,N_44221);
and U47686 (N_47686,N_45436,N_44120);
and U47687 (N_47687,N_45298,N_44461);
or U47688 (N_47688,N_45407,N_44887);
xnor U47689 (N_47689,N_45841,N_44014);
nor U47690 (N_47690,N_45341,N_44195);
xnor U47691 (N_47691,N_45161,N_44359);
or U47692 (N_47692,N_45004,N_45974);
or U47693 (N_47693,N_45208,N_45014);
and U47694 (N_47694,N_44290,N_45219);
or U47695 (N_47695,N_44233,N_45009);
xor U47696 (N_47696,N_45337,N_44243);
nand U47697 (N_47697,N_45528,N_44967);
xnor U47698 (N_47698,N_44857,N_45950);
xor U47699 (N_47699,N_44844,N_44427);
xor U47700 (N_47700,N_45368,N_45592);
nor U47701 (N_47701,N_44133,N_44045);
xnor U47702 (N_47702,N_44856,N_44627);
or U47703 (N_47703,N_45893,N_45760);
nor U47704 (N_47704,N_45560,N_44758);
xor U47705 (N_47705,N_44154,N_44344);
nor U47706 (N_47706,N_45653,N_45263);
nor U47707 (N_47707,N_45502,N_44310);
and U47708 (N_47708,N_45847,N_45732);
and U47709 (N_47709,N_45781,N_45799);
xor U47710 (N_47710,N_45229,N_44823);
xor U47711 (N_47711,N_44713,N_45182);
and U47712 (N_47712,N_44626,N_45275);
nor U47713 (N_47713,N_45527,N_44009);
xor U47714 (N_47714,N_44624,N_45897);
or U47715 (N_47715,N_44955,N_44251);
xor U47716 (N_47716,N_45783,N_44094);
xor U47717 (N_47717,N_44665,N_45359);
nor U47718 (N_47718,N_45178,N_45491);
xor U47719 (N_47719,N_44399,N_45320);
nand U47720 (N_47720,N_44337,N_44260);
nor U47721 (N_47721,N_44148,N_44244);
and U47722 (N_47722,N_44951,N_44830);
nor U47723 (N_47723,N_44827,N_44460);
xor U47724 (N_47724,N_45286,N_45431);
nor U47725 (N_47725,N_45480,N_44112);
or U47726 (N_47726,N_44440,N_44465);
or U47727 (N_47727,N_45835,N_44243);
nor U47728 (N_47728,N_44703,N_44689);
nand U47729 (N_47729,N_45344,N_44504);
nand U47730 (N_47730,N_45208,N_44306);
nand U47731 (N_47731,N_44740,N_45242);
and U47732 (N_47732,N_45570,N_44250);
nand U47733 (N_47733,N_45706,N_44749);
nor U47734 (N_47734,N_45511,N_44737);
nand U47735 (N_47735,N_45401,N_44852);
or U47736 (N_47736,N_44636,N_44507);
or U47737 (N_47737,N_44690,N_44309);
xor U47738 (N_47738,N_44254,N_45368);
or U47739 (N_47739,N_45903,N_44413);
or U47740 (N_47740,N_45736,N_45743);
nand U47741 (N_47741,N_45389,N_45254);
nand U47742 (N_47742,N_44461,N_45678);
and U47743 (N_47743,N_44675,N_45793);
nor U47744 (N_47744,N_45443,N_44297);
nor U47745 (N_47745,N_45141,N_44229);
xor U47746 (N_47746,N_45090,N_44314);
and U47747 (N_47747,N_44988,N_45200);
nand U47748 (N_47748,N_45571,N_44435);
nand U47749 (N_47749,N_44439,N_45022);
nor U47750 (N_47750,N_44937,N_45455);
nand U47751 (N_47751,N_45468,N_45131);
and U47752 (N_47752,N_45265,N_44936);
xor U47753 (N_47753,N_44954,N_45610);
or U47754 (N_47754,N_45835,N_44184);
nand U47755 (N_47755,N_44921,N_45702);
and U47756 (N_47756,N_44469,N_45214);
and U47757 (N_47757,N_45776,N_45671);
nor U47758 (N_47758,N_45067,N_44434);
nand U47759 (N_47759,N_45713,N_45758);
xnor U47760 (N_47760,N_45027,N_45091);
and U47761 (N_47761,N_45739,N_44802);
nand U47762 (N_47762,N_44434,N_44989);
xnor U47763 (N_47763,N_45135,N_45629);
or U47764 (N_47764,N_45054,N_45655);
and U47765 (N_47765,N_44927,N_45091);
or U47766 (N_47766,N_45294,N_44796);
or U47767 (N_47767,N_45098,N_45124);
nand U47768 (N_47768,N_44638,N_45663);
or U47769 (N_47769,N_44985,N_44686);
nor U47770 (N_47770,N_44146,N_45385);
nor U47771 (N_47771,N_44716,N_45096);
xor U47772 (N_47772,N_45178,N_45223);
xor U47773 (N_47773,N_44907,N_45389);
xnor U47774 (N_47774,N_45278,N_45092);
nand U47775 (N_47775,N_45441,N_44054);
nand U47776 (N_47776,N_45580,N_44109);
nand U47777 (N_47777,N_44045,N_44484);
and U47778 (N_47778,N_44870,N_45986);
nor U47779 (N_47779,N_44211,N_44033);
xnor U47780 (N_47780,N_44604,N_45099);
and U47781 (N_47781,N_44108,N_44770);
xor U47782 (N_47782,N_45150,N_44682);
nor U47783 (N_47783,N_44489,N_45134);
nand U47784 (N_47784,N_44800,N_44462);
xor U47785 (N_47785,N_44551,N_44946);
xor U47786 (N_47786,N_44749,N_45963);
nor U47787 (N_47787,N_44493,N_44868);
nand U47788 (N_47788,N_45328,N_44726);
nor U47789 (N_47789,N_45677,N_44366);
and U47790 (N_47790,N_44632,N_45553);
nand U47791 (N_47791,N_44774,N_44207);
and U47792 (N_47792,N_44151,N_44303);
and U47793 (N_47793,N_44834,N_45439);
or U47794 (N_47794,N_44660,N_44733);
xnor U47795 (N_47795,N_45933,N_44829);
or U47796 (N_47796,N_44609,N_45205);
nand U47797 (N_47797,N_44437,N_44471);
xnor U47798 (N_47798,N_45331,N_44879);
nor U47799 (N_47799,N_44293,N_45532);
nand U47800 (N_47800,N_45138,N_44441);
xnor U47801 (N_47801,N_45157,N_44899);
nor U47802 (N_47802,N_45300,N_44353);
nand U47803 (N_47803,N_44848,N_44337);
nor U47804 (N_47804,N_45858,N_45260);
and U47805 (N_47805,N_44552,N_45283);
nand U47806 (N_47806,N_44523,N_45312);
and U47807 (N_47807,N_45936,N_45069);
or U47808 (N_47808,N_44044,N_44118);
xor U47809 (N_47809,N_45656,N_44363);
nand U47810 (N_47810,N_44212,N_45389);
xor U47811 (N_47811,N_45676,N_45348);
nor U47812 (N_47812,N_44301,N_44243);
nand U47813 (N_47813,N_44249,N_44528);
nand U47814 (N_47814,N_45672,N_45749);
or U47815 (N_47815,N_44895,N_44749);
nor U47816 (N_47816,N_45526,N_45026);
and U47817 (N_47817,N_44162,N_45023);
nor U47818 (N_47818,N_44224,N_44160);
or U47819 (N_47819,N_44419,N_44152);
nor U47820 (N_47820,N_44824,N_45228);
or U47821 (N_47821,N_44691,N_45597);
or U47822 (N_47822,N_44376,N_45818);
nor U47823 (N_47823,N_44441,N_44229);
nand U47824 (N_47824,N_45918,N_45965);
nand U47825 (N_47825,N_44355,N_45702);
nor U47826 (N_47826,N_44560,N_44906);
and U47827 (N_47827,N_44549,N_44852);
or U47828 (N_47828,N_45069,N_44971);
and U47829 (N_47829,N_44176,N_45616);
xnor U47830 (N_47830,N_44454,N_45135);
and U47831 (N_47831,N_44343,N_44526);
nand U47832 (N_47832,N_44672,N_45750);
or U47833 (N_47833,N_44872,N_44321);
or U47834 (N_47834,N_44343,N_44815);
nor U47835 (N_47835,N_45601,N_45583);
nand U47836 (N_47836,N_44078,N_45807);
nand U47837 (N_47837,N_45121,N_45623);
xnor U47838 (N_47838,N_45088,N_45187);
nand U47839 (N_47839,N_44543,N_45109);
nand U47840 (N_47840,N_44140,N_44616);
or U47841 (N_47841,N_45851,N_45374);
nor U47842 (N_47842,N_44764,N_45182);
nand U47843 (N_47843,N_45095,N_45166);
xnor U47844 (N_47844,N_44414,N_44614);
and U47845 (N_47845,N_45799,N_45560);
nor U47846 (N_47846,N_44781,N_45747);
and U47847 (N_47847,N_44478,N_45458);
and U47848 (N_47848,N_45836,N_45314);
nor U47849 (N_47849,N_44288,N_45605);
or U47850 (N_47850,N_45169,N_44915);
nand U47851 (N_47851,N_44857,N_45090);
nor U47852 (N_47852,N_45300,N_45480);
nor U47853 (N_47853,N_45039,N_45573);
nand U47854 (N_47854,N_45125,N_45756);
xnor U47855 (N_47855,N_44539,N_45331);
and U47856 (N_47856,N_45247,N_45590);
or U47857 (N_47857,N_45457,N_45971);
or U47858 (N_47858,N_44100,N_45338);
nand U47859 (N_47859,N_45321,N_45860);
and U47860 (N_47860,N_45691,N_44881);
and U47861 (N_47861,N_45187,N_44493);
nand U47862 (N_47862,N_45173,N_45353);
nor U47863 (N_47863,N_44433,N_44341);
xnor U47864 (N_47864,N_45444,N_44663);
nor U47865 (N_47865,N_45387,N_44976);
nor U47866 (N_47866,N_45211,N_45606);
or U47867 (N_47867,N_44175,N_44729);
or U47868 (N_47868,N_45105,N_44553);
or U47869 (N_47869,N_44520,N_44919);
nand U47870 (N_47870,N_45232,N_44095);
nor U47871 (N_47871,N_45143,N_45661);
xnor U47872 (N_47872,N_45688,N_45884);
and U47873 (N_47873,N_45394,N_45513);
or U47874 (N_47874,N_44365,N_45253);
xnor U47875 (N_47875,N_45342,N_45749);
nand U47876 (N_47876,N_44698,N_44245);
and U47877 (N_47877,N_44019,N_44093);
or U47878 (N_47878,N_44703,N_45559);
and U47879 (N_47879,N_45341,N_44567);
nor U47880 (N_47880,N_45696,N_45050);
nor U47881 (N_47881,N_45230,N_44817);
nor U47882 (N_47882,N_44435,N_44228);
and U47883 (N_47883,N_45232,N_44972);
or U47884 (N_47884,N_45847,N_44389);
or U47885 (N_47885,N_45374,N_44494);
or U47886 (N_47886,N_44025,N_45980);
or U47887 (N_47887,N_44506,N_44760);
and U47888 (N_47888,N_44169,N_45970);
nor U47889 (N_47889,N_44877,N_44954);
or U47890 (N_47890,N_45013,N_45288);
nor U47891 (N_47891,N_45212,N_45004);
nand U47892 (N_47892,N_45362,N_44584);
nand U47893 (N_47893,N_45321,N_44941);
nand U47894 (N_47894,N_45031,N_45388);
nand U47895 (N_47895,N_45549,N_44563);
xor U47896 (N_47896,N_45264,N_44805);
nor U47897 (N_47897,N_45390,N_45259);
nor U47898 (N_47898,N_44816,N_44316);
nand U47899 (N_47899,N_45646,N_45386);
or U47900 (N_47900,N_44784,N_45060);
xnor U47901 (N_47901,N_45591,N_45095);
xor U47902 (N_47902,N_44809,N_44397);
nand U47903 (N_47903,N_44504,N_45235);
or U47904 (N_47904,N_45590,N_44803);
nand U47905 (N_47905,N_45430,N_45807);
or U47906 (N_47906,N_45297,N_45776);
nor U47907 (N_47907,N_45516,N_44201);
nor U47908 (N_47908,N_44298,N_44328);
or U47909 (N_47909,N_44787,N_44083);
nor U47910 (N_47910,N_44992,N_45348);
nor U47911 (N_47911,N_45933,N_44837);
nand U47912 (N_47912,N_44068,N_44004);
or U47913 (N_47913,N_44319,N_45486);
xnor U47914 (N_47914,N_44787,N_45237);
nor U47915 (N_47915,N_44047,N_44235);
nand U47916 (N_47916,N_45608,N_45900);
or U47917 (N_47917,N_44297,N_45904);
nand U47918 (N_47918,N_45231,N_45486);
or U47919 (N_47919,N_45747,N_44914);
or U47920 (N_47920,N_45023,N_44105);
or U47921 (N_47921,N_45277,N_45508);
or U47922 (N_47922,N_45572,N_45995);
and U47923 (N_47923,N_45998,N_45010);
or U47924 (N_47924,N_45176,N_45595);
and U47925 (N_47925,N_45261,N_45798);
xnor U47926 (N_47926,N_44169,N_44120);
nor U47927 (N_47927,N_44333,N_45554);
nand U47928 (N_47928,N_44846,N_45548);
nor U47929 (N_47929,N_44241,N_44805);
nor U47930 (N_47930,N_45361,N_44305);
or U47931 (N_47931,N_44581,N_45468);
and U47932 (N_47932,N_45973,N_45234);
nor U47933 (N_47933,N_44928,N_44238);
xor U47934 (N_47934,N_44465,N_44552);
or U47935 (N_47935,N_45993,N_44836);
xor U47936 (N_47936,N_44886,N_45119);
nor U47937 (N_47937,N_44135,N_44532);
xnor U47938 (N_47938,N_45345,N_44763);
nor U47939 (N_47939,N_44456,N_45770);
nand U47940 (N_47940,N_45417,N_44785);
and U47941 (N_47941,N_45815,N_44632);
xor U47942 (N_47942,N_44721,N_45224);
and U47943 (N_47943,N_44750,N_45219);
and U47944 (N_47944,N_45876,N_45946);
xor U47945 (N_47945,N_44782,N_45005);
and U47946 (N_47946,N_45397,N_45079);
or U47947 (N_47947,N_44260,N_45832);
or U47948 (N_47948,N_45561,N_44555);
or U47949 (N_47949,N_44655,N_44498);
xor U47950 (N_47950,N_44700,N_45336);
nor U47951 (N_47951,N_45249,N_44075);
or U47952 (N_47952,N_45261,N_44547);
or U47953 (N_47953,N_44081,N_44870);
nor U47954 (N_47954,N_44132,N_44514);
or U47955 (N_47955,N_44650,N_44868);
nand U47956 (N_47956,N_44041,N_44465);
nor U47957 (N_47957,N_45142,N_45140);
and U47958 (N_47958,N_44389,N_45866);
and U47959 (N_47959,N_44861,N_45663);
nor U47960 (N_47960,N_44958,N_45493);
and U47961 (N_47961,N_45623,N_45238);
nor U47962 (N_47962,N_45290,N_44887);
nand U47963 (N_47963,N_44300,N_45582);
xnor U47964 (N_47964,N_44311,N_45713);
nand U47965 (N_47965,N_45476,N_45065);
and U47966 (N_47966,N_45764,N_45727);
nor U47967 (N_47967,N_44945,N_45067);
nor U47968 (N_47968,N_44030,N_44191);
and U47969 (N_47969,N_45712,N_44148);
nor U47970 (N_47970,N_44375,N_45881);
nand U47971 (N_47971,N_44234,N_44675);
or U47972 (N_47972,N_44956,N_45047);
and U47973 (N_47973,N_44916,N_45613);
and U47974 (N_47974,N_45182,N_45362);
xnor U47975 (N_47975,N_44394,N_44861);
or U47976 (N_47976,N_45098,N_44069);
nand U47977 (N_47977,N_44788,N_45569);
nor U47978 (N_47978,N_45457,N_44550);
or U47979 (N_47979,N_45905,N_45950);
nor U47980 (N_47980,N_45934,N_44134);
or U47981 (N_47981,N_44594,N_44831);
nand U47982 (N_47982,N_44017,N_45662);
or U47983 (N_47983,N_44821,N_45039);
nand U47984 (N_47984,N_45759,N_45608);
nand U47985 (N_47985,N_45919,N_44069);
nor U47986 (N_47986,N_45814,N_44803);
nand U47987 (N_47987,N_45795,N_44580);
or U47988 (N_47988,N_45678,N_44770);
nand U47989 (N_47989,N_45628,N_44140);
and U47990 (N_47990,N_44441,N_45630);
xnor U47991 (N_47991,N_44458,N_45180);
or U47992 (N_47992,N_44050,N_45857);
nor U47993 (N_47993,N_44589,N_45863);
nor U47994 (N_47994,N_45205,N_45076);
nor U47995 (N_47995,N_45579,N_44278);
xor U47996 (N_47996,N_45379,N_45179);
nor U47997 (N_47997,N_44333,N_44159);
or U47998 (N_47998,N_44308,N_44375);
xor U47999 (N_47999,N_44220,N_45317);
and U48000 (N_48000,N_47421,N_47030);
and U48001 (N_48001,N_46031,N_47326);
or U48002 (N_48002,N_47060,N_47607);
nand U48003 (N_48003,N_46892,N_46678);
or U48004 (N_48004,N_46394,N_47138);
and U48005 (N_48005,N_47951,N_46554);
and U48006 (N_48006,N_47630,N_47396);
nand U48007 (N_48007,N_46188,N_46160);
and U48008 (N_48008,N_46714,N_46341);
and U48009 (N_48009,N_46896,N_47589);
and U48010 (N_48010,N_46638,N_47472);
and U48011 (N_48011,N_47841,N_47389);
or U48012 (N_48012,N_47545,N_46481);
xor U48013 (N_48013,N_46475,N_46017);
nor U48014 (N_48014,N_46075,N_47122);
nor U48015 (N_48015,N_46456,N_47853);
and U48016 (N_48016,N_46817,N_46921);
nor U48017 (N_48017,N_46329,N_47787);
nor U48018 (N_48018,N_46052,N_46322);
xnor U48019 (N_48019,N_46957,N_46081);
or U48020 (N_48020,N_46589,N_46376);
or U48021 (N_48021,N_46254,N_46506);
and U48022 (N_48022,N_46266,N_47916);
nand U48023 (N_48023,N_47790,N_47897);
or U48024 (N_48024,N_47331,N_46455);
and U48025 (N_48025,N_47145,N_47211);
or U48026 (N_48026,N_47987,N_46545);
xnor U48027 (N_48027,N_47686,N_47656);
nand U48028 (N_48028,N_47792,N_47891);
xnor U48029 (N_48029,N_46599,N_46229);
and U48030 (N_48030,N_46020,N_46588);
nand U48031 (N_48031,N_47579,N_46163);
nor U48032 (N_48032,N_47536,N_46606);
and U48033 (N_48033,N_47104,N_46038);
and U48034 (N_48034,N_47873,N_46916);
and U48035 (N_48035,N_47480,N_47203);
and U48036 (N_48036,N_46507,N_47007);
nor U48037 (N_48037,N_47142,N_46856);
nand U48038 (N_48038,N_47912,N_47105);
or U48039 (N_48039,N_46985,N_47143);
xnor U48040 (N_48040,N_46468,N_46291);
xnor U48041 (N_48041,N_47188,N_46926);
nor U48042 (N_48042,N_47923,N_46209);
or U48043 (N_48043,N_47931,N_47309);
and U48044 (N_48044,N_47922,N_46919);
nor U48045 (N_48045,N_47412,N_47023);
xor U48046 (N_48046,N_47198,N_46812);
or U48047 (N_48047,N_46251,N_46739);
nand U48048 (N_48048,N_47055,N_46256);
xnor U48049 (N_48049,N_46460,N_47748);
nand U48050 (N_48050,N_47302,N_46126);
or U48051 (N_48051,N_46218,N_47471);
or U48052 (N_48052,N_47084,N_47561);
nand U48053 (N_48053,N_46575,N_47521);
or U48054 (N_48054,N_47982,N_46009);
or U48055 (N_48055,N_47557,N_46718);
xnor U48056 (N_48056,N_47720,N_46012);
and U48057 (N_48057,N_46186,N_46899);
nand U48058 (N_48058,N_46294,N_47868);
nand U48059 (N_48059,N_46267,N_46463);
and U48060 (N_48060,N_46814,N_46767);
nor U48061 (N_48061,N_47469,N_47348);
nand U48062 (N_48062,N_46122,N_47524);
and U48063 (N_48063,N_47542,N_47422);
nand U48064 (N_48064,N_47051,N_46312);
xnor U48065 (N_48065,N_46519,N_46295);
or U48066 (N_48066,N_46411,N_47864);
or U48067 (N_48067,N_46906,N_47675);
xnor U48068 (N_48068,N_47628,N_46712);
nand U48069 (N_48069,N_47018,N_46986);
nand U48070 (N_48070,N_46960,N_47929);
nor U48071 (N_48071,N_47565,N_47419);
nor U48072 (N_48072,N_46366,N_47266);
or U48073 (N_48073,N_47443,N_46726);
nor U48074 (N_48074,N_46103,N_46841);
xnor U48075 (N_48075,N_46947,N_46752);
and U48076 (N_48076,N_47091,N_46168);
or U48077 (N_48077,N_47103,N_46583);
and U48078 (N_48078,N_47593,N_46059);
or U48079 (N_48079,N_46477,N_46318);
or U48080 (N_48080,N_47505,N_47726);
nor U48081 (N_48081,N_46962,N_46269);
nor U48082 (N_48082,N_47235,N_46998);
nand U48083 (N_48083,N_47898,N_46166);
xor U48084 (N_48084,N_47242,N_46696);
or U48085 (N_48085,N_47282,N_46040);
and U48086 (N_48086,N_46508,N_47642);
and U48087 (N_48087,N_46895,N_46239);
xor U48088 (N_48088,N_47756,N_46848);
xnor U48089 (N_48089,N_46368,N_46334);
nor U48090 (N_48090,N_47059,N_47394);
nand U48091 (N_48091,N_46815,N_46014);
or U48092 (N_48092,N_46244,N_47612);
or U48093 (N_48093,N_47402,N_47121);
nor U48094 (N_48094,N_46340,N_47076);
nand U48095 (N_48095,N_47381,N_46721);
and U48096 (N_48096,N_46129,N_47681);
xor U48097 (N_48097,N_46442,N_47174);
and U48098 (N_48098,N_47273,N_47118);
nor U48099 (N_48099,N_46749,N_47786);
nand U48100 (N_48100,N_46236,N_47383);
nand U48101 (N_48101,N_46661,N_46203);
nor U48102 (N_48102,N_47872,N_47942);
nor U48103 (N_48103,N_47563,N_46610);
and U48104 (N_48104,N_47894,N_46622);
and U48105 (N_48105,N_46479,N_47695);
xor U48106 (N_48106,N_47090,N_47517);
nor U48107 (N_48107,N_46922,N_47011);
nor U48108 (N_48108,N_46478,N_46959);
xnor U48109 (N_48109,N_46805,N_47149);
and U48110 (N_48110,N_46383,N_46082);
and U48111 (N_48111,N_46655,N_46104);
or U48112 (N_48112,N_46711,N_47291);
or U48113 (N_48113,N_46046,N_47719);
nor U48114 (N_48114,N_47155,N_47353);
and U48115 (N_48115,N_46543,N_46220);
or U48116 (N_48116,N_46204,N_47346);
or U48117 (N_48117,N_46375,N_46769);
nor U48118 (N_48118,N_46894,N_47647);
nor U48119 (N_48119,N_47233,N_46728);
xnor U48120 (N_48120,N_46932,N_46015);
nand U48121 (N_48121,N_47807,N_46772);
and U48122 (N_48122,N_47026,N_46564);
nand U48123 (N_48123,N_46471,N_47403);
and U48124 (N_48124,N_47655,N_47514);
and U48125 (N_48125,N_47566,N_46145);
nand U48126 (N_48126,N_46307,N_46346);
xor U48127 (N_48127,N_47967,N_46142);
nand U48128 (N_48128,N_47540,N_47013);
and U48129 (N_48129,N_47312,N_46883);
or U48130 (N_48130,N_46620,N_47519);
xnor U48131 (N_48131,N_46450,N_47310);
nor U48132 (N_48132,N_47861,N_47602);
xor U48133 (N_48133,N_46045,N_46582);
and U48134 (N_48134,N_46779,N_46541);
or U48135 (N_48135,N_46434,N_47515);
or U48136 (N_48136,N_46466,N_47371);
xnor U48137 (N_48137,N_46022,N_47307);
xor U48138 (N_48138,N_46486,N_46314);
nand U48139 (N_48139,N_47523,N_46461);
nand U48140 (N_48140,N_46987,N_47496);
nor U48141 (N_48141,N_47042,N_46816);
nor U48142 (N_48142,N_46200,N_47718);
xor U48143 (N_48143,N_47328,N_46303);
nor U48144 (N_48144,N_46968,N_47771);
or U48145 (N_48145,N_47934,N_46953);
and U48146 (N_48146,N_47603,N_47061);
or U48147 (N_48147,N_47003,N_46654);
and U48148 (N_48148,N_46969,N_47140);
nor U48149 (N_48149,N_46219,N_46097);
nand U48150 (N_48150,N_47116,N_46156);
or U48151 (N_48151,N_47658,N_47054);
nand U48152 (N_48152,N_46139,N_47028);
and U48153 (N_48153,N_46289,N_47795);
and U48154 (N_48154,N_47859,N_46143);
and U48155 (N_48155,N_46195,N_47458);
and U48156 (N_48156,N_46401,N_46268);
nor U48157 (N_48157,N_46591,N_46021);
xnor U48158 (N_48158,N_47509,N_46994);
nand U48159 (N_48159,N_47993,N_46601);
nor U48160 (N_48160,N_47989,N_46860);
xnor U48161 (N_48161,N_47345,N_46474);
nand U48162 (N_48162,N_46647,N_47966);
xnor U48163 (N_48163,N_46652,N_46955);
nand U48164 (N_48164,N_46003,N_47087);
nand U48165 (N_48165,N_47665,N_47941);
or U48166 (N_48166,N_46345,N_46578);
xnor U48167 (N_48167,N_46516,N_46153);
or U48168 (N_48168,N_47313,N_46646);
xnor U48169 (N_48169,N_47288,N_47560);
nand U48170 (N_48170,N_47330,N_46886);
or U48171 (N_48171,N_47991,N_46207);
nor U48172 (N_48172,N_46349,N_46447);
and U48173 (N_48173,N_46996,N_46213);
nand U48174 (N_48174,N_47337,N_47914);
nand U48175 (N_48175,N_46874,N_47881);
and U48176 (N_48176,N_47144,N_47927);
xnor U48177 (N_48177,N_46786,N_47713);
or U48178 (N_48178,N_46644,N_47865);
or U48179 (N_48179,N_46290,N_47161);
and U48180 (N_48180,N_47193,N_47315);
nor U48181 (N_48181,N_46065,N_46077);
and U48182 (N_48182,N_47549,N_46808);
and U48183 (N_48183,N_46016,N_47744);
xor U48184 (N_48184,N_47796,N_47216);
or U48185 (N_48185,N_46183,N_47685);
and U48186 (N_48186,N_46927,N_47308);
and U48187 (N_48187,N_46458,N_47433);
or U48188 (N_48188,N_47928,N_47298);
or U48189 (N_48189,N_46199,N_46540);
xnor U48190 (N_48190,N_47449,N_47210);
xor U48191 (N_48191,N_46399,N_46073);
or U48192 (N_48192,N_47910,N_47268);
nand U48193 (N_48193,N_46497,N_46277);
and U48194 (N_48194,N_46148,N_47283);
or U48195 (N_48195,N_46058,N_46400);
nand U48196 (N_48196,N_46514,N_47390);
xnor U48197 (N_48197,N_46804,N_46370);
nand U48198 (N_48198,N_46760,N_46252);
or U48199 (N_48199,N_47279,N_47503);
xnor U48200 (N_48200,N_46175,N_46102);
xor U48201 (N_48201,N_47812,N_46595);
or U48202 (N_48202,N_46337,N_46305);
or U48203 (N_48203,N_46558,N_47624);
and U48204 (N_48204,N_47583,N_46748);
and U48205 (N_48205,N_46264,N_46547);
xnor U48206 (N_48206,N_47250,N_46690);
or U48207 (N_48207,N_47270,N_47772);
or U48208 (N_48208,N_46286,N_46941);
nor U48209 (N_48209,N_47866,N_46071);
xor U48210 (N_48210,N_46823,N_47730);
xor U48211 (N_48211,N_47318,N_46887);
and U48212 (N_48212,N_46884,N_47276);
or U48213 (N_48213,N_47271,N_47305);
and U48214 (N_48214,N_46768,N_46745);
nor U48215 (N_48215,N_47552,N_47543);
nand U48216 (N_48216,N_46181,N_46951);
xnor U48217 (N_48217,N_46611,N_46320);
and U48218 (N_48218,N_47435,N_46417);
or U48219 (N_48219,N_47473,N_46873);
and U48220 (N_48220,N_47454,N_47842);
nand U48221 (N_48221,N_47654,N_46544);
or U48222 (N_48222,N_47219,N_46348);
nor U48223 (N_48223,N_47366,N_46490);
or U48224 (N_48224,N_47754,N_47578);
and U48225 (N_48225,N_47907,N_46722);
nand U48226 (N_48226,N_47431,N_46327);
nor U48227 (N_48227,N_46352,N_47662);
and U48228 (N_48228,N_46720,N_46433);
and U48229 (N_48229,N_47277,N_46551);
nand U48230 (N_48230,N_46628,N_47014);
nor U48231 (N_48231,N_47025,N_46282);
or U48232 (N_48232,N_47339,N_47320);
and U48233 (N_48233,N_47901,N_46250);
nand U48234 (N_48234,N_46005,N_47836);
nand U48235 (N_48235,N_46579,N_46988);
nor U48236 (N_48236,N_47078,N_46942);
xor U48237 (N_48237,N_47159,N_47732);
xor U48238 (N_48238,N_46862,N_47797);
nand U48239 (N_48239,N_47102,N_47869);
nand U48240 (N_48240,N_46078,N_46571);
and U48241 (N_48241,N_46882,N_47939);
nor U48242 (N_48242,N_47213,N_46840);
xnor U48243 (N_48243,N_46574,N_46495);
nor U48244 (N_48244,N_46758,N_46441);
and U48245 (N_48245,N_47166,N_47997);
nor U48246 (N_48246,N_46997,N_47132);
nand U48247 (N_48247,N_47971,N_47676);
nor U48248 (N_48248,N_47251,N_46934);
or U48249 (N_48249,N_47915,N_47131);
or U48250 (N_48250,N_46662,N_47349);
xor U48251 (N_48251,N_46083,N_46432);
or U48252 (N_48252,N_47197,N_47892);
and U48253 (N_48253,N_46018,N_47538);
and U48254 (N_48254,N_47553,N_46824);
xnor U48255 (N_48255,N_46271,N_47810);
and U48256 (N_48256,N_46134,N_46469);
or U48257 (N_48257,N_47697,N_46794);
and U48258 (N_48258,N_47176,N_46624);
and U48259 (N_48259,N_47906,N_47506);
nand U48260 (N_48260,N_46671,N_47809);
nand U48261 (N_48261,N_47491,N_47024);
nand U48262 (N_48262,N_47937,N_47784);
xnor U48263 (N_48263,N_46037,N_46948);
or U48264 (N_48264,N_46563,N_47187);
nor U48265 (N_48265,N_47010,N_47860);
nor U48266 (N_48266,N_46636,N_47564);
and U48267 (N_48267,N_47246,N_46167);
nand U48268 (N_48268,N_46498,N_46585);
xor U48269 (N_48269,N_46053,N_47293);
nand U48270 (N_48270,N_46502,N_46092);
and U48271 (N_48271,N_47021,N_46773);
xor U48272 (N_48272,N_47640,N_46827);
nand U48273 (N_48273,N_47970,N_47779);
or U48274 (N_48274,N_46245,N_47284);
nor U48275 (N_48275,N_47992,N_47370);
xor U48276 (N_48276,N_47481,N_47386);
nand U48277 (N_48277,N_47848,N_47043);
or U48278 (N_48278,N_47633,N_46424);
nand U48279 (N_48279,N_47526,N_47067);
nand U48280 (N_48280,N_47262,N_47113);
xnor U48281 (N_48281,N_47759,N_47767);
and U48282 (N_48282,N_47816,N_46706);
and U48283 (N_48283,N_47033,N_46384);
xor U48284 (N_48284,N_47889,N_46499);
and U48285 (N_48285,N_46914,N_47582);
or U48286 (N_48286,N_47500,N_47813);
or U48287 (N_48287,N_46913,N_47005);
nor U48288 (N_48288,N_47199,N_47379);
and U48289 (N_48289,N_46136,N_47782);
nor U48290 (N_48290,N_47334,N_47414);
or U48291 (N_48291,N_47350,N_46697);
and U48292 (N_48292,N_47008,N_46623);
xor U48293 (N_48293,N_47287,N_46033);
and U48294 (N_48294,N_47064,N_47747);
or U48295 (N_48295,N_47996,N_46422);
nor U48296 (N_48296,N_46556,N_46284);
and U48297 (N_48297,N_46496,N_46235);
nor U48298 (N_48298,N_47446,N_47548);
nor U48299 (N_48299,N_46803,N_47027);
or U48300 (N_48300,N_46945,N_47998);
nand U48301 (N_48301,N_47380,N_46179);
xor U48302 (N_48302,N_46665,N_46965);
nand U48303 (N_48303,N_46673,N_46421);
nor U48304 (N_48304,N_46858,N_47688);
nand U48305 (N_48305,N_47776,N_47858);
nand U48306 (N_48306,N_46263,N_46023);
xnor U48307 (N_48307,N_46609,N_47344);
and U48308 (N_48308,N_46656,N_47252);
or U48309 (N_48309,N_46682,N_47728);
xor U48310 (N_48310,N_47227,N_46797);
and U48311 (N_48311,N_47306,N_46691);
nand U48312 (N_48312,N_47743,N_47236);
nand U48313 (N_48313,N_46783,N_47206);
and U48314 (N_48314,N_47527,N_46249);
nor U48315 (N_48315,N_47530,N_47200);
and U48316 (N_48316,N_47333,N_47314);
nor U48317 (N_48317,N_47365,N_46465);
and U48318 (N_48318,N_46643,N_46403);
nor U48319 (N_48319,N_46389,N_47913);
and U48320 (N_48320,N_47444,N_47887);
nor U48321 (N_48321,N_47494,N_46522);
xor U48322 (N_48322,N_47762,N_47099);
and U48323 (N_48323,N_46231,N_47399);
nor U48324 (N_48324,N_47677,N_46576);
or U48325 (N_48325,N_47512,N_46889);
xnor U48326 (N_48326,N_46626,N_46049);
or U48327 (N_48327,N_47826,N_47832);
nand U48328 (N_48328,N_47173,N_47324);
and U48329 (N_48329,N_46190,N_46449);
nand U48330 (N_48330,N_47755,N_46790);
or U48331 (N_48331,N_47715,N_47946);
nand U48332 (N_48332,N_46736,N_46750);
nor U48333 (N_48333,N_47031,N_47294);
nand U48334 (N_48334,N_47709,N_47725);
xnor U48335 (N_48335,N_47332,N_46822);
or U48336 (N_48336,N_47053,N_47664);
nor U48337 (N_48337,N_47046,N_46171);
and U48338 (N_48338,N_46146,N_47855);
xnor U48339 (N_48339,N_46358,N_46215);
or U48340 (N_48340,N_46866,N_47554);
or U48341 (N_48341,N_46339,N_46119);
xnor U48342 (N_48342,N_47511,N_46299);
and U48343 (N_48343,N_47650,N_46637);
nor U48344 (N_48344,N_46388,N_47740);
xor U48345 (N_48345,N_46517,N_46331);
and U48346 (N_48346,N_46351,N_46128);
xnor U48347 (N_48347,N_47479,N_47232);
or U48348 (N_48348,N_47184,N_46310);
or U48349 (N_48349,N_47663,N_47299);
nor U48350 (N_48350,N_47995,N_46741);
and U48351 (N_48351,N_47608,N_47735);
nor U48352 (N_48352,N_46679,N_46048);
and U48353 (N_48353,N_46801,N_46127);
or U48354 (N_48354,N_46344,N_46831);
nand U48355 (N_48355,N_46857,N_47958);
or U48356 (N_48356,N_47595,N_46683);
and U48357 (N_48357,N_47351,N_46616);
nand U48358 (N_48358,N_47979,N_47115);
xnor U48359 (N_48359,N_47611,N_47933);
xor U48360 (N_48360,N_46864,N_47625);
and U48361 (N_48361,N_46629,N_47632);
xnor U48362 (N_48362,N_46854,N_46660);
nor U48363 (N_48363,N_47034,N_47867);
or U48364 (N_48364,N_47671,N_46381);
or U48365 (N_48365,N_46954,N_47101);
nor U48366 (N_48366,N_47151,N_47097);
xnor U48367 (N_48367,N_47134,N_46505);
nor U48368 (N_48368,N_46253,N_47824);
or U48369 (N_48369,N_47154,N_46030);
nand U48370 (N_48370,N_46285,N_46118);
nor U48371 (N_48371,N_47167,N_46323);
and U48372 (N_48372,N_47172,N_46642);
or U48373 (N_48373,N_46255,N_46710);
xnor U48374 (N_48374,N_46648,N_46905);
xor U48375 (N_48375,N_47082,N_46311);
nor U48376 (N_48376,N_47004,N_46765);
xnor U48377 (N_48377,N_47965,N_46594);
xnor U48378 (N_48378,N_46419,N_47201);
or U48379 (N_48379,N_46100,N_47501);
nand U48380 (N_48380,N_47918,N_46759);
xor U48381 (N_48381,N_47150,N_47765);
nand U48382 (N_48382,N_47890,N_46977);
and U48383 (N_48383,N_47190,N_47609);
nand U48384 (N_48384,N_46843,N_46792);
nor U48385 (N_48385,N_47111,N_46566);
and U48386 (N_48386,N_46933,N_46708);
xor U48387 (N_48387,N_47799,N_46261);
and U48388 (N_48388,N_46799,N_47168);
and U48389 (N_48389,N_47645,N_46839);
nor U48390 (N_48390,N_46232,N_47228);
xor U48391 (N_48391,N_47217,N_47610);
nor U48392 (N_48392,N_46774,N_47094);
xnor U48393 (N_48393,N_46632,N_47035);
xnor U48394 (N_48394,N_47462,N_46230);
xor U48395 (N_48395,N_47420,N_46151);
nand U48396 (N_48396,N_47237,N_46451);
xnor U48397 (N_48397,N_47849,N_47146);
xor U48398 (N_48398,N_47050,N_46832);
or U48399 (N_48399,N_46004,N_46374);
nand U48400 (N_48400,N_46452,N_47470);
nand U48401 (N_48401,N_47475,N_47830);
or U48402 (N_48402,N_47802,N_47729);
and U48403 (N_48403,N_46859,N_47823);
xnor U48404 (N_48404,N_47773,N_47518);
xnor U48405 (N_48405,N_47428,N_46061);
or U48406 (N_48406,N_47065,N_46723);
and U48407 (N_48407,N_46732,N_46108);
or U48408 (N_48408,N_46523,N_47960);
or U48409 (N_48409,N_46740,N_47120);
or U48410 (N_48410,N_46670,N_46747);
nor U48411 (N_48411,N_46068,N_47940);
or U48412 (N_48412,N_47562,N_47874);
nand U48413 (N_48413,N_47834,N_47944);
nand U48414 (N_48414,N_46354,N_46343);
nand U48415 (N_48415,N_46630,N_46810);
and U48416 (N_48416,N_47281,N_46762);
or U48417 (N_48417,N_47418,N_46568);
nand U48418 (N_48418,N_46426,N_47264);
or U48419 (N_48419,N_47147,N_47999);
nand U48420 (N_48420,N_47751,N_47788);
nor U48421 (N_48421,N_46182,N_47077);
xor U48422 (N_48422,N_46373,N_46995);
nor U48423 (N_48423,N_46993,N_46006);
or U48424 (N_48424,N_46818,N_47988);
or U48425 (N_48425,N_46000,N_47136);
xnor U48426 (N_48426,N_46482,N_47429);
nand U48427 (N_48427,N_47207,N_47949);
and U48428 (N_48428,N_47800,N_47300);
nand U48429 (N_48429,N_47930,N_47905);
or U48430 (N_48430,N_47378,N_47592);
or U48431 (N_48431,N_47356,N_46570);
nand U48432 (N_48432,N_46243,N_46970);
or U48433 (N_48433,N_47617,N_47598);
xor U48434 (N_48434,N_47156,N_47653);
xnor U48435 (N_48435,N_46846,N_46332);
nand U48436 (N_48436,N_47742,N_47037);
or U48437 (N_48437,N_46042,N_46333);
or U48438 (N_48438,N_46435,N_47727);
xnor U48439 (N_48439,N_47362,N_47416);
and U48440 (N_48440,N_47845,N_46980);
nor U48441 (N_48441,N_47107,N_46789);
nand U48442 (N_48442,N_47620,N_47627);
nor U48443 (N_48443,N_46174,N_47485);
or U48444 (N_48444,N_46027,N_47857);
xor U48445 (N_48445,N_46111,N_47885);
or U48446 (N_48446,N_47466,N_46501);
nor U48447 (N_48447,N_47649,N_47581);
nand U48448 (N_48448,N_46743,N_46084);
and U48449 (N_48449,N_46001,N_47497);
and U48450 (N_48450,N_46444,N_47130);
and U48451 (N_48451,N_47089,N_47781);
nor U48452 (N_48452,N_47192,N_46353);
or U48453 (N_48453,N_47408,N_46380);
nand U48454 (N_48454,N_46565,N_47423);
nor U48455 (N_48455,N_47701,N_46173);
nand U48456 (N_48456,N_46855,N_47070);
nand U48457 (N_48457,N_46237,N_46276);
and U48458 (N_48458,N_47019,N_47002);
and U48459 (N_48459,N_46764,N_47483);
or U48460 (N_48460,N_46511,N_46695);
nand U48461 (N_48461,N_46110,N_46713);
or U48462 (N_48462,N_46437,N_47261);
nand U48463 (N_48463,N_47708,N_46292);
or U48464 (N_48464,N_47106,N_47793);
or U48465 (N_48465,N_47057,N_47241);
and U48466 (N_48466,N_47680,N_46079);
or U48467 (N_48467,N_47733,N_46106);
or U48468 (N_48468,N_46725,N_47798);
and U48469 (N_48469,N_46095,N_47202);
and U48470 (N_48470,N_47690,N_46260);
and U48471 (N_48471,N_46169,N_46135);
nand U48472 (N_48472,N_47917,N_47811);
xor U48473 (N_48473,N_46775,N_47432);
nand U48474 (N_48474,N_46597,N_46819);
nand U48475 (N_48475,N_47181,N_47691);
and U48476 (N_48476,N_46372,N_47818);
and U48477 (N_48477,N_47407,N_46029);
or U48478 (N_48478,N_47259,N_47777);
nor U48479 (N_48479,N_47182,N_47248);
xnor U48480 (N_48480,N_47577,N_46067);
or U48481 (N_48481,N_46144,N_46569);
nand U48482 (N_48482,N_46115,N_47978);
or U48483 (N_48483,N_46089,N_47001);
xnor U48484 (N_48484,N_46013,N_46216);
or U48485 (N_48485,N_47945,N_47133);
or U48486 (N_48486,N_47705,N_46653);
nand U48487 (N_48487,N_47038,N_46724);
xor U48488 (N_48488,N_46192,N_46367);
xnor U48489 (N_48489,N_46915,N_47597);
and U48490 (N_48490,N_46055,N_47731);
nand U48491 (N_48491,N_47975,N_46771);
nor U48492 (N_48492,N_46807,N_47706);
or U48493 (N_48493,N_47178,N_47616);
or U48494 (N_48494,N_46635,N_46602);
nand U48495 (N_48495,N_47170,N_47534);
or U48496 (N_48496,N_47072,N_46709);
nand U48497 (N_48497,N_46850,N_47096);
nor U48498 (N_48498,N_47763,N_47212);
nand U48499 (N_48499,N_46793,N_47343);
nand U48500 (N_48500,N_46315,N_46596);
nor U48501 (N_48501,N_46929,N_46931);
xor U48502 (N_48502,N_46705,N_46178);
xor U48503 (N_48503,N_46076,N_46909);
xor U48504 (N_48504,N_46761,N_47840);
and U48505 (N_48505,N_47081,N_47039);
nand U48506 (N_48506,N_46639,N_47977);
nor U48507 (N_48507,N_46211,N_46088);
and U48508 (N_48508,N_46800,N_47438);
nor U48509 (N_48509,N_46716,N_47126);
xnor U48510 (N_48510,N_46967,N_47477);
or U48511 (N_48511,N_47492,N_47532);
and U48512 (N_48512,N_47376,N_47738);
xor U48513 (N_48513,N_47162,N_47135);
or U48514 (N_48514,N_47764,N_46844);
and U48515 (N_48515,N_47714,N_47938);
and U48516 (N_48516,N_46227,N_47240);
nor U48517 (N_48517,N_46757,N_46246);
nand U48518 (N_48518,N_46008,N_47619);
xnor U48519 (N_48519,N_47392,N_46233);
nand U48520 (N_48520,N_46537,N_46476);
and U48521 (N_48521,N_46542,N_46520);
nand U48522 (N_48522,N_47425,N_46838);
nand U48523 (N_48523,N_47745,N_46270);
nor U48524 (N_48524,N_47643,N_47157);
or U48525 (N_48525,N_46885,N_47789);
xnor U48526 (N_48526,N_46123,N_46694);
or U48527 (N_48527,N_47639,N_47817);
nor U48528 (N_48528,N_47158,N_47434);
nand U48529 (N_48529,N_47879,N_47447);
and U48530 (N_48530,N_46409,N_47086);
or U48531 (N_48531,N_47336,N_46763);
nor U48532 (N_48532,N_46193,N_47635);
nor U48533 (N_48533,N_47179,N_47098);
or U48534 (N_48534,N_46335,N_47244);
xnor U48535 (N_48535,N_46689,N_46438);
or U48536 (N_48536,N_46615,N_46707);
nand U48537 (N_48537,N_47510,N_47606);
nor U48538 (N_48538,N_47904,N_46090);
nor U48539 (N_48539,N_46613,N_46238);
and U48540 (N_48540,N_46420,N_47405);
or U48541 (N_48541,N_47388,N_47631);
xor U48542 (N_48542,N_47785,N_46872);
nand U48543 (N_48543,N_46754,N_46319);
nand U48544 (N_48544,N_46901,N_47100);
or U48545 (N_48545,N_47095,N_47358);
xor U48546 (N_48546,N_46669,N_46666);
xor U48547 (N_48547,N_46064,N_47504);
and U48548 (N_48548,N_47794,N_47783);
nor U48549 (N_48549,N_46105,N_46494);
nor U48550 (N_48550,N_47588,N_47361);
nand U48551 (N_48551,N_47531,N_46676);
nand U48552 (N_48552,N_46198,N_47976);
xnor U48553 (N_48553,N_47292,N_47736);
nand U48554 (N_48554,N_47225,N_46555);
and U48555 (N_48555,N_47016,N_46984);
nor U48556 (N_48556,N_47660,N_47382);
nor U48557 (N_48557,N_47445,N_47301);
nor U48558 (N_48558,N_47075,N_47994);
nor U48559 (N_48559,N_46159,N_47460);
nor U48560 (N_48560,N_47068,N_46663);
or U48561 (N_48561,N_46778,N_46043);
or U48562 (N_48562,N_46503,N_46036);
and U48563 (N_48563,N_47029,N_47770);
or U48564 (N_48564,N_46539,N_46687);
xor U48565 (N_48565,N_47613,N_46313);
nor U48566 (N_48566,N_46412,N_47049);
nand U48567 (N_48567,N_46436,N_47417);
or U48568 (N_48568,N_46133,N_47123);
and U48569 (N_48569,N_46212,N_46521);
xnor U48570 (N_48570,N_46457,N_46274);
nor U48571 (N_48571,N_47226,N_47956);
and U48572 (N_48572,N_46698,N_47629);
and U48573 (N_48573,N_47924,N_46668);
and U48574 (N_48574,N_46464,N_46280);
and U48575 (N_48575,N_46950,N_47805);
nand U48576 (N_48576,N_47260,N_47963);
and U48577 (N_48577,N_46205,N_46904);
or U48578 (N_48578,N_46184,N_47766);
or U48579 (N_48579,N_47615,N_47015);
nand U48580 (N_48580,N_46631,N_47384);
or U48581 (N_48581,N_47195,N_46378);
xor U48582 (N_48582,N_46881,N_47846);
nor U48583 (N_48583,N_47490,N_46228);
xor U48584 (N_48584,N_46066,N_47591);
nor U48585 (N_48585,N_47265,N_47245);
nand U48586 (N_48586,N_47911,N_47700);
nand U48587 (N_48587,N_47400,N_47231);
nand U48588 (N_48588,N_47902,N_47644);
xor U48589 (N_48589,N_46869,N_47452);
nand U48590 (N_48590,N_47875,N_47363);
or U48591 (N_48591,N_46693,N_46137);
or U48592 (N_48592,N_46928,N_47541);
or U48593 (N_48593,N_46060,N_46492);
nor U48594 (N_48594,N_46484,N_47843);
xnor U48595 (N_48595,N_47856,N_47450);
or U48596 (N_48596,N_47218,N_46584);
xnor U48597 (N_48597,N_47451,N_46811);
or U48598 (N_48598,N_46019,N_47909);
and U48599 (N_48599,N_47208,N_46273);
nor U48600 (N_48600,N_46937,N_47364);
nor U48601 (N_48601,N_46991,N_47249);
nor U48602 (N_48602,N_46350,N_46524);
xnor U48603 (N_48603,N_47711,N_47621);
nand U48604 (N_48604,N_46470,N_46158);
xnor U48605 (N_48605,N_47837,N_46363);
nand U48606 (N_48606,N_46301,N_46480);
xor U48607 (N_48607,N_47636,N_47406);
and U48608 (N_48608,N_46491,N_46397);
and U48609 (N_48609,N_46870,N_47585);
and U48610 (N_48610,N_46776,N_47883);
nor U48611 (N_48611,N_46918,N_46217);
and U48612 (N_48612,N_47436,N_47893);
nor U48613 (N_48613,N_47397,N_47269);
and U48614 (N_48614,N_47669,N_47368);
xor U48615 (N_48615,N_47804,N_46891);
or U48616 (N_48616,N_46784,N_46080);
and U48617 (N_48617,N_47550,N_47441);
nor U48618 (N_48618,N_47572,N_46258);
nor U48619 (N_48619,N_46391,N_47476);
nand U48620 (N_48620,N_46956,N_47164);
nor U48621 (N_48621,N_47153,N_47646);
nand U48622 (N_48622,N_46828,N_47952);
and U48623 (N_48623,N_47508,N_47223);
nand U48624 (N_48624,N_47539,N_47255);
nand U48625 (N_48625,N_46347,N_46034);
nand U48626 (N_48626,N_46429,N_46510);
or U48627 (N_48627,N_47215,N_47373);
nand U48628 (N_48628,N_46974,N_46262);
or U48629 (N_48629,N_47876,N_46924);
or U48630 (N_48630,N_47465,N_47862);
nor U48631 (N_48631,N_46070,N_46658);
nand U48632 (N_48632,N_46113,N_46098);
or U48633 (N_48633,N_46672,N_47835);
or U48634 (N_48634,N_47574,N_47413);
nand U48635 (N_48635,N_47833,N_47605);
or U48636 (N_48636,N_47604,N_47984);
or U48637 (N_48637,N_46050,N_46590);
nor U48638 (N_48638,N_47575,N_46109);
and U48639 (N_48639,N_47185,N_47461);
nor U48640 (N_48640,N_46701,N_47129);
xor U48641 (N_48641,N_47768,N_46733);
or U48642 (N_48642,N_46051,N_47175);
xor U48643 (N_48643,N_47814,N_47297);
nand U48644 (N_48644,N_46172,N_47827);
xnor U48645 (N_48645,N_46608,N_46737);
nand U48646 (N_48646,N_46296,N_46911);
or U48647 (N_48647,N_46283,N_47243);
or U48648 (N_48648,N_46085,N_47753);
and U48649 (N_48649,N_47478,N_46527);
nor U48650 (N_48650,N_46826,N_47495);
nor U48651 (N_48651,N_47074,N_46925);
or U48652 (N_48652,N_47325,N_46485);
xnor U48653 (N_48653,N_47045,N_46324);
nand U48654 (N_48654,N_47186,N_47704);
nand U48655 (N_48655,N_46963,N_47110);
and U48656 (N_48656,N_46112,N_46785);
nor U48657 (N_48657,N_47032,N_47831);
nand U48658 (N_48658,N_46880,N_46493);
or U48659 (N_48659,N_46650,N_47224);
nor U48660 (N_48660,N_46851,N_47278);
or U48661 (N_48661,N_46852,N_47442);
nand U48662 (N_48662,N_47377,N_46336);
or U48663 (N_48663,N_46820,N_46154);
nor U48664 (N_48664,N_46699,N_46281);
or U48665 (N_48665,N_47626,N_46140);
or U48666 (N_48666,N_46356,N_47815);
xor U48667 (N_48667,N_47806,N_46062);
nor U48668 (N_48668,N_46096,N_46330);
nand U48669 (N_48669,N_46861,N_47555);
or U48670 (N_48670,N_47707,N_47600);
or U48671 (N_48671,N_47069,N_47637);
and U48672 (N_48672,N_47844,N_46257);
and U48673 (N_48673,N_46504,N_47296);
or U48674 (N_48674,N_46386,N_46187);
xnor U48675 (N_48675,N_46338,N_47171);
and U48676 (N_48676,N_46007,N_47694);
or U48677 (N_48677,N_47000,N_46413);
nor U48678 (N_48678,N_47903,N_47821);
nand U48679 (N_48679,N_46530,N_47319);
nor U48680 (N_48680,N_47659,N_47528);
nor U48681 (N_48681,N_47758,N_47239);
and U48682 (N_48682,N_47180,N_47870);
nand U48683 (N_48683,N_46893,N_46964);
nand U48684 (N_48684,N_46645,N_46813);
and U48685 (N_48685,N_46234,N_47369);
xnor U48686 (N_48686,N_47969,N_47899);
and U48687 (N_48687,N_46972,N_47056);
or U48688 (N_48688,N_46056,N_46536);
or U48689 (N_48689,N_47424,N_46526);
or U48690 (N_48690,N_46548,N_47258);
or U48691 (N_48691,N_47499,N_46845);
nor U48692 (N_48692,N_46259,N_47295);
xor U48693 (N_48693,N_46396,N_46297);
and U48694 (N_48694,N_46035,N_46221);
nand U48695 (N_48695,N_46912,N_46382);
and U48696 (N_48696,N_46715,N_47457);
and U48697 (N_48697,N_46462,N_46483);
and U48698 (N_48698,N_46835,N_47974);
nand U48699 (N_48699,N_46439,N_47229);
xnor U48700 (N_48700,N_46935,N_47954);
nor U48701 (N_48701,N_47367,N_46719);
nor U48702 (N_48702,N_46917,N_46971);
xnor U48703 (N_48703,N_46500,N_47290);
xnor U48704 (N_48704,N_46528,N_46605);
and U48705 (N_48705,N_46738,N_47327);
or U48706 (N_48706,N_46057,N_46120);
nor U48707 (N_48707,N_46703,N_46164);
or U48708 (N_48708,N_47822,N_47769);
xor U48709 (N_48709,N_46727,N_47040);
nand U48710 (N_48710,N_47017,N_47455);
xor U48711 (N_48711,N_46361,N_46300);
xor U48712 (N_48712,N_46240,N_47329);
nand U48713 (N_48713,N_46572,N_47657);
nand U48714 (N_48714,N_47234,N_46976);
and U48715 (N_48715,N_47682,N_46879);
nand U48716 (N_48716,N_47571,N_46560);
xnor U48717 (N_48717,N_46074,N_47749);
or U48718 (N_48718,N_47453,N_46063);
nor U48719 (N_48719,N_46125,N_47652);
nor U48720 (N_48720,N_46293,N_46952);
and U48721 (N_48721,N_46897,N_47972);
xnor U48722 (N_48722,N_46930,N_47558);
or U48723 (N_48723,N_47439,N_47689);
and U48724 (N_48724,N_46999,N_47482);
and U48725 (N_48725,N_46044,N_47009);
and U48726 (N_48726,N_46940,N_46407);
nor U48727 (N_48727,N_46979,N_47486);
and U48728 (N_48728,N_47119,N_47648);
nand U48729 (N_48729,N_46405,N_47774);
and U48730 (N_48730,N_46002,N_46821);
or U48731 (N_48731,N_47177,N_46448);
nand U48732 (N_48732,N_46362,N_47169);
and U48733 (N_48733,N_46751,N_47791);
or U48734 (N_48734,N_46410,N_47638);
nand U48735 (N_48735,N_46586,N_47474);
xnor U48736 (N_48736,N_46011,N_47983);
nand U48737 (N_48737,N_47529,N_46659);
and U48738 (N_48738,N_46241,N_47340);
or U48739 (N_48739,N_46834,N_46598);
xnor U48740 (N_48740,N_47570,N_47973);
and U48741 (N_48741,N_46753,N_46944);
nand U48742 (N_48742,N_47522,N_47839);
nand U48743 (N_48743,N_47253,N_46387);
or U48744 (N_48744,N_46453,N_46700);
and U48745 (N_48745,N_47886,N_47036);
xnor U48746 (N_48746,N_47775,N_46177);
or U48747 (N_48747,N_47702,N_47684);
nor U48748 (N_48748,N_47267,N_47062);
and U48749 (N_48749,N_47847,N_47851);
xor U48750 (N_48750,N_46430,N_47880);
nor U48751 (N_48751,N_47568,N_47047);
nand U48752 (N_48752,N_47569,N_46321);
nand U48753 (N_48753,N_46640,N_47196);
nand U48754 (N_48754,N_46958,N_46214);
xor U48755 (N_48755,N_47670,N_47257);
nand U48756 (N_48756,N_47341,N_47012);
nor U48757 (N_48757,N_47354,N_47651);
and U48758 (N_48758,N_46981,N_47066);
nand U48759 (N_48759,N_47547,N_46559);
or U48760 (N_48760,N_46357,N_46875);
nor U48761 (N_48761,N_46157,N_46603);
and U48762 (N_48762,N_46392,N_46202);
or U48763 (N_48763,N_47112,N_47335);
nand U48764 (N_48764,N_46416,N_47194);
nand U48765 (N_48765,N_46116,N_46535);
or U48766 (N_48766,N_47238,N_47535);
and U48767 (N_48767,N_47165,N_47667);
and U48768 (N_48768,N_47962,N_46842);
nand U48769 (N_48769,N_47721,N_46047);
and U48770 (N_48770,N_46900,N_46890);
nand U48771 (N_48771,N_47668,N_46729);
nand U48772 (N_48772,N_46593,N_47189);
and U48773 (N_48773,N_47311,N_46978);
or U48774 (N_48774,N_47778,N_46117);
xnor U48775 (N_48775,N_46194,N_46876);
or U48776 (N_48776,N_47634,N_47430);
and U48777 (N_48777,N_46121,N_46101);
xor U48778 (N_48778,N_47863,N_46306);
or U48779 (N_48779,N_46625,N_47693);
or U48780 (N_48780,N_47520,N_47489);
and U48781 (N_48781,N_46371,N_47968);
xnor U48782 (N_48782,N_46686,N_46853);
or U48783 (N_48783,N_46210,N_46731);
nor U48784 (N_48784,N_46675,N_47352);
xnor U48785 (N_48785,N_47085,N_46730);
nor U48786 (N_48786,N_46684,N_46406);
and U48787 (N_48787,N_47580,N_46788);
nand U48788 (N_48788,N_46489,N_47359);
and U48789 (N_48789,N_47020,N_46222);
and U48790 (N_48790,N_46360,N_46717);
and U48791 (N_48791,N_47355,N_46734);
or U48792 (N_48792,N_46054,N_46830);
nand U48793 (N_48793,N_46275,N_47947);
or U48794 (N_48794,N_47594,N_46201);
xor U48795 (N_48795,N_46445,N_46533);
nand U48796 (N_48796,N_47537,N_47985);
nand U48797 (N_48797,N_46242,N_46086);
and U48798 (N_48798,N_47819,N_46278);
nand U48799 (N_48799,N_46390,N_47507);
or U48800 (N_48800,N_46617,N_47401);
or U48801 (N_48801,N_46580,N_47404);
nor U48802 (N_48802,N_46248,N_47936);
and U48803 (N_48803,N_46744,N_47828);
and U48804 (N_48804,N_46777,N_47109);
and U48805 (N_48805,N_46170,N_47209);
or U48806 (N_48806,N_47525,N_46992);
nor U48807 (N_48807,N_46402,N_46518);
xnor U48808 (N_48808,N_46039,N_46032);
and U48809 (N_48809,N_47920,N_47838);
or U48810 (N_48810,N_47556,N_46132);
and U48811 (N_48811,N_47493,N_47551);
xor U48812 (N_48812,N_47780,N_47926);
xnor U48813 (N_48813,N_47052,N_46226);
nand U48814 (N_48814,N_47925,N_47596);
nor U48815 (N_48815,N_46910,N_47573);
nor U48816 (N_48816,N_47125,N_46865);
xor U48817 (N_48817,N_47878,N_47426);
or U48818 (N_48818,N_46619,N_47761);
or U48819 (N_48819,N_46155,N_46641);
and U48820 (N_48820,N_46627,N_47280);
xor U48821 (N_48821,N_47342,N_46847);
or U48822 (N_48822,N_47374,N_47908);
and U48823 (N_48823,N_46836,N_46304);
nor U48824 (N_48824,N_46966,N_47882);
nand U48825 (N_48825,N_46868,N_46780);
and U48826 (N_48826,N_46791,N_46604);
nor U48827 (N_48827,N_47641,N_47221);
nand U48828 (N_48828,N_47205,N_47895);
nand U48829 (N_48829,N_47114,N_47080);
xor U48830 (N_48830,N_47440,N_46990);
or U48831 (N_48831,N_46983,N_46531);
or U48832 (N_48832,N_46552,N_46902);
xor U48833 (N_48833,N_46829,N_47666);
nor U48834 (N_48834,N_46467,N_47437);
nand U48835 (N_48835,N_46557,N_47073);
xor U48836 (N_48836,N_47124,N_47459);
nand U48837 (N_48837,N_47163,N_47673);
and U48838 (N_48838,N_47955,N_46787);
nand U48839 (N_48839,N_47272,N_46208);
xor U48840 (N_48840,N_46587,N_47502);
xor U48841 (N_48841,N_47141,N_46428);
or U48842 (N_48842,N_47559,N_46224);
and U48843 (N_48843,N_46425,N_47183);
nand U48844 (N_48844,N_47398,N_47567);
or U48845 (N_48845,N_46196,N_47623);
nor U48846 (N_48846,N_46664,N_46141);
and U48847 (N_48847,N_46946,N_47411);
nor U48848 (N_48848,N_47943,N_46355);
or U48849 (N_48849,N_47716,N_46364);
or U48850 (N_48850,N_46600,N_46379);
xnor U48851 (N_48851,N_46685,N_47393);
and U48852 (N_48852,N_47387,N_46404);
nand U48853 (N_48853,N_46796,N_47092);
and U48854 (N_48854,N_46287,N_47980);
nand U48855 (N_48855,N_47304,N_46026);
and U48856 (N_48856,N_47587,N_46509);
xor U48857 (N_48857,N_46472,N_46692);
nor U48858 (N_48858,N_46573,N_47322);
xnor U48859 (N_48859,N_46581,N_46431);
or U48860 (N_48860,N_46091,N_47919);
and U48861 (N_48861,N_46621,N_46782);
nand U48862 (N_48862,N_46878,N_46180);
nand U48863 (N_48863,N_47063,N_46592);
and U48864 (N_48864,N_47083,N_46440);
nor U48865 (N_48865,N_47750,N_46825);
nand U48866 (N_48866,N_46443,N_47222);
xor U48867 (N_48867,N_46550,N_46325);
and U48868 (N_48868,N_47964,N_47884);
nand U48869 (N_48869,N_47739,N_46704);
and U48870 (N_48870,N_47484,N_47986);
nand U48871 (N_48871,N_46920,N_47959);
and U48872 (N_48872,N_46446,N_47896);
and U48873 (N_48873,N_46735,N_47071);
nor U48874 (N_48874,N_47679,N_47357);
or U48875 (N_48875,N_47214,N_46415);
xor U48876 (N_48876,N_46114,N_47760);
nor U48877 (N_48877,N_46365,N_47139);
nand U48878 (N_48878,N_47850,N_47712);
nand U48879 (N_48879,N_47692,N_46418);
and U48880 (N_48880,N_47710,N_46408);
nor U48881 (N_48881,N_46898,N_47256);
xor U48882 (N_48882,N_46328,N_46657);
and U48883 (N_48883,N_46010,N_47093);
nor U48884 (N_48884,N_47950,N_47323);
nor U48885 (N_48885,N_47360,N_47801);
xor U48886 (N_48886,N_47752,N_47317);
and U48887 (N_48887,N_47128,N_47614);
and U48888 (N_48888,N_46532,N_46185);
or U48889 (N_48889,N_47516,N_47696);
and U48890 (N_48890,N_46534,N_46206);
nand U48891 (N_48891,N_47338,N_46342);
nor U48892 (N_48892,N_47672,N_46131);
and U48893 (N_48893,N_47274,N_47079);
xnor U48894 (N_48894,N_46833,N_46124);
nor U48895 (N_48895,N_47852,N_46265);
xnor U48896 (N_48896,N_46863,N_46756);
or U48897 (N_48897,N_46567,N_46150);
nand U48898 (N_48898,N_47703,N_47990);
or U48899 (N_48899,N_46680,N_47191);
and U48900 (N_48900,N_46546,N_47599);
or U48901 (N_48901,N_46223,N_46798);
or U48902 (N_48902,N_46427,N_46538);
nand U48903 (N_48903,N_46908,N_46487);
or U48904 (N_48904,N_46024,N_47044);
nand U48905 (N_48905,N_46982,N_47395);
or U48906 (N_48906,N_47464,N_46755);
nor U48907 (N_48907,N_46316,N_47127);
and U48908 (N_48908,N_47372,N_47160);
or U48909 (N_48909,N_46488,N_47415);
and U48910 (N_48910,N_47618,N_47498);
and U48911 (N_48911,N_47467,N_46975);
and U48912 (N_48912,N_47347,N_47058);
nor U48913 (N_48913,N_46176,N_47820);
and U48914 (N_48914,N_46562,N_46302);
xor U48915 (N_48915,N_47088,N_47391);
nor U48916 (N_48916,N_46152,N_46888);
nor U48917 (N_48917,N_47678,N_47275);
nor U48918 (N_48918,N_47900,N_46867);
or U48919 (N_48919,N_46308,N_47385);
nand U48920 (N_48920,N_47204,N_46189);
nand U48921 (N_48921,N_46087,N_46877);
xnor U48922 (N_48922,N_46423,N_46191);
and U48923 (N_48923,N_46949,N_46529);
and U48924 (N_48924,N_47448,N_46612);
nand U48925 (N_48925,N_46688,N_46414);
or U48926 (N_48926,N_47285,N_46025);
or U48927 (N_48927,N_46459,N_47463);
nor U48928 (N_48928,N_46041,N_46938);
xor U48929 (N_48929,N_46513,N_47871);
nand U48930 (N_48930,N_47041,N_47601);
xor U48931 (N_48931,N_47757,N_47022);
nand U48932 (N_48932,N_46770,N_46681);
xor U48933 (N_48933,N_46359,N_47661);
xor U48934 (N_48934,N_46961,N_46871);
xor U48935 (N_48935,N_46225,N_47152);
and U48936 (N_48936,N_46781,N_47006);
xor U48937 (N_48937,N_46943,N_46165);
or U48938 (N_48938,N_46288,N_46395);
nor U48939 (N_48939,N_47932,N_47584);
nor U48940 (N_48940,N_46607,N_46667);
nand U48941 (N_48941,N_46674,N_47953);
or U48942 (N_48942,N_46147,N_46279);
nor U48943 (N_48943,N_46746,N_46149);
and U48944 (N_48944,N_47263,N_46107);
nand U48945 (N_48945,N_46028,N_47303);
and U48946 (N_48946,N_47957,N_47289);
xnor U48947 (N_48947,N_46162,N_47734);
xnor U48948 (N_48948,N_47888,N_46099);
xnor U48949 (N_48949,N_46553,N_47487);
and U48950 (N_48950,N_47829,N_46298);
xor U48951 (N_48951,N_47456,N_47687);
nand U48952 (N_48952,N_47513,N_46634);
xnor U48953 (N_48953,N_46614,N_46369);
and U48954 (N_48954,N_46272,N_46795);
and U48955 (N_48955,N_47247,N_47948);
and U48956 (N_48956,N_46802,N_47674);
nand U48957 (N_48957,N_47546,N_46973);
or U48958 (N_48958,N_46473,N_46525);
and U48959 (N_48959,N_46385,N_46069);
xor U48960 (N_48960,N_47590,N_46515);
nor U48961 (N_48961,N_46677,N_47488);
xnor U48962 (N_48962,N_46454,N_47137);
nand U48963 (N_48963,N_47544,N_46072);
or U48964 (N_48964,N_46197,N_47803);
or U48965 (N_48965,N_47316,N_47723);
and U48966 (N_48966,N_47746,N_46939);
xor U48967 (N_48967,N_47724,N_47108);
and U48968 (N_48968,N_46649,N_46809);
nor U48969 (N_48969,N_47698,N_46130);
nand U48970 (N_48970,N_46989,N_46393);
xor U48971 (N_48971,N_46309,N_46633);
xor U48972 (N_48972,N_46247,N_46094);
and U48973 (N_48973,N_47622,N_47220);
or U48974 (N_48974,N_46577,N_47683);
and U48975 (N_48975,N_47737,N_46561);
xor U48976 (N_48976,N_46326,N_46398);
xor U48977 (N_48977,N_47117,N_47808);
or U48978 (N_48978,N_47148,N_46837);
xor U48979 (N_48979,N_47375,N_47409);
xor U48980 (N_48980,N_47877,N_47286);
and U48981 (N_48981,N_47854,N_47935);
nand U48982 (N_48982,N_46317,N_46923);
nand U48983 (N_48983,N_46512,N_46093);
nor U48984 (N_48984,N_47717,N_47321);
nor U48985 (N_48985,N_47427,N_46849);
nor U48986 (N_48986,N_47699,N_47741);
and U48987 (N_48987,N_47981,N_47533);
or U48988 (N_48988,N_47586,N_46618);
and U48989 (N_48989,N_46806,N_47921);
and U48990 (N_48990,N_47254,N_47722);
or U48991 (N_48991,N_46651,N_46702);
or U48992 (N_48992,N_47230,N_46138);
or U48993 (N_48993,N_47825,N_47468);
nor U48994 (N_48994,N_47961,N_47576);
nand U48995 (N_48995,N_46377,N_47048);
and U48996 (N_48996,N_46766,N_46907);
nand U48997 (N_48997,N_47410,N_46161);
nand U48998 (N_48998,N_46549,N_46903);
or U48999 (N_48999,N_46936,N_46742);
or U49000 (N_49000,N_46962,N_47886);
nand U49001 (N_49001,N_47613,N_47207);
xor U49002 (N_49002,N_47147,N_47434);
and U49003 (N_49003,N_46901,N_47390);
nand U49004 (N_49004,N_47246,N_47277);
or U49005 (N_49005,N_47444,N_46956);
nand U49006 (N_49006,N_46637,N_47224);
and U49007 (N_49007,N_47039,N_46571);
or U49008 (N_49008,N_47557,N_47865);
and U49009 (N_49009,N_46883,N_47475);
nand U49010 (N_49010,N_47545,N_47115);
xnor U49011 (N_49011,N_46055,N_47003);
nand U49012 (N_49012,N_47511,N_46917);
nand U49013 (N_49013,N_47025,N_47393);
and U49014 (N_49014,N_47589,N_47044);
nor U49015 (N_49015,N_47954,N_46281);
nand U49016 (N_49016,N_46386,N_47176);
or U49017 (N_49017,N_47660,N_46959);
nor U49018 (N_49018,N_47956,N_46754);
nand U49019 (N_49019,N_46919,N_47810);
or U49020 (N_49020,N_46967,N_46137);
and U49021 (N_49021,N_46859,N_46515);
nor U49022 (N_49022,N_46356,N_46652);
and U49023 (N_49023,N_46287,N_47782);
or U49024 (N_49024,N_47074,N_46492);
nor U49025 (N_49025,N_47151,N_47848);
nor U49026 (N_49026,N_46003,N_46024);
nand U49027 (N_49027,N_46293,N_47017);
or U49028 (N_49028,N_47433,N_47929);
nand U49029 (N_49029,N_47721,N_46377);
nor U49030 (N_49030,N_47543,N_46761);
nor U49031 (N_49031,N_47497,N_47771);
or U49032 (N_49032,N_46149,N_47499);
and U49033 (N_49033,N_46824,N_46863);
nor U49034 (N_49034,N_47544,N_47750);
and U49035 (N_49035,N_46260,N_46920);
or U49036 (N_49036,N_47197,N_46678);
nor U49037 (N_49037,N_47928,N_46152);
nor U49038 (N_49038,N_46188,N_47821);
xnor U49039 (N_49039,N_46859,N_47015);
or U49040 (N_49040,N_47881,N_47542);
or U49041 (N_49041,N_47827,N_46974);
nor U49042 (N_49042,N_46188,N_47720);
or U49043 (N_49043,N_47437,N_46192);
and U49044 (N_49044,N_47917,N_46422);
nor U49045 (N_49045,N_47868,N_46620);
or U49046 (N_49046,N_46162,N_46572);
nand U49047 (N_49047,N_46765,N_47453);
or U49048 (N_49048,N_47587,N_46434);
nand U49049 (N_49049,N_46130,N_47796);
xnor U49050 (N_49050,N_46599,N_46181);
and U49051 (N_49051,N_47363,N_47133);
and U49052 (N_49052,N_46947,N_47488);
nand U49053 (N_49053,N_46799,N_47889);
xor U49054 (N_49054,N_47678,N_47936);
or U49055 (N_49055,N_46049,N_47763);
and U49056 (N_49056,N_47600,N_46678);
xnor U49057 (N_49057,N_47058,N_47668);
nand U49058 (N_49058,N_47361,N_46686);
xnor U49059 (N_49059,N_47878,N_47356);
and U49060 (N_49060,N_47017,N_47168);
xnor U49061 (N_49061,N_46425,N_46272);
xor U49062 (N_49062,N_47936,N_47928);
and U49063 (N_49063,N_46194,N_46775);
nand U49064 (N_49064,N_47424,N_47849);
or U49065 (N_49065,N_47784,N_46229);
nand U49066 (N_49066,N_47099,N_46416);
xor U49067 (N_49067,N_46794,N_46552);
nand U49068 (N_49068,N_47120,N_46367);
xor U49069 (N_49069,N_47201,N_47041);
nand U49070 (N_49070,N_47924,N_46627);
nand U49071 (N_49071,N_47638,N_46723);
nor U49072 (N_49072,N_46332,N_47952);
or U49073 (N_49073,N_47162,N_46384);
or U49074 (N_49074,N_47182,N_47520);
nand U49075 (N_49075,N_46088,N_47891);
or U49076 (N_49076,N_46087,N_47705);
nand U49077 (N_49077,N_46766,N_46862);
nor U49078 (N_49078,N_47724,N_46330);
or U49079 (N_49079,N_47211,N_46989);
and U49080 (N_49080,N_47040,N_46573);
nor U49081 (N_49081,N_46353,N_46607);
nand U49082 (N_49082,N_47157,N_46371);
nand U49083 (N_49083,N_47816,N_46508);
nor U49084 (N_49084,N_47803,N_47398);
or U49085 (N_49085,N_47489,N_46804);
or U49086 (N_49086,N_47696,N_47164);
xnor U49087 (N_49087,N_47025,N_47488);
or U49088 (N_49088,N_46883,N_47064);
and U49089 (N_49089,N_47613,N_47208);
and U49090 (N_49090,N_46614,N_46526);
nor U49091 (N_49091,N_46600,N_47595);
nand U49092 (N_49092,N_47567,N_47992);
nor U49093 (N_49093,N_46389,N_47292);
xor U49094 (N_49094,N_46649,N_47287);
or U49095 (N_49095,N_47767,N_47351);
and U49096 (N_49096,N_47919,N_47226);
nand U49097 (N_49097,N_46324,N_46131);
and U49098 (N_49098,N_46718,N_47525);
and U49099 (N_49099,N_46626,N_47479);
xnor U49100 (N_49100,N_47948,N_47334);
nor U49101 (N_49101,N_46581,N_47739);
and U49102 (N_49102,N_46162,N_47131);
and U49103 (N_49103,N_47172,N_46664);
or U49104 (N_49104,N_47372,N_47846);
and U49105 (N_49105,N_46520,N_47290);
nor U49106 (N_49106,N_46630,N_47823);
xor U49107 (N_49107,N_46795,N_47917);
and U49108 (N_49108,N_46542,N_46458);
and U49109 (N_49109,N_46013,N_46391);
nor U49110 (N_49110,N_46337,N_46451);
and U49111 (N_49111,N_46843,N_47155);
nor U49112 (N_49112,N_46021,N_46274);
and U49113 (N_49113,N_47130,N_47052);
and U49114 (N_49114,N_46962,N_47732);
and U49115 (N_49115,N_46430,N_46750);
and U49116 (N_49116,N_47099,N_47899);
and U49117 (N_49117,N_47249,N_47977);
or U49118 (N_49118,N_46881,N_46109);
and U49119 (N_49119,N_46543,N_46345);
nor U49120 (N_49120,N_46969,N_47279);
nand U49121 (N_49121,N_47361,N_47821);
xnor U49122 (N_49122,N_46204,N_47265);
nor U49123 (N_49123,N_47042,N_46653);
nor U49124 (N_49124,N_47520,N_46560);
nor U49125 (N_49125,N_46405,N_46803);
and U49126 (N_49126,N_46932,N_46323);
xnor U49127 (N_49127,N_46369,N_47962);
nor U49128 (N_49128,N_47333,N_46032);
xnor U49129 (N_49129,N_47077,N_47655);
and U49130 (N_49130,N_47960,N_47645);
nor U49131 (N_49131,N_47875,N_46381);
xnor U49132 (N_49132,N_46954,N_46198);
xor U49133 (N_49133,N_46562,N_46703);
or U49134 (N_49134,N_46016,N_46780);
nor U49135 (N_49135,N_47402,N_46476);
or U49136 (N_49136,N_46366,N_46604);
nor U49137 (N_49137,N_46107,N_47049);
or U49138 (N_49138,N_47303,N_47783);
and U49139 (N_49139,N_46355,N_47508);
nor U49140 (N_49140,N_46090,N_47971);
and U49141 (N_49141,N_47734,N_46089);
xnor U49142 (N_49142,N_46541,N_46408);
xnor U49143 (N_49143,N_47625,N_46101);
nor U49144 (N_49144,N_47393,N_47274);
and U49145 (N_49145,N_46094,N_46187);
and U49146 (N_49146,N_47178,N_46000);
and U49147 (N_49147,N_46316,N_46286);
xor U49148 (N_49148,N_47213,N_46119);
nor U49149 (N_49149,N_47843,N_46698);
and U49150 (N_49150,N_46212,N_47074);
nand U49151 (N_49151,N_47378,N_46463);
and U49152 (N_49152,N_47552,N_47700);
and U49153 (N_49153,N_47550,N_46728);
and U49154 (N_49154,N_46576,N_46712);
and U49155 (N_49155,N_47386,N_47394);
nand U49156 (N_49156,N_46886,N_46824);
and U49157 (N_49157,N_46442,N_46659);
and U49158 (N_49158,N_46796,N_47553);
nand U49159 (N_49159,N_46461,N_47436);
xor U49160 (N_49160,N_47804,N_47801);
or U49161 (N_49161,N_47180,N_46812);
nor U49162 (N_49162,N_46513,N_46731);
xnor U49163 (N_49163,N_46347,N_47507);
nor U49164 (N_49164,N_46396,N_46399);
or U49165 (N_49165,N_46035,N_46282);
and U49166 (N_49166,N_47001,N_46641);
nand U49167 (N_49167,N_46314,N_47704);
nor U49168 (N_49168,N_47193,N_46282);
nor U49169 (N_49169,N_47313,N_47799);
or U49170 (N_49170,N_46749,N_47574);
nor U49171 (N_49171,N_46216,N_46916);
xnor U49172 (N_49172,N_46842,N_47584);
or U49173 (N_49173,N_47026,N_46340);
nand U49174 (N_49174,N_47481,N_46170);
or U49175 (N_49175,N_46916,N_47573);
xnor U49176 (N_49176,N_47721,N_47292);
nor U49177 (N_49177,N_46244,N_47709);
nor U49178 (N_49178,N_47165,N_47685);
xnor U49179 (N_49179,N_47558,N_46854);
xnor U49180 (N_49180,N_47961,N_47632);
nor U49181 (N_49181,N_46013,N_47623);
or U49182 (N_49182,N_46786,N_47190);
and U49183 (N_49183,N_47327,N_47348);
or U49184 (N_49184,N_46593,N_47067);
nand U49185 (N_49185,N_46640,N_46534);
xor U49186 (N_49186,N_46833,N_46435);
and U49187 (N_49187,N_46912,N_46735);
and U49188 (N_49188,N_47613,N_46572);
or U49189 (N_49189,N_46024,N_46826);
nor U49190 (N_49190,N_47553,N_46599);
or U49191 (N_49191,N_46566,N_47718);
xor U49192 (N_49192,N_46521,N_47036);
nand U49193 (N_49193,N_46150,N_47629);
xor U49194 (N_49194,N_47326,N_47101);
and U49195 (N_49195,N_46517,N_47687);
nand U49196 (N_49196,N_47584,N_47267);
xor U49197 (N_49197,N_47668,N_46062);
nand U49198 (N_49198,N_46420,N_47916);
xor U49199 (N_49199,N_46157,N_46801);
xnor U49200 (N_49200,N_47017,N_47712);
or U49201 (N_49201,N_46909,N_46136);
and U49202 (N_49202,N_46082,N_47345);
xnor U49203 (N_49203,N_46588,N_47534);
xor U49204 (N_49204,N_46848,N_47860);
nor U49205 (N_49205,N_46250,N_47377);
xor U49206 (N_49206,N_46366,N_47540);
xor U49207 (N_49207,N_47617,N_47160);
nand U49208 (N_49208,N_46658,N_47335);
xor U49209 (N_49209,N_47447,N_47243);
nor U49210 (N_49210,N_47100,N_46286);
xnor U49211 (N_49211,N_47776,N_46940);
nand U49212 (N_49212,N_47082,N_47495);
nor U49213 (N_49213,N_47199,N_46823);
or U49214 (N_49214,N_47473,N_46172);
nor U49215 (N_49215,N_47314,N_46041);
nor U49216 (N_49216,N_47162,N_47636);
nand U49217 (N_49217,N_46846,N_47507);
nand U49218 (N_49218,N_47042,N_46682);
nor U49219 (N_49219,N_46900,N_47968);
or U49220 (N_49220,N_47800,N_47175);
xor U49221 (N_49221,N_46108,N_47801);
nor U49222 (N_49222,N_46738,N_47925);
and U49223 (N_49223,N_46136,N_47212);
nor U49224 (N_49224,N_47426,N_46173);
and U49225 (N_49225,N_47206,N_47119);
nor U49226 (N_49226,N_47984,N_46567);
xor U49227 (N_49227,N_46798,N_47124);
xnor U49228 (N_49228,N_46137,N_46592);
nor U49229 (N_49229,N_47074,N_47614);
or U49230 (N_49230,N_47517,N_47217);
and U49231 (N_49231,N_46558,N_46086);
nand U49232 (N_49232,N_47602,N_46598);
and U49233 (N_49233,N_47797,N_47125);
nand U49234 (N_49234,N_47106,N_46421);
or U49235 (N_49235,N_47561,N_47466);
or U49236 (N_49236,N_47067,N_46244);
nor U49237 (N_49237,N_46385,N_47794);
nor U49238 (N_49238,N_46706,N_47712);
xnor U49239 (N_49239,N_47604,N_47614);
and U49240 (N_49240,N_47018,N_46636);
or U49241 (N_49241,N_47367,N_47793);
and U49242 (N_49242,N_46416,N_47464);
nand U49243 (N_49243,N_46853,N_47470);
nand U49244 (N_49244,N_47485,N_46069);
nand U49245 (N_49245,N_46423,N_46127);
nand U49246 (N_49246,N_47300,N_47411);
nor U49247 (N_49247,N_47479,N_47803);
nand U49248 (N_49248,N_46460,N_47432);
xor U49249 (N_49249,N_47145,N_46219);
nand U49250 (N_49250,N_46306,N_47060);
or U49251 (N_49251,N_47844,N_46381);
nor U49252 (N_49252,N_46669,N_47046);
xnor U49253 (N_49253,N_46766,N_46863);
and U49254 (N_49254,N_47711,N_46710);
and U49255 (N_49255,N_46531,N_46064);
or U49256 (N_49256,N_46066,N_47658);
or U49257 (N_49257,N_46605,N_46021);
or U49258 (N_49258,N_46942,N_47383);
nand U49259 (N_49259,N_46982,N_46127);
xnor U49260 (N_49260,N_46713,N_46006);
nand U49261 (N_49261,N_46570,N_46170);
nand U49262 (N_49262,N_46812,N_46040);
or U49263 (N_49263,N_47627,N_47763);
and U49264 (N_49264,N_46161,N_46289);
nor U49265 (N_49265,N_46286,N_46047);
and U49266 (N_49266,N_46524,N_47820);
xnor U49267 (N_49267,N_46191,N_47731);
or U49268 (N_49268,N_46399,N_47630);
or U49269 (N_49269,N_47487,N_47921);
and U49270 (N_49270,N_47355,N_46322);
nand U49271 (N_49271,N_47116,N_47224);
xor U49272 (N_49272,N_46929,N_46843);
or U49273 (N_49273,N_46530,N_47128);
and U49274 (N_49274,N_47302,N_47543);
and U49275 (N_49275,N_47291,N_47186);
nand U49276 (N_49276,N_46736,N_47534);
or U49277 (N_49277,N_46705,N_47588);
xor U49278 (N_49278,N_46156,N_46860);
and U49279 (N_49279,N_47840,N_46953);
or U49280 (N_49280,N_47751,N_47048);
xnor U49281 (N_49281,N_46452,N_46818);
or U49282 (N_49282,N_47426,N_47218);
xnor U49283 (N_49283,N_47683,N_47445);
nand U49284 (N_49284,N_47591,N_46753);
xor U49285 (N_49285,N_47085,N_47991);
and U49286 (N_49286,N_47511,N_47321);
or U49287 (N_49287,N_46779,N_46780);
or U49288 (N_49288,N_47753,N_47800);
xor U49289 (N_49289,N_46517,N_47958);
nor U49290 (N_49290,N_47034,N_47872);
and U49291 (N_49291,N_46105,N_47794);
xor U49292 (N_49292,N_47165,N_47130);
nor U49293 (N_49293,N_46553,N_46835);
and U49294 (N_49294,N_47699,N_47931);
nand U49295 (N_49295,N_47150,N_47252);
xnor U49296 (N_49296,N_46790,N_47554);
and U49297 (N_49297,N_46041,N_47982);
or U49298 (N_49298,N_47209,N_46729);
nand U49299 (N_49299,N_47849,N_47137);
or U49300 (N_49300,N_47330,N_47654);
xnor U49301 (N_49301,N_47273,N_47767);
or U49302 (N_49302,N_47296,N_47569);
or U49303 (N_49303,N_46407,N_47673);
nand U49304 (N_49304,N_47035,N_46309);
and U49305 (N_49305,N_47062,N_47526);
or U49306 (N_49306,N_46900,N_46579);
nor U49307 (N_49307,N_46293,N_46557);
xnor U49308 (N_49308,N_47033,N_46336);
and U49309 (N_49309,N_46558,N_47653);
nor U49310 (N_49310,N_47426,N_46120);
nor U49311 (N_49311,N_47209,N_46266);
and U49312 (N_49312,N_47137,N_46028);
nor U49313 (N_49313,N_47981,N_46513);
nor U49314 (N_49314,N_46713,N_47176);
xnor U49315 (N_49315,N_46108,N_46269);
nand U49316 (N_49316,N_46534,N_47378);
and U49317 (N_49317,N_46467,N_47061);
or U49318 (N_49318,N_46208,N_47003);
nor U49319 (N_49319,N_47272,N_47593);
xnor U49320 (N_49320,N_46123,N_46732);
nand U49321 (N_49321,N_46542,N_47652);
or U49322 (N_49322,N_47107,N_46632);
and U49323 (N_49323,N_47112,N_46337);
and U49324 (N_49324,N_46801,N_46767);
or U49325 (N_49325,N_47338,N_46018);
nor U49326 (N_49326,N_46283,N_47855);
or U49327 (N_49327,N_47415,N_47904);
xor U49328 (N_49328,N_46511,N_46144);
xor U49329 (N_49329,N_47611,N_47380);
nand U49330 (N_49330,N_47076,N_46179);
nor U49331 (N_49331,N_46390,N_47321);
or U49332 (N_49332,N_47483,N_46768);
nand U49333 (N_49333,N_47316,N_46034);
or U49334 (N_49334,N_46297,N_47183);
xnor U49335 (N_49335,N_46584,N_46370);
or U49336 (N_49336,N_46239,N_47596);
and U49337 (N_49337,N_47976,N_47923);
nor U49338 (N_49338,N_47255,N_47450);
nor U49339 (N_49339,N_46628,N_47925);
nand U49340 (N_49340,N_47892,N_46224);
xnor U49341 (N_49341,N_47981,N_47517);
or U49342 (N_49342,N_46715,N_46076);
or U49343 (N_49343,N_47362,N_46265);
and U49344 (N_49344,N_47763,N_47193);
and U49345 (N_49345,N_47043,N_46226);
xnor U49346 (N_49346,N_46638,N_47050);
xor U49347 (N_49347,N_47664,N_46780);
or U49348 (N_49348,N_46695,N_46576);
nor U49349 (N_49349,N_47548,N_46997);
or U49350 (N_49350,N_46578,N_47706);
and U49351 (N_49351,N_46504,N_47044);
and U49352 (N_49352,N_46043,N_46593);
nand U49353 (N_49353,N_47148,N_46037);
xor U49354 (N_49354,N_47658,N_46634);
xnor U49355 (N_49355,N_47757,N_46577);
nand U49356 (N_49356,N_47277,N_46688);
or U49357 (N_49357,N_46454,N_47301);
nand U49358 (N_49358,N_47083,N_46144);
nand U49359 (N_49359,N_46688,N_47398);
and U49360 (N_49360,N_46366,N_46174);
xor U49361 (N_49361,N_47183,N_46871);
nand U49362 (N_49362,N_47913,N_47382);
or U49363 (N_49363,N_47754,N_46843);
xor U49364 (N_49364,N_47114,N_46677);
and U49365 (N_49365,N_47063,N_47366);
nor U49366 (N_49366,N_47646,N_46635);
xnor U49367 (N_49367,N_47748,N_47148);
or U49368 (N_49368,N_46107,N_47811);
nand U49369 (N_49369,N_47102,N_47521);
or U49370 (N_49370,N_46406,N_47802);
nand U49371 (N_49371,N_47794,N_46427);
and U49372 (N_49372,N_47370,N_47260);
nand U49373 (N_49373,N_46998,N_47238);
xnor U49374 (N_49374,N_46860,N_46744);
nor U49375 (N_49375,N_47826,N_46500);
xnor U49376 (N_49376,N_46764,N_47449);
or U49377 (N_49377,N_47325,N_46462);
and U49378 (N_49378,N_47181,N_47730);
and U49379 (N_49379,N_47927,N_47638);
nor U49380 (N_49380,N_47024,N_46592);
nand U49381 (N_49381,N_47053,N_47143);
nor U49382 (N_49382,N_46008,N_47451);
nand U49383 (N_49383,N_46764,N_46047);
nand U49384 (N_49384,N_46024,N_47215);
xnor U49385 (N_49385,N_46067,N_46671);
nor U49386 (N_49386,N_46605,N_47497);
nand U49387 (N_49387,N_47783,N_46235);
or U49388 (N_49388,N_46553,N_46220);
nand U49389 (N_49389,N_46924,N_47984);
and U49390 (N_49390,N_46932,N_47373);
xor U49391 (N_49391,N_47387,N_46063);
nor U49392 (N_49392,N_46920,N_47672);
xnor U49393 (N_49393,N_46848,N_47128);
and U49394 (N_49394,N_46902,N_46428);
nand U49395 (N_49395,N_46574,N_47063);
nand U49396 (N_49396,N_47521,N_47418);
nor U49397 (N_49397,N_47329,N_46861);
or U49398 (N_49398,N_47819,N_47297);
nor U49399 (N_49399,N_46391,N_47821);
nor U49400 (N_49400,N_46480,N_47979);
or U49401 (N_49401,N_47041,N_46472);
nor U49402 (N_49402,N_47929,N_47581);
nand U49403 (N_49403,N_47375,N_46809);
xnor U49404 (N_49404,N_46835,N_47427);
nor U49405 (N_49405,N_46070,N_46993);
and U49406 (N_49406,N_46007,N_47769);
and U49407 (N_49407,N_46631,N_46414);
or U49408 (N_49408,N_47958,N_46262);
nand U49409 (N_49409,N_46072,N_47917);
or U49410 (N_49410,N_47324,N_46850);
xor U49411 (N_49411,N_46560,N_47044);
nand U49412 (N_49412,N_47602,N_46319);
nand U49413 (N_49413,N_47152,N_47381);
nand U49414 (N_49414,N_47960,N_47525);
nor U49415 (N_49415,N_47274,N_47940);
or U49416 (N_49416,N_46980,N_47596);
xor U49417 (N_49417,N_47809,N_47517);
xnor U49418 (N_49418,N_47259,N_47280);
xor U49419 (N_49419,N_46754,N_47199);
or U49420 (N_49420,N_47014,N_46976);
nor U49421 (N_49421,N_47269,N_47473);
nand U49422 (N_49422,N_46859,N_47196);
or U49423 (N_49423,N_47067,N_46050);
nand U49424 (N_49424,N_47112,N_47483);
and U49425 (N_49425,N_46704,N_47424);
nor U49426 (N_49426,N_46488,N_46373);
nor U49427 (N_49427,N_47047,N_46372);
xor U49428 (N_49428,N_47223,N_47581);
xnor U49429 (N_49429,N_46551,N_46345);
nor U49430 (N_49430,N_46986,N_46597);
and U49431 (N_49431,N_46340,N_46189);
nand U49432 (N_49432,N_47149,N_46285);
nor U49433 (N_49433,N_47454,N_46734);
xnor U49434 (N_49434,N_46745,N_46485);
nor U49435 (N_49435,N_46469,N_46132);
and U49436 (N_49436,N_46394,N_46112);
or U49437 (N_49437,N_46585,N_46704);
or U49438 (N_49438,N_47064,N_46533);
or U49439 (N_49439,N_47994,N_46957);
nand U49440 (N_49440,N_47455,N_46618);
nand U49441 (N_49441,N_46462,N_47210);
nor U49442 (N_49442,N_46623,N_47144);
and U49443 (N_49443,N_46889,N_47185);
xor U49444 (N_49444,N_46338,N_46194);
nor U49445 (N_49445,N_46931,N_46726);
nand U49446 (N_49446,N_47487,N_46282);
or U49447 (N_49447,N_47375,N_47643);
nor U49448 (N_49448,N_47920,N_47586);
nor U49449 (N_49449,N_46854,N_46847);
and U49450 (N_49450,N_46078,N_46382);
and U49451 (N_49451,N_47006,N_46714);
nand U49452 (N_49452,N_47862,N_47202);
nor U49453 (N_49453,N_47459,N_46875);
nand U49454 (N_49454,N_47918,N_47693);
nor U49455 (N_49455,N_46886,N_46412);
and U49456 (N_49456,N_47788,N_46832);
nor U49457 (N_49457,N_47967,N_46795);
nor U49458 (N_49458,N_47770,N_46613);
or U49459 (N_49459,N_47326,N_47759);
nand U49460 (N_49460,N_46527,N_46810);
xor U49461 (N_49461,N_47116,N_47579);
and U49462 (N_49462,N_46896,N_46525);
or U49463 (N_49463,N_47744,N_46932);
and U49464 (N_49464,N_46740,N_47065);
or U49465 (N_49465,N_47556,N_47528);
nor U49466 (N_49466,N_47077,N_47602);
nand U49467 (N_49467,N_46682,N_47717);
xnor U49468 (N_49468,N_47190,N_47422);
and U49469 (N_49469,N_46552,N_46089);
nand U49470 (N_49470,N_46527,N_47056);
and U49471 (N_49471,N_47711,N_47109);
xor U49472 (N_49472,N_47223,N_46325);
or U49473 (N_49473,N_46635,N_47449);
and U49474 (N_49474,N_47964,N_46700);
xnor U49475 (N_49475,N_46459,N_46232);
nor U49476 (N_49476,N_47307,N_47883);
nand U49477 (N_49477,N_47777,N_47537);
xnor U49478 (N_49478,N_46697,N_46588);
nor U49479 (N_49479,N_47102,N_47442);
nor U49480 (N_49480,N_46134,N_47256);
nor U49481 (N_49481,N_47086,N_47416);
xor U49482 (N_49482,N_47459,N_47354);
or U49483 (N_49483,N_46250,N_46468);
or U49484 (N_49484,N_46487,N_47749);
and U49485 (N_49485,N_46688,N_47065);
nor U49486 (N_49486,N_46469,N_47064);
or U49487 (N_49487,N_47117,N_46460);
xor U49488 (N_49488,N_46962,N_47312);
or U49489 (N_49489,N_47961,N_47406);
xor U49490 (N_49490,N_46033,N_46460);
or U49491 (N_49491,N_46960,N_47008);
nor U49492 (N_49492,N_46087,N_46377);
and U49493 (N_49493,N_47550,N_46467);
and U49494 (N_49494,N_47284,N_47762);
xor U49495 (N_49495,N_47671,N_47120);
or U49496 (N_49496,N_46859,N_46484);
and U49497 (N_49497,N_46894,N_47680);
xnor U49498 (N_49498,N_47159,N_46209);
xnor U49499 (N_49499,N_46002,N_47493);
nor U49500 (N_49500,N_46407,N_46916);
and U49501 (N_49501,N_46419,N_47972);
or U49502 (N_49502,N_46592,N_47124);
or U49503 (N_49503,N_47374,N_46872);
and U49504 (N_49504,N_46277,N_47428);
nand U49505 (N_49505,N_47512,N_47242);
xor U49506 (N_49506,N_47337,N_46052);
nor U49507 (N_49507,N_46386,N_46291);
or U49508 (N_49508,N_46285,N_46203);
nand U49509 (N_49509,N_47557,N_46432);
nand U49510 (N_49510,N_47043,N_46946);
or U49511 (N_49511,N_46943,N_47617);
and U49512 (N_49512,N_47149,N_46767);
and U49513 (N_49513,N_46132,N_46673);
xor U49514 (N_49514,N_46714,N_46711);
nor U49515 (N_49515,N_46294,N_46908);
or U49516 (N_49516,N_46002,N_46454);
nor U49517 (N_49517,N_47766,N_47777);
nor U49518 (N_49518,N_47626,N_47848);
and U49519 (N_49519,N_46202,N_46608);
nor U49520 (N_49520,N_47954,N_46023);
nor U49521 (N_49521,N_47825,N_46667);
and U49522 (N_49522,N_46446,N_46797);
and U49523 (N_49523,N_47258,N_46930);
or U49524 (N_49524,N_46648,N_46366);
or U49525 (N_49525,N_47616,N_47031);
and U49526 (N_49526,N_47933,N_47012);
nor U49527 (N_49527,N_47239,N_47146);
nor U49528 (N_49528,N_47121,N_47009);
nand U49529 (N_49529,N_46432,N_46869);
nand U49530 (N_49530,N_47536,N_47012);
nand U49531 (N_49531,N_46247,N_46142);
nand U49532 (N_49532,N_47970,N_47674);
xor U49533 (N_49533,N_47241,N_46278);
nor U49534 (N_49534,N_46041,N_47376);
or U49535 (N_49535,N_46030,N_46873);
or U49536 (N_49536,N_47658,N_47304);
or U49537 (N_49537,N_47598,N_47043);
and U49538 (N_49538,N_47944,N_47682);
nor U49539 (N_49539,N_47715,N_46921);
and U49540 (N_49540,N_47482,N_46373);
nand U49541 (N_49541,N_47974,N_46034);
or U49542 (N_49542,N_46718,N_46403);
xnor U49543 (N_49543,N_47046,N_47773);
xnor U49544 (N_49544,N_46106,N_47339);
nor U49545 (N_49545,N_46453,N_47437);
nor U49546 (N_49546,N_46639,N_47573);
nand U49547 (N_49547,N_46381,N_46727);
nand U49548 (N_49548,N_47226,N_46569);
nor U49549 (N_49549,N_47436,N_46768);
nand U49550 (N_49550,N_47719,N_47760);
and U49551 (N_49551,N_46943,N_47037);
nor U49552 (N_49552,N_47102,N_46717);
or U49553 (N_49553,N_46402,N_46317);
or U49554 (N_49554,N_47119,N_46362);
nand U49555 (N_49555,N_47398,N_47115);
and U49556 (N_49556,N_46568,N_47452);
or U49557 (N_49557,N_47882,N_46202);
nand U49558 (N_49558,N_46470,N_46397);
nand U49559 (N_49559,N_46842,N_47647);
or U49560 (N_49560,N_46489,N_47382);
nor U49561 (N_49561,N_47942,N_46121);
nand U49562 (N_49562,N_46705,N_46403);
nand U49563 (N_49563,N_46492,N_46444);
nand U49564 (N_49564,N_46126,N_46066);
nand U49565 (N_49565,N_47195,N_47905);
nor U49566 (N_49566,N_46034,N_46640);
nor U49567 (N_49567,N_46058,N_46380);
xor U49568 (N_49568,N_47773,N_47039);
xnor U49569 (N_49569,N_46264,N_46640);
or U49570 (N_49570,N_46672,N_47327);
nand U49571 (N_49571,N_47635,N_46602);
and U49572 (N_49572,N_46826,N_47344);
and U49573 (N_49573,N_46757,N_47795);
or U49574 (N_49574,N_46340,N_47665);
xor U49575 (N_49575,N_46839,N_46627);
or U49576 (N_49576,N_47981,N_47456);
nor U49577 (N_49577,N_46144,N_47859);
and U49578 (N_49578,N_46769,N_47387);
nand U49579 (N_49579,N_46960,N_46373);
or U49580 (N_49580,N_46719,N_46932);
and U49581 (N_49581,N_46215,N_46677);
nand U49582 (N_49582,N_46371,N_46857);
nand U49583 (N_49583,N_46625,N_46936);
and U49584 (N_49584,N_46712,N_47305);
nand U49585 (N_49585,N_47283,N_47638);
or U49586 (N_49586,N_47312,N_46998);
nand U49587 (N_49587,N_46510,N_46068);
nor U49588 (N_49588,N_47453,N_47592);
nor U49589 (N_49589,N_46301,N_46947);
or U49590 (N_49590,N_47634,N_47178);
and U49591 (N_49591,N_47659,N_47814);
xnor U49592 (N_49592,N_46348,N_47350);
and U49593 (N_49593,N_47435,N_47744);
and U49594 (N_49594,N_47428,N_46444);
or U49595 (N_49595,N_47605,N_47565);
nand U49596 (N_49596,N_47640,N_46771);
nand U49597 (N_49597,N_47931,N_47997);
nor U49598 (N_49598,N_46287,N_47864);
xnor U49599 (N_49599,N_46561,N_46589);
nand U49600 (N_49600,N_47236,N_46531);
nor U49601 (N_49601,N_46652,N_47491);
or U49602 (N_49602,N_47838,N_46212);
or U49603 (N_49603,N_47063,N_46933);
and U49604 (N_49604,N_47316,N_46989);
nor U49605 (N_49605,N_47129,N_46130);
nor U49606 (N_49606,N_46147,N_47975);
and U49607 (N_49607,N_46863,N_46552);
and U49608 (N_49608,N_47430,N_46413);
nand U49609 (N_49609,N_46629,N_46822);
or U49610 (N_49610,N_46693,N_46395);
nand U49611 (N_49611,N_47249,N_46480);
nand U49612 (N_49612,N_47023,N_47477);
xor U49613 (N_49613,N_47357,N_46682);
and U49614 (N_49614,N_47742,N_46561);
and U49615 (N_49615,N_46814,N_46610);
nor U49616 (N_49616,N_47999,N_46797);
or U49617 (N_49617,N_46231,N_46844);
or U49618 (N_49618,N_47862,N_46806);
xnor U49619 (N_49619,N_47258,N_46592);
and U49620 (N_49620,N_47047,N_47311);
nand U49621 (N_49621,N_47543,N_47181);
xnor U49622 (N_49622,N_47255,N_46955);
nor U49623 (N_49623,N_46097,N_46375);
nand U49624 (N_49624,N_46346,N_46721);
nor U49625 (N_49625,N_47880,N_47504);
xor U49626 (N_49626,N_47062,N_46304);
and U49627 (N_49627,N_46591,N_47576);
nor U49628 (N_49628,N_46832,N_46984);
nor U49629 (N_49629,N_46262,N_46191);
or U49630 (N_49630,N_46639,N_47931);
or U49631 (N_49631,N_46754,N_47103);
nor U49632 (N_49632,N_46041,N_46363);
xor U49633 (N_49633,N_46124,N_47912);
or U49634 (N_49634,N_47061,N_47422);
xor U49635 (N_49635,N_46466,N_47497);
nand U49636 (N_49636,N_46797,N_47996);
nor U49637 (N_49637,N_46515,N_46453);
nor U49638 (N_49638,N_47464,N_46829);
xor U49639 (N_49639,N_47494,N_46666);
nand U49640 (N_49640,N_47488,N_46406);
and U49641 (N_49641,N_46467,N_46310);
and U49642 (N_49642,N_47207,N_47948);
nand U49643 (N_49643,N_47723,N_46802);
nor U49644 (N_49644,N_46852,N_47079);
or U49645 (N_49645,N_46361,N_46054);
nor U49646 (N_49646,N_46042,N_46246);
and U49647 (N_49647,N_46073,N_46359);
xor U49648 (N_49648,N_46783,N_47971);
and U49649 (N_49649,N_47270,N_47217);
nand U49650 (N_49650,N_47642,N_46154);
or U49651 (N_49651,N_46675,N_46765);
xor U49652 (N_49652,N_46704,N_46334);
or U49653 (N_49653,N_47991,N_46206);
or U49654 (N_49654,N_46381,N_46914);
nand U49655 (N_49655,N_46270,N_47445);
nand U49656 (N_49656,N_46940,N_47537);
nor U49657 (N_49657,N_46685,N_47346);
nor U49658 (N_49658,N_46437,N_47600);
nor U49659 (N_49659,N_46644,N_47870);
nand U49660 (N_49660,N_47158,N_47124);
xnor U49661 (N_49661,N_47716,N_47615);
or U49662 (N_49662,N_46677,N_46611);
nor U49663 (N_49663,N_46296,N_47810);
nand U49664 (N_49664,N_46777,N_46993);
and U49665 (N_49665,N_47011,N_46985);
xnor U49666 (N_49666,N_46003,N_46121);
nand U49667 (N_49667,N_47400,N_47570);
nand U49668 (N_49668,N_47157,N_47158);
xnor U49669 (N_49669,N_46729,N_46548);
xnor U49670 (N_49670,N_46860,N_46592);
xnor U49671 (N_49671,N_46727,N_47945);
or U49672 (N_49672,N_46985,N_46048);
xnor U49673 (N_49673,N_47085,N_46735);
nand U49674 (N_49674,N_46138,N_47797);
nand U49675 (N_49675,N_46094,N_46836);
or U49676 (N_49676,N_46182,N_47558);
nor U49677 (N_49677,N_46425,N_47411);
nand U49678 (N_49678,N_46570,N_46119);
nor U49679 (N_49679,N_46099,N_47828);
and U49680 (N_49680,N_46488,N_46624);
nor U49681 (N_49681,N_46199,N_47911);
or U49682 (N_49682,N_46957,N_46282);
nand U49683 (N_49683,N_46872,N_47071);
and U49684 (N_49684,N_46259,N_46659);
xnor U49685 (N_49685,N_47535,N_46457);
or U49686 (N_49686,N_47309,N_46559);
nor U49687 (N_49687,N_46938,N_46392);
and U49688 (N_49688,N_46180,N_47563);
nand U49689 (N_49689,N_46557,N_47469);
xor U49690 (N_49690,N_46756,N_46800);
xnor U49691 (N_49691,N_46540,N_46453);
xnor U49692 (N_49692,N_46766,N_46925);
nand U49693 (N_49693,N_46905,N_47301);
nand U49694 (N_49694,N_46507,N_46563);
and U49695 (N_49695,N_46961,N_47500);
and U49696 (N_49696,N_46046,N_47281);
or U49697 (N_49697,N_46435,N_47281);
nor U49698 (N_49698,N_46267,N_46031);
xnor U49699 (N_49699,N_47334,N_47102);
xor U49700 (N_49700,N_46219,N_47272);
or U49701 (N_49701,N_46927,N_46358);
or U49702 (N_49702,N_46326,N_47079);
xor U49703 (N_49703,N_47716,N_46603);
xnor U49704 (N_49704,N_46392,N_46830);
xnor U49705 (N_49705,N_46337,N_47241);
and U49706 (N_49706,N_46307,N_46392);
xor U49707 (N_49707,N_47383,N_47709);
and U49708 (N_49708,N_47449,N_47294);
or U49709 (N_49709,N_47245,N_47689);
nor U49710 (N_49710,N_47739,N_47370);
nor U49711 (N_49711,N_46157,N_47238);
or U49712 (N_49712,N_47607,N_46802);
and U49713 (N_49713,N_46510,N_46255);
nand U49714 (N_49714,N_47927,N_46400);
and U49715 (N_49715,N_46640,N_46524);
and U49716 (N_49716,N_47633,N_46749);
nor U49717 (N_49717,N_46760,N_46587);
or U49718 (N_49718,N_46348,N_47328);
nand U49719 (N_49719,N_46151,N_46091);
nor U49720 (N_49720,N_47358,N_47112);
nand U49721 (N_49721,N_47823,N_47603);
nor U49722 (N_49722,N_46953,N_46150);
or U49723 (N_49723,N_47877,N_46354);
or U49724 (N_49724,N_47083,N_47289);
xnor U49725 (N_49725,N_47502,N_46996);
or U49726 (N_49726,N_47300,N_47900);
nand U49727 (N_49727,N_46960,N_47558);
and U49728 (N_49728,N_47130,N_46977);
nor U49729 (N_49729,N_47663,N_46903);
nor U49730 (N_49730,N_47920,N_46284);
and U49731 (N_49731,N_46393,N_46389);
and U49732 (N_49732,N_47796,N_47343);
xnor U49733 (N_49733,N_47478,N_46052);
or U49734 (N_49734,N_47517,N_47430);
nand U49735 (N_49735,N_47903,N_47438);
nor U49736 (N_49736,N_46569,N_46322);
nand U49737 (N_49737,N_47157,N_47075);
nand U49738 (N_49738,N_46248,N_46787);
nor U49739 (N_49739,N_47360,N_47967);
nor U49740 (N_49740,N_47454,N_47912);
nand U49741 (N_49741,N_47666,N_46953);
and U49742 (N_49742,N_46224,N_47619);
nor U49743 (N_49743,N_47463,N_47937);
xnor U49744 (N_49744,N_47671,N_46728);
or U49745 (N_49745,N_46200,N_47406);
or U49746 (N_49746,N_46900,N_46488);
or U49747 (N_49747,N_47387,N_46261);
nand U49748 (N_49748,N_47032,N_47463);
xnor U49749 (N_49749,N_47213,N_47569);
and U49750 (N_49750,N_47213,N_46533);
and U49751 (N_49751,N_46448,N_46587);
nor U49752 (N_49752,N_47000,N_47591);
xor U49753 (N_49753,N_47186,N_46274);
or U49754 (N_49754,N_47283,N_47866);
and U49755 (N_49755,N_47433,N_46570);
nor U49756 (N_49756,N_47016,N_46220);
or U49757 (N_49757,N_46116,N_47649);
and U49758 (N_49758,N_46220,N_47309);
xnor U49759 (N_49759,N_47101,N_47972);
nor U49760 (N_49760,N_47733,N_46930);
nor U49761 (N_49761,N_46757,N_46520);
nor U49762 (N_49762,N_46464,N_46977);
or U49763 (N_49763,N_46341,N_46640);
nor U49764 (N_49764,N_46684,N_46271);
nand U49765 (N_49765,N_46957,N_47526);
xor U49766 (N_49766,N_46706,N_47040);
or U49767 (N_49767,N_47005,N_46580);
nor U49768 (N_49768,N_47165,N_47220);
nand U49769 (N_49769,N_46449,N_47242);
nand U49770 (N_49770,N_46446,N_47592);
nand U49771 (N_49771,N_47170,N_47748);
nor U49772 (N_49772,N_46928,N_46567);
nand U49773 (N_49773,N_47345,N_47392);
xnor U49774 (N_49774,N_46809,N_46902);
or U49775 (N_49775,N_46299,N_46943);
and U49776 (N_49776,N_47574,N_47008);
or U49777 (N_49777,N_47005,N_47916);
nand U49778 (N_49778,N_46947,N_46080);
or U49779 (N_49779,N_47717,N_47470);
nor U49780 (N_49780,N_47130,N_46177);
nand U49781 (N_49781,N_47542,N_47135);
xnor U49782 (N_49782,N_47227,N_47272);
nand U49783 (N_49783,N_47020,N_47886);
nor U49784 (N_49784,N_47944,N_46409);
xor U49785 (N_49785,N_46645,N_47202);
or U49786 (N_49786,N_46597,N_47937);
xnor U49787 (N_49787,N_46717,N_47439);
or U49788 (N_49788,N_46402,N_46376);
and U49789 (N_49789,N_47515,N_47417);
nor U49790 (N_49790,N_46344,N_47165);
xor U49791 (N_49791,N_47042,N_46025);
and U49792 (N_49792,N_46342,N_47109);
nand U49793 (N_49793,N_46545,N_46042);
nand U49794 (N_49794,N_46351,N_46078);
xor U49795 (N_49795,N_47210,N_47820);
or U49796 (N_49796,N_47361,N_47294);
xor U49797 (N_49797,N_47336,N_47381);
or U49798 (N_49798,N_47186,N_47697);
and U49799 (N_49799,N_47739,N_47860);
or U49800 (N_49800,N_47720,N_46791);
or U49801 (N_49801,N_46394,N_47530);
or U49802 (N_49802,N_47589,N_46924);
or U49803 (N_49803,N_46877,N_47916);
nor U49804 (N_49804,N_46019,N_46816);
xnor U49805 (N_49805,N_46628,N_46537);
xnor U49806 (N_49806,N_47756,N_46295);
or U49807 (N_49807,N_46374,N_47647);
nor U49808 (N_49808,N_47916,N_47637);
nor U49809 (N_49809,N_47147,N_46926);
nor U49810 (N_49810,N_47351,N_46045);
nor U49811 (N_49811,N_47616,N_46241);
and U49812 (N_49812,N_46433,N_46790);
nor U49813 (N_49813,N_47220,N_46502);
or U49814 (N_49814,N_46781,N_47883);
or U49815 (N_49815,N_46451,N_47528);
xor U49816 (N_49816,N_46903,N_46634);
and U49817 (N_49817,N_46139,N_47065);
and U49818 (N_49818,N_46491,N_46712);
nor U49819 (N_49819,N_47545,N_47256);
xor U49820 (N_49820,N_46984,N_47895);
nand U49821 (N_49821,N_46820,N_46923);
xor U49822 (N_49822,N_46595,N_47646);
xor U49823 (N_49823,N_47584,N_46601);
xnor U49824 (N_49824,N_47356,N_46392);
xor U49825 (N_49825,N_46725,N_47499);
and U49826 (N_49826,N_47208,N_47395);
nand U49827 (N_49827,N_47061,N_46421);
and U49828 (N_49828,N_46180,N_46880);
nor U49829 (N_49829,N_47638,N_47695);
nor U49830 (N_49830,N_46933,N_46561);
or U49831 (N_49831,N_46373,N_47756);
nor U49832 (N_49832,N_46589,N_47838);
nand U49833 (N_49833,N_46688,N_46078);
nand U49834 (N_49834,N_46029,N_47979);
and U49835 (N_49835,N_47828,N_46956);
and U49836 (N_49836,N_47144,N_47663);
xnor U49837 (N_49837,N_47345,N_47998);
or U49838 (N_49838,N_46470,N_46239);
nand U49839 (N_49839,N_47713,N_46728);
xnor U49840 (N_49840,N_46344,N_47958);
or U49841 (N_49841,N_46544,N_46419);
or U49842 (N_49842,N_46056,N_47541);
nand U49843 (N_49843,N_46365,N_47206);
or U49844 (N_49844,N_47798,N_47220);
and U49845 (N_49845,N_46199,N_47452);
or U49846 (N_49846,N_46042,N_46178);
nor U49847 (N_49847,N_47473,N_46595);
and U49848 (N_49848,N_47072,N_47933);
or U49849 (N_49849,N_47074,N_47062);
xnor U49850 (N_49850,N_47278,N_47150);
and U49851 (N_49851,N_47457,N_47164);
or U49852 (N_49852,N_47636,N_46160);
or U49853 (N_49853,N_46353,N_46369);
or U49854 (N_49854,N_46398,N_46557);
nor U49855 (N_49855,N_46947,N_47405);
or U49856 (N_49856,N_46975,N_46757);
nand U49857 (N_49857,N_46027,N_47748);
xnor U49858 (N_49858,N_46611,N_47412);
xnor U49859 (N_49859,N_47730,N_47755);
nand U49860 (N_49860,N_47807,N_46036);
or U49861 (N_49861,N_47993,N_47725);
nor U49862 (N_49862,N_46261,N_46974);
nand U49863 (N_49863,N_47764,N_47375);
xnor U49864 (N_49864,N_46375,N_47511);
and U49865 (N_49865,N_46801,N_46320);
xnor U49866 (N_49866,N_47502,N_46264);
xor U49867 (N_49867,N_46750,N_46767);
nand U49868 (N_49868,N_46586,N_46969);
nand U49869 (N_49869,N_46939,N_47867);
or U49870 (N_49870,N_46560,N_47403);
or U49871 (N_49871,N_46092,N_46620);
nand U49872 (N_49872,N_46895,N_47796);
and U49873 (N_49873,N_47681,N_47781);
nor U49874 (N_49874,N_46475,N_47063);
nand U49875 (N_49875,N_46493,N_46847);
xor U49876 (N_49876,N_46483,N_47888);
and U49877 (N_49877,N_47324,N_47155);
and U49878 (N_49878,N_47425,N_47706);
xnor U49879 (N_49879,N_46755,N_46729);
and U49880 (N_49880,N_46966,N_46885);
or U49881 (N_49881,N_47636,N_46127);
and U49882 (N_49882,N_46195,N_47719);
or U49883 (N_49883,N_47847,N_46695);
and U49884 (N_49884,N_46736,N_47276);
and U49885 (N_49885,N_47917,N_47027);
nand U49886 (N_49886,N_46620,N_47532);
or U49887 (N_49887,N_46289,N_46891);
nand U49888 (N_49888,N_46939,N_46770);
and U49889 (N_49889,N_47183,N_47434);
and U49890 (N_49890,N_46174,N_47148);
nand U49891 (N_49891,N_47421,N_46490);
and U49892 (N_49892,N_47624,N_47842);
xor U49893 (N_49893,N_46322,N_47716);
nand U49894 (N_49894,N_47620,N_46016);
and U49895 (N_49895,N_46183,N_47614);
and U49896 (N_49896,N_46248,N_47272);
nand U49897 (N_49897,N_46689,N_47340);
or U49898 (N_49898,N_46458,N_46116);
xor U49899 (N_49899,N_46064,N_46902);
nor U49900 (N_49900,N_47312,N_46924);
xnor U49901 (N_49901,N_47433,N_46707);
nor U49902 (N_49902,N_47473,N_46043);
and U49903 (N_49903,N_46904,N_47075);
xnor U49904 (N_49904,N_47277,N_47191);
xnor U49905 (N_49905,N_47444,N_46486);
and U49906 (N_49906,N_46448,N_46865);
nand U49907 (N_49907,N_47721,N_46294);
nor U49908 (N_49908,N_46675,N_46170);
nand U49909 (N_49909,N_47191,N_47223);
and U49910 (N_49910,N_46482,N_47584);
nand U49911 (N_49911,N_47531,N_47302);
or U49912 (N_49912,N_46084,N_46646);
or U49913 (N_49913,N_46998,N_47914);
or U49914 (N_49914,N_47773,N_47622);
and U49915 (N_49915,N_47823,N_46254);
or U49916 (N_49916,N_47359,N_47551);
nor U49917 (N_49917,N_47119,N_46738);
nand U49918 (N_49918,N_47074,N_46062);
nor U49919 (N_49919,N_47330,N_46597);
xor U49920 (N_49920,N_46918,N_46314);
nand U49921 (N_49921,N_47807,N_46833);
or U49922 (N_49922,N_47433,N_46497);
or U49923 (N_49923,N_47101,N_46581);
nor U49924 (N_49924,N_46351,N_46364);
xor U49925 (N_49925,N_47259,N_46350);
or U49926 (N_49926,N_46318,N_46492);
xnor U49927 (N_49927,N_46048,N_47593);
nor U49928 (N_49928,N_46817,N_46541);
or U49929 (N_49929,N_47005,N_46050);
and U49930 (N_49930,N_46108,N_46624);
and U49931 (N_49931,N_47929,N_46504);
or U49932 (N_49932,N_46591,N_47255);
and U49933 (N_49933,N_46214,N_46879);
nand U49934 (N_49934,N_47693,N_46037);
nor U49935 (N_49935,N_47357,N_47900);
or U49936 (N_49936,N_46508,N_46486);
or U49937 (N_49937,N_47667,N_47003);
nor U49938 (N_49938,N_46020,N_47095);
or U49939 (N_49939,N_46434,N_47046);
nand U49940 (N_49940,N_46120,N_46848);
nand U49941 (N_49941,N_46182,N_47490);
or U49942 (N_49942,N_47506,N_46096);
nand U49943 (N_49943,N_47808,N_47501);
and U49944 (N_49944,N_46292,N_46634);
nand U49945 (N_49945,N_46578,N_46600);
nand U49946 (N_49946,N_47199,N_46191);
nand U49947 (N_49947,N_46749,N_47991);
nor U49948 (N_49948,N_46627,N_47212);
and U49949 (N_49949,N_47434,N_47966);
and U49950 (N_49950,N_46681,N_46745);
and U49951 (N_49951,N_46292,N_47144);
xor U49952 (N_49952,N_47514,N_46412);
and U49953 (N_49953,N_46579,N_47110);
or U49954 (N_49954,N_47951,N_47498);
nor U49955 (N_49955,N_47597,N_46760);
xor U49956 (N_49956,N_46051,N_47795);
or U49957 (N_49957,N_46372,N_46386);
and U49958 (N_49958,N_46615,N_47054);
and U49959 (N_49959,N_47812,N_46937);
xor U49960 (N_49960,N_47801,N_47735);
nor U49961 (N_49961,N_47343,N_47242);
or U49962 (N_49962,N_47675,N_47852);
and U49963 (N_49963,N_46048,N_46767);
nand U49964 (N_49964,N_46517,N_47465);
xnor U49965 (N_49965,N_47224,N_46305);
or U49966 (N_49966,N_46409,N_47750);
nand U49967 (N_49967,N_46943,N_46164);
xnor U49968 (N_49968,N_47670,N_46530);
and U49969 (N_49969,N_47296,N_46980);
xor U49970 (N_49970,N_47411,N_46169);
and U49971 (N_49971,N_47908,N_46231);
xnor U49972 (N_49972,N_46253,N_46371);
nand U49973 (N_49973,N_46726,N_46557);
and U49974 (N_49974,N_47059,N_46428);
xnor U49975 (N_49975,N_46368,N_47550);
xor U49976 (N_49976,N_47922,N_46454);
nor U49977 (N_49977,N_47647,N_47930);
xor U49978 (N_49978,N_47460,N_46191);
nand U49979 (N_49979,N_47315,N_47020);
nand U49980 (N_49980,N_47253,N_47071);
or U49981 (N_49981,N_46495,N_46851);
and U49982 (N_49982,N_46129,N_46872);
xnor U49983 (N_49983,N_46459,N_46005);
nor U49984 (N_49984,N_47084,N_47286);
xor U49985 (N_49985,N_47916,N_46529);
xor U49986 (N_49986,N_47153,N_46706);
nor U49987 (N_49987,N_47483,N_47714);
nand U49988 (N_49988,N_46343,N_47812);
nand U49989 (N_49989,N_46545,N_47778);
xnor U49990 (N_49990,N_47573,N_46874);
or U49991 (N_49991,N_47256,N_47571);
nor U49992 (N_49992,N_46004,N_47177);
and U49993 (N_49993,N_46753,N_46340);
and U49994 (N_49994,N_46072,N_46447);
and U49995 (N_49995,N_47287,N_47050);
and U49996 (N_49996,N_46392,N_47511);
nor U49997 (N_49997,N_46675,N_47047);
and U49998 (N_49998,N_46930,N_47764);
nor U49999 (N_49999,N_47900,N_46818);
nor UO_0 (O_0,N_48694,N_48072);
xor UO_1 (O_1,N_48675,N_48106);
and UO_2 (O_2,N_48282,N_49851);
nand UO_3 (O_3,N_48595,N_49198);
xnor UO_4 (O_4,N_48091,N_48894);
and UO_5 (O_5,N_48334,N_48364);
and UO_6 (O_6,N_48351,N_48197);
or UO_7 (O_7,N_49462,N_48882);
xnor UO_8 (O_8,N_49140,N_48909);
nor UO_9 (O_9,N_48752,N_48021);
or UO_10 (O_10,N_49664,N_49449);
and UO_11 (O_11,N_48766,N_49305);
xnor UO_12 (O_12,N_49836,N_48388);
nor UO_13 (O_13,N_48058,N_49719);
nand UO_14 (O_14,N_48070,N_49456);
and UO_15 (O_15,N_49620,N_48137);
and UO_16 (O_16,N_48528,N_49020);
and UO_17 (O_17,N_49961,N_49364);
nand UO_18 (O_18,N_49375,N_48973);
or UO_19 (O_19,N_49983,N_49991);
or UO_20 (O_20,N_49967,N_48158);
and UO_21 (O_21,N_48862,N_49532);
xnor UO_22 (O_22,N_48448,N_48564);
nand UO_23 (O_23,N_49731,N_48858);
xor UO_24 (O_24,N_48193,N_49433);
or UO_25 (O_25,N_49776,N_48823);
nor UO_26 (O_26,N_49277,N_48370);
xnor UO_27 (O_27,N_49469,N_48573);
nor UO_28 (O_28,N_48793,N_49885);
xnor UO_29 (O_29,N_48235,N_49622);
nor UO_30 (O_30,N_48553,N_49012);
or UO_31 (O_31,N_48611,N_49679);
or UO_32 (O_32,N_49058,N_48105);
nor UO_33 (O_33,N_49199,N_48969);
nand UO_34 (O_34,N_48727,N_49412);
or UO_35 (O_35,N_48183,N_49924);
nand UO_36 (O_36,N_48957,N_49558);
nor UO_37 (O_37,N_49554,N_49130);
or UO_38 (O_38,N_49703,N_49709);
nand UO_39 (O_39,N_48166,N_48508);
xnor UO_40 (O_40,N_48265,N_48861);
and UO_41 (O_41,N_48311,N_48459);
and UO_42 (O_42,N_48309,N_49318);
or UO_43 (O_43,N_49208,N_49292);
xor UO_44 (O_44,N_48250,N_48246);
nor UO_45 (O_45,N_49011,N_48118);
or UO_46 (O_46,N_49100,N_48418);
or UO_47 (O_47,N_49215,N_49720);
nor UO_48 (O_48,N_48652,N_48913);
nor UO_49 (O_49,N_49518,N_49394);
nand UO_50 (O_50,N_48542,N_49704);
and UO_51 (O_51,N_48147,N_49181);
nor UO_52 (O_52,N_49945,N_49052);
and UO_53 (O_53,N_48164,N_48461);
or UO_54 (O_54,N_49396,N_48980);
nand UO_55 (O_55,N_48574,N_49284);
nand UO_56 (O_56,N_48159,N_49663);
and UO_57 (O_57,N_48324,N_49116);
nor UO_58 (O_58,N_48753,N_48240);
nor UO_59 (O_59,N_49701,N_49085);
or UO_60 (O_60,N_48667,N_48067);
xnor UO_61 (O_61,N_49438,N_49078);
nor UO_62 (O_62,N_48956,N_48839);
and UO_63 (O_63,N_48682,N_49949);
nand UO_64 (O_64,N_49227,N_48502);
nand UO_65 (O_65,N_48944,N_49503);
and UO_66 (O_66,N_48500,N_48920);
xnor UO_67 (O_67,N_49281,N_49539);
nand UO_68 (O_68,N_49311,N_48884);
and UO_69 (O_69,N_49398,N_48199);
or UO_70 (O_70,N_49033,N_48571);
nand UO_71 (O_71,N_49431,N_48084);
and UO_72 (O_72,N_48287,N_49549);
xnor UO_73 (O_73,N_49126,N_48340);
or UO_74 (O_74,N_48840,N_48192);
or UO_75 (O_75,N_49470,N_49905);
and UO_76 (O_76,N_48045,N_48128);
nor UO_77 (O_77,N_48593,N_48748);
and UO_78 (O_78,N_48307,N_49040);
nor UO_79 (O_79,N_49948,N_49101);
xor UO_80 (O_80,N_48776,N_48316);
nand UO_81 (O_81,N_49560,N_48998);
nor UO_82 (O_82,N_49471,N_49342);
and UO_83 (O_83,N_49635,N_49441);
or UO_84 (O_84,N_49045,N_49128);
xnor UO_85 (O_85,N_48172,N_49520);
or UO_86 (O_86,N_48942,N_49804);
and UO_87 (O_87,N_48342,N_49616);
xnor UO_88 (O_88,N_49098,N_48229);
or UO_89 (O_89,N_49690,N_49829);
nor UO_90 (O_90,N_48296,N_48236);
or UO_91 (O_91,N_48596,N_48294);
xnor UO_92 (O_92,N_48297,N_49749);
nor UO_93 (O_93,N_48721,N_48904);
nor UO_94 (O_94,N_49504,N_48702);
nor UO_95 (O_95,N_48256,N_48946);
and UO_96 (O_96,N_48977,N_49397);
and UO_97 (O_97,N_48405,N_49510);
and UO_98 (O_98,N_49071,N_48962);
nand UO_99 (O_99,N_49573,N_48339);
or UO_100 (O_100,N_49632,N_49009);
nand UO_101 (O_101,N_49666,N_48640);
nand UO_102 (O_102,N_49958,N_48472);
nor UO_103 (O_103,N_48000,N_49330);
or UO_104 (O_104,N_48581,N_49337);
nand UO_105 (O_105,N_49737,N_49834);
nand UO_106 (O_106,N_49468,N_49132);
or UO_107 (O_107,N_49036,N_48919);
or UO_108 (O_108,N_48353,N_48313);
or UO_109 (O_109,N_49094,N_49800);
xnor UO_110 (O_110,N_49385,N_48486);
nor UO_111 (O_111,N_49773,N_49463);
nor UO_112 (O_112,N_48634,N_48974);
nor UO_113 (O_113,N_49236,N_48203);
nand UO_114 (O_114,N_48109,N_48756);
xnor UO_115 (O_115,N_49826,N_48444);
or UO_116 (O_116,N_49677,N_48874);
xor UO_117 (O_117,N_48879,N_48175);
nand UO_118 (O_118,N_48865,N_48781);
and UO_119 (O_119,N_49386,N_49741);
nor UO_120 (O_120,N_49574,N_48083);
xor UO_121 (O_121,N_48231,N_49321);
nor UO_122 (O_122,N_49575,N_49478);
nand UO_123 (O_123,N_48310,N_48018);
nor UO_124 (O_124,N_48849,N_49861);
xnor UO_125 (O_125,N_49700,N_48982);
nand UO_126 (O_126,N_49372,N_49633);
nand UO_127 (O_127,N_48411,N_49570);
nor UO_128 (O_128,N_48868,N_49395);
or UO_129 (O_129,N_49237,N_49524);
or UO_130 (O_130,N_49550,N_48619);
xor UO_131 (O_131,N_49498,N_48216);
and UO_132 (O_132,N_48715,N_49920);
nor UO_133 (O_133,N_49008,N_49260);
and UO_134 (O_134,N_48488,N_49147);
nor UO_135 (O_135,N_49043,N_48420);
nand UO_136 (O_136,N_48071,N_49895);
xnor UO_137 (O_137,N_48677,N_49336);
or UO_138 (O_138,N_49380,N_49865);
or UO_139 (O_139,N_49927,N_48419);
or UO_140 (O_140,N_49642,N_48037);
and UO_141 (O_141,N_49276,N_48271);
or UO_142 (O_142,N_48968,N_49686);
nand UO_143 (O_143,N_48487,N_49297);
and UO_144 (O_144,N_48604,N_49450);
or UO_145 (O_145,N_48774,N_49345);
nor UO_146 (O_146,N_48699,N_49367);
and UO_147 (O_147,N_49930,N_48632);
nor UO_148 (O_148,N_49087,N_49211);
nor UO_149 (O_149,N_48492,N_49073);
nand UO_150 (O_150,N_49739,N_49623);
nand UO_151 (O_151,N_48932,N_49628);
xnor UO_152 (O_152,N_49497,N_48556);
nand UO_153 (O_153,N_48538,N_49408);
nand UO_154 (O_154,N_49902,N_48790);
nor UO_155 (O_155,N_48938,N_48001);
and UO_156 (O_156,N_48114,N_49602);
nor UO_157 (O_157,N_49593,N_49348);
xor UO_158 (O_158,N_48269,N_49429);
xnor UO_159 (O_159,N_49951,N_49658);
and UO_160 (O_160,N_48559,N_48154);
or UO_161 (O_161,N_48377,N_48255);
nand UO_162 (O_162,N_49963,N_48941);
or UO_163 (O_163,N_49080,N_48873);
and UO_164 (O_164,N_49459,N_48156);
and UO_165 (O_165,N_49178,N_49555);
nand UO_166 (O_166,N_49840,N_49279);
nor UO_167 (O_167,N_48275,N_48078);
and UO_168 (O_168,N_48844,N_49392);
nor UO_169 (O_169,N_48964,N_49411);
nor UO_170 (O_170,N_49378,N_49577);
xnor UO_171 (O_171,N_48724,N_48767);
xor UO_172 (O_172,N_49695,N_48304);
nor UO_173 (O_173,N_49821,N_48945);
xor UO_174 (O_174,N_48856,N_48788);
xor UO_175 (O_175,N_48100,N_48253);
or UO_176 (O_176,N_48741,N_48952);
nor UO_177 (O_177,N_48585,N_49893);
and UO_178 (O_178,N_49476,N_48760);
nor UO_179 (O_179,N_48068,N_49979);
nor UO_180 (O_180,N_48273,N_48646);
nand UO_181 (O_181,N_49723,N_49494);
nor UO_182 (O_182,N_48155,N_48171);
xnor UO_183 (O_183,N_49377,N_49446);
xnor UO_184 (O_184,N_49595,N_49406);
xor UO_185 (O_185,N_48227,N_49886);
nor UO_186 (O_186,N_49047,N_49638);
and UO_187 (O_187,N_49858,N_49225);
xor UO_188 (O_188,N_49023,N_49994);
and UO_189 (O_189,N_48586,N_48570);
nand UO_190 (O_190,N_49486,N_49030);
nand UO_191 (O_191,N_49221,N_48030);
xnor UO_192 (O_192,N_49320,N_49822);
or UO_193 (O_193,N_48552,N_48055);
and UO_194 (O_194,N_49872,N_48117);
xnor UO_195 (O_195,N_49597,N_48582);
or UO_196 (O_196,N_49475,N_49598);
and UO_197 (O_197,N_49585,N_49608);
xnor UO_198 (O_198,N_49996,N_48735);
xnor UO_199 (O_199,N_48103,N_48771);
xnor UO_200 (O_200,N_48412,N_48916);
nor UO_201 (O_201,N_49485,N_48270);
xnor UO_202 (O_202,N_49940,N_48743);
nand UO_203 (O_203,N_49669,N_49452);
xnor UO_204 (O_204,N_49888,N_49261);
xnor UO_205 (O_205,N_49496,N_49136);
nor UO_206 (O_206,N_49481,N_49464);
nand UO_207 (O_207,N_49135,N_49877);
nor UO_208 (O_208,N_48762,N_48057);
and UO_209 (O_209,N_48807,N_48544);
xor UO_210 (O_210,N_48174,N_48140);
xnor UO_211 (O_211,N_48031,N_49744);
and UO_212 (O_212,N_49578,N_49247);
and UO_213 (O_213,N_48496,N_49767);
or UO_214 (O_214,N_49978,N_49316);
xnor UO_215 (O_215,N_49010,N_49420);
nand UO_216 (O_216,N_49892,N_48809);
and UO_217 (O_217,N_48098,N_48814);
and UO_218 (O_218,N_49610,N_48181);
nand UO_219 (O_219,N_48299,N_48643);
nand UO_220 (O_220,N_48734,N_48277);
xor UO_221 (O_221,N_48173,N_48737);
and UO_222 (O_222,N_49552,N_48020);
nor UO_223 (O_223,N_49519,N_48825);
or UO_224 (O_224,N_49137,N_49918);
and UO_225 (O_225,N_48097,N_49534);
xor UO_226 (O_226,N_48378,N_49661);
xor UO_227 (O_227,N_48723,N_48332);
or UO_228 (O_228,N_48738,N_48725);
nor UO_229 (O_229,N_49322,N_48579);
or UO_230 (O_230,N_49736,N_48594);
or UO_231 (O_231,N_49084,N_49809);
nor UO_232 (O_232,N_49748,N_49210);
xor UO_233 (O_233,N_49007,N_48708);
or UO_234 (O_234,N_48951,N_48575);
xnor UO_235 (O_235,N_49814,N_49625);
nor UO_236 (O_236,N_49454,N_48006);
nor UO_237 (O_237,N_49060,N_48930);
and UO_238 (O_238,N_49203,N_48426);
and UO_239 (O_239,N_48900,N_48428);
or UO_240 (O_240,N_49442,N_48606);
nand UO_241 (O_241,N_49989,N_48955);
nor UO_242 (O_242,N_48744,N_48683);
nand UO_243 (O_243,N_49567,N_49296);
xor UO_244 (O_244,N_48292,N_49660);
or UO_245 (O_245,N_49358,N_48341);
nand UO_246 (O_246,N_48794,N_48061);
nand UO_247 (O_247,N_48323,N_48449);
nor UO_248 (O_248,N_49584,N_49880);
nor UO_249 (O_249,N_48495,N_48222);
nand UO_250 (O_250,N_48731,N_49238);
or UO_251 (O_251,N_48751,N_49618);
xor UO_252 (O_252,N_48090,N_48554);
nor UO_253 (O_253,N_48764,N_49097);
xnor UO_254 (O_254,N_48934,N_48518);
xor UO_255 (O_255,N_49752,N_48303);
xor UO_256 (O_256,N_48654,N_49190);
nand UO_257 (O_257,N_49769,N_48168);
xnor UO_258 (O_258,N_48805,N_49721);
and UO_259 (O_259,N_48536,N_49757);
and UO_260 (O_260,N_48293,N_48681);
or UO_261 (O_261,N_49415,N_48890);
and UO_262 (O_262,N_48750,N_48369);
and UO_263 (O_263,N_48550,N_48950);
or UO_264 (O_264,N_48626,N_48434);
or UO_265 (O_265,N_49304,N_48600);
and UO_266 (O_266,N_48186,N_48768);
and UO_267 (O_267,N_48129,N_48692);
and UO_268 (O_268,N_49547,N_48926);
xor UO_269 (O_269,N_49566,N_49131);
and UO_270 (O_270,N_49596,N_49802);
nor UO_271 (O_271,N_49477,N_48792);
nand UO_272 (O_272,N_48623,N_49425);
nand UO_273 (O_273,N_49689,N_49646);
or UO_274 (O_274,N_49985,N_49529);
xnor UO_275 (O_275,N_49158,N_49956);
nor UO_276 (O_276,N_49545,N_49421);
nor UO_277 (O_277,N_49604,N_48985);
or UO_278 (O_278,N_49779,N_48897);
nand UO_279 (O_279,N_49523,N_48824);
or UO_280 (O_280,N_49806,N_48659);
nor UO_281 (O_281,N_49067,N_49670);
nor UO_282 (O_282,N_48565,N_48927);
and UO_283 (O_283,N_49344,N_48661);
xor UO_284 (O_284,N_49540,N_48870);
nand UO_285 (O_285,N_48679,N_48960);
nor UO_286 (O_286,N_49022,N_49359);
nor UO_287 (O_287,N_48249,N_49817);
or UO_288 (O_288,N_48170,N_48245);
nor UO_289 (O_289,N_49090,N_49837);
nand UO_290 (O_290,N_49460,N_49671);
and UO_291 (O_291,N_48241,N_49624);
xnor UO_292 (O_292,N_48772,N_48213);
xnor UO_293 (O_293,N_49026,N_48687);
and UO_294 (O_294,N_49838,N_49245);
nand UO_295 (O_295,N_48943,N_48330);
xnor UO_296 (O_296,N_49495,N_49059);
or UO_297 (O_297,N_49055,N_48069);
xor UO_298 (O_298,N_49995,N_49218);
nand UO_299 (O_299,N_49546,N_49946);
and UO_300 (O_300,N_48462,N_48288);
nand UO_301 (O_301,N_49735,N_48637);
and UO_302 (O_302,N_49264,N_48470);
and UO_303 (O_303,N_49964,N_48371);
or UO_304 (O_304,N_48163,N_48049);
and UO_305 (O_305,N_48456,N_49976);
nand UO_306 (O_306,N_48322,N_49650);
nor UO_307 (O_307,N_49465,N_49404);
xnor UO_308 (O_308,N_48473,N_48445);
and UO_309 (O_309,N_49427,N_48522);
or UO_310 (O_310,N_49751,N_48423);
and UO_311 (O_311,N_48655,N_48548);
xor UO_312 (O_312,N_49269,N_48914);
and UO_313 (O_313,N_48169,N_49122);
and UO_314 (O_314,N_49506,N_49353);
nand UO_315 (O_315,N_48523,N_49423);
nor UO_316 (O_316,N_48479,N_48491);
and UO_317 (O_317,N_49790,N_49799);
xnor UO_318 (O_318,N_49066,N_48123);
nor UO_319 (O_319,N_49298,N_48828);
and UO_320 (O_320,N_48628,N_49847);
nand UO_321 (O_321,N_48641,N_48335);
nor UO_322 (O_322,N_48736,N_49254);
nand UO_323 (O_323,N_48259,N_48427);
xor UO_324 (O_324,N_49244,N_48471);
or UO_325 (O_325,N_49656,N_48389);
nor UO_326 (O_326,N_49863,N_49490);
or UO_327 (O_327,N_49246,N_49416);
and UO_328 (O_328,N_48366,N_49160);
xnor UO_329 (O_329,N_48953,N_49763);
or UO_330 (O_330,N_49091,N_48887);
or UO_331 (O_331,N_48002,N_48132);
xor UO_332 (O_332,N_49301,N_48664);
xor UO_333 (O_333,N_49474,N_48875);
nand UO_334 (O_334,N_49157,N_48136);
nor UO_335 (O_335,N_48698,N_48223);
or UO_336 (O_336,N_49306,N_49874);
nand UO_337 (O_337,N_49155,N_48690);
nand UO_338 (O_338,N_48424,N_48761);
and UO_339 (O_339,N_48185,N_48546);
nand UO_340 (O_340,N_49017,N_48886);
or UO_341 (O_341,N_48688,N_48124);
or UO_342 (O_342,N_48605,N_48179);
nand UO_343 (O_343,N_48669,N_49413);
nor UO_344 (O_344,N_49729,N_49226);
nor UO_345 (O_345,N_48896,N_49070);
nor UO_346 (O_346,N_49370,N_49213);
and UO_347 (O_347,N_48379,N_48922);
or UO_348 (O_348,N_49734,N_48326);
nand UO_349 (O_349,N_48798,N_49876);
and UO_350 (O_350,N_48384,N_48499);
xor UO_351 (O_351,N_49207,N_49913);
and UO_352 (O_352,N_49232,N_49867);
or UO_353 (O_353,N_49031,N_49115);
or UO_354 (O_354,N_48120,N_48162);
nor UO_355 (O_355,N_48662,N_49681);
xnor UO_356 (O_356,N_49493,N_49153);
or UO_357 (O_357,N_48142,N_49069);
nor UO_358 (O_358,N_49326,N_49580);
nor UO_359 (O_359,N_49149,N_48407);
xnor UO_360 (O_360,N_49350,N_48622);
xor UO_361 (O_361,N_48718,N_48657);
nor UO_362 (O_362,N_49673,N_49038);
and UO_363 (O_363,N_48618,N_48693);
nand UO_364 (O_364,N_48048,N_49535);
and UO_365 (O_365,N_49630,N_49119);
nor UO_366 (O_366,N_48096,N_49708);
and UO_367 (O_367,N_48385,N_49177);
xor UO_368 (O_368,N_49592,N_49204);
xnor UO_369 (O_369,N_49166,N_49500);
nor UO_370 (O_370,N_48452,N_49252);
or UO_371 (O_371,N_49722,N_49374);
nand UO_372 (O_372,N_48433,N_48806);
or UO_373 (O_373,N_49368,N_49076);
nor UO_374 (O_374,N_49013,N_48054);
and UO_375 (O_375,N_49445,N_48242);
nand UO_376 (O_376,N_49791,N_48510);
nor UO_377 (O_377,N_49621,N_48355);
and UO_378 (O_378,N_49855,N_48899);
and UO_379 (O_379,N_48535,N_48838);
nand UO_380 (O_380,N_48613,N_48947);
nor UO_381 (O_381,N_48872,N_48075);
nor UO_382 (O_382,N_48441,N_49505);
and UO_383 (O_383,N_49201,N_48372);
or UO_384 (O_384,N_48961,N_49750);
and UO_385 (O_385,N_48810,N_49189);
xnor UO_386 (O_386,N_48220,N_48983);
xnor UO_387 (O_387,N_49228,N_48918);
and UO_388 (O_388,N_49113,N_48435);
or UO_389 (O_389,N_48547,N_48024);
or UO_390 (O_390,N_49167,N_48867);
xnor UO_391 (O_391,N_48038,N_48190);
xnor UO_392 (O_392,N_49600,N_49347);
xnor UO_393 (O_393,N_49831,N_48016);
nand UO_394 (O_394,N_48394,N_48328);
or UO_395 (O_395,N_49082,N_48134);
xnor UO_396 (O_396,N_48089,N_48033);
or UO_397 (O_397,N_48453,N_49356);
and UO_398 (O_398,N_48852,N_48785);
xnor UO_399 (O_399,N_49641,N_48184);
or UO_400 (O_400,N_49928,N_48976);
nor UO_401 (O_401,N_48144,N_48217);
xor UO_402 (O_402,N_49143,N_48885);
nand UO_403 (O_403,N_48836,N_49842);
nand UO_404 (O_404,N_49507,N_49125);
or UO_405 (O_405,N_48374,N_48397);
xnor UO_406 (O_406,N_48521,N_49962);
nand UO_407 (O_407,N_49453,N_49601);
or UO_408 (O_408,N_48381,N_49824);
nor UO_409 (O_409,N_48442,N_48315);
xor UO_410 (O_410,N_49970,N_48850);
or UO_411 (O_411,N_48759,N_49915);
nand UO_412 (O_412,N_49194,N_48300);
nand UO_413 (O_413,N_48219,N_49410);
nor UO_414 (O_414,N_49564,N_49127);
xor UO_415 (O_415,N_48940,N_49192);
xor UO_416 (O_416,N_49676,N_48795);
nand UO_417 (O_417,N_48458,N_49114);
xor UO_418 (O_418,N_49903,N_49340);
nor UO_419 (O_419,N_48933,N_49294);
and UO_420 (O_420,N_48221,N_49953);
and UO_421 (O_421,N_48531,N_49738);
nor UO_422 (O_422,N_48555,N_49852);
and UO_423 (O_423,N_48178,N_49175);
nor UO_424 (O_424,N_48333,N_49988);
nor UO_425 (O_425,N_49916,N_49768);
and UO_426 (O_426,N_48399,N_48032);
and UO_427 (O_427,N_49807,N_49662);
nand UO_428 (O_428,N_49401,N_49200);
nand UO_429 (O_429,N_49933,N_48653);
and UO_430 (O_430,N_49048,N_48530);
and UO_431 (O_431,N_49788,N_48029);
and UO_432 (O_432,N_48509,N_49846);
nor UO_433 (O_433,N_48023,N_49095);
xor UO_434 (O_434,N_48212,N_49766);
and UO_435 (O_435,N_49765,N_48966);
nand UO_436 (O_436,N_49243,N_48676);
xnor UO_437 (O_437,N_49212,N_48148);
nor UO_438 (O_438,N_49384,N_49430);
or UO_439 (O_439,N_49891,N_49096);
or UO_440 (O_440,N_48802,N_48855);
xor UO_441 (O_441,N_48276,N_48717);
nor UO_442 (O_442,N_49900,N_48046);
nor UO_443 (O_443,N_48770,N_48396);
and UO_444 (O_444,N_49382,N_49182);
or UO_445 (O_445,N_48638,N_48597);
and UO_446 (O_446,N_48714,N_49993);
nor UO_447 (O_447,N_48112,N_49636);
xnor UO_448 (O_448,N_48898,N_48232);
nand UO_449 (O_449,N_49492,N_49606);
xor UO_450 (O_450,N_48642,N_48505);
nor UO_451 (O_451,N_48912,N_48811);
nand UO_452 (O_452,N_48060,N_49974);
nor UO_453 (O_453,N_48414,N_49667);
nor UO_454 (O_454,N_48188,N_49777);
xnor UO_455 (O_455,N_48799,N_48206);
or UO_456 (O_456,N_48846,N_48413);
or UO_457 (O_457,N_48577,N_48077);
xor UO_458 (O_458,N_48895,N_49312);
nand UO_459 (O_459,N_48286,N_48877);
nor UO_460 (O_460,N_48258,N_49857);
nand UO_461 (O_461,N_48285,N_49527);
and UO_462 (O_462,N_48338,N_49141);
or UO_463 (O_463,N_49357,N_48238);
nand UO_464 (O_464,N_49883,N_48262);
xor UO_465 (O_465,N_48290,N_48935);
and UO_466 (O_466,N_48674,N_48254);
and UO_467 (O_467,N_49668,N_49742);
or UO_468 (O_468,N_48380,N_48189);
and UO_469 (O_469,N_48907,N_48549);
and UO_470 (O_470,N_49461,N_48678);
nand UO_471 (O_471,N_49145,N_49849);
xor UO_472 (O_472,N_48819,N_48387);
nand UO_473 (O_473,N_48386,N_49925);
and UO_474 (O_474,N_48383,N_49705);
nand UO_475 (O_475,N_48972,N_49890);
xor UO_476 (O_476,N_49665,N_49909);
nand UO_477 (O_477,N_48150,N_49025);
nand UO_478 (O_478,N_49004,N_49755);
xnor UO_479 (O_479,N_48636,N_49691);
and UO_480 (O_480,N_48513,N_48398);
nor UO_481 (O_481,N_48975,N_48589);
or UO_482 (O_482,N_49794,N_49054);
xor UO_483 (O_483,N_49583,N_48019);
nand UO_484 (O_484,N_49714,N_48620);
nand UO_485 (O_485,N_48039,N_48527);
and UO_486 (O_486,N_48517,N_48152);
nand UO_487 (O_487,N_48345,N_48034);
xnor UO_488 (O_488,N_48146,N_49812);
nand UO_489 (O_489,N_49062,N_49006);
xor UO_490 (O_490,N_48797,N_49365);
xnor UO_491 (O_491,N_48610,N_49980);
nand UO_492 (O_492,N_49869,N_49403);
and UO_493 (O_493,N_48247,N_48911);
and UO_494 (O_494,N_49936,N_49117);
nor UO_495 (O_495,N_48515,N_48291);
or UO_496 (O_496,N_48218,N_48337);
xor UO_497 (O_497,N_49355,N_49882);
and UO_498 (O_498,N_48466,N_49860);
xnor UO_499 (O_499,N_48194,N_48064);
nand UO_500 (O_500,N_48712,N_48161);
and UO_501 (O_501,N_48432,N_48463);
nor UO_502 (O_502,N_49309,N_48765);
and UO_503 (O_503,N_49253,N_49363);
and UO_504 (O_504,N_49576,N_48436);
xor UO_505 (O_505,N_49841,N_48325);
xnor UO_506 (O_506,N_48689,N_49693);
xor UO_507 (O_507,N_49144,N_48837);
xor UO_508 (O_508,N_49862,N_48889);
and UO_509 (O_509,N_49556,N_49816);
and UO_510 (O_510,N_49015,N_49644);
xor UO_511 (O_511,N_49557,N_48971);
or UO_512 (O_512,N_49609,N_48248);
nor UO_513 (O_513,N_48670,N_48431);
nand UO_514 (O_514,N_48393,N_48263);
nand UO_515 (O_515,N_49362,N_48214);
nor UO_516 (O_516,N_48780,N_48004);
and UO_517 (O_517,N_48860,N_48660);
and UO_518 (O_518,N_48949,N_48954);
nand UO_519 (O_519,N_48228,N_48126);
and UO_520 (O_520,N_48901,N_48005);
nor UO_521 (O_521,N_48224,N_48368);
nor UO_522 (O_522,N_49997,N_49255);
and UO_523 (O_523,N_48588,N_48131);
and UO_524 (O_524,N_49151,N_49832);
or UO_525 (O_525,N_48056,N_49057);
and UO_526 (O_526,N_48684,N_48994);
xor UO_527 (O_527,N_48503,N_49315);
xnor UO_528 (O_528,N_49267,N_49286);
xor UO_529 (O_529,N_48893,N_48672);
nor UO_530 (O_530,N_48314,N_48121);
nor UO_531 (O_531,N_49762,N_48266);
xnor UO_532 (O_532,N_49544,N_49195);
and UO_533 (O_533,N_48857,N_49634);
nor UO_534 (O_534,N_48821,N_48421);
and UO_535 (O_535,N_49789,N_48996);
xnor UO_536 (O_536,N_49103,N_49046);
xnor UO_537 (O_537,N_49682,N_49270);
or UO_538 (O_538,N_49110,N_49491);
nand UO_539 (O_539,N_48635,N_48864);
or UO_540 (O_540,N_48783,N_49850);
or UO_541 (O_541,N_49290,N_48361);
xor UO_542 (O_542,N_48826,N_48959);
nand UO_543 (O_543,N_49629,N_49075);
nor UO_544 (O_544,N_48784,N_48317);
xnor UO_545 (O_545,N_49399,N_48408);
and UO_546 (O_546,N_48696,N_48406);
and UO_547 (O_547,N_49257,N_49064);
and UO_548 (O_548,N_48451,N_48921);
or UO_549 (O_549,N_49698,N_48673);
nor UO_550 (O_550,N_49482,N_49121);
or UO_551 (O_551,N_48603,N_48624);
nor UO_552 (O_552,N_48382,N_48331);
or UO_553 (O_553,N_49922,N_48493);
and UO_554 (O_554,N_49639,N_49818);
nand UO_555 (O_555,N_48279,N_48177);
or UO_556 (O_556,N_49447,N_48481);
nand UO_557 (O_557,N_48167,N_48541);
or UO_558 (O_558,N_49265,N_49923);
nand UO_559 (O_559,N_49654,N_49259);
or UO_560 (O_560,N_48569,N_49473);
and UO_561 (O_561,N_48028,N_49907);
xor UO_562 (O_562,N_48835,N_48025);
and UO_563 (O_563,N_49233,N_48832);
nand UO_564 (O_564,N_48543,N_49917);
or UO_565 (O_565,N_49051,N_48373);
nand UO_566 (O_566,N_49581,N_48483);
xor UO_567 (O_567,N_48079,N_48252);
xnor UO_568 (O_568,N_48719,N_48349);
nand UO_569 (O_569,N_49152,N_48308);
nand UO_570 (O_570,N_48746,N_49437);
nand UO_571 (O_571,N_48022,N_49898);
nand UO_572 (O_572,N_48346,N_49754);
xor UO_573 (O_573,N_48376,N_49266);
nand UO_574 (O_574,N_48356,N_48512);
or UO_575 (O_575,N_49904,N_49934);
nor UO_576 (O_576,N_49422,N_48113);
xnor UO_577 (O_577,N_48145,N_48732);
or UO_578 (O_578,N_49373,N_48400);
and UO_579 (O_579,N_48602,N_48557);
nor UO_580 (O_580,N_48507,N_49439);
or UO_581 (O_581,N_49123,N_48409);
nand UO_582 (O_582,N_49513,N_48475);
xor UO_583 (O_583,N_49230,N_49746);
nand UO_584 (O_584,N_49220,N_48668);
xor UO_585 (O_585,N_48525,N_48931);
or UO_586 (O_586,N_49146,N_49740);
and UO_587 (O_587,N_48416,N_49998);
or UO_588 (O_588,N_49056,N_49548);
and UO_589 (O_589,N_49393,N_49982);
nor UO_590 (O_590,N_49615,N_48707);
nor UO_591 (O_591,N_49288,N_49448);
xnor UO_592 (O_592,N_48085,N_48576);
nand UO_593 (O_593,N_49165,N_49029);
and UO_594 (O_594,N_49972,N_48514);
nor UO_595 (O_595,N_49124,N_49896);
or UO_596 (O_596,N_49521,N_49879);
xnor UO_597 (O_597,N_48501,N_48474);
xnor UO_598 (O_598,N_49516,N_48281);
or UO_599 (O_599,N_49483,N_48990);
or UO_600 (O_600,N_48443,N_48243);
xor UO_601 (O_601,N_49018,N_49389);
nor UO_602 (O_602,N_49553,N_48995);
and UO_603 (O_603,N_48722,N_49436);
xor UO_604 (O_604,N_49159,N_49647);
xnor UO_605 (O_605,N_48204,N_49685);
xor UO_606 (O_606,N_49349,N_49835);
nor UO_607 (O_607,N_49955,N_49409);
nor UO_608 (O_608,N_49833,N_48730);
or UO_609 (O_609,N_49987,N_48711);
nand UO_610 (O_610,N_49875,N_49914);
xnor UO_611 (O_611,N_48319,N_48815);
or UO_612 (O_612,N_48239,N_49327);
and UO_613 (O_613,N_48978,N_48562);
and UO_614 (O_614,N_49037,N_48467);
nand UO_615 (O_615,N_48869,N_49263);
and UO_616 (O_616,N_49161,N_48305);
and UO_617 (O_617,N_49761,N_49783);
xor UO_618 (O_618,N_49774,N_48460);
xor UO_619 (O_619,N_49522,N_48320);
nor UO_620 (O_620,N_48430,N_49391);
or UO_621 (O_621,N_49871,N_49455);
nor UO_622 (O_622,N_48014,N_48534);
nor UO_623 (O_623,N_48043,N_49343);
nand UO_624 (O_624,N_49072,N_48631);
or UO_625 (O_625,N_49104,N_48524);
or UO_626 (O_626,N_48745,N_49889);
nor UO_627 (O_627,N_49319,N_48520);
and UO_628 (O_628,N_49919,N_48274);
nand UO_629 (O_629,N_48991,N_49371);
or UO_630 (O_630,N_48415,N_48044);
xor UO_631 (O_631,N_49688,N_49050);
and UO_632 (O_632,N_48205,N_49543);
or UO_633 (O_633,N_49614,N_48429);
and UO_634 (O_634,N_49792,N_48800);
nand UO_635 (O_635,N_49479,N_48648);
or UO_636 (O_636,N_49426,N_48110);
or UO_637 (O_637,N_48076,N_48257);
or UO_638 (O_638,N_49986,N_48260);
nand UO_639 (O_639,N_49517,N_49303);
xor UO_640 (O_640,N_49588,N_48011);
nand UO_641 (O_641,N_49659,N_48686);
or UO_642 (O_642,N_49133,N_49333);
nor UO_643 (O_643,N_48561,N_49864);
and UO_644 (O_644,N_49787,N_48695);
and UO_645 (O_645,N_49718,N_49901);
nor UO_646 (O_646,N_49960,N_48680);
or UO_647 (O_647,N_49106,N_49224);
or UO_648 (O_648,N_49950,N_49784);
and UO_649 (O_649,N_48560,N_48697);
xnor UO_650 (O_650,N_49981,N_49912);
and UO_651 (O_651,N_49275,N_49743);
and UO_652 (O_652,N_48758,N_49268);
xnor UO_653 (O_653,N_48883,N_48801);
nor UO_654 (O_654,N_48834,N_49713);
nand UO_655 (O_655,N_48244,N_48133);
nor UO_656 (O_656,N_49820,N_48348);
nand UO_657 (O_657,N_48747,N_48851);
or UO_658 (O_658,N_49331,N_48545);
and UO_659 (O_659,N_49188,N_49329);
and UO_660 (O_660,N_49771,N_49759);
nor UO_661 (O_661,N_48347,N_49458);
or UO_662 (O_662,N_48321,N_48958);
nor UO_663 (O_663,N_49262,N_49248);
and UO_664 (O_664,N_48970,N_48003);
xor UO_665 (O_665,N_48749,N_49594);
or UO_666 (O_666,N_48042,N_49674);
xnor UO_667 (O_667,N_49323,N_48876);
or UO_668 (O_668,N_48040,N_48568);
or UO_669 (O_669,N_49990,N_48902);
or UO_670 (O_670,N_49092,N_49354);
xnor UO_671 (O_671,N_48280,N_49590);
xnor UO_672 (O_672,N_48127,N_49702);
or UO_673 (O_673,N_48357,N_48139);
nand UO_674 (O_674,N_49587,N_48650);
or UO_675 (O_675,N_49139,N_48592);
and UO_676 (O_676,N_48656,N_48504);
xor UO_677 (O_677,N_49308,N_48352);
nand UO_678 (O_678,N_49250,N_49484);
xor UO_679 (O_679,N_48818,N_49241);
xor UO_680 (O_680,N_49489,N_49341);
xnor UO_681 (O_681,N_49870,N_49369);
and UO_682 (O_682,N_49651,N_49088);
nor UO_683 (O_683,N_49699,N_49339);
and UO_684 (O_684,N_49808,N_48583);
nand UO_685 (O_685,N_48306,N_49223);
nand UO_686 (O_686,N_48925,N_48842);
or UO_687 (O_687,N_49786,N_49440);
or UO_688 (O_688,N_48301,N_48122);
and UO_689 (O_689,N_48539,N_49878);
or UO_690 (O_690,N_48629,N_48267);
or UO_691 (O_691,N_49179,N_49335);
nand UO_692 (O_692,N_48666,N_49648);
and UO_693 (O_693,N_49801,N_48350);
nand UO_694 (O_694,N_49191,N_48910);
nor UO_695 (O_695,N_49003,N_49240);
xnor UO_696 (O_696,N_49525,N_48989);
xor UO_697 (O_697,N_48395,N_48278);
or UO_698 (O_698,N_49068,N_48465);
nand UO_699 (O_699,N_48027,N_49586);
or UO_700 (O_700,N_48295,N_48843);
or UO_701 (O_701,N_49512,N_48272);
and UO_702 (O_702,N_49019,N_49613);
and UO_703 (O_703,N_49351,N_49400);
nor UO_704 (O_704,N_48086,N_49005);
nor UO_705 (O_705,N_49291,N_49839);
and UO_706 (O_706,N_49111,N_49242);
xor UO_707 (O_707,N_48685,N_49039);
nor UO_708 (O_708,N_49280,N_49142);
xor UO_709 (O_709,N_48808,N_49173);
and UO_710 (O_710,N_49000,N_49187);
nor UO_711 (O_711,N_48391,N_48454);
or UO_712 (O_712,N_49387,N_48052);
and UO_713 (O_713,N_48477,N_49712);
nor UO_714 (O_714,N_49083,N_49845);
nand UO_715 (O_715,N_49637,N_49684);
nand UO_716 (O_716,N_48312,N_49795);
and UO_717 (O_717,N_48264,N_49197);
xnor UO_718 (O_718,N_49171,N_49944);
or UO_719 (O_719,N_49563,N_49844);
or UO_720 (O_720,N_48621,N_48180);
nor UO_721 (O_721,N_49533,N_48082);
and UO_722 (O_722,N_48095,N_49272);
nor UO_723 (O_723,N_48455,N_48967);
or UO_724 (O_724,N_49134,N_49383);
or UO_725 (O_725,N_48012,N_49975);
nor UO_726 (O_726,N_49725,N_49717);
xor UO_727 (O_727,N_49034,N_48644);
or UO_728 (O_728,N_48365,N_49065);
and UO_729 (O_729,N_48438,N_49672);
and UO_730 (O_730,N_48987,N_48859);
and UO_731 (O_731,N_48803,N_48208);
or UO_732 (O_732,N_48892,N_49899);
nor UO_733 (O_733,N_48363,N_48115);
nor UO_734 (O_734,N_48013,N_48820);
xor UO_735 (O_735,N_49172,N_49715);
nand UO_736 (O_736,N_48401,N_48529);
nand UO_737 (O_737,N_48237,N_48906);
nand UO_738 (O_738,N_48209,N_49764);
nand UO_739 (O_739,N_49617,N_49467);
nor UO_740 (O_740,N_48087,N_48074);
xnor UO_741 (O_741,N_49028,N_48187);
xor UO_742 (O_742,N_48457,N_48796);
and UO_743 (O_743,N_48567,N_49938);
nor UO_744 (O_744,N_49959,N_49696);
xnor UO_745 (O_745,N_49108,N_49174);
nand UO_746 (O_746,N_49234,N_49607);
nor UO_747 (O_747,N_48390,N_49079);
nor UO_748 (O_748,N_48062,N_48786);
nand UO_749 (O_749,N_48609,N_49655);
nor UO_750 (O_750,N_49205,N_48201);
and UO_751 (O_751,N_48773,N_49770);
or UO_752 (O_752,N_48367,N_49405);
or UO_753 (O_753,N_48354,N_49541);
nand UO_754 (O_754,N_49381,N_49077);
xnor UO_755 (O_755,N_48630,N_48791);
xnor UO_756 (O_756,N_49873,N_48234);
xor UO_757 (O_757,N_49217,N_49388);
nand UO_758 (O_758,N_48866,N_48404);
xor UO_759 (O_759,N_49251,N_49631);
xnor UO_760 (O_760,N_49733,N_49049);
and UO_761 (O_761,N_49813,N_49760);
nand UO_762 (O_762,N_49952,N_48847);
and UO_763 (O_763,N_49780,N_49605);
nor UO_764 (O_764,N_48489,N_48584);
and UO_765 (O_765,N_49680,N_49569);
or UO_766 (O_766,N_48817,N_49435);
nand UO_767 (O_767,N_49156,N_49035);
nand UO_768 (O_768,N_48986,N_49235);
and UO_769 (O_769,N_48871,N_48041);
nor UO_770 (O_770,N_49063,N_48997);
and UO_771 (O_771,N_48497,N_49118);
or UO_772 (O_772,N_49256,N_49775);
nand UO_773 (O_773,N_48853,N_49571);
or UO_774 (O_774,N_48706,N_48948);
or UO_775 (O_775,N_49612,N_49361);
nor UO_776 (O_776,N_48480,N_49216);
xor UO_777 (O_777,N_49848,N_48599);
or UO_778 (O_778,N_48739,N_48053);
or UO_779 (O_779,N_49120,N_49032);
nor UO_780 (O_780,N_48587,N_48880);
nor UO_781 (O_781,N_49856,N_48939);
xnor UO_782 (O_782,N_48563,N_48829);
xnor UO_783 (O_783,N_49793,N_48403);
xnor UO_784 (O_784,N_49154,N_49021);
nand UO_785 (O_785,N_48289,N_49678);
nor UO_786 (O_786,N_48035,N_48226);
or UO_787 (O_787,N_49511,N_48065);
and UO_788 (O_788,N_48375,N_49293);
or UO_789 (O_789,N_48813,N_49781);
xor UO_790 (O_790,N_48468,N_48268);
and UO_791 (O_791,N_49551,N_48111);
or UO_792 (O_792,N_49107,N_49697);
and UO_793 (O_793,N_49603,N_49488);
nor UO_794 (O_794,N_48963,N_49214);
or UO_795 (O_795,N_49390,N_48936);
nand UO_796 (O_796,N_49027,N_48908);
nor UO_797 (O_797,N_48905,N_49169);
or UO_798 (O_798,N_49324,N_49992);
xor UO_799 (O_799,N_49977,N_48537);
xor UO_800 (O_800,N_49501,N_49853);
or UO_801 (O_801,N_49528,N_48200);
nor UO_802 (O_802,N_48073,N_49163);
or UO_803 (O_803,N_49024,N_48845);
xor UO_804 (O_804,N_49745,N_49758);
xnor UO_805 (O_805,N_48720,N_49170);
nand UO_806 (O_806,N_49376,N_49530);
xnor UO_807 (O_807,N_49334,N_49536);
or UO_808 (O_808,N_49797,N_48733);
xor UO_809 (O_809,N_49942,N_48612);
nand UO_810 (O_810,N_48558,N_48318);
or UO_811 (O_811,N_49828,N_49999);
nand UO_812 (O_812,N_49911,N_49652);
and UO_813 (O_813,N_48782,N_49906);
or UO_814 (O_814,N_48233,N_48425);
xor UO_815 (O_815,N_48482,N_48437);
xor UO_816 (O_816,N_48284,N_49129);
and UO_817 (O_817,N_48165,N_49278);
or UO_818 (O_818,N_49868,N_49968);
nor UO_819 (O_819,N_48713,N_49803);
or UO_820 (O_820,N_48854,N_48026);
xnor UO_821 (O_821,N_49332,N_49640);
xor UO_822 (O_822,N_49014,N_49531);
and UO_823 (O_823,N_49089,N_49728);
xnor UO_824 (O_824,N_49526,N_49825);
xor UO_825 (O_825,N_48700,N_49202);
or UO_826 (O_826,N_49657,N_49407);
nor UO_827 (O_827,N_49138,N_48440);
and UO_828 (O_828,N_48891,N_48742);
nand UO_829 (O_829,N_48446,N_49086);
and UO_830 (O_830,N_48716,N_49105);
or UO_831 (O_831,N_49965,N_48965);
or UO_832 (O_832,N_48763,N_49894);
nor UO_833 (O_833,N_48775,N_48066);
nor UO_834 (O_834,N_49093,N_49307);
or UO_835 (O_835,N_48225,N_49074);
xnor UO_836 (O_836,N_49866,N_49206);
and UO_837 (O_837,N_48007,N_48017);
or UO_838 (O_838,N_48777,N_49249);
or UO_839 (O_839,N_49184,N_49694);
nand UO_840 (O_840,N_48494,N_48757);
xnor UO_841 (O_841,N_48207,N_49001);
and UO_842 (O_842,N_49346,N_49258);
and UO_843 (O_843,N_48848,N_48344);
and UO_844 (O_844,N_48080,N_48984);
xor UO_845 (O_845,N_49611,N_48081);
xnor UO_846 (O_846,N_48726,N_48691);
nor UO_847 (O_847,N_48615,N_48108);
or UO_848 (O_848,N_48362,N_49325);
or UO_849 (O_849,N_48130,N_48647);
or UO_850 (O_850,N_48476,N_48703);
or UO_851 (O_851,N_49941,N_49626);
nand UO_852 (O_852,N_48094,N_49957);
and UO_853 (O_853,N_49379,N_49414);
nor UO_854 (O_854,N_48093,N_49289);
nor UO_855 (O_855,N_48616,N_49823);
xor UO_856 (O_856,N_48625,N_49724);
xnor UO_857 (O_857,N_49772,N_48671);
nand UO_858 (O_858,N_48580,N_49675);
nor UO_859 (O_859,N_49061,N_49811);
or UO_860 (O_860,N_48658,N_49239);
xor UO_861 (O_861,N_49931,N_49854);
xnor UO_862 (O_862,N_49572,N_48804);
and UO_863 (O_863,N_48572,N_48816);
and UO_864 (O_864,N_48336,N_48215);
xor UO_865 (O_865,N_48063,N_48135);
or UO_866 (O_866,N_48511,N_48182);
nor UO_867 (O_867,N_49285,N_49538);
and UO_868 (O_868,N_49314,N_49711);
or UO_869 (O_869,N_48779,N_48450);
nand UO_870 (O_870,N_49317,N_49947);
nand UO_871 (O_871,N_48729,N_49559);
or UO_872 (O_872,N_49537,N_49428);
or UO_873 (O_873,N_48261,N_49683);
xnor UO_874 (O_874,N_49910,N_48036);
nand UO_875 (O_875,N_49271,N_49935);
nand UO_876 (O_876,N_48447,N_48211);
or UO_877 (O_877,N_48047,N_48532);
and UO_878 (O_878,N_48051,N_48519);
nor UO_879 (O_879,N_48059,N_49112);
and UO_880 (O_880,N_49109,N_49732);
and UO_881 (O_881,N_49599,N_48099);
nand UO_882 (O_882,N_48198,N_48981);
nor UO_883 (O_883,N_48651,N_49984);
nor UO_884 (O_884,N_49041,N_48009);
and UO_885 (O_885,N_49499,N_49451);
nor UO_886 (O_886,N_49619,N_49219);
nand UO_887 (O_887,N_49196,N_49810);
nor UO_888 (O_888,N_49418,N_48088);
nor UO_889 (O_889,N_49487,N_49884);
and UO_890 (O_890,N_49222,N_49706);
and UO_891 (O_891,N_49366,N_49419);
and UO_892 (O_892,N_48881,N_49360);
or UO_893 (O_893,N_49778,N_49726);
xor UO_894 (O_894,N_49424,N_48485);
and UO_895 (O_895,N_48464,N_48812);
nand UO_896 (O_896,N_49053,N_48993);
or UO_897 (O_897,N_48841,N_49627);
and UO_898 (O_898,N_49502,N_49582);
nand UO_899 (O_899,N_49148,N_48010);
xnor UO_900 (O_900,N_49649,N_49932);
or UO_901 (O_901,N_48551,N_48402);
xor UO_902 (O_902,N_49273,N_49282);
or UO_903 (O_903,N_48608,N_48329);
nor UO_904 (O_904,N_48822,N_49937);
xor UO_905 (O_905,N_49565,N_48104);
nand UO_906 (O_906,N_48705,N_48778);
nand UO_907 (O_907,N_49162,N_49186);
nor UO_908 (O_908,N_49287,N_48915);
xnor UO_909 (O_909,N_49954,N_48141);
xor UO_910 (O_910,N_48863,N_48665);
nand UO_911 (O_911,N_48138,N_49042);
xor UO_912 (O_912,N_48498,N_49231);
and UO_913 (O_913,N_49881,N_49645);
and UO_914 (O_914,N_48302,N_48283);
or UO_915 (O_915,N_49710,N_49589);
xnor UO_916 (O_916,N_49444,N_48143);
or UO_917 (O_917,N_49081,N_48903);
nand UO_918 (O_918,N_49542,N_48191);
and UO_919 (O_919,N_49859,N_48417);
and UO_920 (O_920,N_49747,N_48917);
and UO_921 (O_921,N_49908,N_48831);
xor UO_922 (O_922,N_49727,N_48359);
and UO_923 (O_923,N_49782,N_48789);
and UO_924 (O_924,N_49568,N_48639);
or UO_925 (O_925,N_49164,N_49302);
and UO_926 (O_926,N_48533,N_49209);
or UO_927 (O_927,N_48578,N_49313);
or UO_928 (O_928,N_49274,N_48929);
or UO_929 (O_929,N_49796,N_49310);
nand UO_930 (O_930,N_48422,N_49798);
nor UO_931 (O_931,N_49643,N_49328);
or UO_932 (O_932,N_48478,N_48526);
nand UO_933 (O_933,N_48710,N_48878);
and UO_934 (O_934,N_49515,N_49753);
and UO_935 (O_935,N_48119,N_49338);
or UO_936 (O_936,N_49352,N_49168);
xor UO_937 (O_937,N_48704,N_48540);
or UO_938 (O_938,N_49480,N_49843);
xor UO_939 (O_939,N_49176,N_49002);
nor UO_940 (O_940,N_49707,N_49508);
nor UO_941 (O_941,N_48092,N_48210);
xor UO_942 (O_942,N_49819,N_48649);
or UO_943 (O_943,N_48769,N_48728);
nor UO_944 (O_944,N_48196,N_49579);
and UO_945 (O_945,N_49939,N_49815);
nor UO_946 (O_946,N_48614,N_48627);
nor UO_947 (O_947,N_48251,N_48999);
nor UO_948 (O_948,N_49830,N_49099);
or UO_949 (O_949,N_49102,N_49562);
or UO_950 (O_950,N_48015,N_48992);
nor UO_951 (O_951,N_48153,N_48101);
or UO_952 (O_952,N_49785,N_49971);
and UO_953 (O_953,N_48358,N_48195);
or UO_954 (O_954,N_48833,N_48392);
nand UO_955 (O_955,N_49150,N_49756);
and UO_956 (O_956,N_48343,N_48924);
nand UO_957 (O_957,N_49966,N_49283);
nand UO_958 (O_958,N_49457,N_48360);
and UO_959 (O_959,N_48102,N_48591);
or UO_960 (O_960,N_48125,N_49591);
and UO_961 (O_961,N_49653,N_49417);
and UO_962 (O_962,N_49300,N_48230);
xnor UO_963 (O_963,N_48107,N_49185);
xor UO_964 (O_964,N_48590,N_48116);
xnor UO_965 (O_965,N_49687,N_48008);
nor UO_966 (O_966,N_49509,N_48157);
nor UO_967 (O_967,N_48506,N_48202);
and UO_968 (O_968,N_49443,N_49434);
or UO_969 (O_969,N_48701,N_48327);
or UO_970 (O_970,N_49514,N_48645);
xnor UO_971 (O_971,N_49943,N_48988);
or UO_972 (O_972,N_48709,N_49299);
xnor UO_973 (O_973,N_49193,N_48923);
nor UO_974 (O_974,N_48888,N_48937);
and UO_975 (O_975,N_48663,N_49183);
nor UO_976 (O_976,N_48830,N_49432);
xnor UO_977 (O_977,N_48160,N_48298);
xor UO_978 (O_978,N_49921,N_49716);
xnor UO_979 (O_979,N_48439,N_48787);
or UO_980 (O_980,N_49929,N_49016);
or UO_981 (O_981,N_49926,N_48633);
nor UO_982 (O_982,N_48176,N_48050);
and UO_983 (O_983,N_49472,N_49044);
and UO_984 (O_984,N_49466,N_48490);
nor UO_985 (O_985,N_49692,N_48469);
nor UO_986 (O_986,N_48740,N_49730);
nand UO_987 (O_987,N_48928,N_49887);
nor UO_988 (O_988,N_48566,N_48410);
nor UO_989 (O_989,N_48484,N_48151);
xnor UO_990 (O_990,N_49180,N_48601);
and UO_991 (O_991,N_49973,N_49969);
and UO_992 (O_992,N_49827,N_49229);
and UO_993 (O_993,N_49561,N_48755);
nand UO_994 (O_994,N_48617,N_48149);
nand UO_995 (O_995,N_49295,N_49402);
or UO_996 (O_996,N_48827,N_49897);
or UO_997 (O_997,N_48979,N_48607);
or UO_998 (O_998,N_48754,N_48598);
nor UO_999 (O_999,N_49805,N_48516);
xnor UO_1000 (O_1000,N_48665,N_48116);
or UO_1001 (O_1001,N_48759,N_48188);
or UO_1002 (O_1002,N_49397,N_49274);
or UO_1003 (O_1003,N_49502,N_49038);
or UO_1004 (O_1004,N_48304,N_48007);
xor UO_1005 (O_1005,N_48351,N_48224);
or UO_1006 (O_1006,N_48643,N_48528);
and UO_1007 (O_1007,N_48617,N_49277);
xor UO_1008 (O_1008,N_48361,N_49514);
nor UO_1009 (O_1009,N_49417,N_49126);
and UO_1010 (O_1010,N_48070,N_48065);
or UO_1011 (O_1011,N_48454,N_49870);
nor UO_1012 (O_1012,N_49015,N_48209);
and UO_1013 (O_1013,N_48811,N_49108);
xnor UO_1014 (O_1014,N_48456,N_48245);
or UO_1015 (O_1015,N_48375,N_49112);
or UO_1016 (O_1016,N_48345,N_49331);
nor UO_1017 (O_1017,N_49643,N_49414);
xor UO_1018 (O_1018,N_49933,N_48538);
nand UO_1019 (O_1019,N_49403,N_49509);
nor UO_1020 (O_1020,N_49445,N_49664);
or UO_1021 (O_1021,N_48986,N_49608);
and UO_1022 (O_1022,N_48474,N_49163);
or UO_1023 (O_1023,N_49640,N_49249);
xor UO_1024 (O_1024,N_48281,N_48720);
or UO_1025 (O_1025,N_48857,N_49186);
nand UO_1026 (O_1026,N_49189,N_49209);
and UO_1027 (O_1027,N_49007,N_48791);
nor UO_1028 (O_1028,N_48521,N_48107);
xor UO_1029 (O_1029,N_49996,N_48521);
or UO_1030 (O_1030,N_48871,N_48547);
nand UO_1031 (O_1031,N_48671,N_48794);
nand UO_1032 (O_1032,N_48388,N_49303);
nor UO_1033 (O_1033,N_49014,N_49927);
or UO_1034 (O_1034,N_49727,N_49776);
nand UO_1035 (O_1035,N_49195,N_49509);
xnor UO_1036 (O_1036,N_48647,N_49287);
nor UO_1037 (O_1037,N_49286,N_48231);
xor UO_1038 (O_1038,N_48106,N_48694);
nor UO_1039 (O_1039,N_49442,N_49102);
xnor UO_1040 (O_1040,N_48227,N_48867);
xor UO_1041 (O_1041,N_49823,N_48816);
nor UO_1042 (O_1042,N_48094,N_49482);
or UO_1043 (O_1043,N_49709,N_49947);
or UO_1044 (O_1044,N_48058,N_49152);
xor UO_1045 (O_1045,N_48683,N_48660);
or UO_1046 (O_1046,N_48401,N_48691);
xor UO_1047 (O_1047,N_48294,N_49359);
or UO_1048 (O_1048,N_49679,N_49636);
nand UO_1049 (O_1049,N_49661,N_48259);
and UO_1050 (O_1050,N_49477,N_49577);
or UO_1051 (O_1051,N_49755,N_48283);
and UO_1052 (O_1052,N_48888,N_48701);
nand UO_1053 (O_1053,N_49610,N_48510);
nand UO_1054 (O_1054,N_49133,N_49856);
and UO_1055 (O_1055,N_49599,N_48030);
nand UO_1056 (O_1056,N_48412,N_48066);
xor UO_1057 (O_1057,N_48263,N_48760);
nand UO_1058 (O_1058,N_49994,N_49108);
nand UO_1059 (O_1059,N_49434,N_49433);
or UO_1060 (O_1060,N_48742,N_49952);
nor UO_1061 (O_1061,N_49489,N_49457);
nand UO_1062 (O_1062,N_49533,N_48812);
nor UO_1063 (O_1063,N_48367,N_49279);
and UO_1064 (O_1064,N_48137,N_49869);
nand UO_1065 (O_1065,N_48313,N_48603);
xor UO_1066 (O_1066,N_49513,N_49059);
xnor UO_1067 (O_1067,N_48870,N_49951);
or UO_1068 (O_1068,N_49763,N_48033);
xnor UO_1069 (O_1069,N_49421,N_48532);
nor UO_1070 (O_1070,N_48158,N_49120);
nand UO_1071 (O_1071,N_49850,N_49365);
and UO_1072 (O_1072,N_48771,N_49361);
nor UO_1073 (O_1073,N_49905,N_48764);
or UO_1074 (O_1074,N_48321,N_48366);
nor UO_1075 (O_1075,N_49525,N_49892);
and UO_1076 (O_1076,N_49590,N_48108);
and UO_1077 (O_1077,N_48814,N_48292);
and UO_1078 (O_1078,N_49494,N_48770);
nor UO_1079 (O_1079,N_48862,N_48311);
nor UO_1080 (O_1080,N_48352,N_49888);
nand UO_1081 (O_1081,N_48922,N_48338);
nor UO_1082 (O_1082,N_49185,N_48375);
or UO_1083 (O_1083,N_48673,N_48550);
and UO_1084 (O_1084,N_48200,N_49204);
xnor UO_1085 (O_1085,N_48820,N_48158);
or UO_1086 (O_1086,N_49680,N_48213);
nand UO_1087 (O_1087,N_49125,N_48361);
nand UO_1088 (O_1088,N_48873,N_49310);
xor UO_1089 (O_1089,N_49064,N_49470);
nor UO_1090 (O_1090,N_48389,N_48494);
nand UO_1091 (O_1091,N_49497,N_48434);
nor UO_1092 (O_1092,N_49828,N_48097);
xnor UO_1093 (O_1093,N_49715,N_49807);
nand UO_1094 (O_1094,N_49490,N_49325);
xor UO_1095 (O_1095,N_49069,N_49635);
nand UO_1096 (O_1096,N_49196,N_49822);
and UO_1097 (O_1097,N_49428,N_49463);
or UO_1098 (O_1098,N_48102,N_49296);
xnor UO_1099 (O_1099,N_48419,N_48163);
xor UO_1100 (O_1100,N_48872,N_49685);
xor UO_1101 (O_1101,N_48200,N_48832);
nand UO_1102 (O_1102,N_48335,N_48929);
or UO_1103 (O_1103,N_49805,N_48120);
nor UO_1104 (O_1104,N_48260,N_49969);
or UO_1105 (O_1105,N_48602,N_49727);
or UO_1106 (O_1106,N_49245,N_48787);
or UO_1107 (O_1107,N_49481,N_49973);
and UO_1108 (O_1108,N_48848,N_48773);
xor UO_1109 (O_1109,N_48084,N_49020);
xnor UO_1110 (O_1110,N_48902,N_49654);
and UO_1111 (O_1111,N_49922,N_48770);
and UO_1112 (O_1112,N_48538,N_49508);
and UO_1113 (O_1113,N_49790,N_49876);
xnor UO_1114 (O_1114,N_48584,N_49228);
xnor UO_1115 (O_1115,N_48904,N_48718);
and UO_1116 (O_1116,N_48310,N_49064);
nor UO_1117 (O_1117,N_49615,N_49965);
or UO_1118 (O_1118,N_48802,N_49231);
and UO_1119 (O_1119,N_49914,N_49159);
or UO_1120 (O_1120,N_48448,N_48748);
nor UO_1121 (O_1121,N_49474,N_48368);
or UO_1122 (O_1122,N_49634,N_49309);
and UO_1123 (O_1123,N_49360,N_49425);
or UO_1124 (O_1124,N_48868,N_48688);
nand UO_1125 (O_1125,N_48768,N_48683);
nor UO_1126 (O_1126,N_48032,N_49985);
xor UO_1127 (O_1127,N_49528,N_48956);
xor UO_1128 (O_1128,N_49771,N_49988);
or UO_1129 (O_1129,N_49332,N_49177);
nand UO_1130 (O_1130,N_48279,N_48903);
nand UO_1131 (O_1131,N_49799,N_49970);
and UO_1132 (O_1132,N_49189,N_49153);
and UO_1133 (O_1133,N_48868,N_48042);
xor UO_1134 (O_1134,N_48043,N_49968);
xnor UO_1135 (O_1135,N_49075,N_49339);
nand UO_1136 (O_1136,N_48629,N_49909);
nor UO_1137 (O_1137,N_48274,N_48158);
or UO_1138 (O_1138,N_48832,N_48674);
or UO_1139 (O_1139,N_48467,N_48382);
or UO_1140 (O_1140,N_48980,N_48869);
and UO_1141 (O_1141,N_48174,N_49122);
nor UO_1142 (O_1142,N_48944,N_49173);
xnor UO_1143 (O_1143,N_49886,N_48187);
nand UO_1144 (O_1144,N_49150,N_48113);
nor UO_1145 (O_1145,N_48105,N_48225);
xnor UO_1146 (O_1146,N_48861,N_48530);
xnor UO_1147 (O_1147,N_48697,N_48520);
xnor UO_1148 (O_1148,N_48607,N_48757);
xnor UO_1149 (O_1149,N_48762,N_48140);
and UO_1150 (O_1150,N_48362,N_48993);
nand UO_1151 (O_1151,N_49971,N_49960);
or UO_1152 (O_1152,N_48080,N_49472);
nor UO_1153 (O_1153,N_48704,N_49848);
nor UO_1154 (O_1154,N_49399,N_49457);
and UO_1155 (O_1155,N_49479,N_49597);
nor UO_1156 (O_1156,N_49509,N_48659);
or UO_1157 (O_1157,N_49270,N_48524);
and UO_1158 (O_1158,N_48711,N_49944);
nor UO_1159 (O_1159,N_48827,N_49840);
or UO_1160 (O_1160,N_49589,N_49648);
nor UO_1161 (O_1161,N_49845,N_48605);
nand UO_1162 (O_1162,N_49421,N_48544);
nand UO_1163 (O_1163,N_49004,N_48687);
xnor UO_1164 (O_1164,N_48154,N_48181);
xnor UO_1165 (O_1165,N_49079,N_49311);
or UO_1166 (O_1166,N_48427,N_49505);
nor UO_1167 (O_1167,N_48840,N_49768);
nor UO_1168 (O_1168,N_49788,N_49396);
nand UO_1169 (O_1169,N_49876,N_49826);
nand UO_1170 (O_1170,N_49847,N_48236);
nand UO_1171 (O_1171,N_49477,N_48401);
xor UO_1172 (O_1172,N_48540,N_48899);
nor UO_1173 (O_1173,N_48059,N_49073);
xnor UO_1174 (O_1174,N_48022,N_49385);
or UO_1175 (O_1175,N_49727,N_48254);
xor UO_1176 (O_1176,N_49034,N_48994);
and UO_1177 (O_1177,N_48628,N_49851);
xnor UO_1178 (O_1178,N_49539,N_49959);
nor UO_1179 (O_1179,N_49348,N_49212);
and UO_1180 (O_1180,N_49558,N_49294);
and UO_1181 (O_1181,N_49059,N_49435);
or UO_1182 (O_1182,N_49225,N_48875);
or UO_1183 (O_1183,N_49575,N_48476);
nand UO_1184 (O_1184,N_49644,N_48142);
and UO_1185 (O_1185,N_48061,N_48588);
xnor UO_1186 (O_1186,N_49796,N_48686);
nand UO_1187 (O_1187,N_48541,N_48506);
xnor UO_1188 (O_1188,N_48054,N_49571);
and UO_1189 (O_1189,N_49591,N_48885);
nand UO_1190 (O_1190,N_49722,N_48577);
xor UO_1191 (O_1191,N_49235,N_48453);
xor UO_1192 (O_1192,N_49090,N_49791);
xnor UO_1193 (O_1193,N_48542,N_49673);
xnor UO_1194 (O_1194,N_48180,N_48619);
and UO_1195 (O_1195,N_49401,N_48024);
nor UO_1196 (O_1196,N_48189,N_48616);
and UO_1197 (O_1197,N_48501,N_49084);
nand UO_1198 (O_1198,N_48588,N_49283);
nand UO_1199 (O_1199,N_48905,N_48127);
and UO_1200 (O_1200,N_49090,N_48759);
and UO_1201 (O_1201,N_49033,N_49307);
or UO_1202 (O_1202,N_48425,N_48175);
nor UO_1203 (O_1203,N_48471,N_49993);
and UO_1204 (O_1204,N_49720,N_49730);
xor UO_1205 (O_1205,N_48025,N_48127);
and UO_1206 (O_1206,N_48245,N_49175);
or UO_1207 (O_1207,N_48922,N_48106);
or UO_1208 (O_1208,N_48955,N_48518);
and UO_1209 (O_1209,N_48396,N_49225);
nand UO_1210 (O_1210,N_48356,N_48608);
or UO_1211 (O_1211,N_48992,N_49347);
and UO_1212 (O_1212,N_48473,N_49772);
xnor UO_1213 (O_1213,N_49721,N_49379);
xor UO_1214 (O_1214,N_49811,N_49671);
and UO_1215 (O_1215,N_48052,N_48773);
nand UO_1216 (O_1216,N_48348,N_49660);
xnor UO_1217 (O_1217,N_48314,N_49609);
nand UO_1218 (O_1218,N_48431,N_49143);
or UO_1219 (O_1219,N_49152,N_49573);
xnor UO_1220 (O_1220,N_48022,N_48773);
xor UO_1221 (O_1221,N_49315,N_49558);
and UO_1222 (O_1222,N_48074,N_49375);
or UO_1223 (O_1223,N_48954,N_48767);
xor UO_1224 (O_1224,N_48048,N_48036);
nand UO_1225 (O_1225,N_48191,N_49132);
and UO_1226 (O_1226,N_49506,N_48600);
xnor UO_1227 (O_1227,N_48101,N_49817);
nand UO_1228 (O_1228,N_48752,N_48665);
nor UO_1229 (O_1229,N_49988,N_48073);
or UO_1230 (O_1230,N_49432,N_48360);
or UO_1231 (O_1231,N_48034,N_48733);
or UO_1232 (O_1232,N_48448,N_49190);
or UO_1233 (O_1233,N_49462,N_49319);
xnor UO_1234 (O_1234,N_49044,N_48551);
and UO_1235 (O_1235,N_48085,N_49379);
xnor UO_1236 (O_1236,N_49539,N_49890);
or UO_1237 (O_1237,N_49952,N_49951);
xnor UO_1238 (O_1238,N_49984,N_48006);
nor UO_1239 (O_1239,N_48217,N_48392);
and UO_1240 (O_1240,N_48846,N_49361);
xor UO_1241 (O_1241,N_49415,N_49524);
nor UO_1242 (O_1242,N_49726,N_49958);
xnor UO_1243 (O_1243,N_49605,N_48208);
and UO_1244 (O_1244,N_48469,N_48385);
xnor UO_1245 (O_1245,N_48766,N_49292);
nor UO_1246 (O_1246,N_49360,N_49368);
xor UO_1247 (O_1247,N_48008,N_48531);
and UO_1248 (O_1248,N_49763,N_48702);
nor UO_1249 (O_1249,N_49154,N_49923);
nor UO_1250 (O_1250,N_49028,N_49797);
nor UO_1251 (O_1251,N_48551,N_49620);
or UO_1252 (O_1252,N_49892,N_49391);
nor UO_1253 (O_1253,N_48412,N_48206);
and UO_1254 (O_1254,N_49538,N_49800);
or UO_1255 (O_1255,N_49168,N_49162);
xnor UO_1256 (O_1256,N_48897,N_49822);
nand UO_1257 (O_1257,N_48976,N_49064);
nor UO_1258 (O_1258,N_48619,N_49255);
nor UO_1259 (O_1259,N_48556,N_49504);
nand UO_1260 (O_1260,N_48657,N_48559);
nand UO_1261 (O_1261,N_49781,N_49596);
xnor UO_1262 (O_1262,N_48742,N_49933);
or UO_1263 (O_1263,N_48100,N_49980);
nor UO_1264 (O_1264,N_49493,N_49686);
xor UO_1265 (O_1265,N_49771,N_48035);
xor UO_1266 (O_1266,N_48340,N_48425);
and UO_1267 (O_1267,N_48693,N_49434);
or UO_1268 (O_1268,N_48281,N_49920);
and UO_1269 (O_1269,N_48115,N_48204);
and UO_1270 (O_1270,N_49412,N_48787);
xnor UO_1271 (O_1271,N_49654,N_49711);
or UO_1272 (O_1272,N_48482,N_48069);
nor UO_1273 (O_1273,N_49441,N_49861);
xnor UO_1274 (O_1274,N_48081,N_48747);
xnor UO_1275 (O_1275,N_48671,N_49748);
xnor UO_1276 (O_1276,N_48824,N_48383);
or UO_1277 (O_1277,N_48553,N_48445);
nand UO_1278 (O_1278,N_48365,N_49706);
and UO_1279 (O_1279,N_48213,N_49645);
or UO_1280 (O_1280,N_48551,N_48716);
xnor UO_1281 (O_1281,N_49623,N_48077);
nand UO_1282 (O_1282,N_48944,N_49809);
xor UO_1283 (O_1283,N_49722,N_49602);
or UO_1284 (O_1284,N_48284,N_49342);
or UO_1285 (O_1285,N_49625,N_48360);
nand UO_1286 (O_1286,N_49150,N_49675);
and UO_1287 (O_1287,N_49507,N_49523);
and UO_1288 (O_1288,N_49225,N_48991);
nor UO_1289 (O_1289,N_49398,N_48103);
nand UO_1290 (O_1290,N_49569,N_48417);
nand UO_1291 (O_1291,N_48513,N_48184);
and UO_1292 (O_1292,N_49910,N_48602);
and UO_1293 (O_1293,N_49524,N_49023);
nand UO_1294 (O_1294,N_48587,N_49205);
or UO_1295 (O_1295,N_49054,N_49776);
or UO_1296 (O_1296,N_49430,N_48943);
or UO_1297 (O_1297,N_48105,N_48900);
and UO_1298 (O_1298,N_48391,N_49704);
and UO_1299 (O_1299,N_48666,N_48091);
xnor UO_1300 (O_1300,N_49946,N_48307);
nand UO_1301 (O_1301,N_49207,N_48349);
nor UO_1302 (O_1302,N_49666,N_48610);
or UO_1303 (O_1303,N_48602,N_48673);
or UO_1304 (O_1304,N_48863,N_48164);
nor UO_1305 (O_1305,N_49845,N_48052);
or UO_1306 (O_1306,N_49277,N_48049);
nand UO_1307 (O_1307,N_49587,N_48278);
nand UO_1308 (O_1308,N_49714,N_49165);
xnor UO_1309 (O_1309,N_49257,N_48547);
and UO_1310 (O_1310,N_48062,N_49602);
and UO_1311 (O_1311,N_48517,N_49931);
xnor UO_1312 (O_1312,N_48883,N_48531);
nand UO_1313 (O_1313,N_48740,N_48892);
nor UO_1314 (O_1314,N_49204,N_48287);
and UO_1315 (O_1315,N_49685,N_49183);
nand UO_1316 (O_1316,N_49529,N_48992);
or UO_1317 (O_1317,N_49798,N_48515);
and UO_1318 (O_1318,N_49827,N_49936);
nor UO_1319 (O_1319,N_48333,N_49119);
or UO_1320 (O_1320,N_49984,N_48170);
and UO_1321 (O_1321,N_49717,N_49485);
and UO_1322 (O_1322,N_49982,N_49128);
xnor UO_1323 (O_1323,N_49493,N_49924);
and UO_1324 (O_1324,N_48779,N_48471);
and UO_1325 (O_1325,N_49107,N_48265);
and UO_1326 (O_1326,N_49750,N_48845);
xnor UO_1327 (O_1327,N_49515,N_48007);
and UO_1328 (O_1328,N_48135,N_49307);
or UO_1329 (O_1329,N_48458,N_48317);
and UO_1330 (O_1330,N_49894,N_48153);
nor UO_1331 (O_1331,N_49163,N_49629);
xnor UO_1332 (O_1332,N_48582,N_48475);
xor UO_1333 (O_1333,N_48737,N_49697);
and UO_1334 (O_1334,N_49028,N_48807);
or UO_1335 (O_1335,N_48808,N_49650);
nor UO_1336 (O_1336,N_48542,N_48457);
nand UO_1337 (O_1337,N_48449,N_48877);
nor UO_1338 (O_1338,N_48597,N_49301);
nand UO_1339 (O_1339,N_48922,N_48988);
nand UO_1340 (O_1340,N_49583,N_49543);
xor UO_1341 (O_1341,N_49147,N_48224);
nor UO_1342 (O_1342,N_48755,N_48200);
nor UO_1343 (O_1343,N_48058,N_49924);
and UO_1344 (O_1344,N_49247,N_48628);
xnor UO_1345 (O_1345,N_48493,N_49519);
and UO_1346 (O_1346,N_49405,N_48450);
or UO_1347 (O_1347,N_48960,N_49820);
nor UO_1348 (O_1348,N_48314,N_49304);
or UO_1349 (O_1349,N_49822,N_49399);
or UO_1350 (O_1350,N_49725,N_48900);
nor UO_1351 (O_1351,N_48409,N_48359);
nor UO_1352 (O_1352,N_49552,N_49092);
xnor UO_1353 (O_1353,N_48254,N_48350);
and UO_1354 (O_1354,N_48152,N_49744);
nand UO_1355 (O_1355,N_49322,N_49495);
xor UO_1356 (O_1356,N_49479,N_49770);
nand UO_1357 (O_1357,N_48439,N_49255);
nand UO_1358 (O_1358,N_49308,N_48664);
nand UO_1359 (O_1359,N_48531,N_48158);
nand UO_1360 (O_1360,N_48061,N_48119);
or UO_1361 (O_1361,N_49086,N_49750);
xor UO_1362 (O_1362,N_49690,N_48488);
nor UO_1363 (O_1363,N_49637,N_48018);
xnor UO_1364 (O_1364,N_48134,N_48529);
nor UO_1365 (O_1365,N_48640,N_49539);
nand UO_1366 (O_1366,N_48465,N_49784);
xnor UO_1367 (O_1367,N_48091,N_48367);
nand UO_1368 (O_1368,N_48319,N_49365);
xnor UO_1369 (O_1369,N_48302,N_48446);
and UO_1370 (O_1370,N_48633,N_49847);
or UO_1371 (O_1371,N_49470,N_49077);
and UO_1372 (O_1372,N_49741,N_49055);
and UO_1373 (O_1373,N_48927,N_48097);
nor UO_1374 (O_1374,N_49787,N_49183);
or UO_1375 (O_1375,N_49627,N_49737);
nand UO_1376 (O_1376,N_49777,N_48706);
nand UO_1377 (O_1377,N_48941,N_48538);
or UO_1378 (O_1378,N_48493,N_48302);
or UO_1379 (O_1379,N_49499,N_48599);
nor UO_1380 (O_1380,N_48299,N_48541);
or UO_1381 (O_1381,N_48379,N_48853);
nor UO_1382 (O_1382,N_49848,N_49796);
nand UO_1383 (O_1383,N_48956,N_49592);
xnor UO_1384 (O_1384,N_48714,N_49280);
xnor UO_1385 (O_1385,N_49101,N_49713);
xnor UO_1386 (O_1386,N_49830,N_49078);
nor UO_1387 (O_1387,N_49683,N_49305);
nor UO_1388 (O_1388,N_48021,N_48581);
and UO_1389 (O_1389,N_49072,N_48997);
xnor UO_1390 (O_1390,N_49213,N_48111);
xnor UO_1391 (O_1391,N_49323,N_48489);
nor UO_1392 (O_1392,N_48630,N_48215);
and UO_1393 (O_1393,N_49663,N_48498);
and UO_1394 (O_1394,N_48272,N_49466);
nand UO_1395 (O_1395,N_48831,N_48303);
nor UO_1396 (O_1396,N_48184,N_48394);
or UO_1397 (O_1397,N_49335,N_48682);
nor UO_1398 (O_1398,N_49353,N_49747);
nor UO_1399 (O_1399,N_49675,N_48824);
and UO_1400 (O_1400,N_49843,N_49055);
and UO_1401 (O_1401,N_48882,N_48486);
or UO_1402 (O_1402,N_49108,N_49283);
xor UO_1403 (O_1403,N_48236,N_48558);
and UO_1404 (O_1404,N_49352,N_49026);
xor UO_1405 (O_1405,N_48879,N_49326);
nand UO_1406 (O_1406,N_49171,N_49867);
and UO_1407 (O_1407,N_49674,N_49638);
and UO_1408 (O_1408,N_48016,N_48987);
or UO_1409 (O_1409,N_48431,N_49575);
or UO_1410 (O_1410,N_48979,N_49628);
and UO_1411 (O_1411,N_48295,N_48258);
xor UO_1412 (O_1412,N_49127,N_48759);
and UO_1413 (O_1413,N_48987,N_49866);
xnor UO_1414 (O_1414,N_49384,N_48578);
and UO_1415 (O_1415,N_49260,N_49244);
or UO_1416 (O_1416,N_48696,N_49043);
nand UO_1417 (O_1417,N_48962,N_49121);
xnor UO_1418 (O_1418,N_48678,N_49537);
nand UO_1419 (O_1419,N_49727,N_48856);
or UO_1420 (O_1420,N_48218,N_49259);
or UO_1421 (O_1421,N_49640,N_48943);
or UO_1422 (O_1422,N_48931,N_48046);
nand UO_1423 (O_1423,N_48560,N_49881);
and UO_1424 (O_1424,N_49679,N_49575);
xnor UO_1425 (O_1425,N_49041,N_48022);
nor UO_1426 (O_1426,N_49948,N_49493);
nor UO_1427 (O_1427,N_49765,N_48471);
or UO_1428 (O_1428,N_49741,N_48575);
nand UO_1429 (O_1429,N_49109,N_48848);
nor UO_1430 (O_1430,N_48265,N_48353);
nand UO_1431 (O_1431,N_49673,N_48640);
nor UO_1432 (O_1432,N_49183,N_49594);
or UO_1433 (O_1433,N_48127,N_49070);
nor UO_1434 (O_1434,N_48632,N_49152);
or UO_1435 (O_1435,N_48618,N_49618);
or UO_1436 (O_1436,N_48674,N_48480);
xnor UO_1437 (O_1437,N_49642,N_48492);
nand UO_1438 (O_1438,N_48106,N_48467);
or UO_1439 (O_1439,N_49408,N_49389);
nor UO_1440 (O_1440,N_49806,N_48865);
nor UO_1441 (O_1441,N_49759,N_49077);
nand UO_1442 (O_1442,N_49608,N_48944);
nor UO_1443 (O_1443,N_48427,N_48057);
nor UO_1444 (O_1444,N_49910,N_49960);
xor UO_1445 (O_1445,N_49673,N_49361);
and UO_1446 (O_1446,N_49719,N_49641);
xor UO_1447 (O_1447,N_49928,N_48999);
and UO_1448 (O_1448,N_49568,N_49990);
nor UO_1449 (O_1449,N_48513,N_48782);
xor UO_1450 (O_1450,N_49139,N_48801);
nor UO_1451 (O_1451,N_48241,N_49274);
and UO_1452 (O_1452,N_48015,N_49456);
or UO_1453 (O_1453,N_48286,N_49677);
or UO_1454 (O_1454,N_48124,N_48100);
nor UO_1455 (O_1455,N_48370,N_49574);
xnor UO_1456 (O_1456,N_49362,N_49596);
and UO_1457 (O_1457,N_48490,N_49989);
nand UO_1458 (O_1458,N_48094,N_48406);
xnor UO_1459 (O_1459,N_49119,N_49843);
and UO_1460 (O_1460,N_48918,N_49190);
or UO_1461 (O_1461,N_48250,N_48090);
or UO_1462 (O_1462,N_49532,N_48230);
and UO_1463 (O_1463,N_48838,N_48871);
nand UO_1464 (O_1464,N_49754,N_49849);
xor UO_1465 (O_1465,N_49765,N_49965);
nor UO_1466 (O_1466,N_49820,N_49692);
and UO_1467 (O_1467,N_48362,N_48806);
and UO_1468 (O_1468,N_48710,N_49087);
and UO_1469 (O_1469,N_49367,N_48375);
and UO_1470 (O_1470,N_48180,N_49772);
or UO_1471 (O_1471,N_49711,N_48637);
or UO_1472 (O_1472,N_49087,N_49584);
and UO_1473 (O_1473,N_48430,N_49578);
nor UO_1474 (O_1474,N_49367,N_48507);
and UO_1475 (O_1475,N_48730,N_49449);
nor UO_1476 (O_1476,N_48958,N_49670);
nor UO_1477 (O_1477,N_48679,N_49968);
nand UO_1478 (O_1478,N_48767,N_49060);
xnor UO_1479 (O_1479,N_49226,N_49107);
xor UO_1480 (O_1480,N_48804,N_49706);
nor UO_1481 (O_1481,N_48104,N_49843);
or UO_1482 (O_1482,N_48206,N_49631);
and UO_1483 (O_1483,N_49107,N_48833);
or UO_1484 (O_1484,N_49480,N_49146);
nand UO_1485 (O_1485,N_48387,N_49107);
nand UO_1486 (O_1486,N_49147,N_49588);
nor UO_1487 (O_1487,N_49761,N_49047);
xor UO_1488 (O_1488,N_48411,N_48739);
nand UO_1489 (O_1489,N_49409,N_48780);
nor UO_1490 (O_1490,N_49449,N_49431);
or UO_1491 (O_1491,N_48890,N_49987);
and UO_1492 (O_1492,N_49125,N_48384);
nand UO_1493 (O_1493,N_49824,N_48932);
nand UO_1494 (O_1494,N_49934,N_49899);
nor UO_1495 (O_1495,N_48881,N_49942);
or UO_1496 (O_1496,N_48826,N_48926);
nand UO_1497 (O_1497,N_48232,N_49848);
xor UO_1498 (O_1498,N_49895,N_49561);
and UO_1499 (O_1499,N_48449,N_49858);
and UO_1500 (O_1500,N_48491,N_48321);
nor UO_1501 (O_1501,N_49233,N_49264);
nand UO_1502 (O_1502,N_48137,N_48906);
nor UO_1503 (O_1503,N_49837,N_49308);
and UO_1504 (O_1504,N_49459,N_48629);
nor UO_1505 (O_1505,N_49486,N_48388);
nor UO_1506 (O_1506,N_48947,N_49430);
and UO_1507 (O_1507,N_49303,N_48684);
nor UO_1508 (O_1508,N_49175,N_48040);
and UO_1509 (O_1509,N_48898,N_49610);
and UO_1510 (O_1510,N_48039,N_48882);
nand UO_1511 (O_1511,N_48168,N_49688);
nor UO_1512 (O_1512,N_49172,N_48928);
xnor UO_1513 (O_1513,N_48953,N_49899);
and UO_1514 (O_1514,N_49287,N_49470);
xnor UO_1515 (O_1515,N_49684,N_48157);
or UO_1516 (O_1516,N_48357,N_48988);
or UO_1517 (O_1517,N_49138,N_48917);
or UO_1518 (O_1518,N_48951,N_48408);
and UO_1519 (O_1519,N_49603,N_48820);
or UO_1520 (O_1520,N_48413,N_49868);
nor UO_1521 (O_1521,N_48082,N_49709);
nor UO_1522 (O_1522,N_49755,N_49588);
or UO_1523 (O_1523,N_49913,N_49476);
nor UO_1524 (O_1524,N_49191,N_49755);
nor UO_1525 (O_1525,N_49161,N_49656);
and UO_1526 (O_1526,N_49906,N_49593);
xnor UO_1527 (O_1527,N_48477,N_48677);
nand UO_1528 (O_1528,N_49947,N_48310);
or UO_1529 (O_1529,N_49840,N_49749);
or UO_1530 (O_1530,N_49156,N_48268);
or UO_1531 (O_1531,N_48838,N_48178);
nor UO_1532 (O_1532,N_49858,N_49871);
and UO_1533 (O_1533,N_48166,N_49885);
nor UO_1534 (O_1534,N_49710,N_48945);
nand UO_1535 (O_1535,N_48881,N_49794);
xor UO_1536 (O_1536,N_49142,N_49417);
nor UO_1537 (O_1537,N_48374,N_49771);
and UO_1538 (O_1538,N_49748,N_49104);
nor UO_1539 (O_1539,N_49534,N_48330);
and UO_1540 (O_1540,N_48344,N_49077);
and UO_1541 (O_1541,N_48741,N_48071);
and UO_1542 (O_1542,N_48574,N_48895);
nor UO_1543 (O_1543,N_49588,N_48860);
or UO_1544 (O_1544,N_49962,N_49888);
xnor UO_1545 (O_1545,N_49790,N_49448);
nor UO_1546 (O_1546,N_48732,N_49889);
and UO_1547 (O_1547,N_49155,N_48156);
and UO_1548 (O_1548,N_48824,N_48112);
and UO_1549 (O_1549,N_48139,N_49814);
and UO_1550 (O_1550,N_48430,N_49532);
and UO_1551 (O_1551,N_49653,N_48242);
or UO_1552 (O_1552,N_49767,N_48334);
nand UO_1553 (O_1553,N_48743,N_49335);
nor UO_1554 (O_1554,N_49571,N_48596);
or UO_1555 (O_1555,N_49927,N_48740);
or UO_1556 (O_1556,N_48948,N_49968);
or UO_1557 (O_1557,N_48101,N_48306);
xor UO_1558 (O_1558,N_49193,N_48902);
nand UO_1559 (O_1559,N_48027,N_49477);
and UO_1560 (O_1560,N_49135,N_49652);
and UO_1561 (O_1561,N_48832,N_48490);
nand UO_1562 (O_1562,N_48107,N_49041);
xor UO_1563 (O_1563,N_48174,N_49019);
or UO_1564 (O_1564,N_48067,N_48356);
and UO_1565 (O_1565,N_48778,N_49682);
nor UO_1566 (O_1566,N_48803,N_49538);
nor UO_1567 (O_1567,N_48332,N_49691);
xor UO_1568 (O_1568,N_49474,N_48638);
nand UO_1569 (O_1569,N_49573,N_48153);
nor UO_1570 (O_1570,N_49619,N_48674);
and UO_1571 (O_1571,N_49537,N_49674);
or UO_1572 (O_1572,N_49884,N_49008);
nand UO_1573 (O_1573,N_48781,N_48943);
nand UO_1574 (O_1574,N_48576,N_49363);
xor UO_1575 (O_1575,N_49123,N_48457);
xor UO_1576 (O_1576,N_48229,N_49184);
nor UO_1577 (O_1577,N_48002,N_49440);
or UO_1578 (O_1578,N_48833,N_48890);
or UO_1579 (O_1579,N_48825,N_48347);
xor UO_1580 (O_1580,N_49728,N_48707);
or UO_1581 (O_1581,N_49739,N_48282);
nor UO_1582 (O_1582,N_48842,N_49230);
xor UO_1583 (O_1583,N_49286,N_49906);
or UO_1584 (O_1584,N_48050,N_49049);
nand UO_1585 (O_1585,N_49922,N_48779);
and UO_1586 (O_1586,N_49646,N_49503);
xnor UO_1587 (O_1587,N_49040,N_49041);
or UO_1588 (O_1588,N_48535,N_48086);
nor UO_1589 (O_1589,N_48179,N_48244);
or UO_1590 (O_1590,N_49241,N_49056);
and UO_1591 (O_1591,N_49046,N_48098);
or UO_1592 (O_1592,N_49842,N_49313);
and UO_1593 (O_1593,N_48576,N_49376);
xnor UO_1594 (O_1594,N_49307,N_48501);
nand UO_1595 (O_1595,N_49781,N_48208);
xnor UO_1596 (O_1596,N_48723,N_48925);
xor UO_1597 (O_1597,N_49259,N_48767);
or UO_1598 (O_1598,N_48907,N_48776);
xor UO_1599 (O_1599,N_48019,N_48993);
nor UO_1600 (O_1600,N_48345,N_48813);
xnor UO_1601 (O_1601,N_49066,N_49235);
nor UO_1602 (O_1602,N_49348,N_48790);
xor UO_1603 (O_1603,N_48625,N_48531);
or UO_1604 (O_1604,N_48883,N_49456);
and UO_1605 (O_1605,N_48132,N_48547);
xnor UO_1606 (O_1606,N_48598,N_49475);
nand UO_1607 (O_1607,N_48521,N_49880);
nor UO_1608 (O_1608,N_48839,N_48164);
and UO_1609 (O_1609,N_48853,N_49092);
xor UO_1610 (O_1610,N_49444,N_49834);
and UO_1611 (O_1611,N_48152,N_49862);
or UO_1612 (O_1612,N_48506,N_49266);
or UO_1613 (O_1613,N_49316,N_49072);
xor UO_1614 (O_1614,N_48166,N_49248);
nand UO_1615 (O_1615,N_49113,N_49032);
nand UO_1616 (O_1616,N_48462,N_48565);
or UO_1617 (O_1617,N_48071,N_48223);
nand UO_1618 (O_1618,N_48898,N_49457);
nand UO_1619 (O_1619,N_49795,N_49114);
nand UO_1620 (O_1620,N_48074,N_48000);
nor UO_1621 (O_1621,N_49648,N_48615);
or UO_1622 (O_1622,N_48381,N_48027);
xor UO_1623 (O_1623,N_48508,N_48595);
and UO_1624 (O_1624,N_48434,N_48374);
or UO_1625 (O_1625,N_49103,N_48343);
nor UO_1626 (O_1626,N_49711,N_48363);
nor UO_1627 (O_1627,N_49826,N_48269);
xor UO_1628 (O_1628,N_49845,N_49288);
and UO_1629 (O_1629,N_48358,N_49141);
or UO_1630 (O_1630,N_49638,N_49274);
nand UO_1631 (O_1631,N_48719,N_48683);
xnor UO_1632 (O_1632,N_49804,N_49026);
xnor UO_1633 (O_1633,N_48382,N_48551);
nand UO_1634 (O_1634,N_48014,N_49680);
nand UO_1635 (O_1635,N_48181,N_49383);
and UO_1636 (O_1636,N_48214,N_48253);
and UO_1637 (O_1637,N_48829,N_49303);
nor UO_1638 (O_1638,N_48956,N_49288);
xor UO_1639 (O_1639,N_48138,N_49062);
or UO_1640 (O_1640,N_48246,N_48830);
xor UO_1641 (O_1641,N_48754,N_49021);
or UO_1642 (O_1642,N_49160,N_48151);
xor UO_1643 (O_1643,N_49209,N_49450);
or UO_1644 (O_1644,N_48435,N_48540);
and UO_1645 (O_1645,N_48624,N_48348);
xnor UO_1646 (O_1646,N_48397,N_48736);
or UO_1647 (O_1647,N_49050,N_48941);
nand UO_1648 (O_1648,N_49855,N_48349);
and UO_1649 (O_1649,N_49478,N_48111);
xnor UO_1650 (O_1650,N_49640,N_49270);
xor UO_1651 (O_1651,N_49045,N_48225);
xnor UO_1652 (O_1652,N_48773,N_49226);
xnor UO_1653 (O_1653,N_48932,N_48255);
xnor UO_1654 (O_1654,N_48957,N_48753);
xnor UO_1655 (O_1655,N_48692,N_49280);
nand UO_1656 (O_1656,N_49975,N_49482);
nand UO_1657 (O_1657,N_48991,N_49266);
nor UO_1658 (O_1658,N_48566,N_48105);
or UO_1659 (O_1659,N_48741,N_48713);
and UO_1660 (O_1660,N_49183,N_49341);
nand UO_1661 (O_1661,N_49065,N_49651);
nand UO_1662 (O_1662,N_48239,N_48541);
nand UO_1663 (O_1663,N_48157,N_49739);
or UO_1664 (O_1664,N_49691,N_48451);
nand UO_1665 (O_1665,N_48796,N_48036);
nand UO_1666 (O_1666,N_49889,N_49245);
nor UO_1667 (O_1667,N_48247,N_48372);
or UO_1668 (O_1668,N_49542,N_48380);
nor UO_1669 (O_1669,N_49426,N_49455);
nand UO_1670 (O_1670,N_48525,N_49848);
nand UO_1671 (O_1671,N_49038,N_49631);
and UO_1672 (O_1672,N_49355,N_49898);
and UO_1673 (O_1673,N_48375,N_49775);
nand UO_1674 (O_1674,N_48169,N_49656);
and UO_1675 (O_1675,N_49445,N_48463);
xnor UO_1676 (O_1676,N_48843,N_49814);
and UO_1677 (O_1677,N_48142,N_49176);
or UO_1678 (O_1678,N_49074,N_48157);
or UO_1679 (O_1679,N_49002,N_48812);
nor UO_1680 (O_1680,N_49115,N_49056);
nor UO_1681 (O_1681,N_48201,N_49354);
or UO_1682 (O_1682,N_49355,N_49141);
or UO_1683 (O_1683,N_49417,N_49357);
xnor UO_1684 (O_1684,N_48411,N_48003);
and UO_1685 (O_1685,N_49906,N_48440);
or UO_1686 (O_1686,N_49943,N_48748);
nor UO_1687 (O_1687,N_49076,N_48645);
xnor UO_1688 (O_1688,N_48473,N_49171);
and UO_1689 (O_1689,N_48858,N_48357);
nor UO_1690 (O_1690,N_48030,N_48448);
and UO_1691 (O_1691,N_48613,N_49161);
nor UO_1692 (O_1692,N_49789,N_48079);
nor UO_1693 (O_1693,N_48177,N_48499);
and UO_1694 (O_1694,N_48348,N_49541);
or UO_1695 (O_1695,N_48550,N_49215);
nor UO_1696 (O_1696,N_48484,N_48117);
nor UO_1697 (O_1697,N_49152,N_49394);
nand UO_1698 (O_1698,N_49264,N_49716);
xor UO_1699 (O_1699,N_48839,N_49818);
or UO_1700 (O_1700,N_48880,N_48916);
or UO_1701 (O_1701,N_49929,N_48726);
xor UO_1702 (O_1702,N_49747,N_48613);
or UO_1703 (O_1703,N_48681,N_48014);
nand UO_1704 (O_1704,N_49038,N_48488);
xnor UO_1705 (O_1705,N_49305,N_49026);
nor UO_1706 (O_1706,N_48135,N_48924);
nand UO_1707 (O_1707,N_49711,N_49141);
nand UO_1708 (O_1708,N_49965,N_49102);
nor UO_1709 (O_1709,N_49917,N_48808);
and UO_1710 (O_1710,N_49988,N_48490);
nand UO_1711 (O_1711,N_49616,N_48480);
nor UO_1712 (O_1712,N_49064,N_48526);
and UO_1713 (O_1713,N_48399,N_49974);
or UO_1714 (O_1714,N_48382,N_49729);
nor UO_1715 (O_1715,N_49368,N_49671);
or UO_1716 (O_1716,N_48635,N_48923);
xor UO_1717 (O_1717,N_49860,N_49106);
nand UO_1718 (O_1718,N_48495,N_48003);
nor UO_1719 (O_1719,N_49462,N_49461);
xor UO_1720 (O_1720,N_48667,N_49872);
and UO_1721 (O_1721,N_49322,N_49005);
and UO_1722 (O_1722,N_48082,N_48596);
xor UO_1723 (O_1723,N_49442,N_49620);
xor UO_1724 (O_1724,N_48629,N_49402);
nand UO_1725 (O_1725,N_49592,N_48152);
nor UO_1726 (O_1726,N_48159,N_48323);
nand UO_1727 (O_1727,N_49972,N_49488);
nand UO_1728 (O_1728,N_48951,N_49502);
nand UO_1729 (O_1729,N_48302,N_48325);
xnor UO_1730 (O_1730,N_48888,N_49148);
xor UO_1731 (O_1731,N_49020,N_49759);
or UO_1732 (O_1732,N_49463,N_48044);
or UO_1733 (O_1733,N_48689,N_49577);
or UO_1734 (O_1734,N_48969,N_48987);
xor UO_1735 (O_1735,N_48240,N_48196);
nor UO_1736 (O_1736,N_49757,N_48570);
xnor UO_1737 (O_1737,N_48026,N_49220);
and UO_1738 (O_1738,N_49760,N_48756);
or UO_1739 (O_1739,N_48126,N_49306);
xor UO_1740 (O_1740,N_49072,N_48258);
or UO_1741 (O_1741,N_49781,N_48233);
xnor UO_1742 (O_1742,N_49409,N_48153);
and UO_1743 (O_1743,N_49713,N_48255);
nor UO_1744 (O_1744,N_48545,N_48443);
nand UO_1745 (O_1745,N_48651,N_49772);
or UO_1746 (O_1746,N_48474,N_48388);
and UO_1747 (O_1747,N_49318,N_48524);
or UO_1748 (O_1748,N_48224,N_49075);
or UO_1749 (O_1749,N_48282,N_49953);
or UO_1750 (O_1750,N_49325,N_48845);
and UO_1751 (O_1751,N_48608,N_49721);
and UO_1752 (O_1752,N_48600,N_48359);
nand UO_1753 (O_1753,N_48191,N_48330);
or UO_1754 (O_1754,N_49369,N_49344);
nand UO_1755 (O_1755,N_48306,N_49407);
xor UO_1756 (O_1756,N_49522,N_49663);
or UO_1757 (O_1757,N_48414,N_49824);
nand UO_1758 (O_1758,N_49111,N_48855);
nor UO_1759 (O_1759,N_49628,N_48119);
nand UO_1760 (O_1760,N_48907,N_49108);
nand UO_1761 (O_1761,N_48251,N_48667);
xnor UO_1762 (O_1762,N_49606,N_48911);
and UO_1763 (O_1763,N_48190,N_49728);
or UO_1764 (O_1764,N_48286,N_48949);
xnor UO_1765 (O_1765,N_48974,N_49966);
nor UO_1766 (O_1766,N_49317,N_49458);
and UO_1767 (O_1767,N_49779,N_49772);
and UO_1768 (O_1768,N_48170,N_49005);
or UO_1769 (O_1769,N_49534,N_49553);
nand UO_1770 (O_1770,N_49253,N_49163);
or UO_1771 (O_1771,N_48793,N_49948);
xor UO_1772 (O_1772,N_48031,N_49313);
xor UO_1773 (O_1773,N_48392,N_48972);
xor UO_1774 (O_1774,N_48385,N_48229);
xor UO_1775 (O_1775,N_49071,N_48243);
nand UO_1776 (O_1776,N_48759,N_49167);
or UO_1777 (O_1777,N_48804,N_48508);
nand UO_1778 (O_1778,N_48016,N_49549);
nand UO_1779 (O_1779,N_48206,N_48857);
nand UO_1780 (O_1780,N_48082,N_49519);
or UO_1781 (O_1781,N_48356,N_48415);
nor UO_1782 (O_1782,N_48785,N_48603);
nor UO_1783 (O_1783,N_48159,N_49932);
nand UO_1784 (O_1784,N_49644,N_48003);
nor UO_1785 (O_1785,N_49616,N_49041);
and UO_1786 (O_1786,N_49834,N_49179);
and UO_1787 (O_1787,N_49236,N_49010);
nand UO_1788 (O_1788,N_49149,N_49105);
and UO_1789 (O_1789,N_48180,N_48368);
or UO_1790 (O_1790,N_49498,N_48364);
and UO_1791 (O_1791,N_48626,N_49752);
nand UO_1792 (O_1792,N_49169,N_49143);
nor UO_1793 (O_1793,N_49102,N_48898);
and UO_1794 (O_1794,N_49017,N_49290);
and UO_1795 (O_1795,N_48210,N_49464);
nand UO_1796 (O_1796,N_49625,N_49502);
or UO_1797 (O_1797,N_49245,N_49165);
nand UO_1798 (O_1798,N_49642,N_49954);
xor UO_1799 (O_1799,N_48436,N_49009);
nand UO_1800 (O_1800,N_49944,N_48472);
nand UO_1801 (O_1801,N_49388,N_48706);
nor UO_1802 (O_1802,N_49730,N_49695);
nand UO_1803 (O_1803,N_49094,N_48573);
nand UO_1804 (O_1804,N_49532,N_48562);
xor UO_1805 (O_1805,N_48916,N_49492);
nor UO_1806 (O_1806,N_49866,N_48747);
and UO_1807 (O_1807,N_49315,N_48861);
and UO_1808 (O_1808,N_49038,N_48305);
and UO_1809 (O_1809,N_48706,N_49243);
xnor UO_1810 (O_1810,N_49519,N_49840);
and UO_1811 (O_1811,N_49678,N_48223);
nor UO_1812 (O_1812,N_49778,N_48292);
nand UO_1813 (O_1813,N_48260,N_48118);
and UO_1814 (O_1814,N_49374,N_48013);
nand UO_1815 (O_1815,N_49365,N_48943);
xor UO_1816 (O_1816,N_49462,N_49976);
nor UO_1817 (O_1817,N_49443,N_49634);
xnor UO_1818 (O_1818,N_48818,N_49727);
nor UO_1819 (O_1819,N_49341,N_48381);
nand UO_1820 (O_1820,N_48737,N_49616);
nand UO_1821 (O_1821,N_48097,N_49811);
xnor UO_1822 (O_1822,N_49478,N_48026);
and UO_1823 (O_1823,N_48800,N_49062);
and UO_1824 (O_1824,N_48364,N_49447);
xnor UO_1825 (O_1825,N_48388,N_49959);
xor UO_1826 (O_1826,N_48576,N_48496);
and UO_1827 (O_1827,N_48077,N_48671);
xor UO_1828 (O_1828,N_49787,N_49936);
xor UO_1829 (O_1829,N_48147,N_48096);
or UO_1830 (O_1830,N_49309,N_48009);
and UO_1831 (O_1831,N_48269,N_49835);
or UO_1832 (O_1832,N_48612,N_49225);
and UO_1833 (O_1833,N_49909,N_48923);
and UO_1834 (O_1834,N_49150,N_48747);
xnor UO_1835 (O_1835,N_49535,N_49645);
xor UO_1836 (O_1836,N_48668,N_49866);
or UO_1837 (O_1837,N_48803,N_48022);
nor UO_1838 (O_1838,N_48094,N_49564);
and UO_1839 (O_1839,N_48062,N_49768);
and UO_1840 (O_1840,N_48412,N_49444);
and UO_1841 (O_1841,N_49359,N_49997);
and UO_1842 (O_1842,N_48474,N_49892);
nor UO_1843 (O_1843,N_49444,N_48741);
and UO_1844 (O_1844,N_49337,N_49370);
nor UO_1845 (O_1845,N_48984,N_49463);
and UO_1846 (O_1846,N_48041,N_49005);
xor UO_1847 (O_1847,N_48471,N_49502);
and UO_1848 (O_1848,N_48028,N_48722);
and UO_1849 (O_1849,N_49436,N_48966);
or UO_1850 (O_1850,N_49639,N_49610);
or UO_1851 (O_1851,N_48507,N_49189);
nor UO_1852 (O_1852,N_48737,N_48160);
and UO_1853 (O_1853,N_49494,N_49737);
or UO_1854 (O_1854,N_49623,N_49848);
xor UO_1855 (O_1855,N_49811,N_48517);
nor UO_1856 (O_1856,N_48117,N_49057);
nand UO_1857 (O_1857,N_49900,N_49263);
or UO_1858 (O_1858,N_48776,N_48259);
or UO_1859 (O_1859,N_49142,N_48479);
nor UO_1860 (O_1860,N_48971,N_49857);
nor UO_1861 (O_1861,N_48545,N_48318);
xnor UO_1862 (O_1862,N_49918,N_48456);
nand UO_1863 (O_1863,N_48257,N_49738);
and UO_1864 (O_1864,N_49772,N_49143);
xnor UO_1865 (O_1865,N_48532,N_49311);
nor UO_1866 (O_1866,N_49661,N_49699);
nor UO_1867 (O_1867,N_49801,N_49837);
nand UO_1868 (O_1868,N_48311,N_48864);
nor UO_1869 (O_1869,N_49652,N_49326);
nor UO_1870 (O_1870,N_48431,N_48473);
xor UO_1871 (O_1871,N_49754,N_48656);
nor UO_1872 (O_1872,N_48584,N_48630);
nand UO_1873 (O_1873,N_49279,N_49752);
or UO_1874 (O_1874,N_48771,N_49038);
nand UO_1875 (O_1875,N_49321,N_49362);
and UO_1876 (O_1876,N_49399,N_48472);
xor UO_1877 (O_1877,N_48661,N_48390);
nand UO_1878 (O_1878,N_48375,N_49769);
nand UO_1879 (O_1879,N_48042,N_49500);
nand UO_1880 (O_1880,N_49446,N_49032);
nand UO_1881 (O_1881,N_49471,N_49881);
and UO_1882 (O_1882,N_48060,N_48158);
nor UO_1883 (O_1883,N_49908,N_48273);
xor UO_1884 (O_1884,N_48408,N_49739);
and UO_1885 (O_1885,N_49809,N_48018);
nor UO_1886 (O_1886,N_48447,N_48042);
nand UO_1887 (O_1887,N_49821,N_49323);
or UO_1888 (O_1888,N_48808,N_49453);
nand UO_1889 (O_1889,N_48850,N_49673);
nand UO_1890 (O_1890,N_48293,N_49074);
or UO_1891 (O_1891,N_49827,N_49688);
nand UO_1892 (O_1892,N_48723,N_49106);
xnor UO_1893 (O_1893,N_48282,N_49872);
nand UO_1894 (O_1894,N_48386,N_49661);
nand UO_1895 (O_1895,N_49805,N_48781);
nand UO_1896 (O_1896,N_48786,N_48839);
or UO_1897 (O_1897,N_48143,N_48434);
and UO_1898 (O_1898,N_48395,N_48134);
and UO_1899 (O_1899,N_49783,N_48536);
nor UO_1900 (O_1900,N_49251,N_48159);
and UO_1901 (O_1901,N_49199,N_48799);
or UO_1902 (O_1902,N_48544,N_49375);
and UO_1903 (O_1903,N_48254,N_48742);
and UO_1904 (O_1904,N_49398,N_48234);
xnor UO_1905 (O_1905,N_48466,N_49741);
and UO_1906 (O_1906,N_48382,N_48073);
xor UO_1907 (O_1907,N_49812,N_48803);
nand UO_1908 (O_1908,N_49129,N_49116);
nand UO_1909 (O_1909,N_49952,N_49493);
or UO_1910 (O_1910,N_49540,N_48380);
or UO_1911 (O_1911,N_49811,N_48554);
xnor UO_1912 (O_1912,N_48740,N_49631);
nand UO_1913 (O_1913,N_49701,N_49151);
nor UO_1914 (O_1914,N_49115,N_48640);
nor UO_1915 (O_1915,N_49377,N_49170);
nand UO_1916 (O_1916,N_48251,N_48185);
nand UO_1917 (O_1917,N_49239,N_48636);
or UO_1918 (O_1918,N_49867,N_48561);
or UO_1919 (O_1919,N_49237,N_49705);
or UO_1920 (O_1920,N_49497,N_49812);
or UO_1921 (O_1921,N_49574,N_48133);
nand UO_1922 (O_1922,N_48637,N_48693);
nor UO_1923 (O_1923,N_49239,N_49624);
or UO_1924 (O_1924,N_48877,N_48735);
xor UO_1925 (O_1925,N_48607,N_49056);
xnor UO_1926 (O_1926,N_49731,N_48793);
xnor UO_1927 (O_1927,N_48908,N_48246);
nand UO_1928 (O_1928,N_48407,N_49433);
or UO_1929 (O_1929,N_48993,N_49764);
xor UO_1930 (O_1930,N_49664,N_49193);
xor UO_1931 (O_1931,N_48662,N_49358);
or UO_1932 (O_1932,N_49216,N_49505);
or UO_1933 (O_1933,N_49079,N_49922);
and UO_1934 (O_1934,N_48691,N_49354);
and UO_1935 (O_1935,N_49229,N_48480);
nor UO_1936 (O_1936,N_48782,N_49019);
xnor UO_1937 (O_1937,N_48260,N_49441);
nor UO_1938 (O_1938,N_49725,N_49040);
or UO_1939 (O_1939,N_49683,N_49969);
nor UO_1940 (O_1940,N_48607,N_49019);
xor UO_1941 (O_1941,N_49365,N_49171);
nand UO_1942 (O_1942,N_49541,N_49086);
or UO_1943 (O_1943,N_49672,N_49751);
nand UO_1944 (O_1944,N_49486,N_49412);
and UO_1945 (O_1945,N_49657,N_49354);
xor UO_1946 (O_1946,N_48345,N_49795);
or UO_1947 (O_1947,N_48807,N_48983);
or UO_1948 (O_1948,N_48046,N_48080);
xor UO_1949 (O_1949,N_48845,N_48958);
nor UO_1950 (O_1950,N_49033,N_49617);
nand UO_1951 (O_1951,N_48648,N_49059);
xnor UO_1952 (O_1952,N_48377,N_48280);
xnor UO_1953 (O_1953,N_49299,N_48465);
nand UO_1954 (O_1954,N_49756,N_48980);
and UO_1955 (O_1955,N_48898,N_49965);
and UO_1956 (O_1956,N_48300,N_49818);
nor UO_1957 (O_1957,N_49790,N_49310);
nand UO_1958 (O_1958,N_49476,N_48353);
xor UO_1959 (O_1959,N_49697,N_48131);
and UO_1960 (O_1960,N_48042,N_48004);
and UO_1961 (O_1961,N_48465,N_48422);
nand UO_1962 (O_1962,N_49594,N_49799);
xor UO_1963 (O_1963,N_48903,N_48516);
and UO_1964 (O_1964,N_49225,N_48087);
nor UO_1965 (O_1965,N_49579,N_48283);
and UO_1966 (O_1966,N_48132,N_49814);
nand UO_1967 (O_1967,N_49761,N_48952);
and UO_1968 (O_1968,N_49271,N_49712);
and UO_1969 (O_1969,N_48037,N_48878);
nand UO_1970 (O_1970,N_48656,N_49612);
nand UO_1971 (O_1971,N_49367,N_49894);
and UO_1972 (O_1972,N_48069,N_48417);
xnor UO_1973 (O_1973,N_48086,N_49859);
and UO_1974 (O_1974,N_48497,N_48841);
or UO_1975 (O_1975,N_49756,N_48158);
and UO_1976 (O_1976,N_48197,N_48861);
nor UO_1977 (O_1977,N_48789,N_48419);
nor UO_1978 (O_1978,N_48217,N_48440);
nand UO_1979 (O_1979,N_48137,N_49175);
and UO_1980 (O_1980,N_48298,N_48457);
nand UO_1981 (O_1981,N_48125,N_49020);
or UO_1982 (O_1982,N_48045,N_48334);
xnor UO_1983 (O_1983,N_49960,N_48908);
or UO_1984 (O_1984,N_48361,N_48307);
or UO_1985 (O_1985,N_48568,N_49138);
or UO_1986 (O_1986,N_49592,N_49015);
nor UO_1987 (O_1987,N_49206,N_48528);
or UO_1988 (O_1988,N_49723,N_49831);
nor UO_1989 (O_1989,N_48887,N_49665);
nand UO_1990 (O_1990,N_49047,N_48189);
and UO_1991 (O_1991,N_48845,N_48070);
xnor UO_1992 (O_1992,N_49493,N_49515);
or UO_1993 (O_1993,N_49919,N_49071);
or UO_1994 (O_1994,N_49917,N_48491);
nor UO_1995 (O_1995,N_48271,N_48507);
and UO_1996 (O_1996,N_48754,N_48566);
xor UO_1997 (O_1997,N_49433,N_48656);
or UO_1998 (O_1998,N_48107,N_49769);
nand UO_1999 (O_1999,N_49755,N_49678);
xnor UO_2000 (O_2000,N_49553,N_48972);
or UO_2001 (O_2001,N_48867,N_48514);
and UO_2002 (O_2002,N_49620,N_48488);
nand UO_2003 (O_2003,N_49060,N_49993);
nor UO_2004 (O_2004,N_48654,N_49032);
and UO_2005 (O_2005,N_48965,N_49234);
xnor UO_2006 (O_2006,N_49253,N_49329);
or UO_2007 (O_2007,N_49690,N_48980);
xor UO_2008 (O_2008,N_49223,N_49494);
or UO_2009 (O_2009,N_49112,N_49405);
nand UO_2010 (O_2010,N_49827,N_49655);
and UO_2011 (O_2011,N_48677,N_48300);
or UO_2012 (O_2012,N_48005,N_49647);
and UO_2013 (O_2013,N_48991,N_49745);
and UO_2014 (O_2014,N_49725,N_48785);
nor UO_2015 (O_2015,N_48158,N_48104);
and UO_2016 (O_2016,N_48224,N_49642);
nand UO_2017 (O_2017,N_49614,N_49160);
and UO_2018 (O_2018,N_48459,N_49170);
xnor UO_2019 (O_2019,N_48833,N_48756);
nor UO_2020 (O_2020,N_48848,N_48252);
nor UO_2021 (O_2021,N_48050,N_49567);
xnor UO_2022 (O_2022,N_49637,N_49648);
and UO_2023 (O_2023,N_48841,N_48577);
nor UO_2024 (O_2024,N_49176,N_48330);
or UO_2025 (O_2025,N_48540,N_48938);
nand UO_2026 (O_2026,N_49206,N_49791);
nand UO_2027 (O_2027,N_48807,N_49819);
nand UO_2028 (O_2028,N_49197,N_48368);
or UO_2029 (O_2029,N_49648,N_49357);
or UO_2030 (O_2030,N_48837,N_49991);
and UO_2031 (O_2031,N_48412,N_48386);
nand UO_2032 (O_2032,N_48007,N_48080);
nor UO_2033 (O_2033,N_49485,N_49278);
nand UO_2034 (O_2034,N_48808,N_48645);
nand UO_2035 (O_2035,N_49967,N_49408);
nor UO_2036 (O_2036,N_48566,N_49515);
or UO_2037 (O_2037,N_48632,N_49990);
or UO_2038 (O_2038,N_49045,N_48249);
nand UO_2039 (O_2039,N_49237,N_48272);
xnor UO_2040 (O_2040,N_49399,N_48984);
xor UO_2041 (O_2041,N_49238,N_49314);
and UO_2042 (O_2042,N_48932,N_49033);
or UO_2043 (O_2043,N_49601,N_48764);
nor UO_2044 (O_2044,N_49158,N_48502);
nand UO_2045 (O_2045,N_48029,N_49544);
nand UO_2046 (O_2046,N_49837,N_49104);
nand UO_2047 (O_2047,N_48852,N_49768);
xnor UO_2048 (O_2048,N_49146,N_49883);
or UO_2049 (O_2049,N_48060,N_48748);
nand UO_2050 (O_2050,N_49212,N_48151);
nand UO_2051 (O_2051,N_48611,N_49797);
nand UO_2052 (O_2052,N_49401,N_49170);
nand UO_2053 (O_2053,N_48393,N_49336);
or UO_2054 (O_2054,N_49907,N_48565);
nand UO_2055 (O_2055,N_49861,N_49147);
nand UO_2056 (O_2056,N_49115,N_49626);
xor UO_2057 (O_2057,N_49109,N_48766);
nand UO_2058 (O_2058,N_48101,N_48790);
nor UO_2059 (O_2059,N_48717,N_49421);
nand UO_2060 (O_2060,N_49206,N_48674);
nor UO_2061 (O_2061,N_48887,N_49356);
or UO_2062 (O_2062,N_49598,N_48952);
nand UO_2063 (O_2063,N_49604,N_49053);
xnor UO_2064 (O_2064,N_49218,N_48309);
nand UO_2065 (O_2065,N_48596,N_48709);
and UO_2066 (O_2066,N_48261,N_49310);
nor UO_2067 (O_2067,N_48520,N_48722);
nor UO_2068 (O_2068,N_48177,N_48504);
nand UO_2069 (O_2069,N_49175,N_49057);
nand UO_2070 (O_2070,N_48152,N_49059);
and UO_2071 (O_2071,N_48553,N_49411);
nor UO_2072 (O_2072,N_49336,N_49053);
xor UO_2073 (O_2073,N_49615,N_49223);
nor UO_2074 (O_2074,N_49488,N_48372);
xnor UO_2075 (O_2075,N_48299,N_48748);
or UO_2076 (O_2076,N_49548,N_48114);
nand UO_2077 (O_2077,N_49998,N_49262);
or UO_2078 (O_2078,N_49997,N_48536);
nand UO_2079 (O_2079,N_49610,N_48430);
nor UO_2080 (O_2080,N_49013,N_49393);
nand UO_2081 (O_2081,N_48677,N_48546);
nand UO_2082 (O_2082,N_49899,N_49160);
and UO_2083 (O_2083,N_48812,N_49435);
nand UO_2084 (O_2084,N_49330,N_48923);
xnor UO_2085 (O_2085,N_49256,N_49531);
or UO_2086 (O_2086,N_48143,N_49543);
or UO_2087 (O_2087,N_48523,N_49125);
nor UO_2088 (O_2088,N_48508,N_49525);
or UO_2089 (O_2089,N_49784,N_49524);
nor UO_2090 (O_2090,N_49046,N_48500);
nor UO_2091 (O_2091,N_49467,N_48266);
or UO_2092 (O_2092,N_48210,N_49211);
and UO_2093 (O_2093,N_49498,N_49127);
xor UO_2094 (O_2094,N_48965,N_49026);
nor UO_2095 (O_2095,N_48755,N_48177);
nand UO_2096 (O_2096,N_48221,N_48485);
xnor UO_2097 (O_2097,N_49688,N_49926);
or UO_2098 (O_2098,N_48232,N_48358);
and UO_2099 (O_2099,N_49606,N_49133);
xnor UO_2100 (O_2100,N_49007,N_49983);
nor UO_2101 (O_2101,N_49903,N_48888);
nand UO_2102 (O_2102,N_49654,N_48857);
nor UO_2103 (O_2103,N_49205,N_48348);
and UO_2104 (O_2104,N_48149,N_49974);
nor UO_2105 (O_2105,N_48914,N_49027);
xor UO_2106 (O_2106,N_48063,N_49557);
and UO_2107 (O_2107,N_48035,N_48612);
xnor UO_2108 (O_2108,N_48637,N_49470);
and UO_2109 (O_2109,N_49943,N_48739);
nand UO_2110 (O_2110,N_48161,N_48225);
or UO_2111 (O_2111,N_48316,N_48675);
and UO_2112 (O_2112,N_49242,N_48640);
nor UO_2113 (O_2113,N_48143,N_49520);
nand UO_2114 (O_2114,N_48925,N_48347);
and UO_2115 (O_2115,N_48859,N_48208);
and UO_2116 (O_2116,N_49314,N_49872);
nand UO_2117 (O_2117,N_48140,N_49986);
and UO_2118 (O_2118,N_49662,N_48822);
and UO_2119 (O_2119,N_48713,N_48686);
or UO_2120 (O_2120,N_48954,N_49254);
and UO_2121 (O_2121,N_48628,N_48906);
xnor UO_2122 (O_2122,N_49000,N_49129);
or UO_2123 (O_2123,N_48008,N_49208);
nor UO_2124 (O_2124,N_48478,N_48218);
nand UO_2125 (O_2125,N_48543,N_49553);
or UO_2126 (O_2126,N_48157,N_48836);
and UO_2127 (O_2127,N_48339,N_49297);
nor UO_2128 (O_2128,N_49410,N_48457);
or UO_2129 (O_2129,N_49987,N_49324);
or UO_2130 (O_2130,N_49334,N_48153);
nor UO_2131 (O_2131,N_48206,N_49256);
or UO_2132 (O_2132,N_48608,N_48337);
xor UO_2133 (O_2133,N_49792,N_49672);
or UO_2134 (O_2134,N_49900,N_49001);
nand UO_2135 (O_2135,N_48591,N_49598);
xor UO_2136 (O_2136,N_48160,N_48177);
xor UO_2137 (O_2137,N_49948,N_49868);
nor UO_2138 (O_2138,N_48530,N_48517);
nand UO_2139 (O_2139,N_49768,N_48009);
or UO_2140 (O_2140,N_48435,N_49463);
nor UO_2141 (O_2141,N_49005,N_48183);
nor UO_2142 (O_2142,N_48400,N_49443);
and UO_2143 (O_2143,N_48326,N_48216);
or UO_2144 (O_2144,N_48066,N_49875);
nand UO_2145 (O_2145,N_49556,N_48816);
nand UO_2146 (O_2146,N_48482,N_49711);
or UO_2147 (O_2147,N_49074,N_49201);
nor UO_2148 (O_2148,N_48139,N_48893);
and UO_2149 (O_2149,N_48243,N_48012);
nor UO_2150 (O_2150,N_49842,N_48014);
xor UO_2151 (O_2151,N_48273,N_48874);
nand UO_2152 (O_2152,N_48043,N_48871);
xnor UO_2153 (O_2153,N_49219,N_48901);
xor UO_2154 (O_2154,N_49944,N_48646);
nand UO_2155 (O_2155,N_48192,N_48070);
xnor UO_2156 (O_2156,N_49601,N_48063);
and UO_2157 (O_2157,N_49649,N_49332);
nand UO_2158 (O_2158,N_49965,N_48296);
or UO_2159 (O_2159,N_49708,N_48568);
nand UO_2160 (O_2160,N_48247,N_49850);
nand UO_2161 (O_2161,N_49270,N_48560);
nor UO_2162 (O_2162,N_48606,N_49814);
and UO_2163 (O_2163,N_48329,N_49985);
and UO_2164 (O_2164,N_48401,N_49174);
nor UO_2165 (O_2165,N_48418,N_48139);
nor UO_2166 (O_2166,N_48227,N_48150);
xnor UO_2167 (O_2167,N_48349,N_48503);
xnor UO_2168 (O_2168,N_48110,N_49488);
nor UO_2169 (O_2169,N_48442,N_49278);
or UO_2170 (O_2170,N_48934,N_48099);
and UO_2171 (O_2171,N_49397,N_49280);
nor UO_2172 (O_2172,N_48693,N_49655);
and UO_2173 (O_2173,N_49851,N_48501);
nor UO_2174 (O_2174,N_48100,N_49279);
nand UO_2175 (O_2175,N_48564,N_48007);
and UO_2176 (O_2176,N_49576,N_48246);
nand UO_2177 (O_2177,N_48995,N_49323);
or UO_2178 (O_2178,N_48086,N_49600);
nand UO_2179 (O_2179,N_48251,N_49784);
or UO_2180 (O_2180,N_48609,N_49976);
nand UO_2181 (O_2181,N_49333,N_48594);
and UO_2182 (O_2182,N_49268,N_48982);
nand UO_2183 (O_2183,N_49207,N_48375);
nand UO_2184 (O_2184,N_49505,N_48330);
or UO_2185 (O_2185,N_49695,N_48210);
xor UO_2186 (O_2186,N_48770,N_49017);
nand UO_2187 (O_2187,N_48696,N_49429);
xor UO_2188 (O_2188,N_48290,N_49826);
xnor UO_2189 (O_2189,N_48777,N_49690);
xnor UO_2190 (O_2190,N_49051,N_49541);
or UO_2191 (O_2191,N_49511,N_49888);
nor UO_2192 (O_2192,N_48423,N_48139);
or UO_2193 (O_2193,N_48771,N_49175);
and UO_2194 (O_2194,N_49113,N_49633);
or UO_2195 (O_2195,N_48975,N_48202);
and UO_2196 (O_2196,N_48919,N_49203);
or UO_2197 (O_2197,N_49835,N_48421);
xnor UO_2198 (O_2198,N_49492,N_49150);
and UO_2199 (O_2199,N_48798,N_49003);
or UO_2200 (O_2200,N_48854,N_49184);
nand UO_2201 (O_2201,N_48349,N_48227);
and UO_2202 (O_2202,N_48706,N_49585);
nand UO_2203 (O_2203,N_48954,N_49292);
or UO_2204 (O_2204,N_48481,N_48641);
nor UO_2205 (O_2205,N_49629,N_48351);
and UO_2206 (O_2206,N_49556,N_49520);
or UO_2207 (O_2207,N_48946,N_48015);
xnor UO_2208 (O_2208,N_49032,N_48353);
xnor UO_2209 (O_2209,N_49582,N_48906);
nand UO_2210 (O_2210,N_48608,N_48889);
nor UO_2211 (O_2211,N_48699,N_48057);
or UO_2212 (O_2212,N_48693,N_48228);
and UO_2213 (O_2213,N_48035,N_48569);
or UO_2214 (O_2214,N_48674,N_48955);
xor UO_2215 (O_2215,N_48314,N_48481);
or UO_2216 (O_2216,N_48621,N_48056);
and UO_2217 (O_2217,N_48196,N_49460);
nand UO_2218 (O_2218,N_48341,N_49726);
or UO_2219 (O_2219,N_49745,N_48684);
xnor UO_2220 (O_2220,N_49624,N_48169);
and UO_2221 (O_2221,N_49721,N_49936);
nor UO_2222 (O_2222,N_48123,N_49514);
xnor UO_2223 (O_2223,N_48800,N_48206);
xor UO_2224 (O_2224,N_48559,N_49234);
or UO_2225 (O_2225,N_49380,N_48138);
xor UO_2226 (O_2226,N_48402,N_49403);
xnor UO_2227 (O_2227,N_49878,N_48376);
or UO_2228 (O_2228,N_48197,N_49606);
and UO_2229 (O_2229,N_48149,N_48597);
nand UO_2230 (O_2230,N_48632,N_49708);
or UO_2231 (O_2231,N_49698,N_48887);
xnor UO_2232 (O_2232,N_48301,N_49247);
and UO_2233 (O_2233,N_49019,N_49307);
nand UO_2234 (O_2234,N_48896,N_49038);
xor UO_2235 (O_2235,N_49453,N_48365);
nor UO_2236 (O_2236,N_48872,N_48984);
and UO_2237 (O_2237,N_49014,N_48297);
xnor UO_2238 (O_2238,N_48733,N_48029);
and UO_2239 (O_2239,N_49413,N_48645);
nor UO_2240 (O_2240,N_48367,N_49833);
nand UO_2241 (O_2241,N_49889,N_49097);
xor UO_2242 (O_2242,N_48877,N_49390);
and UO_2243 (O_2243,N_48057,N_48537);
and UO_2244 (O_2244,N_48481,N_49408);
nor UO_2245 (O_2245,N_49486,N_48649);
nand UO_2246 (O_2246,N_49553,N_49470);
nor UO_2247 (O_2247,N_48975,N_48270);
or UO_2248 (O_2248,N_49751,N_48623);
nand UO_2249 (O_2249,N_49474,N_48797);
or UO_2250 (O_2250,N_49605,N_49037);
nor UO_2251 (O_2251,N_48226,N_49362);
xor UO_2252 (O_2252,N_49377,N_49036);
nand UO_2253 (O_2253,N_48734,N_49204);
and UO_2254 (O_2254,N_49983,N_49343);
xnor UO_2255 (O_2255,N_49865,N_48502);
and UO_2256 (O_2256,N_49159,N_49982);
nor UO_2257 (O_2257,N_49246,N_48317);
nor UO_2258 (O_2258,N_48528,N_48547);
xnor UO_2259 (O_2259,N_48206,N_49526);
nor UO_2260 (O_2260,N_49410,N_48023);
nand UO_2261 (O_2261,N_49630,N_48469);
nor UO_2262 (O_2262,N_49962,N_48654);
nor UO_2263 (O_2263,N_48410,N_48920);
nor UO_2264 (O_2264,N_49341,N_49097);
nand UO_2265 (O_2265,N_48726,N_49386);
xor UO_2266 (O_2266,N_49197,N_48049);
or UO_2267 (O_2267,N_48142,N_49529);
or UO_2268 (O_2268,N_48948,N_49100);
nor UO_2269 (O_2269,N_49028,N_49286);
nand UO_2270 (O_2270,N_49212,N_49906);
nor UO_2271 (O_2271,N_48480,N_49225);
nor UO_2272 (O_2272,N_49442,N_48292);
nand UO_2273 (O_2273,N_48800,N_48939);
nor UO_2274 (O_2274,N_49246,N_49223);
nand UO_2275 (O_2275,N_48176,N_49743);
xnor UO_2276 (O_2276,N_48295,N_48782);
or UO_2277 (O_2277,N_48376,N_49566);
nor UO_2278 (O_2278,N_49388,N_49357);
xnor UO_2279 (O_2279,N_48519,N_49663);
xnor UO_2280 (O_2280,N_48327,N_49521);
xor UO_2281 (O_2281,N_48733,N_48420);
nor UO_2282 (O_2282,N_48418,N_48241);
nand UO_2283 (O_2283,N_49320,N_48896);
and UO_2284 (O_2284,N_48383,N_49682);
nor UO_2285 (O_2285,N_48235,N_48424);
nand UO_2286 (O_2286,N_48118,N_48677);
and UO_2287 (O_2287,N_48950,N_49638);
xnor UO_2288 (O_2288,N_48114,N_49970);
nand UO_2289 (O_2289,N_49503,N_49084);
nor UO_2290 (O_2290,N_48313,N_49325);
xor UO_2291 (O_2291,N_49666,N_48801);
xnor UO_2292 (O_2292,N_49728,N_48620);
xor UO_2293 (O_2293,N_49698,N_48555);
nand UO_2294 (O_2294,N_48296,N_48097);
nand UO_2295 (O_2295,N_49502,N_49460);
nand UO_2296 (O_2296,N_48343,N_49956);
nor UO_2297 (O_2297,N_49348,N_49050);
or UO_2298 (O_2298,N_49144,N_48892);
nand UO_2299 (O_2299,N_49876,N_48329);
nand UO_2300 (O_2300,N_48481,N_49305);
and UO_2301 (O_2301,N_48386,N_48499);
xor UO_2302 (O_2302,N_48236,N_48992);
xnor UO_2303 (O_2303,N_48996,N_48617);
and UO_2304 (O_2304,N_48616,N_48939);
nor UO_2305 (O_2305,N_48905,N_48518);
nor UO_2306 (O_2306,N_48364,N_49307);
or UO_2307 (O_2307,N_49062,N_48757);
xnor UO_2308 (O_2308,N_48553,N_49423);
and UO_2309 (O_2309,N_49493,N_49148);
nand UO_2310 (O_2310,N_48388,N_49628);
xor UO_2311 (O_2311,N_49658,N_48118);
nor UO_2312 (O_2312,N_48525,N_48675);
and UO_2313 (O_2313,N_49345,N_48554);
and UO_2314 (O_2314,N_49870,N_48492);
and UO_2315 (O_2315,N_49593,N_49384);
or UO_2316 (O_2316,N_49405,N_48910);
and UO_2317 (O_2317,N_49170,N_48538);
or UO_2318 (O_2318,N_48199,N_49808);
nor UO_2319 (O_2319,N_48949,N_49527);
or UO_2320 (O_2320,N_49587,N_48094);
and UO_2321 (O_2321,N_48526,N_48425);
nand UO_2322 (O_2322,N_49470,N_48648);
and UO_2323 (O_2323,N_48880,N_49034);
and UO_2324 (O_2324,N_48448,N_48508);
xor UO_2325 (O_2325,N_48758,N_49757);
and UO_2326 (O_2326,N_48373,N_49003);
xnor UO_2327 (O_2327,N_49395,N_48397);
xor UO_2328 (O_2328,N_48000,N_48606);
and UO_2329 (O_2329,N_49469,N_48752);
xor UO_2330 (O_2330,N_48777,N_48968);
or UO_2331 (O_2331,N_48220,N_48556);
and UO_2332 (O_2332,N_48964,N_49514);
xnor UO_2333 (O_2333,N_49954,N_48861);
nor UO_2334 (O_2334,N_49046,N_48382);
nand UO_2335 (O_2335,N_48263,N_48508);
or UO_2336 (O_2336,N_48624,N_49780);
or UO_2337 (O_2337,N_49408,N_48999);
or UO_2338 (O_2338,N_49757,N_49258);
nor UO_2339 (O_2339,N_48123,N_49092);
and UO_2340 (O_2340,N_48409,N_49569);
nor UO_2341 (O_2341,N_48425,N_48044);
or UO_2342 (O_2342,N_49186,N_48471);
xor UO_2343 (O_2343,N_49739,N_49720);
and UO_2344 (O_2344,N_49243,N_49953);
xor UO_2345 (O_2345,N_48380,N_48197);
and UO_2346 (O_2346,N_48289,N_49971);
or UO_2347 (O_2347,N_48433,N_49564);
nand UO_2348 (O_2348,N_49044,N_48137);
nor UO_2349 (O_2349,N_49062,N_48113);
xor UO_2350 (O_2350,N_49989,N_49790);
xor UO_2351 (O_2351,N_48095,N_48697);
xnor UO_2352 (O_2352,N_49320,N_49808);
or UO_2353 (O_2353,N_49711,N_49235);
xnor UO_2354 (O_2354,N_48334,N_48175);
and UO_2355 (O_2355,N_49196,N_48880);
xnor UO_2356 (O_2356,N_48910,N_49806);
and UO_2357 (O_2357,N_48713,N_48949);
and UO_2358 (O_2358,N_48649,N_49718);
xnor UO_2359 (O_2359,N_48998,N_49871);
or UO_2360 (O_2360,N_49048,N_48831);
xor UO_2361 (O_2361,N_48675,N_48968);
nor UO_2362 (O_2362,N_49904,N_48984);
nor UO_2363 (O_2363,N_49392,N_48444);
or UO_2364 (O_2364,N_48597,N_49291);
and UO_2365 (O_2365,N_48427,N_48853);
nand UO_2366 (O_2366,N_48855,N_49103);
nor UO_2367 (O_2367,N_49028,N_48792);
xor UO_2368 (O_2368,N_49100,N_48029);
and UO_2369 (O_2369,N_49889,N_49401);
xnor UO_2370 (O_2370,N_48054,N_49637);
and UO_2371 (O_2371,N_48551,N_48315);
or UO_2372 (O_2372,N_49685,N_48828);
nor UO_2373 (O_2373,N_49597,N_48826);
xnor UO_2374 (O_2374,N_48548,N_48296);
nor UO_2375 (O_2375,N_49156,N_49921);
or UO_2376 (O_2376,N_48453,N_49857);
xnor UO_2377 (O_2377,N_48824,N_49634);
nand UO_2378 (O_2378,N_48325,N_48971);
nand UO_2379 (O_2379,N_48155,N_49263);
xnor UO_2380 (O_2380,N_48351,N_49954);
xor UO_2381 (O_2381,N_49893,N_48348);
xor UO_2382 (O_2382,N_48780,N_49118);
and UO_2383 (O_2383,N_49982,N_49149);
and UO_2384 (O_2384,N_49082,N_49125);
nand UO_2385 (O_2385,N_48914,N_49963);
nand UO_2386 (O_2386,N_48191,N_49189);
nand UO_2387 (O_2387,N_49572,N_49534);
and UO_2388 (O_2388,N_49255,N_48146);
nor UO_2389 (O_2389,N_49342,N_49769);
nor UO_2390 (O_2390,N_48456,N_48020);
and UO_2391 (O_2391,N_49451,N_48813);
and UO_2392 (O_2392,N_49951,N_49039);
nor UO_2393 (O_2393,N_48734,N_49996);
nor UO_2394 (O_2394,N_49912,N_49449);
and UO_2395 (O_2395,N_49978,N_48408);
nor UO_2396 (O_2396,N_49785,N_49623);
xor UO_2397 (O_2397,N_49539,N_48202);
xor UO_2398 (O_2398,N_49641,N_49705);
or UO_2399 (O_2399,N_49979,N_48283);
or UO_2400 (O_2400,N_48819,N_48104);
or UO_2401 (O_2401,N_49775,N_48099);
xor UO_2402 (O_2402,N_48271,N_48468);
xnor UO_2403 (O_2403,N_49476,N_49023);
nand UO_2404 (O_2404,N_48057,N_49488);
nor UO_2405 (O_2405,N_48102,N_48325);
xnor UO_2406 (O_2406,N_49837,N_49255);
and UO_2407 (O_2407,N_48491,N_48604);
or UO_2408 (O_2408,N_49799,N_48414);
nor UO_2409 (O_2409,N_49444,N_48194);
and UO_2410 (O_2410,N_48135,N_48727);
nand UO_2411 (O_2411,N_48617,N_48690);
nor UO_2412 (O_2412,N_48288,N_48667);
nor UO_2413 (O_2413,N_49004,N_49877);
or UO_2414 (O_2414,N_48578,N_48314);
nor UO_2415 (O_2415,N_48427,N_49314);
and UO_2416 (O_2416,N_49169,N_48004);
and UO_2417 (O_2417,N_48710,N_48272);
nor UO_2418 (O_2418,N_48261,N_48194);
nor UO_2419 (O_2419,N_48201,N_49214);
or UO_2420 (O_2420,N_49223,N_49852);
nand UO_2421 (O_2421,N_49875,N_49330);
nand UO_2422 (O_2422,N_49094,N_49337);
or UO_2423 (O_2423,N_48500,N_48736);
or UO_2424 (O_2424,N_49704,N_48965);
nor UO_2425 (O_2425,N_49377,N_49963);
and UO_2426 (O_2426,N_48596,N_49829);
or UO_2427 (O_2427,N_48623,N_48982);
or UO_2428 (O_2428,N_49263,N_49605);
nand UO_2429 (O_2429,N_49979,N_48026);
xor UO_2430 (O_2430,N_49605,N_48630);
nor UO_2431 (O_2431,N_49993,N_49797);
nand UO_2432 (O_2432,N_49950,N_49313);
and UO_2433 (O_2433,N_49716,N_48724);
and UO_2434 (O_2434,N_48844,N_49553);
or UO_2435 (O_2435,N_48893,N_48685);
and UO_2436 (O_2436,N_49577,N_48069);
nor UO_2437 (O_2437,N_48175,N_48103);
nand UO_2438 (O_2438,N_48332,N_48685);
xor UO_2439 (O_2439,N_49817,N_48219);
and UO_2440 (O_2440,N_48204,N_48039);
xnor UO_2441 (O_2441,N_49911,N_48379);
or UO_2442 (O_2442,N_48670,N_49689);
and UO_2443 (O_2443,N_49558,N_48446);
nor UO_2444 (O_2444,N_49104,N_48073);
xnor UO_2445 (O_2445,N_49199,N_49408);
or UO_2446 (O_2446,N_49358,N_48391);
xnor UO_2447 (O_2447,N_48592,N_49900);
xor UO_2448 (O_2448,N_48071,N_49279);
nand UO_2449 (O_2449,N_48709,N_49605);
nor UO_2450 (O_2450,N_49338,N_49477);
or UO_2451 (O_2451,N_49112,N_48302);
xor UO_2452 (O_2452,N_49676,N_48617);
or UO_2453 (O_2453,N_49508,N_48590);
and UO_2454 (O_2454,N_48077,N_48013);
nor UO_2455 (O_2455,N_49963,N_49872);
xor UO_2456 (O_2456,N_48275,N_49667);
and UO_2457 (O_2457,N_49820,N_48677);
or UO_2458 (O_2458,N_48962,N_48887);
xnor UO_2459 (O_2459,N_49206,N_48137);
nand UO_2460 (O_2460,N_49030,N_48003);
nand UO_2461 (O_2461,N_49334,N_49513);
nand UO_2462 (O_2462,N_48380,N_48907);
nor UO_2463 (O_2463,N_48053,N_48753);
nand UO_2464 (O_2464,N_48900,N_48586);
or UO_2465 (O_2465,N_48207,N_49000);
or UO_2466 (O_2466,N_48039,N_48910);
and UO_2467 (O_2467,N_48533,N_48772);
nand UO_2468 (O_2468,N_48444,N_49014);
xor UO_2469 (O_2469,N_49339,N_48991);
nand UO_2470 (O_2470,N_49385,N_48359);
nand UO_2471 (O_2471,N_49652,N_49427);
xor UO_2472 (O_2472,N_48633,N_49302);
xnor UO_2473 (O_2473,N_49638,N_49104);
and UO_2474 (O_2474,N_48473,N_48302);
or UO_2475 (O_2475,N_48231,N_49812);
and UO_2476 (O_2476,N_49531,N_48124);
or UO_2477 (O_2477,N_49482,N_49964);
xnor UO_2478 (O_2478,N_48120,N_49634);
or UO_2479 (O_2479,N_49914,N_48909);
nand UO_2480 (O_2480,N_49761,N_48109);
xor UO_2481 (O_2481,N_48265,N_49295);
and UO_2482 (O_2482,N_49049,N_49906);
xor UO_2483 (O_2483,N_48113,N_49443);
or UO_2484 (O_2484,N_49759,N_49401);
xnor UO_2485 (O_2485,N_49170,N_49293);
nand UO_2486 (O_2486,N_48866,N_48720);
and UO_2487 (O_2487,N_48186,N_48838);
nor UO_2488 (O_2488,N_49226,N_49786);
xor UO_2489 (O_2489,N_48640,N_49373);
xnor UO_2490 (O_2490,N_48286,N_48858);
nand UO_2491 (O_2491,N_48771,N_49725);
nand UO_2492 (O_2492,N_48828,N_48420);
or UO_2493 (O_2493,N_48548,N_49292);
and UO_2494 (O_2494,N_49253,N_48527);
or UO_2495 (O_2495,N_49283,N_49243);
or UO_2496 (O_2496,N_48902,N_48114);
xor UO_2497 (O_2497,N_48267,N_48496);
xor UO_2498 (O_2498,N_49701,N_48274);
and UO_2499 (O_2499,N_48967,N_48394);
or UO_2500 (O_2500,N_49664,N_49909);
nand UO_2501 (O_2501,N_49806,N_49089);
nor UO_2502 (O_2502,N_49803,N_48311);
or UO_2503 (O_2503,N_48439,N_48014);
nor UO_2504 (O_2504,N_48119,N_48860);
xnor UO_2505 (O_2505,N_49074,N_49782);
nor UO_2506 (O_2506,N_48197,N_48921);
xor UO_2507 (O_2507,N_49881,N_49996);
and UO_2508 (O_2508,N_48733,N_48851);
nor UO_2509 (O_2509,N_48392,N_49668);
xor UO_2510 (O_2510,N_49736,N_48925);
and UO_2511 (O_2511,N_49390,N_49299);
and UO_2512 (O_2512,N_49981,N_48040);
xor UO_2513 (O_2513,N_48392,N_48750);
nand UO_2514 (O_2514,N_49934,N_49553);
or UO_2515 (O_2515,N_48030,N_48487);
xnor UO_2516 (O_2516,N_48176,N_48259);
or UO_2517 (O_2517,N_49578,N_48007);
xor UO_2518 (O_2518,N_49870,N_49690);
nand UO_2519 (O_2519,N_49503,N_49340);
xnor UO_2520 (O_2520,N_49102,N_49331);
nor UO_2521 (O_2521,N_49011,N_49331);
xnor UO_2522 (O_2522,N_48188,N_48939);
or UO_2523 (O_2523,N_48433,N_49438);
nor UO_2524 (O_2524,N_49904,N_48607);
nor UO_2525 (O_2525,N_48997,N_49824);
or UO_2526 (O_2526,N_49390,N_48287);
nor UO_2527 (O_2527,N_48045,N_48485);
nand UO_2528 (O_2528,N_48417,N_49133);
or UO_2529 (O_2529,N_48499,N_48852);
xor UO_2530 (O_2530,N_48335,N_48299);
nand UO_2531 (O_2531,N_49923,N_48784);
or UO_2532 (O_2532,N_49451,N_49712);
nand UO_2533 (O_2533,N_48400,N_48346);
nor UO_2534 (O_2534,N_49211,N_49059);
xnor UO_2535 (O_2535,N_48397,N_49568);
or UO_2536 (O_2536,N_48373,N_48781);
nand UO_2537 (O_2537,N_49963,N_49321);
nor UO_2538 (O_2538,N_48180,N_49190);
nor UO_2539 (O_2539,N_49848,N_49252);
or UO_2540 (O_2540,N_48440,N_49386);
xor UO_2541 (O_2541,N_49139,N_48827);
nand UO_2542 (O_2542,N_48515,N_49633);
xor UO_2543 (O_2543,N_49908,N_48089);
and UO_2544 (O_2544,N_49291,N_48579);
nor UO_2545 (O_2545,N_48674,N_49332);
nand UO_2546 (O_2546,N_49036,N_48762);
nand UO_2547 (O_2547,N_49104,N_49253);
xnor UO_2548 (O_2548,N_48684,N_49765);
or UO_2549 (O_2549,N_49556,N_48646);
nor UO_2550 (O_2550,N_48977,N_49205);
xor UO_2551 (O_2551,N_48393,N_48824);
or UO_2552 (O_2552,N_48568,N_49574);
and UO_2553 (O_2553,N_48981,N_49191);
nor UO_2554 (O_2554,N_48078,N_48771);
and UO_2555 (O_2555,N_49591,N_48300);
or UO_2556 (O_2556,N_49021,N_49868);
nand UO_2557 (O_2557,N_48770,N_48181);
nor UO_2558 (O_2558,N_49666,N_49581);
nand UO_2559 (O_2559,N_48100,N_49688);
or UO_2560 (O_2560,N_48911,N_49738);
xnor UO_2561 (O_2561,N_49318,N_48338);
and UO_2562 (O_2562,N_49885,N_49188);
xnor UO_2563 (O_2563,N_48334,N_49283);
nand UO_2564 (O_2564,N_49647,N_48596);
nand UO_2565 (O_2565,N_48942,N_48198);
xor UO_2566 (O_2566,N_48246,N_49846);
nor UO_2567 (O_2567,N_49206,N_48235);
nand UO_2568 (O_2568,N_48632,N_48037);
and UO_2569 (O_2569,N_49615,N_48194);
nand UO_2570 (O_2570,N_49568,N_49751);
or UO_2571 (O_2571,N_49895,N_49160);
and UO_2572 (O_2572,N_49502,N_49051);
or UO_2573 (O_2573,N_48384,N_49668);
and UO_2574 (O_2574,N_48039,N_49639);
or UO_2575 (O_2575,N_49032,N_48326);
or UO_2576 (O_2576,N_49939,N_49628);
xnor UO_2577 (O_2577,N_49286,N_48352);
xor UO_2578 (O_2578,N_49733,N_49280);
nand UO_2579 (O_2579,N_49613,N_49448);
nor UO_2580 (O_2580,N_48585,N_48320);
nand UO_2581 (O_2581,N_48556,N_49555);
nand UO_2582 (O_2582,N_49690,N_49705);
xor UO_2583 (O_2583,N_49768,N_48079);
nor UO_2584 (O_2584,N_49252,N_49216);
nor UO_2585 (O_2585,N_49103,N_49227);
nor UO_2586 (O_2586,N_48379,N_48884);
nand UO_2587 (O_2587,N_49744,N_49909);
and UO_2588 (O_2588,N_49401,N_48034);
nor UO_2589 (O_2589,N_49216,N_48519);
nor UO_2590 (O_2590,N_48062,N_49417);
xnor UO_2591 (O_2591,N_48209,N_49564);
nor UO_2592 (O_2592,N_48761,N_49271);
nand UO_2593 (O_2593,N_48888,N_48277);
and UO_2594 (O_2594,N_49270,N_48995);
or UO_2595 (O_2595,N_49326,N_48479);
and UO_2596 (O_2596,N_49100,N_49555);
and UO_2597 (O_2597,N_49866,N_49210);
or UO_2598 (O_2598,N_49249,N_49771);
xnor UO_2599 (O_2599,N_48203,N_49307);
nor UO_2600 (O_2600,N_48564,N_49847);
nand UO_2601 (O_2601,N_49119,N_48913);
and UO_2602 (O_2602,N_48324,N_49388);
xor UO_2603 (O_2603,N_49663,N_49940);
xor UO_2604 (O_2604,N_49227,N_49042);
nor UO_2605 (O_2605,N_48713,N_49323);
xor UO_2606 (O_2606,N_49013,N_49947);
nor UO_2607 (O_2607,N_48805,N_49446);
xor UO_2608 (O_2608,N_48052,N_49430);
xor UO_2609 (O_2609,N_48768,N_49842);
and UO_2610 (O_2610,N_49720,N_48789);
nand UO_2611 (O_2611,N_49143,N_48763);
nor UO_2612 (O_2612,N_48401,N_48049);
nand UO_2613 (O_2613,N_48913,N_48637);
xnor UO_2614 (O_2614,N_48658,N_48194);
xnor UO_2615 (O_2615,N_49158,N_48751);
and UO_2616 (O_2616,N_49563,N_49295);
nand UO_2617 (O_2617,N_48867,N_49238);
xor UO_2618 (O_2618,N_49707,N_48518);
nand UO_2619 (O_2619,N_48675,N_48412);
and UO_2620 (O_2620,N_49230,N_48503);
or UO_2621 (O_2621,N_49383,N_48344);
nand UO_2622 (O_2622,N_48841,N_48360);
nand UO_2623 (O_2623,N_49066,N_49471);
and UO_2624 (O_2624,N_49169,N_48792);
or UO_2625 (O_2625,N_48447,N_48835);
or UO_2626 (O_2626,N_49517,N_48404);
or UO_2627 (O_2627,N_49429,N_49003);
or UO_2628 (O_2628,N_49820,N_49958);
nor UO_2629 (O_2629,N_49714,N_48567);
or UO_2630 (O_2630,N_48163,N_49049);
nor UO_2631 (O_2631,N_49843,N_49146);
and UO_2632 (O_2632,N_48200,N_49789);
xor UO_2633 (O_2633,N_48977,N_48388);
nand UO_2634 (O_2634,N_48556,N_49010);
and UO_2635 (O_2635,N_48505,N_49982);
nor UO_2636 (O_2636,N_48377,N_48923);
nor UO_2637 (O_2637,N_48945,N_48479);
nand UO_2638 (O_2638,N_48398,N_48862);
nor UO_2639 (O_2639,N_48566,N_49863);
xor UO_2640 (O_2640,N_49929,N_48510);
nor UO_2641 (O_2641,N_49500,N_49045);
and UO_2642 (O_2642,N_49774,N_49270);
nand UO_2643 (O_2643,N_48318,N_48396);
nand UO_2644 (O_2644,N_49560,N_49366);
xor UO_2645 (O_2645,N_49675,N_48114);
xor UO_2646 (O_2646,N_49158,N_48781);
xor UO_2647 (O_2647,N_48496,N_48028);
or UO_2648 (O_2648,N_49413,N_48756);
nor UO_2649 (O_2649,N_49432,N_48568);
or UO_2650 (O_2650,N_49102,N_49860);
nor UO_2651 (O_2651,N_48170,N_49171);
nor UO_2652 (O_2652,N_49508,N_49346);
or UO_2653 (O_2653,N_48742,N_48744);
nand UO_2654 (O_2654,N_48772,N_48064);
nor UO_2655 (O_2655,N_48857,N_49350);
or UO_2656 (O_2656,N_49454,N_48322);
nand UO_2657 (O_2657,N_48039,N_48764);
nor UO_2658 (O_2658,N_48332,N_48954);
xor UO_2659 (O_2659,N_48501,N_48530);
nor UO_2660 (O_2660,N_48957,N_48037);
and UO_2661 (O_2661,N_49720,N_49776);
nand UO_2662 (O_2662,N_48076,N_49817);
and UO_2663 (O_2663,N_49868,N_49488);
nand UO_2664 (O_2664,N_48589,N_49588);
nor UO_2665 (O_2665,N_49795,N_49002);
nor UO_2666 (O_2666,N_48713,N_48787);
nor UO_2667 (O_2667,N_49336,N_49440);
nor UO_2668 (O_2668,N_49364,N_48339);
and UO_2669 (O_2669,N_49584,N_49524);
nor UO_2670 (O_2670,N_48330,N_49235);
and UO_2671 (O_2671,N_49252,N_49167);
or UO_2672 (O_2672,N_49946,N_48632);
xnor UO_2673 (O_2673,N_49711,N_48589);
and UO_2674 (O_2674,N_49670,N_49700);
or UO_2675 (O_2675,N_48164,N_48907);
xnor UO_2676 (O_2676,N_48014,N_48007);
nor UO_2677 (O_2677,N_48430,N_48772);
nand UO_2678 (O_2678,N_49972,N_49125);
and UO_2679 (O_2679,N_48199,N_49275);
nor UO_2680 (O_2680,N_49974,N_49105);
nor UO_2681 (O_2681,N_49729,N_49115);
nor UO_2682 (O_2682,N_49475,N_49862);
nand UO_2683 (O_2683,N_48020,N_48003);
xnor UO_2684 (O_2684,N_49069,N_48017);
and UO_2685 (O_2685,N_49461,N_49053);
nor UO_2686 (O_2686,N_49636,N_48242);
and UO_2687 (O_2687,N_49537,N_49134);
and UO_2688 (O_2688,N_48549,N_49660);
xor UO_2689 (O_2689,N_48371,N_48070);
nor UO_2690 (O_2690,N_48852,N_49906);
xor UO_2691 (O_2691,N_48401,N_48454);
or UO_2692 (O_2692,N_49459,N_48296);
or UO_2693 (O_2693,N_49936,N_49678);
or UO_2694 (O_2694,N_48696,N_48706);
nand UO_2695 (O_2695,N_49774,N_49747);
nor UO_2696 (O_2696,N_48827,N_48577);
nor UO_2697 (O_2697,N_49066,N_49123);
xor UO_2698 (O_2698,N_48953,N_48302);
nand UO_2699 (O_2699,N_48356,N_48849);
nor UO_2700 (O_2700,N_48503,N_48679);
or UO_2701 (O_2701,N_49138,N_48350);
nand UO_2702 (O_2702,N_48106,N_49193);
and UO_2703 (O_2703,N_49372,N_49344);
xor UO_2704 (O_2704,N_49803,N_49203);
nor UO_2705 (O_2705,N_48612,N_49715);
nand UO_2706 (O_2706,N_49587,N_48625);
xnor UO_2707 (O_2707,N_49586,N_48819);
xor UO_2708 (O_2708,N_49949,N_49927);
xnor UO_2709 (O_2709,N_48735,N_49705);
nand UO_2710 (O_2710,N_48096,N_48872);
and UO_2711 (O_2711,N_48176,N_48800);
nor UO_2712 (O_2712,N_48203,N_48313);
or UO_2713 (O_2713,N_48587,N_48153);
and UO_2714 (O_2714,N_49715,N_49459);
xnor UO_2715 (O_2715,N_48176,N_48036);
and UO_2716 (O_2716,N_49362,N_49035);
xor UO_2717 (O_2717,N_48227,N_49120);
nor UO_2718 (O_2718,N_48092,N_49570);
nor UO_2719 (O_2719,N_48604,N_48881);
or UO_2720 (O_2720,N_49412,N_49112);
nand UO_2721 (O_2721,N_49464,N_49739);
xor UO_2722 (O_2722,N_49446,N_49305);
and UO_2723 (O_2723,N_49653,N_48889);
xor UO_2724 (O_2724,N_48581,N_49726);
or UO_2725 (O_2725,N_48734,N_49902);
and UO_2726 (O_2726,N_49184,N_48222);
nor UO_2727 (O_2727,N_48874,N_49355);
and UO_2728 (O_2728,N_49083,N_48585);
nand UO_2729 (O_2729,N_49744,N_49676);
and UO_2730 (O_2730,N_49933,N_48433);
or UO_2731 (O_2731,N_49626,N_49276);
or UO_2732 (O_2732,N_48179,N_48236);
and UO_2733 (O_2733,N_49841,N_48242);
and UO_2734 (O_2734,N_48678,N_49800);
nor UO_2735 (O_2735,N_49819,N_48156);
or UO_2736 (O_2736,N_48989,N_49163);
and UO_2737 (O_2737,N_48284,N_49084);
nand UO_2738 (O_2738,N_49609,N_48869);
and UO_2739 (O_2739,N_49013,N_49436);
or UO_2740 (O_2740,N_49298,N_49717);
nand UO_2741 (O_2741,N_48886,N_48447);
or UO_2742 (O_2742,N_48590,N_49603);
nand UO_2743 (O_2743,N_49825,N_48969);
xnor UO_2744 (O_2744,N_49539,N_48857);
or UO_2745 (O_2745,N_48533,N_49872);
and UO_2746 (O_2746,N_48730,N_49683);
nand UO_2747 (O_2747,N_49853,N_48228);
xnor UO_2748 (O_2748,N_49842,N_49698);
nand UO_2749 (O_2749,N_48412,N_49866);
and UO_2750 (O_2750,N_48785,N_49160);
or UO_2751 (O_2751,N_49902,N_49747);
nand UO_2752 (O_2752,N_48507,N_48005);
nand UO_2753 (O_2753,N_49738,N_49115);
nor UO_2754 (O_2754,N_49590,N_49559);
nand UO_2755 (O_2755,N_48498,N_48379);
xnor UO_2756 (O_2756,N_48805,N_49530);
and UO_2757 (O_2757,N_48174,N_49060);
nand UO_2758 (O_2758,N_48311,N_48978);
nor UO_2759 (O_2759,N_49039,N_49452);
nor UO_2760 (O_2760,N_48356,N_48730);
nand UO_2761 (O_2761,N_49222,N_48838);
nand UO_2762 (O_2762,N_48195,N_49810);
or UO_2763 (O_2763,N_48374,N_49393);
nand UO_2764 (O_2764,N_48458,N_49908);
xnor UO_2765 (O_2765,N_48587,N_49663);
nand UO_2766 (O_2766,N_48171,N_49412);
nand UO_2767 (O_2767,N_49372,N_48039);
xnor UO_2768 (O_2768,N_48915,N_49197);
and UO_2769 (O_2769,N_48134,N_48136);
and UO_2770 (O_2770,N_49695,N_49096);
or UO_2771 (O_2771,N_49636,N_48977);
xnor UO_2772 (O_2772,N_49834,N_49901);
and UO_2773 (O_2773,N_48455,N_49125);
xor UO_2774 (O_2774,N_49105,N_48249);
or UO_2775 (O_2775,N_48714,N_49890);
xnor UO_2776 (O_2776,N_49876,N_48663);
nand UO_2777 (O_2777,N_48015,N_49592);
xnor UO_2778 (O_2778,N_48775,N_48655);
or UO_2779 (O_2779,N_49384,N_48604);
nor UO_2780 (O_2780,N_48101,N_49540);
and UO_2781 (O_2781,N_49097,N_49713);
and UO_2782 (O_2782,N_48026,N_49838);
nor UO_2783 (O_2783,N_48966,N_49894);
or UO_2784 (O_2784,N_49798,N_49521);
nand UO_2785 (O_2785,N_49718,N_49421);
nor UO_2786 (O_2786,N_48292,N_49631);
nor UO_2787 (O_2787,N_49355,N_49592);
or UO_2788 (O_2788,N_49642,N_49091);
xor UO_2789 (O_2789,N_49731,N_49027);
nor UO_2790 (O_2790,N_49343,N_48812);
or UO_2791 (O_2791,N_48304,N_48268);
and UO_2792 (O_2792,N_48647,N_48053);
xor UO_2793 (O_2793,N_49877,N_48284);
and UO_2794 (O_2794,N_48613,N_49926);
nand UO_2795 (O_2795,N_48381,N_48855);
nor UO_2796 (O_2796,N_49010,N_48534);
or UO_2797 (O_2797,N_48107,N_49353);
nor UO_2798 (O_2798,N_49379,N_48908);
nand UO_2799 (O_2799,N_49109,N_49253);
nor UO_2800 (O_2800,N_48649,N_48326);
and UO_2801 (O_2801,N_49323,N_49125);
and UO_2802 (O_2802,N_48544,N_49305);
nor UO_2803 (O_2803,N_49974,N_48603);
and UO_2804 (O_2804,N_49398,N_48884);
nand UO_2805 (O_2805,N_49773,N_49485);
and UO_2806 (O_2806,N_48693,N_49444);
nor UO_2807 (O_2807,N_49523,N_49205);
nand UO_2808 (O_2808,N_48684,N_48593);
nand UO_2809 (O_2809,N_49712,N_48833);
and UO_2810 (O_2810,N_48520,N_49598);
and UO_2811 (O_2811,N_49680,N_49242);
and UO_2812 (O_2812,N_48838,N_49641);
nor UO_2813 (O_2813,N_48181,N_48674);
or UO_2814 (O_2814,N_48089,N_48388);
or UO_2815 (O_2815,N_49216,N_48336);
or UO_2816 (O_2816,N_48835,N_48511);
xnor UO_2817 (O_2817,N_48686,N_48920);
or UO_2818 (O_2818,N_49604,N_49849);
xnor UO_2819 (O_2819,N_48430,N_48967);
and UO_2820 (O_2820,N_48820,N_49349);
nor UO_2821 (O_2821,N_49372,N_48321);
nand UO_2822 (O_2822,N_49095,N_49385);
or UO_2823 (O_2823,N_49114,N_49159);
or UO_2824 (O_2824,N_48371,N_49883);
or UO_2825 (O_2825,N_48953,N_49436);
nand UO_2826 (O_2826,N_48356,N_48933);
or UO_2827 (O_2827,N_49138,N_48135);
nand UO_2828 (O_2828,N_48413,N_48420);
nor UO_2829 (O_2829,N_49397,N_48004);
or UO_2830 (O_2830,N_49839,N_48397);
nor UO_2831 (O_2831,N_48767,N_49657);
xor UO_2832 (O_2832,N_48185,N_49470);
and UO_2833 (O_2833,N_48176,N_48559);
nand UO_2834 (O_2834,N_49499,N_48786);
or UO_2835 (O_2835,N_48485,N_49364);
xor UO_2836 (O_2836,N_49748,N_48165);
xnor UO_2837 (O_2837,N_48084,N_48306);
or UO_2838 (O_2838,N_48727,N_49967);
nor UO_2839 (O_2839,N_49143,N_48218);
or UO_2840 (O_2840,N_48443,N_48814);
nand UO_2841 (O_2841,N_48398,N_49135);
xnor UO_2842 (O_2842,N_48210,N_49816);
nand UO_2843 (O_2843,N_48812,N_49589);
and UO_2844 (O_2844,N_48724,N_48560);
and UO_2845 (O_2845,N_48435,N_49101);
xnor UO_2846 (O_2846,N_49804,N_48691);
nor UO_2847 (O_2847,N_48891,N_49820);
and UO_2848 (O_2848,N_48335,N_49922);
nor UO_2849 (O_2849,N_48898,N_48461);
nand UO_2850 (O_2850,N_48911,N_49847);
nor UO_2851 (O_2851,N_48610,N_48805);
xor UO_2852 (O_2852,N_48475,N_48991);
nor UO_2853 (O_2853,N_49502,N_49457);
and UO_2854 (O_2854,N_49564,N_49786);
xor UO_2855 (O_2855,N_49381,N_49084);
nor UO_2856 (O_2856,N_48696,N_49712);
or UO_2857 (O_2857,N_48023,N_48745);
or UO_2858 (O_2858,N_49190,N_49125);
or UO_2859 (O_2859,N_48320,N_48016);
nand UO_2860 (O_2860,N_49928,N_48442);
or UO_2861 (O_2861,N_49550,N_48365);
nand UO_2862 (O_2862,N_48898,N_48423);
or UO_2863 (O_2863,N_49125,N_48958);
or UO_2864 (O_2864,N_49130,N_49914);
and UO_2865 (O_2865,N_48317,N_49947);
and UO_2866 (O_2866,N_48669,N_48037);
nor UO_2867 (O_2867,N_49276,N_48415);
xor UO_2868 (O_2868,N_48190,N_49215);
or UO_2869 (O_2869,N_48487,N_49630);
and UO_2870 (O_2870,N_48570,N_49364);
and UO_2871 (O_2871,N_48637,N_48529);
nand UO_2872 (O_2872,N_49956,N_48602);
nand UO_2873 (O_2873,N_49224,N_48861);
nand UO_2874 (O_2874,N_49027,N_49421);
or UO_2875 (O_2875,N_49413,N_49928);
or UO_2876 (O_2876,N_49777,N_49553);
nand UO_2877 (O_2877,N_49317,N_49208);
nor UO_2878 (O_2878,N_48382,N_48804);
nor UO_2879 (O_2879,N_48147,N_49439);
nand UO_2880 (O_2880,N_48114,N_49754);
and UO_2881 (O_2881,N_49135,N_49574);
nor UO_2882 (O_2882,N_49872,N_49824);
or UO_2883 (O_2883,N_48032,N_48305);
nor UO_2884 (O_2884,N_49948,N_49163);
nand UO_2885 (O_2885,N_49646,N_48232);
xnor UO_2886 (O_2886,N_49366,N_49060);
nand UO_2887 (O_2887,N_49140,N_49157);
xnor UO_2888 (O_2888,N_48824,N_49625);
or UO_2889 (O_2889,N_48350,N_49562);
or UO_2890 (O_2890,N_48186,N_48805);
nor UO_2891 (O_2891,N_48821,N_49228);
or UO_2892 (O_2892,N_49588,N_49724);
and UO_2893 (O_2893,N_49508,N_49520);
or UO_2894 (O_2894,N_49945,N_49766);
or UO_2895 (O_2895,N_48953,N_49453);
and UO_2896 (O_2896,N_48204,N_48690);
nand UO_2897 (O_2897,N_48272,N_48286);
nand UO_2898 (O_2898,N_49297,N_49661);
xnor UO_2899 (O_2899,N_48017,N_48605);
nand UO_2900 (O_2900,N_48361,N_49018);
nor UO_2901 (O_2901,N_48872,N_49096);
nand UO_2902 (O_2902,N_49618,N_48912);
nor UO_2903 (O_2903,N_49720,N_48820);
nand UO_2904 (O_2904,N_49582,N_48458);
nor UO_2905 (O_2905,N_49956,N_48116);
and UO_2906 (O_2906,N_48010,N_48623);
or UO_2907 (O_2907,N_48120,N_48430);
nand UO_2908 (O_2908,N_48876,N_49809);
nor UO_2909 (O_2909,N_48148,N_48622);
xor UO_2910 (O_2910,N_48825,N_48579);
and UO_2911 (O_2911,N_48844,N_49671);
nand UO_2912 (O_2912,N_48248,N_49959);
or UO_2913 (O_2913,N_49200,N_48761);
and UO_2914 (O_2914,N_49315,N_48996);
xnor UO_2915 (O_2915,N_48645,N_48908);
xnor UO_2916 (O_2916,N_48599,N_48862);
xnor UO_2917 (O_2917,N_49367,N_49476);
xnor UO_2918 (O_2918,N_49829,N_48433);
or UO_2919 (O_2919,N_48058,N_49740);
nor UO_2920 (O_2920,N_49744,N_48220);
nor UO_2921 (O_2921,N_49091,N_48973);
nor UO_2922 (O_2922,N_48832,N_48933);
xnor UO_2923 (O_2923,N_48963,N_48558);
nor UO_2924 (O_2924,N_48732,N_49842);
and UO_2925 (O_2925,N_48136,N_49426);
nor UO_2926 (O_2926,N_48866,N_48275);
xor UO_2927 (O_2927,N_48249,N_49992);
or UO_2928 (O_2928,N_49101,N_48069);
or UO_2929 (O_2929,N_48600,N_49494);
nand UO_2930 (O_2930,N_49766,N_48558);
or UO_2931 (O_2931,N_48179,N_49202);
xnor UO_2932 (O_2932,N_48013,N_49715);
nor UO_2933 (O_2933,N_49066,N_49437);
and UO_2934 (O_2934,N_49141,N_48770);
nor UO_2935 (O_2935,N_48427,N_49845);
or UO_2936 (O_2936,N_48682,N_48959);
xor UO_2937 (O_2937,N_49214,N_48006);
nor UO_2938 (O_2938,N_49254,N_48726);
xnor UO_2939 (O_2939,N_48914,N_49893);
or UO_2940 (O_2940,N_48030,N_48463);
nor UO_2941 (O_2941,N_49729,N_48989);
and UO_2942 (O_2942,N_48182,N_49061);
and UO_2943 (O_2943,N_48807,N_48811);
and UO_2944 (O_2944,N_48580,N_48735);
and UO_2945 (O_2945,N_49049,N_48333);
or UO_2946 (O_2946,N_49648,N_48576);
xnor UO_2947 (O_2947,N_49599,N_48853);
nor UO_2948 (O_2948,N_48086,N_49608);
and UO_2949 (O_2949,N_48564,N_49736);
or UO_2950 (O_2950,N_49419,N_49659);
nor UO_2951 (O_2951,N_48078,N_48126);
xor UO_2952 (O_2952,N_49111,N_48489);
or UO_2953 (O_2953,N_48158,N_49518);
nor UO_2954 (O_2954,N_48804,N_49559);
and UO_2955 (O_2955,N_48157,N_48547);
and UO_2956 (O_2956,N_48652,N_49525);
xnor UO_2957 (O_2957,N_49409,N_49158);
or UO_2958 (O_2958,N_49126,N_48416);
nor UO_2959 (O_2959,N_48146,N_48541);
nand UO_2960 (O_2960,N_49970,N_49862);
nand UO_2961 (O_2961,N_49955,N_48215);
or UO_2962 (O_2962,N_48687,N_49449);
and UO_2963 (O_2963,N_48241,N_49963);
or UO_2964 (O_2964,N_49792,N_48991);
and UO_2965 (O_2965,N_49453,N_48340);
or UO_2966 (O_2966,N_48132,N_48134);
xor UO_2967 (O_2967,N_48845,N_49064);
nand UO_2968 (O_2968,N_49414,N_49973);
and UO_2969 (O_2969,N_48773,N_48866);
and UO_2970 (O_2970,N_49839,N_49673);
and UO_2971 (O_2971,N_48234,N_48679);
or UO_2972 (O_2972,N_49775,N_48232);
or UO_2973 (O_2973,N_49530,N_49861);
nor UO_2974 (O_2974,N_49683,N_49104);
and UO_2975 (O_2975,N_49768,N_48941);
and UO_2976 (O_2976,N_49068,N_49507);
nand UO_2977 (O_2977,N_48435,N_48664);
and UO_2978 (O_2978,N_49656,N_49281);
nand UO_2979 (O_2979,N_49137,N_49262);
and UO_2980 (O_2980,N_49433,N_48945);
nor UO_2981 (O_2981,N_49472,N_49479);
nor UO_2982 (O_2982,N_49900,N_48314);
nor UO_2983 (O_2983,N_49260,N_49549);
nor UO_2984 (O_2984,N_48854,N_48866);
and UO_2985 (O_2985,N_49761,N_48046);
xor UO_2986 (O_2986,N_48594,N_49593);
or UO_2987 (O_2987,N_48790,N_48278);
xnor UO_2988 (O_2988,N_49455,N_48070);
and UO_2989 (O_2989,N_48666,N_48243);
nor UO_2990 (O_2990,N_49618,N_49910);
xnor UO_2991 (O_2991,N_49177,N_48715);
nor UO_2992 (O_2992,N_49355,N_49425);
or UO_2993 (O_2993,N_48530,N_49587);
nor UO_2994 (O_2994,N_49085,N_48042);
and UO_2995 (O_2995,N_49699,N_48500);
or UO_2996 (O_2996,N_48780,N_49659);
nand UO_2997 (O_2997,N_48886,N_48307);
nand UO_2998 (O_2998,N_48125,N_48621);
and UO_2999 (O_2999,N_49011,N_48292);
nor UO_3000 (O_3000,N_49031,N_48497);
and UO_3001 (O_3001,N_49522,N_48351);
or UO_3002 (O_3002,N_49390,N_49116);
xor UO_3003 (O_3003,N_49590,N_48068);
or UO_3004 (O_3004,N_48763,N_49686);
and UO_3005 (O_3005,N_48723,N_49652);
or UO_3006 (O_3006,N_49610,N_48243);
nand UO_3007 (O_3007,N_49323,N_48077);
nand UO_3008 (O_3008,N_49008,N_49152);
or UO_3009 (O_3009,N_49987,N_48502);
or UO_3010 (O_3010,N_48206,N_49136);
nor UO_3011 (O_3011,N_49825,N_49604);
and UO_3012 (O_3012,N_48214,N_49736);
nor UO_3013 (O_3013,N_49703,N_49652);
xor UO_3014 (O_3014,N_48537,N_48940);
nand UO_3015 (O_3015,N_48053,N_49221);
and UO_3016 (O_3016,N_48691,N_48835);
nand UO_3017 (O_3017,N_49848,N_49482);
or UO_3018 (O_3018,N_49391,N_48916);
and UO_3019 (O_3019,N_49224,N_48637);
or UO_3020 (O_3020,N_48802,N_48196);
nand UO_3021 (O_3021,N_49693,N_48025);
or UO_3022 (O_3022,N_48149,N_48226);
and UO_3023 (O_3023,N_49245,N_49192);
nor UO_3024 (O_3024,N_48973,N_49098);
xnor UO_3025 (O_3025,N_49925,N_49294);
xnor UO_3026 (O_3026,N_48308,N_49492);
and UO_3027 (O_3027,N_49857,N_48643);
nor UO_3028 (O_3028,N_49726,N_49632);
nor UO_3029 (O_3029,N_48098,N_48235);
or UO_3030 (O_3030,N_49237,N_49393);
or UO_3031 (O_3031,N_48846,N_48276);
nand UO_3032 (O_3032,N_48728,N_49023);
xor UO_3033 (O_3033,N_49762,N_49054);
xnor UO_3034 (O_3034,N_48243,N_48552);
and UO_3035 (O_3035,N_48234,N_48457);
nor UO_3036 (O_3036,N_49258,N_48089);
nor UO_3037 (O_3037,N_49167,N_48642);
xor UO_3038 (O_3038,N_49207,N_48076);
xnor UO_3039 (O_3039,N_49703,N_49523);
xor UO_3040 (O_3040,N_49104,N_49399);
or UO_3041 (O_3041,N_48648,N_48850);
nor UO_3042 (O_3042,N_49160,N_49555);
or UO_3043 (O_3043,N_49030,N_48313);
nor UO_3044 (O_3044,N_48275,N_48939);
nand UO_3045 (O_3045,N_48151,N_49996);
or UO_3046 (O_3046,N_48536,N_48029);
xor UO_3047 (O_3047,N_48402,N_48024);
nand UO_3048 (O_3048,N_48735,N_49387);
nand UO_3049 (O_3049,N_49000,N_49265);
nor UO_3050 (O_3050,N_48610,N_48398);
nor UO_3051 (O_3051,N_49907,N_49430);
and UO_3052 (O_3052,N_49953,N_48470);
xnor UO_3053 (O_3053,N_48935,N_48177);
nand UO_3054 (O_3054,N_49247,N_48954);
nand UO_3055 (O_3055,N_49778,N_48333);
nor UO_3056 (O_3056,N_48786,N_49306);
or UO_3057 (O_3057,N_49081,N_48482);
xor UO_3058 (O_3058,N_49297,N_48021);
nor UO_3059 (O_3059,N_49457,N_48857);
xnor UO_3060 (O_3060,N_49557,N_48714);
and UO_3061 (O_3061,N_49735,N_48243);
or UO_3062 (O_3062,N_48592,N_49632);
and UO_3063 (O_3063,N_49344,N_48884);
and UO_3064 (O_3064,N_48364,N_49668);
and UO_3065 (O_3065,N_49599,N_48443);
xor UO_3066 (O_3066,N_48529,N_48309);
xnor UO_3067 (O_3067,N_49569,N_48638);
nand UO_3068 (O_3068,N_48414,N_49760);
xor UO_3069 (O_3069,N_48044,N_49377);
or UO_3070 (O_3070,N_49617,N_48013);
or UO_3071 (O_3071,N_48372,N_48248);
nand UO_3072 (O_3072,N_49314,N_49019);
nor UO_3073 (O_3073,N_48915,N_49193);
nor UO_3074 (O_3074,N_49730,N_48454);
nand UO_3075 (O_3075,N_49832,N_48918);
and UO_3076 (O_3076,N_48650,N_49963);
nand UO_3077 (O_3077,N_48988,N_49668);
nand UO_3078 (O_3078,N_48331,N_49799);
xnor UO_3079 (O_3079,N_48072,N_48355);
or UO_3080 (O_3080,N_49170,N_48930);
xnor UO_3081 (O_3081,N_49915,N_49950);
and UO_3082 (O_3082,N_48840,N_48652);
nand UO_3083 (O_3083,N_49832,N_49824);
nor UO_3084 (O_3084,N_48262,N_48395);
xor UO_3085 (O_3085,N_48878,N_49506);
nand UO_3086 (O_3086,N_48204,N_48030);
nand UO_3087 (O_3087,N_49586,N_48882);
nor UO_3088 (O_3088,N_49879,N_48750);
xnor UO_3089 (O_3089,N_49416,N_49677);
nand UO_3090 (O_3090,N_49026,N_49647);
and UO_3091 (O_3091,N_49601,N_48377);
nor UO_3092 (O_3092,N_48102,N_48518);
or UO_3093 (O_3093,N_49053,N_48349);
or UO_3094 (O_3094,N_49886,N_49565);
nand UO_3095 (O_3095,N_48060,N_48916);
or UO_3096 (O_3096,N_49210,N_49055);
and UO_3097 (O_3097,N_49061,N_48037);
and UO_3098 (O_3098,N_48085,N_48049);
nor UO_3099 (O_3099,N_48099,N_49251);
or UO_3100 (O_3100,N_48573,N_49940);
xor UO_3101 (O_3101,N_49816,N_48450);
xor UO_3102 (O_3102,N_48593,N_49818);
nand UO_3103 (O_3103,N_49837,N_48215);
xor UO_3104 (O_3104,N_49394,N_48888);
and UO_3105 (O_3105,N_49354,N_49339);
xnor UO_3106 (O_3106,N_48809,N_49170);
and UO_3107 (O_3107,N_49010,N_49605);
nand UO_3108 (O_3108,N_49745,N_48878);
nand UO_3109 (O_3109,N_49167,N_49266);
nor UO_3110 (O_3110,N_48745,N_48717);
nand UO_3111 (O_3111,N_49908,N_48123);
and UO_3112 (O_3112,N_49814,N_48457);
nor UO_3113 (O_3113,N_49764,N_48834);
or UO_3114 (O_3114,N_49836,N_49108);
xor UO_3115 (O_3115,N_49925,N_49943);
nand UO_3116 (O_3116,N_49901,N_48167);
nand UO_3117 (O_3117,N_48961,N_48170);
nand UO_3118 (O_3118,N_49483,N_49922);
and UO_3119 (O_3119,N_48096,N_48204);
or UO_3120 (O_3120,N_48397,N_49359);
xor UO_3121 (O_3121,N_49688,N_48707);
nand UO_3122 (O_3122,N_48352,N_49824);
xnor UO_3123 (O_3123,N_48238,N_48745);
xnor UO_3124 (O_3124,N_48101,N_49525);
nor UO_3125 (O_3125,N_48131,N_49468);
xnor UO_3126 (O_3126,N_49168,N_49676);
xor UO_3127 (O_3127,N_48702,N_49481);
and UO_3128 (O_3128,N_49516,N_48536);
nand UO_3129 (O_3129,N_49029,N_49749);
xor UO_3130 (O_3130,N_49017,N_48784);
xor UO_3131 (O_3131,N_49784,N_49788);
nor UO_3132 (O_3132,N_48565,N_49055);
nor UO_3133 (O_3133,N_48232,N_48899);
xnor UO_3134 (O_3134,N_48251,N_48011);
or UO_3135 (O_3135,N_49205,N_48761);
and UO_3136 (O_3136,N_48426,N_49396);
nor UO_3137 (O_3137,N_49116,N_48421);
and UO_3138 (O_3138,N_49424,N_48314);
or UO_3139 (O_3139,N_49117,N_48565);
nor UO_3140 (O_3140,N_49508,N_48280);
nor UO_3141 (O_3141,N_48635,N_49841);
nand UO_3142 (O_3142,N_48208,N_49352);
xor UO_3143 (O_3143,N_48985,N_49260);
xnor UO_3144 (O_3144,N_48506,N_48722);
xor UO_3145 (O_3145,N_49709,N_48059);
nand UO_3146 (O_3146,N_48695,N_49413);
nor UO_3147 (O_3147,N_49662,N_49736);
nand UO_3148 (O_3148,N_49324,N_48643);
nand UO_3149 (O_3149,N_49442,N_49078);
xor UO_3150 (O_3150,N_48728,N_49140);
and UO_3151 (O_3151,N_48900,N_49812);
or UO_3152 (O_3152,N_49057,N_48427);
nand UO_3153 (O_3153,N_49417,N_48571);
nand UO_3154 (O_3154,N_49624,N_49685);
xnor UO_3155 (O_3155,N_49540,N_49172);
nor UO_3156 (O_3156,N_48768,N_48484);
xnor UO_3157 (O_3157,N_49212,N_48036);
nand UO_3158 (O_3158,N_48895,N_48147);
or UO_3159 (O_3159,N_49654,N_48813);
nor UO_3160 (O_3160,N_49465,N_48930);
nand UO_3161 (O_3161,N_48458,N_49244);
nor UO_3162 (O_3162,N_49421,N_49502);
or UO_3163 (O_3163,N_48267,N_49279);
and UO_3164 (O_3164,N_48797,N_48083);
nor UO_3165 (O_3165,N_48802,N_49965);
and UO_3166 (O_3166,N_48977,N_49927);
nand UO_3167 (O_3167,N_48969,N_49345);
or UO_3168 (O_3168,N_48768,N_48356);
or UO_3169 (O_3169,N_48582,N_49926);
nand UO_3170 (O_3170,N_49984,N_48219);
nor UO_3171 (O_3171,N_48264,N_49507);
nand UO_3172 (O_3172,N_49368,N_48976);
xor UO_3173 (O_3173,N_48656,N_48160);
nand UO_3174 (O_3174,N_49997,N_49800);
nor UO_3175 (O_3175,N_49666,N_48211);
and UO_3176 (O_3176,N_48658,N_48483);
xor UO_3177 (O_3177,N_49469,N_48036);
nand UO_3178 (O_3178,N_48862,N_48251);
xor UO_3179 (O_3179,N_49052,N_48764);
xor UO_3180 (O_3180,N_49469,N_48280);
and UO_3181 (O_3181,N_49037,N_49910);
or UO_3182 (O_3182,N_49484,N_49469);
nor UO_3183 (O_3183,N_48926,N_48810);
xor UO_3184 (O_3184,N_48521,N_49799);
nor UO_3185 (O_3185,N_49912,N_48900);
nand UO_3186 (O_3186,N_49485,N_48086);
xnor UO_3187 (O_3187,N_49947,N_49788);
nand UO_3188 (O_3188,N_48462,N_48135);
xnor UO_3189 (O_3189,N_48976,N_48787);
or UO_3190 (O_3190,N_48194,N_49543);
or UO_3191 (O_3191,N_48016,N_49555);
xor UO_3192 (O_3192,N_48704,N_49945);
xor UO_3193 (O_3193,N_49136,N_48338);
xor UO_3194 (O_3194,N_48528,N_49746);
nor UO_3195 (O_3195,N_48236,N_49007);
xnor UO_3196 (O_3196,N_48547,N_49696);
xnor UO_3197 (O_3197,N_48604,N_48456);
nor UO_3198 (O_3198,N_49489,N_49286);
xnor UO_3199 (O_3199,N_48047,N_48628);
xnor UO_3200 (O_3200,N_49329,N_48960);
xnor UO_3201 (O_3201,N_48604,N_49195);
nor UO_3202 (O_3202,N_49423,N_48473);
and UO_3203 (O_3203,N_48220,N_48964);
nand UO_3204 (O_3204,N_48472,N_48021);
nor UO_3205 (O_3205,N_48902,N_48589);
nand UO_3206 (O_3206,N_48113,N_48522);
xnor UO_3207 (O_3207,N_49255,N_49341);
xor UO_3208 (O_3208,N_49216,N_48793);
and UO_3209 (O_3209,N_48030,N_48710);
nand UO_3210 (O_3210,N_49256,N_48741);
nor UO_3211 (O_3211,N_49232,N_49141);
nand UO_3212 (O_3212,N_48386,N_49243);
and UO_3213 (O_3213,N_48595,N_49871);
nor UO_3214 (O_3214,N_48898,N_48163);
xnor UO_3215 (O_3215,N_49772,N_48959);
nand UO_3216 (O_3216,N_49915,N_49856);
and UO_3217 (O_3217,N_49317,N_49489);
or UO_3218 (O_3218,N_49451,N_49491);
nor UO_3219 (O_3219,N_49045,N_48561);
or UO_3220 (O_3220,N_48011,N_49758);
and UO_3221 (O_3221,N_48138,N_48083);
and UO_3222 (O_3222,N_49189,N_48263);
nor UO_3223 (O_3223,N_49754,N_49123);
xnor UO_3224 (O_3224,N_48175,N_48036);
xor UO_3225 (O_3225,N_49486,N_49766);
nand UO_3226 (O_3226,N_49332,N_48340);
or UO_3227 (O_3227,N_48175,N_48404);
and UO_3228 (O_3228,N_49438,N_48766);
xnor UO_3229 (O_3229,N_49450,N_49291);
and UO_3230 (O_3230,N_48478,N_49691);
nor UO_3231 (O_3231,N_49181,N_49591);
xor UO_3232 (O_3232,N_48716,N_49073);
and UO_3233 (O_3233,N_48204,N_49466);
and UO_3234 (O_3234,N_48684,N_48216);
nand UO_3235 (O_3235,N_49388,N_48222);
and UO_3236 (O_3236,N_49002,N_48610);
and UO_3237 (O_3237,N_48894,N_48852);
or UO_3238 (O_3238,N_49844,N_48488);
or UO_3239 (O_3239,N_48569,N_48244);
nor UO_3240 (O_3240,N_48961,N_49059);
nor UO_3241 (O_3241,N_49111,N_48607);
xnor UO_3242 (O_3242,N_48461,N_48227);
nand UO_3243 (O_3243,N_49770,N_48406);
nand UO_3244 (O_3244,N_49430,N_48709);
xor UO_3245 (O_3245,N_48184,N_48623);
xnor UO_3246 (O_3246,N_48684,N_49574);
xor UO_3247 (O_3247,N_49337,N_49187);
xor UO_3248 (O_3248,N_48881,N_48996);
nand UO_3249 (O_3249,N_49121,N_48240);
xnor UO_3250 (O_3250,N_49210,N_48110);
and UO_3251 (O_3251,N_49987,N_48535);
xnor UO_3252 (O_3252,N_48365,N_49800);
xnor UO_3253 (O_3253,N_49505,N_48394);
or UO_3254 (O_3254,N_48643,N_49637);
nor UO_3255 (O_3255,N_49788,N_48884);
xnor UO_3256 (O_3256,N_48435,N_48762);
xor UO_3257 (O_3257,N_48588,N_49681);
nand UO_3258 (O_3258,N_49715,N_49444);
nand UO_3259 (O_3259,N_49186,N_49064);
or UO_3260 (O_3260,N_48644,N_49430);
or UO_3261 (O_3261,N_48159,N_49668);
or UO_3262 (O_3262,N_49163,N_49615);
xnor UO_3263 (O_3263,N_48349,N_48284);
nand UO_3264 (O_3264,N_48988,N_49438);
nor UO_3265 (O_3265,N_49157,N_48843);
nand UO_3266 (O_3266,N_49544,N_48982);
nor UO_3267 (O_3267,N_48171,N_48049);
or UO_3268 (O_3268,N_48575,N_48541);
or UO_3269 (O_3269,N_48707,N_49766);
and UO_3270 (O_3270,N_49715,N_49711);
and UO_3271 (O_3271,N_49674,N_49681);
xor UO_3272 (O_3272,N_48382,N_49513);
nand UO_3273 (O_3273,N_49096,N_49148);
nand UO_3274 (O_3274,N_48656,N_49421);
and UO_3275 (O_3275,N_49248,N_48432);
xnor UO_3276 (O_3276,N_49440,N_49085);
nor UO_3277 (O_3277,N_49298,N_49731);
nand UO_3278 (O_3278,N_48672,N_48364);
and UO_3279 (O_3279,N_48052,N_49717);
or UO_3280 (O_3280,N_48146,N_48097);
and UO_3281 (O_3281,N_49725,N_48638);
nand UO_3282 (O_3282,N_49406,N_49710);
nor UO_3283 (O_3283,N_48753,N_48689);
xor UO_3284 (O_3284,N_49681,N_49334);
nor UO_3285 (O_3285,N_48779,N_49423);
nand UO_3286 (O_3286,N_49450,N_49598);
or UO_3287 (O_3287,N_49919,N_48868);
nand UO_3288 (O_3288,N_48793,N_49927);
nor UO_3289 (O_3289,N_48306,N_49478);
and UO_3290 (O_3290,N_48218,N_48473);
or UO_3291 (O_3291,N_49402,N_48247);
nor UO_3292 (O_3292,N_49641,N_49723);
nor UO_3293 (O_3293,N_48251,N_49795);
nand UO_3294 (O_3294,N_49235,N_48022);
or UO_3295 (O_3295,N_49821,N_49905);
nand UO_3296 (O_3296,N_48953,N_48256);
or UO_3297 (O_3297,N_48762,N_49184);
or UO_3298 (O_3298,N_49497,N_48330);
and UO_3299 (O_3299,N_49273,N_48471);
nor UO_3300 (O_3300,N_49255,N_48559);
nor UO_3301 (O_3301,N_49621,N_48849);
xor UO_3302 (O_3302,N_48676,N_49965);
xnor UO_3303 (O_3303,N_48877,N_49033);
and UO_3304 (O_3304,N_49632,N_48612);
nor UO_3305 (O_3305,N_49081,N_48162);
or UO_3306 (O_3306,N_48106,N_49047);
nor UO_3307 (O_3307,N_49065,N_49656);
xor UO_3308 (O_3308,N_49237,N_48165);
nor UO_3309 (O_3309,N_48622,N_49200);
nor UO_3310 (O_3310,N_48904,N_49718);
nand UO_3311 (O_3311,N_49860,N_49201);
nor UO_3312 (O_3312,N_49696,N_49898);
xor UO_3313 (O_3313,N_49642,N_48312);
nand UO_3314 (O_3314,N_48458,N_48398);
nor UO_3315 (O_3315,N_49203,N_48653);
and UO_3316 (O_3316,N_49095,N_48925);
xnor UO_3317 (O_3317,N_48879,N_48080);
and UO_3318 (O_3318,N_48961,N_49637);
nor UO_3319 (O_3319,N_48690,N_48524);
xor UO_3320 (O_3320,N_49534,N_48319);
and UO_3321 (O_3321,N_48521,N_48210);
nand UO_3322 (O_3322,N_48160,N_49551);
or UO_3323 (O_3323,N_48759,N_49662);
xor UO_3324 (O_3324,N_48020,N_48291);
nand UO_3325 (O_3325,N_49975,N_48444);
or UO_3326 (O_3326,N_49038,N_48294);
nor UO_3327 (O_3327,N_49174,N_48940);
xnor UO_3328 (O_3328,N_48687,N_48537);
nor UO_3329 (O_3329,N_48296,N_48538);
or UO_3330 (O_3330,N_48337,N_48230);
and UO_3331 (O_3331,N_49675,N_48708);
or UO_3332 (O_3332,N_49318,N_49393);
xnor UO_3333 (O_3333,N_48899,N_48588);
nand UO_3334 (O_3334,N_49766,N_49735);
or UO_3335 (O_3335,N_48813,N_48880);
and UO_3336 (O_3336,N_49333,N_49959);
and UO_3337 (O_3337,N_49012,N_48603);
or UO_3338 (O_3338,N_49487,N_48384);
nand UO_3339 (O_3339,N_48112,N_49718);
nand UO_3340 (O_3340,N_49006,N_49862);
nand UO_3341 (O_3341,N_49425,N_48744);
nor UO_3342 (O_3342,N_49834,N_48381);
nand UO_3343 (O_3343,N_49734,N_48349);
nor UO_3344 (O_3344,N_48149,N_49381);
nor UO_3345 (O_3345,N_48274,N_49407);
and UO_3346 (O_3346,N_48592,N_49529);
or UO_3347 (O_3347,N_49070,N_49193);
xor UO_3348 (O_3348,N_48225,N_49244);
and UO_3349 (O_3349,N_49617,N_48222);
xor UO_3350 (O_3350,N_48062,N_48504);
xor UO_3351 (O_3351,N_48354,N_49523);
nand UO_3352 (O_3352,N_48196,N_48959);
and UO_3353 (O_3353,N_48114,N_49722);
xor UO_3354 (O_3354,N_49652,N_49730);
nand UO_3355 (O_3355,N_49512,N_48677);
nor UO_3356 (O_3356,N_48578,N_48201);
xnor UO_3357 (O_3357,N_48851,N_48778);
nand UO_3358 (O_3358,N_49838,N_49107);
nand UO_3359 (O_3359,N_49062,N_48556);
and UO_3360 (O_3360,N_48029,N_49528);
xor UO_3361 (O_3361,N_49923,N_48242);
or UO_3362 (O_3362,N_48917,N_49168);
or UO_3363 (O_3363,N_49190,N_48321);
xor UO_3364 (O_3364,N_48587,N_49718);
nor UO_3365 (O_3365,N_49255,N_48428);
nand UO_3366 (O_3366,N_49539,N_48686);
nand UO_3367 (O_3367,N_49366,N_49280);
and UO_3368 (O_3368,N_49883,N_49615);
or UO_3369 (O_3369,N_49697,N_49899);
xnor UO_3370 (O_3370,N_49439,N_48450);
nor UO_3371 (O_3371,N_48944,N_49059);
or UO_3372 (O_3372,N_48182,N_48572);
and UO_3373 (O_3373,N_49432,N_48288);
or UO_3374 (O_3374,N_49482,N_49297);
nand UO_3375 (O_3375,N_48629,N_49239);
xor UO_3376 (O_3376,N_48714,N_48793);
or UO_3377 (O_3377,N_49245,N_48024);
xor UO_3378 (O_3378,N_48522,N_48208);
nand UO_3379 (O_3379,N_48643,N_48979);
xnor UO_3380 (O_3380,N_49156,N_48035);
or UO_3381 (O_3381,N_48764,N_49347);
nor UO_3382 (O_3382,N_49081,N_49505);
or UO_3383 (O_3383,N_48088,N_49740);
nor UO_3384 (O_3384,N_49498,N_48404);
nand UO_3385 (O_3385,N_49313,N_48441);
xor UO_3386 (O_3386,N_48555,N_48986);
or UO_3387 (O_3387,N_49334,N_48000);
xnor UO_3388 (O_3388,N_48007,N_48022);
and UO_3389 (O_3389,N_49890,N_48072);
or UO_3390 (O_3390,N_49151,N_48837);
and UO_3391 (O_3391,N_49351,N_48959);
or UO_3392 (O_3392,N_48621,N_49529);
or UO_3393 (O_3393,N_49398,N_48506);
nand UO_3394 (O_3394,N_49977,N_49224);
nand UO_3395 (O_3395,N_49917,N_48893);
xor UO_3396 (O_3396,N_49135,N_48600);
xor UO_3397 (O_3397,N_49434,N_49759);
nand UO_3398 (O_3398,N_49425,N_49812);
and UO_3399 (O_3399,N_48483,N_48365);
nor UO_3400 (O_3400,N_49554,N_49470);
nand UO_3401 (O_3401,N_48757,N_48382);
or UO_3402 (O_3402,N_48931,N_48613);
nand UO_3403 (O_3403,N_48102,N_48152);
xor UO_3404 (O_3404,N_48335,N_49132);
xor UO_3405 (O_3405,N_49621,N_48708);
and UO_3406 (O_3406,N_48264,N_49168);
nand UO_3407 (O_3407,N_49159,N_48753);
nand UO_3408 (O_3408,N_48943,N_49291);
and UO_3409 (O_3409,N_49813,N_49846);
nor UO_3410 (O_3410,N_49693,N_48484);
or UO_3411 (O_3411,N_49161,N_49274);
and UO_3412 (O_3412,N_49617,N_48577);
nand UO_3413 (O_3413,N_49270,N_48407);
xor UO_3414 (O_3414,N_49505,N_49135);
and UO_3415 (O_3415,N_49886,N_49523);
xor UO_3416 (O_3416,N_49919,N_49680);
xor UO_3417 (O_3417,N_48896,N_48311);
or UO_3418 (O_3418,N_48460,N_49867);
xor UO_3419 (O_3419,N_48769,N_49828);
or UO_3420 (O_3420,N_49935,N_48059);
and UO_3421 (O_3421,N_48598,N_49770);
xnor UO_3422 (O_3422,N_49675,N_49345);
nor UO_3423 (O_3423,N_48304,N_49905);
nand UO_3424 (O_3424,N_48170,N_48995);
xnor UO_3425 (O_3425,N_48320,N_48458);
or UO_3426 (O_3426,N_48966,N_48358);
or UO_3427 (O_3427,N_49886,N_49045);
or UO_3428 (O_3428,N_49022,N_49510);
xnor UO_3429 (O_3429,N_48126,N_48421);
nand UO_3430 (O_3430,N_48946,N_48348);
nand UO_3431 (O_3431,N_48845,N_49945);
nand UO_3432 (O_3432,N_48031,N_48579);
and UO_3433 (O_3433,N_49236,N_49321);
or UO_3434 (O_3434,N_49215,N_49120);
nor UO_3435 (O_3435,N_49402,N_49768);
nor UO_3436 (O_3436,N_48425,N_49194);
or UO_3437 (O_3437,N_49876,N_48014);
nand UO_3438 (O_3438,N_48126,N_49400);
and UO_3439 (O_3439,N_48427,N_49839);
and UO_3440 (O_3440,N_48503,N_49080);
and UO_3441 (O_3441,N_49942,N_48040);
or UO_3442 (O_3442,N_48724,N_48363);
or UO_3443 (O_3443,N_48521,N_49877);
and UO_3444 (O_3444,N_49027,N_48563);
xnor UO_3445 (O_3445,N_48752,N_49150);
and UO_3446 (O_3446,N_48028,N_48411);
and UO_3447 (O_3447,N_49623,N_49344);
and UO_3448 (O_3448,N_48707,N_48002);
and UO_3449 (O_3449,N_49283,N_49597);
xnor UO_3450 (O_3450,N_49170,N_48750);
or UO_3451 (O_3451,N_48443,N_48068);
nor UO_3452 (O_3452,N_49009,N_49873);
and UO_3453 (O_3453,N_48702,N_48800);
nand UO_3454 (O_3454,N_49556,N_48517);
and UO_3455 (O_3455,N_49061,N_49492);
nand UO_3456 (O_3456,N_48994,N_49269);
nand UO_3457 (O_3457,N_48149,N_48797);
nor UO_3458 (O_3458,N_49946,N_49954);
nor UO_3459 (O_3459,N_49373,N_48100);
nand UO_3460 (O_3460,N_48240,N_49601);
nand UO_3461 (O_3461,N_49866,N_49599);
xor UO_3462 (O_3462,N_49987,N_48458);
nand UO_3463 (O_3463,N_48952,N_48684);
and UO_3464 (O_3464,N_49380,N_49019);
nor UO_3465 (O_3465,N_48654,N_49749);
and UO_3466 (O_3466,N_49665,N_49809);
nor UO_3467 (O_3467,N_48403,N_48529);
and UO_3468 (O_3468,N_48606,N_48149);
and UO_3469 (O_3469,N_49711,N_48127);
nand UO_3470 (O_3470,N_48070,N_48009);
nand UO_3471 (O_3471,N_48407,N_48450);
or UO_3472 (O_3472,N_48522,N_48814);
and UO_3473 (O_3473,N_49962,N_48422);
nand UO_3474 (O_3474,N_48250,N_49250);
xor UO_3475 (O_3475,N_49044,N_49124);
xor UO_3476 (O_3476,N_49152,N_48384);
and UO_3477 (O_3477,N_49187,N_48187);
xnor UO_3478 (O_3478,N_49164,N_48098);
and UO_3479 (O_3479,N_49912,N_49076);
nor UO_3480 (O_3480,N_48311,N_48540);
nor UO_3481 (O_3481,N_48034,N_49225);
nor UO_3482 (O_3482,N_49122,N_48318);
xor UO_3483 (O_3483,N_48545,N_48218);
nor UO_3484 (O_3484,N_48666,N_48180);
nor UO_3485 (O_3485,N_48787,N_49924);
xnor UO_3486 (O_3486,N_49553,N_48817);
nor UO_3487 (O_3487,N_48964,N_48131);
nor UO_3488 (O_3488,N_49089,N_48381);
and UO_3489 (O_3489,N_48341,N_48072);
xor UO_3490 (O_3490,N_49513,N_48326);
xor UO_3491 (O_3491,N_49375,N_49767);
xor UO_3492 (O_3492,N_48566,N_49700);
and UO_3493 (O_3493,N_49499,N_48866);
nor UO_3494 (O_3494,N_48632,N_49740);
xor UO_3495 (O_3495,N_49942,N_48517);
nand UO_3496 (O_3496,N_48046,N_48039);
nand UO_3497 (O_3497,N_49101,N_48052);
nor UO_3498 (O_3498,N_48290,N_49059);
nor UO_3499 (O_3499,N_48112,N_49268);
nor UO_3500 (O_3500,N_49740,N_48576);
and UO_3501 (O_3501,N_49714,N_48584);
and UO_3502 (O_3502,N_49891,N_49468);
or UO_3503 (O_3503,N_49850,N_49355);
xnor UO_3504 (O_3504,N_48845,N_49221);
xor UO_3505 (O_3505,N_48038,N_49049);
xor UO_3506 (O_3506,N_48391,N_48059);
nand UO_3507 (O_3507,N_48359,N_48170);
or UO_3508 (O_3508,N_49817,N_48273);
and UO_3509 (O_3509,N_49889,N_48740);
xor UO_3510 (O_3510,N_48590,N_48584);
xor UO_3511 (O_3511,N_49265,N_48248);
nor UO_3512 (O_3512,N_49126,N_49293);
nor UO_3513 (O_3513,N_48579,N_49988);
nand UO_3514 (O_3514,N_48012,N_49844);
nor UO_3515 (O_3515,N_49809,N_49173);
nor UO_3516 (O_3516,N_48329,N_49001);
nor UO_3517 (O_3517,N_49616,N_49305);
nand UO_3518 (O_3518,N_48413,N_48430);
xnor UO_3519 (O_3519,N_49146,N_48944);
nand UO_3520 (O_3520,N_49454,N_48087);
or UO_3521 (O_3521,N_48240,N_48376);
and UO_3522 (O_3522,N_48005,N_49849);
xnor UO_3523 (O_3523,N_49808,N_49514);
nor UO_3524 (O_3524,N_48410,N_48953);
and UO_3525 (O_3525,N_48850,N_48263);
nand UO_3526 (O_3526,N_48730,N_48625);
nor UO_3527 (O_3527,N_49049,N_48608);
xnor UO_3528 (O_3528,N_49098,N_48802);
or UO_3529 (O_3529,N_49040,N_48709);
and UO_3530 (O_3530,N_49767,N_49060);
nand UO_3531 (O_3531,N_48183,N_49199);
xnor UO_3532 (O_3532,N_49970,N_48070);
nor UO_3533 (O_3533,N_48024,N_49892);
nand UO_3534 (O_3534,N_48036,N_48811);
or UO_3535 (O_3535,N_48689,N_48299);
nor UO_3536 (O_3536,N_49051,N_48810);
nand UO_3537 (O_3537,N_49344,N_49927);
nor UO_3538 (O_3538,N_48297,N_48640);
and UO_3539 (O_3539,N_49608,N_48788);
or UO_3540 (O_3540,N_48473,N_48540);
or UO_3541 (O_3541,N_49803,N_48373);
xnor UO_3542 (O_3542,N_48101,N_49572);
or UO_3543 (O_3543,N_48915,N_48174);
nand UO_3544 (O_3544,N_49007,N_49919);
nand UO_3545 (O_3545,N_48433,N_49125);
nor UO_3546 (O_3546,N_48611,N_49041);
or UO_3547 (O_3547,N_48196,N_48556);
or UO_3548 (O_3548,N_49348,N_48990);
or UO_3549 (O_3549,N_49971,N_48122);
nor UO_3550 (O_3550,N_49214,N_49369);
or UO_3551 (O_3551,N_49859,N_49676);
and UO_3552 (O_3552,N_49027,N_48628);
nand UO_3553 (O_3553,N_49229,N_48869);
nand UO_3554 (O_3554,N_49673,N_49729);
or UO_3555 (O_3555,N_49718,N_49376);
nor UO_3556 (O_3556,N_49132,N_49012);
and UO_3557 (O_3557,N_49682,N_48361);
nor UO_3558 (O_3558,N_48018,N_49760);
or UO_3559 (O_3559,N_48658,N_48724);
and UO_3560 (O_3560,N_49647,N_48437);
or UO_3561 (O_3561,N_49876,N_48779);
or UO_3562 (O_3562,N_49142,N_49614);
nand UO_3563 (O_3563,N_48725,N_48459);
xnor UO_3564 (O_3564,N_49793,N_49643);
and UO_3565 (O_3565,N_49047,N_48646);
nor UO_3566 (O_3566,N_48596,N_48371);
xor UO_3567 (O_3567,N_48698,N_49775);
xor UO_3568 (O_3568,N_48080,N_49547);
xor UO_3569 (O_3569,N_48854,N_48649);
or UO_3570 (O_3570,N_49178,N_49317);
nor UO_3571 (O_3571,N_49571,N_49298);
nand UO_3572 (O_3572,N_49064,N_49797);
xor UO_3573 (O_3573,N_48962,N_49792);
and UO_3574 (O_3574,N_48411,N_49280);
and UO_3575 (O_3575,N_49883,N_49689);
xnor UO_3576 (O_3576,N_49353,N_49382);
xnor UO_3577 (O_3577,N_49815,N_49226);
nand UO_3578 (O_3578,N_48241,N_49799);
nor UO_3579 (O_3579,N_48709,N_48405);
and UO_3580 (O_3580,N_49661,N_48000);
and UO_3581 (O_3581,N_48244,N_48895);
xor UO_3582 (O_3582,N_49540,N_49575);
nor UO_3583 (O_3583,N_49023,N_49722);
xor UO_3584 (O_3584,N_48740,N_49553);
or UO_3585 (O_3585,N_49049,N_49259);
or UO_3586 (O_3586,N_49637,N_48330);
and UO_3587 (O_3587,N_49610,N_48591);
nand UO_3588 (O_3588,N_49495,N_49274);
or UO_3589 (O_3589,N_49123,N_48397);
xor UO_3590 (O_3590,N_48607,N_49334);
nor UO_3591 (O_3591,N_48734,N_49681);
and UO_3592 (O_3592,N_49034,N_49864);
or UO_3593 (O_3593,N_49159,N_49098);
xnor UO_3594 (O_3594,N_48647,N_49144);
nand UO_3595 (O_3595,N_48651,N_49580);
and UO_3596 (O_3596,N_48996,N_49616);
nor UO_3597 (O_3597,N_49822,N_48813);
nor UO_3598 (O_3598,N_49259,N_49525);
nor UO_3599 (O_3599,N_49864,N_49851);
nor UO_3600 (O_3600,N_49300,N_49252);
or UO_3601 (O_3601,N_48924,N_48945);
nand UO_3602 (O_3602,N_49526,N_49135);
or UO_3603 (O_3603,N_48911,N_49596);
nand UO_3604 (O_3604,N_49540,N_48074);
xor UO_3605 (O_3605,N_49327,N_49844);
xnor UO_3606 (O_3606,N_48062,N_49885);
or UO_3607 (O_3607,N_49077,N_48617);
nor UO_3608 (O_3608,N_48360,N_48056);
nor UO_3609 (O_3609,N_49570,N_48536);
nand UO_3610 (O_3610,N_48112,N_49448);
and UO_3611 (O_3611,N_49349,N_49508);
and UO_3612 (O_3612,N_48060,N_49404);
nand UO_3613 (O_3613,N_49076,N_48294);
or UO_3614 (O_3614,N_49106,N_49936);
xnor UO_3615 (O_3615,N_48864,N_49389);
and UO_3616 (O_3616,N_49599,N_49358);
or UO_3617 (O_3617,N_48747,N_49541);
and UO_3618 (O_3618,N_49578,N_49710);
nand UO_3619 (O_3619,N_48506,N_48604);
xor UO_3620 (O_3620,N_48192,N_49299);
nand UO_3621 (O_3621,N_49535,N_49442);
nand UO_3622 (O_3622,N_49566,N_48295);
nor UO_3623 (O_3623,N_48944,N_48505);
nand UO_3624 (O_3624,N_49640,N_49975);
nor UO_3625 (O_3625,N_49854,N_48511);
and UO_3626 (O_3626,N_48478,N_49028);
nand UO_3627 (O_3627,N_49126,N_48105);
xor UO_3628 (O_3628,N_49569,N_48365);
xnor UO_3629 (O_3629,N_49186,N_48016);
or UO_3630 (O_3630,N_49295,N_49475);
and UO_3631 (O_3631,N_48509,N_49766);
or UO_3632 (O_3632,N_49509,N_49932);
nand UO_3633 (O_3633,N_48110,N_49089);
and UO_3634 (O_3634,N_49224,N_48707);
and UO_3635 (O_3635,N_48825,N_49731);
xnor UO_3636 (O_3636,N_48723,N_49300);
nand UO_3637 (O_3637,N_49368,N_49534);
and UO_3638 (O_3638,N_48501,N_49298);
and UO_3639 (O_3639,N_48748,N_48235);
xnor UO_3640 (O_3640,N_48591,N_48162);
and UO_3641 (O_3641,N_48834,N_49097);
xor UO_3642 (O_3642,N_49244,N_49232);
xor UO_3643 (O_3643,N_49439,N_49677);
nand UO_3644 (O_3644,N_48728,N_48408);
nor UO_3645 (O_3645,N_49427,N_48350);
nor UO_3646 (O_3646,N_49102,N_49228);
nand UO_3647 (O_3647,N_49737,N_49552);
or UO_3648 (O_3648,N_48698,N_48998);
nor UO_3649 (O_3649,N_49347,N_49397);
or UO_3650 (O_3650,N_49443,N_49264);
nor UO_3651 (O_3651,N_49161,N_48611);
and UO_3652 (O_3652,N_48181,N_48146);
or UO_3653 (O_3653,N_49959,N_48227);
xnor UO_3654 (O_3654,N_48576,N_49425);
and UO_3655 (O_3655,N_49722,N_49334);
nand UO_3656 (O_3656,N_49852,N_49698);
nor UO_3657 (O_3657,N_49109,N_48433);
xor UO_3658 (O_3658,N_49388,N_48813);
xnor UO_3659 (O_3659,N_48140,N_49416);
or UO_3660 (O_3660,N_48695,N_49189);
xnor UO_3661 (O_3661,N_49979,N_49159);
nor UO_3662 (O_3662,N_48685,N_48765);
xnor UO_3663 (O_3663,N_49868,N_48224);
or UO_3664 (O_3664,N_49327,N_49211);
xor UO_3665 (O_3665,N_49334,N_49630);
xor UO_3666 (O_3666,N_49895,N_49077);
nor UO_3667 (O_3667,N_48739,N_48292);
and UO_3668 (O_3668,N_49841,N_48674);
nand UO_3669 (O_3669,N_49447,N_49224);
xor UO_3670 (O_3670,N_48907,N_49608);
and UO_3671 (O_3671,N_48217,N_48863);
or UO_3672 (O_3672,N_48488,N_48793);
xnor UO_3673 (O_3673,N_49660,N_48665);
nand UO_3674 (O_3674,N_48294,N_48627);
xor UO_3675 (O_3675,N_49961,N_48924);
nand UO_3676 (O_3676,N_49075,N_49959);
and UO_3677 (O_3677,N_49966,N_48803);
xnor UO_3678 (O_3678,N_48888,N_49670);
or UO_3679 (O_3679,N_48392,N_49848);
or UO_3680 (O_3680,N_48501,N_48201);
xnor UO_3681 (O_3681,N_48766,N_49813);
xor UO_3682 (O_3682,N_48823,N_48778);
nor UO_3683 (O_3683,N_49943,N_49217);
and UO_3684 (O_3684,N_49016,N_49439);
xor UO_3685 (O_3685,N_49209,N_49705);
xnor UO_3686 (O_3686,N_48151,N_49789);
or UO_3687 (O_3687,N_48391,N_49524);
or UO_3688 (O_3688,N_48079,N_49265);
and UO_3689 (O_3689,N_48428,N_49863);
nand UO_3690 (O_3690,N_49299,N_49910);
nand UO_3691 (O_3691,N_49955,N_48126);
nor UO_3692 (O_3692,N_49535,N_48290);
or UO_3693 (O_3693,N_49957,N_49250);
and UO_3694 (O_3694,N_49974,N_48509);
nand UO_3695 (O_3695,N_48847,N_49081);
or UO_3696 (O_3696,N_49809,N_49292);
or UO_3697 (O_3697,N_49763,N_48644);
nand UO_3698 (O_3698,N_48089,N_49093);
nand UO_3699 (O_3699,N_48869,N_49765);
xnor UO_3700 (O_3700,N_49694,N_48773);
and UO_3701 (O_3701,N_49021,N_49148);
and UO_3702 (O_3702,N_49742,N_49849);
nor UO_3703 (O_3703,N_48076,N_48520);
nand UO_3704 (O_3704,N_49327,N_49613);
or UO_3705 (O_3705,N_48785,N_49717);
xor UO_3706 (O_3706,N_49348,N_49311);
xor UO_3707 (O_3707,N_48246,N_49804);
or UO_3708 (O_3708,N_49892,N_49956);
or UO_3709 (O_3709,N_49199,N_48004);
nor UO_3710 (O_3710,N_48862,N_49234);
or UO_3711 (O_3711,N_48652,N_49026);
nand UO_3712 (O_3712,N_49571,N_49695);
nor UO_3713 (O_3713,N_48639,N_48485);
xor UO_3714 (O_3714,N_48171,N_48528);
or UO_3715 (O_3715,N_49396,N_49275);
nand UO_3716 (O_3716,N_48331,N_49529);
xor UO_3717 (O_3717,N_48798,N_49303);
xnor UO_3718 (O_3718,N_48198,N_48041);
nand UO_3719 (O_3719,N_48712,N_49112);
and UO_3720 (O_3720,N_48473,N_48037);
nand UO_3721 (O_3721,N_48863,N_49420);
or UO_3722 (O_3722,N_48724,N_48504);
or UO_3723 (O_3723,N_48586,N_49550);
nand UO_3724 (O_3724,N_49210,N_49379);
or UO_3725 (O_3725,N_49892,N_48210);
or UO_3726 (O_3726,N_48174,N_48144);
xnor UO_3727 (O_3727,N_48761,N_49523);
xnor UO_3728 (O_3728,N_49843,N_49712);
nor UO_3729 (O_3729,N_49919,N_48015);
nand UO_3730 (O_3730,N_49710,N_48308);
and UO_3731 (O_3731,N_48148,N_48596);
xnor UO_3732 (O_3732,N_49133,N_48009);
nand UO_3733 (O_3733,N_48988,N_49612);
xnor UO_3734 (O_3734,N_48577,N_49964);
or UO_3735 (O_3735,N_49148,N_48114);
or UO_3736 (O_3736,N_49245,N_48485);
xnor UO_3737 (O_3737,N_49468,N_48659);
or UO_3738 (O_3738,N_48849,N_48923);
nor UO_3739 (O_3739,N_48442,N_49100);
nand UO_3740 (O_3740,N_48486,N_49744);
or UO_3741 (O_3741,N_49954,N_49698);
nand UO_3742 (O_3742,N_48858,N_49520);
nand UO_3743 (O_3743,N_48435,N_48240);
and UO_3744 (O_3744,N_48929,N_49661);
nand UO_3745 (O_3745,N_48772,N_49755);
and UO_3746 (O_3746,N_49918,N_48187);
and UO_3747 (O_3747,N_49078,N_49372);
xnor UO_3748 (O_3748,N_48302,N_48037);
nor UO_3749 (O_3749,N_49281,N_49344);
and UO_3750 (O_3750,N_48904,N_49864);
and UO_3751 (O_3751,N_49428,N_49409);
and UO_3752 (O_3752,N_48202,N_49469);
or UO_3753 (O_3753,N_48681,N_49159);
xor UO_3754 (O_3754,N_49201,N_49240);
nand UO_3755 (O_3755,N_49604,N_48939);
nor UO_3756 (O_3756,N_49406,N_48366);
nor UO_3757 (O_3757,N_48236,N_48973);
or UO_3758 (O_3758,N_48878,N_49299);
and UO_3759 (O_3759,N_48610,N_49530);
and UO_3760 (O_3760,N_48553,N_49556);
nand UO_3761 (O_3761,N_49809,N_49356);
or UO_3762 (O_3762,N_48783,N_48963);
or UO_3763 (O_3763,N_49901,N_48707);
nand UO_3764 (O_3764,N_48575,N_49341);
xor UO_3765 (O_3765,N_49744,N_48876);
nand UO_3766 (O_3766,N_49771,N_49825);
or UO_3767 (O_3767,N_48152,N_48575);
and UO_3768 (O_3768,N_48199,N_48063);
and UO_3769 (O_3769,N_48006,N_49413);
or UO_3770 (O_3770,N_48130,N_49157);
nand UO_3771 (O_3771,N_49698,N_49607);
xor UO_3772 (O_3772,N_49944,N_49159);
nand UO_3773 (O_3773,N_48777,N_48381);
and UO_3774 (O_3774,N_49378,N_48863);
xor UO_3775 (O_3775,N_48349,N_49526);
nor UO_3776 (O_3776,N_49604,N_49435);
and UO_3777 (O_3777,N_49433,N_49529);
or UO_3778 (O_3778,N_48710,N_48472);
nand UO_3779 (O_3779,N_48335,N_48221);
nor UO_3780 (O_3780,N_49690,N_48229);
xnor UO_3781 (O_3781,N_48823,N_48473);
nand UO_3782 (O_3782,N_49211,N_48696);
nand UO_3783 (O_3783,N_49197,N_48236);
nand UO_3784 (O_3784,N_49256,N_49823);
xor UO_3785 (O_3785,N_48562,N_49609);
nand UO_3786 (O_3786,N_49001,N_49806);
and UO_3787 (O_3787,N_49607,N_48163);
xor UO_3788 (O_3788,N_48443,N_48859);
or UO_3789 (O_3789,N_49671,N_48099);
and UO_3790 (O_3790,N_49712,N_49582);
nand UO_3791 (O_3791,N_49810,N_49177);
or UO_3792 (O_3792,N_49454,N_48443);
nand UO_3793 (O_3793,N_48777,N_49246);
and UO_3794 (O_3794,N_49633,N_48473);
nor UO_3795 (O_3795,N_48147,N_48660);
and UO_3796 (O_3796,N_49613,N_48022);
or UO_3797 (O_3797,N_49488,N_49292);
nand UO_3798 (O_3798,N_48271,N_49055);
or UO_3799 (O_3799,N_48377,N_49425);
and UO_3800 (O_3800,N_48794,N_49608);
nor UO_3801 (O_3801,N_48401,N_48459);
and UO_3802 (O_3802,N_48850,N_48413);
xnor UO_3803 (O_3803,N_49153,N_48650);
and UO_3804 (O_3804,N_48570,N_48284);
nor UO_3805 (O_3805,N_48349,N_48189);
xnor UO_3806 (O_3806,N_49845,N_48107);
xnor UO_3807 (O_3807,N_49888,N_49814);
xor UO_3808 (O_3808,N_48121,N_49618);
xor UO_3809 (O_3809,N_49041,N_48379);
or UO_3810 (O_3810,N_48349,N_48507);
or UO_3811 (O_3811,N_48457,N_49670);
nor UO_3812 (O_3812,N_49948,N_48238);
nand UO_3813 (O_3813,N_48592,N_48187);
or UO_3814 (O_3814,N_49425,N_48955);
and UO_3815 (O_3815,N_48049,N_48154);
or UO_3816 (O_3816,N_49948,N_49221);
or UO_3817 (O_3817,N_48926,N_49699);
or UO_3818 (O_3818,N_49919,N_49958);
nand UO_3819 (O_3819,N_49522,N_49257);
or UO_3820 (O_3820,N_49722,N_48749);
and UO_3821 (O_3821,N_48442,N_48821);
or UO_3822 (O_3822,N_49077,N_48455);
nand UO_3823 (O_3823,N_48268,N_48151);
or UO_3824 (O_3824,N_49464,N_49098);
xor UO_3825 (O_3825,N_49278,N_49755);
nand UO_3826 (O_3826,N_49638,N_48963);
nand UO_3827 (O_3827,N_48826,N_48510);
and UO_3828 (O_3828,N_48046,N_48852);
or UO_3829 (O_3829,N_48003,N_49542);
xnor UO_3830 (O_3830,N_48363,N_48474);
xnor UO_3831 (O_3831,N_48982,N_49886);
nor UO_3832 (O_3832,N_49646,N_49973);
and UO_3833 (O_3833,N_49274,N_49617);
xor UO_3834 (O_3834,N_49528,N_49233);
and UO_3835 (O_3835,N_48083,N_48934);
nor UO_3836 (O_3836,N_48099,N_48354);
nor UO_3837 (O_3837,N_48829,N_49564);
or UO_3838 (O_3838,N_49389,N_49874);
or UO_3839 (O_3839,N_48586,N_49108);
nand UO_3840 (O_3840,N_48538,N_49110);
xor UO_3841 (O_3841,N_49415,N_49864);
or UO_3842 (O_3842,N_49945,N_49730);
xor UO_3843 (O_3843,N_48660,N_49208);
xnor UO_3844 (O_3844,N_48168,N_49130);
xor UO_3845 (O_3845,N_48546,N_49957);
or UO_3846 (O_3846,N_48652,N_48623);
and UO_3847 (O_3847,N_48461,N_48099);
nor UO_3848 (O_3848,N_48536,N_48366);
or UO_3849 (O_3849,N_49852,N_48429);
or UO_3850 (O_3850,N_48557,N_48158);
and UO_3851 (O_3851,N_48660,N_48231);
xor UO_3852 (O_3852,N_49555,N_48472);
nor UO_3853 (O_3853,N_48887,N_49197);
or UO_3854 (O_3854,N_48834,N_49266);
nor UO_3855 (O_3855,N_48417,N_49734);
and UO_3856 (O_3856,N_48934,N_48038);
nor UO_3857 (O_3857,N_49998,N_49371);
xor UO_3858 (O_3858,N_48694,N_49348);
nor UO_3859 (O_3859,N_49214,N_48888);
nor UO_3860 (O_3860,N_48670,N_48666);
nand UO_3861 (O_3861,N_49496,N_49601);
nor UO_3862 (O_3862,N_49191,N_48350);
xnor UO_3863 (O_3863,N_48826,N_48910);
and UO_3864 (O_3864,N_48595,N_48278);
xnor UO_3865 (O_3865,N_49726,N_49310);
nand UO_3866 (O_3866,N_49960,N_48892);
xor UO_3867 (O_3867,N_49669,N_49358);
and UO_3868 (O_3868,N_48663,N_49964);
nor UO_3869 (O_3869,N_48465,N_49260);
xnor UO_3870 (O_3870,N_48597,N_49123);
or UO_3871 (O_3871,N_48325,N_49700);
nor UO_3872 (O_3872,N_48078,N_48375);
xor UO_3873 (O_3873,N_49903,N_49849);
and UO_3874 (O_3874,N_48955,N_48250);
nand UO_3875 (O_3875,N_48949,N_49352);
and UO_3876 (O_3876,N_49163,N_48910);
or UO_3877 (O_3877,N_49902,N_48050);
or UO_3878 (O_3878,N_49058,N_49236);
or UO_3879 (O_3879,N_49259,N_48506);
or UO_3880 (O_3880,N_48180,N_48324);
or UO_3881 (O_3881,N_48080,N_49709);
and UO_3882 (O_3882,N_49067,N_48936);
nand UO_3883 (O_3883,N_48165,N_49718);
and UO_3884 (O_3884,N_48316,N_49192);
and UO_3885 (O_3885,N_49000,N_49297);
or UO_3886 (O_3886,N_48228,N_48523);
nor UO_3887 (O_3887,N_48738,N_48079);
xor UO_3888 (O_3888,N_49157,N_49160);
or UO_3889 (O_3889,N_49475,N_48136);
or UO_3890 (O_3890,N_48923,N_48367);
nor UO_3891 (O_3891,N_48721,N_49497);
and UO_3892 (O_3892,N_48894,N_49062);
and UO_3893 (O_3893,N_49077,N_49291);
nand UO_3894 (O_3894,N_49136,N_49430);
or UO_3895 (O_3895,N_48388,N_49991);
xor UO_3896 (O_3896,N_49739,N_49521);
or UO_3897 (O_3897,N_49339,N_48695);
nor UO_3898 (O_3898,N_49046,N_48343);
nor UO_3899 (O_3899,N_49637,N_48494);
xor UO_3900 (O_3900,N_49719,N_48391);
or UO_3901 (O_3901,N_48688,N_48871);
nand UO_3902 (O_3902,N_48129,N_48150);
or UO_3903 (O_3903,N_49351,N_49756);
and UO_3904 (O_3904,N_48290,N_48063);
and UO_3905 (O_3905,N_49639,N_49850);
or UO_3906 (O_3906,N_48520,N_49453);
or UO_3907 (O_3907,N_49703,N_48244);
nand UO_3908 (O_3908,N_49278,N_48098);
xor UO_3909 (O_3909,N_48367,N_48601);
xor UO_3910 (O_3910,N_49115,N_48394);
or UO_3911 (O_3911,N_48504,N_48077);
xor UO_3912 (O_3912,N_49299,N_49781);
xor UO_3913 (O_3913,N_49291,N_48865);
and UO_3914 (O_3914,N_49009,N_49214);
nor UO_3915 (O_3915,N_49125,N_48731);
and UO_3916 (O_3916,N_49799,N_49506);
and UO_3917 (O_3917,N_48167,N_49622);
nor UO_3918 (O_3918,N_48414,N_48023);
or UO_3919 (O_3919,N_48861,N_49967);
nor UO_3920 (O_3920,N_48230,N_49763);
or UO_3921 (O_3921,N_49119,N_49450);
and UO_3922 (O_3922,N_49305,N_48459);
and UO_3923 (O_3923,N_49276,N_49713);
or UO_3924 (O_3924,N_49304,N_49415);
nand UO_3925 (O_3925,N_48817,N_49227);
xnor UO_3926 (O_3926,N_48946,N_48421);
nand UO_3927 (O_3927,N_48817,N_49733);
xor UO_3928 (O_3928,N_49979,N_48325);
nand UO_3929 (O_3929,N_48364,N_49360);
nor UO_3930 (O_3930,N_48926,N_49195);
and UO_3931 (O_3931,N_49828,N_49567);
nor UO_3932 (O_3932,N_48300,N_49113);
nand UO_3933 (O_3933,N_49605,N_48075);
xor UO_3934 (O_3934,N_49960,N_49114);
and UO_3935 (O_3935,N_48164,N_49837);
and UO_3936 (O_3936,N_49027,N_48574);
nor UO_3937 (O_3937,N_49721,N_49449);
nor UO_3938 (O_3938,N_49292,N_49686);
nand UO_3939 (O_3939,N_48547,N_48426);
or UO_3940 (O_3940,N_49931,N_49151);
and UO_3941 (O_3941,N_49880,N_48567);
or UO_3942 (O_3942,N_48638,N_49909);
xor UO_3943 (O_3943,N_48973,N_49093);
xor UO_3944 (O_3944,N_49451,N_48915);
xnor UO_3945 (O_3945,N_48030,N_48398);
and UO_3946 (O_3946,N_49341,N_48866);
nor UO_3947 (O_3947,N_49618,N_49408);
and UO_3948 (O_3948,N_48998,N_49308);
or UO_3949 (O_3949,N_48793,N_48346);
nor UO_3950 (O_3950,N_49192,N_49090);
xnor UO_3951 (O_3951,N_48622,N_48865);
and UO_3952 (O_3952,N_49887,N_48418);
nor UO_3953 (O_3953,N_48963,N_49685);
xor UO_3954 (O_3954,N_48671,N_48965);
xor UO_3955 (O_3955,N_49941,N_48398);
or UO_3956 (O_3956,N_49489,N_49471);
and UO_3957 (O_3957,N_48698,N_49470);
xnor UO_3958 (O_3958,N_48579,N_48639);
nand UO_3959 (O_3959,N_48262,N_48188);
or UO_3960 (O_3960,N_48002,N_49428);
nor UO_3961 (O_3961,N_48358,N_48980);
nor UO_3962 (O_3962,N_48556,N_49561);
nand UO_3963 (O_3963,N_49150,N_48540);
nor UO_3964 (O_3964,N_48822,N_48792);
xnor UO_3965 (O_3965,N_48513,N_49662);
and UO_3966 (O_3966,N_49627,N_48746);
nor UO_3967 (O_3967,N_49649,N_48462);
or UO_3968 (O_3968,N_48643,N_48682);
or UO_3969 (O_3969,N_49313,N_49760);
or UO_3970 (O_3970,N_49687,N_49353);
nor UO_3971 (O_3971,N_48141,N_48122);
xnor UO_3972 (O_3972,N_49968,N_49358);
xor UO_3973 (O_3973,N_48794,N_49453);
xnor UO_3974 (O_3974,N_48606,N_48366);
or UO_3975 (O_3975,N_48728,N_48041);
xnor UO_3976 (O_3976,N_48433,N_48934);
xnor UO_3977 (O_3977,N_49106,N_48248);
or UO_3978 (O_3978,N_48024,N_49385);
and UO_3979 (O_3979,N_48753,N_49847);
nor UO_3980 (O_3980,N_48530,N_48889);
or UO_3981 (O_3981,N_48567,N_48420);
and UO_3982 (O_3982,N_49665,N_49483);
nand UO_3983 (O_3983,N_49005,N_49003);
nand UO_3984 (O_3984,N_48713,N_49481);
and UO_3985 (O_3985,N_48008,N_49315);
nand UO_3986 (O_3986,N_49174,N_48608);
nand UO_3987 (O_3987,N_49812,N_48427);
xnor UO_3988 (O_3988,N_49872,N_48458);
xor UO_3989 (O_3989,N_49164,N_48723);
xor UO_3990 (O_3990,N_48107,N_48933);
nor UO_3991 (O_3991,N_49429,N_49838);
and UO_3992 (O_3992,N_48348,N_48305);
nor UO_3993 (O_3993,N_49203,N_48100);
xor UO_3994 (O_3994,N_49669,N_48750);
nor UO_3995 (O_3995,N_48986,N_49318);
xnor UO_3996 (O_3996,N_49634,N_48231);
or UO_3997 (O_3997,N_49923,N_49297);
or UO_3998 (O_3998,N_48335,N_49098);
or UO_3999 (O_3999,N_49824,N_48796);
nor UO_4000 (O_4000,N_48939,N_48582);
nor UO_4001 (O_4001,N_49321,N_48774);
or UO_4002 (O_4002,N_49673,N_48750);
nor UO_4003 (O_4003,N_48949,N_48195);
or UO_4004 (O_4004,N_49357,N_49206);
or UO_4005 (O_4005,N_48348,N_48088);
or UO_4006 (O_4006,N_49770,N_48559);
nor UO_4007 (O_4007,N_49074,N_48129);
or UO_4008 (O_4008,N_48985,N_49099);
xnor UO_4009 (O_4009,N_48215,N_49808);
nand UO_4010 (O_4010,N_49554,N_48721);
or UO_4011 (O_4011,N_49346,N_49288);
nand UO_4012 (O_4012,N_49335,N_49425);
and UO_4013 (O_4013,N_49787,N_49738);
nand UO_4014 (O_4014,N_49438,N_48239);
and UO_4015 (O_4015,N_49011,N_49199);
and UO_4016 (O_4016,N_48133,N_49612);
and UO_4017 (O_4017,N_49376,N_48259);
nand UO_4018 (O_4018,N_48492,N_48235);
or UO_4019 (O_4019,N_48456,N_48832);
xor UO_4020 (O_4020,N_48000,N_48648);
nand UO_4021 (O_4021,N_48074,N_48932);
xor UO_4022 (O_4022,N_49961,N_48358);
and UO_4023 (O_4023,N_49719,N_48098);
and UO_4024 (O_4024,N_49751,N_49498);
or UO_4025 (O_4025,N_49048,N_49513);
xor UO_4026 (O_4026,N_48154,N_48388);
or UO_4027 (O_4027,N_49894,N_48481);
and UO_4028 (O_4028,N_49528,N_49022);
nand UO_4029 (O_4029,N_49607,N_48240);
xnor UO_4030 (O_4030,N_48975,N_48205);
or UO_4031 (O_4031,N_48942,N_48675);
nand UO_4032 (O_4032,N_48006,N_49300);
xor UO_4033 (O_4033,N_48461,N_48767);
nor UO_4034 (O_4034,N_49649,N_48731);
nand UO_4035 (O_4035,N_49316,N_48556);
and UO_4036 (O_4036,N_48853,N_48780);
and UO_4037 (O_4037,N_49106,N_49105);
nand UO_4038 (O_4038,N_48769,N_48623);
and UO_4039 (O_4039,N_48524,N_49151);
and UO_4040 (O_4040,N_48352,N_49202);
xor UO_4041 (O_4041,N_48577,N_49313);
nor UO_4042 (O_4042,N_49702,N_48030);
xnor UO_4043 (O_4043,N_49273,N_49298);
nand UO_4044 (O_4044,N_48010,N_49072);
and UO_4045 (O_4045,N_49582,N_49207);
and UO_4046 (O_4046,N_48168,N_49241);
and UO_4047 (O_4047,N_49269,N_48036);
and UO_4048 (O_4048,N_49141,N_48762);
and UO_4049 (O_4049,N_49703,N_48519);
nor UO_4050 (O_4050,N_49617,N_48630);
nand UO_4051 (O_4051,N_48455,N_48386);
nand UO_4052 (O_4052,N_49698,N_49901);
xnor UO_4053 (O_4053,N_48622,N_49923);
or UO_4054 (O_4054,N_48038,N_48194);
nand UO_4055 (O_4055,N_49314,N_49547);
nand UO_4056 (O_4056,N_48715,N_49785);
nor UO_4057 (O_4057,N_48799,N_48914);
and UO_4058 (O_4058,N_48725,N_49842);
or UO_4059 (O_4059,N_49249,N_49715);
or UO_4060 (O_4060,N_49784,N_49411);
nand UO_4061 (O_4061,N_48472,N_49658);
nand UO_4062 (O_4062,N_49538,N_49918);
and UO_4063 (O_4063,N_49143,N_48343);
nand UO_4064 (O_4064,N_48861,N_48994);
nand UO_4065 (O_4065,N_48619,N_49319);
nand UO_4066 (O_4066,N_49256,N_49673);
or UO_4067 (O_4067,N_48279,N_49227);
and UO_4068 (O_4068,N_48008,N_48456);
xor UO_4069 (O_4069,N_48178,N_49832);
or UO_4070 (O_4070,N_48179,N_49629);
or UO_4071 (O_4071,N_49938,N_49189);
nor UO_4072 (O_4072,N_49093,N_49316);
xor UO_4073 (O_4073,N_49046,N_48095);
and UO_4074 (O_4074,N_48592,N_49665);
or UO_4075 (O_4075,N_48787,N_49138);
xnor UO_4076 (O_4076,N_48421,N_49056);
xor UO_4077 (O_4077,N_48138,N_49058);
nand UO_4078 (O_4078,N_48214,N_48049);
nor UO_4079 (O_4079,N_48299,N_48672);
or UO_4080 (O_4080,N_49065,N_49149);
and UO_4081 (O_4081,N_48092,N_49518);
nor UO_4082 (O_4082,N_48296,N_49563);
and UO_4083 (O_4083,N_48582,N_48867);
nor UO_4084 (O_4084,N_49190,N_48551);
or UO_4085 (O_4085,N_49867,N_49411);
xnor UO_4086 (O_4086,N_49326,N_49104);
and UO_4087 (O_4087,N_48220,N_49700);
nor UO_4088 (O_4088,N_49025,N_48664);
xor UO_4089 (O_4089,N_48593,N_48722);
or UO_4090 (O_4090,N_48678,N_49335);
nand UO_4091 (O_4091,N_48947,N_49253);
or UO_4092 (O_4092,N_49037,N_49122);
nor UO_4093 (O_4093,N_48615,N_49220);
xnor UO_4094 (O_4094,N_49870,N_49899);
xnor UO_4095 (O_4095,N_48516,N_49165);
and UO_4096 (O_4096,N_48370,N_49148);
nor UO_4097 (O_4097,N_48432,N_49483);
and UO_4098 (O_4098,N_48897,N_49121);
nand UO_4099 (O_4099,N_49124,N_49507);
xor UO_4100 (O_4100,N_48104,N_48955);
nand UO_4101 (O_4101,N_48385,N_49744);
xor UO_4102 (O_4102,N_48425,N_48477);
and UO_4103 (O_4103,N_49458,N_48859);
nand UO_4104 (O_4104,N_48782,N_48670);
or UO_4105 (O_4105,N_48164,N_49823);
xor UO_4106 (O_4106,N_49954,N_49667);
xnor UO_4107 (O_4107,N_48586,N_48124);
nand UO_4108 (O_4108,N_48782,N_48983);
and UO_4109 (O_4109,N_48366,N_49283);
xnor UO_4110 (O_4110,N_48727,N_49348);
nor UO_4111 (O_4111,N_49469,N_48175);
or UO_4112 (O_4112,N_49713,N_48016);
and UO_4113 (O_4113,N_49010,N_48167);
nor UO_4114 (O_4114,N_48021,N_48913);
nand UO_4115 (O_4115,N_49733,N_49638);
nor UO_4116 (O_4116,N_49200,N_48520);
or UO_4117 (O_4117,N_49295,N_49370);
nand UO_4118 (O_4118,N_49487,N_49107);
or UO_4119 (O_4119,N_48632,N_49153);
xnor UO_4120 (O_4120,N_49257,N_49259);
nor UO_4121 (O_4121,N_49916,N_49528);
nand UO_4122 (O_4122,N_48033,N_49722);
or UO_4123 (O_4123,N_48939,N_48776);
nand UO_4124 (O_4124,N_48484,N_49871);
nand UO_4125 (O_4125,N_48120,N_48006);
or UO_4126 (O_4126,N_49159,N_49419);
and UO_4127 (O_4127,N_48069,N_49873);
nor UO_4128 (O_4128,N_48354,N_49244);
or UO_4129 (O_4129,N_48608,N_48345);
or UO_4130 (O_4130,N_49417,N_49898);
and UO_4131 (O_4131,N_49046,N_49379);
nand UO_4132 (O_4132,N_49506,N_48262);
and UO_4133 (O_4133,N_48714,N_48439);
nand UO_4134 (O_4134,N_49442,N_48016);
and UO_4135 (O_4135,N_48478,N_48613);
nor UO_4136 (O_4136,N_49888,N_49664);
and UO_4137 (O_4137,N_48796,N_49694);
nand UO_4138 (O_4138,N_49651,N_48141);
xor UO_4139 (O_4139,N_49335,N_48599);
or UO_4140 (O_4140,N_48735,N_49682);
and UO_4141 (O_4141,N_49830,N_48005);
and UO_4142 (O_4142,N_49444,N_49265);
xnor UO_4143 (O_4143,N_48369,N_48598);
nand UO_4144 (O_4144,N_49442,N_49835);
and UO_4145 (O_4145,N_49824,N_49256);
xor UO_4146 (O_4146,N_49333,N_49738);
nand UO_4147 (O_4147,N_49401,N_49683);
and UO_4148 (O_4148,N_49970,N_48352);
xnor UO_4149 (O_4149,N_49145,N_48532);
or UO_4150 (O_4150,N_49027,N_49201);
nor UO_4151 (O_4151,N_48471,N_49861);
nor UO_4152 (O_4152,N_48141,N_49022);
or UO_4153 (O_4153,N_48498,N_48368);
and UO_4154 (O_4154,N_49679,N_49394);
nand UO_4155 (O_4155,N_48693,N_49758);
or UO_4156 (O_4156,N_48939,N_49225);
or UO_4157 (O_4157,N_49034,N_49062);
nand UO_4158 (O_4158,N_48787,N_48874);
and UO_4159 (O_4159,N_49594,N_49176);
nor UO_4160 (O_4160,N_48488,N_48782);
nand UO_4161 (O_4161,N_49558,N_49963);
and UO_4162 (O_4162,N_48353,N_49980);
nor UO_4163 (O_4163,N_49446,N_49854);
or UO_4164 (O_4164,N_49857,N_49668);
nand UO_4165 (O_4165,N_49414,N_48437);
and UO_4166 (O_4166,N_48027,N_48423);
or UO_4167 (O_4167,N_49699,N_49243);
or UO_4168 (O_4168,N_49413,N_49554);
nor UO_4169 (O_4169,N_48399,N_48485);
or UO_4170 (O_4170,N_48111,N_48292);
nand UO_4171 (O_4171,N_48746,N_48393);
nand UO_4172 (O_4172,N_49211,N_49110);
xor UO_4173 (O_4173,N_48819,N_49061);
nor UO_4174 (O_4174,N_48686,N_49995);
and UO_4175 (O_4175,N_49376,N_48632);
xor UO_4176 (O_4176,N_48328,N_48142);
nand UO_4177 (O_4177,N_48383,N_49530);
nand UO_4178 (O_4178,N_48656,N_48731);
or UO_4179 (O_4179,N_48582,N_49306);
nor UO_4180 (O_4180,N_48548,N_48848);
and UO_4181 (O_4181,N_48392,N_48200);
or UO_4182 (O_4182,N_48585,N_49000);
nor UO_4183 (O_4183,N_49633,N_48457);
nor UO_4184 (O_4184,N_49396,N_48560);
nand UO_4185 (O_4185,N_49873,N_48672);
and UO_4186 (O_4186,N_49153,N_48543);
xnor UO_4187 (O_4187,N_48682,N_48415);
nand UO_4188 (O_4188,N_49128,N_49085);
xor UO_4189 (O_4189,N_49178,N_49965);
or UO_4190 (O_4190,N_48331,N_48153);
and UO_4191 (O_4191,N_48999,N_49818);
or UO_4192 (O_4192,N_48802,N_48806);
nand UO_4193 (O_4193,N_49953,N_49998);
nand UO_4194 (O_4194,N_49467,N_48763);
nor UO_4195 (O_4195,N_48772,N_49694);
nor UO_4196 (O_4196,N_49778,N_49690);
or UO_4197 (O_4197,N_49288,N_49393);
xnor UO_4198 (O_4198,N_49970,N_49538);
xor UO_4199 (O_4199,N_49476,N_48121);
nand UO_4200 (O_4200,N_48146,N_48497);
and UO_4201 (O_4201,N_48475,N_48331);
and UO_4202 (O_4202,N_48080,N_48638);
nor UO_4203 (O_4203,N_48228,N_49347);
nor UO_4204 (O_4204,N_48918,N_48600);
nand UO_4205 (O_4205,N_48234,N_49386);
and UO_4206 (O_4206,N_49096,N_49022);
or UO_4207 (O_4207,N_49874,N_48302);
and UO_4208 (O_4208,N_48652,N_48680);
or UO_4209 (O_4209,N_48422,N_49048);
nor UO_4210 (O_4210,N_48102,N_48017);
nand UO_4211 (O_4211,N_48023,N_48799);
xor UO_4212 (O_4212,N_49712,N_49589);
or UO_4213 (O_4213,N_49406,N_49274);
or UO_4214 (O_4214,N_49075,N_49467);
nor UO_4215 (O_4215,N_48361,N_49949);
or UO_4216 (O_4216,N_48671,N_48273);
nand UO_4217 (O_4217,N_49369,N_49514);
nand UO_4218 (O_4218,N_48722,N_49022);
xnor UO_4219 (O_4219,N_48775,N_49912);
and UO_4220 (O_4220,N_49585,N_49614);
xnor UO_4221 (O_4221,N_48255,N_48743);
nor UO_4222 (O_4222,N_49136,N_49694);
nor UO_4223 (O_4223,N_49740,N_49951);
nor UO_4224 (O_4224,N_48253,N_48590);
nand UO_4225 (O_4225,N_48815,N_49665);
nand UO_4226 (O_4226,N_49076,N_49803);
nor UO_4227 (O_4227,N_48989,N_49416);
and UO_4228 (O_4228,N_48943,N_49609);
and UO_4229 (O_4229,N_49683,N_48524);
and UO_4230 (O_4230,N_49738,N_49435);
xor UO_4231 (O_4231,N_49561,N_49327);
nor UO_4232 (O_4232,N_48447,N_48047);
nand UO_4233 (O_4233,N_49529,N_49728);
or UO_4234 (O_4234,N_48683,N_48406);
nor UO_4235 (O_4235,N_48680,N_48768);
nor UO_4236 (O_4236,N_49938,N_49200);
or UO_4237 (O_4237,N_48250,N_48717);
xor UO_4238 (O_4238,N_48575,N_49901);
nor UO_4239 (O_4239,N_49701,N_49572);
nor UO_4240 (O_4240,N_48029,N_49303);
nor UO_4241 (O_4241,N_49948,N_48647);
and UO_4242 (O_4242,N_49571,N_49289);
nor UO_4243 (O_4243,N_49241,N_48942);
nor UO_4244 (O_4244,N_48765,N_49440);
nand UO_4245 (O_4245,N_49836,N_49981);
or UO_4246 (O_4246,N_49436,N_48456);
xnor UO_4247 (O_4247,N_48289,N_48577);
nor UO_4248 (O_4248,N_48062,N_48218);
or UO_4249 (O_4249,N_49110,N_48412);
and UO_4250 (O_4250,N_48752,N_49549);
nor UO_4251 (O_4251,N_48743,N_48779);
and UO_4252 (O_4252,N_49898,N_49893);
or UO_4253 (O_4253,N_48914,N_48676);
nand UO_4254 (O_4254,N_48019,N_49530);
or UO_4255 (O_4255,N_48321,N_49405);
xor UO_4256 (O_4256,N_48598,N_48636);
xnor UO_4257 (O_4257,N_49167,N_49159);
and UO_4258 (O_4258,N_48024,N_48591);
nand UO_4259 (O_4259,N_48995,N_49316);
nor UO_4260 (O_4260,N_49378,N_48273);
nand UO_4261 (O_4261,N_48824,N_48078);
nand UO_4262 (O_4262,N_49604,N_49613);
nand UO_4263 (O_4263,N_48597,N_48957);
and UO_4264 (O_4264,N_49252,N_49763);
and UO_4265 (O_4265,N_48055,N_48890);
nor UO_4266 (O_4266,N_49299,N_49067);
and UO_4267 (O_4267,N_48955,N_49536);
or UO_4268 (O_4268,N_49906,N_49030);
and UO_4269 (O_4269,N_48724,N_48619);
or UO_4270 (O_4270,N_48192,N_48406);
xor UO_4271 (O_4271,N_48562,N_48468);
xnor UO_4272 (O_4272,N_49521,N_48727);
and UO_4273 (O_4273,N_49064,N_48171);
and UO_4274 (O_4274,N_49867,N_48461);
and UO_4275 (O_4275,N_49848,N_49768);
or UO_4276 (O_4276,N_48465,N_48526);
and UO_4277 (O_4277,N_48080,N_49759);
and UO_4278 (O_4278,N_49721,N_49311);
xor UO_4279 (O_4279,N_48881,N_49698);
xnor UO_4280 (O_4280,N_48966,N_48509);
nor UO_4281 (O_4281,N_49085,N_48543);
and UO_4282 (O_4282,N_49032,N_49826);
nor UO_4283 (O_4283,N_49194,N_48235);
nor UO_4284 (O_4284,N_48152,N_49671);
nor UO_4285 (O_4285,N_48950,N_49207);
and UO_4286 (O_4286,N_48891,N_49109);
xnor UO_4287 (O_4287,N_48355,N_49434);
nor UO_4288 (O_4288,N_49152,N_49614);
nor UO_4289 (O_4289,N_49855,N_49715);
and UO_4290 (O_4290,N_48093,N_48187);
xnor UO_4291 (O_4291,N_48002,N_48961);
nand UO_4292 (O_4292,N_49818,N_48570);
nand UO_4293 (O_4293,N_48985,N_48915);
nand UO_4294 (O_4294,N_49210,N_48247);
or UO_4295 (O_4295,N_49994,N_48138);
nand UO_4296 (O_4296,N_48564,N_48061);
xor UO_4297 (O_4297,N_48129,N_49864);
nor UO_4298 (O_4298,N_49817,N_48586);
nand UO_4299 (O_4299,N_48236,N_49086);
or UO_4300 (O_4300,N_49454,N_49575);
and UO_4301 (O_4301,N_49607,N_48116);
xor UO_4302 (O_4302,N_49276,N_49620);
nor UO_4303 (O_4303,N_48071,N_48984);
nor UO_4304 (O_4304,N_49340,N_49331);
nor UO_4305 (O_4305,N_48509,N_49926);
nor UO_4306 (O_4306,N_49518,N_49345);
nand UO_4307 (O_4307,N_49191,N_49359);
xnor UO_4308 (O_4308,N_49770,N_48169);
nor UO_4309 (O_4309,N_49994,N_48484);
nand UO_4310 (O_4310,N_49113,N_49561);
xor UO_4311 (O_4311,N_49730,N_49642);
xor UO_4312 (O_4312,N_48427,N_49735);
nor UO_4313 (O_4313,N_49934,N_49198);
or UO_4314 (O_4314,N_49494,N_48926);
and UO_4315 (O_4315,N_48311,N_49749);
nand UO_4316 (O_4316,N_49698,N_48359);
and UO_4317 (O_4317,N_49802,N_48466);
nor UO_4318 (O_4318,N_48736,N_49734);
nor UO_4319 (O_4319,N_49754,N_49096);
or UO_4320 (O_4320,N_48715,N_49975);
or UO_4321 (O_4321,N_49924,N_49580);
or UO_4322 (O_4322,N_49051,N_48286);
xnor UO_4323 (O_4323,N_48897,N_49018);
xnor UO_4324 (O_4324,N_48795,N_48530);
nand UO_4325 (O_4325,N_49002,N_48254);
nand UO_4326 (O_4326,N_49034,N_49706);
xnor UO_4327 (O_4327,N_48080,N_49075);
nand UO_4328 (O_4328,N_48810,N_49800);
nor UO_4329 (O_4329,N_49126,N_49691);
nor UO_4330 (O_4330,N_49957,N_48298);
and UO_4331 (O_4331,N_49927,N_48445);
or UO_4332 (O_4332,N_49636,N_48960);
nand UO_4333 (O_4333,N_48985,N_49710);
xor UO_4334 (O_4334,N_49946,N_49511);
nand UO_4335 (O_4335,N_48127,N_48489);
nand UO_4336 (O_4336,N_49915,N_49923);
nor UO_4337 (O_4337,N_49830,N_49487);
and UO_4338 (O_4338,N_49338,N_49935);
or UO_4339 (O_4339,N_48877,N_49973);
nand UO_4340 (O_4340,N_48566,N_48790);
or UO_4341 (O_4341,N_49784,N_48904);
xor UO_4342 (O_4342,N_48467,N_49495);
and UO_4343 (O_4343,N_48012,N_48636);
nor UO_4344 (O_4344,N_48352,N_48747);
nand UO_4345 (O_4345,N_48707,N_48335);
nand UO_4346 (O_4346,N_48294,N_48349);
xnor UO_4347 (O_4347,N_49910,N_49088);
xnor UO_4348 (O_4348,N_49586,N_49872);
nor UO_4349 (O_4349,N_48471,N_49935);
and UO_4350 (O_4350,N_48867,N_48813);
nor UO_4351 (O_4351,N_49998,N_48320);
nor UO_4352 (O_4352,N_49291,N_48731);
nand UO_4353 (O_4353,N_48716,N_48415);
and UO_4354 (O_4354,N_48265,N_49933);
nor UO_4355 (O_4355,N_49195,N_48950);
xor UO_4356 (O_4356,N_48680,N_49706);
or UO_4357 (O_4357,N_48449,N_49016);
and UO_4358 (O_4358,N_49304,N_49919);
nand UO_4359 (O_4359,N_49081,N_48364);
and UO_4360 (O_4360,N_49160,N_49371);
or UO_4361 (O_4361,N_48290,N_49657);
xor UO_4362 (O_4362,N_49211,N_49964);
or UO_4363 (O_4363,N_49454,N_49277);
nand UO_4364 (O_4364,N_49960,N_49535);
or UO_4365 (O_4365,N_48914,N_48054);
and UO_4366 (O_4366,N_49997,N_48635);
or UO_4367 (O_4367,N_48559,N_48145);
or UO_4368 (O_4368,N_48484,N_49920);
xnor UO_4369 (O_4369,N_48588,N_48619);
and UO_4370 (O_4370,N_48861,N_49087);
xnor UO_4371 (O_4371,N_48425,N_49327);
xor UO_4372 (O_4372,N_48589,N_49782);
and UO_4373 (O_4373,N_49899,N_48314);
nor UO_4374 (O_4374,N_48232,N_49710);
nor UO_4375 (O_4375,N_49915,N_48882);
xor UO_4376 (O_4376,N_48619,N_48301);
nand UO_4377 (O_4377,N_48250,N_49029);
and UO_4378 (O_4378,N_48200,N_48133);
and UO_4379 (O_4379,N_49479,N_48599);
or UO_4380 (O_4380,N_48724,N_48535);
or UO_4381 (O_4381,N_49220,N_48873);
and UO_4382 (O_4382,N_48529,N_49810);
or UO_4383 (O_4383,N_49285,N_49257);
and UO_4384 (O_4384,N_49007,N_48452);
xnor UO_4385 (O_4385,N_48383,N_48958);
and UO_4386 (O_4386,N_48994,N_49036);
nor UO_4387 (O_4387,N_49278,N_49012);
or UO_4388 (O_4388,N_48372,N_49677);
or UO_4389 (O_4389,N_48536,N_48470);
or UO_4390 (O_4390,N_48463,N_49604);
and UO_4391 (O_4391,N_48136,N_49696);
and UO_4392 (O_4392,N_49266,N_49267);
xor UO_4393 (O_4393,N_49664,N_48189);
nor UO_4394 (O_4394,N_48292,N_48641);
xnor UO_4395 (O_4395,N_48810,N_48068);
xor UO_4396 (O_4396,N_48485,N_48864);
nor UO_4397 (O_4397,N_48979,N_49321);
xor UO_4398 (O_4398,N_49733,N_48159);
and UO_4399 (O_4399,N_48027,N_48253);
and UO_4400 (O_4400,N_49706,N_48267);
or UO_4401 (O_4401,N_49518,N_49440);
nor UO_4402 (O_4402,N_48414,N_49432);
or UO_4403 (O_4403,N_48349,N_49699);
xor UO_4404 (O_4404,N_49952,N_48355);
nand UO_4405 (O_4405,N_49020,N_48104);
xnor UO_4406 (O_4406,N_48425,N_49050);
or UO_4407 (O_4407,N_48975,N_48165);
or UO_4408 (O_4408,N_48984,N_48955);
xor UO_4409 (O_4409,N_48513,N_49680);
xnor UO_4410 (O_4410,N_49986,N_49105);
nor UO_4411 (O_4411,N_48412,N_48048);
nand UO_4412 (O_4412,N_48497,N_48153);
nand UO_4413 (O_4413,N_48847,N_49176);
nor UO_4414 (O_4414,N_49876,N_48800);
nor UO_4415 (O_4415,N_48457,N_49525);
nor UO_4416 (O_4416,N_48802,N_48307);
xor UO_4417 (O_4417,N_49946,N_48962);
and UO_4418 (O_4418,N_49740,N_49631);
nor UO_4419 (O_4419,N_48212,N_48502);
xnor UO_4420 (O_4420,N_48261,N_48620);
or UO_4421 (O_4421,N_48494,N_48645);
or UO_4422 (O_4422,N_48060,N_48089);
or UO_4423 (O_4423,N_48163,N_48651);
or UO_4424 (O_4424,N_48240,N_48484);
nor UO_4425 (O_4425,N_48784,N_48094);
xnor UO_4426 (O_4426,N_49557,N_48526);
xnor UO_4427 (O_4427,N_49276,N_49022);
xor UO_4428 (O_4428,N_49308,N_48887);
nor UO_4429 (O_4429,N_49692,N_49490);
nor UO_4430 (O_4430,N_49142,N_49320);
or UO_4431 (O_4431,N_49175,N_49848);
and UO_4432 (O_4432,N_49957,N_49230);
and UO_4433 (O_4433,N_49454,N_48778);
or UO_4434 (O_4434,N_49988,N_48096);
and UO_4435 (O_4435,N_49634,N_49679);
and UO_4436 (O_4436,N_48143,N_48684);
nor UO_4437 (O_4437,N_48076,N_48094);
and UO_4438 (O_4438,N_48886,N_48568);
nand UO_4439 (O_4439,N_48452,N_48198);
nor UO_4440 (O_4440,N_49705,N_48117);
nand UO_4441 (O_4441,N_49046,N_48369);
or UO_4442 (O_4442,N_48118,N_48741);
or UO_4443 (O_4443,N_49656,N_48522);
nand UO_4444 (O_4444,N_48206,N_49528);
nor UO_4445 (O_4445,N_49956,N_49636);
or UO_4446 (O_4446,N_49324,N_48636);
nor UO_4447 (O_4447,N_48120,N_49464);
or UO_4448 (O_4448,N_49893,N_49990);
nor UO_4449 (O_4449,N_48119,N_49858);
and UO_4450 (O_4450,N_48974,N_49834);
and UO_4451 (O_4451,N_49515,N_48845);
and UO_4452 (O_4452,N_48687,N_49207);
and UO_4453 (O_4453,N_49211,N_49306);
or UO_4454 (O_4454,N_48449,N_48908);
nand UO_4455 (O_4455,N_49597,N_48361);
and UO_4456 (O_4456,N_48959,N_48936);
and UO_4457 (O_4457,N_49996,N_48374);
and UO_4458 (O_4458,N_48336,N_48827);
nand UO_4459 (O_4459,N_48046,N_49442);
and UO_4460 (O_4460,N_48117,N_48893);
nand UO_4461 (O_4461,N_49637,N_48363);
or UO_4462 (O_4462,N_49491,N_49809);
and UO_4463 (O_4463,N_49447,N_49101);
nand UO_4464 (O_4464,N_49579,N_48155);
nor UO_4465 (O_4465,N_49165,N_48328);
or UO_4466 (O_4466,N_49364,N_48434);
and UO_4467 (O_4467,N_48800,N_49221);
xnor UO_4468 (O_4468,N_49776,N_49902);
or UO_4469 (O_4469,N_48793,N_49389);
and UO_4470 (O_4470,N_48721,N_49546);
xnor UO_4471 (O_4471,N_49439,N_48511);
and UO_4472 (O_4472,N_49321,N_49493);
or UO_4473 (O_4473,N_48685,N_49517);
nand UO_4474 (O_4474,N_49481,N_48952);
nand UO_4475 (O_4475,N_48227,N_49373);
nor UO_4476 (O_4476,N_48815,N_48860);
nor UO_4477 (O_4477,N_49569,N_49150);
nor UO_4478 (O_4478,N_49851,N_48522);
nor UO_4479 (O_4479,N_48906,N_48572);
or UO_4480 (O_4480,N_48403,N_48910);
or UO_4481 (O_4481,N_49373,N_49387);
xnor UO_4482 (O_4482,N_49335,N_48518);
nand UO_4483 (O_4483,N_49839,N_48258);
nor UO_4484 (O_4484,N_49005,N_49976);
nor UO_4485 (O_4485,N_49476,N_48422);
xor UO_4486 (O_4486,N_49723,N_48764);
or UO_4487 (O_4487,N_48896,N_48789);
xor UO_4488 (O_4488,N_49986,N_49501);
and UO_4489 (O_4489,N_49360,N_48038);
xor UO_4490 (O_4490,N_48981,N_48872);
and UO_4491 (O_4491,N_49942,N_48021);
nor UO_4492 (O_4492,N_48240,N_48034);
xor UO_4493 (O_4493,N_48243,N_48851);
or UO_4494 (O_4494,N_49070,N_48354);
xor UO_4495 (O_4495,N_48932,N_48909);
nor UO_4496 (O_4496,N_48979,N_48715);
nor UO_4497 (O_4497,N_49735,N_49707);
or UO_4498 (O_4498,N_49387,N_48523);
nor UO_4499 (O_4499,N_48048,N_48382);
or UO_4500 (O_4500,N_48186,N_48572);
nor UO_4501 (O_4501,N_48640,N_48953);
and UO_4502 (O_4502,N_48198,N_48335);
nor UO_4503 (O_4503,N_48570,N_48048);
and UO_4504 (O_4504,N_49121,N_48834);
and UO_4505 (O_4505,N_48926,N_49094);
nand UO_4506 (O_4506,N_48455,N_49147);
and UO_4507 (O_4507,N_49317,N_49012);
and UO_4508 (O_4508,N_48975,N_48639);
xnor UO_4509 (O_4509,N_49819,N_48990);
and UO_4510 (O_4510,N_49150,N_48277);
and UO_4511 (O_4511,N_48147,N_49566);
or UO_4512 (O_4512,N_48331,N_49833);
xnor UO_4513 (O_4513,N_49614,N_49731);
and UO_4514 (O_4514,N_48226,N_49850);
nand UO_4515 (O_4515,N_49394,N_49945);
xnor UO_4516 (O_4516,N_49849,N_49118);
nand UO_4517 (O_4517,N_49114,N_48372);
nand UO_4518 (O_4518,N_48036,N_49192);
nor UO_4519 (O_4519,N_48694,N_48488);
nor UO_4520 (O_4520,N_48658,N_49315);
xor UO_4521 (O_4521,N_48000,N_49730);
nor UO_4522 (O_4522,N_48982,N_49219);
or UO_4523 (O_4523,N_49644,N_49356);
and UO_4524 (O_4524,N_49689,N_48468);
and UO_4525 (O_4525,N_49714,N_48921);
and UO_4526 (O_4526,N_48234,N_48073);
nand UO_4527 (O_4527,N_48987,N_49666);
nor UO_4528 (O_4528,N_49623,N_48820);
nand UO_4529 (O_4529,N_49371,N_49553);
nor UO_4530 (O_4530,N_48021,N_49832);
nor UO_4531 (O_4531,N_49222,N_48141);
xnor UO_4532 (O_4532,N_48488,N_49772);
nand UO_4533 (O_4533,N_49495,N_48295);
and UO_4534 (O_4534,N_49835,N_49947);
and UO_4535 (O_4535,N_49393,N_49271);
xor UO_4536 (O_4536,N_48202,N_49713);
nand UO_4537 (O_4537,N_48568,N_48013);
nand UO_4538 (O_4538,N_48371,N_49383);
and UO_4539 (O_4539,N_49940,N_48181);
nand UO_4540 (O_4540,N_48823,N_48340);
nand UO_4541 (O_4541,N_48267,N_49935);
and UO_4542 (O_4542,N_48133,N_48317);
and UO_4543 (O_4543,N_48184,N_49510);
nor UO_4544 (O_4544,N_49583,N_48252);
nand UO_4545 (O_4545,N_49103,N_48568);
xor UO_4546 (O_4546,N_48403,N_49692);
xor UO_4547 (O_4547,N_48530,N_49811);
or UO_4548 (O_4548,N_49628,N_49897);
or UO_4549 (O_4549,N_49691,N_49222);
nand UO_4550 (O_4550,N_48721,N_48085);
xor UO_4551 (O_4551,N_49759,N_48741);
xor UO_4552 (O_4552,N_49512,N_49471);
nand UO_4553 (O_4553,N_49087,N_49557);
xnor UO_4554 (O_4554,N_48796,N_48085);
nor UO_4555 (O_4555,N_48624,N_49661);
nor UO_4556 (O_4556,N_49845,N_48991);
nand UO_4557 (O_4557,N_48045,N_49711);
nor UO_4558 (O_4558,N_48543,N_48687);
xor UO_4559 (O_4559,N_49611,N_49024);
nand UO_4560 (O_4560,N_49651,N_48002);
xor UO_4561 (O_4561,N_48170,N_49285);
and UO_4562 (O_4562,N_49571,N_49639);
xnor UO_4563 (O_4563,N_49663,N_48710);
nor UO_4564 (O_4564,N_49972,N_49167);
nand UO_4565 (O_4565,N_48830,N_48408);
nand UO_4566 (O_4566,N_48955,N_48729);
xor UO_4567 (O_4567,N_48479,N_48585);
xor UO_4568 (O_4568,N_49123,N_49434);
nor UO_4569 (O_4569,N_49888,N_48736);
or UO_4570 (O_4570,N_48789,N_49188);
and UO_4571 (O_4571,N_48995,N_48033);
and UO_4572 (O_4572,N_49104,N_48051);
nand UO_4573 (O_4573,N_48970,N_48549);
and UO_4574 (O_4574,N_49096,N_48114);
nor UO_4575 (O_4575,N_48197,N_48895);
nor UO_4576 (O_4576,N_48844,N_48840);
or UO_4577 (O_4577,N_48501,N_49452);
nand UO_4578 (O_4578,N_49170,N_48845);
nor UO_4579 (O_4579,N_48527,N_48906);
xor UO_4580 (O_4580,N_48269,N_48436);
or UO_4581 (O_4581,N_49121,N_49897);
nor UO_4582 (O_4582,N_48199,N_48396);
and UO_4583 (O_4583,N_49223,N_48546);
xnor UO_4584 (O_4584,N_49155,N_49003);
xnor UO_4585 (O_4585,N_48244,N_49514);
and UO_4586 (O_4586,N_49709,N_48542);
and UO_4587 (O_4587,N_48788,N_49498);
nand UO_4588 (O_4588,N_49181,N_49290);
xnor UO_4589 (O_4589,N_49026,N_49706);
and UO_4590 (O_4590,N_48003,N_48811);
nand UO_4591 (O_4591,N_49267,N_49643);
nand UO_4592 (O_4592,N_48294,N_48246);
nor UO_4593 (O_4593,N_49505,N_49601);
or UO_4594 (O_4594,N_48422,N_48844);
nand UO_4595 (O_4595,N_48563,N_49933);
or UO_4596 (O_4596,N_49844,N_48477);
and UO_4597 (O_4597,N_48892,N_49818);
nand UO_4598 (O_4598,N_49742,N_49901);
and UO_4599 (O_4599,N_49925,N_48837);
xnor UO_4600 (O_4600,N_48853,N_48515);
or UO_4601 (O_4601,N_48760,N_49942);
or UO_4602 (O_4602,N_48074,N_48500);
or UO_4603 (O_4603,N_48278,N_48203);
nor UO_4604 (O_4604,N_48816,N_48047);
and UO_4605 (O_4605,N_48131,N_49118);
xnor UO_4606 (O_4606,N_49263,N_48885);
xor UO_4607 (O_4607,N_49787,N_48619);
nor UO_4608 (O_4608,N_49201,N_48424);
nor UO_4609 (O_4609,N_48917,N_49536);
xor UO_4610 (O_4610,N_48148,N_48034);
nand UO_4611 (O_4611,N_49059,N_49816);
and UO_4612 (O_4612,N_48445,N_48798);
and UO_4613 (O_4613,N_48421,N_48303);
nor UO_4614 (O_4614,N_48056,N_48207);
and UO_4615 (O_4615,N_48889,N_48083);
xnor UO_4616 (O_4616,N_48359,N_48751);
nand UO_4617 (O_4617,N_48061,N_48908);
and UO_4618 (O_4618,N_49072,N_49865);
nor UO_4619 (O_4619,N_49850,N_48462);
or UO_4620 (O_4620,N_48368,N_49389);
xor UO_4621 (O_4621,N_48206,N_49025);
nand UO_4622 (O_4622,N_48200,N_49067);
nand UO_4623 (O_4623,N_48657,N_48916);
and UO_4624 (O_4624,N_49643,N_48151);
xor UO_4625 (O_4625,N_49637,N_48652);
or UO_4626 (O_4626,N_48503,N_49122);
xor UO_4627 (O_4627,N_49192,N_48948);
and UO_4628 (O_4628,N_49559,N_49371);
and UO_4629 (O_4629,N_49183,N_48726);
and UO_4630 (O_4630,N_48022,N_49685);
xor UO_4631 (O_4631,N_49917,N_49380);
or UO_4632 (O_4632,N_49705,N_48235);
xnor UO_4633 (O_4633,N_49143,N_48426);
or UO_4634 (O_4634,N_49854,N_49541);
and UO_4635 (O_4635,N_48171,N_48047);
or UO_4636 (O_4636,N_49281,N_48938);
or UO_4637 (O_4637,N_49517,N_48564);
nor UO_4638 (O_4638,N_48141,N_49838);
or UO_4639 (O_4639,N_49691,N_48097);
or UO_4640 (O_4640,N_48496,N_48093);
xor UO_4641 (O_4641,N_49242,N_48988);
nor UO_4642 (O_4642,N_48021,N_48116);
nand UO_4643 (O_4643,N_49057,N_48190);
nand UO_4644 (O_4644,N_49768,N_49660);
nand UO_4645 (O_4645,N_49565,N_49750);
xor UO_4646 (O_4646,N_49045,N_49770);
and UO_4647 (O_4647,N_48566,N_48642);
xor UO_4648 (O_4648,N_49010,N_48328);
xnor UO_4649 (O_4649,N_48742,N_49415);
nor UO_4650 (O_4650,N_48163,N_48351);
nand UO_4651 (O_4651,N_49629,N_48492);
or UO_4652 (O_4652,N_49805,N_49095);
xnor UO_4653 (O_4653,N_49605,N_48441);
nor UO_4654 (O_4654,N_48823,N_49298);
and UO_4655 (O_4655,N_49009,N_48834);
xnor UO_4656 (O_4656,N_48793,N_48066);
nor UO_4657 (O_4657,N_49162,N_48504);
nand UO_4658 (O_4658,N_48493,N_48004);
and UO_4659 (O_4659,N_49393,N_49123);
nand UO_4660 (O_4660,N_48870,N_48049);
nand UO_4661 (O_4661,N_49105,N_48670);
nor UO_4662 (O_4662,N_48678,N_49312);
or UO_4663 (O_4663,N_48662,N_49655);
and UO_4664 (O_4664,N_48921,N_48124);
nor UO_4665 (O_4665,N_48418,N_49604);
and UO_4666 (O_4666,N_49937,N_49316);
and UO_4667 (O_4667,N_49451,N_49433);
and UO_4668 (O_4668,N_49643,N_48747);
nand UO_4669 (O_4669,N_49613,N_49088);
xnor UO_4670 (O_4670,N_48644,N_48796);
xnor UO_4671 (O_4671,N_49477,N_48565);
nor UO_4672 (O_4672,N_49901,N_49156);
and UO_4673 (O_4673,N_48980,N_49505);
xor UO_4674 (O_4674,N_49355,N_48538);
nand UO_4675 (O_4675,N_49888,N_49965);
xnor UO_4676 (O_4676,N_49267,N_48439);
xnor UO_4677 (O_4677,N_49500,N_48294);
nor UO_4678 (O_4678,N_49669,N_49254);
or UO_4679 (O_4679,N_48854,N_49401);
nor UO_4680 (O_4680,N_49653,N_48456);
xor UO_4681 (O_4681,N_49075,N_49589);
and UO_4682 (O_4682,N_49324,N_49179);
nand UO_4683 (O_4683,N_48459,N_48192);
and UO_4684 (O_4684,N_49984,N_48465);
or UO_4685 (O_4685,N_49581,N_48416);
and UO_4686 (O_4686,N_48579,N_48075);
and UO_4687 (O_4687,N_49974,N_49699);
and UO_4688 (O_4688,N_48765,N_49082);
xnor UO_4689 (O_4689,N_48079,N_48203);
or UO_4690 (O_4690,N_49334,N_48924);
xnor UO_4691 (O_4691,N_48866,N_48259);
or UO_4692 (O_4692,N_48935,N_49076);
nor UO_4693 (O_4693,N_49272,N_49207);
and UO_4694 (O_4694,N_49233,N_48664);
xnor UO_4695 (O_4695,N_48903,N_48657);
xnor UO_4696 (O_4696,N_48775,N_49447);
and UO_4697 (O_4697,N_48774,N_49742);
or UO_4698 (O_4698,N_49481,N_48188);
nor UO_4699 (O_4699,N_49617,N_48471);
or UO_4700 (O_4700,N_49880,N_48759);
xnor UO_4701 (O_4701,N_49874,N_48521);
xor UO_4702 (O_4702,N_48299,N_49007);
and UO_4703 (O_4703,N_48995,N_48912);
or UO_4704 (O_4704,N_49665,N_49652);
nand UO_4705 (O_4705,N_48148,N_49134);
xor UO_4706 (O_4706,N_48481,N_48811);
or UO_4707 (O_4707,N_49122,N_49855);
or UO_4708 (O_4708,N_49060,N_48050);
nor UO_4709 (O_4709,N_48563,N_49446);
xnor UO_4710 (O_4710,N_49753,N_48210);
and UO_4711 (O_4711,N_49555,N_49234);
nand UO_4712 (O_4712,N_48662,N_48882);
or UO_4713 (O_4713,N_49826,N_48912);
and UO_4714 (O_4714,N_48897,N_48714);
and UO_4715 (O_4715,N_49029,N_48404);
nor UO_4716 (O_4716,N_48513,N_49354);
nor UO_4717 (O_4717,N_49812,N_49056);
or UO_4718 (O_4718,N_49307,N_49397);
xnor UO_4719 (O_4719,N_48497,N_48985);
xor UO_4720 (O_4720,N_48516,N_48485);
nor UO_4721 (O_4721,N_49260,N_48405);
nor UO_4722 (O_4722,N_48022,N_48748);
nand UO_4723 (O_4723,N_49292,N_48357);
and UO_4724 (O_4724,N_49269,N_48176);
nor UO_4725 (O_4725,N_49730,N_48874);
nand UO_4726 (O_4726,N_49064,N_49265);
nand UO_4727 (O_4727,N_49044,N_48886);
nor UO_4728 (O_4728,N_49102,N_49213);
or UO_4729 (O_4729,N_48435,N_48330);
xor UO_4730 (O_4730,N_48020,N_49937);
and UO_4731 (O_4731,N_48161,N_48063);
nor UO_4732 (O_4732,N_48380,N_48166);
nand UO_4733 (O_4733,N_48708,N_49344);
xor UO_4734 (O_4734,N_49724,N_49117);
or UO_4735 (O_4735,N_49765,N_48093);
and UO_4736 (O_4736,N_48373,N_48952);
nand UO_4737 (O_4737,N_49948,N_49895);
xnor UO_4738 (O_4738,N_48224,N_49963);
nand UO_4739 (O_4739,N_49721,N_48071);
nor UO_4740 (O_4740,N_48199,N_48813);
and UO_4741 (O_4741,N_48685,N_49013);
or UO_4742 (O_4742,N_49898,N_49683);
or UO_4743 (O_4743,N_48704,N_48905);
xnor UO_4744 (O_4744,N_49337,N_49521);
and UO_4745 (O_4745,N_49285,N_49889);
and UO_4746 (O_4746,N_48638,N_48242);
and UO_4747 (O_4747,N_49043,N_49734);
or UO_4748 (O_4748,N_49894,N_48328);
xor UO_4749 (O_4749,N_48962,N_49787);
or UO_4750 (O_4750,N_49954,N_48920);
nand UO_4751 (O_4751,N_48184,N_48060);
nor UO_4752 (O_4752,N_49861,N_48685);
xor UO_4753 (O_4753,N_48344,N_49370);
nand UO_4754 (O_4754,N_48233,N_49296);
nor UO_4755 (O_4755,N_48524,N_48728);
and UO_4756 (O_4756,N_48043,N_48267);
and UO_4757 (O_4757,N_48276,N_48070);
or UO_4758 (O_4758,N_48535,N_49352);
or UO_4759 (O_4759,N_48620,N_48531);
xnor UO_4760 (O_4760,N_49855,N_49095);
or UO_4761 (O_4761,N_49243,N_48468);
xnor UO_4762 (O_4762,N_48139,N_49090);
xnor UO_4763 (O_4763,N_49217,N_49648);
nand UO_4764 (O_4764,N_48310,N_48405);
and UO_4765 (O_4765,N_49726,N_48053);
and UO_4766 (O_4766,N_48612,N_48783);
xor UO_4767 (O_4767,N_48263,N_49234);
xnor UO_4768 (O_4768,N_49940,N_48590);
nand UO_4769 (O_4769,N_48384,N_49477);
xnor UO_4770 (O_4770,N_48929,N_48027);
or UO_4771 (O_4771,N_48791,N_48323);
xnor UO_4772 (O_4772,N_49546,N_48488);
nand UO_4773 (O_4773,N_48229,N_48613);
or UO_4774 (O_4774,N_49123,N_49694);
nor UO_4775 (O_4775,N_49439,N_49091);
xnor UO_4776 (O_4776,N_48994,N_49057);
nor UO_4777 (O_4777,N_49458,N_49509);
and UO_4778 (O_4778,N_48134,N_48372);
nor UO_4779 (O_4779,N_49801,N_48874);
nand UO_4780 (O_4780,N_49838,N_49946);
nand UO_4781 (O_4781,N_48667,N_49506);
or UO_4782 (O_4782,N_49489,N_49766);
nand UO_4783 (O_4783,N_48195,N_48253);
or UO_4784 (O_4784,N_48453,N_49072);
nand UO_4785 (O_4785,N_48312,N_48757);
nor UO_4786 (O_4786,N_49432,N_49738);
xor UO_4787 (O_4787,N_49532,N_48675);
nor UO_4788 (O_4788,N_49659,N_48212);
and UO_4789 (O_4789,N_48053,N_49057);
nor UO_4790 (O_4790,N_48411,N_48875);
nor UO_4791 (O_4791,N_48780,N_49572);
nor UO_4792 (O_4792,N_49858,N_49608);
or UO_4793 (O_4793,N_48889,N_48626);
nand UO_4794 (O_4794,N_48684,N_49165);
and UO_4795 (O_4795,N_49605,N_49837);
nor UO_4796 (O_4796,N_48691,N_48562);
xor UO_4797 (O_4797,N_49841,N_49711);
xnor UO_4798 (O_4798,N_48020,N_49472);
nor UO_4799 (O_4799,N_49137,N_49403);
nand UO_4800 (O_4800,N_49101,N_49139);
or UO_4801 (O_4801,N_49770,N_48264);
or UO_4802 (O_4802,N_49110,N_49844);
or UO_4803 (O_4803,N_48186,N_48922);
nand UO_4804 (O_4804,N_48896,N_49037);
xor UO_4805 (O_4805,N_48816,N_49364);
nand UO_4806 (O_4806,N_48179,N_48761);
xnor UO_4807 (O_4807,N_49334,N_49875);
or UO_4808 (O_4808,N_48890,N_49602);
or UO_4809 (O_4809,N_48438,N_48966);
or UO_4810 (O_4810,N_48221,N_49138);
and UO_4811 (O_4811,N_48751,N_49863);
nor UO_4812 (O_4812,N_49592,N_48801);
xnor UO_4813 (O_4813,N_49556,N_48919);
and UO_4814 (O_4814,N_48022,N_49384);
xnor UO_4815 (O_4815,N_48049,N_49703);
and UO_4816 (O_4816,N_48617,N_49120);
and UO_4817 (O_4817,N_49573,N_48503);
and UO_4818 (O_4818,N_48190,N_49603);
nor UO_4819 (O_4819,N_48144,N_49248);
and UO_4820 (O_4820,N_48984,N_48082);
nor UO_4821 (O_4821,N_49733,N_48358);
xnor UO_4822 (O_4822,N_49512,N_49792);
nor UO_4823 (O_4823,N_49909,N_49004);
or UO_4824 (O_4824,N_48166,N_49264);
xor UO_4825 (O_4825,N_49136,N_49913);
and UO_4826 (O_4826,N_48660,N_49170);
xor UO_4827 (O_4827,N_48274,N_48920);
and UO_4828 (O_4828,N_48052,N_48861);
and UO_4829 (O_4829,N_48485,N_49592);
and UO_4830 (O_4830,N_48435,N_49803);
and UO_4831 (O_4831,N_48143,N_49871);
xor UO_4832 (O_4832,N_49443,N_48372);
xnor UO_4833 (O_4833,N_48471,N_49924);
xor UO_4834 (O_4834,N_49466,N_48252);
xnor UO_4835 (O_4835,N_48475,N_48254);
xnor UO_4836 (O_4836,N_49293,N_49321);
or UO_4837 (O_4837,N_48627,N_49857);
nor UO_4838 (O_4838,N_48697,N_48892);
and UO_4839 (O_4839,N_49106,N_49392);
and UO_4840 (O_4840,N_49166,N_48575);
nand UO_4841 (O_4841,N_49406,N_48438);
xnor UO_4842 (O_4842,N_49039,N_49512);
nor UO_4843 (O_4843,N_48426,N_48285);
and UO_4844 (O_4844,N_49452,N_49688);
nand UO_4845 (O_4845,N_49256,N_48336);
and UO_4846 (O_4846,N_48537,N_49818);
xor UO_4847 (O_4847,N_49894,N_49452);
or UO_4848 (O_4848,N_49407,N_49962);
xor UO_4849 (O_4849,N_49007,N_49239);
nand UO_4850 (O_4850,N_48111,N_49560);
nor UO_4851 (O_4851,N_48224,N_49450);
xnor UO_4852 (O_4852,N_49737,N_48818);
xor UO_4853 (O_4853,N_48508,N_49518);
or UO_4854 (O_4854,N_49115,N_49394);
or UO_4855 (O_4855,N_49419,N_48180);
nand UO_4856 (O_4856,N_48937,N_48619);
and UO_4857 (O_4857,N_49086,N_49397);
nand UO_4858 (O_4858,N_48984,N_49590);
and UO_4859 (O_4859,N_48755,N_48901);
xor UO_4860 (O_4860,N_49059,N_49740);
xnor UO_4861 (O_4861,N_49277,N_49012);
and UO_4862 (O_4862,N_49984,N_49485);
xor UO_4863 (O_4863,N_49038,N_49898);
and UO_4864 (O_4864,N_49172,N_49681);
xor UO_4865 (O_4865,N_48064,N_48636);
or UO_4866 (O_4866,N_48718,N_48218);
nor UO_4867 (O_4867,N_49937,N_49893);
and UO_4868 (O_4868,N_48029,N_49222);
and UO_4869 (O_4869,N_48332,N_49635);
nor UO_4870 (O_4870,N_49465,N_48851);
or UO_4871 (O_4871,N_48476,N_49650);
xnor UO_4872 (O_4872,N_49675,N_48030);
nand UO_4873 (O_4873,N_49682,N_48475);
and UO_4874 (O_4874,N_49179,N_49976);
xor UO_4875 (O_4875,N_49146,N_48771);
nand UO_4876 (O_4876,N_48369,N_48745);
nor UO_4877 (O_4877,N_49842,N_49522);
xnor UO_4878 (O_4878,N_49641,N_49009);
nor UO_4879 (O_4879,N_49082,N_48332);
and UO_4880 (O_4880,N_48579,N_49154);
or UO_4881 (O_4881,N_48642,N_48120);
nor UO_4882 (O_4882,N_48681,N_49897);
nand UO_4883 (O_4883,N_49623,N_49320);
xnor UO_4884 (O_4884,N_49498,N_48802);
or UO_4885 (O_4885,N_49585,N_49606);
nor UO_4886 (O_4886,N_49197,N_48987);
and UO_4887 (O_4887,N_48008,N_49834);
nand UO_4888 (O_4888,N_48095,N_48862);
or UO_4889 (O_4889,N_49105,N_48165);
xnor UO_4890 (O_4890,N_49020,N_48964);
and UO_4891 (O_4891,N_48056,N_49211);
xnor UO_4892 (O_4892,N_49478,N_48934);
nand UO_4893 (O_4893,N_48814,N_48375);
or UO_4894 (O_4894,N_48995,N_48249);
nand UO_4895 (O_4895,N_49676,N_48825);
nand UO_4896 (O_4896,N_49615,N_49649);
xnor UO_4897 (O_4897,N_49621,N_49651);
and UO_4898 (O_4898,N_49488,N_48813);
or UO_4899 (O_4899,N_48919,N_48158);
and UO_4900 (O_4900,N_48566,N_49147);
xor UO_4901 (O_4901,N_49040,N_49217);
nand UO_4902 (O_4902,N_49640,N_48860);
nand UO_4903 (O_4903,N_49455,N_49883);
xor UO_4904 (O_4904,N_49463,N_49032);
or UO_4905 (O_4905,N_49641,N_48453);
xnor UO_4906 (O_4906,N_48132,N_48777);
xnor UO_4907 (O_4907,N_48195,N_49695);
xor UO_4908 (O_4908,N_49944,N_48126);
nor UO_4909 (O_4909,N_48640,N_48560);
xor UO_4910 (O_4910,N_48602,N_48943);
nor UO_4911 (O_4911,N_48870,N_49987);
nand UO_4912 (O_4912,N_49228,N_48846);
xor UO_4913 (O_4913,N_48080,N_48699);
xnor UO_4914 (O_4914,N_49595,N_49264);
nand UO_4915 (O_4915,N_49859,N_48014);
xor UO_4916 (O_4916,N_49012,N_49992);
or UO_4917 (O_4917,N_48903,N_49270);
and UO_4918 (O_4918,N_48128,N_49753);
nand UO_4919 (O_4919,N_49583,N_48157);
xnor UO_4920 (O_4920,N_48998,N_49854);
nor UO_4921 (O_4921,N_48477,N_48528);
nor UO_4922 (O_4922,N_48648,N_48359);
nor UO_4923 (O_4923,N_48822,N_48493);
nand UO_4924 (O_4924,N_49904,N_48284);
xor UO_4925 (O_4925,N_49255,N_49567);
xnor UO_4926 (O_4926,N_49188,N_49000);
nor UO_4927 (O_4927,N_48880,N_49611);
nand UO_4928 (O_4928,N_48987,N_49555);
xor UO_4929 (O_4929,N_49854,N_49989);
and UO_4930 (O_4930,N_49041,N_48943);
xor UO_4931 (O_4931,N_48156,N_49026);
and UO_4932 (O_4932,N_48694,N_48791);
xnor UO_4933 (O_4933,N_48530,N_48825);
or UO_4934 (O_4934,N_49277,N_49395);
or UO_4935 (O_4935,N_48971,N_49008);
or UO_4936 (O_4936,N_49719,N_48255);
xnor UO_4937 (O_4937,N_48644,N_49242);
nand UO_4938 (O_4938,N_48381,N_49933);
nor UO_4939 (O_4939,N_49964,N_48331);
nand UO_4940 (O_4940,N_48561,N_48702);
nor UO_4941 (O_4941,N_48392,N_49885);
nor UO_4942 (O_4942,N_48468,N_49668);
xnor UO_4943 (O_4943,N_48329,N_49578);
and UO_4944 (O_4944,N_49271,N_48790);
or UO_4945 (O_4945,N_49726,N_48013);
xor UO_4946 (O_4946,N_48872,N_49802);
xor UO_4947 (O_4947,N_49479,N_49548);
and UO_4948 (O_4948,N_48970,N_48190);
nand UO_4949 (O_4949,N_49082,N_48306);
nand UO_4950 (O_4950,N_49895,N_48311);
nor UO_4951 (O_4951,N_48537,N_49699);
or UO_4952 (O_4952,N_48625,N_48029);
nor UO_4953 (O_4953,N_48827,N_48695);
nand UO_4954 (O_4954,N_49055,N_49557);
nand UO_4955 (O_4955,N_48028,N_49733);
and UO_4956 (O_4956,N_49243,N_48834);
or UO_4957 (O_4957,N_48895,N_48713);
and UO_4958 (O_4958,N_49598,N_48894);
xor UO_4959 (O_4959,N_49702,N_49281);
nor UO_4960 (O_4960,N_49934,N_48712);
and UO_4961 (O_4961,N_49407,N_49857);
or UO_4962 (O_4962,N_48928,N_48766);
nor UO_4963 (O_4963,N_49378,N_49351);
nand UO_4964 (O_4964,N_48468,N_48183);
nand UO_4965 (O_4965,N_49840,N_49691);
nor UO_4966 (O_4966,N_49895,N_48855);
nor UO_4967 (O_4967,N_49661,N_48714);
xnor UO_4968 (O_4968,N_49111,N_48272);
and UO_4969 (O_4969,N_48424,N_49982);
xor UO_4970 (O_4970,N_49478,N_48771);
xor UO_4971 (O_4971,N_48257,N_49528);
nor UO_4972 (O_4972,N_48230,N_48848);
or UO_4973 (O_4973,N_48325,N_48726);
and UO_4974 (O_4974,N_48902,N_49872);
xnor UO_4975 (O_4975,N_48853,N_49601);
nor UO_4976 (O_4976,N_48795,N_49804);
and UO_4977 (O_4977,N_48662,N_49467);
and UO_4978 (O_4978,N_49910,N_48605);
nand UO_4979 (O_4979,N_48831,N_49813);
or UO_4980 (O_4980,N_49546,N_49572);
nand UO_4981 (O_4981,N_49593,N_49231);
xor UO_4982 (O_4982,N_48783,N_49589);
nor UO_4983 (O_4983,N_49458,N_48279);
nor UO_4984 (O_4984,N_49991,N_49097);
nor UO_4985 (O_4985,N_48366,N_49914);
or UO_4986 (O_4986,N_49828,N_48545);
or UO_4987 (O_4987,N_49656,N_49664);
nor UO_4988 (O_4988,N_48246,N_49870);
and UO_4989 (O_4989,N_49326,N_48154);
xor UO_4990 (O_4990,N_48269,N_49145);
or UO_4991 (O_4991,N_49058,N_49718);
and UO_4992 (O_4992,N_49667,N_48370);
xor UO_4993 (O_4993,N_48197,N_49816);
nand UO_4994 (O_4994,N_48401,N_49660);
xor UO_4995 (O_4995,N_49889,N_49581);
and UO_4996 (O_4996,N_48260,N_49786);
or UO_4997 (O_4997,N_49821,N_49886);
nand UO_4998 (O_4998,N_48053,N_49546);
xnor UO_4999 (O_4999,N_48159,N_48362);
endmodule