module basic_2500_25000_3000_10_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nand U0 (N_0,In_974,In_260);
nor U1 (N_1,In_468,In_2224);
xor U2 (N_2,In_1344,In_1604);
or U3 (N_3,In_409,In_736);
xor U4 (N_4,In_669,In_2012);
nor U5 (N_5,In_1273,In_2464);
or U6 (N_6,In_1529,In_789);
and U7 (N_7,In_382,In_1536);
xor U8 (N_8,In_1620,In_828);
and U9 (N_9,In_1929,In_725);
or U10 (N_10,In_1833,In_2136);
nor U11 (N_11,In_2159,In_301);
or U12 (N_12,In_1678,In_1413);
and U13 (N_13,In_227,In_378);
xor U14 (N_14,In_1790,In_788);
and U15 (N_15,In_1939,In_2269);
and U16 (N_16,In_503,In_1417);
nor U17 (N_17,In_792,In_1108);
xnor U18 (N_18,In_1290,In_2027);
nand U19 (N_19,In_2015,In_2454);
nand U20 (N_20,In_380,In_1200);
xnor U21 (N_21,In_573,In_2069);
and U22 (N_22,In_1466,In_1071);
nand U23 (N_23,In_1325,In_2452);
or U24 (N_24,In_2161,In_2302);
or U25 (N_25,In_1803,In_1767);
and U26 (N_26,In_1192,In_1483);
nor U27 (N_27,In_2184,In_1927);
xnor U28 (N_28,In_593,In_1120);
nand U29 (N_29,In_2,In_2429);
xnor U30 (N_30,In_502,In_614);
or U31 (N_31,In_1625,In_1098);
nor U32 (N_32,In_553,In_1188);
nor U33 (N_33,In_2203,In_727);
and U34 (N_34,In_1133,In_1690);
nor U35 (N_35,In_1855,In_21);
xor U36 (N_36,In_2005,In_578);
and U37 (N_37,In_75,In_909);
xnor U38 (N_38,In_1713,In_2442);
nor U39 (N_39,In_1706,In_1135);
or U40 (N_40,In_1952,In_1011);
nand U41 (N_41,In_37,In_1172);
nand U42 (N_42,In_1727,In_918);
or U43 (N_43,In_2228,In_1209);
nand U44 (N_44,In_2384,In_979);
or U45 (N_45,In_2091,In_1680);
nor U46 (N_46,In_2309,In_1942);
nand U47 (N_47,In_1672,In_2474);
nand U48 (N_48,In_238,In_1136);
or U49 (N_49,In_371,In_1180);
nor U50 (N_50,In_747,In_1720);
nand U51 (N_51,In_2191,In_2242);
xnor U52 (N_52,In_256,In_1474);
nor U53 (N_53,In_667,In_726);
or U54 (N_54,In_293,In_1069);
xor U55 (N_55,In_1637,In_848);
and U56 (N_56,In_1844,In_1065);
nor U57 (N_57,In_29,In_2339);
and U58 (N_58,In_407,In_2077);
and U59 (N_59,In_749,In_2476);
nand U60 (N_60,In_560,In_2400);
or U61 (N_61,In_274,In_200);
and U62 (N_62,In_68,In_2209);
or U63 (N_63,In_517,In_1579);
nand U64 (N_64,In_2483,In_1428);
nand U65 (N_65,In_2223,In_1208);
xor U66 (N_66,In_2185,In_2214);
nor U67 (N_67,In_990,In_1350);
or U68 (N_68,In_510,In_2222);
xnor U69 (N_69,In_2215,In_1828);
nor U70 (N_70,In_719,In_2252);
nor U71 (N_71,In_2107,In_1718);
nand U72 (N_72,In_1294,In_1392);
and U73 (N_73,In_2248,In_2092);
or U74 (N_74,In_1326,In_2492);
nand U75 (N_75,In_1997,In_69);
nand U76 (N_76,In_1207,In_2084);
and U77 (N_77,In_152,In_800);
nand U78 (N_78,In_2162,In_988);
or U79 (N_79,In_169,In_529);
nor U80 (N_80,In_2102,In_1731);
or U81 (N_81,In_1534,In_1151);
and U82 (N_82,In_756,In_616);
nor U83 (N_83,In_760,In_1259);
and U84 (N_84,In_426,In_693);
and U85 (N_85,In_937,In_246);
nor U86 (N_86,In_1850,In_507);
xnor U87 (N_87,In_2180,In_1772);
nor U88 (N_88,In_1859,In_2381);
and U89 (N_89,In_1056,In_1184);
nand U90 (N_90,In_2078,In_2168);
nand U91 (N_91,In_1475,In_184);
xnor U92 (N_92,In_711,In_700);
nand U93 (N_93,In_189,In_1429);
or U94 (N_94,In_818,In_1610);
xnor U95 (N_95,In_427,In_154);
and U96 (N_96,In_1182,In_977);
nand U97 (N_97,In_420,In_251);
and U98 (N_98,In_316,In_1091);
xnor U99 (N_99,In_527,In_554);
or U100 (N_100,In_2221,In_561);
or U101 (N_101,In_2484,In_1492);
and U102 (N_102,In_2469,In_1682);
and U103 (N_103,In_42,In_2468);
and U104 (N_104,In_1478,In_1359);
nor U105 (N_105,In_414,In_932);
nand U106 (N_106,In_2439,In_2262);
nand U107 (N_107,In_226,In_1365);
xor U108 (N_108,In_992,In_2139);
and U109 (N_109,In_972,In_1078);
nor U110 (N_110,In_1622,In_2227);
nand U111 (N_111,In_2040,In_2048);
xnor U112 (N_112,In_743,In_322);
or U113 (N_113,In_197,In_1203);
and U114 (N_114,In_1097,In_998);
nor U115 (N_115,In_281,In_1452);
and U116 (N_116,In_34,In_1277);
or U117 (N_117,In_1112,In_1967);
or U118 (N_118,In_660,In_982);
xnor U119 (N_119,In_2423,In_1535);
nand U120 (N_120,In_1702,In_45);
nor U121 (N_121,In_54,In_2033);
xnor U122 (N_122,In_2275,In_803);
xnor U123 (N_123,In_1261,In_1132);
xnor U124 (N_124,In_2175,In_1827);
or U125 (N_125,In_213,In_359);
nor U126 (N_126,In_753,In_1571);
nand U127 (N_127,In_1383,In_526);
xnor U128 (N_128,In_1219,In_1079);
nor U129 (N_129,In_2019,In_1846);
nor U130 (N_130,In_910,In_2194);
nand U131 (N_131,In_941,In_1334);
xor U132 (N_132,In_1490,In_396);
or U133 (N_133,In_2082,In_1212);
nand U134 (N_134,In_858,In_185);
and U135 (N_135,In_1698,In_1746);
xor U136 (N_136,In_1569,In_2402);
nand U137 (N_137,In_1064,In_1020);
or U138 (N_138,In_1304,In_354);
nand U139 (N_139,In_110,In_417);
nor U140 (N_140,In_2499,In_1373);
nand U141 (N_141,In_1499,In_1287);
xor U142 (N_142,In_1444,In_2494);
xnor U143 (N_143,In_841,In_2325);
and U144 (N_144,In_1046,In_1454);
nor U145 (N_145,In_1934,In_366);
xnor U146 (N_146,In_2441,In_1202);
nand U147 (N_147,In_1119,In_897);
or U148 (N_148,In_2448,In_595);
nand U149 (N_149,In_1728,In_1494);
nor U150 (N_150,In_1531,In_934);
or U151 (N_151,In_1856,In_1761);
nor U152 (N_152,In_2308,In_437);
nand U153 (N_153,In_1305,In_576);
and U154 (N_154,In_1694,In_1804);
or U155 (N_155,In_239,In_2100);
nor U156 (N_156,In_597,In_2287);
xnor U157 (N_157,In_1652,In_1247);
or U158 (N_158,In_2213,In_97);
and U159 (N_159,In_1456,In_141);
nand U160 (N_160,In_1303,In_266);
or U161 (N_161,In_1745,In_41);
and U162 (N_162,In_583,In_1381);
nor U163 (N_163,In_477,In_892);
xor U164 (N_164,In_2349,In_400);
xor U165 (N_165,In_496,In_744);
and U166 (N_166,In_1817,In_2150);
xnor U167 (N_167,In_1530,In_1852);
nand U168 (N_168,In_1195,In_1029);
xnor U169 (N_169,In_2461,In_1440);
or U170 (N_170,In_1606,In_271);
xnor U171 (N_171,In_847,In_397);
or U172 (N_172,In_1236,In_1461);
nand U173 (N_173,In_108,In_1560);
xor U174 (N_174,In_5,In_938);
nand U175 (N_175,In_863,In_1051);
or U176 (N_176,In_1324,In_524);
or U177 (N_177,In_900,In_1962);
and U178 (N_178,In_2270,In_406);
and U179 (N_179,In_883,In_2394);
nand U180 (N_180,In_203,In_2080);
nor U181 (N_181,In_1345,In_484);
or U182 (N_182,In_1353,In_632);
xor U183 (N_183,In_2288,In_1991);
or U184 (N_184,In_2493,In_1221);
or U185 (N_185,In_1235,In_2202);
or U186 (N_186,In_544,In_133);
nor U187 (N_187,In_543,In_1885);
nor U188 (N_188,In_1960,In_882);
nor U189 (N_189,In_1544,In_1403);
or U190 (N_190,In_1282,In_1793);
and U191 (N_191,In_304,In_673);
or U192 (N_192,In_1214,In_1216);
and U193 (N_193,In_1917,In_43);
nor U194 (N_194,In_249,In_1555);
nor U195 (N_195,In_986,In_2419);
and U196 (N_196,In_369,In_2260);
nor U197 (N_197,In_2427,In_12);
nand U198 (N_198,In_757,In_1559);
xor U199 (N_199,In_1557,In_2052);
and U200 (N_200,In_1588,In_1027);
nor U201 (N_201,In_1522,In_209);
nor U202 (N_202,In_1600,In_646);
or U203 (N_203,In_2137,In_1425);
or U204 (N_204,In_1564,In_1455);
nand U205 (N_205,In_2146,In_2183);
nand U206 (N_206,In_334,In_2096);
nor U207 (N_207,In_1757,In_1969);
and U208 (N_208,In_2407,In_651);
nor U209 (N_209,In_1111,In_822);
and U210 (N_210,In_2356,In_443);
or U211 (N_211,In_2197,In_525);
xnor U212 (N_212,In_2470,In_27);
nor U213 (N_213,In_1408,In_2271);
nand U214 (N_214,In_175,In_621);
or U215 (N_215,In_1271,In_323);
and U216 (N_216,In_402,In_1603);
nand U217 (N_217,In_1882,In_1187);
nor U218 (N_218,In_1930,In_1217);
and U219 (N_219,In_1460,In_149);
nor U220 (N_220,In_1580,In_2031);
xor U221 (N_221,In_1193,In_2064);
nor U222 (N_222,In_124,In_2119);
or U223 (N_223,In_2389,In_1224);
xnor U224 (N_224,In_2436,In_665);
nor U225 (N_225,In_855,In_1986);
xnor U226 (N_226,In_1060,In_501);
nand U227 (N_227,In_729,In_2028);
xor U228 (N_228,In_2174,In_1080);
nor U229 (N_229,In_440,In_868);
nor U230 (N_230,In_1007,In_1178);
nand U231 (N_231,In_1329,In_2170);
nor U232 (N_232,In_2296,In_658);
and U233 (N_233,In_1726,In_2473);
xnor U234 (N_234,In_625,In_1031);
nand U235 (N_235,In_2061,In_288);
nor U236 (N_236,In_1375,In_2085);
or U237 (N_237,In_1553,In_1511);
or U238 (N_238,In_2334,In_338);
and U239 (N_239,In_1465,In_1124);
nand U240 (N_240,In_688,In_1890);
or U241 (N_241,In_1218,In_1122);
and U242 (N_242,In_2272,In_1293);
and U243 (N_243,In_123,In_1512);
nand U244 (N_244,In_257,In_1342);
xnor U245 (N_245,In_1558,In_1059);
and U246 (N_246,In_1707,In_664);
nor U247 (N_247,In_411,In_999);
nor U248 (N_248,In_1436,In_2313);
and U249 (N_249,In_2188,In_2243);
or U250 (N_250,In_1109,In_2340);
nor U251 (N_251,In_70,In_856);
or U252 (N_252,In_1158,In_1016);
xor U253 (N_253,In_423,In_1343);
and U254 (N_254,In_2290,In_691);
and U255 (N_255,In_1086,In_125);
xnor U256 (N_256,In_1909,In_1493);
nor U257 (N_257,In_408,In_733);
and U258 (N_258,In_2481,In_836);
and U259 (N_259,In_1479,In_709);
or U260 (N_260,In_1738,In_1094);
xor U261 (N_261,In_1264,In_1675);
nor U262 (N_262,In_1538,In_1156);
nand U263 (N_263,In_2018,In_547);
xnor U264 (N_264,In_2336,In_1575);
or U265 (N_265,In_585,In_1751);
nor U266 (N_266,In_2383,In_2433);
nor U267 (N_267,In_2006,In_2392);
nor U268 (N_268,In_1181,In_824);
nand U269 (N_269,In_105,In_532);
nand U270 (N_270,In_2259,In_603);
nor U271 (N_271,In_1813,In_2196);
nand U272 (N_272,In_1496,In_2014);
or U273 (N_273,In_1627,In_40);
or U274 (N_274,In_1647,In_145);
or U275 (N_275,In_214,In_1581);
or U276 (N_276,In_137,In_158);
nand U277 (N_277,In_1599,In_1858);
xnor U278 (N_278,In_857,In_920);
and U279 (N_279,In_2047,In_1765);
and U280 (N_280,In_568,In_280);
xnor U281 (N_281,In_1570,In_784);
xnor U282 (N_282,In_946,In_1777);
and U283 (N_283,In_2358,In_1352);
and U284 (N_284,In_1651,In_619);
nor U285 (N_285,In_319,In_1521);
and U286 (N_286,In_1543,In_1228);
or U287 (N_287,In_166,In_87);
xnor U288 (N_288,In_2479,In_1724);
xnor U289 (N_289,In_1023,In_22);
xnor U290 (N_290,In_1926,In_1470);
xnor U291 (N_291,In_1835,In_2432);
and U292 (N_292,In_707,In_1500);
and U293 (N_293,In_1129,In_1340);
nand U294 (N_294,In_1319,In_143);
and U295 (N_295,In_1337,In_1561);
and U296 (N_296,In_2003,In_1286);
nand U297 (N_297,In_126,In_1387);
nand U298 (N_298,In_550,In_113);
xor U299 (N_299,In_1306,In_235);
xnor U300 (N_300,In_710,In_331);
nand U301 (N_301,In_1307,In_686);
nand U302 (N_302,In_2333,In_1632);
and U303 (N_303,In_513,In_829);
xnor U304 (N_304,In_2330,In_2201);
nand U305 (N_305,In_1585,In_2477);
xor U306 (N_306,In_2059,In_33);
or U307 (N_307,In_773,In_146);
or U308 (N_308,In_2123,In_1696);
or U309 (N_309,In_2301,In_1809);
nand U310 (N_310,In_404,In_48);
nor U311 (N_311,In_1422,In_1635);
nor U312 (N_312,In_1223,In_1090);
nand U313 (N_313,In_1655,In_1262);
nor U314 (N_314,In_1710,In_2128);
and U315 (N_315,In_2486,In_499);
nand U316 (N_316,In_2368,In_2241);
and U317 (N_317,In_916,In_891);
xnor U318 (N_318,In_1315,In_1431);
nand U319 (N_319,In_1592,In_675);
xnor U320 (N_320,In_395,In_65);
xor U321 (N_321,In_2354,In_1398);
or U322 (N_322,In_655,In_1626);
or U323 (N_323,In_914,In_2387);
nand U324 (N_324,In_2025,In_1222);
xor U325 (N_325,In_357,In_365);
and U326 (N_326,In_1177,In_85);
nand U327 (N_327,In_1053,In_630);
xor U328 (N_328,In_970,In_571);
nand U329 (N_329,In_1684,In_2357);
nor U330 (N_330,In_38,In_1275);
or U331 (N_331,In_1054,In_1002);
xnor U332 (N_332,In_456,In_332);
and U333 (N_333,In_2446,In_802);
or U334 (N_334,In_1915,In_307);
xor U335 (N_335,In_204,In_292);
nand U336 (N_336,In_253,In_430);
xor U337 (N_337,In_845,In_295);
xnor U338 (N_338,In_1965,In_2366);
or U339 (N_339,In_1910,In_644);
xnor U340 (N_340,In_2478,In_1605);
nand U341 (N_341,In_2424,In_2253);
and U342 (N_342,In_210,In_2403);
xor U343 (N_343,In_52,In_2236);
xnor U344 (N_344,In_73,In_486);
or U345 (N_345,In_2449,In_61);
nand U346 (N_346,In_1577,In_1669);
or U347 (N_347,In_1831,In_95);
xor U348 (N_348,In_1643,In_261);
nand U349 (N_349,In_1593,In_771);
xnor U350 (N_350,In_1704,In_1732);
xnor U351 (N_351,In_564,In_1541);
nand U352 (N_352,In_1439,In_2007);
nand U353 (N_353,In_2435,In_1829);
nor U354 (N_354,In_1781,In_1049);
and U355 (N_355,In_966,In_627);
or U356 (N_356,In_721,In_91);
xor U357 (N_357,In_1658,In_305);
nand U358 (N_358,In_2495,In_1780);
nor U359 (N_359,In_790,In_1185);
xor U360 (N_360,In_572,In_88);
xnor U361 (N_361,In_1485,In_14);
and U362 (N_362,In_2193,In_1723);
nand U363 (N_363,In_83,In_864);
nor U364 (N_364,In_964,In_1442);
and U365 (N_365,In_391,In_1113);
xnor U366 (N_366,In_2192,In_2093);
nand U367 (N_367,In_718,In_755);
xor U368 (N_368,In_1895,In_874);
or U369 (N_369,In_2133,In_886);
nor U370 (N_370,In_1232,In_850);
and U371 (N_371,In_767,In_1339);
or U372 (N_372,In_649,In_642);
nor U373 (N_373,In_2022,In_942);
nor U374 (N_374,In_121,In_1378);
nand U375 (N_375,In_2276,In_1333);
nor U376 (N_376,In_1611,In_939);
nand U377 (N_377,In_201,In_2086);
or U378 (N_378,In_816,In_1887);
or U379 (N_379,In_894,In_2010);
nor U380 (N_380,In_264,In_1811);
or U381 (N_381,In_1115,In_1405);
nand U382 (N_382,In_860,In_866);
nor U383 (N_383,In_2051,In_796);
or U384 (N_384,In_1384,In_2053);
and U385 (N_385,In_958,In_351);
and U386 (N_386,In_1869,In_1504);
or U387 (N_387,In_361,In_350);
nand U388 (N_388,In_324,In_799);
or U389 (N_389,In_678,In_963);
xor U390 (N_390,In_1331,In_96);
and U391 (N_391,In_140,In_290);
and U392 (N_392,In_2362,In_2380);
nand U393 (N_393,In_1668,In_2447);
nor U394 (N_394,In_17,In_1379);
xor U395 (N_395,In_1285,In_1101);
nand U396 (N_396,In_2134,In_1576);
or U397 (N_397,In_2303,In_1041);
nor U398 (N_398,In_1750,In_1782);
and U399 (N_399,In_1545,In_1074);
nor U400 (N_400,In_340,In_1523);
xnor U401 (N_401,In_2285,In_155);
and U402 (N_402,In_392,In_1432);
or U403 (N_403,In_509,In_1248);
nand U404 (N_404,In_263,In_1154);
and U405 (N_405,In_381,In_1587);
and U406 (N_406,In_216,In_1533);
or U407 (N_407,In_738,In_666);
or U408 (N_408,In_1351,In_242);
and U409 (N_409,In_785,In_1372);
xor U410 (N_410,In_740,In_2067);
xor U411 (N_411,In_714,In_1471);
nand U412 (N_412,In_1888,In_1058);
and U413 (N_413,In_434,In_1240);
nor U414 (N_414,In_1875,In_663);
nor U415 (N_415,In_1367,In_383);
nand U416 (N_416,In_1584,In_1096);
or U417 (N_417,In_577,In_1001);
or U418 (N_418,In_2190,In_2050);
or U419 (N_419,In_310,In_1316);
nor U420 (N_420,In_314,In_2250);
or U421 (N_421,In_358,In_1540);
xnor U422 (N_422,In_2462,In_1088);
nor U423 (N_423,In_1100,In_814);
and U424 (N_424,In_2239,In_2391);
xnor U425 (N_425,In_821,In_1527);
or U426 (N_426,In_1872,In_1666);
and U427 (N_427,In_1601,In_1970);
nand U428 (N_428,In_849,In_1671);
and U429 (N_429,In_2471,In_2158);
nand U430 (N_430,In_893,In_89);
and U431 (N_431,In_1640,In_495);
nor U432 (N_432,In_565,In_2002);
nor U433 (N_433,In_62,In_162);
or U434 (N_434,In_1874,In_1725);
and U435 (N_435,In_705,In_840);
nand U436 (N_436,In_1018,In_1977);
or U437 (N_437,In_1328,In_929);
and U438 (N_438,In_794,In_2322);
nand U439 (N_439,In_2324,In_374);
nor U440 (N_440,In_432,In_168);
nand U441 (N_441,In_661,In_1255);
xnor U442 (N_442,In_1532,In_1902);
nor U443 (N_443,In_2127,In_1820);
or U444 (N_444,In_247,In_1589);
nand U445 (N_445,In_1225,In_1595);
or U446 (N_446,In_1737,In_1314);
nand U447 (N_447,In_2360,In_1194);
or U448 (N_448,In_1899,In_869);
and U449 (N_449,In_1267,In_1254);
nand U450 (N_450,In_450,In_1520);
or U451 (N_451,In_770,In_1841);
and U452 (N_452,In_442,In_1);
nor U453 (N_453,In_708,In_1994);
and U454 (N_454,In_2295,In_1019);
nand U455 (N_455,In_1562,In_438);
or U456 (N_456,In_1931,In_2345);
xor U457 (N_457,In_1574,In_1961);
and U458 (N_458,In_1839,In_1947);
or U459 (N_459,In_606,In_379);
or U460 (N_460,In_1130,In_1840);
and U461 (N_461,In_2109,In_530);
xor U462 (N_462,In_312,In_436);
nand U463 (N_463,In_2004,In_1061);
or U464 (N_464,In_2038,In_1760);
or U465 (N_465,In_1636,In_1884);
nor U466 (N_466,In_1701,In_741);
xor U467 (N_467,In_735,In_921);
or U468 (N_468,In_1369,In_701);
and U469 (N_469,In_1489,In_2099);
nand U470 (N_470,In_1443,In_2412);
nand U471 (N_471,In_2316,In_2140);
nor U472 (N_472,In_813,In_853);
and U473 (N_473,In_275,In_491);
nand U474 (N_474,In_925,In_1099);
or U475 (N_475,In_1693,In_1688);
xor U476 (N_476,In_1396,In_2042);
nand U477 (N_477,In_1318,In_940);
nand U478 (N_478,In_1972,In_580);
nor U479 (N_479,In_46,In_1799);
and U480 (N_480,In_132,In_1477);
and U481 (N_481,In_1983,In_1176);
nand U482 (N_482,In_556,In_602);
nor U483 (N_483,In_2444,In_2244);
nor U484 (N_484,In_2044,In_190);
xnor U485 (N_485,In_833,In_480);
nor U486 (N_486,In_1515,In_1753);
or U487 (N_487,In_245,In_1419);
or U488 (N_488,In_867,In_1513);
nand U489 (N_489,In_1362,In_2066);
nor U490 (N_490,In_2171,In_948);
or U491 (N_491,In_924,In_1729);
nand U492 (N_492,In_460,In_111);
and U493 (N_493,In_2312,In_1870);
nand U494 (N_494,In_763,In_533);
and U495 (N_495,In_1778,In_1245);
nor U496 (N_496,In_81,In_1998);
xnor U497 (N_497,In_10,In_498);
and U498 (N_498,In_278,In_78);
xor U499 (N_499,In_2320,In_1506);
or U500 (N_500,In_1137,In_2106);
xor U501 (N_501,In_333,In_2088);
or U502 (N_502,In_629,In_2315);
xnor U503 (N_503,In_1763,In_1618);
or U504 (N_504,In_255,In_1648);
nand U505 (N_505,In_224,In_552);
xor U506 (N_506,In_0,In_67);
and U507 (N_507,In_1276,In_2347);
nor U508 (N_508,In_471,In_1434);
xor U509 (N_509,In_2068,In_1191);
nor U510 (N_510,In_2135,In_1118);
nand U511 (N_511,In_2154,In_601);
nand U512 (N_512,In_151,In_1692);
xnor U513 (N_513,In_363,In_1186);
nand U514 (N_514,In_1025,In_1215);
or U515 (N_515,In_1292,In_1665);
nor U516 (N_516,In_960,In_823);
xor U517 (N_517,In_1518,In_2293);
or U518 (N_518,In_1774,In_368);
nor U519 (N_519,In_1048,In_2371);
nor U520 (N_520,In_588,In_1987);
or U521 (N_521,In_1551,In_782);
or U522 (N_522,In_862,In_1301);
or U523 (N_523,In_1982,In_2013);
nand U524 (N_524,In_902,In_1773);
nand U525 (N_525,In_712,In_959);
and U526 (N_526,In_273,In_90);
nor U527 (N_527,In_945,In_804);
nor U528 (N_528,In_1573,In_1166);
or U529 (N_529,In_1213,In_1338);
nand U530 (N_530,In_208,In_1451);
nand U531 (N_531,In_265,In_720);
and U532 (N_532,In_1903,In_2129);
xnor U533 (N_533,In_464,In_2212);
nand U534 (N_534,In_1596,In_1144);
xnor U535 (N_535,In_2480,In_49);
xor U536 (N_536,In_180,In_405);
nor U537 (N_537,In_682,In_1806);
xor U538 (N_538,In_876,In_807);
nand U539 (N_539,In_1299,In_1807);
xor U540 (N_540,In_2124,In_134);
or U541 (N_541,In_895,In_996);
xnor U542 (N_542,In_2445,In_1448);
nor U543 (N_543,In_1615,In_2342);
nand U544 (N_544,In_2155,In_2410);
nand U545 (N_545,In_1243,In_2409);
xor U546 (N_546,In_1689,In_2265);
nand U547 (N_547,In_1566,In_2103);
nand U548 (N_548,In_2310,In_35);
or U549 (N_549,In_1995,In_1582);
or U550 (N_550,In_742,In_871);
nand U551 (N_551,In_444,In_2405);
or U552 (N_552,In_587,In_2206);
or U553 (N_553,In_51,In_607);
or U554 (N_554,In_980,In_71);
or U555 (N_555,In_1220,In_177);
xnor U556 (N_556,In_1360,In_1568);
or U557 (N_557,In_1013,In_793);
xor U558 (N_558,In_2343,In_1653);
and U559 (N_559,In_1481,In_645);
nor U560 (N_560,In_1845,In_2177);
nand U561 (N_561,In_386,In_1586);
nor U562 (N_562,In_254,In_86);
xor U563 (N_563,In_419,In_952);
and U564 (N_564,In_540,In_1040);
or U565 (N_565,In_1837,In_1722);
and U566 (N_566,In_1968,In_1893);
or U567 (N_567,In_1958,In_26);
nor U568 (N_568,In_2251,In_697);
or U569 (N_569,In_689,In_336);
nand U570 (N_570,In_1183,In_993);
nor U571 (N_571,In_1676,In_1567);
or U572 (N_572,In_1873,In_1357);
nor U573 (N_573,In_172,In_2426);
and U574 (N_574,In_1528,In_1169);
and U575 (N_575,In_615,In_2497);
nand U576 (N_576,In_1883,In_1252);
or U577 (N_577,In_313,In_2087);
or U578 (N_578,In_983,In_1412);
or U579 (N_579,In_1851,In_2151);
nor U580 (N_580,In_2249,In_2034);
nor U581 (N_581,In_1095,In_1291);
xor U582 (N_582,In_1280,In_2122);
nand U583 (N_583,In_1085,In_412);
or U584 (N_584,In_1067,In_1450);
nor U585 (N_585,In_2267,In_2169);
or U586 (N_586,In_1445,In_1775);
nor U587 (N_587,In_1152,In_965);
or U588 (N_588,In_58,In_1681);
and U589 (N_589,In_1795,In_724);
xor U590 (N_590,In_2465,In_1755);
and U591 (N_591,In_1764,In_9);
and U592 (N_592,In_173,In_1548);
nor U593 (N_593,In_765,In_1552);
or U594 (N_594,In_706,In_622);
nand U595 (N_595,In_390,In_639);
nand U596 (N_596,In_971,In_157);
xor U597 (N_597,In_551,In_1789);
nor U598 (N_598,In_39,In_1736);
nor U599 (N_599,In_1009,In_1714);
and U600 (N_600,In_234,In_832);
or U601 (N_601,In_1393,In_1949);
nand U602 (N_602,In_2011,In_1649);
nand U603 (N_603,In_291,In_57);
nor U604 (N_604,In_566,In_2152);
nor U605 (N_605,In_489,In_953);
and U606 (N_606,In_1853,In_759);
nor U607 (N_607,In_912,In_20);
xor U608 (N_608,In_1128,In_318);
xor U609 (N_609,In_1519,In_1106);
xor U610 (N_610,In_1864,In_1971);
nor U611 (N_611,In_492,In_1230);
nand U612 (N_612,In_684,In_2001);
nor U613 (N_613,In_325,In_303);
xor U614 (N_614,In_1556,In_1289);
and U615 (N_615,In_752,In_812);
or U616 (N_616,In_648,In_817);
and U617 (N_617,In_1641,In_2142);
nor U618 (N_618,In_453,In_2189);
xnor U619 (N_619,In_928,In_1346);
nand U620 (N_620,In_320,In_2431);
xnor U621 (N_621,In_768,In_193);
nor U622 (N_622,In_259,In_1818);
or U623 (N_623,In_435,In_1539);
nor U624 (N_624,In_150,In_2437);
nor U625 (N_625,In_1925,In_2046);
nor U626 (N_626,In_2463,In_981);
nor U627 (N_627,In_2024,In_674);
and U628 (N_628,In_1231,In_978);
or U629 (N_629,In_2167,In_722);
or U630 (N_630,In_353,In_680);
nor U631 (N_631,In_1646,In_2365);
nor U632 (N_632,In_605,In_539);
and U633 (N_633,In_198,In_1937);
xnor U634 (N_634,In_2331,In_922);
or U635 (N_635,In_1721,In_563);
nor U636 (N_636,In_1487,In_452);
or U637 (N_637,In_1932,In_1488);
nand U638 (N_638,In_2237,In_538);
and U639 (N_639,In_2143,In_2459);
or U640 (N_640,In_1038,In_1629);
xnor U641 (N_641,In_236,In_2070);
nor U642 (N_642,In_1614,In_1685);
or U643 (N_643,In_1358,In_919);
nor U644 (N_644,In_2408,In_687);
or U645 (N_645,In_1612,In_1006);
or U646 (N_646,In_2238,In_944);
and U647 (N_647,In_1347,In_2318);
nand U648 (N_648,In_2351,In_129);
xnor U649 (N_649,In_737,In_461);
or U650 (N_650,In_163,In_99);
xnor U651 (N_651,In_2043,In_915);
or U652 (N_652,In_1457,In_2029);
or U653 (N_653,In_2186,In_2130);
xnor U654 (N_654,In_458,In_1748);
or U655 (N_655,In_2198,In_2363);
and U656 (N_656,In_2187,In_1758);
nor U657 (N_657,In_449,In_954);
nand U658 (N_658,In_762,In_2338);
nand U659 (N_659,In_1792,In_327);
and U660 (N_660,In_1628,In_520);
xnor U661 (N_661,In_167,In_1321);
nand U662 (N_662,In_653,In_2160);
nand U663 (N_663,In_1480,In_557);
or U664 (N_664,In_715,In_490);
xor U665 (N_665,In_512,In_683);
or U666 (N_666,In_626,In_1598);
and U667 (N_667,In_879,In_1238);
and U668 (N_668,In_1313,In_1662);
xnor U669 (N_669,In_1368,In_1389);
or U670 (N_670,In_1590,In_2335);
xor U671 (N_671,In_1210,In_2216);
and U672 (N_672,In_1786,In_1857);
xor U673 (N_673,In_537,In_248);
and U674 (N_674,In_877,In_1740);
and U675 (N_675,In_1270,In_114);
nor U676 (N_676,In_1976,In_2311);
nand U677 (N_677,In_300,In_1103);
nor U678 (N_678,In_885,In_176);
nand U679 (N_679,In_469,In_1905);
and U680 (N_680,In_652,In_1674);
nor U681 (N_681,In_1102,In_282);
xnor U682 (N_682,In_1784,In_835);
and U683 (N_683,In_115,In_1955);
or U684 (N_684,In_2467,In_2035);
and U685 (N_685,In_1406,In_2057);
nor U686 (N_686,In_223,In_2297);
nand U687 (N_687,In_2370,In_2438);
or U688 (N_688,In_306,In_973);
and U689 (N_689,In_1476,In_1400);
or U690 (N_690,In_1410,In_72);
xnor U691 (N_691,In_846,In_1123);
nor U692 (N_692,In_2420,In_1715);
and U693 (N_693,In_1012,In_815);
xnor U694 (N_694,In_232,In_685);
and U695 (N_695,In_2173,In_138);
and U696 (N_696,In_1139,In_933);
and U697 (N_697,In_1394,In_1988);
or U698 (N_698,In_2353,In_2341);
nor U699 (N_699,In_2373,In_2414);
and U700 (N_700,In_2097,In_1447);
or U701 (N_701,In_1826,In_308);
nor U702 (N_702,In_2211,In_2229);
xnor U703 (N_703,In_1848,In_160);
nand U704 (N_704,In_838,In_2226);
and U705 (N_705,In_776,In_889);
xnor U706 (N_706,In_2182,In_805);
nor U707 (N_707,In_2294,In_2329);
or U708 (N_708,In_769,In_1825);
nand U709 (N_709,In_1950,In_346);
and U710 (N_710,In_1933,In_1411);
nor U711 (N_711,In_410,In_1922);
nor U712 (N_712,In_1657,In_429);
nand U713 (N_713,In_182,In_1798);
xnor U714 (N_714,In_2041,In_1791);
nor U715 (N_715,In_1973,In_335);
nand U716 (N_716,In_2071,In_192);
nor U717 (N_717,In_1954,In_859);
xnor U718 (N_718,In_545,In_1162);
nand U719 (N_719,In_594,In_590);
nand U720 (N_720,In_1549,In_1380);
nand U721 (N_721,In_1089,In_1525);
nand U722 (N_722,In_1940,In_1125);
nor U723 (N_723,In_1309,In_865);
and U724 (N_724,In_732,In_240);
or U725 (N_725,In_2210,In_2113);
or U726 (N_726,In_636,In_1322);
xnor U727 (N_727,In_1226,In_106);
and U728 (N_728,In_1140,In_315);
and U729 (N_729,In_1946,In_2132);
nor U730 (N_730,In_355,In_2062);
or U731 (N_731,In_328,In_2350);
xnor U732 (N_732,In_120,In_692);
nor U733 (N_733,In_2063,In_294);
xnor U734 (N_734,In_1776,In_739);
or U735 (N_735,In_63,In_2379);
xor U736 (N_736,In_1057,In_668);
and U737 (N_737,In_1503,In_713);
xnor U738 (N_738,In_1537,In_2147);
nor U739 (N_739,In_2291,In_2299);
nand U740 (N_740,In_2039,In_2496);
or U741 (N_741,In_1708,In_244);
xor U742 (N_742,In_1768,In_463);
nand U743 (N_743,In_936,In_2443);
nand U744 (N_744,In_2149,In_518);
nand U745 (N_745,In_1148,In_1608);
or U746 (N_746,In_654,In_523);
nand U747 (N_747,In_1762,In_1805);
or U748 (N_748,In_1695,In_1189);
xor U749 (N_749,In_1117,In_1142);
or U750 (N_750,In_2021,In_2395);
or U751 (N_751,In_296,In_462);
xor U752 (N_752,In_811,In_575);
or U753 (N_753,In_1068,In_995);
xor U754 (N_754,In_696,In_887);
xor U755 (N_755,In_2388,In_927);
or U756 (N_756,In_1458,In_906);
or U757 (N_757,In_1022,In_795);
and U758 (N_758,In_2413,In_2156);
xnor U759 (N_759,In_1514,In_2264);
and U760 (N_760,In_704,In_1063);
nand U761 (N_761,In_233,In_1242);
nor U762 (N_762,In_875,In_505);
and U763 (N_763,In_347,In_1055);
nor U764 (N_764,In_1004,In_1127);
xor U765 (N_765,In_962,In_1823);
or U766 (N_766,In_142,In_1664);
nor U767 (N_767,In_2458,In_1866);
and U768 (N_768,In_425,In_1993);
xor U769 (N_769,In_1174,In_2450);
nand U770 (N_770,In_1484,In_957);
xor U771 (N_771,In_1036,In_1370);
xnor U772 (N_772,In_1935,In_728);
nor U773 (N_773,In_506,In_2153);
nor U774 (N_774,In_558,In_1959);
xor U775 (N_775,In_2282,In_231);
xnor U776 (N_776,In_640,In_1633);
or U777 (N_777,In_1043,In_2049);
xor U778 (N_778,In_1167,In_2307);
xnor U779 (N_779,In_1591,In_466);
or U780 (N_780,In_1747,In_445);
nand U781 (N_781,In_677,In_535);
xor U782 (N_782,In_473,In_1660);
xor U783 (N_783,In_1822,In_1310);
nand U784 (N_784,In_131,In_161);
and U785 (N_785,In_2026,In_761);
nand U786 (N_786,In_903,In_1409);
and U787 (N_787,In_1821,In_1157);
nor U788 (N_788,In_439,In_1510);
xor U789 (N_789,In_1834,In_2263);
or U790 (N_790,In_2268,In_2466);
xor U791 (N_791,In_2289,In_2475);
xnor U792 (N_792,In_1110,In_384);
and U793 (N_793,In_1361,In_801);
and U794 (N_794,In_299,In_1371);
xor U795 (N_795,In_479,In_2032);
nand U796 (N_796,In_1516,In_1912);
nor U797 (N_797,In_387,In_2460);
nand U798 (N_798,In_1638,In_1941);
nand U799 (N_799,In_2178,In_2488);
and U800 (N_800,In_1469,In_1868);
or U801 (N_801,In_385,In_165);
and U802 (N_802,In_100,In_1257);
and U803 (N_803,In_1034,In_446);
nand U804 (N_804,In_1052,In_79);
or U805 (N_805,In_1801,In_2045);
xnor U806 (N_806,In_2482,In_116);
nor U807 (N_807,In_344,In_1382);
nand U808 (N_808,In_1974,In_326);
nor U809 (N_809,In_1634,In_1945);
or U810 (N_810,In_1010,In_2118);
nand U811 (N_811,In_2247,In_342);
nand U812 (N_812,In_657,In_989);
nand U813 (N_813,In_1861,In_1075);
nor U814 (N_814,In_2218,In_2359);
or U815 (N_815,In_2396,In_777);
nand U816 (N_816,In_1482,In_2323);
nand U817 (N_817,In_516,In_1673);
nor U818 (N_818,In_2422,In_118);
xor U819 (N_819,In_317,In_1146);
xnor U820 (N_820,In_702,In_2281);
and U821 (N_821,In_967,In_64);
nor U822 (N_822,In_1743,In_399);
or U823 (N_823,In_1205,In_1880);
or U824 (N_824,In_1263,In_2286);
nor U825 (N_825,In_504,In_2498);
nor U826 (N_826,In_55,In_1501);
xnor U827 (N_827,In_1026,In_1796);
or U828 (N_828,In_229,In_44);
and U829 (N_829,In_2157,In_1249);
and U830 (N_830,In_2207,In_2205);
xnor U831 (N_831,In_1832,In_598);
and U832 (N_832,In_94,In_311);
and U833 (N_833,In_775,In_930);
or U834 (N_834,In_2399,In_956);
and U835 (N_835,In_1234,In_1847);
nor U836 (N_836,In_531,In_1390);
nor U837 (N_837,In_1901,In_1072);
nand U838 (N_838,In_2453,In_2377);
xnor U839 (N_839,In_1705,In_221);
and U840 (N_840,In_2060,In_542);
and U841 (N_841,In_935,In_2376);
and U842 (N_842,In_2319,In_2163);
nor U843 (N_843,In_555,In_611);
or U844 (N_844,In_1168,In_1697);
xor U845 (N_845,In_330,In_1891);
and U846 (N_846,In_2234,In_717);
xnor U847 (N_847,In_745,In_2321);
nand U848 (N_848,In_1794,In_1246);
xnor U849 (N_849,In_1104,In_1126);
nand U850 (N_850,In_488,In_415);
and U851 (N_851,In_362,In_2235);
nand U852 (N_852,In_764,In_1913);
nand U853 (N_853,In_424,In_2017);
nor U854 (N_854,In_59,In_2305);
and U855 (N_855,In_1143,In_1816);
nor U856 (N_856,In_1486,In_56);
or U857 (N_857,In_1975,In_1082);
xor U858 (N_858,In_1679,In_377);
and U859 (N_859,In_494,In_596);
xor U860 (N_860,In_451,In_276);
xnor U861 (N_861,In_250,In_207);
or U862 (N_862,In_283,In_534);
nor U863 (N_863,In_1045,In_1039);
or U864 (N_864,In_731,In_2245);
or U865 (N_865,In_76,In_482);
nand U866 (N_866,In_1631,In_1810);
nand U867 (N_867,In_153,In_1550);
nor U868 (N_868,In_1517,In_851);
xnor U869 (N_869,In_1990,In_159);
or U870 (N_870,In_1349,In_2054);
or U871 (N_871,In_798,In_1138);
nor U872 (N_872,In_1712,In_16);
nor U873 (N_873,In_77,In_2300);
and U874 (N_874,In_1297,In_917);
nor U875 (N_875,In_1160,In_1388);
nand U876 (N_876,In_1563,In_2327);
nor U877 (N_877,In_783,In_1363);
and U878 (N_878,In_104,In_195);
or U879 (N_879,In_1597,In_205);
xor U880 (N_880,In_1630,In_243);
xor U881 (N_881,In_119,In_2037);
nor U882 (N_882,In_360,In_202);
xnor U883 (N_883,In_1734,In_1526);
xnor U884 (N_884,In_2138,In_2165);
and U885 (N_885,In_2240,In_196);
or U886 (N_886,In_581,In_1005);
or U887 (N_887,In_1812,In_628);
or U888 (N_888,In_2233,In_93);
or U889 (N_889,In_758,In_650);
and U890 (N_890,In_2141,In_194);
nand U891 (N_891,In_1035,In_2009);
nor U892 (N_892,In_188,In_716);
nand U893 (N_893,In_2490,In_2417);
nor U894 (N_894,In_1609,In_212);
or U895 (N_895,In_1024,In_1876);
or U896 (N_896,In_376,In_1956);
and U897 (N_897,In_262,In_1260);
or U898 (N_898,In_1502,In_2098);
and U899 (N_899,In_222,In_750);
or U900 (N_900,In_98,In_1149);
nand U901 (N_901,In_1415,In_1317);
xnor U902 (N_902,In_1906,In_401);
or U903 (N_903,In_1206,In_1716);
or U904 (N_904,In_2274,In_1433);
nand U905 (N_905,In_1266,In_1744);
and U906 (N_906,In_1756,In_634);
or U907 (N_907,In_1081,In_11);
and U908 (N_908,In_1467,In_579);
xnor U909 (N_909,In_211,In_2030);
or U910 (N_910,In_1284,In_1879);
and U911 (N_911,In_457,In_662);
or U912 (N_912,In_1227,In_1897);
and U913 (N_913,In_1015,In_997);
xor U914 (N_914,In_703,In_754);
and U915 (N_915,In_1241,In_428);
or U916 (N_916,In_269,In_2075);
nor U917 (N_917,In_969,In_1427);
nand U918 (N_918,In_2090,In_1421);
or U919 (N_919,In_631,In_1377);
and U920 (N_920,In_1401,In_2081);
nor U921 (N_921,In_1703,In_1497);
nand U922 (N_922,In_1546,In_441);
xnor U923 (N_923,In_1274,In_101);
or U924 (N_924,In_2172,In_2393);
nand U925 (N_925,In_1179,In_1944);
or U926 (N_926,In_1659,In_1860);
nand U927 (N_927,In_2055,In_1924);
xor U928 (N_928,In_2352,In_774);
or U929 (N_929,In_2390,In_28);
nand U930 (N_930,In_1867,In_2375);
nand U931 (N_931,In_2131,In_968);
nor U932 (N_932,In_643,In_584);
or U933 (N_933,In_1295,In_2440);
nand U934 (N_934,In_1918,In_1278);
or U935 (N_935,In_1000,In_612);
xnor U936 (N_936,In_1376,In_1237);
xnor U937 (N_937,In_1843,In_780);
xor U938 (N_938,In_25,In_1258);
nor U939 (N_939,In_830,In_2101);
nor U940 (N_940,In_2083,In_2114);
and U941 (N_941,In_1607,In_1802);
or U942 (N_942,In_2074,In_1889);
nand U943 (N_943,In_2425,In_1449);
or U944 (N_944,In_1892,In_955);
or U945 (N_945,In_2116,In_421);
or U946 (N_946,In_1914,In_102);
and U947 (N_947,In_1639,In_975);
nand U948 (N_948,In_2200,In_356);
nor U949 (N_949,In_1283,In_225);
or U950 (N_950,In_2261,In_1468);
xnor U951 (N_951,In_416,In_1815);
nor U952 (N_952,In_178,In_1779);
nor U953 (N_953,In_2348,In_472);
nand U954 (N_954,In_837,In_994);
nand U955 (N_955,In_136,In_2411);
and U956 (N_956,In_1711,In_926);
xnor U957 (N_957,In_1268,In_2277);
and U958 (N_958,In_373,In_797);
or U959 (N_959,In_831,In_1021);
or U960 (N_960,In_2144,In_2428);
nand U961 (N_961,In_2121,In_2430);
and U962 (N_962,In_1121,In_1814);
or U963 (N_963,In_2166,In_348);
nand U964 (N_964,In_1865,In_825);
or U965 (N_965,In_191,In_1770);
or U966 (N_966,In_148,In_1300);
nand U967 (N_967,In_230,In_447);
xnor U968 (N_968,In_1175,In_536);
xor U969 (N_969,In_459,In_2337);
or U970 (N_970,In_1281,In_884);
xnor U971 (N_971,In_827,In_2220);
xor U972 (N_972,In_826,In_681);
or U973 (N_973,In_298,In_1981);
xnor U974 (N_974,In_2231,In_219);
nor U975 (N_975,In_228,In_890);
or U976 (N_976,In_592,In_1509);
xor U977 (N_977,In_1050,In_1087);
xnor U978 (N_978,In_549,In_187);
nand U979 (N_979,In_734,In_2023);
xor U980 (N_980,In_267,In_1155);
xor U981 (N_981,In_1733,In_215);
nand U982 (N_982,In_1759,In_633);
or U983 (N_983,In_1854,In_475);
or U984 (N_984,In_515,In_2284);
or U985 (N_985,In_1037,In_206);
and U986 (N_986,In_1923,In_199);
or U987 (N_987,In_1107,In_2256);
nor U988 (N_988,In_1886,In_258);
xor U989 (N_989,In_985,In_284);
and U990 (N_990,In_272,In_1594);
nand U991 (N_991,In_2416,In_1014);
xor U992 (N_992,In_1402,In_1265);
or U993 (N_993,In_1709,In_1524);
nand U994 (N_994,In_1364,In_1754);
or U995 (N_995,In_809,In_899);
xor U996 (N_996,In_394,In_1907);
and U997 (N_997,In_1699,In_24);
or U998 (N_998,In_478,In_130);
xor U999 (N_999,In_372,In_1819);
and U1000 (N_1000,In_2181,In_1908);
nor U1001 (N_1001,In_1948,In_888);
and U1002 (N_1002,In_1613,In_1769);
or U1003 (N_1003,In_2421,In_610);
and U1004 (N_1004,In_1399,In_1964);
nor U1005 (N_1005,In_1996,In_541);
and U1006 (N_1006,In_1687,In_1979);
xor U1007 (N_1007,In_1161,In_1204);
nand U1008 (N_1008,In_987,In_1171);
nand U1009 (N_1009,In_1288,In_1938);
or U1010 (N_1010,In_1644,In_1332);
or U1011 (N_1011,In_1145,In_2176);
and U1012 (N_1012,In_1830,In_1735);
nand U1013 (N_1013,In_950,In_1032);
and U1014 (N_1014,In_1749,In_519);
nor U1015 (N_1015,In_1131,In_1507);
and U1016 (N_1016,In_676,In_1771);
or U1017 (N_1017,In_2314,In_128);
xnor U1018 (N_1018,In_2398,In_1311);
nor U1019 (N_1019,In_481,In_2386);
xnor U1020 (N_1020,In_1323,In_2217);
xor U1021 (N_1021,In_600,In_2367);
and U1022 (N_1022,In_951,In_2404);
and U1023 (N_1023,In_1619,In_881);
xnor U1024 (N_1024,In_3,In_1498);
nand U1025 (N_1025,In_2115,In_723);
xnor U1026 (N_1026,In_1395,In_1312);
and U1027 (N_1027,In_1070,In_1201);
xnor U1028 (N_1028,In_670,In_367);
or U1029 (N_1029,In_1916,In_1253);
xor U1030 (N_1030,In_1446,In_1335);
and U1031 (N_1031,In_1686,In_1272);
or U1032 (N_1032,In_1943,In_567);
nand U1033 (N_1033,In_1547,In_2382);
nand U1034 (N_1034,In_2378,In_2491);
nand U1035 (N_1035,In_1153,In_393);
or U1036 (N_1036,In_2199,In_2397);
nand U1037 (N_1037,In_1453,In_1366);
xnor U1038 (N_1038,In_672,In_2472);
or U1039 (N_1039,In_1302,In_84);
nor U1040 (N_1040,In_844,In_574);
nand U1041 (N_1041,In_1391,In_2104);
nand U1042 (N_1042,In_252,In_74);
nor U1043 (N_1043,In_1170,In_1250);
or U1044 (N_1044,In_493,In_1003);
nor U1045 (N_1045,In_1197,In_18);
nor U1046 (N_1046,In_931,In_1824);
nor U1047 (N_1047,In_834,In_820);
and U1048 (N_1048,In_1957,In_66);
and U1049 (N_1049,In_418,In_1642);
or U1050 (N_1050,In_1985,In_984);
and U1051 (N_1051,In_1730,In_1298);
nand U1052 (N_1052,In_2016,In_1650);
and U1053 (N_1053,In_1404,In_297);
or U1054 (N_1054,In_521,In_1073);
or U1055 (N_1055,In_1894,In_2415);
nand U1056 (N_1056,In_1565,In_1330);
and U1057 (N_1057,In_1992,In_641);
and U1058 (N_1058,In_339,In_843);
and U1059 (N_1059,In_286,In_279);
or U1060 (N_1060,In_528,In_2246);
or U1061 (N_1061,In_2385,In_321);
xor U1062 (N_1062,In_2036,In_103);
or U1063 (N_1063,In_1491,In_454);
xor U1064 (N_1064,In_690,In_1911);
or U1065 (N_1065,In_2273,In_1435);
xnor U1066 (N_1066,In_343,In_2306);
or U1067 (N_1067,In_15,In_748);
and U1068 (N_1068,In_1047,In_1953);
and U1069 (N_1069,In_819,In_2126);
xnor U1070 (N_1070,In_2326,In_2111);
and U1071 (N_1071,In_109,In_904);
or U1072 (N_1072,In_117,In_349);
nand U1073 (N_1073,In_1583,In_1416);
or U1074 (N_1074,In_1423,In_624);
nand U1075 (N_1075,In_2089,In_522);
nand U1076 (N_1076,In_2148,In_1386);
nor U1077 (N_1077,In_183,In_1966);
and U1078 (N_1078,In_2332,In_808);
and U1079 (N_1079,In_1199,In_1356);
nand U1080 (N_1080,In_1374,In_695);
and U1081 (N_1081,In_2364,In_287);
nor U1082 (N_1082,In_144,In_901);
or U1083 (N_1083,In_1785,In_2225);
nand U1084 (N_1084,In_1900,In_991);
nor U1085 (N_1085,In_329,In_1437);
xnor U1086 (N_1086,In_2401,In_433);
xor U1087 (N_1087,In_1898,In_487);
nand U1088 (N_1088,In_164,In_147);
xnor U1089 (N_1089,In_2056,In_2179);
or U1090 (N_1090,In_751,In_1505);
nand U1091 (N_1091,In_170,In_1719);
nor U1092 (N_1092,In_1229,In_364);
nor U1093 (N_1093,In_1921,In_604);
nand U1094 (N_1094,In_7,In_2076);
nor U1095 (N_1095,In_309,In_1083);
xnor U1096 (N_1096,In_1008,In_1989);
xnor U1097 (N_1097,In_1667,In_880);
and U1098 (N_1098,In_2110,In_898);
nand U1099 (N_1099,In_2489,In_2125);
nor U1100 (N_1100,In_2112,In_2292);
nor U1101 (N_1101,In_2094,In_2008);
xnor U1102 (N_1102,In_878,In_341);
nor U1103 (N_1103,In_608,In_647);
nor U1104 (N_1104,In_1084,In_671);
or U1105 (N_1105,In_1269,In_1742);
nand U1106 (N_1106,In_1741,In_1116);
nand U1107 (N_1107,In_1430,In_60);
xnor U1108 (N_1108,In_431,In_778);
nand U1109 (N_1109,In_476,In_2328);
and U1110 (N_1110,In_1928,In_2487);
or U1111 (N_1111,In_872,In_2065);
nor U1112 (N_1112,In_485,In_2355);
xor U1113 (N_1113,In_302,In_50);
and U1114 (N_1114,In_1602,In_1542);
and U1115 (N_1115,In_2258,In_1624);
or U1116 (N_1116,In_943,In_949);
or U1117 (N_1117,In_47,In_370);
nor U1118 (N_1118,In_609,In_635);
nor U1119 (N_1119,In_1919,In_1354);
nor U1120 (N_1120,In_508,In_6);
nand U1121 (N_1121,In_1385,In_1341);
or U1122 (N_1122,In_1920,In_1279);
xor U1123 (N_1123,In_923,In_413);
xnor U1124 (N_1124,In_613,In_2257);
nand U1125 (N_1125,In_1420,In_746);
xnor U1126 (N_1126,In_2164,In_2485);
and U1127 (N_1127,In_1030,In_174);
nand U1128 (N_1128,In_659,In_1426);
nand U1129 (N_1129,In_854,In_2020);
and U1130 (N_1130,In_2058,In_1800);
nor U1131 (N_1131,In_171,In_30);
nor U1132 (N_1132,In_31,In_1251);
nor U1133 (N_1133,In_2095,In_791);
xnor U1134 (N_1134,In_1670,In_112);
xnor U1135 (N_1135,In_961,In_217);
nor U1136 (N_1136,In_2072,In_2451);
and U1137 (N_1137,In_1877,In_2346);
nor U1138 (N_1138,In_1397,In_2361);
nor U1139 (N_1139,In_1508,In_2145);
nor U1140 (N_1140,In_1788,In_1623);
or U1141 (N_1141,In_1438,In_2073);
nand U1142 (N_1142,In_1836,In_1963);
or U1143 (N_1143,In_500,In_1783);
xnor U1144 (N_1144,In_1691,In_13);
nor U1145 (N_1145,In_1717,In_19);
nand U1146 (N_1146,In_2204,In_32);
and U1147 (N_1147,In_179,In_1092);
nand U1148 (N_1148,In_786,In_1896);
and U1149 (N_1149,In_1441,In_2117);
nor U1150 (N_1150,In_2230,In_2079);
xor U1151 (N_1151,In_679,In_694);
nand U1152 (N_1152,In_1766,In_546);
nor U1153 (N_1153,In_398,In_1159);
or U1154 (N_1154,In_1980,In_92);
nor U1155 (N_1155,In_1077,In_1871);
nand U1156 (N_1156,In_1244,In_1093);
or U1157 (N_1157,In_870,In_1105);
xnor U1158 (N_1158,In_1797,In_1677);
nand U1159 (N_1159,In_1463,In_907);
nand U1160 (N_1160,In_559,In_122);
nor U1161 (N_1161,In_1141,In_569);
nand U1162 (N_1162,In_562,In_1114);
nand U1163 (N_1163,In_913,In_589);
nand U1164 (N_1164,In_1787,In_623);
nor U1165 (N_1165,In_422,In_1808);
xnor U1166 (N_1166,In_1700,In_1578);
nand U1167 (N_1167,In_599,In_2000);
and U1168 (N_1168,In_766,In_218);
and U1169 (N_1169,In_511,In_1147);
nor U1170 (N_1170,In_1863,In_1616);
xor U1171 (N_1171,In_617,In_1473);
xor U1172 (N_1172,In_135,In_2108);
xnor U1173 (N_1173,In_448,In_1418);
nand U1174 (N_1174,In_497,In_1661);
or U1175 (N_1175,In_2120,In_586);
xnor U1176 (N_1176,In_810,In_2283);
and U1177 (N_1177,In_620,In_2304);
and U1178 (N_1178,In_2105,In_514);
nand U1179 (N_1179,In_2219,In_1838);
nand U1180 (N_1180,In_947,In_806);
nand U1181 (N_1181,In_1978,In_1459);
and U1182 (N_1182,In_1999,In_1196);
or U1183 (N_1183,In_1028,In_1296);
or U1184 (N_1184,In_699,In_1327);
or U1185 (N_1185,In_474,In_1663);
xnor U1186 (N_1186,In_698,In_2455);
nor U1187 (N_1187,In_470,In_1062);
xnor U1188 (N_1188,In_1066,In_2195);
nand U1189 (N_1189,In_139,In_1984);
and U1190 (N_1190,In_1165,In_1654);
nor U1191 (N_1191,In_905,In_285);
nor U1192 (N_1192,In_237,In_787);
and U1193 (N_1193,In_2418,In_1173);
nor U1194 (N_1194,In_656,In_1233);
or U1195 (N_1195,In_852,In_1150);
or U1196 (N_1196,In_730,In_375);
nor U1197 (N_1197,In_241,In_1424);
xor U1198 (N_1198,In_352,In_1462);
nor U1199 (N_1199,In_911,In_2317);
or U1200 (N_1200,In_638,In_2232);
nor U1201 (N_1201,In_1190,In_779);
xor U1202 (N_1202,In_127,In_1495);
and U1203 (N_1203,In_772,In_36);
or U1204 (N_1204,In_1017,In_1211);
and U1205 (N_1205,In_1904,In_1407);
xnor U1206 (N_1206,In_2372,In_1656);
xor U1207 (N_1207,In_1645,In_268);
and U1208 (N_1208,In_896,In_1320);
nand U1209 (N_1209,In_1554,In_1198);
nand U1210 (N_1210,In_1336,In_1472);
nand U1211 (N_1211,In_483,In_637);
and U1212 (N_1212,In_1042,In_1878);
or U1213 (N_1213,In_465,In_2344);
and U1214 (N_1214,In_1414,In_2374);
and U1215 (N_1215,In_186,In_2369);
nor U1216 (N_1216,In_270,In_1752);
and U1217 (N_1217,In_455,In_220);
xor U1218 (N_1218,In_80,In_1256);
and U1219 (N_1219,In_389,In_2255);
nor U1220 (N_1220,In_277,In_2457);
nand U1221 (N_1221,In_781,In_2456);
nor U1222 (N_1222,In_1076,In_1239);
and U1223 (N_1223,In_1134,In_53);
xor U1224 (N_1224,In_1033,In_2254);
and U1225 (N_1225,In_861,In_2208);
and U1226 (N_1226,In_289,In_8);
xor U1227 (N_1227,In_976,In_1164);
nor U1228 (N_1228,In_1044,In_1308);
nand U1229 (N_1229,In_548,In_156);
or U1230 (N_1230,In_2434,In_1572);
or U1231 (N_1231,In_337,In_591);
and U1232 (N_1232,In_1464,In_873);
xnor U1233 (N_1233,In_618,In_388);
and U1234 (N_1234,In_839,In_1621);
nor U1235 (N_1235,In_1849,In_4);
and U1236 (N_1236,In_1951,In_2279);
nor U1237 (N_1237,In_403,In_107);
nand U1238 (N_1238,In_2406,In_582);
nand U1239 (N_1239,In_345,In_842);
nor U1240 (N_1240,In_1617,In_1936);
nor U1241 (N_1241,In_1163,In_1842);
or U1242 (N_1242,In_2280,In_1683);
nor U1243 (N_1243,In_2278,In_23);
nor U1244 (N_1244,In_82,In_2266);
nand U1245 (N_1245,In_181,In_1862);
nor U1246 (N_1246,In_1881,In_1355);
or U1247 (N_1247,In_1739,In_908);
nor U1248 (N_1248,In_1348,In_467);
and U1249 (N_1249,In_570,In_2298);
or U1250 (N_1250,In_1905,In_47);
xor U1251 (N_1251,In_1761,In_2401);
nor U1252 (N_1252,In_13,In_1597);
or U1253 (N_1253,In_874,In_264);
and U1254 (N_1254,In_1191,In_2351);
xor U1255 (N_1255,In_1639,In_1543);
and U1256 (N_1256,In_683,In_889);
xor U1257 (N_1257,In_1319,In_2116);
nand U1258 (N_1258,In_1185,In_967);
xor U1259 (N_1259,In_2246,In_195);
nand U1260 (N_1260,In_2055,In_2203);
xnor U1261 (N_1261,In_1092,In_2388);
and U1262 (N_1262,In_2028,In_1553);
nor U1263 (N_1263,In_469,In_1390);
xnor U1264 (N_1264,In_282,In_192);
nor U1265 (N_1265,In_1917,In_992);
xnor U1266 (N_1266,In_1148,In_453);
xnor U1267 (N_1267,In_637,In_2165);
nor U1268 (N_1268,In_847,In_905);
or U1269 (N_1269,In_1625,In_556);
or U1270 (N_1270,In_2134,In_1154);
nor U1271 (N_1271,In_2103,In_300);
nor U1272 (N_1272,In_1849,In_681);
or U1273 (N_1273,In_1806,In_1570);
or U1274 (N_1274,In_1921,In_1668);
xor U1275 (N_1275,In_279,In_2253);
and U1276 (N_1276,In_1614,In_1169);
and U1277 (N_1277,In_943,In_1011);
nor U1278 (N_1278,In_1098,In_640);
and U1279 (N_1279,In_1353,In_2244);
and U1280 (N_1280,In_720,In_289);
nor U1281 (N_1281,In_1564,In_1304);
xnor U1282 (N_1282,In_889,In_799);
nand U1283 (N_1283,In_1303,In_1443);
nor U1284 (N_1284,In_1768,In_195);
or U1285 (N_1285,In_1084,In_932);
nor U1286 (N_1286,In_186,In_893);
nand U1287 (N_1287,In_660,In_1893);
nor U1288 (N_1288,In_174,In_2206);
and U1289 (N_1289,In_2293,In_668);
nor U1290 (N_1290,In_2426,In_2092);
and U1291 (N_1291,In_588,In_1873);
and U1292 (N_1292,In_1017,In_1758);
or U1293 (N_1293,In_1593,In_973);
nor U1294 (N_1294,In_725,In_293);
nor U1295 (N_1295,In_636,In_736);
or U1296 (N_1296,In_483,In_119);
or U1297 (N_1297,In_1872,In_1452);
nand U1298 (N_1298,In_1025,In_243);
or U1299 (N_1299,In_2423,In_1402);
and U1300 (N_1300,In_122,In_933);
or U1301 (N_1301,In_824,In_1421);
nor U1302 (N_1302,In_2450,In_922);
nor U1303 (N_1303,In_1026,In_2229);
or U1304 (N_1304,In_1768,In_1925);
nor U1305 (N_1305,In_245,In_1234);
nor U1306 (N_1306,In_1418,In_299);
nor U1307 (N_1307,In_312,In_1113);
nand U1308 (N_1308,In_1434,In_819);
or U1309 (N_1309,In_694,In_624);
nand U1310 (N_1310,In_2369,In_2198);
nand U1311 (N_1311,In_146,In_2332);
xor U1312 (N_1312,In_1979,In_1147);
xor U1313 (N_1313,In_2204,In_102);
and U1314 (N_1314,In_1719,In_1121);
nor U1315 (N_1315,In_2024,In_1558);
or U1316 (N_1316,In_976,In_1904);
or U1317 (N_1317,In_1055,In_1620);
xor U1318 (N_1318,In_261,In_1717);
xnor U1319 (N_1319,In_1547,In_1382);
and U1320 (N_1320,In_1593,In_380);
or U1321 (N_1321,In_514,In_600);
nand U1322 (N_1322,In_578,In_1421);
nor U1323 (N_1323,In_183,In_1816);
nand U1324 (N_1324,In_339,In_508);
nor U1325 (N_1325,In_48,In_979);
nor U1326 (N_1326,In_2319,In_154);
xor U1327 (N_1327,In_1408,In_2290);
nand U1328 (N_1328,In_1356,In_1402);
or U1329 (N_1329,In_112,In_1786);
nor U1330 (N_1330,In_1947,In_481);
nand U1331 (N_1331,In_522,In_334);
or U1332 (N_1332,In_2219,In_182);
nor U1333 (N_1333,In_1015,In_423);
or U1334 (N_1334,In_411,In_559);
nor U1335 (N_1335,In_1839,In_83);
xnor U1336 (N_1336,In_298,In_714);
or U1337 (N_1337,In_1052,In_136);
xor U1338 (N_1338,In_1483,In_827);
or U1339 (N_1339,In_1899,In_1412);
and U1340 (N_1340,In_482,In_762);
nor U1341 (N_1341,In_2340,In_222);
nand U1342 (N_1342,In_939,In_777);
and U1343 (N_1343,In_2103,In_759);
or U1344 (N_1344,In_2397,In_464);
xnor U1345 (N_1345,In_556,In_1724);
nand U1346 (N_1346,In_796,In_777);
nand U1347 (N_1347,In_182,In_1339);
xnor U1348 (N_1348,In_1834,In_1543);
nand U1349 (N_1349,In_1159,In_1802);
nand U1350 (N_1350,In_1907,In_540);
nor U1351 (N_1351,In_1854,In_1545);
nand U1352 (N_1352,In_1520,In_1051);
and U1353 (N_1353,In_1249,In_1133);
or U1354 (N_1354,In_586,In_2007);
xor U1355 (N_1355,In_1878,In_1898);
or U1356 (N_1356,In_355,In_2382);
nand U1357 (N_1357,In_955,In_2246);
and U1358 (N_1358,In_2491,In_424);
xor U1359 (N_1359,In_29,In_24);
nor U1360 (N_1360,In_948,In_1615);
nand U1361 (N_1361,In_410,In_430);
xor U1362 (N_1362,In_178,In_2108);
nand U1363 (N_1363,In_411,In_2139);
and U1364 (N_1364,In_618,In_82);
xor U1365 (N_1365,In_1421,In_2079);
nand U1366 (N_1366,In_874,In_2114);
and U1367 (N_1367,In_310,In_272);
and U1368 (N_1368,In_135,In_183);
nor U1369 (N_1369,In_1511,In_2084);
and U1370 (N_1370,In_1547,In_1149);
nand U1371 (N_1371,In_2365,In_2426);
nand U1372 (N_1372,In_344,In_543);
or U1373 (N_1373,In_1894,In_123);
nand U1374 (N_1374,In_1675,In_810);
nand U1375 (N_1375,In_1267,In_2330);
or U1376 (N_1376,In_1487,In_897);
xor U1377 (N_1377,In_2217,In_1059);
xnor U1378 (N_1378,In_1839,In_1230);
nand U1379 (N_1379,In_186,In_2262);
and U1380 (N_1380,In_451,In_496);
nand U1381 (N_1381,In_1326,In_165);
or U1382 (N_1382,In_1718,In_1186);
or U1383 (N_1383,In_2275,In_1277);
xnor U1384 (N_1384,In_1716,In_1526);
nor U1385 (N_1385,In_151,In_1390);
xnor U1386 (N_1386,In_1686,In_2226);
xnor U1387 (N_1387,In_2492,In_1012);
nand U1388 (N_1388,In_930,In_1391);
xnor U1389 (N_1389,In_986,In_1619);
xnor U1390 (N_1390,In_114,In_1611);
and U1391 (N_1391,In_1518,In_1137);
and U1392 (N_1392,In_2079,In_1943);
xor U1393 (N_1393,In_1437,In_1542);
nand U1394 (N_1394,In_887,In_1088);
nor U1395 (N_1395,In_415,In_993);
xnor U1396 (N_1396,In_1450,In_2012);
xor U1397 (N_1397,In_994,In_2151);
nor U1398 (N_1398,In_1845,In_840);
and U1399 (N_1399,In_1517,In_393);
or U1400 (N_1400,In_1728,In_2335);
nand U1401 (N_1401,In_1869,In_1776);
nand U1402 (N_1402,In_1741,In_2018);
or U1403 (N_1403,In_620,In_1007);
or U1404 (N_1404,In_1922,In_1484);
xor U1405 (N_1405,In_326,In_2287);
xor U1406 (N_1406,In_1827,In_1869);
xnor U1407 (N_1407,In_2196,In_237);
or U1408 (N_1408,In_2008,In_2429);
nand U1409 (N_1409,In_1603,In_724);
nand U1410 (N_1410,In_2239,In_1410);
nor U1411 (N_1411,In_434,In_1689);
or U1412 (N_1412,In_1669,In_1637);
xnor U1413 (N_1413,In_598,In_1717);
and U1414 (N_1414,In_1251,In_359);
or U1415 (N_1415,In_1825,In_102);
nand U1416 (N_1416,In_1020,In_844);
nand U1417 (N_1417,In_374,In_756);
nor U1418 (N_1418,In_357,In_458);
xnor U1419 (N_1419,In_255,In_596);
xor U1420 (N_1420,In_1938,In_1081);
or U1421 (N_1421,In_2016,In_239);
xor U1422 (N_1422,In_2213,In_29);
or U1423 (N_1423,In_1000,In_2412);
nand U1424 (N_1424,In_2214,In_855);
nand U1425 (N_1425,In_90,In_1625);
xnor U1426 (N_1426,In_1903,In_1996);
or U1427 (N_1427,In_584,In_666);
and U1428 (N_1428,In_34,In_143);
or U1429 (N_1429,In_988,In_134);
nand U1430 (N_1430,In_30,In_1383);
or U1431 (N_1431,In_465,In_516);
xor U1432 (N_1432,In_820,In_2473);
or U1433 (N_1433,In_2160,In_1492);
and U1434 (N_1434,In_1252,In_1751);
and U1435 (N_1435,In_566,In_2498);
or U1436 (N_1436,In_824,In_1547);
and U1437 (N_1437,In_755,In_463);
or U1438 (N_1438,In_1667,In_2468);
xor U1439 (N_1439,In_2235,In_1927);
nor U1440 (N_1440,In_1077,In_2392);
nand U1441 (N_1441,In_1830,In_1345);
xor U1442 (N_1442,In_2049,In_2493);
nor U1443 (N_1443,In_1014,In_2159);
xnor U1444 (N_1444,In_1737,In_342);
or U1445 (N_1445,In_1521,In_308);
xor U1446 (N_1446,In_933,In_1127);
nor U1447 (N_1447,In_1309,In_1264);
and U1448 (N_1448,In_471,In_1363);
and U1449 (N_1449,In_984,In_477);
and U1450 (N_1450,In_1448,In_2108);
nor U1451 (N_1451,In_2436,In_1458);
and U1452 (N_1452,In_2032,In_724);
xnor U1453 (N_1453,In_301,In_952);
or U1454 (N_1454,In_1396,In_1224);
or U1455 (N_1455,In_734,In_1197);
or U1456 (N_1456,In_1862,In_1575);
xor U1457 (N_1457,In_2171,In_2452);
or U1458 (N_1458,In_1185,In_1478);
xnor U1459 (N_1459,In_1201,In_1583);
nor U1460 (N_1460,In_2347,In_1958);
or U1461 (N_1461,In_689,In_763);
or U1462 (N_1462,In_999,In_2384);
xnor U1463 (N_1463,In_354,In_2429);
xnor U1464 (N_1464,In_296,In_836);
nand U1465 (N_1465,In_1252,In_1242);
xnor U1466 (N_1466,In_1395,In_779);
nand U1467 (N_1467,In_197,In_263);
and U1468 (N_1468,In_1948,In_1074);
or U1469 (N_1469,In_1616,In_1416);
or U1470 (N_1470,In_1830,In_1613);
xnor U1471 (N_1471,In_921,In_1034);
nor U1472 (N_1472,In_640,In_2487);
nand U1473 (N_1473,In_109,In_322);
and U1474 (N_1474,In_2351,In_282);
nor U1475 (N_1475,In_2364,In_1093);
nand U1476 (N_1476,In_727,In_162);
and U1477 (N_1477,In_338,In_1389);
and U1478 (N_1478,In_478,In_1839);
or U1479 (N_1479,In_763,In_779);
or U1480 (N_1480,In_1756,In_2012);
and U1481 (N_1481,In_2106,In_608);
nor U1482 (N_1482,In_51,In_2253);
and U1483 (N_1483,In_1727,In_2096);
nor U1484 (N_1484,In_2042,In_31);
nand U1485 (N_1485,In_1423,In_1970);
nor U1486 (N_1486,In_2211,In_1233);
and U1487 (N_1487,In_621,In_746);
xnor U1488 (N_1488,In_1273,In_1639);
or U1489 (N_1489,In_1868,In_1306);
and U1490 (N_1490,In_2497,In_2429);
xor U1491 (N_1491,In_265,In_1354);
nor U1492 (N_1492,In_152,In_525);
and U1493 (N_1493,In_963,In_2132);
xor U1494 (N_1494,In_2248,In_781);
nor U1495 (N_1495,In_768,In_744);
nand U1496 (N_1496,In_422,In_2150);
or U1497 (N_1497,In_1822,In_105);
and U1498 (N_1498,In_2094,In_376);
or U1499 (N_1499,In_382,In_554);
nor U1500 (N_1500,In_1741,In_1515);
or U1501 (N_1501,In_2128,In_919);
nor U1502 (N_1502,In_435,In_51);
and U1503 (N_1503,In_1133,In_202);
and U1504 (N_1504,In_399,In_2334);
or U1505 (N_1505,In_1843,In_2077);
xor U1506 (N_1506,In_543,In_274);
xnor U1507 (N_1507,In_1161,In_350);
xnor U1508 (N_1508,In_1412,In_1085);
nand U1509 (N_1509,In_301,In_2402);
and U1510 (N_1510,In_1015,In_1379);
nor U1511 (N_1511,In_1304,In_426);
xnor U1512 (N_1512,In_221,In_2047);
and U1513 (N_1513,In_2032,In_976);
or U1514 (N_1514,In_1826,In_1283);
nand U1515 (N_1515,In_926,In_1188);
and U1516 (N_1516,In_420,In_2234);
nor U1517 (N_1517,In_442,In_746);
xnor U1518 (N_1518,In_449,In_418);
nor U1519 (N_1519,In_1349,In_271);
and U1520 (N_1520,In_206,In_4);
or U1521 (N_1521,In_2121,In_1751);
or U1522 (N_1522,In_219,In_626);
and U1523 (N_1523,In_470,In_935);
or U1524 (N_1524,In_1877,In_578);
nand U1525 (N_1525,In_345,In_1980);
xnor U1526 (N_1526,In_930,In_1887);
nand U1527 (N_1527,In_727,In_2419);
xnor U1528 (N_1528,In_1792,In_1116);
xor U1529 (N_1529,In_1904,In_1584);
or U1530 (N_1530,In_48,In_1828);
nand U1531 (N_1531,In_37,In_648);
xor U1532 (N_1532,In_2289,In_810);
and U1533 (N_1533,In_2221,In_2372);
and U1534 (N_1534,In_1296,In_1074);
and U1535 (N_1535,In_13,In_765);
or U1536 (N_1536,In_686,In_2239);
nor U1537 (N_1537,In_720,In_2453);
nor U1538 (N_1538,In_1777,In_2243);
nand U1539 (N_1539,In_1784,In_1414);
nand U1540 (N_1540,In_686,In_1012);
nand U1541 (N_1541,In_2060,In_465);
and U1542 (N_1542,In_1531,In_962);
nand U1543 (N_1543,In_1999,In_2305);
nor U1544 (N_1544,In_1326,In_474);
xor U1545 (N_1545,In_24,In_264);
nand U1546 (N_1546,In_1070,In_2477);
nor U1547 (N_1547,In_2428,In_715);
nand U1548 (N_1548,In_277,In_2374);
or U1549 (N_1549,In_112,In_2200);
xnor U1550 (N_1550,In_1683,In_1697);
xor U1551 (N_1551,In_1486,In_1091);
xor U1552 (N_1552,In_2353,In_2132);
nor U1553 (N_1553,In_1107,In_358);
or U1554 (N_1554,In_1369,In_1636);
and U1555 (N_1555,In_1975,In_2045);
or U1556 (N_1556,In_2137,In_847);
nor U1557 (N_1557,In_1657,In_1588);
nand U1558 (N_1558,In_864,In_1181);
and U1559 (N_1559,In_2411,In_889);
nor U1560 (N_1560,In_2357,In_57);
or U1561 (N_1561,In_1236,In_2310);
and U1562 (N_1562,In_2208,In_418);
or U1563 (N_1563,In_471,In_826);
nand U1564 (N_1564,In_2147,In_1472);
xnor U1565 (N_1565,In_1328,In_2067);
xor U1566 (N_1566,In_1168,In_1252);
and U1567 (N_1567,In_966,In_157);
or U1568 (N_1568,In_2205,In_2061);
nand U1569 (N_1569,In_2418,In_2382);
xnor U1570 (N_1570,In_201,In_312);
xnor U1571 (N_1571,In_1187,In_1832);
xor U1572 (N_1572,In_2359,In_219);
nor U1573 (N_1573,In_1159,In_1925);
or U1574 (N_1574,In_2230,In_2433);
xnor U1575 (N_1575,In_2451,In_1621);
xor U1576 (N_1576,In_1374,In_194);
nand U1577 (N_1577,In_690,In_2021);
nor U1578 (N_1578,In_1,In_1168);
and U1579 (N_1579,In_2289,In_1264);
or U1580 (N_1580,In_1282,In_840);
and U1581 (N_1581,In_451,In_2448);
or U1582 (N_1582,In_1880,In_1048);
or U1583 (N_1583,In_2385,In_1129);
and U1584 (N_1584,In_2427,In_2391);
xor U1585 (N_1585,In_1993,In_356);
or U1586 (N_1586,In_1726,In_2351);
and U1587 (N_1587,In_1231,In_1319);
xnor U1588 (N_1588,In_1201,In_2015);
and U1589 (N_1589,In_492,In_659);
nand U1590 (N_1590,In_195,In_178);
or U1591 (N_1591,In_788,In_1193);
xnor U1592 (N_1592,In_1720,In_457);
xnor U1593 (N_1593,In_836,In_1795);
nor U1594 (N_1594,In_1913,In_1675);
and U1595 (N_1595,In_1744,In_2048);
nor U1596 (N_1596,In_1207,In_1903);
xor U1597 (N_1597,In_1101,In_1994);
xor U1598 (N_1598,In_1486,In_599);
nor U1599 (N_1599,In_849,In_332);
and U1600 (N_1600,In_1074,In_1336);
xor U1601 (N_1601,In_2494,In_2487);
nand U1602 (N_1602,In_1733,In_187);
nand U1603 (N_1603,In_598,In_2328);
and U1604 (N_1604,In_977,In_506);
xnor U1605 (N_1605,In_1949,In_1754);
or U1606 (N_1606,In_589,In_127);
and U1607 (N_1607,In_1304,In_1354);
nand U1608 (N_1608,In_1850,In_491);
nor U1609 (N_1609,In_1444,In_1419);
nand U1610 (N_1610,In_2340,In_1019);
nand U1611 (N_1611,In_1644,In_1069);
nor U1612 (N_1612,In_828,In_2365);
nor U1613 (N_1613,In_1550,In_1773);
xor U1614 (N_1614,In_1559,In_1084);
and U1615 (N_1615,In_1002,In_2322);
or U1616 (N_1616,In_871,In_1645);
and U1617 (N_1617,In_2179,In_972);
and U1618 (N_1618,In_652,In_1523);
nor U1619 (N_1619,In_1362,In_968);
nand U1620 (N_1620,In_1045,In_1789);
nor U1621 (N_1621,In_511,In_1226);
or U1622 (N_1622,In_152,In_450);
xor U1623 (N_1623,In_579,In_2048);
or U1624 (N_1624,In_515,In_607);
and U1625 (N_1625,In_1266,In_342);
or U1626 (N_1626,In_1975,In_1436);
nand U1627 (N_1627,In_942,In_789);
and U1628 (N_1628,In_503,In_1137);
nor U1629 (N_1629,In_342,In_1787);
and U1630 (N_1630,In_634,In_2047);
nor U1631 (N_1631,In_928,In_500);
nor U1632 (N_1632,In_589,In_417);
or U1633 (N_1633,In_1213,In_360);
xnor U1634 (N_1634,In_2294,In_1638);
and U1635 (N_1635,In_282,In_346);
xor U1636 (N_1636,In_1794,In_798);
nor U1637 (N_1637,In_2090,In_1445);
and U1638 (N_1638,In_1156,In_1281);
and U1639 (N_1639,In_1875,In_58);
xnor U1640 (N_1640,In_1834,In_27);
and U1641 (N_1641,In_1934,In_1733);
nor U1642 (N_1642,In_2078,In_2462);
nor U1643 (N_1643,In_659,In_329);
or U1644 (N_1644,In_1172,In_2331);
nor U1645 (N_1645,In_761,In_2455);
nand U1646 (N_1646,In_1076,In_665);
nand U1647 (N_1647,In_335,In_1123);
xnor U1648 (N_1648,In_1150,In_1161);
and U1649 (N_1649,In_1693,In_1650);
and U1650 (N_1650,In_1866,In_288);
and U1651 (N_1651,In_141,In_1018);
nor U1652 (N_1652,In_1286,In_2079);
nor U1653 (N_1653,In_644,In_1298);
nor U1654 (N_1654,In_576,In_512);
nor U1655 (N_1655,In_1575,In_2285);
or U1656 (N_1656,In_132,In_2125);
or U1657 (N_1657,In_789,In_316);
xor U1658 (N_1658,In_1502,In_1639);
xnor U1659 (N_1659,In_1051,In_888);
nand U1660 (N_1660,In_873,In_1982);
xor U1661 (N_1661,In_587,In_1189);
and U1662 (N_1662,In_361,In_1190);
nor U1663 (N_1663,In_112,In_1354);
nor U1664 (N_1664,In_1706,In_279);
nor U1665 (N_1665,In_1617,In_1881);
or U1666 (N_1666,In_1562,In_294);
or U1667 (N_1667,In_459,In_13);
xor U1668 (N_1668,In_2428,In_1644);
and U1669 (N_1669,In_668,In_961);
and U1670 (N_1670,In_272,In_1435);
or U1671 (N_1671,In_1114,In_802);
nor U1672 (N_1672,In_2288,In_1069);
xnor U1673 (N_1673,In_837,In_839);
or U1674 (N_1674,In_1147,In_814);
or U1675 (N_1675,In_2288,In_299);
nand U1676 (N_1676,In_358,In_277);
xnor U1677 (N_1677,In_789,In_2361);
and U1678 (N_1678,In_504,In_60);
and U1679 (N_1679,In_1033,In_2450);
xor U1680 (N_1680,In_903,In_550);
and U1681 (N_1681,In_1346,In_955);
nor U1682 (N_1682,In_973,In_1795);
nand U1683 (N_1683,In_1575,In_649);
xor U1684 (N_1684,In_792,In_1730);
and U1685 (N_1685,In_840,In_1981);
nand U1686 (N_1686,In_971,In_1436);
nand U1687 (N_1687,In_1709,In_1537);
xor U1688 (N_1688,In_1854,In_1186);
nand U1689 (N_1689,In_1479,In_177);
nor U1690 (N_1690,In_1857,In_538);
nor U1691 (N_1691,In_1166,In_912);
nand U1692 (N_1692,In_921,In_2126);
nor U1693 (N_1693,In_1452,In_1667);
nor U1694 (N_1694,In_2249,In_2177);
xor U1695 (N_1695,In_623,In_2161);
nand U1696 (N_1696,In_2303,In_924);
nor U1697 (N_1697,In_745,In_2493);
nand U1698 (N_1698,In_711,In_1311);
nor U1699 (N_1699,In_1759,In_2142);
or U1700 (N_1700,In_1964,In_2112);
and U1701 (N_1701,In_643,In_2360);
and U1702 (N_1702,In_2312,In_480);
and U1703 (N_1703,In_1386,In_1842);
and U1704 (N_1704,In_1456,In_2183);
or U1705 (N_1705,In_1542,In_2209);
or U1706 (N_1706,In_1784,In_2301);
and U1707 (N_1707,In_1282,In_23);
nand U1708 (N_1708,In_2115,In_82);
or U1709 (N_1709,In_1379,In_804);
xnor U1710 (N_1710,In_2037,In_2408);
nand U1711 (N_1711,In_1681,In_87);
or U1712 (N_1712,In_330,In_586);
nand U1713 (N_1713,In_1781,In_334);
nor U1714 (N_1714,In_1268,In_297);
nor U1715 (N_1715,In_1603,In_2312);
or U1716 (N_1716,In_1779,In_577);
xnor U1717 (N_1717,In_2212,In_940);
or U1718 (N_1718,In_224,In_569);
or U1719 (N_1719,In_1152,In_1347);
nand U1720 (N_1720,In_1763,In_345);
xnor U1721 (N_1721,In_1154,In_1626);
nand U1722 (N_1722,In_458,In_1333);
nand U1723 (N_1723,In_346,In_666);
and U1724 (N_1724,In_1239,In_412);
xnor U1725 (N_1725,In_871,In_1385);
xor U1726 (N_1726,In_1882,In_2234);
nand U1727 (N_1727,In_1413,In_786);
xor U1728 (N_1728,In_1278,In_132);
xor U1729 (N_1729,In_2462,In_442);
xor U1730 (N_1730,In_1232,In_1887);
nand U1731 (N_1731,In_1761,In_507);
and U1732 (N_1732,In_583,In_242);
xnor U1733 (N_1733,In_564,In_2100);
nand U1734 (N_1734,In_42,In_697);
nand U1735 (N_1735,In_204,In_1757);
or U1736 (N_1736,In_693,In_224);
xnor U1737 (N_1737,In_2223,In_1759);
and U1738 (N_1738,In_1300,In_921);
and U1739 (N_1739,In_229,In_566);
nand U1740 (N_1740,In_1288,In_667);
or U1741 (N_1741,In_1266,In_176);
nand U1742 (N_1742,In_32,In_1242);
and U1743 (N_1743,In_2083,In_971);
and U1744 (N_1744,In_1308,In_258);
and U1745 (N_1745,In_1828,In_1327);
xnor U1746 (N_1746,In_416,In_515);
nand U1747 (N_1747,In_1872,In_1574);
nor U1748 (N_1748,In_1299,In_296);
or U1749 (N_1749,In_1187,In_1030);
and U1750 (N_1750,In_1883,In_2083);
nor U1751 (N_1751,In_693,In_1360);
and U1752 (N_1752,In_1180,In_1050);
nand U1753 (N_1753,In_589,In_386);
and U1754 (N_1754,In_396,In_1626);
or U1755 (N_1755,In_1829,In_908);
nand U1756 (N_1756,In_1016,In_108);
xor U1757 (N_1757,In_350,In_736);
nand U1758 (N_1758,In_1952,In_2491);
nand U1759 (N_1759,In_2229,In_829);
nor U1760 (N_1760,In_2478,In_2310);
nand U1761 (N_1761,In_1279,In_2370);
or U1762 (N_1762,In_890,In_682);
nand U1763 (N_1763,In_584,In_1801);
or U1764 (N_1764,In_23,In_1140);
nand U1765 (N_1765,In_2384,In_2436);
xor U1766 (N_1766,In_516,In_2332);
nand U1767 (N_1767,In_43,In_1049);
nor U1768 (N_1768,In_1201,In_1362);
and U1769 (N_1769,In_1574,In_2061);
and U1770 (N_1770,In_512,In_2019);
xor U1771 (N_1771,In_1055,In_1037);
or U1772 (N_1772,In_2130,In_720);
xnor U1773 (N_1773,In_439,In_1419);
nand U1774 (N_1774,In_1612,In_957);
nand U1775 (N_1775,In_1423,In_252);
and U1776 (N_1776,In_415,In_1654);
or U1777 (N_1777,In_2364,In_1361);
or U1778 (N_1778,In_272,In_2271);
or U1779 (N_1779,In_6,In_178);
or U1780 (N_1780,In_1426,In_1203);
nor U1781 (N_1781,In_20,In_140);
or U1782 (N_1782,In_1350,In_1582);
or U1783 (N_1783,In_780,In_1974);
nor U1784 (N_1784,In_1806,In_387);
nand U1785 (N_1785,In_422,In_1017);
or U1786 (N_1786,In_2324,In_262);
and U1787 (N_1787,In_298,In_1762);
xnor U1788 (N_1788,In_2302,In_2318);
nor U1789 (N_1789,In_2344,In_2368);
xnor U1790 (N_1790,In_1797,In_918);
and U1791 (N_1791,In_1053,In_330);
xor U1792 (N_1792,In_1443,In_2247);
nor U1793 (N_1793,In_226,In_1029);
xor U1794 (N_1794,In_1733,In_1665);
xnor U1795 (N_1795,In_566,In_609);
nand U1796 (N_1796,In_2192,In_1938);
and U1797 (N_1797,In_1233,In_990);
and U1798 (N_1798,In_850,In_390);
and U1799 (N_1799,In_2217,In_2270);
xnor U1800 (N_1800,In_115,In_418);
or U1801 (N_1801,In_2032,In_917);
nand U1802 (N_1802,In_370,In_1203);
and U1803 (N_1803,In_1833,In_2368);
and U1804 (N_1804,In_257,In_2171);
nand U1805 (N_1805,In_1851,In_701);
and U1806 (N_1806,In_40,In_897);
xnor U1807 (N_1807,In_840,In_735);
nor U1808 (N_1808,In_2004,In_2308);
and U1809 (N_1809,In_721,In_1272);
xor U1810 (N_1810,In_854,In_484);
nand U1811 (N_1811,In_101,In_950);
xor U1812 (N_1812,In_993,In_766);
and U1813 (N_1813,In_672,In_1376);
nor U1814 (N_1814,In_189,In_2185);
nand U1815 (N_1815,In_1220,In_2);
nand U1816 (N_1816,In_1822,In_2124);
nand U1817 (N_1817,In_58,In_1264);
and U1818 (N_1818,In_1298,In_1592);
xnor U1819 (N_1819,In_2339,In_1936);
nand U1820 (N_1820,In_1707,In_2417);
and U1821 (N_1821,In_456,In_1026);
and U1822 (N_1822,In_733,In_160);
nand U1823 (N_1823,In_2414,In_2179);
nor U1824 (N_1824,In_31,In_1282);
nor U1825 (N_1825,In_2017,In_2466);
nor U1826 (N_1826,In_600,In_1042);
xor U1827 (N_1827,In_2198,In_1960);
nand U1828 (N_1828,In_1023,In_1523);
and U1829 (N_1829,In_2275,In_747);
and U1830 (N_1830,In_2249,In_1589);
xor U1831 (N_1831,In_828,In_523);
and U1832 (N_1832,In_2064,In_1140);
or U1833 (N_1833,In_1825,In_1589);
nor U1834 (N_1834,In_741,In_1820);
and U1835 (N_1835,In_1992,In_2467);
nor U1836 (N_1836,In_190,In_1463);
or U1837 (N_1837,In_693,In_1216);
nor U1838 (N_1838,In_1060,In_1624);
xnor U1839 (N_1839,In_2269,In_409);
nor U1840 (N_1840,In_2121,In_2008);
nand U1841 (N_1841,In_1612,In_1229);
xor U1842 (N_1842,In_1235,In_1246);
and U1843 (N_1843,In_1191,In_1139);
nor U1844 (N_1844,In_1495,In_885);
nor U1845 (N_1845,In_344,In_1109);
or U1846 (N_1846,In_2323,In_523);
nand U1847 (N_1847,In_2061,In_2316);
and U1848 (N_1848,In_1501,In_2075);
xnor U1849 (N_1849,In_1785,In_1080);
nor U1850 (N_1850,In_1152,In_394);
nor U1851 (N_1851,In_2431,In_470);
xnor U1852 (N_1852,In_1013,In_1626);
or U1853 (N_1853,In_380,In_1508);
nor U1854 (N_1854,In_2295,In_1086);
nand U1855 (N_1855,In_2098,In_2024);
and U1856 (N_1856,In_179,In_198);
nand U1857 (N_1857,In_585,In_1589);
xor U1858 (N_1858,In_2117,In_2375);
nand U1859 (N_1859,In_874,In_162);
xnor U1860 (N_1860,In_1150,In_1276);
nor U1861 (N_1861,In_521,In_2480);
nor U1862 (N_1862,In_1391,In_1904);
nor U1863 (N_1863,In_128,In_662);
or U1864 (N_1864,In_1297,In_172);
nand U1865 (N_1865,In_2319,In_2413);
and U1866 (N_1866,In_1075,In_2156);
or U1867 (N_1867,In_1595,In_567);
or U1868 (N_1868,In_1683,In_1578);
xnor U1869 (N_1869,In_1154,In_1296);
or U1870 (N_1870,In_102,In_2020);
nand U1871 (N_1871,In_615,In_26);
xor U1872 (N_1872,In_2373,In_1004);
nand U1873 (N_1873,In_1779,In_1534);
and U1874 (N_1874,In_235,In_416);
xnor U1875 (N_1875,In_773,In_1150);
nor U1876 (N_1876,In_1040,In_1801);
or U1877 (N_1877,In_1541,In_132);
or U1878 (N_1878,In_248,In_252);
nand U1879 (N_1879,In_899,In_2322);
nor U1880 (N_1880,In_745,In_1395);
xnor U1881 (N_1881,In_201,In_1203);
nor U1882 (N_1882,In_2388,In_552);
or U1883 (N_1883,In_2303,In_2094);
and U1884 (N_1884,In_355,In_2409);
xnor U1885 (N_1885,In_1483,In_798);
and U1886 (N_1886,In_859,In_2490);
and U1887 (N_1887,In_1984,In_178);
xor U1888 (N_1888,In_1813,In_2233);
nor U1889 (N_1889,In_355,In_1634);
and U1890 (N_1890,In_1406,In_454);
xor U1891 (N_1891,In_124,In_1324);
nor U1892 (N_1892,In_1952,In_705);
and U1893 (N_1893,In_1549,In_539);
xor U1894 (N_1894,In_2249,In_1740);
nor U1895 (N_1895,In_48,In_1301);
nor U1896 (N_1896,In_1118,In_952);
xnor U1897 (N_1897,In_1038,In_1568);
xnor U1898 (N_1898,In_658,In_2367);
and U1899 (N_1899,In_2181,In_1972);
nor U1900 (N_1900,In_1299,In_388);
and U1901 (N_1901,In_2041,In_139);
nor U1902 (N_1902,In_1475,In_2401);
and U1903 (N_1903,In_2410,In_297);
xor U1904 (N_1904,In_1570,In_66);
nor U1905 (N_1905,In_1263,In_1095);
nor U1906 (N_1906,In_605,In_517);
xor U1907 (N_1907,In_614,In_813);
nand U1908 (N_1908,In_1812,In_361);
or U1909 (N_1909,In_191,In_2428);
nand U1910 (N_1910,In_2121,In_1307);
xor U1911 (N_1911,In_2442,In_1264);
and U1912 (N_1912,In_1228,In_2083);
or U1913 (N_1913,In_1773,In_2105);
nor U1914 (N_1914,In_1921,In_1362);
or U1915 (N_1915,In_2410,In_2139);
nor U1916 (N_1916,In_1479,In_1009);
nand U1917 (N_1917,In_720,In_787);
and U1918 (N_1918,In_1987,In_535);
nor U1919 (N_1919,In_1204,In_729);
or U1920 (N_1920,In_74,In_33);
xnor U1921 (N_1921,In_864,In_1483);
or U1922 (N_1922,In_2447,In_2236);
nand U1923 (N_1923,In_954,In_2250);
nand U1924 (N_1924,In_579,In_2059);
and U1925 (N_1925,In_1251,In_908);
xnor U1926 (N_1926,In_1288,In_403);
nand U1927 (N_1927,In_478,In_2020);
nand U1928 (N_1928,In_333,In_1722);
or U1929 (N_1929,In_1657,In_625);
xor U1930 (N_1930,In_1173,In_1695);
xor U1931 (N_1931,In_1804,In_2239);
and U1932 (N_1932,In_783,In_205);
nand U1933 (N_1933,In_1756,In_1619);
nor U1934 (N_1934,In_244,In_859);
and U1935 (N_1935,In_250,In_1779);
xor U1936 (N_1936,In_2306,In_1478);
or U1937 (N_1937,In_1037,In_1809);
nand U1938 (N_1938,In_897,In_2461);
xnor U1939 (N_1939,In_2172,In_1336);
nor U1940 (N_1940,In_1230,In_2279);
xnor U1941 (N_1941,In_2097,In_2453);
xor U1942 (N_1942,In_1937,In_2059);
or U1943 (N_1943,In_1387,In_1768);
or U1944 (N_1944,In_2377,In_806);
xnor U1945 (N_1945,In_107,In_1419);
or U1946 (N_1946,In_475,In_1972);
or U1947 (N_1947,In_1445,In_1033);
nor U1948 (N_1948,In_1652,In_1350);
xnor U1949 (N_1949,In_760,In_2243);
xnor U1950 (N_1950,In_118,In_2308);
or U1951 (N_1951,In_581,In_11);
nand U1952 (N_1952,In_145,In_1319);
nor U1953 (N_1953,In_1002,In_1455);
nand U1954 (N_1954,In_1776,In_712);
nand U1955 (N_1955,In_330,In_728);
nand U1956 (N_1956,In_2055,In_23);
xor U1957 (N_1957,In_1953,In_980);
and U1958 (N_1958,In_101,In_1796);
and U1959 (N_1959,In_2112,In_1873);
nor U1960 (N_1960,In_1538,In_717);
nor U1961 (N_1961,In_2006,In_134);
and U1962 (N_1962,In_591,In_518);
xor U1963 (N_1963,In_2095,In_1589);
nand U1964 (N_1964,In_980,In_2497);
xor U1965 (N_1965,In_122,In_1709);
xnor U1966 (N_1966,In_1268,In_1920);
nand U1967 (N_1967,In_1904,In_1836);
or U1968 (N_1968,In_949,In_98);
and U1969 (N_1969,In_1367,In_322);
and U1970 (N_1970,In_510,In_2433);
nor U1971 (N_1971,In_1306,In_252);
and U1972 (N_1972,In_692,In_1182);
xnor U1973 (N_1973,In_11,In_903);
nor U1974 (N_1974,In_778,In_579);
nor U1975 (N_1975,In_487,In_1787);
nand U1976 (N_1976,In_276,In_1216);
xor U1977 (N_1977,In_1222,In_1583);
and U1978 (N_1978,In_2263,In_145);
xor U1979 (N_1979,In_2028,In_2144);
xor U1980 (N_1980,In_2098,In_1386);
or U1981 (N_1981,In_1592,In_2222);
xnor U1982 (N_1982,In_515,In_1165);
xnor U1983 (N_1983,In_2108,In_2163);
or U1984 (N_1984,In_1743,In_2451);
or U1985 (N_1985,In_1291,In_751);
nor U1986 (N_1986,In_966,In_612);
nand U1987 (N_1987,In_360,In_1236);
nand U1988 (N_1988,In_1364,In_975);
or U1989 (N_1989,In_1475,In_960);
or U1990 (N_1990,In_1375,In_1051);
nand U1991 (N_1991,In_1191,In_2314);
or U1992 (N_1992,In_833,In_214);
and U1993 (N_1993,In_2373,In_2);
nor U1994 (N_1994,In_1694,In_1800);
nand U1995 (N_1995,In_1270,In_1761);
xnor U1996 (N_1996,In_1790,In_2499);
xnor U1997 (N_1997,In_1130,In_1384);
nand U1998 (N_1998,In_1495,In_2304);
nand U1999 (N_1999,In_2433,In_2273);
xor U2000 (N_2000,In_1159,In_1166);
nor U2001 (N_2001,In_1402,In_1260);
nand U2002 (N_2002,In_1799,In_1694);
or U2003 (N_2003,In_302,In_579);
or U2004 (N_2004,In_1532,In_1264);
xor U2005 (N_2005,In_1071,In_398);
or U2006 (N_2006,In_2293,In_923);
or U2007 (N_2007,In_1389,In_956);
nor U2008 (N_2008,In_1600,In_1149);
xor U2009 (N_2009,In_0,In_2040);
nor U2010 (N_2010,In_1952,In_2389);
xnor U2011 (N_2011,In_1350,In_2084);
or U2012 (N_2012,In_55,In_114);
and U2013 (N_2013,In_1080,In_2102);
or U2014 (N_2014,In_2106,In_1817);
nor U2015 (N_2015,In_1355,In_503);
or U2016 (N_2016,In_2087,In_1590);
or U2017 (N_2017,In_354,In_1964);
and U2018 (N_2018,In_1605,In_576);
and U2019 (N_2019,In_952,In_2337);
and U2020 (N_2020,In_266,In_864);
nor U2021 (N_2021,In_159,In_1663);
nor U2022 (N_2022,In_867,In_410);
nor U2023 (N_2023,In_1688,In_940);
or U2024 (N_2024,In_1966,In_2470);
nand U2025 (N_2025,In_1460,In_1764);
and U2026 (N_2026,In_1844,In_350);
or U2027 (N_2027,In_98,In_2333);
or U2028 (N_2028,In_2227,In_49);
or U2029 (N_2029,In_2370,In_2065);
or U2030 (N_2030,In_2434,In_148);
nor U2031 (N_2031,In_111,In_439);
xnor U2032 (N_2032,In_922,In_938);
xor U2033 (N_2033,In_2103,In_861);
or U2034 (N_2034,In_532,In_729);
nand U2035 (N_2035,In_1232,In_2283);
nand U2036 (N_2036,In_214,In_1031);
or U2037 (N_2037,In_692,In_2454);
and U2038 (N_2038,In_1781,In_2237);
xnor U2039 (N_2039,In_979,In_1668);
nor U2040 (N_2040,In_2055,In_2219);
and U2041 (N_2041,In_199,In_1673);
nor U2042 (N_2042,In_957,In_2029);
and U2043 (N_2043,In_1771,In_868);
or U2044 (N_2044,In_465,In_806);
or U2045 (N_2045,In_1533,In_1510);
and U2046 (N_2046,In_1652,In_1648);
or U2047 (N_2047,In_2356,In_1759);
nor U2048 (N_2048,In_1116,In_1399);
nor U2049 (N_2049,In_969,In_872);
nand U2050 (N_2050,In_667,In_1622);
xor U2051 (N_2051,In_383,In_63);
and U2052 (N_2052,In_1247,In_689);
and U2053 (N_2053,In_1477,In_2298);
or U2054 (N_2054,In_106,In_476);
nand U2055 (N_2055,In_559,In_1732);
xnor U2056 (N_2056,In_2467,In_1873);
nand U2057 (N_2057,In_2445,In_1544);
nand U2058 (N_2058,In_1653,In_556);
and U2059 (N_2059,In_332,In_344);
and U2060 (N_2060,In_1732,In_391);
or U2061 (N_2061,In_2205,In_1340);
xor U2062 (N_2062,In_753,In_120);
xnor U2063 (N_2063,In_2022,In_438);
nand U2064 (N_2064,In_664,In_2041);
nand U2065 (N_2065,In_2067,In_1317);
and U2066 (N_2066,In_1791,In_1536);
and U2067 (N_2067,In_495,In_157);
nand U2068 (N_2068,In_1274,In_2121);
nand U2069 (N_2069,In_1714,In_125);
nor U2070 (N_2070,In_1450,In_1244);
nand U2071 (N_2071,In_161,In_452);
nand U2072 (N_2072,In_78,In_1394);
and U2073 (N_2073,In_669,In_356);
nand U2074 (N_2074,In_1002,In_2150);
or U2075 (N_2075,In_1781,In_665);
and U2076 (N_2076,In_1191,In_2153);
xor U2077 (N_2077,In_859,In_348);
xor U2078 (N_2078,In_904,In_1559);
nor U2079 (N_2079,In_732,In_1179);
and U2080 (N_2080,In_534,In_1679);
nand U2081 (N_2081,In_1981,In_483);
xor U2082 (N_2082,In_192,In_740);
and U2083 (N_2083,In_2036,In_929);
and U2084 (N_2084,In_811,In_1082);
or U2085 (N_2085,In_1920,In_48);
nor U2086 (N_2086,In_1427,In_1528);
xnor U2087 (N_2087,In_1601,In_1982);
nor U2088 (N_2088,In_269,In_539);
nor U2089 (N_2089,In_490,In_867);
nand U2090 (N_2090,In_1053,In_875);
and U2091 (N_2091,In_527,In_2286);
or U2092 (N_2092,In_2404,In_1759);
nor U2093 (N_2093,In_373,In_1804);
and U2094 (N_2094,In_2312,In_2269);
or U2095 (N_2095,In_1729,In_713);
or U2096 (N_2096,In_2427,In_1484);
xor U2097 (N_2097,In_1288,In_741);
xnor U2098 (N_2098,In_404,In_797);
xnor U2099 (N_2099,In_229,In_2131);
or U2100 (N_2100,In_611,In_1259);
nand U2101 (N_2101,In_432,In_652);
nor U2102 (N_2102,In_1680,In_2057);
nor U2103 (N_2103,In_1136,In_774);
xnor U2104 (N_2104,In_1561,In_2010);
xor U2105 (N_2105,In_444,In_1006);
nand U2106 (N_2106,In_1771,In_1529);
xnor U2107 (N_2107,In_291,In_220);
and U2108 (N_2108,In_1929,In_1874);
xnor U2109 (N_2109,In_1109,In_795);
nand U2110 (N_2110,In_1342,In_1207);
nand U2111 (N_2111,In_1843,In_44);
and U2112 (N_2112,In_1318,In_2029);
nor U2113 (N_2113,In_2180,In_2485);
or U2114 (N_2114,In_2104,In_1096);
nand U2115 (N_2115,In_493,In_1616);
or U2116 (N_2116,In_2345,In_640);
xnor U2117 (N_2117,In_307,In_2002);
nor U2118 (N_2118,In_1574,In_1395);
xnor U2119 (N_2119,In_1499,In_813);
or U2120 (N_2120,In_517,In_777);
xnor U2121 (N_2121,In_1213,In_488);
or U2122 (N_2122,In_1260,In_1983);
and U2123 (N_2123,In_189,In_2053);
nand U2124 (N_2124,In_51,In_1612);
and U2125 (N_2125,In_2352,In_1344);
or U2126 (N_2126,In_513,In_680);
xnor U2127 (N_2127,In_1348,In_719);
xnor U2128 (N_2128,In_2264,In_1790);
and U2129 (N_2129,In_2421,In_1206);
nor U2130 (N_2130,In_349,In_1221);
nand U2131 (N_2131,In_1707,In_966);
nor U2132 (N_2132,In_2288,In_86);
and U2133 (N_2133,In_1960,In_488);
or U2134 (N_2134,In_954,In_839);
xor U2135 (N_2135,In_1468,In_1793);
xnor U2136 (N_2136,In_420,In_1717);
nor U2137 (N_2137,In_2403,In_1771);
xor U2138 (N_2138,In_69,In_2493);
nor U2139 (N_2139,In_534,In_455);
and U2140 (N_2140,In_1410,In_2418);
nand U2141 (N_2141,In_2444,In_396);
nand U2142 (N_2142,In_893,In_2135);
nor U2143 (N_2143,In_944,In_640);
or U2144 (N_2144,In_1405,In_79);
and U2145 (N_2145,In_469,In_659);
xnor U2146 (N_2146,In_873,In_1932);
and U2147 (N_2147,In_1532,In_2086);
and U2148 (N_2148,In_1508,In_1554);
and U2149 (N_2149,In_743,In_1268);
nand U2150 (N_2150,In_473,In_175);
or U2151 (N_2151,In_1935,In_48);
and U2152 (N_2152,In_2255,In_2344);
xnor U2153 (N_2153,In_2181,In_894);
nand U2154 (N_2154,In_1128,In_2315);
and U2155 (N_2155,In_289,In_556);
or U2156 (N_2156,In_1785,In_118);
nor U2157 (N_2157,In_1284,In_1844);
xnor U2158 (N_2158,In_2119,In_313);
nand U2159 (N_2159,In_811,In_704);
and U2160 (N_2160,In_1498,In_540);
or U2161 (N_2161,In_935,In_2460);
or U2162 (N_2162,In_1405,In_1806);
xnor U2163 (N_2163,In_1838,In_509);
nand U2164 (N_2164,In_1199,In_438);
nor U2165 (N_2165,In_742,In_1215);
xnor U2166 (N_2166,In_976,In_2341);
nand U2167 (N_2167,In_1172,In_1963);
nand U2168 (N_2168,In_1139,In_1459);
nor U2169 (N_2169,In_1890,In_724);
nor U2170 (N_2170,In_956,In_2471);
nor U2171 (N_2171,In_1433,In_588);
and U2172 (N_2172,In_288,In_572);
or U2173 (N_2173,In_1086,In_83);
nor U2174 (N_2174,In_1712,In_1841);
nand U2175 (N_2175,In_2457,In_2417);
or U2176 (N_2176,In_1329,In_1850);
xnor U2177 (N_2177,In_406,In_1101);
nor U2178 (N_2178,In_286,In_817);
nor U2179 (N_2179,In_423,In_1606);
nor U2180 (N_2180,In_678,In_2197);
and U2181 (N_2181,In_2245,In_1920);
nand U2182 (N_2182,In_423,In_1958);
and U2183 (N_2183,In_940,In_1348);
or U2184 (N_2184,In_1276,In_2274);
or U2185 (N_2185,In_741,In_2165);
nor U2186 (N_2186,In_776,In_1430);
or U2187 (N_2187,In_97,In_2486);
or U2188 (N_2188,In_2067,In_2491);
or U2189 (N_2189,In_2383,In_2415);
and U2190 (N_2190,In_334,In_939);
or U2191 (N_2191,In_1694,In_816);
and U2192 (N_2192,In_179,In_373);
nor U2193 (N_2193,In_1671,In_784);
xor U2194 (N_2194,In_886,In_1876);
nor U2195 (N_2195,In_2358,In_2131);
nor U2196 (N_2196,In_159,In_57);
or U2197 (N_2197,In_448,In_2025);
or U2198 (N_2198,In_958,In_1296);
or U2199 (N_2199,In_2278,In_1828);
nand U2200 (N_2200,In_118,In_349);
and U2201 (N_2201,In_896,In_143);
or U2202 (N_2202,In_2391,In_2443);
xor U2203 (N_2203,In_1729,In_96);
or U2204 (N_2204,In_1881,In_1970);
and U2205 (N_2205,In_1278,In_1390);
xor U2206 (N_2206,In_374,In_1557);
and U2207 (N_2207,In_254,In_2491);
nand U2208 (N_2208,In_1605,In_1882);
nand U2209 (N_2209,In_2178,In_99);
nand U2210 (N_2210,In_174,In_1969);
or U2211 (N_2211,In_303,In_1982);
nand U2212 (N_2212,In_2394,In_1017);
or U2213 (N_2213,In_2369,In_1500);
nor U2214 (N_2214,In_659,In_712);
nand U2215 (N_2215,In_1901,In_1654);
and U2216 (N_2216,In_1984,In_1420);
and U2217 (N_2217,In_1687,In_2062);
or U2218 (N_2218,In_1564,In_824);
and U2219 (N_2219,In_2392,In_2326);
nor U2220 (N_2220,In_893,In_769);
and U2221 (N_2221,In_1010,In_1471);
and U2222 (N_2222,In_1527,In_612);
or U2223 (N_2223,In_2359,In_748);
nor U2224 (N_2224,In_862,In_367);
or U2225 (N_2225,In_1116,In_1098);
xor U2226 (N_2226,In_2149,In_903);
and U2227 (N_2227,In_2161,In_693);
and U2228 (N_2228,In_685,In_1485);
xor U2229 (N_2229,In_309,In_1724);
or U2230 (N_2230,In_1633,In_2228);
xnor U2231 (N_2231,In_266,In_385);
and U2232 (N_2232,In_2415,In_587);
xor U2233 (N_2233,In_1630,In_50);
nor U2234 (N_2234,In_1684,In_2206);
nand U2235 (N_2235,In_868,In_1796);
xor U2236 (N_2236,In_1730,In_2054);
xor U2237 (N_2237,In_728,In_2402);
nor U2238 (N_2238,In_1567,In_805);
and U2239 (N_2239,In_1529,In_770);
nand U2240 (N_2240,In_2150,In_1577);
and U2241 (N_2241,In_542,In_1636);
xnor U2242 (N_2242,In_1679,In_122);
nor U2243 (N_2243,In_1218,In_1043);
and U2244 (N_2244,In_1566,In_708);
nand U2245 (N_2245,In_2085,In_1788);
nor U2246 (N_2246,In_1484,In_2382);
nand U2247 (N_2247,In_1163,In_1529);
xnor U2248 (N_2248,In_2144,In_2205);
xnor U2249 (N_2249,In_1277,In_1306);
xor U2250 (N_2250,In_1623,In_1118);
nor U2251 (N_2251,In_1539,In_1361);
or U2252 (N_2252,In_23,In_2105);
and U2253 (N_2253,In_1842,In_1942);
nand U2254 (N_2254,In_659,In_1782);
and U2255 (N_2255,In_1544,In_138);
xor U2256 (N_2256,In_1285,In_596);
and U2257 (N_2257,In_874,In_1743);
xor U2258 (N_2258,In_89,In_1427);
or U2259 (N_2259,In_589,In_2309);
xor U2260 (N_2260,In_191,In_425);
nor U2261 (N_2261,In_2459,In_1956);
and U2262 (N_2262,In_163,In_866);
and U2263 (N_2263,In_2007,In_802);
xor U2264 (N_2264,In_756,In_1536);
and U2265 (N_2265,In_1209,In_722);
or U2266 (N_2266,In_635,In_1169);
and U2267 (N_2267,In_4,In_1721);
or U2268 (N_2268,In_588,In_1244);
xor U2269 (N_2269,In_99,In_2293);
nand U2270 (N_2270,In_1738,In_1655);
nand U2271 (N_2271,In_2034,In_2047);
or U2272 (N_2272,In_1007,In_296);
nand U2273 (N_2273,In_1786,In_139);
and U2274 (N_2274,In_208,In_2389);
nand U2275 (N_2275,In_482,In_1784);
and U2276 (N_2276,In_2275,In_139);
and U2277 (N_2277,In_1752,In_691);
nand U2278 (N_2278,In_1550,In_2000);
xor U2279 (N_2279,In_1969,In_1283);
xnor U2280 (N_2280,In_1176,In_1134);
and U2281 (N_2281,In_238,In_120);
xor U2282 (N_2282,In_896,In_2221);
xor U2283 (N_2283,In_2275,In_2074);
or U2284 (N_2284,In_1054,In_984);
nor U2285 (N_2285,In_649,In_244);
nand U2286 (N_2286,In_2283,In_2163);
nand U2287 (N_2287,In_2469,In_1683);
and U2288 (N_2288,In_1059,In_767);
and U2289 (N_2289,In_1394,In_348);
and U2290 (N_2290,In_1468,In_1426);
nand U2291 (N_2291,In_52,In_2244);
xnor U2292 (N_2292,In_371,In_1849);
nor U2293 (N_2293,In_982,In_2025);
nand U2294 (N_2294,In_107,In_1718);
and U2295 (N_2295,In_2099,In_1714);
xnor U2296 (N_2296,In_817,In_656);
and U2297 (N_2297,In_1572,In_1028);
nand U2298 (N_2298,In_1553,In_2423);
nand U2299 (N_2299,In_1728,In_708);
nor U2300 (N_2300,In_2347,In_1235);
nand U2301 (N_2301,In_1666,In_1096);
or U2302 (N_2302,In_2432,In_1484);
and U2303 (N_2303,In_543,In_1099);
nor U2304 (N_2304,In_1602,In_1014);
or U2305 (N_2305,In_183,In_2101);
xnor U2306 (N_2306,In_166,In_955);
nand U2307 (N_2307,In_1359,In_104);
xnor U2308 (N_2308,In_860,In_336);
nor U2309 (N_2309,In_2031,In_1788);
or U2310 (N_2310,In_332,In_1617);
and U2311 (N_2311,In_451,In_1653);
nand U2312 (N_2312,In_1908,In_735);
nand U2313 (N_2313,In_1613,In_2106);
or U2314 (N_2314,In_615,In_1810);
and U2315 (N_2315,In_2193,In_775);
or U2316 (N_2316,In_232,In_420);
nand U2317 (N_2317,In_1826,In_837);
nor U2318 (N_2318,In_1081,In_1847);
or U2319 (N_2319,In_376,In_1098);
nand U2320 (N_2320,In_820,In_1542);
nor U2321 (N_2321,In_1147,In_34);
nor U2322 (N_2322,In_28,In_1918);
nand U2323 (N_2323,In_2457,In_513);
xor U2324 (N_2324,In_604,In_1990);
nor U2325 (N_2325,In_64,In_1881);
nand U2326 (N_2326,In_1812,In_911);
xor U2327 (N_2327,In_1971,In_2174);
xor U2328 (N_2328,In_1518,In_92);
nor U2329 (N_2329,In_40,In_1320);
or U2330 (N_2330,In_294,In_397);
xnor U2331 (N_2331,In_1710,In_2204);
or U2332 (N_2332,In_1023,In_2420);
nor U2333 (N_2333,In_545,In_2423);
xor U2334 (N_2334,In_311,In_435);
nand U2335 (N_2335,In_124,In_11);
or U2336 (N_2336,In_721,In_1557);
and U2337 (N_2337,In_617,In_734);
or U2338 (N_2338,In_1445,In_1928);
nand U2339 (N_2339,In_1993,In_1673);
nor U2340 (N_2340,In_2483,In_924);
or U2341 (N_2341,In_2222,In_2067);
nand U2342 (N_2342,In_709,In_2428);
and U2343 (N_2343,In_2032,In_145);
nand U2344 (N_2344,In_1945,In_441);
xnor U2345 (N_2345,In_1687,In_658);
nor U2346 (N_2346,In_1764,In_1581);
or U2347 (N_2347,In_597,In_874);
and U2348 (N_2348,In_2061,In_1987);
xnor U2349 (N_2349,In_328,In_1337);
and U2350 (N_2350,In_1590,In_1421);
or U2351 (N_2351,In_2091,In_245);
nand U2352 (N_2352,In_434,In_1361);
nand U2353 (N_2353,In_461,In_1986);
or U2354 (N_2354,In_1480,In_554);
and U2355 (N_2355,In_366,In_1458);
or U2356 (N_2356,In_624,In_534);
xor U2357 (N_2357,In_633,In_741);
or U2358 (N_2358,In_1054,In_2379);
nor U2359 (N_2359,In_2114,In_1697);
xnor U2360 (N_2360,In_572,In_2251);
xnor U2361 (N_2361,In_190,In_2063);
nor U2362 (N_2362,In_448,In_2463);
nand U2363 (N_2363,In_1259,In_925);
and U2364 (N_2364,In_1386,In_1485);
xnor U2365 (N_2365,In_1331,In_295);
xor U2366 (N_2366,In_1689,In_432);
nor U2367 (N_2367,In_1248,In_244);
or U2368 (N_2368,In_604,In_2382);
or U2369 (N_2369,In_944,In_513);
or U2370 (N_2370,In_1667,In_533);
and U2371 (N_2371,In_271,In_1657);
xor U2372 (N_2372,In_671,In_2341);
nand U2373 (N_2373,In_1164,In_894);
nand U2374 (N_2374,In_484,In_1087);
xor U2375 (N_2375,In_22,In_2323);
xnor U2376 (N_2376,In_1806,In_1242);
xor U2377 (N_2377,In_597,In_1632);
nand U2378 (N_2378,In_2451,In_572);
and U2379 (N_2379,In_892,In_577);
nand U2380 (N_2380,In_864,In_154);
or U2381 (N_2381,In_0,In_17);
nor U2382 (N_2382,In_1513,In_428);
or U2383 (N_2383,In_749,In_1541);
or U2384 (N_2384,In_337,In_1454);
nor U2385 (N_2385,In_255,In_1986);
xnor U2386 (N_2386,In_2037,In_789);
or U2387 (N_2387,In_2091,In_2061);
and U2388 (N_2388,In_1966,In_306);
nor U2389 (N_2389,In_452,In_850);
nand U2390 (N_2390,In_49,In_271);
xnor U2391 (N_2391,In_966,In_1492);
nand U2392 (N_2392,In_2340,In_2141);
nand U2393 (N_2393,In_707,In_2047);
nand U2394 (N_2394,In_918,In_445);
and U2395 (N_2395,In_1613,In_700);
or U2396 (N_2396,In_1952,In_2039);
xor U2397 (N_2397,In_312,In_83);
and U2398 (N_2398,In_25,In_2041);
or U2399 (N_2399,In_1636,In_387);
xor U2400 (N_2400,In_1322,In_94);
xor U2401 (N_2401,In_573,In_710);
and U2402 (N_2402,In_1347,In_2436);
nor U2403 (N_2403,In_1367,In_1720);
and U2404 (N_2404,In_1562,In_326);
nand U2405 (N_2405,In_840,In_745);
or U2406 (N_2406,In_932,In_430);
or U2407 (N_2407,In_2170,In_634);
nor U2408 (N_2408,In_558,In_674);
or U2409 (N_2409,In_1045,In_1929);
nor U2410 (N_2410,In_2073,In_917);
xor U2411 (N_2411,In_2018,In_323);
or U2412 (N_2412,In_2252,In_530);
nand U2413 (N_2413,In_1122,In_1581);
or U2414 (N_2414,In_2251,In_24);
and U2415 (N_2415,In_2000,In_528);
or U2416 (N_2416,In_1778,In_352);
nor U2417 (N_2417,In_2061,In_843);
nor U2418 (N_2418,In_221,In_114);
and U2419 (N_2419,In_874,In_1719);
xnor U2420 (N_2420,In_5,In_287);
xor U2421 (N_2421,In_2284,In_2104);
xnor U2422 (N_2422,In_1833,In_2069);
nor U2423 (N_2423,In_2466,In_1126);
or U2424 (N_2424,In_793,In_452);
and U2425 (N_2425,In_1348,In_1473);
xnor U2426 (N_2426,In_2444,In_542);
or U2427 (N_2427,In_2452,In_2422);
and U2428 (N_2428,In_2168,In_1712);
and U2429 (N_2429,In_593,In_1133);
nand U2430 (N_2430,In_1564,In_1883);
nand U2431 (N_2431,In_108,In_448);
nor U2432 (N_2432,In_933,In_276);
xnor U2433 (N_2433,In_2111,In_654);
or U2434 (N_2434,In_346,In_1374);
and U2435 (N_2435,In_1706,In_1189);
nor U2436 (N_2436,In_808,In_1078);
or U2437 (N_2437,In_884,In_1144);
nor U2438 (N_2438,In_1964,In_1113);
nor U2439 (N_2439,In_2409,In_1630);
nor U2440 (N_2440,In_1146,In_811);
and U2441 (N_2441,In_85,In_960);
nand U2442 (N_2442,In_210,In_2130);
xnor U2443 (N_2443,In_1159,In_2127);
and U2444 (N_2444,In_1926,In_322);
nor U2445 (N_2445,In_843,In_1639);
xnor U2446 (N_2446,In_1090,In_347);
and U2447 (N_2447,In_1904,In_1934);
or U2448 (N_2448,In_387,In_1555);
nor U2449 (N_2449,In_1289,In_552);
xnor U2450 (N_2450,In_2066,In_776);
or U2451 (N_2451,In_851,In_2346);
and U2452 (N_2452,In_658,In_349);
and U2453 (N_2453,In_1184,In_1396);
nand U2454 (N_2454,In_1795,In_2137);
or U2455 (N_2455,In_2453,In_1262);
and U2456 (N_2456,In_913,In_1195);
nor U2457 (N_2457,In_198,In_18);
and U2458 (N_2458,In_1797,In_2142);
or U2459 (N_2459,In_1462,In_976);
or U2460 (N_2460,In_835,In_636);
or U2461 (N_2461,In_1675,In_774);
nand U2462 (N_2462,In_197,In_350);
and U2463 (N_2463,In_1753,In_1549);
xnor U2464 (N_2464,In_1776,In_2323);
xor U2465 (N_2465,In_420,In_740);
and U2466 (N_2466,In_1237,In_1052);
or U2467 (N_2467,In_1468,In_1962);
or U2468 (N_2468,In_1856,In_1968);
nor U2469 (N_2469,In_2249,In_510);
or U2470 (N_2470,In_1068,In_1038);
nor U2471 (N_2471,In_1198,In_362);
nand U2472 (N_2472,In_88,In_591);
nand U2473 (N_2473,In_1773,In_2065);
or U2474 (N_2474,In_1882,In_1221);
and U2475 (N_2475,In_474,In_1728);
and U2476 (N_2476,In_124,In_72);
or U2477 (N_2477,In_633,In_266);
or U2478 (N_2478,In_1430,In_2105);
and U2479 (N_2479,In_218,In_141);
or U2480 (N_2480,In_1837,In_1491);
nor U2481 (N_2481,In_2148,In_1449);
nor U2482 (N_2482,In_867,In_1222);
or U2483 (N_2483,In_2034,In_1064);
or U2484 (N_2484,In_37,In_864);
nand U2485 (N_2485,In_1954,In_885);
xnor U2486 (N_2486,In_148,In_774);
or U2487 (N_2487,In_2249,In_157);
nor U2488 (N_2488,In_1238,In_203);
nand U2489 (N_2489,In_422,In_1453);
or U2490 (N_2490,In_1877,In_1867);
nand U2491 (N_2491,In_1706,In_2069);
nand U2492 (N_2492,In_2243,In_1763);
and U2493 (N_2493,In_688,In_151);
nand U2494 (N_2494,In_22,In_2068);
nand U2495 (N_2495,In_1866,In_1010);
nor U2496 (N_2496,In_1677,In_1867);
nor U2497 (N_2497,In_904,In_986);
nor U2498 (N_2498,In_2480,In_2103);
nand U2499 (N_2499,In_2380,In_410);
and U2500 (N_2500,N_1524,N_2111);
or U2501 (N_2501,N_2149,N_1772);
or U2502 (N_2502,N_112,N_1826);
and U2503 (N_2503,N_1965,N_1843);
or U2504 (N_2504,N_570,N_2235);
nor U2505 (N_2505,N_1445,N_288);
or U2506 (N_2506,N_2433,N_178);
xor U2507 (N_2507,N_680,N_1838);
or U2508 (N_2508,N_1812,N_2252);
xnor U2509 (N_2509,N_1545,N_1743);
nor U2510 (N_2510,N_99,N_2243);
nor U2511 (N_2511,N_2300,N_486);
and U2512 (N_2512,N_690,N_2266);
nand U2513 (N_2513,N_1391,N_850);
nor U2514 (N_2514,N_1976,N_326);
and U2515 (N_2515,N_1907,N_2291);
or U2516 (N_2516,N_1557,N_123);
or U2517 (N_2517,N_678,N_1181);
and U2518 (N_2518,N_615,N_1926);
nand U2519 (N_2519,N_1067,N_1021);
or U2520 (N_2520,N_66,N_724);
or U2521 (N_2521,N_1819,N_103);
nor U2522 (N_2522,N_412,N_1556);
or U2523 (N_2523,N_2466,N_164);
xnor U2524 (N_2524,N_2072,N_1140);
xor U2525 (N_2525,N_682,N_196);
xnor U2526 (N_2526,N_313,N_741);
nand U2527 (N_2527,N_1927,N_1124);
nand U2528 (N_2528,N_723,N_2430);
and U2529 (N_2529,N_28,N_432);
or U2530 (N_2530,N_710,N_247);
nand U2531 (N_2531,N_889,N_2044);
nor U2532 (N_2532,N_906,N_1918);
and U2533 (N_2533,N_1733,N_506);
or U2534 (N_2534,N_21,N_996);
xor U2535 (N_2535,N_2486,N_2454);
nand U2536 (N_2536,N_1368,N_275);
nand U2537 (N_2537,N_1191,N_1861);
nand U2538 (N_2538,N_1254,N_1810);
nand U2539 (N_2539,N_870,N_2267);
nand U2540 (N_2540,N_1063,N_1590);
or U2541 (N_2541,N_117,N_509);
or U2542 (N_2542,N_1880,N_1240);
nor U2543 (N_2543,N_1839,N_2058);
xor U2544 (N_2544,N_1046,N_344);
and U2545 (N_2545,N_1328,N_1916);
or U2546 (N_2546,N_552,N_888);
nand U2547 (N_2547,N_2355,N_556);
and U2548 (N_2548,N_1589,N_1227);
xnor U2549 (N_2549,N_974,N_2398);
nor U2550 (N_2550,N_1239,N_1538);
nand U2551 (N_2551,N_120,N_716);
nand U2552 (N_2552,N_366,N_757);
and U2553 (N_2553,N_12,N_143);
and U2554 (N_2554,N_1206,N_2117);
nor U2555 (N_2555,N_2254,N_1582);
and U2556 (N_2556,N_647,N_330);
and U2557 (N_2557,N_1888,N_1016);
and U2558 (N_2558,N_2459,N_2069);
nand U2559 (N_2559,N_1986,N_2108);
nor U2560 (N_2560,N_407,N_1592);
or U2561 (N_2561,N_2045,N_1648);
or U2562 (N_2562,N_297,N_1152);
xor U2563 (N_2563,N_1494,N_2244);
nor U2564 (N_2564,N_2023,N_141);
nand U2565 (N_2565,N_995,N_2070);
nand U2566 (N_2566,N_2217,N_638);
and U2567 (N_2567,N_1241,N_16);
and U2568 (N_2568,N_2078,N_2320);
or U2569 (N_2569,N_1564,N_2145);
and U2570 (N_2570,N_2008,N_1363);
nand U2571 (N_2571,N_1030,N_1229);
nand U2572 (N_2572,N_1755,N_769);
nand U2573 (N_2573,N_46,N_1774);
and U2574 (N_2574,N_1516,N_2406);
nor U2575 (N_2575,N_1284,N_1497);
nand U2576 (N_2576,N_1272,N_2490);
nor U2577 (N_2577,N_1491,N_1212);
or U2578 (N_2578,N_492,N_1535);
and U2579 (N_2579,N_505,N_583);
or U2580 (N_2580,N_965,N_1773);
and U2581 (N_2581,N_118,N_2193);
nand U2582 (N_2582,N_2160,N_984);
nor U2583 (N_2583,N_1040,N_242);
or U2584 (N_2584,N_1035,N_175);
xnor U2585 (N_2585,N_2002,N_327);
nor U2586 (N_2586,N_1514,N_1257);
xnor U2587 (N_2587,N_2180,N_825);
nor U2588 (N_2588,N_2060,N_1796);
and U2589 (N_2589,N_1584,N_166);
or U2590 (N_2590,N_2182,N_232);
xnor U2591 (N_2591,N_1468,N_1325);
nor U2592 (N_2592,N_1768,N_2250);
and U2593 (N_2593,N_2307,N_476);
xor U2594 (N_2594,N_2453,N_610);
or U2595 (N_2595,N_2034,N_283);
nor U2596 (N_2596,N_1473,N_2049);
nand U2597 (N_2597,N_1388,N_390);
or U2598 (N_2598,N_2068,N_999);
nand U2599 (N_2599,N_1139,N_1218);
nor U2600 (N_2600,N_1578,N_1287);
and U2601 (N_2601,N_1065,N_1381);
or U2602 (N_2602,N_1671,N_1682);
and U2603 (N_2603,N_1946,N_74);
xor U2604 (N_2604,N_567,N_2482);
xnor U2605 (N_2605,N_87,N_2370);
nand U2606 (N_2606,N_466,N_942);
nand U2607 (N_2607,N_738,N_1486);
xnor U2608 (N_2608,N_2374,N_2269);
nand U2609 (N_2609,N_2134,N_1998);
nor U2610 (N_2610,N_382,N_2241);
or U2611 (N_2611,N_11,N_1307);
or U2612 (N_2612,N_1354,N_1247);
xor U2613 (N_2613,N_1052,N_1051);
xor U2614 (N_2614,N_1594,N_2222);
and U2615 (N_2615,N_219,N_1170);
xnor U2616 (N_2616,N_662,N_271);
and U2617 (N_2617,N_1717,N_363);
or U2618 (N_2618,N_833,N_2450);
and U2619 (N_2619,N_1673,N_240);
nor U2620 (N_2620,N_93,N_1698);
xnor U2621 (N_2621,N_1709,N_705);
or U2622 (N_2622,N_1728,N_352);
and U2623 (N_2623,N_935,N_33);
and U2624 (N_2624,N_304,N_2128);
nand U2625 (N_2625,N_670,N_2124);
and U2626 (N_2626,N_537,N_594);
xor U2627 (N_2627,N_1162,N_1908);
nand U2628 (N_2628,N_138,N_1133);
nor U2629 (N_2629,N_1090,N_1281);
or U2630 (N_2630,N_1365,N_548);
nand U2631 (N_2631,N_115,N_1077);
nand U2632 (N_2632,N_477,N_1575);
or U2633 (N_2633,N_1457,N_2027);
xor U2634 (N_2634,N_1807,N_1580);
or U2635 (N_2635,N_694,N_1448);
or U2636 (N_2636,N_2474,N_1741);
xnor U2637 (N_2637,N_712,N_8);
or U2638 (N_2638,N_763,N_1781);
xnor U2639 (N_2639,N_456,N_1657);
xor U2640 (N_2640,N_1945,N_337);
nor U2641 (N_2641,N_1808,N_2437);
nand U2642 (N_2642,N_2326,N_475);
nor U2643 (N_2643,N_377,N_2122);
or U2644 (N_2644,N_245,N_2246);
or U2645 (N_2645,N_639,N_1537);
or U2646 (N_2646,N_2349,N_2133);
and U2647 (N_2647,N_1495,N_436);
or U2648 (N_2648,N_940,N_1964);
and U2649 (N_2649,N_177,N_676);
and U2650 (N_2650,N_643,N_41);
xor U2651 (N_2651,N_105,N_1788);
and U2652 (N_2652,N_1539,N_1729);
nand U2653 (N_2653,N_1528,N_986);
and U2654 (N_2654,N_438,N_2280);
xor U2655 (N_2655,N_2277,N_736);
and U2656 (N_2656,N_564,N_2009);
or U2657 (N_2657,N_1285,N_2356);
xnor U2658 (N_2658,N_1470,N_1425);
nand U2659 (N_2659,N_1342,N_2340);
xnor U2660 (N_2660,N_1695,N_1715);
nand U2661 (N_2661,N_793,N_568);
nor U2662 (N_2662,N_1586,N_701);
nor U2663 (N_2663,N_2396,N_2471);
or U2664 (N_2664,N_1782,N_392);
xor U2665 (N_2665,N_201,N_897);
and U2666 (N_2666,N_836,N_65);
and U2667 (N_2667,N_1422,N_525);
or U2668 (N_2668,N_696,N_1867);
xor U2669 (N_2669,N_2238,N_2228);
and U2670 (N_2670,N_1430,N_2175);
nor U2671 (N_2671,N_530,N_1074);
nor U2672 (N_2672,N_578,N_1231);
xor U2673 (N_2673,N_1544,N_2156);
nor U2674 (N_2674,N_1713,N_931);
or U2675 (N_2675,N_659,N_1332);
xor U2676 (N_2676,N_1453,N_318);
nor U2677 (N_2677,N_1746,N_422);
and U2678 (N_2678,N_406,N_1439);
xor U2679 (N_2679,N_1025,N_2048);
or U2680 (N_2680,N_1460,N_2328);
nand U2681 (N_2681,N_1230,N_268);
nand U2682 (N_2682,N_2348,N_130);
nand U2683 (N_2683,N_214,N_184);
and U2684 (N_2684,N_1959,N_1094);
nand U2685 (N_2685,N_1237,N_223);
nand U2686 (N_2686,N_380,N_584);
nand U2687 (N_2687,N_1656,N_565);
nand U2688 (N_2688,N_1195,N_1968);
nor U2689 (N_2689,N_1747,N_844);
and U2690 (N_2690,N_399,N_619);
nor U2691 (N_2691,N_563,N_895);
xnor U2692 (N_2692,N_1120,N_1103);
nor U2693 (N_2693,N_2299,N_2303);
and U2694 (N_2694,N_424,N_1294);
and U2695 (N_2695,N_485,N_2470);
nor U2696 (N_2696,N_234,N_1409);
or U2697 (N_2697,N_1800,N_129);
nor U2698 (N_2698,N_1655,N_1936);
or U2699 (N_2699,N_616,N_2127);
or U2700 (N_2700,N_461,N_2062);
xor U2701 (N_2701,N_2265,N_1909);
or U2702 (N_2702,N_1121,N_1625);
and U2703 (N_2703,N_1851,N_1361);
xnor U2704 (N_2704,N_902,N_733);
nand U2705 (N_2705,N_1367,N_1441);
and U2706 (N_2706,N_633,N_884);
nand U2707 (N_2707,N_1174,N_2112);
xor U2708 (N_2708,N_2331,N_310);
and U2709 (N_2709,N_1338,N_745);
nor U2710 (N_2710,N_587,N_425);
nor U2711 (N_2711,N_915,N_651);
and U2712 (N_2712,N_677,N_2196);
nand U2713 (N_2713,N_2088,N_2102);
nand U2714 (N_2714,N_1923,N_2093);
nor U2715 (N_2715,N_2408,N_554);
or U2716 (N_2716,N_954,N_2064);
nor U2717 (N_2717,N_987,N_673);
xor U2718 (N_2718,N_9,N_1270);
xnor U2719 (N_2719,N_846,N_797);
nor U2720 (N_2720,N_36,N_2080);
nor U2721 (N_2721,N_286,N_2099);
or U2722 (N_2722,N_1399,N_1670);
nand U2723 (N_2723,N_96,N_347);
and U2724 (N_2724,N_1066,N_17);
nand U2725 (N_2725,N_2157,N_484);
or U2726 (N_2726,N_167,N_2439);
nand U2727 (N_2727,N_1718,N_919);
or U2728 (N_2728,N_2010,N_1394);
and U2729 (N_2729,N_1956,N_146);
or U2730 (N_2730,N_2473,N_722);
nand U2731 (N_2731,N_2065,N_847);
xor U2732 (N_2732,N_887,N_1014);
and U2733 (N_2733,N_86,N_1476);
and U2734 (N_2734,N_2181,N_249);
xor U2735 (N_2735,N_1119,N_1898);
nand U2736 (N_2736,N_2037,N_2493);
nand U2737 (N_2737,N_497,N_1037);
nand U2738 (N_2738,N_1228,N_1147);
and U2739 (N_2739,N_1700,N_1114);
nor U2740 (N_2740,N_1279,N_32);
xor U2741 (N_2741,N_1913,N_898);
nor U2742 (N_2742,N_539,N_758);
nand U2743 (N_2743,N_1532,N_452);
nor U2744 (N_2744,N_629,N_636);
nor U2745 (N_2745,N_307,N_1244);
nor U2746 (N_2746,N_707,N_1322);
nor U2747 (N_2747,N_684,N_2480);
nand U2748 (N_2748,N_2184,N_1737);
and U2749 (N_2749,N_717,N_305);
xor U2750 (N_2750,N_373,N_2361);
and U2751 (N_2751,N_1649,N_838);
nor U2752 (N_2752,N_1263,N_504);
and U2753 (N_2753,N_1804,N_864);
nor U2754 (N_2754,N_613,N_2053);
xor U2755 (N_2755,N_1493,N_470);
xor U2756 (N_2756,N_1496,N_1846);
xor U2757 (N_2757,N_291,N_1500);
and U2758 (N_2758,N_1847,N_1615);
nand U2759 (N_2759,N_1172,N_98);
and U2760 (N_2760,N_2276,N_2239);
xor U2761 (N_2761,N_1568,N_1899);
or U2762 (N_2762,N_1689,N_883);
and U2763 (N_2763,N_1881,N_1204);
nand U2764 (N_2764,N_1901,N_2357);
nand U2765 (N_2765,N_1143,N_1672);
nor U2766 (N_2766,N_315,N_1969);
or U2767 (N_2767,N_2268,N_2342);
xnor U2768 (N_2768,N_1627,N_2046);
nor U2769 (N_2769,N_2118,N_1278);
xnor U2770 (N_2770,N_2264,N_19);
nor U2771 (N_2771,N_2395,N_2467);
nor U2772 (N_2772,N_1640,N_573);
nand U2773 (N_2773,N_1061,N_1803);
xor U2774 (N_2774,N_2358,N_671);
nand U2775 (N_2775,N_725,N_877);
xor U2776 (N_2776,N_926,N_1548);
and U2777 (N_2777,N_1925,N_341);
or U2778 (N_2778,N_2383,N_905);
or U2779 (N_2779,N_159,N_1403);
nor U2780 (N_2780,N_1132,N_56);
nor U2781 (N_2781,N_1166,N_973);
xor U2782 (N_2782,N_1101,N_2123);
nand U2783 (N_2783,N_2248,N_1815);
nand U2784 (N_2784,N_2317,N_1864);
nor U2785 (N_2785,N_1631,N_1857);
nand U2786 (N_2786,N_1771,N_1440);
nand U2787 (N_2787,N_1612,N_2188);
nor U2788 (N_2788,N_1759,N_311);
and U2789 (N_2789,N_100,N_1823);
nor U2790 (N_2790,N_241,N_365);
or U2791 (N_2791,N_1963,N_1082);
or U2792 (N_2792,N_1056,N_1680);
nor U2793 (N_2793,N_1744,N_1975);
and U2794 (N_2794,N_462,N_1326);
or U2795 (N_2795,N_398,N_478);
xor U2796 (N_2796,N_695,N_1396);
or U2797 (N_2797,N_1570,N_1947);
xnor U2798 (N_2798,N_405,N_1748);
or U2799 (N_2799,N_1375,N_2032);
nand U2800 (N_2800,N_59,N_985);
or U2801 (N_2801,N_198,N_2379);
and U2802 (N_2802,N_934,N_2139);
nand U2803 (N_2803,N_2488,N_928);
and U2804 (N_2804,N_1225,N_1297);
nand U2805 (N_2805,N_2022,N_408);
and U2806 (N_2806,N_827,N_384);
or U2807 (N_2807,N_58,N_2234);
nor U2808 (N_2808,N_1232,N_2385);
and U2809 (N_2809,N_1574,N_1252);
nand U2810 (N_2810,N_230,N_1643);
nor U2811 (N_2811,N_635,N_388);
xor U2812 (N_2812,N_1869,N_614);
nand U2813 (N_2813,N_1681,N_1859);
or U2814 (N_2814,N_821,N_322);
and U2815 (N_2815,N_1527,N_1767);
xnor U2816 (N_2816,N_2458,N_1319);
nor U2817 (N_2817,N_852,N_170);
and U2818 (N_2818,N_2067,N_2281);
nor U2819 (N_2819,N_2413,N_1702);
nand U2820 (N_2820,N_1371,N_136);
nor U2821 (N_2821,N_1763,N_1154);
nor U2822 (N_2822,N_1641,N_1666);
xor U2823 (N_2823,N_415,N_239);
nor U2824 (N_2824,N_1993,N_1555);
or U2825 (N_2825,N_1750,N_1012);
or U2826 (N_2826,N_429,N_1531);
xor U2827 (N_2827,N_263,N_618);
or U2828 (N_2828,N_225,N_2015);
nand U2829 (N_2829,N_445,N_1268);
and U2830 (N_2830,N_2227,N_561);
or U2831 (N_2831,N_1156,N_1688);
and U2832 (N_2832,N_2056,N_2272);
and U2833 (N_2833,N_3,N_1290);
xor U2834 (N_2834,N_1086,N_1024);
nor U2835 (N_2835,N_51,N_174);
xnor U2836 (N_2836,N_250,N_2052);
nand U2837 (N_2837,N_1591,N_2463);
and U2838 (N_2838,N_1770,N_2129);
or U2839 (N_2839,N_1006,N_1504);
xor U2840 (N_2840,N_2233,N_545);
or U2841 (N_2841,N_53,N_2420);
nand U2842 (N_2842,N_228,N_1050);
or U2843 (N_2843,N_2350,N_2116);
xnor U2844 (N_2844,N_2114,N_1558);
nand U2845 (N_2845,N_997,N_547);
and U2846 (N_2846,N_845,N_1349);
nor U2847 (N_2847,N_2314,N_939);
xnor U2848 (N_2848,N_2110,N_153);
or U2849 (N_2849,N_1117,N_2381);
xor U2850 (N_2850,N_243,N_2103);
and U2851 (N_2851,N_623,N_516);
nor U2852 (N_2852,N_591,N_389);
or U2853 (N_2853,N_1347,N_592);
or U2854 (N_2854,N_37,N_962);
or U2855 (N_2855,N_1343,N_1811);
nand U2856 (N_2856,N_127,N_1637);
and U2857 (N_2857,N_1484,N_1159);
and U2858 (N_2858,N_819,N_518);
xnor U2859 (N_2859,N_2332,N_994);
xor U2860 (N_2860,N_2362,N_1542);
or U2861 (N_2861,N_84,N_1890);
or U2862 (N_2862,N_1123,N_2445);
nor U2863 (N_2863,N_1663,N_1629);
or U2864 (N_2864,N_191,N_881);
nand U2865 (N_2865,N_218,N_444);
or U2866 (N_2866,N_1685,N_460);
or U2867 (N_2867,N_875,N_1250);
or U2868 (N_2868,N_148,N_593);
xor U2869 (N_2869,N_292,N_1920);
or U2870 (N_2870,N_2018,N_119);
nand U2871 (N_2871,N_822,N_502);
or U2872 (N_2872,N_2092,N_273);
xnor U2873 (N_2873,N_1930,N_576);
xor U2874 (N_2874,N_443,N_1203);
nand U2875 (N_2875,N_1258,N_899);
or U2876 (N_2876,N_1220,N_1188);
xor U2877 (N_2877,N_531,N_395);
nand U2878 (N_2878,N_703,N_179);
and U2879 (N_2879,N_1150,N_1169);
nor U2880 (N_2880,N_1197,N_1828);
or U2881 (N_2881,N_2327,N_15);
nor U2882 (N_2882,N_688,N_1892);
nand U2883 (N_2883,N_1415,N_1337);
or U2884 (N_2884,N_2446,N_1275);
xor U2885 (N_2885,N_1416,N_1340);
and U2886 (N_2886,N_2079,N_2345);
and U2887 (N_2887,N_2016,N_1805);
nand U2888 (N_2888,N_2012,N_2055);
and U2889 (N_2889,N_1632,N_471);
or U2890 (N_2890,N_2429,N_2190);
or U2891 (N_2891,N_744,N_258);
and U2892 (N_2892,N_781,N_417);
xor U2893 (N_2893,N_1224,N_1573);
or U2894 (N_2894,N_1001,N_2298);
xnor U2895 (N_2895,N_1190,N_10);
nor U2896 (N_2896,N_227,N_2013);
nor U2897 (N_2897,N_1299,N_1730);
nand U2898 (N_2898,N_2295,N_588);
xnor U2899 (N_2899,N_732,N_2146);
or U2900 (N_2900,N_801,N_1818);
nor U2901 (N_2901,N_910,N_640);
and U2902 (N_2902,N_2230,N_511);
and U2903 (N_2903,N_437,N_886);
or U2904 (N_2904,N_2212,N_2422);
nand U2905 (N_2905,N_1072,N_1163);
xnor U2906 (N_2906,N_1185,N_287);
nand U2907 (N_2907,N_2364,N_2036);
nand U2908 (N_2908,N_302,N_2485);
or U2909 (N_2909,N_869,N_281);
nand U2910 (N_2910,N_473,N_69);
nand U2911 (N_2911,N_1210,N_829);
nor U2912 (N_2912,N_6,N_1525);
and U2913 (N_2913,N_1981,N_1974);
nor U2914 (N_2914,N_1519,N_1834);
and U2915 (N_2915,N_930,N_2384);
xnor U2916 (N_2916,N_2094,N_1906);
xor U2917 (N_2917,N_1844,N_2158);
or U2918 (N_2918,N_1865,N_121);
and U2919 (N_2919,N_1179,N_2435);
and U2920 (N_2920,N_1585,N_26);
nor U2921 (N_2921,N_1370,N_948);
nor U2922 (N_2922,N_598,N_1602);
nor U2923 (N_2923,N_727,N_1412);
nor U2924 (N_2924,N_807,N_1112);
and U2925 (N_2925,N_1235,N_1321);
and U2926 (N_2926,N_40,N_487);
nand U2927 (N_2927,N_205,N_1509);
or U2928 (N_2928,N_2311,N_2325);
nand U2929 (N_2929,N_1824,N_371);
xor U2930 (N_2930,N_1293,N_2426);
nand U2931 (N_2931,N_152,N_111);
and U2932 (N_2932,N_1928,N_1518);
nand U2933 (N_2933,N_186,N_719);
nor U2934 (N_2934,N_1593,N_1553);
or U2935 (N_2935,N_697,N_1431);
nand U2936 (N_2936,N_189,N_50);
xor U2937 (N_2937,N_1383,N_336);
nor U2938 (N_2938,N_116,N_1026);
xor U2939 (N_2939,N_2313,N_328);
or U2940 (N_2940,N_426,N_1462);
nor U2941 (N_2941,N_2411,N_1825);
nor U2942 (N_2942,N_1380,N_2469);
and U2943 (N_2943,N_581,N_685);
nand U2944 (N_2944,N_1919,N_1511);
nand U2945 (N_2945,N_1633,N_747);
and U2946 (N_2946,N_2087,N_960);
or U2947 (N_2947,N_1078,N_495);
xnor U2948 (N_2948,N_1048,N_2168);
xor U2949 (N_2949,N_2042,N_2143);
nand U2950 (N_2950,N_872,N_1621);
nand U2951 (N_2951,N_1506,N_1871);
nand U2952 (N_2952,N_1855,N_1192);
nand U2953 (N_2953,N_970,N_1683);
xor U2954 (N_2954,N_519,N_767);
or U2955 (N_2955,N_967,N_2095);
nor U2956 (N_2956,N_278,N_862);
nor U2957 (N_2957,N_1038,N_464);
or U2958 (N_2958,N_1093,N_2166);
xnor U2959 (N_2959,N_2059,N_1098);
or U2960 (N_2960,N_180,N_368);
and U2961 (N_2961,N_2165,N_1362);
nand U2962 (N_2962,N_173,N_2199);
or U2963 (N_2963,N_2479,N_946);
nor U2964 (N_2964,N_734,N_491);
or U2965 (N_2965,N_806,N_2121);
nor U2966 (N_2966,N_1414,N_2141);
xnor U2967 (N_2967,N_1317,N_1885);
nor U2968 (N_2968,N_1488,N_1949);
nand U2969 (N_2969,N_2497,N_323);
nand U2970 (N_2970,N_270,N_1189);
or U2971 (N_2971,N_27,N_1148);
nand U2972 (N_2972,N_779,N_2419);
or U2973 (N_2973,N_773,N_1779);
and U2974 (N_2974,N_2278,N_2185);
or U2975 (N_2975,N_1161,N_267);
xor U2976 (N_2976,N_500,N_1485);
or U2977 (N_2977,N_770,N_1233);
nand U2978 (N_2978,N_420,N_1635);
nor U2979 (N_2979,N_1723,N_1018);
nor U2980 (N_2980,N_1786,N_1852);
or U2981 (N_2981,N_663,N_961);
nor U2982 (N_2982,N_2378,N_1401);
nor U2983 (N_2983,N_522,N_809);
xnor U2984 (N_2984,N_1499,N_1820);
xnor U2985 (N_2985,N_162,N_45);
nand U2986 (N_2986,N_2247,N_924);
and U2987 (N_2987,N_252,N_1245);
nand U2988 (N_2988,N_834,N_2271);
or U2989 (N_2989,N_1526,N_360);
nand U2990 (N_2990,N_2063,N_401);
or U2991 (N_2991,N_1647,N_2319);
and U2992 (N_2992,N_1449,N_1075);
and U2993 (N_2993,N_2054,N_549);
nand U2994 (N_2994,N_2414,N_0);
xnor U2995 (N_2995,N_1816,N_2465);
and U2996 (N_2996,N_2179,N_1994);
or U2997 (N_2997,N_2025,N_1171);
nand U2998 (N_2998,N_597,N_370);
nand U2999 (N_2999,N_2315,N_2390);
xnor U3000 (N_3000,N_1684,N_2392);
nand U3001 (N_3001,N_1896,N_80);
xor U3002 (N_3002,N_1937,N_381);
and U3003 (N_3003,N_2351,N_1251);
and U3004 (N_3004,N_1405,N_2041);
nor U3005 (N_3005,N_1155,N_1438);
nand U3006 (N_3006,N_1756,N_1022);
and U3007 (N_3007,N_1598,N_1356);
xnor U3008 (N_3008,N_193,N_300);
and U3009 (N_3009,N_728,N_558);
nand U3010 (N_3010,N_2462,N_1153);
nand U3011 (N_3011,N_1389,N_2005);
xor U3012 (N_3012,N_2119,N_2260);
nor U3013 (N_3013,N_718,N_1721);
xnor U3014 (N_3014,N_208,N_1291);
xor U3015 (N_3015,N_866,N_353);
and U3016 (N_3016,N_188,N_1958);
nor U3017 (N_3017,N_666,N_1764);
xnor U3018 (N_3018,N_2073,N_1752);
nor U3019 (N_3019,N_1402,N_885);
or U3020 (N_3020,N_1850,N_1692);
xnor U3021 (N_3021,N_199,N_49);
and U3022 (N_3022,N_559,N_1201);
nand U3023 (N_3023,N_1423,N_1390);
nand U3024 (N_3024,N_192,N_543);
nor U3025 (N_3025,N_1623,N_1384);
or U3026 (N_3026,N_1109,N_2347);
xor U3027 (N_3027,N_1464,N_1809);
nand U3028 (N_3028,N_169,N_465);
xnor U3029 (N_3029,N_1053,N_1127);
nor U3030 (N_3030,N_858,N_463);
nor U3031 (N_3031,N_1679,N_603);
nor U3032 (N_3032,N_2296,N_2039);
nor U3033 (N_3033,N_1406,N_35);
nor U3034 (N_3034,N_409,N_2232);
and U3035 (N_3035,N_799,N_78);
or U3036 (N_3036,N_1795,N_938);
xor U3037 (N_3037,N_1044,N_2262);
xor U3038 (N_3038,N_1853,N_1020);
or U3039 (N_3039,N_362,N_1034);
nand U3040 (N_3040,N_413,N_1407);
xnor U3041 (N_3041,N_1434,N_1207);
nor U3042 (N_3042,N_1492,N_1364);
or U3043 (N_3043,N_364,N_1707);
and U3044 (N_3044,N_731,N_715);
nand U3045 (N_3045,N_1706,N_237);
or U3046 (N_3046,N_1142,N_990);
nand U3047 (N_3047,N_79,N_171);
nor U3048 (N_3048,N_29,N_1638);
nor U3049 (N_3049,N_1213,N_1953);
nor U3050 (N_3050,N_1595,N_194);
or U3051 (N_3051,N_2033,N_1107);
xor U3052 (N_3052,N_1960,N_873);
nor U3053 (N_3053,N_144,N_1696);
nand U3054 (N_3054,N_2293,N_324);
and U3055 (N_3055,N_923,N_1259);
and U3056 (N_3056,N_1830,N_952);
nor U3057 (N_3057,N_1734,N_2401);
or U3058 (N_3058,N_1099,N_290);
and U3059 (N_3059,N_1104,N_295);
and U3060 (N_3060,N_1650,N_2394);
nand U3061 (N_3061,N_1134,N_83);
nor U3062 (N_3062,N_1199,N_1942);
nand U3063 (N_3063,N_501,N_828);
nor U3064 (N_3064,N_2498,N_2148);
xor U3065 (N_3065,N_532,N_953);
or U3066 (N_3066,N_2404,N_1551);
and U3067 (N_3067,N_868,N_963);
and U3068 (N_3068,N_713,N_1693);
nor U3069 (N_3069,N_251,N_361);
and U3070 (N_3070,N_1205,N_514);
or U3071 (N_3071,N_1561,N_2416);
nor U3072 (N_3072,N_451,N_2290);
nor U3073 (N_3073,N_1599,N_1606);
nor U3074 (N_3074,N_1286,N_776);
or U3075 (N_3075,N_1587,N_383);
xnor U3076 (N_3076,N_742,N_699);
nand U3077 (N_3077,N_2224,N_1984);
or U3078 (N_3078,N_2031,N_2057);
nor U3079 (N_3079,N_544,N_865);
xor U3080 (N_3080,N_1262,N_669);
nor U3081 (N_3081,N_319,N_977);
xor U3082 (N_3082,N_1863,N_102);
xnor U3083 (N_3083,N_1995,N_726);
xnor U3084 (N_3084,N_608,N_71);
nand U3085 (N_3085,N_2284,N_1105);
nand U3086 (N_3086,N_1611,N_1450);
or U3087 (N_3087,N_1879,N_2417);
nor U3088 (N_3088,N_400,N_1057);
nor U3089 (N_3089,N_1889,N_1616);
and U3090 (N_3090,N_766,N_1860);
nor U3091 (N_3091,N_2407,N_1661);
nand U3092 (N_3092,N_1541,N_929);
xor U3093 (N_3093,N_761,N_1353);
xnor U3094 (N_3094,N_958,N_1003);
nor U3095 (N_3095,N_2135,N_2275);
nor U3096 (N_3096,N_2255,N_2090);
and U3097 (N_3097,N_282,N_2209);
and U3098 (N_3098,N_1111,N_520);
nor U3099 (N_3099,N_908,N_2442);
nor U3100 (N_3100,N_2363,N_982);
or U3101 (N_3101,N_916,N_950);
nor U3102 (N_3102,N_2100,N_434);
or U3103 (N_3103,N_1128,N_2189);
or U3104 (N_3104,N_308,N_386);
or U3105 (N_3105,N_2304,N_2322);
nor U3106 (N_3106,N_569,N_1331);
nand U3107 (N_3107,N_1221,N_1130);
or U3108 (N_3108,N_2494,N_2402);
or U3109 (N_3109,N_1791,N_2);
and U3110 (N_3110,N_24,N_346);
xor U3111 (N_3111,N_1938,N_1358);
nor U3112 (N_3112,N_279,N_756);
or U3113 (N_3113,N_1515,N_612);
or U3114 (N_3114,N_1979,N_269);
nand U3115 (N_3115,N_1842,N_1991);
nand U3116 (N_3116,N_1822,N_2173);
or U3117 (N_3117,N_342,N_34);
xor U3118 (N_3118,N_992,N_2483);
or U3119 (N_3119,N_2201,N_190);
or U3120 (N_3120,N_527,N_1437);
and U3121 (N_3121,N_771,N_837);
xor U3122 (N_3122,N_312,N_376);
or U3123 (N_3123,N_1392,N_221);
nand U3124 (N_3124,N_1665,N_2472);
or U3125 (N_3125,N_2302,N_972);
xnor U3126 (N_3126,N_320,N_2169);
and U3127 (N_3127,N_2155,N_2152);
nand U3128 (N_3128,N_1565,N_914);
xor U3129 (N_3129,N_2258,N_762);
xor U3130 (N_3130,N_2153,N_772);
xnor U3131 (N_3131,N_602,N_1543);
nor U3132 (N_3132,N_702,N_1265);
nor U3133 (N_3133,N_2024,N_1794);
or U3134 (N_3134,N_2171,N_978);
or U3135 (N_3135,N_1714,N_1690);
or U3136 (N_3136,N_652,N_1735);
and U3137 (N_3137,N_1778,N_912);
xor U3138 (N_3138,N_1878,N_1675);
and U3139 (N_3139,N_945,N_1653);
nand U3140 (N_3140,N_1883,N_2273);
xnor U3141 (N_3141,N_654,N_2231);
nor U3142 (N_3142,N_555,N_1626);
xor U3143 (N_3143,N_743,N_2226);
nand U3144 (N_3144,N_1084,N_1990);
and U3145 (N_3145,N_835,N_1187);
or U3146 (N_3146,N_1442,N_1292);
xor U3147 (N_3147,N_1145,N_1039);
nor U3148 (N_3148,N_1324,N_468);
nor U3149 (N_3149,N_2225,N_1775);
xor U3150 (N_3150,N_2206,N_1100);
xnor U3151 (N_3151,N_1298,N_430);
or U3152 (N_3152,N_325,N_1978);
xor U3153 (N_3153,N_4,N_158);
or U3154 (N_3154,N_1397,N_687);
xnor U3155 (N_3155,N_1761,N_1295);
xor U3156 (N_3156,N_1549,N_753);
or U3157 (N_3157,N_2263,N_458);
nand U3158 (N_3158,N_752,N_2329);
nand U3159 (N_3159,N_2221,N_2257);
and U3160 (N_3160,N_675,N_1939);
xor U3161 (N_3161,N_256,N_1002);
xnor U3162 (N_3162,N_1313,N_1821);
nor U3163 (N_3163,N_2026,N_440);
nor U3164 (N_3164,N_1530,N_2105);
xor U3165 (N_3165,N_686,N_1428);
and U3166 (N_3166,N_795,N_2334);
or U3167 (N_3167,N_2489,N_2339);
or U3168 (N_3168,N_944,N_244);
nor U3169 (N_3169,N_1760,N_991);
or U3170 (N_3170,N_2415,N_1005);
nand U3171 (N_3171,N_861,N_257);
nand U3172 (N_3172,N_1421,N_2220);
or U3173 (N_3173,N_843,N_1944);
or U3174 (N_3174,N_983,N_1379);
xnor U3175 (N_3175,N_200,N_1601);
nand U3176 (N_3176,N_2424,N_260);
and U3177 (N_3177,N_1917,N_2274);
nand U3178 (N_3178,N_108,N_577);
xor U3179 (N_3179,N_951,N_1766);
xnor U3180 (N_3180,N_1957,N_1588);
nor U3181 (N_3181,N_1467,N_1977);
xnor U3182 (N_3182,N_604,N_1636);
xor U3183 (N_3183,N_794,N_2287);
xor U3184 (N_3184,N_1572,N_441);
and U3185 (N_3185,N_674,N_1691);
nor U3186 (N_3186,N_2030,N_1668);
nor U3187 (N_3187,N_1424,N_882);
or U3188 (N_3188,N_541,N_1674);
xnor U3189 (N_3189,N_515,N_1862);
nor U3190 (N_3190,N_1856,N_1008);
nand U3191 (N_3191,N_1455,N_1508);
xnor U3192 (N_3192,N_2359,N_708);
and U3193 (N_3193,N_1886,N_841);
and U3194 (N_3194,N_131,N_1320);
nor U3195 (N_3195,N_655,N_1070);
and U3196 (N_3196,N_1533,N_1654);
nand U3197 (N_3197,N_871,N_755);
xor U3198 (N_3198,N_630,N_735);
or U3199 (N_3199,N_1316,N_2183);
xor U3200 (N_3200,N_1724,N_601);
or U3201 (N_3201,N_1973,N_1922);
xor U3202 (N_3202,N_660,N_1083);
nand U3203 (N_3203,N_2371,N_798);
nor U3204 (N_3204,N_2400,N_433);
or U3205 (N_3205,N_1465,N_2464);
and U3206 (N_3206,N_2343,N_1610);
and U3207 (N_3207,N_1427,N_2035);
and U3208 (N_3208,N_749,N_480);
or U3209 (N_3209,N_1983,N_932);
xor U3210 (N_3210,N_2447,N_1534);
and U3211 (N_3211,N_2147,N_1149);
or U3212 (N_3212,N_1502,N_2191);
nor U3213 (N_3213,N_272,N_317);
nor U3214 (N_3214,N_1837,N_823);
nand U3215 (N_3215,N_2353,N_1498);
or U3216 (N_3216,N_783,N_1608);
nand U3217 (N_3217,N_306,N_340);
or U3218 (N_3218,N_1315,N_482);
or U3219 (N_3219,N_1047,N_611);
xnor U3220 (N_3220,N_1644,N_1255);
or U3221 (N_3221,N_2423,N_1567);
or U3222 (N_3222,N_1996,N_1129);
nor U3223 (N_3223,N_354,N_217);
nand U3224 (N_3224,N_1605,N_1209);
and U3225 (N_3225,N_309,N_2187);
nand U3226 (N_3226,N_2305,N_374);
xnor U3227 (N_3227,N_202,N_1160);
or U3228 (N_3228,N_472,N_2312);
nor U3229 (N_3229,N_832,N_1178);
or U3230 (N_3230,N_1784,N_1954);
nand U3231 (N_3231,N_796,N_5);
nor U3232 (N_3232,N_447,N_901);
or U3233 (N_3233,N_571,N_816);
nor U3234 (N_3234,N_2249,N_1113);
xor U3235 (N_3235,N_2130,N_1569);
xor U3236 (N_3236,N_879,N_419);
nor U3237 (N_3237,N_2289,N_145);
and U3238 (N_3238,N_54,N_212);
xnor U3239 (N_3239,N_560,N_107);
or U3240 (N_3240,N_595,N_1952);
or U3241 (N_3241,N_1443,N_2210);
nor U3242 (N_3242,N_775,N_729);
nand U3243 (N_3243,N_842,N_298);
or U3244 (N_3244,N_2294,N_2499);
and U3245 (N_3245,N_947,N_557);
xnor U3246 (N_3246,N_2297,N_2306);
nor U3247 (N_3247,N_1481,N_1081);
nor U3248 (N_3248,N_329,N_1962);
or U3249 (N_3249,N_891,N_1176);
or U3250 (N_3250,N_439,N_1208);
nor U3251 (N_3251,N_457,N_1992);
xor U3252 (N_3252,N_1507,N_813);
or U3253 (N_3253,N_774,N_55);
nand U3254 (N_3254,N_1614,N_782);
and U3255 (N_3255,N_880,N_1242);
nand U3256 (N_3256,N_2000,N_421);
nor U3257 (N_3257,N_82,N_1489);
nor U3258 (N_3258,N_2387,N_14);
xnor U3259 (N_3259,N_1302,N_1471);
or U3260 (N_3260,N_627,N_855);
and U3261 (N_3261,N_110,N_1248);
nand U3262 (N_3262,N_280,N_1041);
or U3263 (N_3263,N_276,N_264);
nor U3264 (N_3264,N_1597,N_2215);
or U3265 (N_3265,N_1335,N_1200);
xnor U3266 (N_3266,N_2492,N_1667);
or U3267 (N_3267,N_172,N_2170);
nand U3268 (N_3268,N_2242,N_2288);
xor U3269 (N_3269,N_2077,N_149);
or U3270 (N_3270,N_1799,N_1088);
or U3271 (N_3271,N_168,N_1069);
and U3272 (N_3272,N_851,N_778);
nand U3273 (N_3273,N_2097,N_754);
nor U3274 (N_3274,N_2021,N_921);
nand U3275 (N_3275,N_155,N_1745);
xnor U3276 (N_3276,N_759,N_2321);
or U3277 (N_3277,N_1135,N_1711);
nand U3278 (N_3278,N_2457,N_572);
nor U3279 (N_3279,N_1031,N_1469);
nand U3280 (N_3280,N_2195,N_2085);
xnor U3281 (N_3281,N_2083,N_2397);
and U3282 (N_3282,N_1118,N_1987);
nor U3283 (N_3283,N_1753,N_213);
nor U3284 (N_3284,N_989,N_621);
and U3285 (N_3285,N_246,N_316);
and U3286 (N_3286,N_1742,N_489);
nor U3287 (N_3287,N_72,N_1454);
xnor U3288 (N_3288,N_2427,N_2240);
xnor U3289 (N_3289,N_1897,N_1418);
or U3290 (N_3290,N_1490,N_379);
nand U3291 (N_3291,N_1277,N_450);
nand U3292 (N_3292,N_2393,N_77);
and U3293 (N_3293,N_1419,N_1646);
xor U3294 (N_3294,N_1921,N_30);
or U3295 (N_3295,N_540,N_1552);
or U3296 (N_3296,N_574,N_1997);
nand U3297 (N_3297,N_459,N_1273);
nor U3298 (N_3298,N_706,N_1659);
nor U3299 (N_3299,N_181,N_787);
xor U3300 (N_3300,N_1136,N_709);
xnor U3301 (N_3301,N_1563,N_176);
and U3302 (N_3302,N_299,N_2203);
and U3303 (N_3303,N_2151,N_1776);
and U3304 (N_3304,N_785,N_2438);
nor U3305 (N_3305,N_2354,N_197);
nand U3306 (N_3306,N_2029,N_1662);
and U3307 (N_3307,N_1131,N_453);
xor U3308 (N_3308,N_1676,N_750);
nor U3309 (N_3309,N_1004,N_1341);
nor U3310 (N_3310,N_435,N_1802);
and U3311 (N_3311,N_261,N_1011);
nor U3312 (N_3312,N_526,N_1651);
xnor U3313 (N_3313,N_1583,N_2405);
nand U3314 (N_3314,N_1400,N_209);
xor U3315 (N_3315,N_2449,N_510);
or U3316 (N_3316,N_1613,N_2071);
or U3317 (N_3317,N_2098,N_67);
and U3318 (N_3318,N_679,N_248);
xnor U3319 (N_3319,N_760,N_966);
or U3320 (N_3320,N_1260,N_345);
or U3321 (N_3321,N_937,N_971);
and U3322 (N_3322,N_1604,N_1226);
nor U3323 (N_3323,N_2318,N_1560);
xor U3324 (N_3324,N_1905,N_2285);
xor U3325 (N_3325,N_1451,N_2219);
nor U3326 (N_3326,N_1716,N_1404);
or U3327 (N_3327,N_2120,N_128);
xor U3328 (N_3328,N_1060,N_815);
xor U3329 (N_3329,N_1410,N_1330);
nand U3330 (N_3330,N_1658,N_215);
or U3331 (N_3331,N_1829,N_493);
nand U3332 (N_3332,N_2051,N_52);
nor U3333 (N_3333,N_1282,N_2202);
nor U3334 (N_3334,N_748,N_1783);
nor U3335 (N_3335,N_1789,N_2376);
nor U3336 (N_3336,N_1849,N_1032);
nor U3337 (N_3337,N_1780,N_1452);
xor U3338 (N_3338,N_13,N_968);
nand U3339 (N_3339,N_1466,N_1581);
nand U3340 (N_3340,N_1348,N_631);
nand U3341 (N_3341,N_2101,N_1607);
nand U3342 (N_3342,N_2375,N_114);
nor U3343 (N_3343,N_1787,N_393);
nand U3344 (N_3344,N_135,N_414);
xor U3345 (N_3345,N_2279,N_369);
nor U3346 (N_3346,N_988,N_1678);
or U3347 (N_3347,N_101,N_2308);
and U3348 (N_3348,N_1725,N_1068);
xor U3349 (N_3349,N_1894,N_2440);
or U3350 (N_3350,N_562,N_448);
and U3351 (N_3351,N_2132,N_1196);
and U3352 (N_3352,N_2138,N_2372);
or U3353 (N_3353,N_824,N_1249);
or U3354 (N_3354,N_1475,N_1645);
and U3355 (N_3355,N_1740,N_403);
nor U3356 (N_3356,N_2495,N_226);
or U3357 (N_3357,N_1619,N_449);
nand U3358 (N_3358,N_1660,N_2337);
xnor U3359 (N_3359,N_698,N_1872);
nand U3360 (N_3360,N_1941,N_1017);
or U3361 (N_3361,N_498,N_1216);
and U3362 (N_3362,N_416,N_1064);
nor U3363 (N_3363,N_1043,N_957);
or U3364 (N_3364,N_1948,N_216);
nand U3365 (N_3365,N_333,N_1902);
xor U3366 (N_3366,N_1314,N_1413);
and U3367 (N_3367,N_648,N_1369);
nand U3368 (N_3368,N_641,N_2316);
or U3369 (N_3369,N_1719,N_2066);
and U3370 (N_3370,N_1483,N_1444);
nor U3371 (N_3371,N_1697,N_786);
or U3372 (N_3372,N_2403,N_812);
or U3373 (N_3373,N_126,N_1429);
or U3374 (N_3374,N_1304,N_1769);
and U3375 (N_3375,N_1327,N_1887);
nor U3376 (N_3376,N_1310,N_2074);
nor U3377 (N_3377,N_1344,N_1288);
nand U3378 (N_3378,N_1141,N_182);
or U3379 (N_3379,N_1940,N_1505);
nor U3380 (N_3380,N_637,N_206);
or U3381 (N_3381,N_1432,N_1520);
and U3382 (N_3382,N_1566,N_969);
and U3383 (N_3383,N_789,N_1966);
nand U3384 (N_3384,N_1079,N_1877);
and U3385 (N_3385,N_2144,N_2164);
nand U3386 (N_3386,N_1296,N_876);
and U3387 (N_3387,N_2292,N_2451);
xnor U3388 (N_3388,N_508,N_137);
nor U3389 (N_3389,N_1267,N_358);
nor U3390 (N_3390,N_1398,N_2418);
nand U3391 (N_3391,N_1732,N_913);
xnor U3392 (N_3392,N_62,N_1751);
nand U3393 (N_3393,N_575,N_1708);
nor U3394 (N_3394,N_2399,N_1393);
nor U3395 (N_3395,N_2004,N_1562);
xor U3396 (N_3396,N_863,N_1845);
nand U3397 (N_3397,N_1126,N_1985);
or U3398 (N_3398,N_2207,N_1028);
and U3399 (N_3399,N_1929,N_1146);
or U3400 (N_3400,N_1873,N_1798);
or U3401 (N_3401,N_1091,N_1436);
nand U3402 (N_3402,N_1831,N_1870);
nand U3403 (N_3403,N_109,N_2091);
and U3404 (N_3404,N_1970,N_1318);
and U3405 (N_3405,N_20,N_1875);
and U3406 (N_3406,N_1547,N_1914);
or U3407 (N_3407,N_1276,N_1482);
nor U3408 (N_3408,N_154,N_1087);
nor U3409 (N_3409,N_512,N_488);
or U3410 (N_3410,N_1694,N_551);
xor U3411 (N_3411,N_1080,N_2301);
nor U3412 (N_3412,N_1961,N_2330);
and U3413 (N_3413,N_1013,N_2476);
and U3414 (N_3414,N_1382,N_1463);
nor U3415 (N_3415,N_2109,N_2003);
or U3416 (N_3416,N_44,N_1536);
and U3417 (N_3417,N_467,N_255);
nand U3418 (N_3418,N_91,N_1116);
nor U3419 (N_3419,N_1073,N_1350);
nor U3420 (N_3420,N_1736,N_1882);
nand U3421 (N_3421,N_48,N_2081);
xnor U3422 (N_3422,N_331,N_1333);
nand U3423 (N_3423,N_1895,N_2061);
or U3424 (N_3424,N_1447,N_1357);
xnor U3425 (N_3425,N_1151,N_2107);
xor U3426 (N_3426,N_975,N_2137);
and U3427 (N_3427,N_18,N_2338);
nor U3428 (N_3428,N_1891,N_1007);
xor U3429 (N_3429,N_427,N_2194);
nor U3430 (N_3430,N_1687,N_1703);
xor U3431 (N_3431,N_1814,N_2253);
and U3432 (N_3432,N_220,N_1943);
nor U3433 (N_3433,N_253,N_1334);
nor U3434 (N_3434,N_2475,N_2075);
nor U3435 (N_3435,N_1395,N_88);
nor U3436 (N_3436,N_2017,N_536);
nor U3437 (N_3437,N_689,N_1376);
xnor U3438 (N_3438,N_1426,N_2452);
nand U3439 (N_3439,N_1967,N_1924);
xnor U3440 (N_3440,N_2432,N_1355);
or U3441 (N_3441,N_553,N_1989);
nor U3442 (N_3442,N_410,N_2161);
or U3443 (N_3443,N_849,N_357);
and U3444 (N_3444,N_397,N_2163);
nor U3445 (N_3445,N_2218,N_1183);
xnor U3446 (N_3446,N_372,N_2270);
nor U3447 (N_3447,N_1512,N_1110);
or U3448 (N_3448,N_1329,N_1289);
nand U3449 (N_3449,N_764,N_293);
nand U3450 (N_3450,N_134,N_1704);
nor U3451 (N_3451,N_802,N_617);
nand U3452 (N_3452,N_294,N_1236);
and U3453 (N_3453,N_550,N_1762);
nor U3454 (N_3454,N_156,N_586);
nand U3455 (N_3455,N_1059,N_2441);
xor U3456 (N_3456,N_1433,N_2391);
or U3457 (N_3457,N_856,N_976);
xor U3458 (N_3458,N_254,N_1701);
and U3459 (N_3459,N_1630,N_1000);
and U3460 (N_3460,N_1712,N_1352);
xor U3461 (N_3461,N_920,N_418);
nor U3462 (N_3462,N_622,N_579);
and U3463 (N_3463,N_692,N_1387);
nand U3464 (N_3464,N_157,N_231);
or U3465 (N_3465,N_956,N_2412);
nand U3466 (N_3466,N_1577,N_70);
nor U3467 (N_3467,N_43,N_1836);
xor U3468 (N_3468,N_1617,N_1522);
nor U3469 (N_3469,N_2096,N_1754);
and U3470 (N_3470,N_1603,N_1144);
xor U3471 (N_3471,N_1710,N_1219);
or U3472 (N_3472,N_2468,N_1559);
xnor U3473 (N_3473,N_1177,N_535);
xor U3474 (N_3474,N_1833,N_2076);
and U3475 (N_3475,N_704,N_455);
nor U3476 (N_3476,N_2443,N_38);
xnor U3477 (N_3477,N_442,N_2436);
or U3478 (N_3478,N_289,N_2204);
xnor U3479 (N_3479,N_2192,N_1186);
nor U3480 (N_3480,N_1835,N_224);
nor U3481 (N_3481,N_314,N_494);
xor U3482 (N_3482,N_1312,N_1274);
or U3483 (N_3483,N_1554,N_2197);
nand U3484 (N_3484,N_503,N_1622);
nand U3485 (N_3485,N_1726,N_61);
nor U3486 (N_3486,N_1214,N_2352);
xnor U3487 (N_3487,N_1408,N_507);
and U3488 (N_3488,N_2237,N_1624);
and U3489 (N_3489,N_646,N_596);
xor U3490 (N_3490,N_1071,N_1045);
and U3491 (N_3491,N_546,N_959);
nor U3492 (N_3492,N_1019,N_645);
or U3493 (N_3493,N_42,N_1487);
xnor U3494 (N_3494,N_490,N_1385);
and U3495 (N_3495,N_751,N_1175);
xor U3496 (N_3496,N_332,N_2028);
xnor U3497 (N_3497,N_1982,N_187);
nand U3498 (N_3498,N_185,N_1374);
xor U3499 (N_3499,N_2082,N_1167);
and U3500 (N_3500,N_2336,N_1373);
nand U3501 (N_3501,N_2256,N_301);
nor U3502 (N_3502,N_229,N_351);
or U3503 (N_3503,N_1832,N_711);
nor U3504 (N_3504,N_896,N_661);
nand U3505 (N_3505,N_831,N_1054);
xor U3506 (N_3506,N_303,N_2410);
and U3507 (N_3507,N_1015,N_1731);
nor U3508 (N_3508,N_2282,N_1223);
or U3509 (N_3509,N_1062,N_1868);
nand U3510 (N_3510,N_1972,N_2460);
xor U3511 (N_3511,N_1106,N_1122);
or U3512 (N_3512,N_140,N_1904);
or U3513 (N_3513,N_39,N_1521);
and U3514 (N_3514,N_580,N_780);
xnor U3515 (N_3515,N_1955,N_1474);
and U3516 (N_3516,N_1910,N_1932);
and U3517 (N_3517,N_981,N_2007);
nor U3518 (N_3518,N_2421,N_839);
xor U3519 (N_3519,N_499,N_650);
and U3520 (N_3520,N_2172,N_1765);
and U3521 (N_3521,N_1311,N_1817);
and U3522 (N_3522,N_2360,N_75);
or U3523 (N_3523,N_2444,N_1758);
xnor U3524 (N_3524,N_859,N_933);
and U3525 (N_3525,N_566,N_628);
and U3526 (N_3526,N_2481,N_1988);
and U3527 (N_3527,N_1089,N_1459);
and U3528 (N_3528,N_664,N_1912);
and U3529 (N_3529,N_183,N_1010);
and U3530 (N_3530,N_7,N_81);
or U3531 (N_3531,N_481,N_1377);
or U3532 (N_3532,N_124,N_582);
xor U3533 (N_3533,N_2428,N_2377);
nand U3534 (N_3534,N_917,N_590);
nand U3535 (N_3535,N_765,N_1182);
xnor U3536 (N_3536,N_768,N_1801);
and U3537 (N_3537,N_1900,N_810);
nor U3538 (N_3538,N_1420,N_1720);
nand U3539 (N_3539,N_1903,N_1848);
xor U3540 (N_3540,N_1866,N_791);
and U3541 (N_3541,N_521,N_927);
or U3542 (N_3542,N_534,N_203);
or U3543 (N_3543,N_2344,N_2011);
xnor U3544 (N_3544,N_1458,N_804);
or U3545 (N_3545,N_1550,N_139);
or U3546 (N_3546,N_2496,N_2142);
or U3547 (N_3547,N_339,N_2455);
or U3548 (N_3548,N_60,N_1523);
nor U3549 (N_3549,N_890,N_2150);
and U3550 (N_3550,N_85,N_2131);
nand U3551 (N_3551,N_1478,N_2176);
and U3552 (N_3552,N_1793,N_356);
nor U3553 (N_3553,N_693,N_1345);
or U3554 (N_3554,N_740,N_355);
and U3555 (N_3555,N_262,N_585);
or U3556 (N_3556,N_2159,N_800);
xor U3557 (N_3557,N_125,N_1115);
nor U3558 (N_3558,N_1813,N_391);
nor U3559 (N_3559,N_1164,N_1609);
and U3560 (N_3560,N_469,N_1378);
nand U3561 (N_3561,N_1222,N_90);
and U3562 (N_3562,N_2006,N_1336);
or U3563 (N_3563,N_2477,N_23);
and U3564 (N_3564,N_1705,N_113);
nor U3565 (N_3565,N_266,N_909);
xnor U3566 (N_3566,N_387,N_2178);
and U3567 (N_3567,N_349,N_1360);
and U3568 (N_3568,N_523,N_1933);
and U3569 (N_3569,N_2213,N_2487);
and U3570 (N_3570,N_1076,N_1234);
nand U3571 (N_3571,N_428,N_1727);
nand U3572 (N_3572,N_2089,N_1184);
nand U3573 (N_3573,N_1841,N_1);
nor U3574 (N_3574,N_1461,N_274);
and U3575 (N_3575,N_1246,N_1283);
or U3576 (N_3576,N_857,N_1308);
and U3577 (N_3577,N_238,N_1931);
nand U3578 (N_3578,N_1827,N_1193);
or U3579 (N_3579,N_1510,N_538);
nor U3580 (N_3580,N_1215,N_653);
and U3581 (N_3581,N_63,N_1300);
nor U3582 (N_3582,N_941,N_918);
nand U3583 (N_3583,N_1806,N_423);
or U3584 (N_3584,N_993,N_1173);
xor U3585 (N_3585,N_1571,N_1777);
xnor U3586 (N_3586,N_830,N_632);
and U3587 (N_3587,N_132,N_64);
xnor U3588 (N_3588,N_1102,N_2223);
and U3589 (N_3589,N_73,N_147);
and U3590 (N_3590,N_57,N_922);
xor U3591 (N_3591,N_2140,N_2324);
nor U3592 (N_3592,N_737,N_700);
and U3593 (N_3593,N_2323,N_95);
nor U3594 (N_3594,N_2461,N_606);
and U3595 (N_3595,N_1266,N_277);
or U3596 (N_3596,N_1339,N_68);
xnor U3597 (N_3597,N_1529,N_1874);
and U3598 (N_3598,N_2434,N_721);
xor U3599 (N_3599,N_396,N_642);
nor U3600 (N_3600,N_814,N_903);
xor U3601 (N_3601,N_2047,N_656);
nand U3602 (N_3602,N_1934,N_165);
nand U3603 (N_3603,N_1211,N_925);
and U3604 (N_3604,N_542,N_1198);
nand U3605 (N_3605,N_2478,N_1372);
or U3606 (N_3606,N_31,N_1738);
nand U3607 (N_3607,N_605,N_2126);
nand U3608 (N_3608,N_204,N_2208);
nand U3609 (N_3609,N_911,N_479);
nand U3610 (N_3610,N_2020,N_665);
or U3611 (N_3611,N_860,N_730);
nor U3612 (N_3612,N_2491,N_808);
and U3613 (N_3613,N_1435,N_1634);
nor U3614 (N_3614,N_1785,N_2125);
or U3615 (N_3615,N_1950,N_739);
nor U3616 (N_3616,N_2245,N_122);
nor U3617 (N_3617,N_1256,N_1517);
nor U3618 (N_3618,N_1243,N_820);
nand U3619 (N_3619,N_350,N_2346);
nand U3620 (N_3620,N_1579,N_1280);
and U3621 (N_3621,N_483,N_867);
nand U3622 (N_3622,N_1097,N_211);
or U3623 (N_3623,N_1739,N_1323);
nor U3624 (N_3624,N_892,N_1797);
and U3625 (N_3625,N_620,N_803);
or U3626 (N_3626,N_2115,N_89);
xor U3627 (N_3627,N_1749,N_2380);
and U3628 (N_3628,N_2106,N_1009);
xnor U3629 (N_3629,N_980,N_1359);
nor U3630 (N_3630,N_233,N_2366);
nor U3631 (N_3631,N_1253,N_2333);
nor U3632 (N_3632,N_668,N_2373);
xor U3633 (N_3633,N_1261,N_1884);
nand U3634 (N_3634,N_2367,N_296);
and U3635 (N_3635,N_1576,N_1792);
nand U3636 (N_3636,N_2136,N_2386);
xnor U3637 (N_3637,N_811,N_1722);
or U3638 (N_3638,N_2043,N_1125);
nor U3639 (N_3639,N_1036,N_334);
or U3640 (N_3640,N_454,N_1620);
and U3641 (N_3641,N_1180,N_599);
nor U3642 (N_3642,N_2368,N_338);
xor U3643 (N_3643,N_2425,N_784);
xnor U3644 (N_3644,N_2200,N_402);
nor U3645 (N_3645,N_792,N_2259);
xnor U3646 (N_3646,N_681,N_210);
xor U3647 (N_3647,N_848,N_2040);
nand U3648 (N_3648,N_25,N_609);
nor U3649 (N_3649,N_1999,N_1876);
or U3650 (N_3650,N_150,N_161);
and U3651 (N_3651,N_2484,N_411);
xor U3652 (N_3652,N_607,N_321);
nor U3653 (N_3653,N_1669,N_1513);
xnor U3654 (N_3654,N_1790,N_207);
xor U3655 (N_3655,N_76,N_1446);
xnor U3656 (N_3656,N_625,N_1165);
and U3657 (N_3657,N_367,N_1023);
nor U3658 (N_3658,N_1269,N_900);
xor U3659 (N_3659,N_2261,N_1854);
nand U3660 (N_3660,N_1238,N_284);
and U3661 (N_3661,N_517,N_1202);
xnor U3662 (N_3662,N_904,N_657);
and U3663 (N_3663,N_2001,N_133);
or U3664 (N_3664,N_474,N_667);
nor U3665 (N_3665,N_894,N_1456);
xor U3666 (N_3666,N_907,N_853);
or U3667 (N_3667,N_1472,N_2283);
or U3668 (N_3668,N_2431,N_2286);
nor U3669 (N_3669,N_746,N_2214);
nor U3670 (N_3670,N_2050,N_2019);
nand U3671 (N_3671,N_2086,N_1893);
nand U3672 (N_3672,N_335,N_106);
or U3673 (N_3673,N_235,N_1217);
nand U3674 (N_3674,N_2236,N_236);
xor U3675 (N_3675,N_533,N_1386);
xnor U3676 (N_3676,N_22,N_528);
or U3677 (N_3677,N_431,N_840);
nand U3678 (N_3678,N_854,N_2167);
nor U3679 (N_3679,N_2409,N_1417);
nand U3680 (N_3680,N_1546,N_2154);
and U3681 (N_3681,N_394,N_2198);
xor U3682 (N_3682,N_1540,N_1639);
or U3683 (N_3683,N_1596,N_195);
nor U3684 (N_3684,N_1480,N_1049);
and U3685 (N_3685,N_2205,N_2186);
and U3686 (N_3686,N_878,N_1029);
and U3687 (N_3687,N_496,N_658);
xnor U3688 (N_3688,N_2251,N_160);
and U3689 (N_3689,N_1980,N_359);
or U3690 (N_3690,N_2162,N_1935);
nor U3691 (N_3691,N_1699,N_626);
or U3692 (N_3692,N_2174,N_1301);
xnor U3693 (N_3693,N_404,N_151);
nor U3694 (N_3694,N_1092,N_672);
or U3695 (N_3695,N_378,N_2448);
or U3696 (N_3696,N_2211,N_1501);
nor U3697 (N_3697,N_1194,N_1058);
nand U3698 (N_3698,N_2388,N_1677);
nand U3699 (N_3699,N_720,N_1628);
nor U3700 (N_3700,N_936,N_47);
and U3701 (N_3701,N_1303,N_285);
nor U3702 (N_3702,N_998,N_1951);
nand U3703 (N_3703,N_2038,N_1346);
or U3704 (N_3704,N_2341,N_1600);
or U3705 (N_3705,N_1271,N_1858);
nand U3706 (N_3706,N_1027,N_1055);
nor U3707 (N_3707,N_513,N_1503);
and U3708 (N_3708,N_2310,N_2084);
nand U3709 (N_3709,N_649,N_1477);
nor U3710 (N_3710,N_1168,N_1157);
nand U3711 (N_3711,N_2456,N_1137);
nor U3712 (N_3712,N_1915,N_1840);
or U3713 (N_3713,N_1971,N_104);
xor U3714 (N_3714,N_1264,N_1108);
or U3715 (N_3715,N_1757,N_259);
nand U3716 (N_3716,N_600,N_1096);
or U3717 (N_3717,N_2229,N_1911);
nand U3718 (N_3718,N_265,N_385);
xor U3719 (N_3719,N_446,N_955);
xor U3720 (N_3720,N_2014,N_1411);
xnor U3721 (N_3721,N_964,N_1618);
and U3722 (N_3722,N_644,N_2382);
nor U3723 (N_3723,N_1306,N_805);
or U3724 (N_3724,N_691,N_2369);
and U3725 (N_3725,N_348,N_2216);
nor U3726 (N_3726,N_714,N_826);
nand U3727 (N_3727,N_2104,N_92);
nand U3728 (N_3728,N_1642,N_2365);
or U3729 (N_3729,N_163,N_979);
and U3730 (N_3730,N_1479,N_2113);
nand U3731 (N_3731,N_1042,N_1305);
or U3732 (N_3732,N_529,N_97);
and U3733 (N_3733,N_1366,N_94);
nor U3734 (N_3734,N_1138,N_777);
nor U3735 (N_3735,N_683,N_634);
nand U3736 (N_3736,N_1309,N_624);
nor U3737 (N_3737,N_375,N_1351);
nand U3738 (N_3738,N_1158,N_2335);
or U3739 (N_3739,N_788,N_222);
nand U3740 (N_3740,N_2177,N_524);
nand U3741 (N_3741,N_2389,N_1652);
xor U3742 (N_3742,N_817,N_1085);
or U3743 (N_3743,N_949,N_1686);
xor U3744 (N_3744,N_893,N_1033);
nand U3745 (N_3745,N_589,N_343);
nor U3746 (N_3746,N_1095,N_1664);
and U3747 (N_3747,N_2309,N_943);
nor U3748 (N_3748,N_818,N_790);
nand U3749 (N_3749,N_874,N_142);
xnor U3750 (N_3750,N_122,N_1741);
nand U3751 (N_3751,N_1095,N_716);
and U3752 (N_3752,N_882,N_1487);
or U3753 (N_3753,N_1937,N_1425);
and U3754 (N_3754,N_2365,N_1968);
or U3755 (N_3755,N_2019,N_380);
and U3756 (N_3756,N_586,N_1215);
and U3757 (N_3757,N_164,N_2492);
nor U3758 (N_3758,N_288,N_1098);
nor U3759 (N_3759,N_1913,N_1430);
or U3760 (N_3760,N_382,N_1303);
xor U3761 (N_3761,N_1151,N_656);
nand U3762 (N_3762,N_1108,N_1838);
nor U3763 (N_3763,N_624,N_472);
xor U3764 (N_3764,N_2423,N_1500);
or U3765 (N_3765,N_2223,N_20);
nand U3766 (N_3766,N_1236,N_1010);
or U3767 (N_3767,N_859,N_766);
nor U3768 (N_3768,N_1899,N_1437);
xnor U3769 (N_3769,N_743,N_2270);
or U3770 (N_3770,N_344,N_1192);
and U3771 (N_3771,N_72,N_592);
or U3772 (N_3772,N_639,N_940);
xor U3773 (N_3773,N_1232,N_2023);
and U3774 (N_3774,N_606,N_1701);
and U3775 (N_3775,N_131,N_553);
nor U3776 (N_3776,N_385,N_2379);
xor U3777 (N_3777,N_768,N_1122);
xor U3778 (N_3778,N_1989,N_2098);
nor U3779 (N_3779,N_1675,N_6);
nor U3780 (N_3780,N_1571,N_1109);
nor U3781 (N_3781,N_1310,N_288);
or U3782 (N_3782,N_940,N_172);
nor U3783 (N_3783,N_1108,N_1366);
nand U3784 (N_3784,N_90,N_891);
and U3785 (N_3785,N_198,N_1168);
and U3786 (N_3786,N_212,N_381);
or U3787 (N_3787,N_948,N_730);
xnor U3788 (N_3788,N_175,N_490);
xnor U3789 (N_3789,N_136,N_2228);
nor U3790 (N_3790,N_1646,N_2200);
nor U3791 (N_3791,N_2215,N_943);
nand U3792 (N_3792,N_1740,N_333);
and U3793 (N_3793,N_1908,N_141);
nor U3794 (N_3794,N_1919,N_1622);
nand U3795 (N_3795,N_187,N_1587);
nor U3796 (N_3796,N_486,N_2150);
nor U3797 (N_3797,N_1356,N_228);
xor U3798 (N_3798,N_1851,N_1866);
xor U3799 (N_3799,N_2356,N_2322);
nand U3800 (N_3800,N_524,N_1964);
and U3801 (N_3801,N_220,N_797);
xor U3802 (N_3802,N_1222,N_2342);
or U3803 (N_3803,N_2006,N_560);
nor U3804 (N_3804,N_1902,N_1781);
and U3805 (N_3805,N_2402,N_1441);
nor U3806 (N_3806,N_1430,N_936);
xor U3807 (N_3807,N_2384,N_757);
xor U3808 (N_3808,N_404,N_1123);
nor U3809 (N_3809,N_786,N_2455);
or U3810 (N_3810,N_2057,N_850);
and U3811 (N_3811,N_725,N_1764);
and U3812 (N_3812,N_2194,N_2355);
or U3813 (N_3813,N_2078,N_180);
or U3814 (N_3814,N_1029,N_1877);
or U3815 (N_3815,N_51,N_2471);
nor U3816 (N_3816,N_807,N_1651);
nand U3817 (N_3817,N_1209,N_134);
or U3818 (N_3818,N_1115,N_19);
nand U3819 (N_3819,N_1037,N_595);
xor U3820 (N_3820,N_829,N_2490);
nand U3821 (N_3821,N_818,N_861);
nand U3822 (N_3822,N_361,N_1216);
or U3823 (N_3823,N_746,N_1145);
nand U3824 (N_3824,N_997,N_821);
or U3825 (N_3825,N_697,N_2116);
nand U3826 (N_3826,N_995,N_139);
xor U3827 (N_3827,N_2402,N_2384);
or U3828 (N_3828,N_744,N_1642);
xnor U3829 (N_3829,N_982,N_2266);
nor U3830 (N_3830,N_819,N_913);
xnor U3831 (N_3831,N_900,N_2333);
or U3832 (N_3832,N_2066,N_646);
or U3833 (N_3833,N_2488,N_1505);
or U3834 (N_3834,N_260,N_2209);
nand U3835 (N_3835,N_2416,N_2065);
xnor U3836 (N_3836,N_2152,N_56);
nand U3837 (N_3837,N_2069,N_1236);
xor U3838 (N_3838,N_389,N_1526);
nor U3839 (N_3839,N_97,N_796);
and U3840 (N_3840,N_677,N_2185);
xor U3841 (N_3841,N_74,N_1958);
nor U3842 (N_3842,N_1737,N_1892);
nor U3843 (N_3843,N_1384,N_280);
nor U3844 (N_3844,N_948,N_2403);
nor U3845 (N_3845,N_962,N_1765);
nor U3846 (N_3846,N_938,N_1002);
nand U3847 (N_3847,N_1828,N_2070);
and U3848 (N_3848,N_595,N_2105);
nand U3849 (N_3849,N_1976,N_1974);
nand U3850 (N_3850,N_1992,N_1402);
nand U3851 (N_3851,N_54,N_1275);
and U3852 (N_3852,N_1447,N_1738);
and U3853 (N_3853,N_1077,N_1346);
and U3854 (N_3854,N_1670,N_2447);
or U3855 (N_3855,N_1993,N_1677);
nor U3856 (N_3856,N_2264,N_2466);
and U3857 (N_3857,N_1404,N_2487);
or U3858 (N_3858,N_1506,N_1309);
or U3859 (N_3859,N_1251,N_1012);
xor U3860 (N_3860,N_1693,N_1184);
and U3861 (N_3861,N_557,N_1735);
or U3862 (N_3862,N_51,N_1910);
and U3863 (N_3863,N_2371,N_944);
xnor U3864 (N_3864,N_1604,N_1006);
nor U3865 (N_3865,N_2363,N_381);
or U3866 (N_3866,N_1684,N_430);
nor U3867 (N_3867,N_1316,N_765);
nand U3868 (N_3868,N_1257,N_2090);
xnor U3869 (N_3869,N_1691,N_885);
xnor U3870 (N_3870,N_466,N_1246);
xnor U3871 (N_3871,N_1219,N_989);
and U3872 (N_3872,N_1729,N_515);
nand U3873 (N_3873,N_1982,N_976);
xnor U3874 (N_3874,N_807,N_101);
xnor U3875 (N_3875,N_373,N_655);
nand U3876 (N_3876,N_815,N_2060);
or U3877 (N_3877,N_354,N_814);
nor U3878 (N_3878,N_1150,N_299);
nand U3879 (N_3879,N_1992,N_2003);
xor U3880 (N_3880,N_182,N_11);
nor U3881 (N_3881,N_1480,N_1013);
nand U3882 (N_3882,N_1320,N_1951);
and U3883 (N_3883,N_312,N_1129);
xor U3884 (N_3884,N_340,N_456);
nor U3885 (N_3885,N_542,N_1822);
nor U3886 (N_3886,N_164,N_375);
and U3887 (N_3887,N_946,N_94);
or U3888 (N_3888,N_1188,N_1567);
and U3889 (N_3889,N_139,N_2293);
xnor U3890 (N_3890,N_2208,N_1860);
or U3891 (N_3891,N_1217,N_1051);
xor U3892 (N_3892,N_2030,N_1751);
and U3893 (N_3893,N_531,N_816);
nor U3894 (N_3894,N_2031,N_1057);
nand U3895 (N_3895,N_702,N_66);
nor U3896 (N_3896,N_881,N_1296);
or U3897 (N_3897,N_2190,N_1670);
and U3898 (N_3898,N_669,N_123);
or U3899 (N_3899,N_763,N_1566);
and U3900 (N_3900,N_791,N_448);
xor U3901 (N_3901,N_2429,N_1157);
xnor U3902 (N_3902,N_1449,N_67);
xnor U3903 (N_3903,N_1448,N_1347);
and U3904 (N_3904,N_437,N_472);
nand U3905 (N_3905,N_1387,N_1486);
or U3906 (N_3906,N_2432,N_607);
nand U3907 (N_3907,N_1709,N_219);
or U3908 (N_3908,N_1909,N_531);
xnor U3909 (N_3909,N_1767,N_2280);
nor U3910 (N_3910,N_1348,N_1655);
and U3911 (N_3911,N_1274,N_1627);
and U3912 (N_3912,N_461,N_555);
and U3913 (N_3913,N_2225,N_759);
and U3914 (N_3914,N_2259,N_1194);
xor U3915 (N_3915,N_1270,N_2349);
and U3916 (N_3916,N_684,N_1515);
and U3917 (N_3917,N_289,N_981);
nor U3918 (N_3918,N_1016,N_1853);
nand U3919 (N_3919,N_790,N_1751);
nand U3920 (N_3920,N_1767,N_1980);
xnor U3921 (N_3921,N_595,N_12);
and U3922 (N_3922,N_835,N_1671);
nand U3923 (N_3923,N_1594,N_1207);
nor U3924 (N_3924,N_119,N_632);
or U3925 (N_3925,N_2240,N_1550);
xnor U3926 (N_3926,N_762,N_2240);
nor U3927 (N_3927,N_942,N_1617);
xnor U3928 (N_3928,N_881,N_1630);
or U3929 (N_3929,N_2272,N_612);
nand U3930 (N_3930,N_1901,N_1129);
nand U3931 (N_3931,N_552,N_63);
xor U3932 (N_3932,N_2054,N_2014);
and U3933 (N_3933,N_1048,N_1482);
xnor U3934 (N_3934,N_1152,N_472);
or U3935 (N_3935,N_489,N_1592);
and U3936 (N_3936,N_2027,N_1061);
nand U3937 (N_3937,N_1913,N_2405);
nor U3938 (N_3938,N_1070,N_1773);
and U3939 (N_3939,N_1947,N_1919);
and U3940 (N_3940,N_1295,N_380);
nand U3941 (N_3941,N_1395,N_976);
nor U3942 (N_3942,N_2262,N_2354);
or U3943 (N_3943,N_867,N_603);
nor U3944 (N_3944,N_2222,N_880);
or U3945 (N_3945,N_2305,N_1301);
xor U3946 (N_3946,N_1599,N_522);
or U3947 (N_3947,N_2289,N_2146);
and U3948 (N_3948,N_950,N_2284);
and U3949 (N_3949,N_167,N_1956);
or U3950 (N_3950,N_1725,N_128);
and U3951 (N_3951,N_1973,N_2127);
and U3952 (N_3952,N_2192,N_1062);
nor U3953 (N_3953,N_1719,N_1110);
nor U3954 (N_3954,N_96,N_190);
and U3955 (N_3955,N_2230,N_681);
nand U3956 (N_3956,N_1622,N_546);
nor U3957 (N_3957,N_1433,N_63);
or U3958 (N_3958,N_2299,N_2325);
nor U3959 (N_3959,N_945,N_145);
nand U3960 (N_3960,N_2212,N_306);
xor U3961 (N_3961,N_156,N_2420);
nor U3962 (N_3962,N_1184,N_12);
nand U3963 (N_3963,N_23,N_1386);
nand U3964 (N_3964,N_2492,N_1663);
xor U3965 (N_3965,N_1151,N_1764);
and U3966 (N_3966,N_1459,N_2299);
and U3967 (N_3967,N_2023,N_120);
xor U3968 (N_3968,N_1702,N_267);
xnor U3969 (N_3969,N_2382,N_567);
xor U3970 (N_3970,N_2457,N_2023);
nand U3971 (N_3971,N_2128,N_725);
xnor U3972 (N_3972,N_1825,N_2011);
or U3973 (N_3973,N_636,N_147);
and U3974 (N_3974,N_2224,N_1896);
xnor U3975 (N_3975,N_632,N_2357);
and U3976 (N_3976,N_1978,N_1176);
or U3977 (N_3977,N_830,N_26);
nand U3978 (N_3978,N_341,N_1431);
xor U3979 (N_3979,N_1705,N_2467);
nand U3980 (N_3980,N_1693,N_718);
xnor U3981 (N_3981,N_1414,N_1096);
or U3982 (N_3982,N_173,N_1221);
nand U3983 (N_3983,N_1913,N_2057);
xor U3984 (N_3984,N_1437,N_706);
nor U3985 (N_3985,N_1856,N_96);
and U3986 (N_3986,N_1046,N_2279);
nor U3987 (N_3987,N_2090,N_2446);
nor U3988 (N_3988,N_993,N_970);
and U3989 (N_3989,N_2395,N_88);
nor U3990 (N_3990,N_1659,N_1670);
and U3991 (N_3991,N_2099,N_2192);
or U3992 (N_3992,N_1612,N_370);
nand U3993 (N_3993,N_1845,N_2138);
or U3994 (N_3994,N_1659,N_2296);
nand U3995 (N_3995,N_2024,N_159);
or U3996 (N_3996,N_119,N_2461);
and U3997 (N_3997,N_2397,N_1812);
and U3998 (N_3998,N_2324,N_1185);
and U3999 (N_3999,N_405,N_1958);
nor U4000 (N_4000,N_72,N_1401);
xnor U4001 (N_4001,N_991,N_2328);
nor U4002 (N_4002,N_173,N_1668);
or U4003 (N_4003,N_1170,N_396);
or U4004 (N_4004,N_1711,N_1593);
and U4005 (N_4005,N_2460,N_2493);
or U4006 (N_4006,N_1863,N_484);
and U4007 (N_4007,N_2139,N_1401);
and U4008 (N_4008,N_2205,N_1768);
or U4009 (N_4009,N_2142,N_721);
and U4010 (N_4010,N_145,N_58);
or U4011 (N_4011,N_1791,N_619);
nand U4012 (N_4012,N_636,N_363);
xnor U4013 (N_4013,N_2421,N_1856);
nor U4014 (N_4014,N_1549,N_2196);
nor U4015 (N_4015,N_1804,N_209);
and U4016 (N_4016,N_603,N_1293);
nor U4017 (N_4017,N_2034,N_1687);
or U4018 (N_4018,N_1261,N_1410);
xnor U4019 (N_4019,N_2343,N_2030);
or U4020 (N_4020,N_362,N_691);
xnor U4021 (N_4021,N_273,N_1239);
and U4022 (N_4022,N_449,N_1584);
nand U4023 (N_4023,N_2360,N_362);
and U4024 (N_4024,N_257,N_1443);
and U4025 (N_4025,N_2339,N_162);
and U4026 (N_4026,N_2104,N_1500);
xor U4027 (N_4027,N_1206,N_2160);
nand U4028 (N_4028,N_2365,N_838);
nand U4029 (N_4029,N_385,N_1563);
nor U4030 (N_4030,N_656,N_2310);
and U4031 (N_4031,N_1825,N_1598);
xor U4032 (N_4032,N_1128,N_1584);
or U4033 (N_4033,N_854,N_1280);
nand U4034 (N_4034,N_5,N_2273);
or U4035 (N_4035,N_878,N_1558);
and U4036 (N_4036,N_813,N_721);
nor U4037 (N_4037,N_1474,N_600);
nor U4038 (N_4038,N_1351,N_142);
xnor U4039 (N_4039,N_978,N_514);
or U4040 (N_4040,N_2324,N_1447);
and U4041 (N_4041,N_803,N_2174);
nor U4042 (N_4042,N_2426,N_1247);
or U4043 (N_4043,N_1664,N_1286);
and U4044 (N_4044,N_915,N_931);
nor U4045 (N_4045,N_1511,N_1788);
xnor U4046 (N_4046,N_1518,N_801);
nand U4047 (N_4047,N_256,N_1060);
nand U4048 (N_4048,N_1376,N_436);
nor U4049 (N_4049,N_2078,N_109);
or U4050 (N_4050,N_697,N_1880);
xnor U4051 (N_4051,N_665,N_1590);
nand U4052 (N_4052,N_1982,N_1205);
and U4053 (N_4053,N_1466,N_807);
xnor U4054 (N_4054,N_1438,N_342);
nor U4055 (N_4055,N_1611,N_2006);
nor U4056 (N_4056,N_117,N_2405);
nand U4057 (N_4057,N_196,N_766);
xor U4058 (N_4058,N_1923,N_2055);
nand U4059 (N_4059,N_109,N_672);
nand U4060 (N_4060,N_1170,N_2282);
or U4061 (N_4061,N_2357,N_1896);
nand U4062 (N_4062,N_1774,N_1078);
or U4063 (N_4063,N_828,N_192);
nor U4064 (N_4064,N_1708,N_2029);
nand U4065 (N_4065,N_1524,N_1770);
nor U4066 (N_4066,N_2485,N_275);
or U4067 (N_4067,N_1779,N_251);
and U4068 (N_4068,N_699,N_1774);
and U4069 (N_4069,N_1275,N_1088);
or U4070 (N_4070,N_432,N_2194);
nand U4071 (N_4071,N_696,N_2336);
nand U4072 (N_4072,N_2425,N_1512);
and U4073 (N_4073,N_632,N_1026);
nor U4074 (N_4074,N_1992,N_2425);
or U4075 (N_4075,N_1843,N_2408);
and U4076 (N_4076,N_2294,N_337);
xnor U4077 (N_4077,N_710,N_1654);
nor U4078 (N_4078,N_22,N_1427);
nor U4079 (N_4079,N_2289,N_590);
xor U4080 (N_4080,N_2398,N_672);
and U4081 (N_4081,N_1404,N_105);
xnor U4082 (N_4082,N_523,N_1395);
nor U4083 (N_4083,N_1737,N_2034);
xnor U4084 (N_4084,N_2291,N_2252);
and U4085 (N_4085,N_2341,N_17);
nand U4086 (N_4086,N_1778,N_1472);
xor U4087 (N_4087,N_1685,N_1774);
nor U4088 (N_4088,N_1625,N_2205);
nor U4089 (N_4089,N_1334,N_2114);
nand U4090 (N_4090,N_1484,N_2465);
nor U4091 (N_4091,N_317,N_1597);
nor U4092 (N_4092,N_1649,N_1747);
xnor U4093 (N_4093,N_954,N_1720);
and U4094 (N_4094,N_842,N_1350);
nor U4095 (N_4095,N_254,N_1102);
nand U4096 (N_4096,N_1261,N_1986);
nor U4097 (N_4097,N_2239,N_1699);
or U4098 (N_4098,N_1190,N_1639);
nor U4099 (N_4099,N_2389,N_990);
xor U4100 (N_4100,N_965,N_2198);
xor U4101 (N_4101,N_2396,N_2361);
nor U4102 (N_4102,N_194,N_542);
or U4103 (N_4103,N_47,N_1585);
and U4104 (N_4104,N_2362,N_1767);
nand U4105 (N_4105,N_152,N_1007);
nor U4106 (N_4106,N_1580,N_1890);
nor U4107 (N_4107,N_829,N_1729);
xnor U4108 (N_4108,N_2022,N_1250);
or U4109 (N_4109,N_2383,N_1867);
or U4110 (N_4110,N_1033,N_1057);
and U4111 (N_4111,N_1703,N_513);
or U4112 (N_4112,N_2465,N_265);
nand U4113 (N_4113,N_2460,N_2054);
and U4114 (N_4114,N_313,N_2314);
nor U4115 (N_4115,N_789,N_503);
nor U4116 (N_4116,N_501,N_2282);
nand U4117 (N_4117,N_2187,N_241);
nand U4118 (N_4118,N_403,N_1763);
nand U4119 (N_4119,N_1536,N_1865);
and U4120 (N_4120,N_2421,N_136);
or U4121 (N_4121,N_1621,N_2012);
or U4122 (N_4122,N_1358,N_644);
nor U4123 (N_4123,N_2282,N_1809);
nor U4124 (N_4124,N_1327,N_1301);
or U4125 (N_4125,N_409,N_1315);
or U4126 (N_4126,N_1302,N_1745);
and U4127 (N_4127,N_871,N_2496);
xnor U4128 (N_4128,N_1092,N_1759);
xnor U4129 (N_4129,N_1795,N_1934);
and U4130 (N_4130,N_1114,N_2078);
and U4131 (N_4131,N_513,N_698);
nand U4132 (N_4132,N_1406,N_1716);
nand U4133 (N_4133,N_2280,N_1507);
or U4134 (N_4134,N_762,N_2119);
xor U4135 (N_4135,N_2245,N_206);
nand U4136 (N_4136,N_1959,N_219);
and U4137 (N_4137,N_713,N_406);
or U4138 (N_4138,N_1798,N_1117);
and U4139 (N_4139,N_1062,N_2435);
xor U4140 (N_4140,N_1184,N_1991);
nand U4141 (N_4141,N_2162,N_171);
or U4142 (N_4142,N_1274,N_2182);
and U4143 (N_4143,N_1393,N_2045);
nand U4144 (N_4144,N_766,N_1347);
and U4145 (N_4145,N_627,N_920);
nand U4146 (N_4146,N_1406,N_1727);
or U4147 (N_4147,N_797,N_2380);
or U4148 (N_4148,N_187,N_1342);
nor U4149 (N_4149,N_1581,N_1588);
nor U4150 (N_4150,N_550,N_873);
or U4151 (N_4151,N_503,N_1252);
nand U4152 (N_4152,N_1958,N_28);
nand U4153 (N_4153,N_1351,N_1836);
and U4154 (N_4154,N_1167,N_2035);
and U4155 (N_4155,N_1475,N_411);
and U4156 (N_4156,N_1317,N_1016);
nor U4157 (N_4157,N_1758,N_183);
and U4158 (N_4158,N_2407,N_2252);
nor U4159 (N_4159,N_1828,N_1190);
nand U4160 (N_4160,N_2074,N_631);
nor U4161 (N_4161,N_1778,N_2118);
xnor U4162 (N_4162,N_2092,N_689);
xnor U4163 (N_4163,N_956,N_804);
or U4164 (N_4164,N_2404,N_437);
xor U4165 (N_4165,N_1354,N_1150);
nand U4166 (N_4166,N_1849,N_324);
or U4167 (N_4167,N_2273,N_1800);
nor U4168 (N_4168,N_333,N_827);
or U4169 (N_4169,N_327,N_1481);
xor U4170 (N_4170,N_1589,N_606);
nor U4171 (N_4171,N_457,N_207);
xnor U4172 (N_4172,N_682,N_2389);
nand U4173 (N_4173,N_555,N_2149);
and U4174 (N_4174,N_1550,N_2437);
nor U4175 (N_4175,N_2130,N_908);
nor U4176 (N_4176,N_2174,N_2023);
and U4177 (N_4177,N_20,N_1997);
xor U4178 (N_4178,N_976,N_1387);
nand U4179 (N_4179,N_2351,N_1090);
and U4180 (N_4180,N_38,N_67);
nand U4181 (N_4181,N_1104,N_185);
or U4182 (N_4182,N_1663,N_1880);
xnor U4183 (N_4183,N_1943,N_2472);
xnor U4184 (N_4184,N_29,N_459);
and U4185 (N_4185,N_2386,N_2470);
xnor U4186 (N_4186,N_1572,N_130);
nand U4187 (N_4187,N_1532,N_1951);
and U4188 (N_4188,N_950,N_2378);
nor U4189 (N_4189,N_1592,N_184);
xnor U4190 (N_4190,N_1180,N_1774);
nor U4191 (N_4191,N_1565,N_1001);
or U4192 (N_4192,N_1614,N_1527);
nand U4193 (N_4193,N_476,N_607);
and U4194 (N_4194,N_1588,N_1681);
nor U4195 (N_4195,N_77,N_11);
and U4196 (N_4196,N_794,N_1046);
xor U4197 (N_4197,N_392,N_256);
nor U4198 (N_4198,N_1569,N_1071);
and U4199 (N_4199,N_32,N_2444);
nor U4200 (N_4200,N_982,N_1268);
and U4201 (N_4201,N_1592,N_1128);
nand U4202 (N_4202,N_1199,N_951);
xnor U4203 (N_4203,N_216,N_707);
xnor U4204 (N_4204,N_1794,N_552);
and U4205 (N_4205,N_437,N_2490);
xor U4206 (N_4206,N_923,N_1265);
xnor U4207 (N_4207,N_1427,N_1085);
nor U4208 (N_4208,N_2437,N_694);
nand U4209 (N_4209,N_846,N_99);
or U4210 (N_4210,N_255,N_1174);
or U4211 (N_4211,N_480,N_64);
nor U4212 (N_4212,N_2077,N_558);
and U4213 (N_4213,N_837,N_690);
xnor U4214 (N_4214,N_239,N_1569);
xor U4215 (N_4215,N_1895,N_2457);
xor U4216 (N_4216,N_2451,N_2106);
and U4217 (N_4217,N_0,N_1951);
nand U4218 (N_4218,N_1560,N_2499);
xnor U4219 (N_4219,N_2413,N_1150);
and U4220 (N_4220,N_784,N_1369);
nor U4221 (N_4221,N_1996,N_553);
or U4222 (N_4222,N_682,N_1188);
nor U4223 (N_4223,N_2334,N_551);
xor U4224 (N_4224,N_94,N_281);
or U4225 (N_4225,N_255,N_1196);
nand U4226 (N_4226,N_2306,N_2381);
and U4227 (N_4227,N_2096,N_2485);
xor U4228 (N_4228,N_2458,N_1360);
or U4229 (N_4229,N_1084,N_1738);
and U4230 (N_4230,N_1660,N_897);
xnor U4231 (N_4231,N_1236,N_330);
nand U4232 (N_4232,N_2434,N_2439);
nand U4233 (N_4233,N_1520,N_580);
nor U4234 (N_4234,N_1203,N_2225);
nand U4235 (N_4235,N_1820,N_1907);
xor U4236 (N_4236,N_2408,N_189);
nor U4237 (N_4237,N_446,N_870);
and U4238 (N_4238,N_855,N_281);
xor U4239 (N_4239,N_915,N_436);
and U4240 (N_4240,N_203,N_1387);
or U4241 (N_4241,N_1849,N_1621);
xnor U4242 (N_4242,N_557,N_958);
xnor U4243 (N_4243,N_1170,N_829);
or U4244 (N_4244,N_1518,N_1731);
xnor U4245 (N_4245,N_1228,N_1789);
or U4246 (N_4246,N_195,N_2074);
or U4247 (N_4247,N_1010,N_1380);
xor U4248 (N_4248,N_2463,N_786);
and U4249 (N_4249,N_1059,N_49);
nor U4250 (N_4250,N_1549,N_1322);
or U4251 (N_4251,N_2456,N_2004);
nand U4252 (N_4252,N_1314,N_740);
nor U4253 (N_4253,N_867,N_670);
xor U4254 (N_4254,N_1927,N_781);
xnor U4255 (N_4255,N_1801,N_2315);
or U4256 (N_4256,N_86,N_1890);
and U4257 (N_4257,N_2007,N_1004);
and U4258 (N_4258,N_467,N_643);
and U4259 (N_4259,N_2233,N_1646);
nor U4260 (N_4260,N_827,N_1746);
nand U4261 (N_4261,N_2352,N_1424);
nand U4262 (N_4262,N_1868,N_2481);
xnor U4263 (N_4263,N_1826,N_1837);
and U4264 (N_4264,N_209,N_1054);
xnor U4265 (N_4265,N_578,N_14);
nand U4266 (N_4266,N_1310,N_573);
or U4267 (N_4267,N_2419,N_1632);
nand U4268 (N_4268,N_2288,N_229);
nor U4269 (N_4269,N_34,N_2328);
or U4270 (N_4270,N_1915,N_1246);
and U4271 (N_4271,N_268,N_1780);
nor U4272 (N_4272,N_564,N_716);
nor U4273 (N_4273,N_2060,N_1821);
xor U4274 (N_4274,N_596,N_1084);
xnor U4275 (N_4275,N_1355,N_1847);
or U4276 (N_4276,N_2351,N_1609);
nand U4277 (N_4277,N_1212,N_1879);
nor U4278 (N_4278,N_1173,N_1899);
nor U4279 (N_4279,N_639,N_268);
xor U4280 (N_4280,N_1391,N_1480);
xor U4281 (N_4281,N_68,N_1640);
nand U4282 (N_4282,N_1284,N_1700);
or U4283 (N_4283,N_574,N_2292);
nor U4284 (N_4284,N_603,N_2170);
xor U4285 (N_4285,N_264,N_833);
xnor U4286 (N_4286,N_1093,N_56);
or U4287 (N_4287,N_2357,N_353);
or U4288 (N_4288,N_986,N_1893);
nand U4289 (N_4289,N_289,N_628);
nor U4290 (N_4290,N_737,N_688);
or U4291 (N_4291,N_1455,N_2431);
xnor U4292 (N_4292,N_2321,N_1038);
xor U4293 (N_4293,N_1917,N_948);
xnor U4294 (N_4294,N_2445,N_2190);
or U4295 (N_4295,N_1254,N_1123);
and U4296 (N_4296,N_2294,N_810);
nand U4297 (N_4297,N_2479,N_1115);
or U4298 (N_4298,N_2101,N_391);
nand U4299 (N_4299,N_1722,N_2347);
or U4300 (N_4300,N_1947,N_2423);
nor U4301 (N_4301,N_125,N_881);
or U4302 (N_4302,N_110,N_1592);
and U4303 (N_4303,N_1819,N_2189);
nor U4304 (N_4304,N_298,N_1470);
nand U4305 (N_4305,N_2483,N_986);
and U4306 (N_4306,N_576,N_2437);
nand U4307 (N_4307,N_1039,N_1766);
or U4308 (N_4308,N_1391,N_1052);
xor U4309 (N_4309,N_2181,N_778);
or U4310 (N_4310,N_959,N_827);
or U4311 (N_4311,N_1880,N_1207);
nand U4312 (N_4312,N_1176,N_1079);
nand U4313 (N_4313,N_2161,N_173);
nand U4314 (N_4314,N_2395,N_1236);
nor U4315 (N_4315,N_2141,N_1891);
or U4316 (N_4316,N_2347,N_931);
nand U4317 (N_4317,N_86,N_981);
nand U4318 (N_4318,N_1058,N_168);
and U4319 (N_4319,N_1139,N_1922);
xnor U4320 (N_4320,N_1791,N_1570);
nand U4321 (N_4321,N_2318,N_111);
nor U4322 (N_4322,N_2396,N_699);
and U4323 (N_4323,N_1839,N_1287);
or U4324 (N_4324,N_1039,N_799);
nand U4325 (N_4325,N_2396,N_298);
and U4326 (N_4326,N_135,N_1974);
nor U4327 (N_4327,N_1942,N_2247);
or U4328 (N_4328,N_9,N_113);
nand U4329 (N_4329,N_1980,N_164);
nor U4330 (N_4330,N_1590,N_695);
nor U4331 (N_4331,N_2266,N_1736);
xnor U4332 (N_4332,N_771,N_400);
nor U4333 (N_4333,N_373,N_2454);
and U4334 (N_4334,N_524,N_1376);
xor U4335 (N_4335,N_1425,N_2443);
nor U4336 (N_4336,N_190,N_106);
xor U4337 (N_4337,N_1020,N_106);
nand U4338 (N_4338,N_1336,N_1956);
xnor U4339 (N_4339,N_478,N_667);
xor U4340 (N_4340,N_1751,N_1485);
or U4341 (N_4341,N_1495,N_1419);
or U4342 (N_4342,N_980,N_777);
or U4343 (N_4343,N_870,N_162);
xnor U4344 (N_4344,N_244,N_1328);
or U4345 (N_4345,N_1499,N_508);
xor U4346 (N_4346,N_51,N_2058);
and U4347 (N_4347,N_1440,N_338);
or U4348 (N_4348,N_1852,N_1552);
or U4349 (N_4349,N_397,N_335);
and U4350 (N_4350,N_2288,N_91);
and U4351 (N_4351,N_2214,N_1708);
nor U4352 (N_4352,N_878,N_285);
xor U4353 (N_4353,N_461,N_2492);
nor U4354 (N_4354,N_1435,N_2126);
and U4355 (N_4355,N_611,N_793);
nor U4356 (N_4356,N_1698,N_464);
and U4357 (N_4357,N_209,N_376);
nand U4358 (N_4358,N_1525,N_2401);
and U4359 (N_4359,N_1557,N_1880);
xor U4360 (N_4360,N_1469,N_2459);
nor U4361 (N_4361,N_68,N_1382);
nor U4362 (N_4362,N_145,N_486);
nor U4363 (N_4363,N_1851,N_2364);
and U4364 (N_4364,N_1621,N_2466);
or U4365 (N_4365,N_1465,N_772);
and U4366 (N_4366,N_301,N_2414);
nand U4367 (N_4367,N_2427,N_211);
or U4368 (N_4368,N_1511,N_498);
or U4369 (N_4369,N_2103,N_1707);
nand U4370 (N_4370,N_671,N_1366);
xnor U4371 (N_4371,N_2353,N_1818);
and U4372 (N_4372,N_1127,N_369);
xnor U4373 (N_4373,N_388,N_2252);
xor U4374 (N_4374,N_1954,N_325);
nand U4375 (N_4375,N_707,N_1647);
or U4376 (N_4376,N_601,N_563);
nor U4377 (N_4377,N_2008,N_2142);
nand U4378 (N_4378,N_134,N_1516);
xor U4379 (N_4379,N_1537,N_834);
xnor U4380 (N_4380,N_803,N_1170);
nand U4381 (N_4381,N_827,N_1955);
nor U4382 (N_4382,N_840,N_709);
and U4383 (N_4383,N_946,N_1368);
or U4384 (N_4384,N_43,N_48);
or U4385 (N_4385,N_972,N_1710);
and U4386 (N_4386,N_962,N_1474);
xnor U4387 (N_4387,N_1721,N_2129);
xor U4388 (N_4388,N_1001,N_26);
xnor U4389 (N_4389,N_102,N_427);
nand U4390 (N_4390,N_2104,N_1490);
and U4391 (N_4391,N_507,N_2300);
nand U4392 (N_4392,N_1259,N_1674);
or U4393 (N_4393,N_507,N_602);
and U4394 (N_4394,N_1470,N_1427);
xnor U4395 (N_4395,N_2491,N_711);
xnor U4396 (N_4396,N_1398,N_1467);
or U4397 (N_4397,N_1055,N_2183);
and U4398 (N_4398,N_507,N_1844);
or U4399 (N_4399,N_2349,N_2320);
and U4400 (N_4400,N_1452,N_203);
and U4401 (N_4401,N_373,N_2311);
xnor U4402 (N_4402,N_2196,N_2465);
xor U4403 (N_4403,N_1972,N_1362);
nor U4404 (N_4404,N_597,N_144);
nand U4405 (N_4405,N_1629,N_1100);
xnor U4406 (N_4406,N_360,N_560);
nand U4407 (N_4407,N_77,N_885);
nand U4408 (N_4408,N_1824,N_1914);
or U4409 (N_4409,N_1152,N_233);
or U4410 (N_4410,N_759,N_515);
nor U4411 (N_4411,N_2287,N_718);
nand U4412 (N_4412,N_1739,N_623);
xor U4413 (N_4413,N_1677,N_1101);
nand U4414 (N_4414,N_1874,N_207);
xnor U4415 (N_4415,N_134,N_1926);
and U4416 (N_4416,N_510,N_2452);
nor U4417 (N_4417,N_384,N_235);
nor U4418 (N_4418,N_38,N_809);
xor U4419 (N_4419,N_1611,N_2478);
nand U4420 (N_4420,N_1818,N_1100);
and U4421 (N_4421,N_867,N_2128);
and U4422 (N_4422,N_964,N_1679);
nor U4423 (N_4423,N_374,N_112);
and U4424 (N_4424,N_1674,N_683);
xor U4425 (N_4425,N_1158,N_1287);
or U4426 (N_4426,N_94,N_440);
and U4427 (N_4427,N_1703,N_1831);
nand U4428 (N_4428,N_1567,N_1723);
nor U4429 (N_4429,N_2029,N_522);
nand U4430 (N_4430,N_2005,N_276);
or U4431 (N_4431,N_106,N_987);
xor U4432 (N_4432,N_1054,N_539);
and U4433 (N_4433,N_2289,N_1463);
nor U4434 (N_4434,N_1447,N_1793);
nor U4435 (N_4435,N_1743,N_564);
nand U4436 (N_4436,N_1732,N_2438);
xor U4437 (N_4437,N_2363,N_2085);
or U4438 (N_4438,N_1515,N_1895);
xor U4439 (N_4439,N_22,N_1796);
xor U4440 (N_4440,N_1809,N_1849);
or U4441 (N_4441,N_1990,N_46);
nor U4442 (N_4442,N_75,N_16);
nor U4443 (N_4443,N_1873,N_2120);
xnor U4444 (N_4444,N_1743,N_1054);
nor U4445 (N_4445,N_952,N_112);
or U4446 (N_4446,N_1413,N_1701);
nand U4447 (N_4447,N_2166,N_68);
xnor U4448 (N_4448,N_2222,N_1683);
or U4449 (N_4449,N_751,N_762);
nand U4450 (N_4450,N_2007,N_1268);
nand U4451 (N_4451,N_1083,N_2169);
xor U4452 (N_4452,N_649,N_1457);
and U4453 (N_4453,N_201,N_2118);
and U4454 (N_4454,N_2124,N_1004);
nor U4455 (N_4455,N_1063,N_562);
xor U4456 (N_4456,N_537,N_2048);
xor U4457 (N_4457,N_1938,N_1322);
xor U4458 (N_4458,N_2494,N_21);
nand U4459 (N_4459,N_945,N_2278);
xnor U4460 (N_4460,N_2087,N_965);
xor U4461 (N_4461,N_522,N_2216);
or U4462 (N_4462,N_1231,N_391);
xor U4463 (N_4463,N_2275,N_113);
and U4464 (N_4464,N_907,N_528);
nor U4465 (N_4465,N_532,N_1895);
or U4466 (N_4466,N_974,N_674);
nor U4467 (N_4467,N_2481,N_2111);
and U4468 (N_4468,N_2469,N_560);
nand U4469 (N_4469,N_1485,N_2479);
and U4470 (N_4470,N_1173,N_1262);
or U4471 (N_4471,N_2156,N_1155);
nand U4472 (N_4472,N_1428,N_394);
xor U4473 (N_4473,N_162,N_2111);
and U4474 (N_4474,N_1375,N_1489);
and U4475 (N_4475,N_2181,N_123);
nand U4476 (N_4476,N_1427,N_411);
nor U4477 (N_4477,N_1863,N_1550);
nand U4478 (N_4478,N_1538,N_2294);
xor U4479 (N_4479,N_1625,N_146);
or U4480 (N_4480,N_726,N_1432);
xor U4481 (N_4481,N_1549,N_1119);
and U4482 (N_4482,N_290,N_1750);
or U4483 (N_4483,N_1666,N_1474);
and U4484 (N_4484,N_345,N_1360);
or U4485 (N_4485,N_1671,N_1421);
xnor U4486 (N_4486,N_338,N_1804);
nor U4487 (N_4487,N_570,N_1833);
xnor U4488 (N_4488,N_553,N_2036);
nand U4489 (N_4489,N_1428,N_547);
or U4490 (N_4490,N_2174,N_1213);
or U4491 (N_4491,N_1626,N_2365);
or U4492 (N_4492,N_1641,N_2277);
or U4493 (N_4493,N_827,N_1022);
or U4494 (N_4494,N_562,N_2288);
or U4495 (N_4495,N_1711,N_556);
nor U4496 (N_4496,N_925,N_1370);
and U4497 (N_4497,N_2081,N_1711);
nand U4498 (N_4498,N_2450,N_1409);
nor U4499 (N_4499,N_411,N_692);
or U4500 (N_4500,N_484,N_1114);
nor U4501 (N_4501,N_1207,N_1171);
or U4502 (N_4502,N_833,N_633);
or U4503 (N_4503,N_1103,N_1521);
or U4504 (N_4504,N_2100,N_1518);
xnor U4505 (N_4505,N_401,N_2274);
and U4506 (N_4506,N_1528,N_699);
or U4507 (N_4507,N_464,N_945);
or U4508 (N_4508,N_1869,N_1428);
xor U4509 (N_4509,N_1203,N_1690);
xnor U4510 (N_4510,N_1626,N_1268);
or U4511 (N_4511,N_2076,N_1867);
and U4512 (N_4512,N_1822,N_445);
xnor U4513 (N_4513,N_396,N_1721);
nand U4514 (N_4514,N_595,N_2466);
xor U4515 (N_4515,N_2266,N_823);
or U4516 (N_4516,N_1190,N_1441);
xnor U4517 (N_4517,N_524,N_266);
or U4518 (N_4518,N_1981,N_2140);
xnor U4519 (N_4519,N_1923,N_29);
or U4520 (N_4520,N_2372,N_836);
xnor U4521 (N_4521,N_356,N_2286);
and U4522 (N_4522,N_2384,N_2463);
and U4523 (N_4523,N_2189,N_2068);
and U4524 (N_4524,N_2048,N_1544);
xor U4525 (N_4525,N_1766,N_1894);
nor U4526 (N_4526,N_867,N_325);
xnor U4527 (N_4527,N_105,N_1929);
nor U4528 (N_4528,N_1102,N_913);
or U4529 (N_4529,N_1021,N_485);
and U4530 (N_4530,N_1660,N_1976);
nor U4531 (N_4531,N_1763,N_1115);
nand U4532 (N_4532,N_2403,N_2179);
and U4533 (N_4533,N_1736,N_1602);
or U4534 (N_4534,N_13,N_158);
and U4535 (N_4535,N_1124,N_2271);
or U4536 (N_4536,N_2194,N_493);
xor U4537 (N_4537,N_408,N_305);
or U4538 (N_4538,N_989,N_1391);
nor U4539 (N_4539,N_1293,N_113);
or U4540 (N_4540,N_737,N_1066);
nor U4541 (N_4541,N_1623,N_163);
nor U4542 (N_4542,N_2003,N_301);
xnor U4543 (N_4543,N_679,N_1768);
xnor U4544 (N_4544,N_1860,N_2486);
nor U4545 (N_4545,N_2307,N_1379);
xor U4546 (N_4546,N_738,N_1960);
or U4547 (N_4547,N_346,N_779);
and U4548 (N_4548,N_1850,N_2266);
or U4549 (N_4549,N_186,N_1368);
or U4550 (N_4550,N_526,N_1976);
and U4551 (N_4551,N_915,N_1257);
nand U4552 (N_4552,N_1260,N_420);
or U4553 (N_4553,N_1306,N_1570);
nor U4554 (N_4554,N_2304,N_1139);
xor U4555 (N_4555,N_781,N_2080);
xnor U4556 (N_4556,N_957,N_747);
or U4557 (N_4557,N_242,N_2066);
nand U4558 (N_4558,N_341,N_743);
nor U4559 (N_4559,N_2244,N_1755);
and U4560 (N_4560,N_16,N_785);
nand U4561 (N_4561,N_795,N_248);
or U4562 (N_4562,N_455,N_1998);
nand U4563 (N_4563,N_254,N_2153);
nand U4564 (N_4564,N_173,N_1813);
nand U4565 (N_4565,N_1259,N_678);
nor U4566 (N_4566,N_937,N_1993);
nand U4567 (N_4567,N_855,N_254);
nor U4568 (N_4568,N_911,N_1573);
or U4569 (N_4569,N_1360,N_2466);
and U4570 (N_4570,N_1014,N_1358);
xor U4571 (N_4571,N_119,N_565);
and U4572 (N_4572,N_927,N_1906);
nor U4573 (N_4573,N_1616,N_215);
nor U4574 (N_4574,N_1267,N_572);
nor U4575 (N_4575,N_454,N_2229);
or U4576 (N_4576,N_2044,N_154);
and U4577 (N_4577,N_1008,N_1091);
or U4578 (N_4578,N_432,N_984);
xor U4579 (N_4579,N_1958,N_1605);
nand U4580 (N_4580,N_132,N_1989);
nor U4581 (N_4581,N_20,N_508);
nor U4582 (N_4582,N_583,N_1941);
xor U4583 (N_4583,N_951,N_2039);
or U4584 (N_4584,N_1446,N_957);
xor U4585 (N_4585,N_723,N_563);
and U4586 (N_4586,N_645,N_1486);
nand U4587 (N_4587,N_1667,N_1781);
and U4588 (N_4588,N_187,N_1292);
or U4589 (N_4589,N_1593,N_1579);
nand U4590 (N_4590,N_1494,N_2346);
and U4591 (N_4591,N_1024,N_2449);
xor U4592 (N_4592,N_1139,N_358);
and U4593 (N_4593,N_44,N_2411);
xor U4594 (N_4594,N_2299,N_760);
xor U4595 (N_4595,N_2143,N_943);
nand U4596 (N_4596,N_1746,N_1477);
or U4597 (N_4597,N_1825,N_2330);
xor U4598 (N_4598,N_1684,N_2132);
nor U4599 (N_4599,N_18,N_489);
nand U4600 (N_4600,N_692,N_1884);
xor U4601 (N_4601,N_1400,N_2446);
xnor U4602 (N_4602,N_580,N_2184);
xnor U4603 (N_4603,N_659,N_70);
xor U4604 (N_4604,N_1641,N_2205);
or U4605 (N_4605,N_1994,N_1031);
nand U4606 (N_4606,N_1712,N_684);
xor U4607 (N_4607,N_1300,N_2399);
or U4608 (N_4608,N_2181,N_1084);
or U4609 (N_4609,N_951,N_1261);
or U4610 (N_4610,N_295,N_557);
or U4611 (N_4611,N_587,N_281);
or U4612 (N_4612,N_740,N_1004);
xor U4613 (N_4613,N_2206,N_1428);
nand U4614 (N_4614,N_2169,N_660);
and U4615 (N_4615,N_2297,N_161);
nand U4616 (N_4616,N_846,N_698);
and U4617 (N_4617,N_437,N_2147);
xor U4618 (N_4618,N_1821,N_2290);
nand U4619 (N_4619,N_1544,N_753);
nand U4620 (N_4620,N_896,N_110);
xnor U4621 (N_4621,N_1364,N_2436);
nor U4622 (N_4622,N_365,N_1976);
xor U4623 (N_4623,N_831,N_939);
xor U4624 (N_4624,N_845,N_1493);
nand U4625 (N_4625,N_420,N_2147);
xnor U4626 (N_4626,N_1708,N_1100);
nand U4627 (N_4627,N_1515,N_337);
nor U4628 (N_4628,N_1357,N_1617);
or U4629 (N_4629,N_1687,N_2028);
xnor U4630 (N_4630,N_1397,N_1328);
and U4631 (N_4631,N_1356,N_478);
or U4632 (N_4632,N_340,N_24);
or U4633 (N_4633,N_1240,N_1527);
nor U4634 (N_4634,N_1353,N_341);
xor U4635 (N_4635,N_1498,N_1670);
nand U4636 (N_4636,N_1573,N_649);
and U4637 (N_4637,N_759,N_2335);
or U4638 (N_4638,N_2322,N_773);
nand U4639 (N_4639,N_2324,N_552);
xnor U4640 (N_4640,N_673,N_1815);
and U4641 (N_4641,N_715,N_1727);
or U4642 (N_4642,N_884,N_736);
and U4643 (N_4643,N_2073,N_381);
and U4644 (N_4644,N_917,N_2422);
and U4645 (N_4645,N_942,N_1785);
or U4646 (N_4646,N_1259,N_796);
nand U4647 (N_4647,N_1294,N_1848);
nor U4648 (N_4648,N_1004,N_1532);
or U4649 (N_4649,N_2318,N_193);
nand U4650 (N_4650,N_26,N_1292);
nand U4651 (N_4651,N_74,N_120);
nand U4652 (N_4652,N_2225,N_796);
and U4653 (N_4653,N_2410,N_193);
nor U4654 (N_4654,N_1145,N_2266);
and U4655 (N_4655,N_1939,N_894);
and U4656 (N_4656,N_1043,N_279);
nand U4657 (N_4657,N_1668,N_1847);
or U4658 (N_4658,N_612,N_2391);
and U4659 (N_4659,N_1003,N_1193);
and U4660 (N_4660,N_926,N_334);
nand U4661 (N_4661,N_1518,N_2460);
nand U4662 (N_4662,N_1871,N_826);
nor U4663 (N_4663,N_154,N_1875);
and U4664 (N_4664,N_2491,N_2480);
and U4665 (N_4665,N_2175,N_150);
or U4666 (N_4666,N_1939,N_2391);
xor U4667 (N_4667,N_1765,N_1919);
nor U4668 (N_4668,N_1142,N_1008);
and U4669 (N_4669,N_232,N_2396);
and U4670 (N_4670,N_207,N_47);
nand U4671 (N_4671,N_1974,N_960);
and U4672 (N_4672,N_481,N_1927);
and U4673 (N_4673,N_1736,N_1238);
nand U4674 (N_4674,N_1708,N_796);
and U4675 (N_4675,N_837,N_1975);
nor U4676 (N_4676,N_740,N_934);
and U4677 (N_4677,N_580,N_2005);
xnor U4678 (N_4678,N_589,N_1565);
nor U4679 (N_4679,N_1684,N_1121);
nand U4680 (N_4680,N_1891,N_2158);
and U4681 (N_4681,N_1349,N_290);
xnor U4682 (N_4682,N_165,N_1058);
or U4683 (N_4683,N_911,N_1214);
nor U4684 (N_4684,N_20,N_2445);
nand U4685 (N_4685,N_1672,N_714);
and U4686 (N_4686,N_306,N_394);
or U4687 (N_4687,N_2418,N_2329);
xnor U4688 (N_4688,N_1287,N_2065);
nor U4689 (N_4689,N_1617,N_1100);
and U4690 (N_4690,N_937,N_629);
nand U4691 (N_4691,N_2308,N_1002);
or U4692 (N_4692,N_451,N_1213);
or U4693 (N_4693,N_784,N_76);
xor U4694 (N_4694,N_1072,N_1517);
or U4695 (N_4695,N_2203,N_506);
or U4696 (N_4696,N_2402,N_1021);
or U4697 (N_4697,N_1079,N_1575);
xnor U4698 (N_4698,N_932,N_271);
nor U4699 (N_4699,N_1189,N_1437);
nand U4700 (N_4700,N_1016,N_267);
or U4701 (N_4701,N_554,N_477);
xor U4702 (N_4702,N_726,N_943);
and U4703 (N_4703,N_828,N_503);
nor U4704 (N_4704,N_2248,N_1315);
xnor U4705 (N_4705,N_1317,N_277);
or U4706 (N_4706,N_254,N_215);
nor U4707 (N_4707,N_902,N_1084);
or U4708 (N_4708,N_528,N_271);
nor U4709 (N_4709,N_1617,N_536);
and U4710 (N_4710,N_1458,N_2318);
nor U4711 (N_4711,N_91,N_253);
xnor U4712 (N_4712,N_890,N_159);
and U4713 (N_4713,N_1557,N_1512);
and U4714 (N_4714,N_1227,N_1067);
or U4715 (N_4715,N_2410,N_1234);
nand U4716 (N_4716,N_2453,N_996);
and U4717 (N_4717,N_882,N_1785);
nor U4718 (N_4718,N_849,N_138);
nand U4719 (N_4719,N_550,N_540);
and U4720 (N_4720,N_2322,N_2086);
and U4721 (N_4721,N_534,N_1713);
nor U4722 (N_4722,N_1308,N_304);
or U4723 (N_4723,N_1655,N_327);
nand U4724 (N_4724,N_355,N_273);
xnor U4725 (N_4725,N_1659,N_1260);
and U4726 (N_4726,N_1447,N_456);
nand U4727 (N_4727,N_2471,N_2392);
xor U4728 (N_4728,N_1227,N_2267);
and U4729 (N_4729,N_1588,N_456);
nor U4730 (N_4730,N_2396,N_380);
nand U4731 (N_4731,N_1274,N_353);
and U4732 (N_4732,N_1006,N_232);
nor U4733 (N_4733,N_2341,N_755);
and U4734 (N_4734,N_2207,N_1721);
or U4735 (N_4735,N_2431,N_1275);
xnor U4736 (N_4736,N_2111,N_164);
nor U4737 (N_4737,N_1073,N_523);
xnor U4738 (N_4738,N_856,N_231);
or U4739 (N_4739,N_2432,N_325);
nor U4740 (N_4740,N_2264,N_709);
or U4741 (N_4741,N_1781,N_147);
xnor U4742 (N_4742,N_1450,N_1169);
nand U4743 (N_4743,N_1041,N_2003);
nor U4744 (N_4744,N_2249,N_1955);
nor U4745 (N_4745,N_2405,N_1689);
and U4746 (N_4746,N_1143,N_2389);
nor U4747 (N_4747,N_823,N_1155);
and U4748 (N_4748,N_1012,N_783);
nor U4749 (N_4749,N_148,N_1243);
or U4750 (N_4750,N_526,N_1461);
or U4751 (N_4751,N_1924,N_1790);
or U4752 (N_4752,N_1490,N_371);
nand U4753 (N_4753,N_1450,N_1574);
nand U4754 (N_4754,N_1579,N_1389);
and U4755 (N_4755,N_2377,N_462);
nor U4756 (N_4756,N_331,N_444);
and U4757 (N_4757,N_512,N_1782);
or U4758 (N_4758,N_1408,N_892);
nand U4759 (N_4759,N_2111,N_1302);
or U4760 (N_4760,N_1011,N_2329);
nor U4761 (N_4761,N_2292,N_2059);
and U4762 (N_4762,N_145,N_586);
nor U4763 (N_4763,N_2184,N_1952);
xnor U4764 (N_4764,N_1801,N_2234);
and U4765 (N_4765,N_1990,N_1175);
and U4766 (N_4766,N_549,N_1002);
and U4767 (N_4767,N_229,N_1463);
xnor U4768 (N_4768,N_1313,N_652);
or U4769 (N_4769,N_2388,N_2079);
and U4770 (N_4770,N_1198,N_2034);
nor U4771 (N_4771,N_1593,N_1451);
and U4772 (N_4772,N_770,N_572);
nand U4773 (N_4773,N_1244,N_1775);
nand U4774 (N_4774,N_1130,N_1405);
and U4775 (N_4775,N_231,N_84);
and U4776 (N_4776,N_1245,N_1063);
xor U4777 (N_4777,N_384,N_160);
and U4778 (N_4778,N_1257,N_262);
nor U4779 (N_4779,N_1813,N_2067);
nand U4780 (N_4780,N_1286,N_2222);
xnor U4781 (N_4781,N_900,N_253);
nor U4782 (N_4782,N_1403,N_1369);
nor U4783 (N_4783,N_680,N_2330);
nand U4784 (N_4784,N_2140,N_1059);
nor U4785 (N_4785,N_1726,N_383);
nand U4786 (N_4786,N_990,N_1258);
and U4787 (N_4787,N_1874,N_909);
xnor U4788 (N_4788,N_2209,N_257);
or U4789 (N_4789,N_1024,N_1668);
nand U4790 (N_4790,N_2285,N_1024);
nand U4791 (N_4791,N_2017,N_402);
nand U4792 (N_4792,N_676,N_2135);
or U4793 (N_4793,N_778,N_8);
nand U4794 (N_4794,N_1441,N_1365);
or U4795 (N_4795,N_138,N_1285);
and U4796 (N_4796,N_395,N_1681);
nand U4797 (N_4797,N_295,N_17);
nor U4798 (N_4798,N_1463,N_811);
or U4799 (N_4799,N_126,N_304);
xnor U4800 (N_4800,N_971,N_1544);
or U4801 (N_4801,N_488,N_387);
nand U4802 (N_4802,N_617,N_409);
and U4803 (N_4803,N_915,N_689);
nand U4804 (N_4804,N_1358,N_1285);
and U4805 (N_4805,N_1806,N_1350);
xnor U4806 (N_4806,N_1238,N_1737);
or U4807 (N_4807,N_1516,N_44);
xor U4808 (N_4808,N_2130,N_932);
nor U4809 (N_4809,N_893,N_931);
nor U4810 (N_4810,N_157,N_1918);
or U4811 (N_4811,N_656,N_612);
xor U4812 (N_4812,N_2205,N_1785);
and U4813 (N_4813,N_1971,N_892);
or U4814 (N_4814,N_2236,N_1878);
nor U4815 (N_4815,N_2209,N_1841);
or U4816 (N_4816,N_1215,N_1517);
or U4817 (N_4817,N_2151,N_1901);
xor U4818 (N_4818,N_2058,N_239);
nor U4819 (N_4819,N_1378,N_632);
xor U4820 (N_4820,N_242,N_1569);
and U4821 (N_4821,N_2405,N_1383);
or U4822 (N_4822,N_1893,N_709);
or U4823 (N_4823,N_1084,N_1710);
xor U4824 (N_4824,N_553,N_1557);
and U4825 (N_4825,N_174,N_338);
and U4826 (N_4826,N_1722,N_1526);
nor U4827 (N_4827,N_2467,N_1004);
nand U4828 (N_4828,N_1583,N_1656);
or U4829 (N_4829,N_1228,N_792);
or U4830 (N_4830,N_2409,N_1587);
nor U4831 (N_4831,N_809,N_2000);
nand U4832 (N_4832,N_611,N_1412);
nor U4833 (N_4833,N_113,N_960);
nand U4834 (N_4834,N_9,N_685);
nor U4835 (N_4835,N_1589,N_2160);
nor U4836 (N_4836,N_1248,N_2258);
nor U4837 (N_4837,N_1026,N_1943);
xor U4838 (N_4838,N_92,N_294);
nor U4839 (N_4839,N_1623,N_446);
or U4840 (N_4840,N_1795,N_237);
nand U4841 (N_4841,N_1840,N_1586);
nor U4842 (N_4842,N_1482,N_1144);
xor U4843 (N_4843,N_239,N_534);
or U4844 (N_4844,N_311,N_1764);
and U4845 (N_4845,N_1276,N_1801);
xnor U4846 (N_4846,N_570,N_2042);
nand U4847 (N_4847,N_2408,N_1827);
or U4848 (N_4848,N_1867,N_1329);
or U4849 (N_4849,N_2225,N_943);
xnor U4850 (N_4850,N_1412,N_1027);
nor U4851 (N_4851,N_63,N_1136);
nor U4852 (N_4852,N_156,N_1952);
and U4853 (N_4853,N_2185,N_1235);
xor U4854 (N_4854,N_761,N_1588);
or U4855 (N_4855,N_753,N_1201);
nor U4856 (N_4856,N_1959,N_238);
and U4857 (N_4857,N_913,N_1580);
or U4858 (N_4858,N_1454,N_576);
xor U4859 (N_4859,N_1905,N_402);
nor U4860 (N_4860,N_2292,N_343);
or U4861 (N_4861,N_132,N_1092);
xor U4862 (N_4862,N_913,N_387);
nor U4863 (N_4863,N_2153,N_2322);
nor U4864 (N_4864,N_1976,N_1086);
and U4865 (N_4865,N_1074,N_1513);
nand U4866 (N_4866,N_237,N_763);
nand U4867 (N_4867,N_1091,N_697);
nor U4868 (N_4868,N_828,N_2006);
nor U4869 (N_4869,N_2305,N_42);
nand U4870 (N_4870,N_2194,N_2440);
nor U4871 (N_4871,N_1801,N_158);
or U4872 (N_4872,N_70,N_420);
xnor U4873 (N_4873,N_2053,N_513);
nand U4874 (N_4874,N_1591,N_12);
xnor U4875 (N_4875,N_719,N_1961);
xnor U4876 (N_4876,N_350,N_529);
nor U4877 (N_4877,N_1601,N_1904);
nand U4878 (N_4878,N_2251,N_2319);
or U4879 (N_4879,N_1590,N_887);
nor U4880 (N_4880,N_1750,N_1878);
nor U4881 (N_4881,N_1437,N_2155);
or U4882 (N_4882,N_54,N_2082);
xor U4883 (N_4883,N_2299,N_1084);
nor U4884 (N_4884,N_42,N_588);
or U4885 (N_4885,N_283,N_525);
nor U4886 (N_4886,N_591,N_1241);
nand U4887 (N_4887,N_2059,N_1799);
nor U4888 (N_4888,N_217,N_686);
nor U4889 (N_4889,N_692,N_735);
and U4890 (N_4890,N_2244,N_1289);
and U4891 (N_4891,N_1053,N_2496);
and U4892 (N_4892,N_465,N_112);
and U4893 (N_4893,N_687,N_1354);
or U4894 (N_4894,N_926,N_2242);
xnor U4895 (N_4895,N_543,N_1753);
nand U4896 (N_4896,N_624,N_321);
or U4897 (N_4897,N_1689,N_2383);
xnor U4898 (N_4898,N_377,N_177);
and U4899 (N_4899,N_717,N_2136);
nor U4900 (N_4900,N_1339,N_536);
and U4901 (N_4901,N_456,N_2474);
xnor U4902 (N_4902,N_1161,N_383);
and U4903 (N_4903,N_2494,N_1115);
or U4904 (N_4904,N_1918,N_1788);
nand U4905 (N_4905,N_194,N_707);
and U4906 (N_4906,N_1500,N_2467);
or U4907 (N_4907,N_2338,N_1942);
nor U4908 (N_4908,N_105,N_2214);
nor U4909 (N_4909,N_1954,N_1753);
xnor U4910 (N_4910,N_532,N_1152);
or U4911 (N_4911,N_158,N_386);
or U4912 (N_4912,N_2478,N_1699);
xor U4913 (N_4913,N_2337,N_1055);
nand U4914 (N_4914,N_2205,N_1868);
and U4915 (N_4915,N_960,N_1037);
xor U4916 (N_4916,N_1350,N_1579);
and U4917 (N_4917,N_1924,N_658);
nor U4918 (N_4918,N_1190,N_2062);
and U4919 (N_4919,N_285,N_974);
nor U4920 (N_4920,N_2386,N_51);
nand U4921 (N_4921,N_928,N_1619);
nor U4922 (N_4922,N_2037,N_671);
nor U4923 (N_4923,N_1332,N_2402);
or U4924 (N_4924,N_1237,N_1212);
nand U4925 (N_4925,N_1332,N_1414);
xor U4926 (N_4926,N_558,N_894);
xnor U4927 (N_4927,N_248,N_1446);
or U4928 (N_4928,N_250,N_1441);
or U4929 (N_4929,N_2205,N_919);
xor U4930 (N_4930,N_191,N_2112);
xor U4931 (N_4931,N_414,N_1733);
nor U4932 (N_4932,N_915,N_810);
or U4933 (N_4933,N_1836,N_1223);
nand U4934 (N_4934,N_556,N_721);
and U4935 (N_4935,N_693,N_1707);
and U4936 (N_4936,N_2170,N_1337);
or U4937 (N_4937,N_1351,N_268);
nand U4938 (N_4938,N_1510,N_2202);
and U4939 (N_4939,N_1375,N_1940);
nor U4940 (N_4940,N_2000,N_642);
or U4941 (N_4941,N_1250,N_644);
nor U4942 (N_4942,N_1100,N_915);
nand U4943 (N_4943,N_1550,N_875);
xnor U4944 (N_4944,N_435,N_72);
or U4945 (N_4945,N_809,N_1755);
and U4946 (N_4946,N_1974,N_986);
or U4947 (N_4947,N_1931,N_582);
and U4948 (N_4948,N_2383,N_361);
or U4949 (N_4949,N_2117,N_2279);
nand U4950 (N_4950,N_215,N_2153);
nor U4951 (N_4951,N_2450,N_739);
nand U4952 (N_4952,N_1840,N_959);
or U4953 (N_4953,N_1293,N_1413);
nor U4954 (N_4954,N_352,N_1876);
and U4955 (N_4955,N_655,N_2041);
nand U4956 (N_4956,N_279,N_602);
nand U4957 (N_4957,N_283,N_983);
xor U4958 (N_4958,N_597,N_1662);
nor U4959 (N_4959,N_1951,N_1172);
or U4960 (N_4960,N_1713,N_1944);
and U4961 (N_4961,N_1353,N_1970);
nand U4962 (N_4962,N_446,N_48);
nor U4963 (N_4963,N_1640,N_1258);
nor U4964 (N_4964,N_2099,N_1467);
and U4965 (N_4965,N_1086,N_2457);
or U4966 (N_4966,N_304,N_1148);
or U4967 (N_4967,N_1126,N_1938);
nand U4968 (N_4968,N_28,N_223);
and U4969 (N_4969,N_281,N_1518);
xnor U4970 (N_4970,N_2370,N_2135);
nand U4971 (N_4971,N_434,N_2140);
and U4972 (N_4972,N_933,N_1303);
or U4973 (N_4973,N_211,N_1330);
xnor U4974 (N_4974,N_816,N_1439);
nor U4975 (N_4975,N_1708,N_2304);
xnor U4976 (N_4976,N_29,N_2469);
or U4977 (N_4977,N_1399,N_702);
xor U4978 (N_4978,N_1251,N_1469);
xnor U4979 (N_4979,N_69,N_2439);
nand U4980 (N_4980,N_2241,N_198);
nor U4981 (N_4981,N_1970,N_2041);
and U4982 (N_4982,N_327,N_611);
nor U4983 (N_4983,N_898,N_2280);
nor U4984 (N_4984,N_1687,N_482);
and U4985 (N_4985,N_68,N_1386);
xnor U4986 (N_4986,N_2377,N_1661);
and U4987 (N_4987,N_1086,N_1389);
nor U4988 (N_4988,N_157,N_731);
nor U4989 (N_4989,N_1388,N_2389);
and U4990 (N_4990,N_512,N_434);
or U4991 (N_4991,N_2274,N_1391);
xor U4992 (N_4992,N_1663,N_2173);
or U4993 (N_4993,N_2408,N_26);
and U4994 (N_4994,N_666,N_1463);
nor U4995 (N_4995,N_154,N_2491);
nor U4996 (N_4996,N_76,N_2044);
or U4997 (N_4997,N_643,N_2182);
nand U4998 (N_4998,N_2279,N_1647);
or U4999 (N_4999,N_1689,N_1958);
or U5000 (N_5000,N_4922,N_3079);
and U5001 (N_5001,N_4272,N_4335);
nor U5002 (N_5002,N_2708,N_3509);
nor U5003 (N_5003,N_4844,N_3755);
nand U5004 (N_5004,N_3727,N_4976);
xnor U5005 (N_5005,N_4533,N_3174);
nor U5006 (N_5006,N_3578,N_3183);
or U5007 (N_5007,N_3542,N_4802);
or U5008 (N_5008,N_2907,N_3897);
nor U5009 (N_5009,N_4153,N_4390);
xor U5010 (N_5010,N_4917,N_2727);
and U5011 (N_5011,N_3023,N_4187);
nand U5012 (N_5012,N_4310,N_3389);
xor U5013 (N_5013,N_3355,N_2950);
nand U5014 (N_5014,N_4329,N_3964);
nand U5015 (N_5015,N_4300,N_4258);
nor U5016 (N_5016,N_3979,N_3346);
nand U5017 (N_5017,N_3744,N_2803);
xor U5018 (N_5018,N_2955,N_4018);
xor U5019 (N_5019,N_4352,N_2751);
or U5020 (N_5020,N_3416,N_4124);
nand U5021 (N_5021,N_3114,N_4560);
or U5022 (N_5022,N_3135,N_2783);
nand U5023 (N_5023,N_4102,N_2561);
nor U5024 (N_5024,N_4375,N_4453);
nand U5025 (N_5025,N_4945,N_4376);
xnor U5026 (N_5026,N_3675,N_3638);
nor U5027 (N_5027,N_4367,N_3238);
nor U5028 (N_5028,N_4441,N_2583);
xor U5029 (N_5029,N_4177,N_3863);
xor U5030 (N_5030,N_2892,N_3670);
or U5031 (N_5031,N_4563,N_3586);
or U5032 (N_5032,N_4497,N_4440);
and U5033 (N_5033,N_4055,N_2973);
nand U5034 (N_5034,N_4767,N_4629);
and U5035 (N_5035,N_4506,N_2603);
or U5036 (N_5036,N_2776,N_4206);
xnor U5037 (N_5037,N_3100,N_3039);
nor U5038 (N_5038,N_4630,N_4674);
xor U5039 (N_5039,N_3793,N_3987);
or U5040 (N_5040,N_3071,N_4907);
and U5041 (N_5041,N_3400,N_2936);
nand U5042 (N_5042,N_4387,N_3886);
nor U5043 (N_5043,N_3181,N_2592);
nor U5044 (N_5044,N_2879,N_2582);
nor U5045 (N_5045,N_4848,N_3657);
and U5046 (N_5046,N_3662,N_3557);
and U5047 (N_5047,N_3480,N_2997);
or U5048 (N_5048,N_3568,N_3095);
and U5049 (N_5049,N_4290,N_3397);
nand U5050 (N_5050,N_3093,N_3648);
nor U5051 (N_5051,N_3421,N_4688);
nand U5052 (N_5052,N_3026,N_4150);
or U5053 (N_5053,N_3276,N_2653);
nor U5054 (N_5054,N_2543,N_3001);
or U5055 (N_5055,N_3823,N_2576);
nor U5056 (N_5056,N_4807,N_4333);
and U5057 (N_5057,N_4668,N_4762);
nand U5058 (N_5058,N_3575,N_3185);
or U5059 (N_5059,N_4831,N_4406);
xor U5060 (N_5060,N_3535,N_4701);
and U5061 (N_5061,N_4599,N_3459);
xor U5062 (N_5062,N_3685,N_4667);
and U5063 (N_5063,N_4295,N_3365);
nor U5064 (N_5064,N_4189,N_4442);
nand U5065 (N_5065,N_3443,N_4416);
or U5066 (N_5066,N_2787,N_4895);
or U5067 (N_5067,N_4654,N_2584);
or U5068 (N_5068,N_3497,N_4556);
or U5069 (N_5069,N_2714,N_4618);
or U5070 (N_5070,N_3106,N_4501);
xnor U5071 (N_5071,N_2709,N_4585);
xor U5072 (N_5072,N_2522,N_3414);
or U5073 (N_5073,N_4852,N_2745);
and U5074 (N_5074,N_3850,N_2699);
and U5075 (N_5075,N_3187,N_3462);
nand U5076 (N_5076,N_2986,N_2840);
nor U5077 (N_5077,N_2573,N_2967);
nand U5078 (N_5078,N_4853,N_3013);
nor U5079 (N_5079,N_3028,N_4723);
or U5080 (N_5080,N_2963,N_4357);
xor U5081 (N_5081,N_4545,N_4972);
nor U5082 (N_5082,N_3390,N_3167);
nand U5083 (N_5083,N_3044,N_4386);
or U5084 (N_5084,N_4578,N_3628);
nand U5085 (N_5085,N_4829,N_4604);
xnor U5086 (N_5086,N_4444,N_3605);
or U5087 (N_5087,N_4038,N_2526);
and U5088 (N_5088,N_3452,N_3773);
xor U5089 (N_5089,N_4252,N_4663);
xor U5090 (N_5090,N_3604,N_4135);
nor U5091 (N_5091,N_2876,N_4263);
and U5092 (N_5092,N_2652,N_3884);
and U5093 (N_5093,N_3231,N_4336);
nor U5094 (N_5094,N_3917,N_4472);
nand U5095 (N_5095,N_4240,N_3048);
and U5096 (N_5096,N_4257,N_4374);
or U5097 (N_5097,N_2619,N_4897);
xnor U5098 (N_5098,N_3171,N_3073);
xor U5099 (N_5099,N_4815,N_3213);
xnor U5100 (N_5100,N_4571,N_4638);
nand U5101 (N_5101,N_4940,N_3265);
nand U5102 (N_5102,N_3169,N_4321);
and U5103 (N_5103,N_3247,N_4283);
xnor U5104 (N_5104,N_2921,N_2773);
and U5105 (N_5105,N_4391,N_2664);
or U5106 (N_5106,N_4693,N_2985);
nor U5107 (N_5107,N_4017,N_4096);
nand U5108 (N_5108,N_4180,N_2648);
and U5109 (N_5109,N_2974,N_4652);
nor U5110 (N_5110,N_3970,N_4185);
or U5111 (N_5111,N_3872,N_3740);
xnor U5112 (N_5112,N_4176,N_4388);
or U5113 (N_5113,N_2774,N_3022);
nor U5114 (N_5114,N_3817,N_2646);
nor U5115 (N_5115,N_2737,N_3669);
and U5116 (N_5116,N_4330,N_2639);
nand U5117 (N_5117,N_4265,N_4095);
or U5118 (N_5118,N_4608,N_2855);
nor U5119 (N_5119,N_2697,N_4963);
nand U5120 (N_5120,N_4896,N_3179);
nand U5121 (N_5121,N_3325,N_2909);
or U5122 (N_5122,N_3816,N_3258);
or U5123 (N_5123,N_2743,N_2746);
or U5124 (N_5124,N_4858,N_2707);
nor U5125 (N_5125,N_3966,N_4380);
or U5126 (N_5126,N_3042,N_3960);
xor U5127 (N_5127,N_4314,N_4211);
or U5128 (N_5128,N_4537,N_3889);
or U5129 (N_5129,N_3453,N_2856);
and U5130 (N_5130,N_4019,N_4130);
or U5131 (N_5131,N_4328,N_3328);
and U5132 (N_5132,N_4094,N_3519);
or U5133 (N_5133,N_2849,N_3805);
nand U5134 (N_5134,N_2845,N_4229);
or U5135 (N_5135,N_3874,N_4399);
or U5136 (N_5136,N_2654,N_4226);
nor U5137 (N_5137,N_3650,N_4946);
xor U5138 (N_5138,N_4460,N_4152);
nand U5139 (N_5139,N_2738,N_3762);
xnor U5140 (N_5140,N_4422,N_2869);
nand U5141 (N_5141,N_4043,N_3445);
nor U5142 (N_5142,N_4297,N_4659);
and U5143 (N_5143,N_4632,N_3614);
nand U5144 (N_5144,N_2949,N_4254);
or U5145 (N_5145,N_2863,N_3832);
xor U5146 (N_5146,N_2797,N_4686);
or U5147 (N_5147,N_2719,N_3422);
nand U5148 (N_5148,N_3373,N_3712);
nor U5149 (N_5149,N_3704,N_3565);
nand U5150 (N_5150,N_3348,N_4999);
xor U5151 (N_5151,N_4984,N_2594);
nor U5152 (N_5152,N_2586,N_4170);
or U5153 (N_5153,N_3184,N_3948);
nand U5154 (N_5154,N_4623,N_4093);
xnor U5155 (N_5155,N_2811,N_4732);
nor U5156 (N_5156,N_2994,N_3892);
nand U5157 (N_5157,N_4100,N_3045);
nor U5158 (N_5158,N_3413,N_3386);
or U5159 (N_5159,N_3533,N_3461);
xor U5160 (N_5160,N_3838,N_4727);
and U5161 (N_5161,N_4118,N_3054);
xnor U5162 (N_5162,N_3955,N_2591);
nor U5163 (N_5163,N_2796,N_4910);
nor U5164 (N_5164,N_4395,N_4591);
and U5165 (N_5165,N_3959,N_2813);
xor U5166 (N_5166,N_3715,N_4166);
xor U5167 (N_5167,N_4784,N_3802);
or U5168 (N_5168,N_2739,N_4344);
xor U5169 (N_5169,N_3020,N_4107);
or U5170 (N_5170,N_2640,N_4134);
nor U5171 (N_5171,N_3418,N_2650);
nor U5172 (N_5172,N_4861,N_4332);
and U5173 (N_5173,N_3853,N_2502);
nand U5174 (N_5174,N_3983,N_2509);
nand U5175 (N_5175,N_3063,N_4378);
nand U5176 (N_5176,N_4296,N_4868);
and U5177 (N_5177,N_4553,N_4811);
xnor U5178 (N_5178,N_3719,N_4132);
nand U5179 (N_5179,N_3686,N_4671);
nor U5180 (N_5180,N_3561,N_3653);
or U5181 (N_5181,N_2911,N_3393);
nand U5182 (N_5182,N_3363,N_3009);
xor U5183 (N_5183,N_4916,N_4740);
xnor U5184 (N_5184,N_3556,N_2926);
xnor U5185 (N_5185,N_3278,N_2960);
or U5186 (N_5186,N_3340,N_4745);
and U5187 (N_5187,N_3015,N_4901);
or U5188 (N_5188,N_3043,N_4496);
and U5189 (N_5189,N_2988,N_2516);
nor U5190 (N_5190,N_4982,N_2844);
nor U5191 (N_5191,N_2978,N_4201);
xnor U5192 (N_5192,N_4890,N_4370);
nor U5193 (N_5193,N_4912,N_3763);
nor U5194 (N_5194,N_2725,N_4011);
xor U5195 (N_5195,N_4866,N_4438);
or U5196 (N_5196,N_3087,N_4738);
nand U5197 (N_5197,N_4766,N_4580);
and U5198 (N_5198,N_3350,N_3683);
or U5199 (N_5199,N_3776,N_3842);
nor U5200 (N_5200,N_2989,N_3963);
nand U5201 (N_5201,N_3006,N_3695);
nor U5202 (N_5202,N_3759,N_3896);
nand U5203 (N_5203,N_3941,N_3211);
or U5204 (N_5204,N_4068,N_3320);
and U5205 (N_5205,N_4758,N_3778);
xnor U5206 (N_5206,N_4457,N_3444);
or U5207 (N_5207,N_4516,N_4271);
and U5208 (N_5208,N_2841,N_3146);
and U5209 (N_5209,N_4584,N_4565);
xnor U5210 (N_5210,N_3011,N_4157);
and U5211 (N_5211,N_3293,N_4562);
nand U5212 (N_5212,N_4683,N_4318);
and U5213 (N_5213,N_4347,N_3168);
and U5214 (N_5214,N_4168,N_3699);
xor U5215 (N_5215,N_3016,N_3587);
nor U5216 (N_5216,N_3124,N_3267);
nor U5217 (N_5217,N_3730,N_4803);
nor U5218 (N_5218,N_3195,N_3434);
or U5219 (N_5219,N_3190,N_4892);
nand U5220 (N_5220,N_2517,N_2626);
nand U5221 (N_5221,N_4208,N_3339);
or U5222 (N_5222,N_4951,N_3229);
nand U5223 (N_5223,N_2805,N_3243);
nand U5224 (N_5224,N_3076,N_2730);
xnor U5225 (N_5225,N_2927,N_4010);
xor U5226 (N_5226,N_4718,N_3814);
or U5227 (N_5227,N_3905,N_3924);
and U5228 (N_5228,N_4641,N_3357);
and U5229 (N_5229,N_3919,N_4225);
and U5230 (N_5230,N_3160,N_2683);
nand U5231 (N_5231,N_4586,N_4827);
nand U5232 (N_5232,N_3067,N_4891);
nand U5233 (N_5233,N_4382,N_4221);
or U5234 (N_5234,N_3411,N_4733);
and U5235 (N_5235,N_4883,N_4510);
xor U5236 (N_5236,N_3554,N_4266);
nor U5237 (N_5237,N_4074,N_3965);
nor U5238 (N_5238,N_3780,N_4519);
xor U5239 (N_5239,N_3090,N_4230);
nor U5240 (N_5240,N_3148,N_4601);
xnor U5241 (N_5241,N_3482,N_4577);
and U5242 (N_5242,N_2874,N_3511);
xnor U5243 (N_5243,N_2958,N_4707);
nand U5244 (N_5244,N_3246,N_3860);
and U5245 (N_5245,N_3861,N_3698);
and U5246 (N_5246,N_3985,N_3396);
nor U5247 (N_5247,N_3403,N_2951);
and U5248 (N_5248,N_3037,N_4103);
nor U5249 (N_5249,N_3967,N_2547);
nor U5250 (N_5250,N_2513,N_3399);
and U5251 (N_5251,N_3579,N_3731);
nor U5252 (N_5252,N_4466,N_3585);
nor U5253 (N_5253,N_4870,N_3143);
xor U5254 (N_5254,N_4353,N_4133);
nand U5255 (N_5255,N_3507,N_3757);
or U5256 (N_5256,N_4637,N_3997);
or U5257 (N_5257,N_3379,N_3427);
nor U5258 (N_5258,N_4694,N_4590);
or U5259 (N_5259,N_4280,N_4249);
and U5260 (N_5260,N_3716,N_4840);
xor U5261 (N_5261,N_4343,N_4817);
nand U5262 (N_5262,N_4863,N_3374);
xor U5263 (N_5263,N_2858,N_2784);
xor U5264 (N_5264,N_4731,N_4572);
nor U5265 (N_5265,N_3040,N_4938);
and U5266 (N_5266,N_3818,N_3127);
or U5267 (N_5267,N_4199,N_3259);
or U5268 (N_5268,N_3703,N_3865);
and U5269 (N_5269,N_2802,N_4925);
or U5270 (N_5270,N_3834,N_2638);
and U5271 (N_5271,N_4739,N_3203);
and U5272 (N_5272,N_4903,N_4785);
or U5273 (N_5273,N_3671,N_3639);
nor U5274 (N_5274,N_2546,N_2940);
nor U5275 (N_5275,N_4035,N_3352);
nand U5276 (N_5276,N_3464,N_4575);
nor U5277 (N_5277,N_2672,N_4499);
and U5278 (N_5278,N_4777,N_3223);
xor U5279 (N_5279,N_2530,N_3696);
or U5280 (N_5280,N_4816,N_4613);
and U5281 (N_5281,N_3601,N_4763);
xnor U5282 (N_5282,N_4119,N_3728);
and U5283 (N_5283,N_2663,N_3285);
xor U5284 (N_5284,N_3908,N_4616);
and U5285 (N_5285,N_4915,N_3209);
xnor U5286 (N_5286,N_4692,N_3878);
xor U5287 (N_5287,N_4906,N_2669);
or U5288 (N_5288,N_4626,N_4062);
xnor U5289 (N_5289,N_2612,N_4040);
nor U5290 (N_5290,N_4875,N_3977);
nand U5291 (N_5291,N_4856,N_3361);
nor U5292 (N_5292,N_2637,N_2541);
nor U5293 (N_5293,N_2756,N_3094);
and U5294 (N_5294,N_3688,N_3341);
nor U5295 (N_5295,N_2902,N_3824);
nor U5296 (N_5296,N_4242,N_2815);
nor U5297 (N_5297,N_2624,N_2843);
or U5298 (N_5298,N_3454,N_2712);
nor U5299 (N_5299,N_4358,N_3074);
and U5300 (N_5300,N_3201,N_4712);
and U5301 (N_5301,N_4372,N_3262);
and U5302 (N_5302,N_2760,N_3121);
nand U5303 (N_5303,N_4639,N_4955);
xor U5304 (N_5304,N_2528,N_4800);
xnor U5305 (N_5305,N_3132,N_4798);
xor U5306 (N_5306,N_4022,N_3736);
xor U5307 (N_5307,N_3440,N_3649);
nor U5308 (N_5308,N_3836,N_2539);
and U5309 (N_5309,N_4914,N_3271);
nand U5310 (N_5310,N_4411,N_2941);
xor U5311 (N_5311,N_3110,N_4569);
xnor U5312 (N_5312,N_4085,N_3576);
or U5313 (N_5313,N_2647,N_4685);
nor U5314 (N_5314,N_3909,N_4425);
nand U5315 (N_5315,N_3911,N_3072);
or U5316 (N_5316,N_4106,N_2822);
or U5317 (N_5317,N_2992,N_3947);
nor U5318 (N_5318,N_3172,N_4774);
xor U5319 (N_5319,N_4512,N_3492);
xor U5320 (N_5320,N_3684,N_2548);
xnor U5321 (N_5321,N_3077,N_4084);
and U5322 (N_5322,N_2896,N_4407);
nor U5323 (N_5323,N_2560,N_4541);
or U5324 (N_5324,N_3316,N_3176);
or U5325 (N_5325,N_4480,N_3976);
or U5326 (N_5326,N_3133,N_3558);
and U5327 (N_5327,N_4307,N_4024);
nor U5328 (N_5328,N_2752,N_3939);
and U5329 (N_5329,N_3550,N_3574);
nand U5330 (N_5330,N_4385,N_4636);
nor U5331 (N_5331,N_4463,N_3517);
nand U5332 (N_5332,N_2740,N_3518);
nand U5333 (N_5333,N_3237,N_3333);
nor U5334 (N_5334,N_4924,N_4072);
and U5335 (N_5335,N_2588,N_2657);
or U5336 (N_5336,N_3120,N_4764);
or U5337 (N_5337,N_4465,N_4953);
nand U5338 (N_5338,N_3922,N_2680);
and U5339 (N_5339,N_4851,N_4186);
nand U5340 (N_5340,N_2733,N_4360);
nand U5341 (N_5341,N_2608,N_4483);
nand U5342 (N_5342,N_4319,N_3600);
nand U5343 (N_5343,N_3555,N_4564);
xor U5344 (N_5344,N_4698,N_4841);
nand U5345 (N_5345,N_3282,N_4361);
or U5346 (N_5346,N_3395,N_3809);
and U5347 (N_5347,N_3487,N_4053);
nand U5348 (N_5348,N_4820,N_4989);
and U5349 (N_5349,N_4339,N_4830);
and U5350 (N_5350,N_3900,N_4779);
xor U5351 (N_5351,N_2801,N_3291);
nor U5352 (N_5352,N_4156,N_3980);
xor U5353 (N_5353,N_4042,N_3046);
and U5354 (N_5354,N_3774,N_3761);
xor U5355 (N_5355,N_4056,N_4631);
xnor U5356 (N_5356,N_2627,N_3324);
and U5357 (N_5357,N_3890,N_3580);
and U5358 (N_5358,N_3916,N_4760);
nand U5359 (N_5359,N_3368,N_2939);
and U5360 (N_5360,N_3978,N_3142);
and U5361 (N_5361,N_2836,N_3687);
or U5362 (N_5362,N_3233,N_4143);
or U5363 (N_5363,N_3115,N_3391);
or U5364 (N_5364,N_4838,N_4052);
xnor U5365 (N_5365,N_4801,N_3711);
nor U5366 (N_5366,N_4127,N_4509);
xor U5367 (N_5367,N_4768,N_4369);
or U5368 (N_5368,N_3618,N_3051);
or U5369 (N_5369,N_4928,N_4462);
or U5370 (N_5370,N_3249,N_4467);
xnor U5371 (N_5371,N_3113,N_3111);
and U5372 (N_5372,N_2620,N_4744);
nor U5373 (N_5373,N_4125,N_4859);
or U5374 (N_5374,N_3283,N_4617);
and U5375 (N_5375,N_2574,N_2764);
or U5376 (N_5376,N_3002,N_3027);
nor U5377 (N_5377,N_4862,N_2629);
and U5378 (N_5378,N_3625,N_4413);
and U5379 (N_5379,N_4341,N_3681);
and U5380 (N_5380,N_4684,N_3754);
xor U5381 (N_5381,N_4948,N_4909);
or U5382 (N_5382,N_2670,N_3538);
and U5383 (N_5383,N_4044,N_4126);
nand U5384 (N_5384,N_3629,N_2713);
xnor U5385 (N_5385,N_4155,N_2829);
nand U5386 (N_5386,N_3738,N_4567);
and U5387 (N_5387,N_4342,N_4262);
or U5388 (N_5388,N_2922,N_3645);
xnor U5389 (N_5389,N_3973,N_3366);
xnor U5390 (N_5390,N_4202,N_4819);
nor U5391 (N_5391,N_4792,N_4719);
xnor U5392 (N_5392,N_3024,N_4154);
or U5393 (N_5393,N_2690,N_3470);
and U5394 (N_5394,N_3795,N_4904);
xnor U5395 (N_5395,N_3118,N_3792);
nand U5396 (N_5396,N_3182,N_3253);
nor U5397 (N_5397,N_4525,N_4931);
and U5398 (N_5398,N_3624,N_2865);
xnor U5399 (N_5399,N_4101,N_2930);
or U5400 (N_5400,N_2847,N_2642);
or U5401 (N_5401,N_2655,N_4192);
and U5402 (N_5402,N_4006,N_4089);
nand U5403 (N_5403,N_4888,N_4935);
xor U5404 (N_5404,N_3526,N_4709);
xor U5405 (N_5405,N_2795,N_3989);
nand U5406 (N_5406,N_2970,N_3749);
or U5407 (N_5407,N_4471,N_4818);
and U5408 (N_5408,N_3354,N_2755);
or U5409 (N_5409,N_4970,N_3619);
or U5410 (N_5410,N_4179,N_4047);
nor U5411 (N_5411,N_3796,N_3310);
or U5412 (N_5412,N_3513,N_2693);
xnor U5413 (N_5413,N_4394,N_3982);
or U5414 (N_5414,N_4429,N_3177);
or U5415 (N_5415,N_3129,N_3877);
and U5416 (N_5416,N_3534,N_3153);
nor U5417 (N_5417,N_3777,N_4493);
and U5418 (N_5418,N_3713,N_3827);
nor U5419 (N_5419,N_4786,N_4447);
xor U5420 (N_5420,N_3460,N_4515);
nand U5421 (N_5421,N_2854,N_3197);
nand U5422 (N_5422,N_3990,N_3705);
or U5423 (N_5423,N_3718,N_3577);
and U5424 (N_5424,N_4839,N_3327);
or U5425 (N_5425,N_4433,N_3166);
xor U5426 (N_5426,N_2809,N_3260);
and U5427 (N_5427,N_3737,N_3745);
nor U5428 (N_5428,N_2682,N_4345);
or U5429 (N_5429,N_3199,N_4288);
nor U5430 (N_5430,N_2885,N_3306);
and U5431 (N_5431,N_2534,N_4600);
and U5432 (N_5432,N_3216,N_3164);
or U5433 (N_5433,N_4822,N_3566);
and U5434 (N_5434,N_3017,N_4751);
and U5435 (N_5435,N_4129,N_3104);
xnor U5436 (N_5436,N_3173,N_3584);
xnor U5437 (N_5437,N_2782,N_2991);
nand U5438 (N_5438,N_2744,N_3154);
nand U5439 (N_5439,N_3848,N_2726);
nand U5440 (N_5440,N_2761,N_4197);
nor U5441 (N_5441,N_4427,N_4322);
and U5442 (N_5442,N_4614,N_2819);
nand U5443 (N_5443,N_4079,N_2980);
or U5444 (N_5444,N_3784,N_4003);
nor U5445 (N_5445,N_3899,N_3206);
xor U5446 (N_5446,N_3995,N_4536);
nand U5447 (N_5447,N_2665,N_3170);
or U5448 (N_5448,N_3822,N_4728);
and U5449 (N_5449,N_2750,N_4775);
xor U5450 (N_5450,N_4486,N_4523);
or U5451 (N_5451,N_4412,N_3733);
or U5452 (N_5452,N_3342,N_3956);
xnor U5453 (N_5453,N_3131,N_3607);
nand U5454 (N_5454,N_3813,N_3483);
and U5455 (N_5455,N_3700,N_3934);
nand U5456 (N_5456,N_2536,N_4529);
nand U5457 (N_5457,N_3771,N_4535);
xor U5458 (N_5458,N_4885,N_3918);
xor U5459 (N_5459,N_3564,N_3858);
xnor U5460 (N_5460,N_4611,N_4821);
nand U5461 (N_5461,N_4736,N_4691);
and U5462 (N_5462,N_3597,N_2685);
and U5463 (N_5463,N_4649,N_3972);
nand U5464 (N_5464,N_3062,N_4459);
or U5465 (N_5465,N_4071,N_3943);
or U5466 (N_5466,N_3510,N_4243);
nand U5467 (N_5467,N_3791,N_3192);
nand U5468 (N_5468,N_4308,N_3268);
nor U5469 (N_5469,N_4828,N_4007);
nand U5470 (N_5470,N_3799,N_3904);
and U5471 (N_5471,N_3130,N_4312);
xnor U5472 (N_5472,N_4204,N_2520);
and U5473 (N_5473,N_2570,N_2861);
and U5474 (N_5474,N_3123,N_3086);
nor U5475 (N_5475,N_4514,N_4772);
or U5476 (N_5476,N_2731,N_4362);
nor U5477 (N_5477,N_3212,N_4434);
nor U5478 (N_5478,N_4110,N_2736);
nor U5479 (N_5479,N_4405,N_4610);
xor U5480 (N_5480,N_3204,N_2552);
nor U5481 (N_5481,N_3857,N_3360);
or U5482 (N_5482,N_3021,N_4175);
and U5483 (N_5483,N_4730,N_2928);
and U5484 (N_5484,N_4696,N_4404);
nand U5485 (N_5485,N_3770,N_2812);
nor U5486 (N_5486,N_2614,N_4958);
xor U5487 (N_5487,N_2527,N_4877);
or U5488 (N_5488,N_3615,N_3596);
xnor U5489 (N_5489,N_2643,N_4646);
nor U5490 (N_5490,N_4212,N_2881);
xor U5491 (N_5491,N_3951,N_4146);
xor U5492 (N_5492,N_4568,N_3807);
nor U5493 (N_5493,N_2899,N_4445);
and U5494 (N_5494,N_4690,N_3409);
nor U5495 (N_5495,N_4032,N_2943);
and U5496 (N_5496,N_4066,N_3304);
xor U5497 (N_5497,N_4164,N_3667);
nand U5498 (N_5498,N_2873,N_4228);
nor U5499 (N_5499,N_3066,N_4069);
nor U5500 (N_5500,N_2649,N_3887);
and U5501 (N_5501,N_4880,N_3993);
or U5502 (N_5502,N_2998,N_4936);
xor U5503 (N_5503,N_4356,N_4650);
or U5504 (N_5504,N_2757,N_2914);
nor U5505 (N_5505,N_3288,N_2721);
nand U5506 (N_5506,N_3725,N_4028);
nor U5507 (N_5507,N_4959,N_3830);
nor U5508 (N_5508,N_4408,N_4790);
nor U5509 (N_5509,N_4942,N_3255);
nand U5510 (N_5510,N_3301,N_4911);
and U5511 (N_5511,N_3296,N_4682);
nor U5512 (N_5512,N_2886,N_3849);
nand U5513 (N_5513,N_4437,N_3082);
nor U5514 (N_5514,N_3101,N_3450);
and U5515 (N_5515,N_4544,N_3018);
or U5516 (N_5516,N_3501,N_3481);
and U5517 (N_5517,N_3630,N_4104);
nor U5518 (N_5518,N_4920,N_3250);
or U5519 (N_5519,N_3410,N_3529);
nor U5520 (N_5520,N_4500,N_2607);
and U5521 (N_5521,N_3758,N_4918);
xor U5522 (N_5522,N_3621,N_4021);
xor U5523 (N_5523,N_4464,N_2772);
xnor U5524 (N_5524,N_3835,N_4481);
and U5525 (N_5525,N_4115,N_4207);
nand U5526 (N_5526,N_4583,N_3901);
and U5527 (N_5527,N_3375,N_3547);
xnor U5528 (N_5528,N_3928,N_2827);
nand U5529 (N_5529,N_2722,N_4939);
or U5530 (N_5530,N_2887,N_3846);
or U5531 (N_5531,N_3313,N_3359);
xor U5532 (N_5532,N_3272,N_4039);
or U5533 (N_5533,N_3239,N_3274);
nand U5534 (N_5534,N_4400,N_3091);
xor U5535 (N_5535,N_3936,N_3546);
nor U5536 (N_5536,N_3856,N_3717);
or U5537 (N_5537,N_4770,N_2689);
xnor U5538 (N_5538,N_3563,N_2983);
nor U5539 (N_5539,N_3407,N_2817);
or U5540 (N_5540,N_4398,N_4469);
and U5541 (N_5541,N_3292,N_3378);
xnor U5542 (N_5542,N_2832,N_4304);
and U5543 (N_5543,N_4415,N_3893);
or U5544 (N_5544,N_2593,N_4397);
xor U5545 (N_5545,N_2550,N_3097);
and U5546 (N_5546,N_4814,N_3103);
or U5547 (N_5547,N_4593,N_2523);
xnor U5548 (N_5548,N_3107,N_2590);
or U5549 (N_5549,N_3401,N_3224);
xor U5550 (N_5550,N_4454,N_3752);
nor U5551 (N_5551,N_2505,N_3999);
and U5552 (N_5552,N_3923,N_4991);
nand U5553 (N_5553,N_4507,N_4194);
nand U5554 (N_5554,N_2937,N_2948);
xor U5555 (N_5555,N_4721,N_2686);
or U5556 (N_5556,N_4971,N_2617);
nor U5557 (N_5557,N_3377,N_4051);
and U5558 (N_5558,N_2651,N_3159);
and U5559 (N_5559,N_3242,N_4273);
nand U5560 (N_5560,N_4041,N_4139);
nor U5561 (N_5561,N_2535,N_3380);
or U5562 (N_5562,N_4542,N_3085);
or U5563 (N_5563,N_3996,N_4749);
xor U5564 (N_5564,N_2571,N_3092);
nand U5565 (N_5565,N_2838,N_4091);
or U5566 (N_5566,N_3330,N_4060);
nor U5567 (N_5567,N_3706,N_3641);
nand U5568 (N_5568,N_3196,N_2952);
and U5569 (N_5569,N_3034,N_3828);
xnor U5570 (N_5570,N_3303,N_4582);
and U5571 (N_5571,N_3404,N_4348);
xnor U5572 (N_5572,N_4403,N_4455);
nor U5573 (N_5573,N_4088,N_4145);
and U5574 (N_5574,N_4960,N_3870);
nor U5575 (N_5575,N_4648,N_4527);
or U5576 (N_5576,N_2715,N_4267);
nor U5577 (N_5577,N_4761,N_3147);
nor U5578 (N_5578,N_4276,N_4235);
nor U5579 (N_5579,N_4363,N_3962);
nand U5580 (N_5580,N_4227,N_4350);
and U5581 (N_5581,N_2891,N_4355);
nand U5582 (N_5582,N_4715,N_3797);
xnor U5583 (N_5583,N_3463,N_4876);
xnor U5584 (N_5584,N_4808,N_2645);
and U5585 (N_5585,N_4002,N_3710);
and U5586 (N_5586,N_2599,N_3019);
xnor U5587 (N_5587,N_4245,N_4298);
nor U5588 (N_5588,N_2966,N_2823);
xnor U5589 (N_5589,N_4518,N_3163);
and U5590 (N_5590,N_4217,N_2674);
xnor U5591 (N_5591,N_2673,N_3484);
and U5592 (N_5592,N_4494,N_2898);
and U5593 (N_5593,N_3428,N_2825);
xor U5594 (N_5594,N_3812,N_3611);
nand U5595 (N_5595,N_4393,N_2990);
xnor U5596 (N_5596,N_4969,N_2789);
or U5597 (N_5597,N_3448,N_2723);
nor U5598 (N_5598,N_2565,N_2799);
nand U5599 (N_5599,N_4531,N_2568);
nand U5600 (N_5600,N_4351,N_3831);
and U5601 (N_5601,N_2602,N_4260);
nor U5602 (N_5602,N_2710,N_4780);
xor U5603 (N_5603,N_4773,N_3486);
nand U5604 (N_5604,N_3102,N_4027);
nor U5605 (N_5605,N_3198,N_3290);
and U5606 (N_5606,N_4884,N_4627);
xor U5607 (N_5607,N_2932,N_3854);
xor U5608 (N_5608,N_3490,N_4238);
xnor U5609 (N_5609,N_3261,N_2728);
xnor U5610 (N_5610,N_4128,N_2925);
nor U5611 (N_5611,N_4717,N_2702);
nand U5612 (N_5612,N_4835,N_4420);
xor U5613 (N_5613,N_2906,N_4188);
and U5614 (N_5614,N_3029,N_3504);
xor U5615 (N_5615,N_3867,N_4426);
nand U5616 (N_5616,N_3056,N_3847);
nand U5617 (N_5617,N_4520,N_2540);
and U5618 (N_5618,N_4705,N_2566);
xnor U5619 (N_5619,N_4354,N_4414);
nand U5620 (N_5620,N_2551,N_4033);
or U5621 (N_5621,N_2971,N_3583);
nor U5622 (N_5622,N_4787,N_4476);
or U5623 (N_5623,N_3430,N_3105);
xnor U5624 (N_5624,N_3083,N_3139);
xnor U5625 (N_5625,N_2605,N_3188);
and U5626 (N_5626,N_3851,N_2934);
or U5627 (N_5627,N_3633,N_4753);
nand U5628 (N_5628,N_4561,N_3426);
and U5629 (N_5629,N_2741,N_2946);
nor U5630 (N_5630,N_3898,N_4834);
nor U5631 (N_5631,N_4964,N_4754);
nand U5632 (N_5632,N_4365,N_2701);
nand U5633 (N_5633,N_3408,N_3724);
or U5634 (N_5634,N_4595,N_3895);
nor U5635 (N_5635,N_3808,N_2888);
xnor U5636 (N_5636,N_3299,N_3431);
nor U5637 (N_5637,N_4843,N_4491);
or U5638 (N_5638,N_4148,N_3680);
and U5639 (N_5639,N_3302,N_4700);
and U5640 (N_5640,N_3562,N_4837);
nor U5641 (N_5641,N_3432,N_3286);
xnor U5642 (N_5642,N_3746,N_3220);
xnor U5643 (N_5643,N_2993,N_3753);
nor U5644 (N_5644,N_2883,N_2580);
xnor U5645 (N_5645,N_4058,N_4031);
nor U5646 (N_5646,N_4549,N_2598);
and U5647 (N_5647,N_4001,N_4023);
or U5648 (N_5648,N_3767,N_4451);
nand U5649 (N_5649,N_4796,N_4957);
or U5650 (N_5650,N_3560,N_4366);
and U5651 (N_5651,N_4172,N_4203);
nand U5652 (N_5652,N_4282,N_4759);
and U5653 (N_5653,N_3722,N_3592);
xnor U5654 (N_5654,N_4410,N_2769);
and U5655 (N_5655,N_4277,N_4793);
or U5656 (N_5656,N_3820,N_2575);
or U5657 (N_5657,N_4418,N_3635);
nor U5658 (N_5658,N_3099,N_2601);
or U5659 (N_5659,N_3356,N_3821);
or U5660 (N_5660,N_3968,N_4670);
or U5661 (N_5661,N_4097,N_3559);
nor U5662 (N_5662,N_4286,N_3372);
nor U5663 (N_5663,N_3544,N_3571);
nor U5664 (N_5664,N_4349,N_2717);
xor U5665 (N_5665,N_4540,N_2553);
nand U5666 (N_5666,N_3661,N_3673);
xnor U5667 (N_5667,N_2711,N_3734);
nand U5668 (N_5668,N_3476,N_2600);
nor U5669 (N_5669,N_4324,N_3852);
and U5670 (N_5670,N_3012,N_3981);
or U5671 (N_5671,N_3582,N_3503);
nand U5672 (N_5672,N_4161,N_4847);
xnor U5673 (N_5673,N_3881,N_3050);
and U5674 (N_5674,N_3367,N_2762);
nand U5675 (N_5675,N_3691,N_4665);
nor U5676 (N_5676,N_4594,N_3218);
and U5677 (N_5677,N_4012,N_3868);
nor U5678 (N_5678,N_3709,N_4311);
xnor U5679 (N_5679,N_3998,N_4109);
xor U5680 (N_5680,N_4169,N_4602);
xor U5681 (N_5681,N_3720,N_2518);
or U5682 (N_5682,N_3694,N_4092);
nand U5683 (N_5683,N_3536,N_3642);
xnor U5684 (N_5684,N_2732,N_4105);
xnor U5685 (N_5685,N_2742,N_2691);
or U5686 (N_5686,N_4293,N_2984);
nand U5687 (N_5687,N_4795,N_4713);
and U5688 (N_5688,N_3961,N_4812);
or U5689 (N_5689,N_3141,N_3664);
and U5690 (N_5690,N_4026,N_3277);
nand U5691 (N_5691,N_4981,N_3665);
nor U5692 (N_5692,N_4478,N_4248);
or U5693 (N_5693,N_3210,N_4528);
nor U5694 (N_5694,N_3479,N_3419);
xor U5695 (N_5695,N_3279,N_2976);
nand U5696 (N_5696,N_3194,N_2791);
and U5697 (N_5697,N_4443,N_3766);
nand U5698 (N_5698,N_2634,N_4624);
and U5699 (N_5699,N_2616,N_2954);
nor U5700 (N_5700,N_3004,N_3447);
nor U5701 (N_5701,N_4200,N_4666);
or U5702 (N_5702,N_3569,N_3697);
xnor U5703 (N_5703,N_4923,N_3116);
and U5704 (N_5704,N_4218,N_4269);
nor U5705 (N_5705,N_3644,N_4836);
xor U5706 (N_5706,N_3632,N_2912);
nor U5707 (N_5707,N_3610,N_2857);
nor U5708 (N_5708,N_3112,N_3270);
nand U5709 (N_5709,N_3521,N_2905);
nor U5710 (N_5710,N_3640,N_3888);
nor U5711 (N_5711,N_2904,N_3000);
and U5712 (N_5712,N_4034,N_4016);
or U5713 (N_5713,N_3214,N_4490);
xor U5714 (N_5714,N_2837,N_4210);
or U5715 (N_5715,N_3358,N_2903);
and U5716 (N_5716,N_4219,N_4934);
xor U5717 (N_5717,N_4070,N_4573);
or U5718 (N_5718,N_4259,N_2692);
or U5719 (N_5719,N_3338,N_4664);
xnor U5720 (N_5720,N_4769,N_3287);
or U5721 (N_5721,N_4778,N_4589);
nand U5722 (N_5722,N_2514,N_4538);
and U5723 (N_5723,N_2703,N_4855);
and U5724 (N_5724,N_4198,N_2704);
or U5725 (N_5725,N_4004,N_3402);
and U5726 (N_5726,N_3643,N_4980);
or U5727 (N_5727,N_4592,N_3843);
xor U5728 (N_5728,N_2964,N_4432);
and U5729 (N_5729,N_4908,N_3202);
nor U5730 (N_5730,N_3075,N_2880);
and U5731 (N_5731,N_3760,N_2924);
nor U5732 (N_5732,N_2759,N_4431);
or U5733 (N_5733,N_4927,N_2913);
nor U5734 (N_5734,N_2918,N_3319);
nor U5735 (N_5735,N_3217,N_3289);
nand U5736 (N_5736,N_4882,N_2820);
xnor U5737 (N_5737,N_4281,N_3927);
xor U5738 (N_5738,N_3412,N_3570);
xnor U5739 (N_5739,N_4098,N_2916);
or U5740 (N_5740,N_4487,N_3423);
nor U5741 (N_5741,N_3726,N_2875);
and U5742 (N_5742,N_4452,N_3514);
xnor U5743 (N_5743,N_4458,N_3573);
and U5744 (N_5744,N_4581,N_3775);
or U5745 (N_5745,N_4279,N_3609);
nand U5746 (N_5746,N_4921,N_3469);
or U5747 (N_5747,N_3485,N_3525);
nand U5748 (N_5748,N_3913,N_4669);
xnor U5749 (N_5749,N_4809,N_4570);
xnor U5750 (N_5750,N_4076,N_4975);
nand U5751 (N_5751,N_4231,N_3971);
nand U5752 (N_5752,N_3588,N_2623);
nand U5753 (N_5753,N_3234,N_4233);
nor U5754 (N_5754,N_4241,N_3910);
and U5755 (N_5755,N_2920,N_3438);
nor U5756 (N_5756,N_3474,N_4049);
xor U5757 (N_5757,N_3907,N_2860);
or U5758 (N_5758,N_4237,N_3787);
and U5759 (N_5759,N_2778,N_4061);
nor U5760 (N_5760,N_4930,N_4289);
xor U5761 (N_5761,N_2828,N_3473);
nor U5762 (N_5762,N_3030,N_4635);
nand U5763 (N_5763,N_4409,N_2785);
nor U5764 (N_5764,N_3235,N_3207);
xnor U5765 (N_5765,N_4136,N_4726);
xor U5766 (N_5766,N_2945,N_3747);
xor U5767 (N_5767,N_3508,N_4090);
xor U5768 (N_5768,N_3371,N_3637);
xor U5769 (N_5769,N_4158,N_2641);
or U5770 (N_5770,N_4967,N_2806);
nand U5771 (N_5771,N_3465,N_4687);
nor U5772 (N_5772,N_2770,N_4159);
xnor U5773 (N_5773,N_2999,N_2821);
or U5774 (N_5774,N_3221,N_4505);
xnor U5775 (N_5775,N_3475,N_4392);
nand U5776 (N_5776,N_3953,N_2675);
xnor U5777 (N_5777,N_3729,N_4086);
xnor U5778 (N_5778,N_4655,N_4151);
nand U5779 (N_5779,N_3420,N_2668);
nor U5780 (N_5780,N_2656,N_4913);
or U5781 (N_5781,N_4508,N_4205);
and U5782 (N_5782,N_4498,N_3676);
nand U5783 (N_5783,N_4383,N_2766);
xnor U5784 (N_5784,N_4746,N_2908);
nor U5785 (N_5785,N_3839,N_4482);
nor U5786 (N_5786,N_3708,N_3424);
nand U5787 (N_5787,N_3055,N_4020);
nor U5788 (N_5788,N_3732,N_2567);
nor U5789 (N_5789,N_4430,N_3284);
or U5790 (N_5790,N_4000,N_2779);
nand U5791 (N_5791,N_4195,N_3926);
nand U5792 (N_5792,N_4193,N_2957);
and U5793 (N_5793,N_4952,N_4607);
xor U5794 (N_5794,N_3741,N_3122);
and U5795 (N_5795,N_4346,N_2749);
and U5796 (N_5796,N_2900,N_3879);
xor U5797 (N_5797,N_3433,N_3532);
and U5798 (N_5798,N_4209,N_4111);
and U5799 (N_5799,N_3520,N_2694);
nand U5800 (N_5800,N_4867,N_3608);
nor U5801 (N_5801,N_3398,N_4797);
and U5802 (N_5802,N_3305,N_4902);
nand U5803 (N_5803,N_3527,N_4063);
and U5804 (N_5804,N_2572,N_4521);
or U5805 (N_5805,N_3539,N_4962);
or U5806 (N_5806,N_4301,N_3298);
and U5807 (N_5807,N_4504,N_3531);
nor U5808 (N_5808,N_3940,N_3627);
nor U5809 (N_5809,N_2533,N_3060);
xor U5810 (N_5810,N_3567,N_4702);
or U5811 (N_5811,N_4879,N_4703);
nor U5812 (N_5812,N_3735,N_4402);
and U5813 (N_5813,N_3674,N_2681);
nand U5814 (N_5814,N_2853,N_2633);
nor U5815 (N_5815,N_3178,N_3456);
xnor U5816 (N_5816,N_4900,N_4294);
and U5817 (N_5817,N_3151,N_3468);
nor U5818 (N_5818,N_2910,N_4554);
or U5819 (N_5819,N_3266,N_3227);
xnor U5820 (N_5820,N_4251,N_2577);
or U5821 (N_5821,N_2618,N_2677);
or U5822 (N_5822,N_3679,N_4215);
and U5823 (N_5823,N_2678,N_3788);
nor U5824 (N_5824,N_4087,N_2611);
nor U5825 (N_5825,N_2676,N_3656);
nand U5826 (N_5826,N_2544,N_3590);
and U5827 (N_5827,N_2793,N_4734);
nand U5828 (N_5828,N_2718,N_3659);
or U5829 (N_5829,N_3161,N_2549);
and U5830 (N_5830,N_3902,N_2929);
xor U5831 (N_5831,N_3499,N_3739);
nor U5832 (N_5832,N_3005,N_3041);
nor U5833 (N_5833,N_4337,N_3446);
or U5834 (N_5834,N_4742,N_4147);
or U5835 (N_5835,N_3215,N_3498);
nor U5836 (N_5836,N_4306,N_4933);
or U5837 (N_5837,N_3068,N_4794);
nor U5838 (N_5838,N_4791,N_3294);
nor U5839 (N_5839,N_4824,N_3666);
and U5840 (N_5840,N_3254,N_3949);
or U5841 (N_5841,N_3059,N_3540);
and U5842 (N_5842,N_4944,N_3859);
nor U5843 (N_5843,N_4805,N_3186);
nand U5844 (N_5844,N_4747,N_3308);
and U5845 (N_5845,N_2798,N_4725);
nand U5846 (N_5846,N_2835,N_3353);
nor U5847 (N_5847,N_3701,N_4833);
nor U5848 (N_5848,N_3723,N_2661);
nor U5849 (N_5849,N_4806,N_3543);
and U5850 (N_5850,N_3781,N_2834);
xor U5851 (N_5851,N_2901,N_3455);
nor U5852 (N_5852,N_4080,N_3938);
or U5853 (N_5853,N_2866,N_2846);
nand U5854 (N_5854,N_2833,N_4054);
xnor U5855 (N_5855,N_4899,N_2852);
nor U5856 (N_5856,N_3545,N_3957);
nand U5857 (N_5857,N_3256,N_3047);
and U5858 (N_5858,N_4854,N_4379);
xor U5859 (N_5859,N_3053,N_3875);
nand U5860 (N_5860,N_2788,N_3441);
and U5861 (N_5861,N_4244,N_4886);
nand U5862 (N_5862,N_3156,N_4789);
nor U5863 (N_5863,N_4974,N_4887);
or U5864 (N_5864,N_4943,N_4804);
or U5865 (N_5865,N_4642,N_4160);
nor U5866 (N_5866,N_4678,N_4865);
or U5867 (N_5867,N_2658,N_3668);
nand U5868 (N_5868,N_3458,N_3191);
nand U5869 (N_5869,N_3634,N_3383);
or U5870 (N_5870,N_3636,N_3049);
xnor U5871 (N_5871,N_2679,N_4973);
nand U5872 (N_5872,N_4941,N_3145);
xor U5873 (N_5873,N_4075,N_4547);
nor U5874 (N_5874,N_4653,N_3654);
nor U5875 (N_5875,N_3598,N_4184);
and U5876 (N_5876,N_3032,N_3394);
nand U5877 (N_5877,N_4326,N_2897);
nand U5878 (N_5878,N_4446,N_2581);
xor U5879 (N_5879,N_3945,N_2615);
or U5880 (N_5880,N_2747,N_4048);
or U5881 (N_5881,N_2872,N_3323);
nor U5882 (N_5882,N_3524,N_4679);
xor U5883 (N_5883,N_4174,N_3128);
xor U5884 (N_5884,N_4557,N_3219);
nor U5885 (N_5885,N_3954,N_3317);
and U5886 (N_5886,N_4331,N_2965);
xor U5887 (N_5887,N_4183,N_3014);
nand U5888 (N_5888,N_2804,N_3150);
or U5889 (N_5889,N_3655,N_4640);
nor U5890 (N_5890,N_4711,N_2882);
nand U5891 (N_5891,N_3599,N_4384);
nand U5892 (N_5892,N_3318,N_3273);
nand U5893 (N_5893,N_3647,N_4680);
and U5894 (N_5894,N_4550,N_3158);
or U5895 (N_5895,N_3826,N_3331);
or U5896 (N_5896,N_4622,N_3119);
xor U5897 (N_5897,N_4681,N_2814);
nor U5898 (N_5898,N_2972,N_3658);
and U5899 (N_5899,N_3415,N_4993);
xnor U5900 (N_5900,N_4309,N_4178);
or U5901 (N_5901,N_4724,N_4609);
xor U5902 (N_5902,N_4534,N_4014);
xnor U5903 (N_5903,N_2628,N_4677);
and U5904 (N_5904,N_4223,N_3869);
or U5905 (N_5905,N_2720,N_2842);
or U5906 (N_5906,N_4716,N_4165);
or U5907 (N_5907,N_3885,N_3603);
nor U5908 (N_5908,N_3991,N_4644);
and U5909 (N_5909,N_3810,N_4449);
and U5910 (N_5910,N_3794,N_3435);
nor U5911 (N_5911,N_3523,N_3714);
or U5912 (N_5912,N_2933,N_3882);
nand U5913 (N_5913,N_4597,N_4138);
xnor U5914 (N_5914,N_3088,N_4656);
and U5915 (N_5915,N_4898,N_2792);
nor U5916 (N_5916,N_4013,N_3225);
nand U5917 (N_5917,N_4057,N_4845);
nor U5918 (N_5918,N_3269,N_3806);
or U5919 (N_5919,N_4517,N_3921);
xor U5920 (N_5920,N_3322,N_3958);
and U5921 (N_5921,N_3069,N_3140);
or U5922 (N_5922,N_4113,N_2790);
xnor U5923 (N_5923,N_2559,N_2504);
nor U5924 (N_5924,N_3789,N_2538);
and U5925 (N_5925,N_2839,N_3505);
or U5926 (N_5926,N_3149,N_4932);
and U5927 (N_5927,N_3281,N_4015);
xnor U5928 (N_5928,N_4988,N_2754);
xnor U5929 (N_5929,N_3631,N_4239);
and U5930 (N_5930,N_3314,N_4869);
and U5931 (N_5931,N_3765,N_4628);
and U5932 (N_5932,N_3779,N_4937);
nand U5933 (N_5933,N_3240,N_3311);
nor U5934 (N_5934,N_2688,N_3933);
nor U5935 (N_5935,N_3494,N_2831);
or U5936 (N_5936,N_3528,N_3369);
or U5937 (N_5937,N_2771,N_3626);
nand U5938 (N_5938,N_3010,N_4842);
nand U5939 (N_5939,N_2830,N_2666);
nor U5940 (N_5940,N_2893,N_2500);
nand U5941 (N_5941,N_4256,N_4546);
nor U5942 (N_5942,N_2753,N_3572);
xnor U5943 (N_5943,N_3950,N_3205);
xnor U5944 (N_5944,N_3388,N_4008);
nand U5945 (N_5945,N_3833,N_4246);
and U5946 (N_5946,N_4983,N_3392);
or U5947 (N_5947,N_4735,N_2537);
nor U5948 (N_5948,N_4325,N_3466);
and U5949 (N_5949,N_3031,N_4340);
nor U5950 (N_5950,N_4503,N_2956);
xnor U5951 (N_5951,N_3336,N_3078);
and U5952 (N_5952,N_2532,N_2684);
xor U5953 (N_5953,N_3321,N_4291);
or U5954 (N_5954,N_4619,N_4587);
and U5955 (N_5955,N_4657,N_4530);
xnor U5956 (N_5956,N_4990,N_2931);
and U5957 (N_5957,N_4436,N_4832);
xor U5958 (N_5958,N_3589,N_2758);
nand U5959 (N_5959,N_3495,N_3008);
xor U5960 (N_5960,N_4270,N_4495);
or U5961 (N_5961,N_3864,N_4950);
and U5962 (N_5962,N_4037,N_3772);
nor U5963 (N_5963,N_4522,N_3162);
or U5964 (N_5964,N_2597,N_4846);
nor U5965 (N_5965,N_3189,N_4488);
nor U5966 (N_5966,N_4171,N_3489);
nor U5967 (N_5967,N_2589,N_4558);
nand U5968 (N_5968,N_4756,N_4234);
and U5969 (N_5969,N_2979,N_2889);
and U5970 (N_5970,N_3117,N_3442);
xor U5971 (N_5971,N_3036,N_4788);
nand U5972 (N_5972,N_3530,N_3551);
nand U5973 (N_5973,N_3942,N_4905);
nand U5974 (N_5974,N_3935,N_4551);
or U5975 (N_5975,N_4144,N_4036);
or U5976 (N_5976,N_3660,N_3883);
nor U5977 (N_5977,N_3108,N_3750);
or U5978 (N_5978,N_3512,N_2775);
xor U5979 (N_5979,N_3944,N_3252);
and U5980 (N_5980,N_3007,N_4722);
and U5981 (N_5981,N_2987,N_2519);
nor U5982 (N_5982,N_4706,N_3783);
xnor U5983 (N_5983,N_4633,N_2810);
xnor U5984 (N_5984,N_4673,N_2781);
xnor U5985 (N_5985,N_4236,N_4214);
and U5986 (N_5986,N_2687,N_3903);
nor U5987 (N_5987,N_3344,N_2982);
nor U5988 (N_5988,N_3537,N_2923);
nor U5989 (N_5989,N_2953,N_4949);
or U5990 (N_5990,N_3932,N_3873);
xnor U5991 (N_5991,N_4149,N_3241);
nand U5992 (N_5992,N_3815,N_2780);
or U5993 (N_5993,N_3591,N_4131);
or U5994 (N_5994,N_3975,N_3064);
xor U5995 (N_5995,N_4860,N_4823);
xnor U5996 (N_5996,N_3581,N_3678);
xnor U5997 (N_5997,N_4660,N_3138);
nor U5998 (N_5998,N_2768,N_4612);
nor U5999 (N_5999,N_4323,N_4475);
nand U6000 (N_6000,N_2826,N_3193);
xnor U6001 (N_6001,N_4278,N_2507);
xnor U6002 (N_6002,N_4081,N_4661);
xor U6003 (N_6003,N_4603,N_2895);
nand U6004 (N_6004,N_4588,N_4141);
nor U6005 (N_6005,N_4658,N_2531);
xor U6006 (N_6006,N_2503,N_4566);
nor U6007 (N_6007,N_4511,N_4196);
and U6008 (N_6008,N_3984,N_3244);
nor U6009 (N_6009,N_4647,N_3263);
nand U6010 (N_6010,N_4539,N_3602);
nor U6011 (N_6011,N_4389,N_4708);
or U6012 (N_6012,N_3862,N_2877);
nand U6013 (N_6013,N_3930,N_3080);
xor U6014 (N_6014,N_4699,N_4167);
and U6015 (N_6015,N_2524,N_3595);
or U6016 (N_6016,N_3175,N_3003);
nor U6017 (N_6017,N_4864,N_4073);
nor U6018 (N_6018,N_4030,N_4643);
xnor U6019 (N_6019,N_3471,N_3552);
and U6020 (N_6020,N_4173,N_4428);
nor U6021 (N_6021,N_2521,N_4625);
or U6022 (N_6022,N_4029,N_3663);
nor U6023 (N_6023,N_3721,N_4448);
and U6024 (N_6024,N_4849,N_4526);
or U6025 (N_6025,N_4274,N_4695);
xnor U6026 (N_6026,N_3180,N_3437);
or U6027 (N_6027,N_4994,N_3743);
nand U6028 (N_6028,N_3345,N_2808);
xnor U6029 (N_6029,N_2962,N_3707);
nand U6030 (N_6030,N_3425,N_3364);
xnor U6031 (N_6031,N_4596,N_4025);
or U6032 (N_6032,N_3912,N_3387);
nor U6033 (N_6033,N_4492,N_4985);
nand U6034 (N_6034,N_4381,N_4401);
and U6035 (N_6035,N_4116,N_2563);
nor U6036 (N_6036,N_4714,N_4737);
nand U6037 (N_6037,N_4513,N_4112);
nand U6038 (N_6038,N_3312,N_3620);
xor U6039 (N_6039,N_3622,N_2975);
nand U6040 (N_6040,N_4765,N_3804);
nor U6041 (N_6041,N_3381,N_4373);
and U6042 (N_6042,N_4720,N_2595);
nor U6043 (N_6043,N_2884,N_2968);
nor U6044 (N_6044,N_4137,N_3451);
nand U6045 (N_6045,N_3689,N_3617);
nor U6046 (N_6046,N_4995,N_2859);
or U6047 (N_6047,N_4799,N_3038);
nor U6048 (N_6048,N_3623,N_3946);
and U6049 (N_6049,N_2942,N_4045);
nor U6050 (N_6050,N_2667,N_3769);
and U6051 (N_6051,N_4064,N_3370);
xnor U6052 (N_6052,N_4729,N_3230);
xor U6053 (N_6053,N_3098,N_2525);
nand U6054 (N_6054,N_4748,N_2959);
nor U6055 (N_6055,N_4743,N_4320);
nand U6056 (N_6056,N_4216,N_4305);
or U6057 (N_6057,N_2786,N_2696);
nor U6058 (N_6058,N_3457,N_2938);
nor U6059 (N_6059,N_4689,N_4620);
and U6060 (N_6060,N_4615,N_3871);
or U6061 (N_6061,N_4781,N_3891);
nor U6062 (N_6062,N_4261,N_2700);
or U6063 (N_6063,N_4986,N_3516);
or U6064 (N_6064,N_3152,N_3125);
xor U6065 (N_6065,N_3251,N_3126);
nor U6066 (N_6066,N_4285,N_3144);
nor U6067 (N_6067,N_4470,N_4224);
xor U6068 (N_6068,N_4182,N_2511);
nor U6069 (N_6069,N_4120,N_2995);
nor U6070 (N_6070,N_4334,N_3109);
or U6071 (N_6071,N_3553,N_4077);
and U6072 (N_6072,N_3136,N_2944);
nand U6073 (N_6073,N_3914,N_4083);
or U6074 (N_6074,N_4850,N_3646);
nand U6075 (N_6075,N_4881,N_3876);
nor U6076 (N_6076,N_3840,N_2625);
nor U6077 (N_6077,N_4247,N_3937);
xor U6078 (N_6078,N_3236,N_3866);
or U6079 (N_6079,N_3756,N_3994);
and U6080 (N_6080,N_3081,N_4757);
and U6081 (N_6081,N_4099,N_4302);
nand U6082 (N_6082,N_2777,N_3057);
xor U6083 (N_6083,N_4473,N_4250);
nand U6084 (N_6084,N_2609,N_3988);
nand U6085 (N_6085,N_3351,N_3334);
nand U6086 (N_6086,N_2763,N_2659);
nor U6087 (N_6087,N_4477,N_3522);
nor U6088 (N_6088,N_2915,N_2977);
and U6089 (N_6089,N_3429,N_2508);
and U6090 (N_6090,N_2705,N_4456);
nor U6091 (N_6091,N_3677,N_2510);
and U6092 (N_6092,N_4315,N_4313);
and U6093 (N_6093,N_2596,N_2919);
nand U6094 (N_6094,N_4327,N_4489);
or U6095 (N_6095,N_2878,N_4559);
nand U6096 (N_6096,N_3315,N_3096);
or U6097 (N_6097,N_3548,N_2558);
and U6098 (N_6098,N_2610,N_4697);
and U6099 (N_6099,N_3382,N_4543);
nand U6100 (N_6100,N_3405,N_4826);
nand U6101 (N_6101,N_3329,N_2621);
xnor U6102 (N_6102,N_4552,N_4710);
and U6103 (N_6103,N_4359,N_4461);
nand U6104 (N_6104,N_3952,N_3157);
nor U6105 (N_6105,N_3974,N_4977);
and U6106 (N_6106,N_3280,N_4191);
xor U6107 (N_6107,N_3337,N_2529);
nor U6108 (N_6108,N_4555,N_4998);
or U6109 (N_6109,N_4919,N_3084);
and U6110 (N_6110,N_3033,N_2671);
and U6111 (N_6111,N_2569,N_3800);
xnor U6112 (N_6112,N_4954,N_2501);
or U6113 (N_6113,N_3208,N_4675);
and U6114 (N_6114,N_3228,N_2890);
nand U6115 (N_6115,N_4606,N_4163);
nand U6116 (N_6116,N_3058,N_4997);
xnor U6117 (N_6117,N_4050,N_2587);
xor U6118 (N_6118,N_2585,N_4046);
or U6119 (N_6119,N_2632,N_2631);
nor U6120 (N_6120,N_4377,N_3384);
nand U6121 (N_6121,N_2554,N_2606);
nand U6122 (N_6122,N_4771,N_3929);
and U6123 (N_6123,N_3155,N_4371);
nand U6124 (N_6124,N_4874,N_3764);
and U6125 (N_6125,N_4502,N_3496);
or U6126 (N_6126,N_2961,N_2635);
nand U6127 (N_6127,N_3845,N_4857);
or U6128 (N_6128,N_3844,N_4621);
or U6129 (N_6129,N_3347,N_4338);
or U6130 (N_6130,N_2564,N_2969);
or U6131 (N_6131,N_3309,N_4450);
nand U6132 (N_6132,N_4364,N_2800);
nor U6133 (N_6133,N_3436,N_2660);
nand U6134 (N_6134,N_4532,N_2871);
nand U6135 (N_6135,N_4114,N_3612);
nand U6136 (N_6136,N_2506,N_3692);
nand U6137 (N_6137,N_2729,N_3061);
nor U6138 (N_6138,N_3515,N_4275);
and U6139 (N_6139,N_3549,N_4893);
and U6140 (N_6140,N_2706,N_3500);
nor U6141 (N_6141,N_4929,N_2604);
or U6142 (N_6142,N_2613,N_4978);
or U6143 (N_6143,N_4121,N_4439);
and U6144 (N_6144,N_4961,N_3541);
and U6145 (N_6145,N_3245,N_4059);
or U6146 (N_6146,N_2698,N_4284);
and U6147 (N_6147,N_3417,N_4232);
and U6148 (N_6148,N_2864,N_2542);
nor U6149 (N_6149,N_3506,N_2735);
xnor U6150 (N_6150,N_4992,N_4987);
or U6151 (N_6151,N_4435,N_4750);
and U6152 (N_6152,N_3693,N_2644);
nor U6153 (N_6153,N_4810,N_3931);
or U6154 (N_6154,N_3035,N_2894);
xnor U6155 (N_6155,N_3915,N_2917);
xor U6156 (N_6156,N_3275,N_4220);
or U6157 (N_6157,N_3065,N_4082);
or U6158 (N_6158,N_3782,N_3690);
or U6159 (N_6159,N_4396,N_3593);
or U6160 (N_6160,N_3613,N_4479);
nor U6161 (N_6161,N_3472,N_4117);
nand U6162 (N_6162,N_2622,N_4676);
nor U6163 (N_6163,N_2851,N_2794);
nor U6164 (N_6164,N_3785,N_2630);
and U6165 (N_6165,N_3257,N_4140);
nor U6166 (N_6166,N_4783,N_3478);
nor U6167 (N_6167,N_4579,N_2578);
xor U6168 (N_6168,N_4634,N_4419);
xor U6169 (N_6169,N_4894,N_2695);
and U6170 (N_6170,N_4421,N_3332);
xor U6171 (N_6171,N_3855,N_3362);
xor U6172 (N_6172,N_2870,N_2824);
xor U6173 (N_6173,N_3385,N_3200);
nand U6174 (N_6174,N_4782,N_4872);
xnor U6175 (N_6175,N_4299,N_4968);
or U6176 (N_6176,N_4662,N_3491);
xnor U6177 (N_6177,N_4776,N_2848);
or U6178 (N_6178,N_3742,N_2862);
or U6179 (N_6179,N_3335,N_3969);
or U6180 (N_6180,N_4067,N_2562);
or U6181 (N_6181,N_2981,N_4253);
nor U6182 (N_6182,N_3803,N_3906);
nor U6183 (N_6183,N_3089,N_3439);
nand U6184 (N_6184,N_2816,N_3651);
nor U6185 (N_6185,N_3801,N_3986);
nor U6186 (N_6186,N_3751,N_2512);
or U6187 (N_6187,N_4645,N_4755);
nor U6188 (N_6188,N_3652,N_3025);
and U6189 (N_6189,N_4966,N_4605);
and U6190 (N_6190,N_4065,N_2947);
nand U6191 (N_6191,N_3165,N_3488);
xnor U6192 (N_6192,N_3837,N_3606);
and U6193 (N_6193,N_2734,N_3406);
xnor U6194 (N_6194,N_3798,N_2996);
and U6195 (N_6195,N_4108,N_3137);
or U6196 (N_6196,N_4213,N_2748);
xnor U6197 (N_6197,N_4825,N_3070);
or U6198 (N_6198,N_4965,N_2555);
and U6199 (N_6199,N_2818,N_4576);
and U6200 (N_6200,N_4255,N_4813);
nand U6201 (N_6201,N_4651,N_3349);
nand U6202 (N_6202,N_4704,N_4292);
xnor U6203 (N_6203,N_3829,N_3841);
nand U6204 (N_6204,N_2850,N_4142);
or U6205 (N_6205,N_4524,N_4926);
nand U6206 (N_6206,N_3925,N_3682);
xnor U6207 (N_6207,N_2935,N_4873);
and U6208 (N_6208,N_4598,N_2662);
xor U6209 (N_6209,N_4005,N_3326);
and U6210 (N_6210,N_3702,N_3825);
or U6211 (N_6211,N_3819,N_3232);
or U6212 (N_6212,N_4287,N_3449);
nand U6213 (N_6213,N_3594,N_3811);
nor U6214 (N_6214,N_4947,N_3786);
and U6215 (N_6215,N_3376,N_3297);
and U6216 (N_6216,N_4303,N_2807);
and U6217 (N_6217,N_2556,N_3134);
nand U6218 (N_6218,N_4996,N_4956);
and U6219 (N_6219,N_4979,N_2868);
xnor U6220 (N_6220,N_2724,N_3672);
and U6221 (N_6221,N_2515,N_4181);
nand U6222 (N_6222,N_4123,N_2867);
nor U6223 (N_6223,N_3226,N_4009);
xnor U6224 (N_6224,N_2579,N_4752);
and U6225 (N_6225,N_3748,N_3222);
or U6226 (N_6226,N_2636,N_2765);
or U6227 (N_6227,N_4474,N_3264);
nor U6228 (N_6228,N_4574,N_4368);
and U6229 (N_6229,N_3502,N_4222);
nand U6230 (N_6230,N_2557,N_4424);
or U6231 (N_6231,N_4878,N_3052);
xor U6232 (N_6232,N_4190,N_4417);
xnor U6233 (N_6233,N_4423,N_3992);
nor U6234 (N_6234,N_3295,N_3248);
or U6235 (N_6235,N_4268,N_3477);
nand U6236 (N_6236,N_3493,N_4485);
nor U6237 (N_6237,N_3616,N_4078);
and U6238 (N_6238,N_4871,N_4264);
nand U6239 (N_6239,N_2716,N_4162);
and U6240 (N_6240,N_4741,N_4316);
and U6241 (N_6241,N_3343,N_3920);
nor U6242 (N_6242,N_4548,N_3467);
nor U6243 (N_6243,N_4317,N_4672);
nand U6244 (N_6244,N_4889,N_3894);
xor U6245 (N_6245,N_3300,N_3307);
xnor U6246 (N_6246,N_2545,N_2767);
xnor U6247 (N_6247,N_4468,N_3880);
nand U6248 (N_6248,N_4484,N_3790);
nand U6249 (N_6249,N_3768,N_4122);
xnor U6250 (N_6250,N_4025,N_3034);
nand U6251 (N_6251,N_4586,N_2584);
xnor U6252 (N_6252,N_2611,N_3484);
nand U6253 (N_6253,N_2806,N_3457);
and U6254 (N_6254,N_4923,N_4296);
nor U6255 (N_6255,N_4282,N_3836);
and U6256 (N_6256,N_3784,N_4497);
and U6257 (N_6257,N_2737,N_3118);
nand U6258 (N_6258,N_4832,N_4532);
or U6259 (N_6259,N_4062,N_4409);
xor U6260 (N_6260,N_4596,N_3411);
or U6261 (N_6261,N_3650,N_3330);
or U6262 (N_6262,N_2597,N_4973);
or U6263 (N_6263,N_3486,N_3290);
or U6264 (N_6264,N_3278,N_3830);
or U6265 (N_6265,N_4154,N_4798);
nand U6266 (N_6266,N_4528,N_4116);
xor U6267 (N_6267,N_3031,N_4152);
or U6268 (N_6268,N_3597,N_3710);
nand U6269 (N_6269,N_2992,N_3224);
or U6270 (N_6270,N_3310,N_4637);
or U6271 (N_6271,N_2683,N_2888);
or U6272 (N_6272,N_3718,N_3615);
xnor U6273 (N_6273,N_2721,N_4402);
nor U6274 (N_6274,N_2850,N_3959);
and U6275 (N_6275,N_4699,N_4777);
nand U6276 (N_6276,N_2821,N_4603);
and U6277 (N_6277,N_3705,N_3993);
nand U6278 (N_6278,N_4328,N_3034);
nand U6279 (N_6279,N_3758,N_4622);
nand U6280 (N_6280,N_2949,N_4870);
xor U6281 (N_6281,N_4024,N_2937);
or U6282 (N_6282,N_4160,N_4263);
xnor U6283 (N_6283,N_3309,N_3922);
nand U6284 (N_6284,N_4945,N_3557);
nor U6285 (N_6285,N_3829,N_2882);
xor U6286 (N_6286,N_2864,N_3573);
nand U6287 (N_6287,N_2946,N_3019);
nand U6288 (N_6288,N_3902,N_4335);
and U6289 (N_6289,N_4983,N_4883);
and U6290 (N_6290,N_3054,N_2674);
or U6291 (N_6291,N_4168,N_3356);
and U6292 (N_6292,N_2642,N_4461);
or U6293 (N_6293,N_4452,N_2689);
nand U6294 (N_6294,N_4610,N_4812);
nand U6295 (N_6295,N_4724,N_3188);
xor U6296 (N_6296,N_2644,N_4989);
xnor U6297 (N_6297,N_4449,N_4519);
or U6298 (N_6298,N_3387,N_4271);
nor U6299 (N_6299,N_4431,N_4876);
and U6300 (N_6300,N_2914,N_3508);
nand U6301 (N_6301,N_4208,N_2970);
xor U6302 (N_6302,N_2974,N_3452);
xnor U6303 (N_6303,N_3801,N_4044);
and U6304 (N_6304,N_3411,N_3664);
or U6305 (N_6305,N_4498,N_2712);
nand U6306 (N_6306,N_4719,N_3496);
xor U6307 (N_6307,N_3250,N_2893);
nand U6308 (N_6308,N_3822,N_3500);
or U6309 (N_6309,N_4011,N_3754);
xor U6310 (N_6310,N_2890,N_4681);
and U6311 (N_6311,N_4375,N_3005);
and U6312 (N_6312,N_4143,N_3450);
or U6313 (N_6313,N_3537,N_3349);
nor U6314 (N_6314,N_4111,N_4777);
xor U6315 (N_6315,N_4260,N_3629);
or U6316 (N_6316,N_2726,N_3188);
and U6317 (N_6317,N_3572,N_4031);
nand U6318 (N_6318,N_4297,N_4254);
or U6319 (N_6319,N_3763,N_2828);
xor U6320 (N_6320,N_4964,N_4900);
or U6321 (N_6321,N_2862,N_3003);
and U6322 (N_6322,N_3980,N_4256);
nand U6323 (N_6323,N_4946,N_3895);
nand U6324 (N_6324,N_2781,N_4032);
or U6325 (N_6325,N_4597,N_3225);
nor U6326 (N_6326,N_4397,N_4969);
nand U6327 (N_6327,N_4924,N_4883);
or U6328 (N_6328,N_4099,N_2558);
xnor U6329 (N_6329,N_2528,N_4821);
nand U6330 (N_6330,N_3830,N_4477);
nand U6331 (N_6331,N_2616,N_4449);
nor U6332 (N_6332,N_4326,N_2564);
xor U6333 (N_6333,N_4676,N_4403);
and U6334 (N_6334,N_3833,N_4820);
xnor U6335 (N_6335,N_3907,N_2630);
nand U6336 (N_6336,N_3892,N_4013);
nor U6337 (N_6337,N_4410,N_4012);
nor U6338 (N_6338,N_4844,N_4181);
nand U6339 (N_6339,N_2660,N_3016);
and U6340 (N_6340,N_4703,N_3484);
xor U6341 (N_6341,N_2688,N_4366);
xor U6342 (N_6342,N_2756,N_3592);
nand U6343 (N_6343,N_3073,N_4756);
nor U6344 (N_6344,N_4949,N_2607);
or U6345 (N_6345,N_4471,N_3067);
nor U6346 (N_6346,N_3093,N_3936);
xor U6347 (N_6347,N_3309,N_3859);
nand U6348 (N_6348,N_3023,N_4492);
and U6349 (N_6349,N_4891,N_4993);
nor U6350 (N_6350,N_3400,N_4975);
nor U6351 (N_6351,N_4464,N_4363);
nor U6352 (N_6352,N_4924,N_4012);
and U6353 (N_6353,N_2796,N_4017);
nor U6354 (N_6354,N_4721,N_4309);
xnor U6355 (N_6355,N_4705,N_3014);
or U6356 (N_6356,N_3404,N_2539);
and U6357 (N_6357,N_3346,N_4468);
and U6358 (N_6358,N_3100,N_3038);
nor U6359 (N_6359,N_4734,N_2865);
nand U6360 (N_6360,N_2694,N_3645);
nor U6361 (N_6361,N_4657,N_4654);
nand U6362 (N_6362,N_2655,N_4585);
and U6363 (N_6363,N_3267,N_4099);
nor U6364 (N_6364,N_4009,N_2788);
or U6365 (N_6365,N_3508,N_3698);
xnor U6366 (N_6366,N_3301,N_2947);
xnor U6367 (N_6367,N_4664,N_4769);
nor U6368 (N_6368,N_4286,N_4180);
or U6369 (N_6369,N_2729,N_4899);
nor U6370 (N_6370,N_3462,N_4185);
xnor U6371 (N_6371,N_4671,N_3566);
xor U6372 (N_6372,N_2675,N_4095);
and U6373 (N_6373,N_4487,N_3376);
and U6374 (N_6374,N_3974,N_3165);
or U6375 (N_6375,N_4133,N_3604);
and U6376 (N_6376,N_3629,N_3071);
nand U6377 (N_6377,N_4356,N_4167);
and U6378 (N_6378,N_2704,N_2520);
nor U6379 (N_6379,N_3694,N_3973);
nor U6380 (N_6380,N_4533,N_4442);
and U6381 (N_6381,N_3027,N_4410);
nor U6382 (N_6382,N_4322,N_4944);
nor U6383 (N_6383,N_2501,N_4466);
and U6384 (N_6384,N_3222,N_2661);
nor U6385 (N_6385,N_3270,N_3863);
xor U6386 (N_6386,N_3328,N_3085);
or U6387 (N_6387,N_3039,N_3608);
xnor U6388 (N_6388,N_2727,N_4352);
and U6389 (N_6389,N_4720,N_3022);
xnor U6390 (N_6390,N_3067,N_4867);
nand U6391 (N_6391,N_2745,N_4871);
xnor U6392 (N_6392,N_4228,N_4202);
nand U6393 (N_6393,N_4478,N_4358);
nand U6394 (N_6394,N_4389,N_2597);
or U6395 (N_6395,N_3179,N_3577);
and U6396 (N_6396,N_4557,N_3362);
nand U6397 (N_6397,N_3959,N_4833);
nor U6398 (N_6398,N_4501,N_4481);
or U6399 (N_6399,N_2611,N_3025);
and U6400 (N_6400,N_4280,N_2693);
and U6401 (N_6401,N_2745,N_3998);
nor U6402 (N_6402,N_4115,N_4809);
xnor U6403 (N_6403,N_2567,N_3445);
or U6404 (N_6404,N_4711,N_3526);
xnor U6405 (N_6405,N_4909,N_3820);
nor U6406 (N_6406,N_3776,N_4095);
nor U6407 (N_6407,N_4032,N_4298);
or U6408 (N_6408,N_3409,N_2764);
nand U6409 (N_6409,N_4683,N_4825);
nand U6410 (N_6410,N_4669,N_3647);
xor U6411 (N_6411,N_3966,N_2868);
xor U6412 (N_6412,N_2907,N_3009);
and U6413 (N_6413,N_4066,N_2766);
and U6414 (N_6414,N_2967,N_4988);
or U6415 (N_6415,N_4214,N_3619);
nand U6416 (N_6416,N_3620,N_4750);
nand U6417 (N_6417,N_3655,N_2778);
nor U6418 (N_6418,N_4290,N_3803);
nor U6419 (N_6419,N_2892,N_2645);
nand U6420 (N_6420,N_4298,N_3965);
or U6421 (N_6421,N_4182,N_4836);
xor U6422 (N_6422,N_2807,N_3828);
xor U6423 (N_6423,N_4215,N_4345);
nor U6424 (N_6424,N_2826,N_4384);
or U6425 (N_6425,N_4457,N_3462);
or U6426 (N_6426,N_2933,N_2595);
and U6427 (N_6427,N_3785,N_3443);
and U6428 (N_6428,N_4497,N_2667);
nand U6429 (N_6429,N_3162,N_3811);
or U6430 (N_6430,N_4893,N_4444);
nor U6431 (N_6431,N_4407,N_3205);
or U6432 (N_6432,N_3206,N_4082);
nand U6433 (N_6433,N_3596,N_4582);
xor U6434 (N_6434,N_4575,N_4756);
nand U6435 (N_6435,N_4270,N_3208);
nor U6436 (N_6436,N_3388,N_3600);
nor U6437 (N_6437,N_4270,N_2778);
nor U6438 (N_6438,N_3178,N_3644);
nand U6439 (N_6439,N_4555,N_3755);
or U6440 (N_6440,N_2993,N_3939);
nand U6441 (N_6441,N_2520,N_3587);
and U6442 (N_6442,N_3198,N_4481);
or U6443 (N_6443,N_4327,N_3063);
or U6444 (N_6444,N_3717,N_3926);
nand U6445 (N_6445,N_3451,N_2779);
or U6446 (N_6446,N_4613,N_2503);
and U6447 (N_6447,N_3005,N_3425);
or U6448 (N_6448,N_3773,N_3088);
xor U6449 (N_6449,N_3396,N_4379);
xnor U6450 (N_6450,N_2935,N_2999);
nor U6451 (N_6451,N_3977,N_3727);
or U6452 (N_6452,N_4285,N_4789);
or U6453 (N_6453,N_3556,N_4077);
or U6454 (N_6454,N_4219,N_4070);
xor U6455 (N_6455,N_2904,N_4645);
xnor U6456 (N_6456,N_4123,N_4682);
and U6457 (N_6457,N_4762,N_3217);
or U6458 (N_6458,N_4141,N_3370);
xnor U6459 (N_6459,N_3151,N_4031);
nor U6460 (N_6460,N_4426,N_4563);
xor U6461 (N_6461,N_3529,N_4640);
nor U6462 (N_6462,N_4171,N_3356);
xnor U6463 (N_6463,N_4583,N_4527);
or U6464 (N_6464,N_3951,N_3204);
xor U6465 (N_6465,N_3411,N_3441);
nor U6466 (N_6466,N_4939,N_2690);
nand U6467 (N_6467,N_2536,N_3252);
or U6468 (N_6468,N_4915,N_4127);
nand U6469 (N_6469,N_2509,N_2558);
nor U6470 (N_6470,N_3716,N_3812);
nor U6471 (N_6471,N_3830,N_3039);
and U6472 (N_6472,N_2957,N_4247);
xnor U6473 (N_6473,N_2749,N_3940);
xnor U6474 (N_6474,N_3280,N_3688);
nor U6475 (N_6475,N_3570,N_2741);
nor U6476 (N_6476,N_4286,N_4473);
and U6477 (N_6477,N_3505,N_2538);
or U6478 (N_6478,N_3985,N_4787);
or U6479 (N_6479,N_2544,N_2744);
xor U6480 (N_6480,N_3764,N_4304);
xor U6481 (N_6481,N_3469,N_2952);
nand U6482 (N_6482,N_4431,N_3070);
or U6483 (N_6483,N_4842,N_4267);
xnor U6484 (N_6484,N_3237,N_3641);
xor U6485 (N_6485,N_4651,N_4141);
and U6486 (N_6486,N_2918,N_3288);
nor U6487 (N_6487,N_4950,N_3688);
nand U6488 (N_6488,N_2881,N_3800);
nor U6489 (N_6489,N_2824,N_4579);
or U6490 (N_6490,N_4517,N_2910);
nor U6491 (N_6491,N_4546,N_2907);
and U6492 (N_6492,N_2797,N_2901);
xnor U6493 (N_6493,N_3809,N_3215);
nand U6494 (N_6494,N_3964,N_3922);
and U6495 (N_6495,N_4532,N_4215);
xor U6496 (N_6496,N_2564,N_2649);
xnor U6497 (N_6497,N_3381,N_4601);
xnor U6498 (N_6498,N_3728,N_3635);
and U6499 (N_6499,N_4219,N_3471);
xnor U6500 (N_6500,N_3872,N_4430);
nand U6501 (N_6501,N_4797,N_2619);
nor U6502 (N_6502,N_3158,N_3939);
and U6503 (N_6503,N_3193,N_3605);
or U6504 (N_6504,N_3708,N_4075);
and U6505 (N_6505,N_4591,N_3303);
and U6506 (N_6506,N_4498,N_4218);
or U6507 (N_6507,N_3691,N_3761);
and U6508 (N_6508,N_4829,N_4103);
xor U6509 (N_6509,N_4497,N_4859);
and U6510 (N_6510,N_2662,N_3679);
nand U6511 (N_6511,N_4817,N_3638);
xor U6512 (N_6512,N_4559,N_2709);
nor U6513 (N_6513,N_4908,N_3907);
and U6514 (N_6514,N_4164,N_4485);
nor U6515 (N_6515,N_4687,N_4196);
and U6516 (N_6516,N_4450,N_4642);
or U6517 (N_6517,N_2711,N_2986);
and U6518 (N_6518,N_3032,N_3375);
and U6519 (N_6519,N_4051,N_3329);
nor U6520 (N_6520,N_3054,N_4607);
and U6521 (N_6521,N_3671,N_2578);
and U6522 (N_6522,N_4106,N_4013);
and U6523 (N_6523,N_4973,N_3322);
xor U6524 (N_6524,N_2712,N_2868);
or U6525 (N_6525,N_4193,N_2559);
and U6526 (N_6526,N_3843,N_2776);
and U6527 (N_6527,N_4439,N_2790);
nand U6528 (N_6528,N_4519,N_2540);
nor U6529 (N_6529,N_3827,N_3258);
nand U6530 (N_6530,N_2714,N_3582);
nor U6531 (N_6531,N_2743,N_3813);
nand U6532 (N_6532,N_3343,N_2731);
nor U6533 (N_6533,N_2957,N_2836);
nand U6534 (N_6534,N_4199,N_3361);
nor U6535 (N_6535,N_3470,N_4885);
and U6536 (N_6536,N_4465,N_3447);
xor U6537 (N_6537,N_4572,N_3897);
xnor U6538 (N_6538,N_3063,N_3284);
or U6539 (N_6539,N_3148,N_4855);
and U6540 (N_6540,N_3865,N_4461);
or U6541 (N_6541,N_2978,N_3647);
and U6542 (N_6542,N_3002,N_3220);
xnor U6543 (N_6543,N_3263,N_2943);
xor U6544 (N_6544,N_4935,N_3554);
xor U6545 (N_6545,N_3216,N_4261);
and U6546 (N_6546,N_3213,N_3393);
nor U6547 (N_6547,N_2526,N_3752);
xnor U6548 (N_6548,N_4410,N_2524);
nand U6549 (N_6549,N_4698,N_3163);
and U6550 (N_6550,N_2669,N_3813);
xnor U6551 (N_6551,N_3961,N_3437);
nand U6552 (N_6552,N_4297,N_3134);
and U6553 (N_6553,N_2961,N_3864);
xor U6554 (N_6554,N_2915,N_2787);
or U6555 (N_6555,N_4948,N_4392);
nor U6556 (N_6556,N_4728,N_3061);
nor U6557 (N_6557,N_4545,N_3650);
or U6558 (N_6558,N_2988,N_3042);
nor U6559 (N_6559,N_4934,N_3333);
or U6560 (N_6560,N_4181,N_3539);
and U6561 (N_6561,N_4456,N_4802);
and U6562 (N_6562,N_3721,N_4596);
nand U6563 (N_6563,N_3011,N_3794);
and U6564 (N_6564,N_2928,N_3192);
nor U6565 (N_6565,N_3295,N_4314);
nand U6566 (N_6566,N_3417,N_4781);
and U6567 (N_6567,N_3163,N_4595);
nor U6568 (N_6568,N_3445,N_4659);
nand U6569 (N_6569,N_3349,N_4476);
or U6570 (N_6570,N_4242,N_3229);
xnor U6571 (N_6571,N_4547,N_2562);
or U6572 (N_6572,N_3362,N_2924);
or U6573 (N_6573,N_4097,N_4716);
xnor U6574 (N_6574,N_3961,N_4450);
xnor U6575 (N_6575,N_4526,N_4201);
nor U6576 (N_6576,N_3062,N_4270);
xor U6577 (N_6577,N_4039,N_4984);
or U6578 (N_6578,N_3767,N_3168);
nor U6579 (N_6579,N_3220,N_2923);
nor U6580 (N_6580,N_4083,N_3274);
nor U6581 (N_6581,N_4650,N_4941);
nand U6582 (N_6582,N_3166,N_2910);
xnor U6583 (N_6583,N_3036,N_3123);
nand U6584 (N_6584,N_2863,N_3956);
or U6585 (N_6585,N_4361,N_4035);
xnor U6586 (N_6586,N_2912,N_4428);
and U6587 (N_6587,N_3959,N_3690);
and U6588 (N_6588,N_4629,N_3454);
nand U6589 (N_6589,N_4140,N_3891);
and U6590 (N_6590,N_4108,N_2757);
xnor U6591 (N_6591,N_3285,N_4744);
xnor U6592 (N_6592,N_3024,N_4372);
xor U6593 (N_6593,N_3220,N_2810);
nand U6594 (N_6594,N_2814,N_2711);
nor U6595 (N_6595,N_3651,N_3668);
or U6596 (N_6596,N_4162,N_3600);
xor U6597 (N_6597,N_3275,N_3769);
xnor U6598 (N_6598,N_4409,N_4207);
nand U6599 (N_6599,N_2921,N_4252);
nor U6600 (N_6600,N_2529,N_3524);
or U6601 (N_6601,N_2588,N_4499);
or U6602 (N_6602,N_2861,N_3711);
nor U6603 (N_6603,N_4553,N_3244);
or U6604 (N_6604,N_3788,N_4430);
or U6605 (N_6605,N_4337,N_3923);
xnor U6606 (N_6606,N_4233,N_4185);
nand U6607 (N_6607,N_3712,N_3299);
and U6608 (N_6608,N_3961,N_4469);
xnor U6609 (N_6609,N_2524,N_3488);
xnor U6610 (N_6610,N_4759,N_4262);
or U6611 (N_6611,N_4243,N_3794);
and U6612 (N_6612,N_2566,N_4901);
xnor U6613 (N_6613,N_2742,N_3347);
xnor U6614 (N_6614,N_4628,N_2635);
or U6615 (N_6615,N_3254,N_3347);
and U6616 (N_6616,N_2843,N_3735);
or U6617 (N_6617,N_2762,N_4765);
nand U6618 (N_6618,N_4868,N_2941);
nor U6619 (N_6619,N_3295,N_4247);
and U6620 (N_6620,N_2787,N_4327);
nor U6621 (N_6621,N_3868,N_3130);
or U6622 (N_6622,N_3050,N_2665);
xnor U6623 (N_6623,N_3493,N_3180);
nand U6624 (N_6624,N_3026,N_2990);
and U6625 (N_6625,N_3595,N_4140);
nand U6626 (N_6626,N_3092,N_3372);
nor U6627 (N_6627,N_3391,N_3984);
nor U6628 (N_6628,N_2668,N_4060);
or U6629 (N_6629,N_4035,N_3590);
and U6630 (N_6630,N_3332,N_3989);
xnor U6631 (N_6631,N_2507,N_4265);
xor U6632 (N_6632,N_4773,N_3073);
nor U6633 (N_6633,N_3433,N_2514);
or U6634 (N_6634,N_4976,N_3183);
nor U6635 (N_6635,N_3978,N_4132);
xnor U6636 (N_6636,N_3603,N_3766);
xor U6637 (N_6637,N_3944,N_3652);
or U6638 (N_6638,N_2837,N_3917);
nor U6639 (N_6639,N_2540,N_4564);
nor U6640 (N_6640,N_4630,N_3733);
nor U6641 (N_6641,N_3372,N_2885);
xor U6642 (N_6642,N_4173,N_4649);
or U6643 (N_6643,N_3260,N_4369);
nor U6644 (N_6644,N_3451,N_4918);
nand U6645 (N_6645,N_3590,N_4315);
nand U6646 (N_6646,N_2773,N_3059);
nand U6647 (N_6647,N_3869,N_2598);
nor U6648 (N_6648,N_4783,N_2657);
xor U6649 (N_6649,N_2578,N_4192);
or U6650 (N_6650,N_4205,N_3694);
nor U6651 (N_6651,N_2917,N_4718);
or U6652 (N_6652,N_3570,N_3931);
xor U6653 (N_6653,N_4155,N_4186);
or U6654 (N_6654,N_4574,N_2643);
or U6655 (N_6655,N_3197,N_2663);
xor U6656 (N_6656,N_4211,N_3366);
xor U6657 (N_6657,N_3637,N_4487);
and U6658 (N_6658,N_4114,N_3411);
xor U6659 (N_6659,N_4706,N_4253);
or U6660 (N_6660,N_4446,N_3816);
and U6661 (N_6661,N_4750,N_2652);
and U6662 (N_6662,N_3943,N_3091);
nor U6663 (N_6663,N_2742,N_3275);
nor U6664 (N_6664,N_2614,N_3591);
nor U6665 (N_6665,N_4241,N_3987);
nand U6666 (N_6666,N_4724,N_3235);
and U6667 (N_6667,N_4474,N_4505);
or U6668 (N_6668,N_4896,N_2976);
and U6669 (N_6669,N_3290,N_3001);
or U6670 (N_6670,N_4015,N_4998);
nand U6671 (N_6671,N_4318,N_4338);
xnor U6672 (N_6672,N_3096,N_2984);
nand U6673 (N_6673,N_3121,N_3628);
nand U6674 (N_6674,N_4592,N_2677);
nor U6675 (N_6675,N_2817,N_4197);
nor U6676 (N_6676,N_4014,N_4669);
nand U6677 (N_6677,N_2657,N_4317);
xor U6678 (N_6678,N_3853,N_4334);
nand U6679 (N_6679,N_3506,N_4456);
and U6680 (N_6680,N_3608,N_4302);
and U6681 (N_6681,N_3866,N_4879);
nand U6682 (N_6682,N_4726,N_3963);
nor U6683 (N_6683,N_2742,N_3574);
nand U6684 (N_6684,N_4918,N_4937);
nand U6685 (N_6685,N_3490,N_4068);
nand U6686 (N_6686,N_3028,N_3143);
nand U6687 (N_6687,N_3186,N_4566);
and U6688 (N_6688,N_2926,N_4973);
and U6689 (N_6689,N_2966,N_4503);
nand U6690 (N_6690,N_2700,N_3419);
and U6691 (N_6691,N_3332,N_3626);
or U6692 (N_6692,N_3519,N_3156);
nor U6693 (N_6693,N_3276,N_2619);
nor U6694 (N_6694,N_4044,N_2706);
or U6695 (N_6695,N_3228,N_3671);
xnor U6696 (N_6696,N_2890,N_2638);
xnor U6697 (N_6697,N_4811,N_3295);
nand U6698 (N_6698,N_3754,N_4571);
or U6699 (N_6699,N_4310,N_2844);
nor U6700 (N_6700,N_2763,N_4527);
xor U6701 (N_6701,N_3193,N_3467);
nand U6702 (N_6702,N_3602,N_2584);
nand U6703 (N_6703,N_4215,N_3031);
nand U6704 (N_6704,N_4723,N_3315);
and U6705 (N_6705,N_3942,N_3946);
xor U6706 (N_6706,N_4383,N_4142);
nor U6707 (N_6707,N_2969,N_3117);
nor U6708 (N_6708,N_4126,N_4227);
and U6709 (N_6709,N_2803,N_2881);
xnor U6710 (N_6710,N_2780,N_2652);
and U6711 (N_6711,N_3933,N_3896);
or U6712 (N_6712,N_4461,N_4135);
nor U6713 (N_6713,N_3532,N_4363);
xor U6714 (N_6714,N_2767,N_4823);
xnor U6715 (N_6715,N_3947,N_3080);
and U6716 (N_6716,N_2854,N_2988);
nor U6717 (N_6717,N_4648,N_3780);
nand U6718 (N_6718,N_3131,N_4231);
and U6719 (N_6719,N_3729,N_3541);
xor U6720 (N_6720,N_3384,N_3155);
nand U6721 (N_6721,N_2619,N_4517);
xnor U6722 (N_6722,N_4926,N_4614);
xor U6723 (N_6723,N_4300,N_3707);
and U6724 (N_6724,N_2548,N_2778);
nor U6725 (N_6725,N_2597,N_3953);
xnor U6726 (N_6726,N_4629,N_4197);
xnor U6727 (N_6727,N_2846,N_3203);
or U6728 (N_6728,N_4835,N_3638);
xor U6729 (N_6729,N_4242,N_3507);
nand U6730 (N_6730,N_4475,N_4907);
xnor U6731 (N_6731,N_3448,N_2506);
and U6732 (N_6732,N_3322,N_4726);
xor U6733 (N_6733,N_3516,N_2651);
or U6734 (N_6734,N_4487,N_4154);
nand U6735 (N_6735,N_4916,N_4917);
nor U6736 (N_6736,N_4489,N_4569);
nand U6737 (N_6737,N_2980,N_3160);
xor U6738 (N_6738,N_4081,N_3315);
nor U6739 (N_6739,N_3915,N_3918);
xnor U6740 (N_6740,N_4991,N_4145);
or U6741 (N_6741,N_4747,N_4978);
nand U6742 (N_6742,N_2892,N_4630);
nor U6743 (N_6743,N_3548,N_3612);
xor U6744 (N_6744,N_2957,N_3573);
nand U6745 (N_6745,N_4059,N_4377);
xnor U6746 (N_6746,N_3997,N_4812);
and U6747 (N_6747,N_3071,N_3977);
xor U6748 (N_6748,N_2763,N_4581);
xor U6749 (N_6749,N_3368,N_2646);
and U6750 (N_6750,N_3822,N_3368);
nor U6751 (N_6751,N_4938,N_4198);
and U6752 (N_6752,N_2500,N_3844);
nor U6753 (N_6753,N_3633,N_4933);
nand U6754 (N_6754,N_4724,N_4465);
xnor U6755 (N_6755,N_4405,N_4556);
xnor U6756 (N_6756,N_4533,N_3528);
nor U6757 (N_6757,N_4757,N_4966);
nor U6758 (N_6758,N_4262,N_4315);
or U6759 (N_6759,N_3304,N_2574);
nand U6760 (N_6760,N_4162,N_4595);
nand U6761 (N_6761,N_3117,N_2629);
nand U6762 (N_6762,N_4182,N_3485);
nor U6763 (N_6763,N_4186,N_2751);
or U6764 (N_6764,N_4555,N_4728);
or U6765 (N_6765,N_3899,N_4533);
nor U6766 (N_6766,N_3253,N_2564);
and U6767 (N_6767,N_3135,N_4908);
nor U6768 (N_6768,N_4703,N_4126);
nor U6769 (N_6769,N_4279,N_4880);
xnor U6770 (N_6770,N_2591,N_4270);
and U6771 (N_6771,N_4093,N_3374);
nor U6772 (N_6772,N_3937,N_4381);
nor U6773 (N_6773,N_2912,N_4929);
nor U6774 (N_6774,N_2511,N_3956);
nand U6775 (N_6775,N_4128,N_2588);
and U6776 (N_6776,N_4680,N_4223);
or U6777 (N_6777,N_4277,N_4142);
nor U6778 (N_6778,N_2910,N_4199);
and U6779 (N_6779,N_4317,N_4512);
or U6780 (N_6780,N_3308,N_3377);
and U6781 (N_6781,N_4824,N_3630);
nor U6782 (N_6782,N_3928,N_3355);
nor U6783 (N_6783,N_4091,N_3940);
xor U6784 (N_6784,N_2786,N_4243);
xor U6785 (N_6785,N_2629,N_4778);
or U6786 (N_6786,N_4912,N_3514);
nor U6787 (N_6787,N_3775,N_2631);
nor U6788 (N_6788,N_4232,N_3616);
nand U6789 (N_6789,N_2583,N_4894);
nor U6790 (N_6790,N_4040,N_4758);
or U6791 (N_6791,N_3284,N_4657);
xor U6792 (N_6792,N_2654,N_2562);
xor U6793 (N_6793,N_3765,N_3370);
xnor U6794 (N_6794,N_2831,N_4871);
or U6795 (N_6795,N_3445,N_4272);
or U6796 (N_6796,N_4413,N_2737);
or U6797 (N_6797,N_4844,N_4920);
xor U6798 (N_6798,N_4632,N_4013);
nand U6799 (N_6799,N_3870,N_4127);
and U6800 (N_6800,N_2532,N_3155);
nor U6801 (N_6801,N_4038,N_3864);
or U6802 (N_6802,N_4288,N_2840);
nand U6803 (N_6803,N_2535,N_4836);
nand U6804 (N_6804,N_4447,N_2847);
or U6805 (N_6805,N_4440,N_3859);
nand U6806 (N_6806,N_4956,N_2951);
or U6807 (N_6807,N_4899,N_4637);
nor U6808 (N_6808,N_4490,N_2928);
nor U6809 (N_6809,N_4894,N_4766);
nor U6810 (N_6810,N_3723,N_3090);
xnor U6811 (N_6811,N_4839,N_4486);
nand U6812 (N_6812,N_4582,N_4917);
and U6813 (N_6813,N_4109,N_4302);
xor U6814 (N_6814,N_2711,N_2508);
xor U6815 (N_6815,N_4362,N_2713);
nor U6816 (N_6816,N_2576,N_4179);
nand U6817 (N_6817,N_2838,N_4416);
nor U6818 (N_6818,N_2999,N_3497);
and U6819 (N_6819,N_4138,N_3747);
nor U6820 (N_6820,N_2707,N_4686);
and U6821 (N_6821,N_2558,N_3994);
or U6822 (N_6822,N_4885,N_4911);
xor U6823 (N_6823,N_2932,N_4748);
nor U6824 (N_6824,N_3178,N_3933);
xnor U6825 (N_6825,N_4451,N_4308);
nand U6826 (N_6826,N_4421,N_4314);
nand U6827 (N_6827,N_3466,N_4057);
nand U6828 (N_6828,N_2718,N_4242);
or U6829 (N_6829,N_3528,N_3125);
nand U6830 (N_6830,N_2923,N_4496);
xor U6831 (N_6831,N_2572,N_3369);
or U6832 (N_6832,N_4301,N_4528);
and U6833 (N_6833,N_3078,N_3805);
or U6834 (N_6834,N_2691,N_4252);
nand U6835 (N_6835,N_2749,N_3557);
xor U6836 (N_6836,N_4612,N_4981);
nor U6837 (N_6837,N_3764,N_2560);
or U6838 (N_6838,N_4539,N_2538);
xnor U6839 (N_6839,N_4482,N_4483);
nor U6840 (N_6840,N_4165,N_2836);
xor U6841 (N_6841,N_2814,N_3862);
nor U6842 (N_6842,N_4766,N_4137);
nand U6843 (N_6843,N_4333,N_2745);
xor U6844 (N_6844,N_4069,N_3657);
nor U6845 (N_6845,N_3977,N_3962);
or U6846 (N_6846,N_4009,N_3905);
nand U6847 (N_6847,N_3168,N_2912);
nor U6848 (N_6848,N_4143,N_3821);
xor U6849 (N_6849,N_3740,N_3726);
and U6850 (N_6850,N_4230,N_2724);
or U6851 (N_6851,N_4386,N_3173);
or U6852 (N_6852,N_3485,N_4502);
nand U6853 (N_6853,N_3339,N_3579);
nand U6854 (N_6854,N_4500,N_3828);
or U6855 (N_6855,N_4461,N_2975);
nand U6856 (N_6856,N_4937,N_4725);
or U6857 (N_6857,N_3624,N_4314);
nand U6858 (N_6858,N_4850,N_2773);
nand U6859 (N_6859,N_4825,N_3500);
nor U6860 (N_6860,N_3745,N_2503);
xnor U6861 (N_6861,N_3305,N_2582);
and U6862 (N_6862,N_4305,N_4002);
or U6863 (N_6863,N_4346,N_4429);
xor U6864 (N_6864,N_3269,N_4152);
nand U6865 (N_6865,N_3265,N_4269);
and U6866 (N_6866,N_4892,N_3733);
nand U6867 (N_6867,N_4867,N_3326);
or U6868 (N_6868,N_4715,N_2692);
nor U6869 (N_6869,N_3214,N_3130);
nor U6870 (N_6870,N_4319,N_3106);
and U6871 (N_6871,N_2689,N_4108);
or U6872 (N_6872,N_4189,N_3633);
nor U6873 (N_6873,N_3946,N_3560);
nor U6874 (N_6874,N_3751,N_4426);
and U6875 (N_6875,N_4805,N_4750);
and U6876 (N_6876,N_3096,N_3442);
nor U6877 (N_6877,N_3831,N_3041);
xnor U6878 (N_6878,N_2767,N_4323);
nand U6879 (N_6879,N_4091,N_2743);
xor U6880 (N_6880,N_2626,N_4716);
and U6881 (N_6881,N_2851,N_3822);
nor U6882 (N_6882,N_3318,N_3569);
xor U6883 (N_6883,N_3577,N_2735);
and U6884 (N_6884,N_4942,N_2504);
or U6885 (N_6885,N_2636,N_4011);
or U6886 (N_6886,N_4470,N_3380);
nand U6887 (N_6887,N_4015,N_3403);
or U6888 (N_6888,N_3900,N_4181);
or U6889 (N_6889,N_4239,N_4972);
xor U6890 (N_6890,N_2721,N_3899);
xnor U6891 (N_6891,N_2945,N_3524);
or U6892 (N_6892,N_4278,N_3281);
nor U6893 (N_6893,N_4987,N_2707);
nand U6894 (N_6894,N_2792,N_4521);
xnor U6895 (N_6895,N_3339,N_3108);
nand U6896 (N_6896,N_3723,N_3367);
xnor U6897 (N_6897,N_3382,N_4025);
xor U6898 (N_6898,N_3900,N_4159);
and U6899 (N_6899,N_3582,N_4071);
nand U6900 (N_6900,N_4022,N_3100);
nor U6901 (N_6901,N_4479,N_4104);
and U6902 (N_6902,N_4857,N_4793);
xor U6903 (N_6903,N_4436,N_3058);
and U6904 (N_6904,N_3235,N_3428);
nand U6905 (N_6905,N_4259,N_4857);
or U6906 (N_6906,N_2587,N_2792);
and U6907 (N_6907,N_2834,N_3885);
or U6908 (N_6908,N_4058,N_2808);
xnor U6909 (N_6909,N_3304,N_2650);
or U6910 (N_6910,N_3125,N_3505);
or U6911 (N_6911,N_3238,N_4071);
or U6912 (N_6912,N_3699,N_4834);
nor U6913 (N_6913,N_4135,N_3551);
xor U6914 (N_6914,N_3433,N_3638);
nor U6915 (N_6915,N_3872,N_2945);
nand U6916 (N_6916,N_3603,N_4194);
nor U6917 (N_6917,N_4604,N_4701);
xnor U6918 (N_6918,N_4419,N_3535);
or U6919 (N_6919,N_4398,N_4900);
nand U6920 (N_6920,N_3653,N_4171);
nor U6921 (N_6921,N_3666,N_4851);
nand U6922 (N_6922,N_4584,N_4370);
xor U6923 (N_6923,N_3639,N_3648);
xor U6924 (N_6924,N_2744,N_4894);
and U6925 (N_6925,N_4597,N_3184);
xor U6926 (N_6926,N_4318,N_4673);
nand U6927 (N_6927,N_3532,N_3006);
and U6928 (N_6928,N_2614,N_3079);
nand U6929 (N_6929,N_3489,N_2761);
or U6930 (N_6930,N_4285,N_3704);
xnor U6931 (N_6931,N_3792,N_3751);
and U6932 (N_6932,N_3155,N_2566);
or U6933 (N_6933,N_3318,N_4054);
or U6934 (N_6934,N_3010,N_2511);
xnor U6935 (N_6935,N_2531,N_3222);
xor U6936 (N_6936,N_2976,N_4193);
nand U6937 (N_6937,N_2629,N_3776);
nand U6938 (N_6938,N_2973,N_4956);
and U6939 (N_6939,N_4122,N_2769);
and U6940 (N_6940,N_2582,N_2905);
xnor U6941 (N_6941,N_4946,N_3813);
xnor U6942 (N_6942,N_3568,N_4529);
nand U6943 (N_6943,N_3696,N_4221);
nand U6944 (N_6944,N_4719,N_4464);
nor U6945 (N_6945,N_4662,N_3864);
and U6946 (N_6946,N_2822,N_3710);
nand U6947 (N_6947,N_4334,N_3575);
or U6948 (N_6948,N_3897,N_2912);
nor U6949 (N_6949,N_3480,N_4353);
or U6950 (N_6950,N_4249,N_3081);
and U6951 (N_6951,N_4452,N_4576);
nor U6952 (N_6952,N_3662,N_3074);
nand U6953 (N_6953,N_3144,N_4085);
and U6954 (N_6954,N_4036,N_4395);
and U6955 (N_6955,N_3621,N_3359);
xnor U6956 (N_6956,N_3196,N_3442);
nand U6957 (N_6957,N_3286,N_2950);
xnor U6958 (N_6958,N_3292,N_3669);
nor U6959 (N_6959,N_4426,N_3912);
nor U6960 (N_6960,N_4148,N_4106);
or U6961 (N_6961,N_3710,N_4190);
and U6962 (N_6962,N_3871,N_2714);
or U6963 (N_6963,N_4288,N_3388);
xnor U6964 (N_6964,N_3265,N_2675);
or U6965 (N_6965,N_2748,N_2707);
xnor U6966 (N_6966,N_2810,N_4092);
nor U6967 (N_6967,N_2748,N_3048);
nand U6968 (N_6968,N_4769,N_3612);
and U6969 (N_6969,N_2819,N_3967);
xor U6970 (N_6970,N_2662,N_2543);
nand U6971 (N_6971,N_4074,N_2794);
and U6972 (N_6972,N_2582,N_4212);
or U6973 (N_6973,N_3328,N_2811);
nor U6974 (N_6974,N_3512,N_3254);
and U6975 (N_6975,N_2961,N_2889);
nor U6976 (N_6976,N_2527,N_3256);
and U6977 (N_6977,N_4118,N_4906);
or U6978 (N_6978,N_4533,N_4129);
and U6979 (N_6979,N_4866,N_3875);
nor U6980 (N_6980,N_3631,N_3817);
or U6981 (N_6981,N_2713,N_2962);
and U6982 (N_6982,N_4217,N_2626);
and U6983 (N_6983,N_4375,N_3288);
xor U6984 (N_6984,N_4564,N_3321);
or U6985 (N_6985,N_2971,N_2531);
and U6986 (N_6986,N_3121,N_2852);
and U6987 (N_6987,N_3112,N_2826);
xor U6988 (N_6988,N_4291,N_4597);
nand U6989 (N_6989,N_4357,N_3897);
xor U6990 (N_6990,N_4770,N_3490);
or U6991 (N_6991,N_4566,N_2856);
nor U6992 (N_6992,N_2539,N_2682);
nor U6993 (N_6993,N_3360,N_4297);
nand U6994 (N_6994,N_3854,N_2969);
nor U6995 (N_6995,N_3835,N_4546);
xnor U6996 (N_6996,N_3887,N_3874);
nand U6997 (N_6997,N_4302,N_4884);
and U6998 (N_6998,N_3179,N_4276);
xnor U6999 (N_6999,N_3445,N_3052);
nor U7000 (N_7000,N_3582,N_4434);
and U7001 (N_7001,N_2984,N_3278);
nor U7002 (N_7002,N_2507,N_4690);
or U7003 (N_7003,N_3237,N_4081);
xor U7004 (N_7004,N_4326,N_3879);
nand U7005 (N_7005,N_2741,N_3903);
and U7006 (N_7006,N_3332,N_3862);
and U7007 (N_7007,N_2664,N_3911);
nor U7008 (N_7008,N_3771,N_4449);
nand U7009 (N_7009,N_4825,N_4907);
nor U7010 (N_7010,N_3462,N_3059);
or U7011 (N_7011,N_4657,N_3729);
and U7012 (N_7012,N_4811,N_4589);
nor U7013 (N_7013,N_4352,N_3333);
and U7014 (N_7014,N_3846,N_3918);
nand U7015 (N_7015,N_3543,N_3671);
xor U7016 (N_7016,N_2899,N_4665);
nand U7017 (N_7017,N_4861,N_4881);
nand U7018 (N_7018,N_3730,N_4745);
and U7019 (N_7019,N_4669,N_3179);
xnor U7020 (N_7020,N_2533,N_2809);
or U7021 (N_7021,N_3412,N_4766);
xor U7022 (N_7022,N_2574,N_4382);
nand U7023 (N_7023,N_2779,N_2544);
or U7024 (N_7024,N_3979,N_3574);
nand U7025 (N_7025,N_3019,N_4568);
nand U7026 (N_7026,N_4999,N_4479);
nand U7027 (N_7027,N_4578,N_3873);
and U7028 (N_7028,N_3647,N_3518);
nand U7029 (N_7029,N_4678,N_4001);
nor U7030 (N_7030,N_2860,N_2529);
xnor U7031 (N_7031,N_3744,N_4441);
or U7032 (N_7032,N_4860,N_4610);
and U7033 (N_7033,N_3963,N_4948);
xnor U7034 (N_7034,N_2526,N_2545);
xnor U7035 (N_7035,N_3887,N_4908);
and U7036 (N_7036,N_4818,N_4708);
or U7037 (N_7037,N_4918,N_4460);
xnor U7038 (N_7038,N_2568,N_4438);
nand U7039 (N_7039,N_4099,N_3183);
and U7040 (N_7040,N_4004,N_4193);
nand U7041 (N_7041,N_4716,N_3956);
or U7042 (N_7042,N_3488,N_4329);
or U7043 (N_7043,N_3231,N_4453);
nand U7044 (N_7044,N_4670,N_2865);
nor U7045 (N_7045,N_4120,N_2943);
nand U7046 (N_7046,N_4129,N_3436);
or U7047 (N_7047,N_2720,N_3198);
nor U7048 (N_7048,N_4258,N_4017);
nand U7049 (N_7049,N_2964,N_3659);
nor U7050 (N_7050,N_4075,N_4150);
or U7051 (N_7051,N_3391,N_4698);
xnor U7052 (N_7052,N_3552,N_4328);
nand U7053 (N_7053,N_2625,N_4029);
nor U7054 (N_7054,N_3209,N_3063);
nor U7055 (N_7055,N_2864,N_3309);
nand U7056 (N_7056,N_2569,N_4907);
xnor U7057 (N_7057,N_2572,N_3776);
nand U7058 (N_7058,N_3716,N_4122);
nor U7059 (N_7059,N_3618,N_3860);
or U7060 (N_7060,N_3364,N_4464);
xor U7061 (N_7061,N_3454,N_2990);
and U7062 (N_7062,N_4757,N_4605);
nand U7063 (N_7063,N_2545,N_4743);
xnor U7064 (N_7064,N_3449,N_3957);
xnor U7065 (N_7065,N_4727,N_3478);
and U7066 (N_7066,N_2954,N_3347);
nand U7067 (N_7067,N_3559,N_3008);
or U7068 (N_7068,N_4155,N_3969);
nor U7069 (N_7069,N_3890,N_3560);
nand U7070 (N_7070,N_3605,N_2655);
nand U7071 (N_7071,N_4988,N_4402);
or U7072 (N_7072,N_4613,N_4412);
nand U7073 (N_7073,N_2512,N_3323);
xor U7074 (N_7074,N_4215,N_3692);
nor U7075 (N_7075,N_3209,N_4097);
or U7076 (N_7076,N_2910,N_3959);
nor U7077 (N_7077,N_3463,N_3685);
nand U7078 (N_7078,N_2625,N_4424);
nor U7079 (N_7079,N_4890,N_2731);
and U7080 (N_7080,N_4339,N_3124);
or U7081 (N_7081,N_3273,N_3355);
or U7082 (N_7082,N_3152,N_3715);
and U7083 (N_7083,N_3361,N_3600);
or U7084 (N_7084,N_4505,N_3556);
nor U7085 (N_7085,N_2771,N_4340);
nand U7086 (N_7086,N_4469,N_2854);
or U7087 (N_7087,N_4809,N_3112);
xnor U7088 (N_7088,N_2652,N_3432);
nand U7089 (N_7089,N_3388,N_2761);
and U7090 (N_7090,N_3662,N_2785);
and U7091 (N_7091,N_3534,N_4239);
or U7092 (N_7092,N_3141,N_3648);
or U7093 (N_7093,N_3936,N_3491);
xnor U7094 (N_7094,N_2602,N_3120);
nand U7095 (N_7095,N_4330,N_3890);
xor U7096 (N_7096,N_2987,N_3229);
and U7097 (N_7097,N_4024,N_2508);
and U7098 (N_7098,N_3363,N_3510);
nor U7099 (N_7099,N_2567,N_3457);
or U7100 (N_7100,N_4762,N_3727);
nand U7101 (N_7101,N_2676,N_4284);
xor U7102 (N_7102,N_2797,N_3967);
xor U7103 (N_7103,N_3640,N_2769);
and U7104 (N_7104,N_3232,N_4491);
xnor U7105 (N_7105,N_3475,N_3720);
nand U7106 (N_7106,N_2867,N_4332);
nor U7107 (N_7107,N_3732,N_2549);
nor U7108 (N_7108,N_3971,N_3125);
nand U7109 (N_7109,N_4232,N_2710);
and U7110 (N_7110,N_3773,N_3760);
nor U7111 (N_7111,N_4347,N_3398);
nor U7112 (N_7112,N_2982,N_3575);
nand U7113 (N_7113,N_2632,N_3348);
nand U7114 (N_7114,N_2886,N_3248);
nand U7115 (N_7115,N_3814,N_3629);
xnor U7116 (N_7116,N_3150,N_3848);
nor U7117 (N_7117,N_3312,N_3567);
or U7118 (N_7118,N_3481,N_3469);
nand U7119 (N_7119,N_4857,N_3372);
and U7120 (N_7120,N_4392,N_2791);
and U7121 (N_7121,N_4096,N_2699);
and U7122 (N_7122,N_3379,N_4565);
nand U7123 (N_7123,N_3515,N_3617);
nor U7124 (N_7124,N_4108,N_4332);
nor U7125 (N_7125,N_2662,N_2866);
xor U7126 (N_7126,N_3006,N_2844);
and U7127 (N_7127,N_3564,N_2862);
xnor U7128 (N_7128,N_4307,N_2574);
nor U7129 (N_7129,N_3445,N_2595);
xor U7130 (N_7130,N_2787,N_4049);
and U7131 (N_7131,N_3025,N_4411);
xor U7132 (N_7132,N_4045,N_4541);
and U7133 (N_7133,N_3139,N_3655);
and U7134 (N_7134,N_4442,N_3755);
and U7135 (N_7135,N_4551,N_2872);
and U7136 (N_7136,N_4523,N_3560);
xnor U7137 (N_7137,N_3036,N_3390);
nand U7138 (N_7138,N_3017,N_2692);
nor U7139 (N_7139,N_3825,N_3033);
xor U7140 (N_7140,N_3741,N_4178);
xor U7141 (N_7141,N_4096,N_2628);
xor U7142 (N_7142,N_2610,N_3742);
nor U7143 (N_7143,N_3517,N_3359);
nand U7144 (N_7144,N_4691,N_2985);
nand U7145 (N_7145,N_4253,N_2696);
nand U7146 (N_7146,N_3958,N_4466);
nor U7147 (N_7147,N_4017,N_3685);
and U7148 (N_7148,N_2630,N_4699);
and U7149 (N_7149,N_3689,N_3345);
nand U7150 (N_7150,N_4165,N_4848);
and U7151 (N_7151,N_4513,N_4842);
nand U7152 (N_7152,N_3166,N_4901);
or U7153 (N_7153,N_2720,N_2944);
or U7154 (N_7154,N_3147,N_2909);
xor U7155 (N_7155,N_4129,N_3368);
nor U7156 (N_7156,N_4783,N_3015);
xnor U7157 (N_7157,N_3946,N_2774);
nand U7158 (N_7158,N_2732,N_3685);
nor U7159 (N_7159,N_4434,N_3409);
xor U7160 (N_7160,N_4969,N_4302);
nand U7161 (N_7161,N_4652,N_3328);
nor U7162 (N_7162,N_2651,N_4037);
nand U7163 (N_7163,N_3856,N_3106);
and U7164 (N_7164,N_3520,N_4614);
nand U7165 (N_7165,N_4341,N_3977);
or U7166 (N_7166,N_3927,N_3067);
nor U7167 (N_7167,N_4556,N_3555);
xor U7168 (N_7168,N_3061,N_4883);
and U7169 (N_7169,N_2995,N_3341);
nand U7170 (N_7170,N_4032,N_4344);
and U7171 (N_7171,N_2882,N_2942);
xnor U7172 (N_7172,N_3305,N_2931);
or U7173 (N_7173,N_4592,N_2611);
nand U7174 (N_7174,N_4729,N_2886);
or U7175 (N_7175,N_4547,N_2814);
or U7176 (N_7176,N_3560,N_2918);
and U7177 (N_7177,N_4585,N_3345);
and U7178 (N_7178,N_3518,N_4237);
nand U7179 (N_7179,N_4694,N_3628);
xor U7180 (N_7180,N_3582,N_3006);
nor U7181 (N_7181,N_4308,N_4408);
nor U7182 (N_7182,N_3018,N_2888);
xor U7183 (N_7183,N_4383,N_3292);
and U7184 (N_7184,N_4199,N_3330);
nor U7185 (N_7185,N_4274,N_3652);
nand U7186 (N_7186,N_4360,N_4564);
nand U7187 (N_7187,N_4467,N_3967);
and U7188 (N_7188,N_2963,N_4462);
or U7189 (N_7189,N_3238,N_2632);
or U7190 (N_7190,N_4992,N_4089);
nor U7191 (N_7191,N_3422,N_3170);
and U7192 (N_7192,N_4894,N_2823);
and U7193 (N_7193,N_2836,N_4143);
nand U7194 (N_7194,N_2756,N_3903);
and U7195 (N_7195,N_3824,N_4560);
or U7196 (N_7196,N_4551,N_4741);
nand U7197 (N_7197,N_4580,N_4482);
and U7198 (N_7198,N_3785,N_4020);
and U7199 (N_7199,N_4233,N_4727);
nor U7200 (N_7200,N_4132,N_4557);
and U7201 (N_7201,N_4785,N_4782);
and U7202 (N_7202,N_4176,N_3620);
or U7203 (N_7203,N_2625,N_4586);
or U7204 (N_7204,N_2543,N_2767);
nand U7205 (N_7205,N_3745,N_2523);
nand U7206 (N_7206,N_3548,N_4310);
xnor U7207 (N_7207,N_3175,N_4664);
and U7208 (N_7208,N_4131,N_4560);
nor U7209 (N_7209,N_3515,N_3847);
or U7210 (N_7210,N_4383,N_3353);
and U7211 (N_7211,N_4950,N_4972);
nand U7212 (N_7212,N_3906,N_2540);
and U7213 (N_7213,N_3335,N_3464);
xnor U7214 (N_7214,N_3472,N_4372);
xor U7215 (N_7215,N_4430,N_4214);
or U7216 (N_7216,N_3905,N_2942);
nand U7217 (N_7217,N_4273,N_4483);
xnor U7218 (N_7218,N_4463,N_4634);
nand U7219 (N_7219,N_2666,N_2703);
or U7220 (N_7220,N_4996,N_3340);
xor U7221 (N_7221,N_4652,N_4604);
xnor U7222 (N_7222,N_3148,N_4984);
nand U7223 (N_7223,N_4683,N_4904);
and U7224 (N_7224,N_3265,N_4958);
xnor U7225 (N_7225,N_4967,N_4847);
xor U7226 (N_7226,N_2661,N_3935);
xnor U7227 (N_7227,N_4804,N_2823);
nor U7228 (N_7228,N_4050,N_4345);
xor U7229 (N_7229,N_4530,N_4795);
or U7230 (N_7230,N_4571,N_4629);
and U7231 (N_7231,N_4226,N_3034);
or U7232 (N_7232,N_4806,N_4958);
and U7233 (N_7233,N_4284,N_3859);
nand U7234 (N_7234,N_2841,N_3248);
xnor U7235 (N_7235,N_4410,N_3389);
or U7236 (N_7236,N_3833,N_4075);
nor U7237 (N_7237,N_4335,N_2782);
and U7238 (N_7238,N_4068,N_4692);
nand U7239 (N_7239,N_3559,N_4773);
or U7240 (N_7240,N_4049,N_4800);
xor U7241 (N_7241,N_3224,N_4176);
nor U7242 (N_7242,N_2682,N_4389);
nand U7243 (N_7243,N_2636,N_3190);
xor U7244 (N_7244,N_2699,N_3594);
and U7245 (N_7245,N_4575,N_3263);
xor U7246 (N_7246,N_3232,N_3360);
nand U7247 (N_7247,N_4050,N_3081);
or U7248 (N_7248,N_4732,N_2623);
or U7249 (N_7249,N_2955,N_3254);
xnor U7250 (N_7250,N_4459,N_4487);
and U7251 (N_7251,N_3533,N_4240);
xor U7252 (N_7252,N_3584,N_3833);
or U7253 (N_7253,N_3562,N_3757);
and U7254 (N_7254,N_2519,N_2873);
nor U7255 (N_7255,N_4677,N_2779);
and U7256 (N_7256,N_2797,N_3859);
and U7257 (N_7257,N_3232,N_3591);
or U7258 (N_7258,N_4538,N_3344);
or U7259 (N_7259,N_3907,N_3140);
nand U7260 (N_7260,N_4205,N_4123);
nor U7261 (N_7261,N_4152,N_2603);
nor U7262 (N_7262,N_4802,N_3741);
xor U7263 (N_7263,N_4070,N_3495);
or U7264 (N_7264,N_4573,N_2754);
and U7265 (N_7265,N_3748,N_2980);
and U7266 (N_7266,N_4926,N_3056);
and U7267 (N_7267,N_2687,N_2579);
xor U7268 (N_7268,N_4461,N_4291);
xor U7269 (N_7269,N_3798,N_3073);
or U7270 (N_7270,N_4129,N_3627);
nor U7271 (N_7271,N_3868,N_3918);
nand U7272 (N_7272,N_4165,N_4339);
and U7273 (N_7273,N_4570,N_4652);
nand U7274 (N_7274,N_4430,N_2927);
xnor U7275 (N_7275,N_3199,N_4176);
nand U7276 (N_7276,N_4994,N_4639);
and U7277 (N_7277,N_4795,N_3565);
xnor U7278 (N_7278,N_4741,N_3785);
nand U7279 (N_7279,N_4232,N_2689);
xor U7280 (N_7280,N_4431,N_3043);
and U7281 (N_7281,N_3088,N_3742);
xor U7282 (N_7282,N_2822,N_4352);
nor U7283 (N_7283,N_4908,N_3978);
nor U7284 (N_7284,N_4019,N_3306);
xnor U7285 (N_7285,N_2798,N_2872);
nand U7286 (N_7286,N_3225,N_4079);
or U7287 (N_7287,N_2968,N_3585);
or U7288 (N_7288,N_3428,N_2620);
nor U7289 (N_7289,N_3723,N_3488);
xor U7290 (N_7290,N_3201,N_3562);
and U7291 (N_7291,N_3331,N_3813);
or U7292 (N_7292,N_3911,N_3675);
nand U7293 (N_7293,N_3623,N_4043);
and U7294 (N_7294,N_4594,N_3839);
or U7295 (N_7295,N_3219,N_3250);
xor U7296 (N_7296,N_4152,N_2723);
or U7297 (N_7297,N_4773,N_4485);
and U7298 (N_7298,N_3898,N_4854);
and U7299 (N_7299,N_3972,N_3535);
or U7300 (N_7300,N_4950,N_2678);
or U7301 (N_7301,N_3409,N_4506);
and U7302 (N_7302,N_2713,N_4807);
xor U7303 (N_7303,N_2807,N_3840);
or U7304 (N_7304,N_4628,N_2879);
nand U7305 (N_7305,N_4677,N_4872);
nor U7306 (N_7306,N_3974,N_3161);
nand U7307 (N_7307,N_2615,N_4539);
nand U7308 (N_7308,N_4674,N_3886);
or U7309 (N_7309,N_2680,N_4879);
or U7310 (N_7310,N_4421,N_4192);
and U7311 (N_7311,N_4487,N_3647);
and U7312 (N_7312,N_4442,N_2876);
and U7313 (N_7313,N_4122,N_3447);
and U7314 (N_7314,N_4000,N_3682);
or U7315 (N_7315,N_2995,N_3526);
nor U7316 (N_7316,N_3659,N_4003);
nor U7317 (N_7317,N_4315,N_4756);
and U7318 (N_7318,N_3203,N_2782);
nor U7319 (N_7319,N_2772,N_3484);
xor U7320 (N_7320,N_4516,N_4855);
xnor U7321 (N_7321,N_2690,N_4731);
and U7322 (N_7322,N_3835,N_4869);
nor U7323 (N_7323,N_2537,N_4189);
and U7324 (N_7324,N_2698,N_3028);
nor U7325 (N_7325,N_4168,N_3807);
nand U7326 (N_7326,N_4977,N_2885);
and U7327 (N_7327,N_3875,N_3529);
and U7328 (N_7328,N_4426,N_3293);
or U7329 (N_7329,N_3281,N_3301);
or U7330 (N_7330,N_4694,N_3594);
or U7331 (N_7331,N_4791,N_4460);
xor U7332 (N_7332,N_4768,N_3214);
and U7333 (N_7333,N_2793,N_2690);
nand U7334 (N_7334,N_4942,N_3354);
and U7335 (N_7335,N_3630,N_2865);
or U7336 (N_7336,N_4709,N_3836);
and U7337 (N_7337,N_4605,N_4361);
nand U7338 (N_7338,N_2716,N_4281);
and U7339 (N_7339,N_3816,N_3770);
nor U7340 (N_7340,N_3645,N_2773);
or U7341 (N_7341,N_4239,N_2992);
nand U7342 (N_7342,N_3354,N_3923);
nand U7343 (N_7343,N_2908,N_4942);
nor U7344 (N_7344,N_2944,N_4202);
or U7345 (N_7345,N_3094,N_3516);
nor U7346 (N_7346,N_3990,N_3474);
nor U7347 (N_7347,N_2883,N_2787);
nand U7348 (N_7348,N_3710,N_3598);
nand U7349 (N_7349,N_4100,N_2514);
nor U7350 (N_7350,N_2947,N_3343);
xor U7351 (N_7351,N_4884,N_4088);
and U7352 (N_7352,N_3126,N_3199);
nor U7353 (N_7353,N_2865,N_3093);
and U7354 (N_7354,N_3148,N_4576);
xnor U7355 (N_7355,N_3258,N_3555);
and U7356 (N_7356,N_2700,N_2799);
nand U7357 (N_7357,N_2662,N_3709);
xor U7358 (N_7358,N_3712,N_3665);
or U7359 (N_7359,N_4313,N_3219);
nand U7360 (N_7360,N_3655,N_3565);
or U7361 (N_7361,N_2830,N_2571);
nor U7362 (N_7362,N_2731,N_2770);
and U7363 (N_7363,N_3659,N_2766);
or U7364 (N_7364,N_4397,N_4206);
nand U7365 (N_7365,N_3091,N_4505);
and U7366 (N_7366,N_2992,N_4112);
nor U7367 (N_7367,N_4442,N_4827);
xnor U7368 (N_7368,N_3067,N_2630);
and U7369 (N_7369,N_3952,N_3313);
and U7370 (N_7370,N_4574,N_3832);
and U7371 (N_7371,N_2880,N_2769);
nand U7372 (N_7372,N_4275,N_3774);
and U7373 (N_7373,N_3795,N_4628);
or U7374 (N_7374,N_3693,N_2778);
nand U7375 (N_7375,N_4209,N_4866);
xor U7376 (N_7376,N_2776,N_3150);
or U7377 (N_7377,N_4590,N_3016);
or U7378 (N_7378,N_2749,N_4354);
or U7379 (N_7379,N_3503,N_3017);
and U7380 (N_7380,N_2765,N_3853);
nor U7381 (N_7381,N_3278,N_3111);
nor U7382 (N_7382,N_2589,N_4932);
or U7383 (N_7383,N_4465,N_3498);
nand U7384 (N_7384,N_4273,N_4963);
or U7385 (N_7385,N_3071,N_2948);
or U7386 (N_7386,N_3511,N_4409);
nand U7387 (N_7387,N_3680,N_4910);
xnor U7388 (N_7388,N_3406,N_3305);
and U7389 (N_7389,N_4293,N_3829);
nor U7390 (N_7390,N_4332,N_4546);
or U7391 (N_7391,N_3163,N_4651);
and U7392 (N_7392,N_4188,N_3731);
or U7393 (N_7393,N_3547,N_2773);
xnor U7394 (N_7394,N_3715,N_3910);
nor U7395 (N_7395,N_4152,N_2607);
nand U7396 (N_7396,N_4241,N_4350);
or U7397 (N_7397,N_3352,N_3491);
or U7398 (N_7398,N_4679,N_2996);
and U7399 (N_7399,N_4286,N_2687);
xnor U7400 (N_7400,N_2790,N_4907);
or U7401 (N_7401,N_3850,N_4836);
nor U7402 (N_7402,N_2620,N_4532);
nand U7403 (N_7403,N_4397,N_3184);
and U7404 (N_7404,N_3985,N_2637);
and U7405 (N_7405,N_4119,N_4185);
and U7406 (N_7406,N_4349,N_4880);
and U7407 (N_7407,N_4107,N_4977);
or U7408 (N_7408,N_2883,N_4423);
and U7409 (N_7409,N_4689,N_4384);
nor U7410 (N_7410,N_3665,N_3250);
or U7411 (N_7411,N_3174,N_3555);
or U7412 (N_7412,N_2823,N_4788);
xnor U7413 (N_7413,N_3464,N_4844);
and U7414 (N_7414,N_3502,N_2873);
or U7415 (N_7415,N_3621,N_4298);
and U7416 (N_7416,N_4574,N_2645);
nor U7417 (N_7417,N_3154,N_4904);
and U7418 (N_7418,N_4645,N_4279);
nand U7419 (N_7419,N_4121,N_2710);
or U7420 (N_7420,N_2629,N_3298);
xnor U7421 (N_7421,N_3486,N_3203);
or U7422 (N_7422,N_3565,N_3126);
nor U7423 (N_7423,N_3822,N_2895);
xor U7424 (N_7424,N_4307,N_4481);
or U7425 (N_7425,N_3664,N_4478);
nand U7426 (N_7426,N_4965,N_4658);
or U7427 (N_7427,N_4924,N_2704);
or U7428 (N_7428,N_3579,N_4022);
and U7429 (N_7429,N_3357,N_3879);
nor U7430 (N_7430,N_3787,N_4581);
and U7431 (N_7431,N_3930,N_3788);
or U7432 (N_7432,N_4931,N_3363);
nand U7433 (N_7433,N_4380,N_3792);
nor U7434 (N_7434,N_4500,N_2734);
nand U7435 (N_7435,N_2525,N_4833);
xor U7436 (N_7436,N_3703,N_4207);
and U7437 (N_7437,N_4864,N_3471);
or U7438 (N_7438,N_4685,N_2730);
nor U7439 (N_7439,N_2685,N_3679);
and U7440 (N_7440,N_4087,N_3275);
nor U7441 (N_7441,N_4356,N_4330);
or U7442 (N_7442,N_3200,N_3041);
and U7443 (N_7443,N_2811,N_3571);
nor U7444 (N_7444,N_4703,N_4010);
nand U7445 (N_7445,N_4884,N_4082);
nand U7446 (N_7446,N_3479,N_2928);
or U7447 (N_7447,N_3729,N_4505);
xnor U7448 (N_7448,N_4747,N_4370);
nand U7449 (N_7449,N_2710,N_4262);
and U7450 (N_7450,N_4299,N_3321);
or U7451 (N_7451,N_4099,N_3288);
and U7452 (N_7452,N_2791,N_4357);
nor U7453 (N_7453,N_3777,N_3913);
nor U7454 (N_7454,N_3741,N_3586);
nor U7455 (N_7455,N_4020,N_3408);
nor U7456 (N_7456,N_4792,N_4479);
or U7457 (N_7457,N_4223,N_3726);
nor U7458 (N_7458,N_4615,N_4477);
nand U7459 (N_7459,N_3681,N_2612);
nor U7460 (N_7460,N_3904,N_3580);
nand U7461 (N_7461,N_4162,N_2962);
nand U7462 (N_7462,N_2867,N_4200);
and U7463 (N_7463,N_2646,N_3401);
and U7464 (N_7464,N_2979,N_4548);
xnor U7465 (N_7465,N_3535,N_3933);
xor U7466 (N_7466,N_4557,N_2953);
nor U7467 (N_7467,N_3054,N_3383);
xnor U7468 (N_7468,N_3655,N_4863);
or U7469 (N_7469,N_3233,N_4261);
xnor U7470 (N_7470,N_4507,N_3875);
xor U7471 (N_7471,N_3519,N_4707);
or U7472 (N_7472,N_3514,N_2723);
and U7473 (N_7473,N_3112,N_2902);
nand U7474 (N_7474,N_4422,N_4556);
and U7475 (N_7475,N_4154,N_3312);
nand U7476 (N_7476,N_2649,N_4330);
and U7477 (N_7477,N_3780,N_2599);
nand U7478 (N_7478,N_3739,N_3986);
and U7479 (N_7479,N_3628,N_2835);
xnor U7480 (N_7480,N_4377,N_3845);
nor U7481 (N_7481,N_3361,N_3426);
xor U7482 (N_7482,N_3398,N_2574);
nand U7483 (N_7483,N_4912,N_3265);
nand U7484 (N_7484,N_4132,N_2711);
nor U7485 (N_7485,N_3136,N_2586);
nand U7486 (N_7486,N_4251,N_3310);
and U7487 (N_7487,N_3074,N_3036);
and U7488 (N_7488,N_4440,N_4823);
nand U7489 (N_7489,N_4758,N_3497);
nand U7490 (N_7490,N_3135,N_3563);
nand U7491 (N_7491,N_3194,N_4192);
nand U7492 (N_7492,N_4722,N_3890);
xor U7493 (N_7493,N_3857,N_4644);
xnor U7494 (N_7494,N_2738,N_3668);
and U7495 (N_7495,N_3460,N_4222);
nand U7496 (N_7496,N_3584,N_2842);
nand U7497 (N_7497,N_3832,N_3727);
nor U7498 (N_7498,N_3243,N_4262);
xnor U7499 (N_7499,N_3171,N_4895);
nand U7500 (N_7500,N_6396,N_5630);
or U7501 (N_7501,N_7218,N_7033);
xor U7502 (N_7502,N_6414,N_6348);
nor U7503 (N_7503,N_5719,N_5832);
xnor U7504 (N_7504,N_5212,N_5107);
xnor U7505 (N_7505,N_7191,N_6022);
xor U7506 (N_7506,N_6755,N_5290);
nor U7507 (N_7507,N_6175,N_6633);
xnor U7508 (N_7508,N_6247,N_5369);
nand U7509 (N_7509,N_6248,N_5269);
xor U7510 (N_7510,N_7392,N_6651);
nand U7511 (N_7511,N_7436,N_6098);
or U7512 (N_7512,N_6983,N_7018);
and U7513 (N_7513,N_6603,N_5318);
xor U7514 (N_7514,N_6044,N_5240);
xnor U7515 (N_7515,N_5271,N_6899);
or U7516 (N_7516,N_7421,N_7031);
nor U7517 (N_7517,N_7341,N_7256);
xor U7518 (N_7518,N_5262,N_6205);
nand U7519 (N_7519,N_7270,N_6407);
nor U7520 (N_7520,N_7054,N_5396);
or U7521 (N_7521,N_5078,N_5321);
nand U7522 (N_7522,N_6187,N_5169);
nor U7523 (N_7523,N_7339,N_5513);
and U7524 (N_7524,N_6274,N_5468);
nor U7525 (N_7525,N_7344,N_6455);
or U7526 (N_7526,N_5586,N_6498);
and U7527 (N_7527,N_6086,N_6554);
and U7528 (N_7528,N_6087,N_7350);
xnor U7529 (N_7529,N_7426,N_6890);
xor U7530 (N_7530,N_6871,N_6045);
and U7531 (N_7531,N_7412,N_6174);
or U7532 (N_7532,N_5579,N_5608);
nand U7533 (N_7533,N_6138,N_7065);
and U7534 (N_7534,N_5744,N_5139);
and U7535 (N_7535,N_6611,N_5814);
or U7536 (N_7536,N_6847,N_6924);
nor U7537 (N_7537,N_6125,N_6804);
or U7538 (N_7538,N_5418,N_6851);
and U7539 (N_7539,N_5201,N_5100);
xnor U7540 (N_7540,N_5215,N_6552);
or U7541 (N_7541,N_6089,N_7414);
and U7542 (N_7542,N_6178,N_5527);
xnor U7543 (N_7543,N_5255,N_6506);
and U7544 (N_7544,N_6989,N_6723);
nand U7545 (N_7545,N_7014,N_5748);
or U7546 (N_7546,N_6293,N_6562);
nand U7547 (N_7547,N_5532,N_5802);
and U7548 (N_7548,N_7021,N_5297);
xor U7549 (N_7549,N_6164,N_5788);
xnor U7550 (N_7550,N_5642,N_5299);
and U7551 (N_7551,N_6672,N_5181);
xnor U7552 (N_7552,N_7486,N_6673);
and U7553 (N_7553,N_5680,N_7429);
nor U7554 (N_7554,N_6535,N_6432);
nand U7555 (N_7555,N_5146,N_6226);
nor U7556 (N_7556,N_5202,N_5332);
and U7557 (N_7557,N_5003,N_7290);
or U7558 (N_7558,N_6343,N_5599);
and U7559 (N_7559,N_6967,N_7069);
xnor U7560 (N_7560,N_6970,N_6576);
or U7561 (N_7561,N_6757,N_6258);
and U7562 (N_7562,N_7485,N_6306);
and U7563 (N_7563,N_7255,N_7276);
and U7564 (N_7564,N_6849,N_5300);
or U7565 (N_7565,N_7376,N_5660);
and U7566 (N_7566,N_5618,N_5995);
nor U7567 (N_7567,N_6077,N_7219);
and U7568 (N_7568,N_6259,N_5307);
nor U7569 (N_7569,N_6331,N_5339);
or U7570 (N_7570,N_6663,N_7390);
xnor U7571 (N_7571,N_6588,N_7280);
or U7572 (N_7572,N_6634,N_6386);
nor U7573 (N_7573,N_7230,N_5090);
or U7574 (N_7574,N_5973,N_7000);
and U7575 (N_7575,N_6971,N_6763);
nand U7576 (N_7576,N_6124,N_5913);
nand U7577 (N_7577,N_7292,N_7066);
xor U7578 (N_7578,N_7316,N_5303);
xor U7579 (N_7579,N_7407,N_5759);
nand U7580 (N_7580,N_7441,N_5121);
xor U7581 (N_7581,N_5356,N_5780);
and U7582 (N_7582,N_6915,N_6188);
and U7583 (N_7583,N_6350,N_5947);
xnor U7584 (N_7584,N_6228,N_6660);
and U7585 (N_7585,N_6405,N_6788);
xnor U7586 (N_7586,N_7439,N_6625);
and U7587 (N_7587,N_7460,N_6520);
and U7588 (N_7588,N_5977,N_7360);
nor U7589 (N_7589,N_6406,N_5923);
xor U7590 (N_7590,N_5274,N_6469);
and U7591 (N_7591,N_7184,N_5849);
nor U7592 (N_7592,N_6713,N_6497);
xnor U7593 (N_7593,N_7196,N_6691);
and U7594 (N_7594,N_5985,N_6215);
nand U7595 (N_7595,N_6919,N_5399);
or U7596 (N_7596,N_5187,N_6627);
xnor U7597 (N_7597,N_6281,N_5697);
nand U7598 (N_7598,N_6769,N_7487);
or U7599 (N_7599,N_5053,N_6093);
nand U7600 (N_7600,N_6954,N_5058);
xor U7601 (N_7601,N_6993,N_5460);
nor U7602 (N_7602,N_7268,N_7083);
and U7603 (N_7603,N_6756,N_5316);
xnor U7604 (N_7604,N_6901,N_5874);
nor U7605 (N_7605,N_6369,N_5253);
nand U7606 (N_7606,N_6282,N_7176);
and U7607 (N_7607,N_6973,N_6298);
or U7608 (N_7608,N_7101,N_6523);
nand U7609 (N_7609,N_5196,N_6488);
and U7610 (N_7610,N_5441,N_5232);
nand U7611 (N_7611,N_5024,N_5711);
or U7612 (N_7612,N_6329,N_6473);
xnor U7613 (N_7613,N_7100,N_5745);
nor U7614 (N_7614,N_6068,N_5669);
xor U7615 (N_7615,N_5508,N_6917);
nor U7616 (N_7616,N_5077,N_7165);
nor U7617 (N_7617,N_7062,N_5765);
nand U7618 (N_7618,N_6796,N_6856);
nand U7619 (N_7619,N_5519,N_5693);
xnor U7620 (N_7620,N_6922,N_5192);
and U7621 (N_7621,N_5151,N_6207);
and U7622 (N_7622,N_5084,N_5966);
and U7623 (N_7623,N_5521,N_5329);
xor U7624 (N_7624,N_7343,N_6938);
xor U7625 (N_7625,N_5541,N_5524);
and U7626 (N_7626,N_5328,N_6083);
or U7627 (N_7627,N_6511,N_6979);
and U7628 (N_7628,N_6618,N_6302);
nor U7629 (N_7629,N_6269,N_6674);
nor U7630 (N_7630,N_6736,N_7384);
nor U7631 (N_7631,N_6437,N_5291);
nor U7632 (N_7632,N_6877,N_6430);
and U7633 (N_7633,N_5739,N_7375);
nand U7634 (N_7634,N_7297,N_5395);
xnor U7635 (N_7635,N_7144,N_6773);
or U7636 (N_7636,N_7468,N_7313);
or U7637 (N_7637,N_5904,N_7007);
and U7638 (N_7638,N_5185,N_6819);
nand U7639 (N_7639,N_7351,N_5437);
or U7640 (N_7640,N_5135,N_5234);
xnor U7641 (N_7641,N_7329,N_5920);
or U7642 (N_7642,N_6664,N_5406);
or U7643 (N_7643,N_5847,N_6047);
nand U7644 (N_7644,N_6295,N_5052);
nand U7645 (N_7645,N_6156,N_7396);
nor U7646 (N_7646,N_5674,N_7078);
and U7647 (N_7647,N_5726,N_6012);
xnor U7648 (N_7648,N_6799,N_6649);
nor U7649 (N_7649,N_5790,N_5081);
nand U7650 (N_7650,N_7273,N_6404);
and U7651 (N_7651,N_5256,N_6793);
xor U7652 (N_7652,N_5403,N_6777);
and U7653 (N_7653,N_6075,N_6543);
or U7654 (N_7654,N_7499,N_5310);
nand U7655 (N_7655,N_5286,N_6900);
nor U7656 (N_7656,N_5385,N_6969);
nor U7657 (N_7657,N_5818,N_7148);
or U7658 (N_7658,N_6885,N_6040);
and U7659 (N_7659,N_6252,N_5701);
or U7660 (N_7660,N_5322,N_7135);
nand U7661 (N_7661,N_7027,N_5806);
or U7662 (N_7662,N_6061,N_6861);
xor U7663 (N_7663,N_5311,N_5512);
nor U7664 (N_7664,N_7498,N_7393);
and U7665 (N_7665,N_5844,N_5800);
nand U7666 (N_7666,N_5917,N_5029);
or U7667 (N_7667,N_6452,N_6641);
or U7668 (N_7668,N_5881,N_6335);
and U7669 (N_7669,N_5539,N_7364);
nor U7670 (N_7670,N_5485,N_7042);
xnor U7671 (N_7671,N_7115,N_5091);
nor U7672 (N_7672,N_6795,N_7046);
nand U7673 (N_7673,N_6460,N_5893);
nand U7674 (N_7674,N_5099,N_6671);
xor U7675 (N_7675,N_6710,N_5775);
or U7676 (N_7676,N_6719,N_5771);
or U7677 (N_7677,N_5547,N_6525);
nand U7678 (N_7678,N_6734,N_6581);
nand U7679 (N_7679,N_7377,N_5622);
or U7680 (N_7680,N_6132,N_6942);
or U7681 (N_7681,N_5333,N_6374);
xnor U7682 (N_7682,N_6017,N_6037);
and U7683 (N_7683,N_6578,N_6679);
nand U7684 (N_7684,N_6830,N_5360);
xnor U7685 (N_7685,N_5469,N_6166);
nand U7686 (N_7686,N_6524,N_5837);
nor U7687 (N_7687,N_6167,N_5383);
xor U7688 (N_7688,N_6957,N_6470);
xor U7689 (N_7689,N_5969,N_5643);
and U7690 (N_7690,N_6112,N_5921);
nand U7691 (N_7691,N_5301,N_7087);
and U7692 (N_7692,N_6889,N_7013);
nor U7693 (N_7693,N_5016,N_6333);
and U7694 (N_7694,N_5857,N_6449);
xor U7695 (N_7695,N_6242,N_6682);
nand U7696 (N_7696,N_7310,N_5431);
xnor U7697 (N_7697,N_6308,N_5955);
xor U7698 (N_7698,N_6782,N_5685);
nor U7699 (N_7699,N_5117,N_5293);
nand U7700 (N_7700,N_5561,N_6468);
or U7701 (N_7701,N_5621,N_5027);
or U7702 (N_7702,N_5957,N_5227);
nand U7703 (N_7703,N_6531,N_7286);
or U7704 (N_7704,N_6192,N_5294);
or U7705 (N_7705,N_5530,N_5822);
and U7706 (N_7706,N_5902,N_7397);
xnor U7707 (N_7707,N_6786,N_7475);
and U7708 (N_7708,N_5639,N_5043);
nor U7709 (N_7709,N_5342,N_7402);
and U7710 (N_7710,N_5900,N_6024);
nor U7711 (N_7711,N_6031,N_5309);
nor U7712 (N_7712,N_6873,N_5390);
nand U7713 (N_7713,N_5148,N_6408);
and U7714 (N_7714,N_5026,N_6324);
xor U7715 (N_7715,N_6735,N_7444);
and U7716 (N_7716,N_5807,N_5064);
nand U7717 (N_7717,N_7025,N_6244);
and U7718 (N_7718,N_6872,N_6920);
nand U7719 (N_7719,N_6463,N_7370);
nor U7720 (N_7720,N_7369,N_5025);
xor U7721 (N_7721,N_5594,N_7020);
nand U7722 (N_7722,N_5125,N_7012);
nor U7723 (N_7723,N_7045,N_5533);
xor U7724 (N_7724,N_5838,N_5314);
xor U7725 (N_7725,N_6139,N_6182);
xor U7726 (N_7726,N_6714,N_6314);
nor U7727 (N_7727,N_6076,N_5796);
or U7728 (N_7728,N_6262,N_7466);
or U7729 (N_7729,N_6636,N_7259);
nand U7730 (N_7730,N_5828,N_7404);
and U7731 (N_7731,N_6709,N_5129);
xnor U7732 (N_7732,N_5762,N_6426);
nand U7733 (N_7733,N_6398,N_5631);
or U7734 (N_7734,N_7332,N_7432);
and U7735 (N_7735,N_5896,N_6360);
or U7736 (N_7736,N_6540,N_5854);
xnor U7737 (N_7737,N_7431,N_5470);
nor U7738 (N_7738,N_5895,N_7320);
nor U7739 (N_7739,N_5228,N_7422);
or U7740 (N_7740,N_6812,N_6276);
xor U7741 (N_7741,N_6655,N_7328);
xor U7742 (N_7742,N_5872,N_7388);
nor U7743 (N_7743,N_5157,N_7401);
xnor U7744 (N_7744,N_5059,N_6949);
xnor U7745 (N_7745,N_6322,N_5218);
nand U7746 (N_7746,N_5067,N_7494);
or U7747 (N_7747,N_6632,N_5382);
or U7748 (N_7748,N_5747,N_6561);
xor U7749 (N_7749,N_5836,N_6806);
xor U7750 (N_7750,N_7127,N_5794);
and U7751 (N_7751,N_5248,N_5563);
nor U7752 (N_7752,N_5213,N_6121);
nand U7753 (N_7753,N_7278,N_6260);
or U7754 (N_7754,N_6574,N_5263);
or U7755 (N_7755,N_6436,N_5420);
and U7756 (N_7756,N_5946,N_5555);
xor U7757 (N_7757,N_6312,N_7039);
or U7758 (N_7758,N_7423,N_7052);
nand U7759 (N_7759,N_7124,N_7009);
nor U7760 (N_7760,N_5753,N_6229);
and U7761 (N_7761,N_6370,N_6748);
nor U7762 (N_7762,N_5534,N_5720);
or U7763 (N_7763,N_6791,N_5104);
xnor U7764 (N_7764,N_7079,N_7128);
nor U7765 (N_7765,N_5149,N_5761);
nand U7766 (N_7766,N_5199,N_5931);
nand U7767 (N_7767,N_7257,N_5503);
xnor U7768 (N_7768,N_7269,N_6986);
nand U7769 (N_7769,N_5646,N_7208);
nand U7770 (N_7770,N_6648,N_7231);
nor U7771 (N_7771,N_6261,N_7195);
xnor U7772 (N_7772,N_6662,N_5672);
nand U7773 (N_7773,N_7489,N_7373);
and U7774 (N_7774,N_6557,N_6150);
or U7775 (N_7775,N_6238,N_6462);
or U7776 (N_7776,N_6771,N_6256);
nor U7777 (N_7777,N_6162,N_5225);
nor U7778 (N_7778,N_5401,N_6667);
or U7779 (N_7779,N_5051,N_6959);
and U7780 (N_7780,N_5284,N_6071);
and U7781 (N_7781,N_6034,N_7188);
nand U7782 (N_7782,N_5531,N_7185);
xor U7783 (N_7783,N_6213,N_6009);
and U7784 (N_7784,N_7178,N_6292);
or U7785 (N_7785,N_5862,N_7319);
or U7786 (N_7786,N_5171,N_5178);
and U7787 (N_7787,N_7482,N_6113);
or U7788 (N_7788,N_6568,N_7287);
or U7789 (N_7789,N_6070,N_5689);
or U7790 (N_7790,N_7266,N_6555);
nor U7791 (N_7791,N_5658,N_7203);
xor U7792 (N_7792,N_5289,N_6999);
xor U7793 (N_7793,N_5870,N_5159);
xor U7794 (N_7794,N_5486,N_6008);
xnor U7795 (N_7795,N_6443,N_6698);
and U7796 (N_7796,N_7177,N_7312);
nand U7797 (N_7797,N_5118,N_5455);
or U7798 (N_7798,N_6413,N_5194);
nand U7799 (N_7799,N_7092,N_6066);
nor U7800 (N_7800,N_5557,N_7238);
and U7801 (N_7801,N_6442,N_5951);
and U7802 (N_7802,N_5548,N_5821);
nand U7803 (N_7803,N_5770,N_6088);
xnor U7804 (N_7804,N_6879,N_6878);
and U7805 (N_7805,N_6082,N_7112);
nor U7806 (N_7806,N_7153,N_6895);
nor U7807 (N_7807,N_5734,N_6645);
or U7808 (N_7808,N_6201,N_5368);
nor U7809 (N_7809,N_6489,N_5281);
and U7810 (N_7810,N_7035,N_6265);
nand U7811 (N_7811,N_7157,N_6241);
or U7812 (N_7812,N_5852,N_7113);
nand U7813 (N_7813,N_7116,N_5145);
xnor U7814 (N_7814,N_6685,N_6270);
xor U7815 (N_7815,N_5285,N_7438);
or U7816 (N_7816,N_6703,N_6422);
or U7817 (N_7817,N_6392,N_5376);
nor U7818 (N_7818,N_7451,N_5447);
xnor U7819 (N_7819,N_7399,N_5959);
nor U7820 (N_7820,N_5371,N_6433);
and U7821 (N_7821,N_6445,N_7166);
and U7822 (N_7822,N_5730,N_6490);
xnor U7823 (N_7823,N_7132,N_7228);
nor U7824 (N_7824,N_5999,N_5438);
nor U7825 (N_7825,N_5699,N_5002);
nor U7826 (N_7826,N_7200,N_5233);
or U7827 (N_7827,N_5186,N_7222);
nand U7828 (N_7828,N_5141,N_6958);
xnor U7829 (N_7829,N_5098,N_6021);
or U7830 (N_7830,N_6079,N_5476);
nand U7831 (N_7831,N_5927,N_6760);
and U7832 (N_7832,N_5130,N_5976);
xnor U7833 (N_7833,N_6728,N_7197);
nor U7834 (N_7834,N_5175,N_5166);
and U7835 (N_7835,N_6739,N_7336);
or U7836 (N_7836,N_5477,N_5434);
nor U7837 (N_7837,N_5811,N_5915);
or U7838 (N_7838,N_5163,N_5123);
nand U7839 (N_7839,N_7029,N_6754);
and U7840 (N_7840,N_5464,N_7194);
xor U7841 (N_7841,N_6368,N_6943);
or U7842 (N_7842,N_7248,N_6690);
or U7843 (N_7843,N_7325,N_5683);
nor U7844 (N_7844,N_5695,N_5848);
and U7845 (N_7845,N_6095,N_6286);
and U7846 (N_7846,N_6599,N_6509);
or U7847 (N_7847,N_7317,N_5346);
nand U7848 (N_7848,N_7235,N_6519);
xnor U7849 (N_7849,N_7352,N_5668);
and U7850 (N_7850,N_6517,N_5535);
nand U7851 (N_7851,N_7395,N_5188);
or U7852 (N_7852,N_5176,N_7229);
nand U7853 (N_7853,N_5808,N_5334);
nand U7854 (N_7854,N_6859,N_5056);
xnor U7855 (N_7855,N_6179,N_7213);
nand U7856 (N_7856,N_5357,N_5912);
or U7857 (N_7857,N_6807,N_6152);
or U7858 (N_7858,N_5882,N_5605);
or U7859 (N_7859,N_7064,N_5840);
and U7860 (N_7860,N_6956,N_5010);
nor U7861 (N_7861,N_6834,N_6571);
or U7862 (N_7862,N_5238,N_7374);
and U7863 (N_7863,N_6210,N_6668);
nand U7864 (N_7864,N_7050,N_6237);
nand U7865 (N_7865,N_6953,N_5978);
or U7866 (N_7866,N_5568,N_5742);
or U7867 (N_7867,N_5362,N_5088);
xnor U7868 (N_7868,N_6518,N_5868);
nor U7869 (N_7869,N_6028,N_5787);
nand U7870 (N_7870,N_5974,N_7179);
or U7871 (N_7871,N_6458,N_7005);
or U7872 (N_7872,N_5195,N_5222);
nor U7873 (N_7873,N_7417,N_6380);
or U7874 (N_7874,N_5861,N_5189);
and U7875 (N_7875,N_5173,N_5466);
nor U7876 (N_7876,N_5552,N_6765);
nor U7877 (N_7877,N_6450,N_5700);
or U7878 (N_7878,N_7207,N_7056);
nor U7879 (N_7879,N_7187,N_5839);
nand U7880 (N_7880,N_6802,N_5254);
nor U7881 (N_7881,N_5797,N_5292);
xor U7882 (N_7882,N_6065,N_7085);
and U7883 (N_7883,N_6078,N_5860);
nand U7884 (N_7884,N_5217,N_7097);
or U7885 (N_7885,N_7372,N_6389);
and U7886 (N_7886,N_6310,N_5649);
xor U7887 (N_7887,N_5393,N_5465);
nor U7888 (N_7888,N_6440,N_6832);
and U7889 (N_7889,N_7470,N_5877);
nor U7890 (N_7890,N_6505,N_5721);
nor U7891 (N_7891,N_5692,N_6512);
nor U7892 (N_7892,N_6816,N_7129);
xnor U7893 (N_7893,N_6052,N_5352);
and U7894 (N_7894,N_7289,N_7354);
or U7895 (N_7895,N_7496,N_6400);
nor U7896 (N_7896,N_5150,N_7300);
nor U7897 (N_7897,N_6912,N_6043);
xnor U7898 (N_7898,N_5691,N_5735);
xor U7899 (N_7899,N_6136,N_5277);
xor U7900 (N_7900,N_6246,N_6173);
and U7901 (N_7901,N_7347,N_5331);
or U7902 (N_7902,N_5161,N_7419);
nand U7903 (N_7903,N_5374,N_7059);
or U7904 (N_7904,N_6332,N_6199);
xnor U7905 (N_7905,N_5496,N_5990);
xnor U7906 (N_7906,N_7149,N_7398);
nor U7907 (N_7907,N_7241,N_5597);
or U7908 (N_7908,N_6344,N_6172);
nor U7909 (N_7909,N_5950,N_5994);
nand U7910 (N_7910,N_5423,N_5515);
nor U7911 (N_7911,N_7172,N_7081);
nor U7912 (N_7912,N_6251,N_6937);
xnor U7913 (N_7913,N_6996,N_6813);
or U7914 (N_7914,N_6930,N_5778);
nor U7915 (N_7915,N_7283,N_5510);
or U7916 (N_7916,N_5389,N_5174);
xnor U7917 (N_7917,N_6725,N_5180);
xnor U7918 (N_7918,N_6821,N_7483);
xnor U7919 (N_7919,N_5115,N_5542);
xor U7920 (N_7920,N_7359,N_6094);
and U7921 (N_7921,N_5598,N_5204);
or U7922 (N_7922,N_5706,N_6475);
xor U7923 (N_7923,N_6140,N_6410);
xor U7924 (N_7924,N_6542,N_6023);
and U7925 (N_7925,N_6250,N_5155);
xnor U7926 (N_7926,N_5550,N_6421);
and U7927 (N_7927,N_7051,N_5591);
and U7928 (N_7928,N_6472,N_6610);
nor U7929 (N_7929,N_5624,N_5670);
or U7930 (N_7930,N_6510,N_6533);
nor U7931 (N_7931,N_5036,N_6701);
nand U7932 (N_7932,N_7002,N_7220);
nor U7933 (N_7933,N_5656,N_5219);
nor U7934 (N_7934,N_5428,N_6235);
nand U7935 (N_7935,N_5940,N_6290);
xor U7936 (N_7936,N_5268,N_5914);
and U7937 (N_7937,N_7293,N_6184);
and U7938 (N_7938,N_5566,N_5640);
nand U7939 (N_7939,N_5251,N_5086);
nor U7940 (N_7940,N_5791,N_5714);
or U7941 (N_7941,N_7413,N_7173);
xor U7942 (N_7942,N_7418,N_5493);
nor U7943 (N_7943,N_6624,N_5784);
or U7944 (N_7944,N_6595,N_6305);
or U7945 (N_7945,N_6761,N_6415);
and U7946 (N_7946,N_6319,N_7119);
xnor U7947 (N_7947,N_5214,N_6619);
nand U7948 (N_7948,N_6666,N_7380);
and U7949 (N_7949,N_6976,N_6397);
nor U7950 (N_7950,N_5878,N_6459);
nor U7951 (N_7951,N_5997,N_7102);
nor U7952 (N_7952,N_5184,N_5338);
and U7953 (N_7953,N_6170,N_6808);
nor U7954 (N_7954,N_5386,N_6658);
nand U7955 (N_7955,N_6020,N_7453);
nand U7956 (N_7956,N_7348,N_7281);
or U7957 (N_7957,N_6965,N_6684);
nand U7958 (N_7958,N_7333,N_6338);
nand U7959 (N_7959,N_6977,N_7314);
and U7960 (N_7960,N_6352,N_5588);
or U7961 (N_7961,N_5952,N_5815);
nor U7962 (N_7962,N_5731,N_6620);
and U7963 (N_7963,N_5035,N_5230);
or U7964 (N_7964,N_7058,N_5265);
nor U7965 (N_7965,N_6718,N_5417);
and U7966 (N_7966,N_5340,N_5305);
nand U7967 (N_7967,N_6893,N_5267);
and U7968 (N_7968,N_5725,N_7201);
nor U7969 (N_7969,N_7488,N_5752);
or U7970 (N_7970,N_5210,N_6740);
and U7971 (N_7971,N_6990,N_5020);
nand U7972 (N_7972,N_7169,N_7038);
nand U7973 (N_7973,N_7143,N_6746);
nor U7974 (N_7974,N_7435,N_6950);
xor U7975 (N_7975,N_6747,N_5671);
xor U7976 (N_7976,N_7240,N_7226);
xnor U7977 (N_7977,N_6361,N_6377);
nand U7978 (N_7978,N_5006,N_5391);
xor U7979 (N_7979,N_6128,N_7246);
or U7980 (N_7980,N_6069,N_6732);
nand U7981 (N_7981,N_7041,N_5687);
xnor U7982 (N_7982,N_6120,N_5907);
nor U7983 (N_7983,N_5526,N_5461);
and U7984 (N_7984,N_5954,N_5569);
nand U7985 (N_7985,N_5453,N_5205);
or U7986 (N_7986,N_5520,N_7049);
and U7987 (N_7987,N_6161,N_6145);
xnor U7988 (N_7988,N_5074,N_5678);
nand U7989 (N_7989,N_5867,N_6067);
and U7990 (N_7990,N_7362,N_6054);
xor U7991 (N_7991,N_5992,N_5536);
nor U7992 (N_7992,N_6716,N_6750);
nand U7993 (N_7993,N_5509,N_5686);
nor U7994 (N_7994,N_7474,N_6617);
or U7995 (N_7995,N_5160,N_5375);
nand U7996 (N_7996,N_5667,N_5087);
nand U7997 (N_7997,N_6863,N_6257);
nand U7998 (N_7998,N_6592,N_5905);
nor U7999 (N_7999,N_6598,N_7309);
nand U8000 (N_8000,N_6211,N_5756);
nand U8001 (N_8001,N_5040,N_6018);
nor U8002 (N_8002,N_6853,N_5203);
nand U8003 (N_8003,N_7326,N_6081);
and U8004 (N_8004,N_5810,N_5529);
or U8005 (N_8005,N_7133,N_7409);
and U8006 (N_8006,N_6902,N_7275);
or U8007 (N_8007,N_7342,N_6538);
nand U8008 (N_8008,N_5945,N_5249);
xor U8009 (N_8009,N_7299,N_5366);
nor U8010 (N_8010,N_6330,N_6232);
and U8011 (N_8011,N_5168,N_5799);
or U8012 (N_8012,N_7428,N_5774);
xnor U8013 (N_8013,N_5073,N_5381);
xor U8014 (N_8014,N_5645,N_7136);
and U8015 (N_8015,N_7096,N_5302);
xor U8016 (N_8016,N_6142,N_6219);
and U8017 (N_8017,N_6850,N_5257);
or U8018 (N_8018,N_7331,N_6590);
xnor U8019 (N_8019,N_5908,N_5517);
and U8020 (N_8020,N_5892,N_7182);
nor U8021 (N_8021,N_7458,N_5120);
or U8022 (N_8022,N_6159,N_7199);
and U8023 (N_8023,N_5103,N_6457);
nor U8024 (N_8024,N_5738,N_5728);
or U8025 (N_8025,N_6704,N_6029);
nand U8026 (N_8026,N_6579,N_5873);
nor U8027 (N_8027,N_6465,N_6194);
nand U8028 (N_8028,N_6321,N_6340);
nor U8029 (N_8029,N_6461,N_6134);
nand U8030 (N_8030,N_7094,N_6016);
xnor U8031 (N_8031,N_5850,N_6809);
nor U8032 (N_8032,N_7424,N_5272);
and U8033 (N_8033,N_6820,N_5456);
or U8034 (N_8034,N_6656,N_6558);
and U8035 (N_8035,N_6615,N_7443);
nand U8036 (N_8036,N_5275,N_7137);
xor U8037 (N_8037,N_5859,N_5936);
and U8038 (N_8038,N_6263,N_6749);
or U8039 (N_8039,N_5540,N_7303);
nand U8040 (N_8040,N_6946,N_6130);
nand U8041 (N_8041,N_6264,N_5712);
or U8042 (N_8042,N_5518,N_6288);
xor U8043 (N_8043,N_7110,N_5446);
nand U8044 (N_8044,N_7104,N_5785);
nand U8045 (N_8045,N_5682,N_5610);
or U8046 (N_8046,N_7106,N_5948);
and U8047 (N_8047,N_6032,N_6589);
nor U8048 (N_8048,N_5266,N_6526);
xnor U8049 (N_8049,N_7252,N_5988);
or U8050 (N_8050,N_6823,N_7415);
and U8051 (N_8051,N_6700,N_6677);
or U8052 (N_8052,N_7335,N_5154);
nand U8053 (N_8053,N_7337,N_7334);
xor U8054 (N_8054,N_6438,N_7430);
and U8055 (N_8055,N_7215,N_5235);
or U8056 (N_8056,N_5938,N_7311);
and U8057 (N_8057,N_6657,N_7154);
nor U8058 (N_8058,N_5191,N_7473);
or U8059 (N_8059,N_6939,N_6100);
nor U8060 (N_8060,N_6935,N_5538);
xnor U8061 (N_8061,N_5336,N_6351);
nand U8062 (N_8062,N_5282,N_6854);
nor U8063 (N_8063,N_6284,N_6243);
and U8064 (N_8064,N_5004,N_6391);
and U8065 (N_8065,N_7262,N_7077);
or U8066 (N_8066,N_6060,N_6474);
nand U8067 (N_8067,N_6171,N_7449);
or U8068 (N_8068,N_6865,N_7161);
xnor U8069 (N_8069,N_5443,N_6266);
xnor U8070 (N_8070,N_5324,N_5260);
or U8071 (N_8071,N_7295,N_6584);
or U8072 (N_8072,N_6737,N_7202);
nand U8073 (N_8073,N_7138,N_5351);
and U8074 (N_8074,N_5312,N_5582);
or U8075 (N_8075,N_6168,N_5491);
nor U8076 (N_8076,N_6116,N_7057);
and U8077 (N_8077,N_6245,N_5412);
or U8078 (N_8078,N_6453,N_5879);
xor U8079 (N_8079,N_5894,N_6287);
and U8080 (N_8080,N_7126,N_6002);
nand U8081 (N_8081,N_7491,N_6191);
and U8082 (N_8082,N_7361,N_5070);
xnor U8083 (N_8083,N_5435,N_5613);
and U8084 (N_8084,N_5962,N_6311);
and U8085 (N_8085,N_6118,N_5918);
or U8086 (N_8086,N_6223,N_5793);
or U8087 (N_8087,N_5792,N_7198);
and U8088 (N_8088,N_5575,N_5544);
xnor U8089 (N_8089,N_7249,N_5991);
and U8090 (N_8090,N_6829,N_5574);
or U8091 (N_8091,N_5065,N_5034);
and U8092 (N_8092,N_6186,N_6940);
and U8093 (N_8093,N_5961,N_5746);
or U8094 (N_8094,N_5049,N_6905);
and U8095 (N_8095,N_6479,N_6280);
xnor U8096 (N_8096,N_5654,N_7459);
nor U8097 (N_8097,N_6357,N_5258);
nand U8098 (N_8098,N_7457,N_5816);
or U8099 (N_8099,N_5452,N_7245);
or U8100 (N_8100,N_7285,N_5664);
nand U8101 (N_8101,N_6217,N_7254);
xor U8102 (N_8102,N_7288,N_6204);
xnor U8103 (N_8103,N_5993,N_7302);
nor U8104 (N_8104,N_6896,N_7095);
nor U8105 (N_8105,N_7405,N_5717);
xnor U8106 (N_8106,N_5819,N_5600);
xor U8107 (N_8107,N_6532,N_5698);
xor U8108 (N_8108,N_7425,N_6354);
or U8109 (N_8109,N_6585,N_5384);
nor U8110 (N_8110,N_5304,N_5072);
and U8111 (N_8111,N_6811,N_6941);
and U8112 (N_8112,N_5288,N_7437);
nor U8113 (N_8113,N_7103,N_7114);
nand U8114 (N_8114,N_6107,N_6926);
xnor U8115 (N_8115,N_6549,N_5498);
and U8116 (N_8116,N_6039,N_6857);
or U8117 (N_8117,N_6692,N_5583);
nor U8118 (N_8118,N_6928,N_6844);
and U8119 (N_8119,N_6968,N_6362);
nand U8120 (N_8120,N_5370,N_6640);
and U8121 (N_8121,N_5278,N_5688);
nand U8122 (N_8122,N_6058,N_7075);
xor U8123 (N_8123,N_6843,N_6200);
nand U8124 (N_8124,N_6342,N_6837);
and U8125 (N_8125,N_5132,N_6486);
nor U8126 (N_8126,N_5089,N_6196);
or U8127 (N_8127,N_5198,N_5856);
and U8128 (N_8128,N_5611,N_6084);
and U8129 (N_8129,N_6604,N_6654);
nor U8130 (N_8130,N_5972,N_6176);
or U8131 (N_8131,N_6347,N_5030);
nand U8132 (N_8132,N_7261,N_6133);
or U8133 (N_8133,N_6514,N_6637);
nand U8134 (N_8134,N_5061,N_5355);
xnor U8135 (N_8135,N_5083,N_6628);
or U8136 (N_8136,N_6399,N_5863);
nand U8137 (N_8137,N_5236,N_6966);
and U8138 (N_8138,N_6062,N_5032);
or U8139 (N_8139,N_5855,N_5743);
xnor U8140 (N_8140,N_6629,N_6814);
nand U8141 (N_8141,N_5623,N_6577);
nor U8142 (N_8142,N_7183,N_5449);
and U8143 (N_8143,N_6491,N_5475);
nand U8144 (N_8144,N_6978,N_5603);
nor U8145 (N_8145,N_7291,N_5888);
nor U8146 (N_8146,N_7497,N_6197);
and U8147 (N_8147,N_6227,N_5944);
xnor U8148 (N_8148,N_5264,N_5377);
and U8149 (N_8149,N_5283,N_5152);
and U8150 (N_8150,N_5935,N_5763);
and U8151 (N_8151,N_7233,N_5459);
nand U8152 (N_8152,N_7464,N_5363);
nand U8153 (N_8153,N_7383,N_6752);
or U8154 (N_8154,N_5853,N_5666);
or U8155 (N_8155,N_5361,N_7223);
or U8156 (N_8156,N_5454,N_6647);
xnor U8157 (N_8157,N_7366,N_5716);
xnor U8158 (N_8158,N_5330,N_7193);
nor U8159 (N_8159,N_5776,N_7452);
nor U8160 (N_8160,N_5392,N_6846);
nor U8161 (N_8161,N_6387,N_7385);
or U8162 (N_8162,N_5562,N_7190);
nand U8163 (N_8163,N_5193,N_6327);
nand U8164 (N_8164,N_5394,N_7322);
xor U8165 (N_8165,N_5108,N_5483);
or U8166 (N_8166,N_7324,N_6035);
nand U8167 (N_8167,N_5956,N_5604);
xnor U8168 (N_8168,N_6195,N_7164);
and U8169 (N_8169,N_6631,N_5876);
nor U8170 (N_8170,N_5097,N_6886);
or U8171 (N_8171,N_6916,N_6800);
xor U8172 (N_8172,N_7479,N_5607);
xor U8173 (N_8173,N_7074,N_6803);
or U8174 (N_8174,N_5295,N_7044);
xnor U8175 (N_8175,N_5045,N_7030);
xor U8176 (N_8176,N_6626,N_5949);
nand U8177 (N_8177,N_7037,N_5335);
nor U8178 (N_8178,N_6997,N_7406);
nand U8179 (N_8179,N_5017,N_7387);
or U8180 (N_8180,N_5242,N_6216);
and U8181 (N_8181,N_6001,N_7118);
and U8182 (N_8182,N_7142,N_7260);
and U8183 (N_8183,N_6742,N_7308);
nor U8184 (N_8184,N_5665,N_5619);
xnor U8185 (N_8185,N_6336,N_7340);
xor U8186 (N_8186,N_5425,N_5968);
nor U8187 (N_8187,N_6537,N_6294);
and U8188 (N_8188,N_6858,N_5831);
nor U8189 (N_8189,N_7253,N_7010);
or U8190 (N_8190,N_7189,N_6780);
or U8191 (N_8191,N_7304,N_6726);
nor U8192 (N_8192,N_5313,N_6101);
xnor U8193 (N_8193,N_6681,N_6818);
xnor U8194 (N_8194,N_5474,N_6564);
or U8195 (N_8195,N_6317,N_5388);
xnor U8196 (N_8196,N_6778,N_6092);
or U8197 (N_8197,N_6254,N_5592);
nor U8198 (N_8198,N_6974,N_6913);
and U8199 (N_8199,N_7234,N_6733);
xor U8200 (N_8200,N_7060,N_6840);
xor U8201 (N_8201,N_7036,N_6955);
or U8202 (N_8202,N_5142,N_7420);
xnor U8203 (N_8203,N_6643,N_7151);
nand U8204 (N_8204,N_6504,N_6927);
and U8205 (N_8205,N_6835,N_5554);
or U8206 (N_8206,N_6817,N_6892);
nand U8207 (N_8207,N_5482,N_6371);
xor U8208 (N_8208,N_6384,N_7363);
and U8209 (N_8209,N_6144,N_6363);
nand U8210 (N_8210,N_6127,N_7477);
xnor U8211 (N_8211,N_5296,N_6447);
nor U8212 (N_8212,N_5546,N_7099);
and U8213 (N_8213,N_7478,N_5564);
nand U8214 (N_8214,N_5359,N_5616);
xnor U8215 (N_8215,N_5044,N_6527);
nand U8216 (N_8216,N_5320,N_5522);
nand U8217 (N_8217,N_6998,N_6309);
nand U8218 (N_8218,N_6379,N_7480);
xor U8219 (N_8219,N_6774,N_5516);
and U8220 (N_8220,N_5337,N_5114);
xnor U8221 (N_8221,N_5581,N_5488);
xor U8222 (N_8222,N_6805,N_5216);
nand U8223 (N_8223,N_5560,N_5929);
nor U8224 (N_8224,N_6569,N_5183);
nand U8225 (N_8225,N_5414,N_6307);
nand U8226 (N_8226,N_6476,N_5694);
or U8227 (N_8227,N_5197,N_5632);
or U8228 (N_8228,N_6596,N_5826);
nand U8229 (N_8229,N_5596,N_6961);
nor U8230 (N_8230,N_6724,N_6160);
or U8231 (N_8231,N_6177,N_6074);
nor U8232 (N_8232,N_6482,N_7086);
and U8233 (N_8233,N_6911,N_6548);
or U8234 (N_8234,N_5400,N_5648);
nand U8235 (N_8235,N_7155,N_5809);
nor U8236 (N_8236,N_6358,N_6304);
nor U8237 (N_8237,N_5805,N_5019);
and U8238 (N_8238,N_6781,N_6972);
or U8239 (N_8239,N_7091,N_5165);
xor U8240 (N_8240,N_6004,N_5634);
nor U8241 (N_8241,N_7284,N_6155);
xor U8242 (N_8242,N_6904,N_6456);
nor U8243 (N_8243,N_6860,N_6867);
or U8244 (N_8244,N_6003,N_5009);
xor U8245 (N_8245,N_6383,N_5824);
or U8246 (N_8246,N_6427,N_5589);
or U8247 (N_8247,N_5653,N_6493);
xnor U8248 (N_8248,N_5939,N_5609);
and U8249 (N_8249,N_5681,N_5750);
or U8250 (N_8250,N_7239,N_7204);
and U8251 (N_8251,N_6480,N_6785);
nor U8252 (N_8252,N_7321,N_5707);
nor U8253 (N_8253,N_5758,N_7225);
or U8254 (N_8254,N_6394,N_6189);
nor U8255 (N_8255,N_5958,N_5781);
nand U8256 (N_8256,N_6945,N_5451);
and U8257 (N_8257,N_6546,N_5378);
nand U8258 (N_8258,N_7244,N_7090);
or U8259 (N_8259,N_5830,N_5373);
and U8260 (N_8260,N_5397,N_5549);
nand U8261 (N_8261,N_5408,N_5317);
nor U8262 (N_8262,N_5804,N_5657);
and U8263 (N_8263,N_5755,N_5573);
nor U8264 (N_8264,N_5585,N_6563);
or U8265 (N_8265,N_6903,N_5795);
nor U8266 (N_8266,N_5841,N_5247);
and U8267 (N_8267,N_6932,N_7353);
nand U8268 (N_8268,N_5500,N_6758);
xor U8269 (N_8269,N_7093,N_7156);
xor U8270 (N_8270,N_5430,N_6508);
and U8271 (N_8271,N_5116,N_7265);
nand U8272 (N_8272,N_6833,N_6137);
nand U8273 (N_8273,N_5684,N_5553);
nor U8274 (N_8274,N_7072,N_6934);
xnor U8275 (N_8275,N_7019,N_5347);
or U8276 (N_8276,N_5037,N_6030);
nand U8277 (N_8277,N_5127,N_7323);
nand U8278 (N_8278,N_7028,N_6594);
nor U8279 (N_8279,N_6206,N_7082);
or U8280 (N_8280,N_5134,N_6117);
nor U8281 (N_8281,N_6221,N_6848);
or U8282 (N_8282,N_5102,N_6367);
and U8283 (N_8283,N_5559,N_6402);
and U8284 (N_8284,N_6776,N_6948);
nor U8285 (N_8285,N_6318,N_6852);
nand U8286 (N_8286,N_5473,N_6921);
and U8287 (N_8287,N_7391,N_7274);
or U8288 (N_8288,N_5737,N_5866);
and U8289 (N_8289,N_7411,N_6798);
xnor U8290 (N_8290,N_6694,N_6059);
and U8291 (N_8291,N_6203,N_6982);
xnor U8292 (N_8292,N_5239,N_5614);
and U8293 (N_8293,N_6425,N_7327);
nor U8294 (N_8294,N_5845,N_6923);
nand U8295 (N_8295,N_5651,N_5367);
or U8296 (N_8296,N_7209,N_5833);
or U8297 (N_8297,N_6881,N_5054);
xor U8298 (N_8298,N_6154,N_5661);
and U8299 (N_8299,N_6249,N_7434);
xor U8300 (N_8300,N_5110,N_5093);
and U8301 (N_8301,N_5101,N_5068);
xnor U8302 (N_8302,N_5537,N_6153);
or U8303 (N_8303,N_7088,N_6964);
or U8304 (N_8304,N_6882,N_7367);
nand U8305 (N_8305,N_6051,N_6696);
xnor U8306 (N_8306,N_5899,N_6722);
nor U8307 (N_8307,N_7123,N_6952);
nand U8308 (N_8308,N_6914,N_5467);
and U8309 (N_8309,N_6420,N_6055);
xor U8310 (N_8310,N_5601,N_5358);
nand U8311 (N_8311,N_6048,N_6233);
nand U8312 (N_8312,N_6271,N_7192);
nand U8313 (N_8313,N_5525,N_6842);
xor U8314 (N_8314,N_5982,N_5063);
nand U8315 (N_8315,N_5612,N_6283);
and U8316 (N_8316,N_6565,N_5875);
nor U8317 (N_8317,N_6158,N_7071);
nor U8318 (N_8318,N_7378,N_6653);
xor U8319 (N_8319,N_7108,N_6467);
nand U8320 (N_8320,N_5506,N_5595);
or U8321 (N_8321,N_7125,N_5137);
xor U8322 (N_8322,N_7017,N_6303);
and U8323 (N_8323,N_7440,N_5308);
xor U8324 (N_8324,N_6015,N_6635);
nand U8325 (N_8325,N_6390,N_6484);
nand U8326 (N_8326,N_6388,N_6253);
or U8327 (N_8327,N_6980,N_5140);
or U8328 (N_8328,N_6669,N_5031);
xor U8329 (N_8329,N_7107,N_5112);
xor U8330 (N_8330,N_6285,N_7298);
xnor U8331 (N_8331,N_5014,N_7175);
xnor U8332 (N_8332,N_5652,N_6296);
nor U8333 (N_8333,N_5528,N_5241);
nor U8334 (N_8334,N_6507,N_7217);
nor U8335 (N_8335,N_6411,N_5062);
nor U8336 (N_8336,N_5764,N_6268);
or U8337 (N_8337,N_6148,N_7145);
or U8338 (N_8338,N_6836,N_5445);
and U8339 (N_8339,N_6320,N_5080);
nor U8340 (N_8340,N_6888,N_5981);
nand U8341 (N_8341,N_7047,N_5835);
or U8342 (N_8342,N_6267,N_5450);
nor U8343 (N_8343,N_5673,N_7186);
nor U8344 (N_8344,N_6234,N_6869);
xor U8345 (N_8345,N_7456,N_5786);
nor U8346 (N_8346,N_6894,N_6109);
xor U8347 (N_8347,N_5011,N_7294);
nor U8348 (N_8348,N_6960,N_5638);
or U8349 (N_8349,N_5928,N_7168);
or U8350 (N_8350,N_7355,N_6011);
and U8351 (N_8351,N_5757,N_7221);
and U8352 (N_8352,N_5986,N_6122);
nand U8353 (N_8353,N_5287,N_6753);
and U8354 (N_8354,N_6775,N_5244);
nor U8355 (N_8355,N_5364,N_5353);
and U8356 (N_8356,N_6454,N_6880);
xnor U8357 (N_8357,N_6721,N_6992);
nand U8358 (N_8358,N_6381,N_6661);
or U8359 (N_8359,N_6481,N_6106);
nor U8360 (N_8360,N_6451,N_7026);
and U8361 (N_8361,N_7271,N_7236);
or U8362 (N_8362,N_5820,N_6135);
nor U8363 (N_8363,N_6884,N_6163);
and U8364 (N_8364,N_5490,N_5572);
and U8365 (N_8365,N_7386,N_6478);
nand U8366 (N_8366,N_5323,N_6147);
nand U8367 (N_8367,N_6090,N_5846);
and U8368 (N_8368,N_6741,N_7462);
xnor U8369 (N_8369,N_5143,N_6573);
nor U8370 (N_8370,N_6695,N_5325);
nand U8371 (N_8371,N_6730,N_7032);
nor U8372 (N_8372,N_5636,N_5413);
nand U8373 (N_8373,N_7379,N_6091);
nand U8374 (N_8374,N_6131,N_6097);
and U8375 (N_8375,N_5941,N_5164);
and U8376 (N_8376,N_7272,N_6534);
and U8377 (N_8377,N_5662,N_6686);
or U8378 (N_8378,N_6855,N_5422);
xor U8379 (N_8379,N_6143,N_5405);
nand U8380 (N_8380,N_6005,N_6706);
and U8381 (N_8381,N_7463,N_5567);
xor U8382 (N_8382,N_6123,N_6630);
nor U8383 (N_8383,N_6409,N_5380);
nand U8384 (N_8384,N_6337,N_5298);
nand U8385 (N_8385,N_7158,N_7264);
xnor U8386 (N_8386,N_5910,N_6236);
xor U8387 (N_8387,N_7282,N_6985);
nand U8388 (N_8388,N_5221,N_7493);
nor U8389 (N_8389,N_6827,N_6770);
xnor U8390 (N_8390,N_6193,N_5457);
nor U8391 (N_8391,N_5484,N_5906);
and U8392 (N_8392,N_6586,N_7338);
xor U8393 (N_8393,N_6208,N_5751);
or U8394 (N_8394,N_7492,N_7001);
nor U8395 (N_8395,N_5615,N_5458);
or U8396 (N_8396,N_6743,N_5109);
xnor U8397 (N_8397,N_7043,N_6670);
nor U8398 (N_8398,N_6652,N_7073);
nor U8399 (N_8399,N_5106,N_6745);
nor U8400 (N_8400,N_6792,N_6103);
nor U8401 (N_8401,N_6621,N_6738);
nor U8402 (N_8402,N_5727,N_5626);
and U8403 (N_8403,N_7427,N_6874);
nand U8404 (N_8404,N_5348,N_7034);
nand U8405 (N_8405,N_5741,N_5644);
xnor U8406 (N_8406,N_5545,N_5177);
and U8407 (N_8407,N_7305,N_7381);
xnor U8408 (N_8408,N_5504,N_6365);
nand U8409 (N_8409,N_6559,N_5489);
nand U8410 (N_8410,N_7122,N_6883);
and U8411 (N_8411,N_6764,N_6085);
and U8412 (N_8412,N_5733,N_6393);
xnor U8413 (N_8413,N_5344,N_6729);
nand U8414 (N_8414,N_5018,N_5479);
nand U8415 (N_8415,N_5007,N_5842);
nand U8416 (N_8416,N_7167,N_6607);
and U8417 (N_8417,N_7070,N_5259);
xnor U8418 (N_8418,N_5979,N_5909);
and U8419 (N_8419,N_5050,N_6545);
and U8420 (N_8420,N_6918,N_6539);
nor U8421 (N_8421,N_5411,N_7227);
or U8422 (N_8422,N_6831,N_6826);
xor U8423 (N_8423,N_7080,N_5349);
and U8424 (N_8424,N_7160,N_6046);
or U8425 (N_8425,N_6181,N_5983);
and U8426 (N_8426,N_6501,N_6272);
nand U8427 (N_8427,N_6705,N_7467);
nand U8428 (N_8428,N_5812,N_5710);
or U8429 (N_8429,N_6580,N_6897);
xnor U8430 (N_8430,N_6300,N_6326);
nand U8431 (N_8431,N_6255,N_6687);
nand U8432 (N_8432,N_5829,N_5372);
nand U8433 (N_8433,N_6566,N_5133);
nand U8434 (N_8434,N_6720,N_5514);
and U8435 (N_8435,N_7368,N_5023);
nand U8436 (N_8436,N_6019,N_6180);
and U8437 (N_8437,N_7174,N_6325);
nand U8438 (N_8438,N_7206,N_6790);
xnor U8439 (N_8439,N_6516,N_6513);
nand U8440 (N_8440,N_5628,N_5000);
nand U8441 (N_8441,N_7159,N_5858);
nor U8442 (N_8442,N_5410,N_5436);
nor U8443 (N_8443,N_6464,N_6471);
nor U8444 (N_8444,N_5076,N_6356);
and U8445 (N_8445,N_6359,N_5156);
and U8446 (N_8446,N_6646,N_5096);
nand U8447 (N_8447,N_5402,N_6057);
xnor U8448 (N_8448,N_5523,N_5379);
xnor U8449 (N_8449,N_6600,N_6291);
or U8450 (N_8450,N_6096,N_6487);
xnor U8451 (N_8451,N_7216,N_5625);
nand U8452 (N_8452,N_7214,N_5172);
nand U8453 (N_8453,N_5766,N_6824);
or U8454 (N_8454,N_7433,N_7134);
nor U8455 (N_8455,N_6676,N_5580);
xor U8456 (N_8456,N_6115,N_5851);
and U8457 (N_8457,N_5495,N_5487);
nand U8458 (N_8458,N_5967,N_6727);
nand U8459 (N_8459,N_6984,N_6925);
nand U8460 (N_8460,N_7301,N_6693);
and U8461 (N_8461,N_5001,N_7471);
xnor U8462 (N_8462,N_6862,N_5419);
and U8463 (N_8463,N_6006,N_7476);
nor U8464 (N_8464,N_5916,N_6828);
xor U8465 (N_8465,N_5798,N_5243);
xnor U8466 (N_8466,N_7181,N_7403);
nor U8467 (N_8467,N_6149,N_6014);
xnor U8468 (N_8468,N_6891,N_7205);
xnor U8469 (N_8469,N_5208,N_5696);
or U8470 (N_8470,N_6049,N_7016);
nor U8471 (N_8471,N_7146,N_6157);
nand U8472 (N_8472,N_5209,N_5069);
nand U8473 (N_8473,N_6378,N_5439);
nand U8474 (N_8474,N_5932,N_6114);
or U8475 (N_8475,N_6126,N_5996);
nor U8476 (N_8476,N_7147,N_5179);
xnor U8477 (N_8477,N_7330,N_6026);
or U8478 (N_8478,N_6702,N_6575);
nor U8479 (N_8479,N_5158,N_6345);
nand U8480 (N_8480,N_6572,N_5182);
nand U8481 (N_8481,N_6275,N_5885);
and U8482 (N_8482,N_7318,N_5754);
nor U8483 (N_8483,N_7371,N_5577);
or U8484 (N_8484,N_6417,N_5898);
xnor U8485 (N_8485,N_7445,N_5650);
nand U8486 (N_8486,N_5768,N_6887);
or U8487 (N_8487,N_5122,N_6212);
nor U8488 (N_8488,N_6364,N_5627);
nand U8489 (N_8489,N_5779,N_7258);
nor U8490 (N_8490,N_6042,N_5620);
and U8491 (N_8491,N_6875,N_5606);
or U8492 (N_8492,N_7150,N_5570);
nand U8493 (N_8493,N_6708,N_6503);
and U8494 (N_8494,N_5729,N_7089);
and U8495 (N_8495,N_7251,N_7067);
or U8496 (N_8496,N_6593,N_5501);
nor U8497 (N_8497,N_5843,N_6372);
nor U8498 (N_8498,N_6815,N_5960);
and U8499 (N_8499,N_6963,N_6936);
and U8500 (N_8500,N_5279,N_5354);
or U8501 (N_8501,N_6313,N_5326);
nand U8502 (N_8502,N_5421,N_6988);
nor U8503 (N_8503,N_7023,N_6731);
or U8504 (N_8504,N_5602,N_7162);
nor U8505 (N_8505,N_5827,N_5736);
or U8506 (N_8506,N_5094,N_5170);
nand U8507 (N_8507,N_5663,N_6056);
and U8508 (N_8508,N_6766,N_5162);
nor U8509 (N_8509,N_5887,N_5276);
or U8510 (N_8510,N_6801,N_5048);
nand U8511 (N_8511,N_6025,N_6416);
or U8512 (N_8512,N_5922,N_6779);
nand U8513 (N_8513,N_6605,N_6597);
and U8514 (N_8514,N_6041,N_6495);
nor U8515 (N_8515,N_6423,N_7454);
xor U8516 (N_8516,N_7105,N_6587);
and U8517 (N_8517,N_5066,N_6339);
or U8518 (N_8518,N_7394,N_5883);
nor U8519 (N_8519,N_6441,N_6680);
and U8520 (N_8520,N_6868,N_6214);
or U8521 (N_8521,N_5492,N_7447);
and U8522 (N_8522,N_5925,N_7171);
or U8523 (N_8523,N_7250,N_7490);
nor U8524 (N_8524,N_5834,N_5767);
xnor U8525 (N_8525,N_5343,N_6315);
xnor U8526 (N_8526,N_6053,N_5409);
xnor U8527 (N_8527,N_7307,N_6787);
nand U8528 (N_8528,N_5718,N_6373);
or U8529 (N_8529,N_6822,N_6010);
nor U8530 (N_8530,N_6080,N_5884);
or U8531 (N_8531,N_5047,N_5629);
nand U8532 (N_8532,N_5478,N_6583);
nor U8533 (N_8533,N_6644,N_5416);
nor U8534 (N_8534,N_6544,N_6898);
nor U8535 (N_8535,N_7450,N_5773);
xnor U8536 (N_8536,N_5033,N_7455);
xor U8537 (N_8537,N_5953,N_7358);
nor U8538 (N_8538,N_5497,N_7098);
and U8539 (N_8539,N_5789,N_6492);
and U8540 (N_8540,N_6063,N_6446);
nor U8541 (N_8541,N_7481,N_5028);
nand U8542 (N_8542,N_5041,N_6104);
or U8543 (N_8543,N_7346,N_6665);
nand U8544 (N_8544,N_5341,N_5584);
nand U8545 (N_8545,N_5507,N_5055);
xor U8546 (N_8546,N_7345,N_6530);
nor U8547 (N_8547,N_6994,N_5722);
and U8548 (N_8548,N_5919,N_5869);
nor U8549 (N_8549,N_5903,N_6064);
nand U8550 (N_8550,N_7237,N_6050);
xor U8551 (N_8551,N_5783,N_5502);
and U8552 (N_8552,N_5481,N_5220);
xor U8553 (N_8553,N_5543,N_7400);
and U8554 (N_8554,N_7006,N_7121);
or U8555 (N_8555,N_6515,N_5984);
nand U8556 (N_8556,N_5637,N_5641);
nand U8557 (N_8557,N_5690,N_5407);
xnor U8558 (N_8558,N_5223,N_6500);
nand U8559 (N_8559,N_5732,N_6908);
nor U8560 (N_8560,N_5245,N_5724);
or U8561 (N_8561,N_6810,N_6616);
or U8562 (N_8562,N_7053,N_7084);
nand U8563 (N_8563,N_5119,N_6536);
nor U8564 (N_8564,N_5675,N_5012);
xnor U8565 (N_8565,N_6870,N_6000);
and U8566 (N_8566,N_6346,N_5593);
xnor U8567 (N_8567,N_6825,N_5825);
xnor U8568 (N_8568,N_5565,N_5440);
xnor U8569 (N_8569,N_5319,N_6876);
nor U8570 (N_8570,N_6466,N_6224);
nor U8571 (N_8571,N_5897,N_6278);
nor U8572 (N_8572,N_5082,N_5415);
or U8573 (N_8573,N_7442,N_5803);
nor U8574 (N_8574,N_6328,N_5206);
and U8575 (N_8575,N_7315,N_7356);
xnor U8576 (N_8576,N_7263,N_6697);
and U8577 (N_8577,N_5740,N_6146);
or U8578 (N_8578,N_6496,N_5617);
and U8579 (N_8579,N_6797,N_5229);
nor U8580 (N_8580,N_5723,N_6036);
xor U8581 (N_8581,N_6499,N_5965);
nand U8582 (N_8582,N_5964,N_6273);
xnor U8583 (N_8583,N_5207,N_6553);
nor U8584 (N_8584,N_5864,N_5777);
or U8585 (N_8585,N_6013,N_5426);
and U8586 (N_8586,N_6231,N_5676);
nor U8587 (N_8587,N_6995,N_5911);
or U8588 (N_8588,N_7210,N_6439);
or U8589 (N_8589,N_6412,N_5113);
nor U8590 (N_8590,N_6550,N_6382);
and U8591 (N_8591,N_6642,N_5273);
or U8592 (N_8592,N_7004,N_6323);
xnor U8593 (N_8593,N_5128,N_6183);
and U8594 (N_8594,N_5131,N_7055);
nor U8595 (N_8595,N_7495,N_6334);
nand U8596 (N_8596,N_5246,N_5511);
and U8597 (N_8597,N_6027,N_5462);
nand U8598 (N_8598,N_6277,N_6418);
nor U8599 (N_8599,N_6712,N_6609);
nand U8600 (N_8600,N_6751,N_6622);
or U8601 (N_8601,N_5365,N_6551);
and U8602 (N_8602,N_6864,N_6355);
nand U8603 (N_8603,N_5153,N_6987);
nand U8604 (N_8604,N_6783,N_6768);
and U8605 (N_8605,N_6435,N_6209);
xor U8606 (N_8606,N_6301,N_5013);
xor U8607 (N_8607,N_6299,N_5444);
and U8608 (N_8608,N_5677,N_5889);
nand U8609 (N_8609,N_5886,N_5306);
xnor U8610 (N_8610,N_5427,N_6689);
or U8611 (N_8611,N_7139,N_6403);
nand U8612 (N_8612,N_6521,N_5022);
nor U8613 (N_8613,N_5703,N_6202);
nor U8614 (N_8614,N_6602,N_6349);
nand U8615 (N_8615,N_6772,N_7170);
nor U8616 (N_8616,N_6699,N_5963);
xor U8617 (N_8617,N_6556,N_6866);
nor U8618 (N_8618,N_6991,N_5760);
xor U8619 (N_8619,N_5924,N_5934);
nand U8620 (N_8620,N_5704,N_7180);
or U8621 (N_8621,N_7416,N_5715);
and U8622 (N_8622,N_5398,N_5980);
xnor U8623 (N_8623,N_6111,N_6639);
or U8624 (N_8624,N_5709,N_7232);
xor U8625 (N_8625,N_6659,N_7247);
and U8626 (N_8626,N_7277,N_5079);
or U8627 (N_8627,N_6072,N_5261);
and U8628 (N_8628,N_5252,N_5989);
nand U8629 (N_8629,N_6707,N_6141);
nor U8630 (N_8630,N_6744,N_5998);
and U8631 (N_8631,N_6606,N_7141);
or U8632 (N_8632,N_6981,N_6541);
nor U8633 (N_8633,N_5190,N_7243);
nor U8634 (N_8634,N_7410,N_7015);
or U8635 (N_8635,N_5971,N_5226);
nand U8636 (N_8636,N_5901,N_5442);
and U8637 (N_8637,N_5327,N_6073);
and U8638 (N_8638,N_6419,N_6962);
and U8639 (N_8639,N_6494,N_5144);
or U8640 (N_8640,N_6151,N_6366);
and U8641 (N_8641,N_6434,N_5138);
or U8642 (N_8642,N_6448,N_5270);
or U8643 (N_8643,N_6477,N_7109);
nor U8644 (N_8644,N_7048,N_5558);
or U8645 (N_8645,N_5817,N_5865);
and U8646 (N_8646,N_5590,N_6395);
nand U8647 (N_8647,N_6929,N_6762);
nor U8648 (N_8648,N_6759,N_5926);
or U8649 (N_8649,N_5085,N_5147);
nand U8650 (N_8650,N_6502,N_6717);
and U8651 (N_8651,N_7011,N_7111);
xnor U8652 (N_8652,N_6522,N_6688);
xor U8653 (N_8653,N_5633,N_7130);
or U8654 (N_8654,N_7461,N_7472);
or U8655 (N_8655,N_7003,N_5702);
nor U8656 (N_8656,N_5749,N_7117);
or U8657 (N_8657,N_5647,N_7152);
xor U8658 (N_8658,N_5200,N_7076);
nand U8659 (N_8659,N_5890,N_6038);
nor U8660 (N_8660,N_7061,N_7131);
xor U8661 (N_8661,N_5772,N_5480);
xor U8662 (N_8662,N_6220,N_7279);
nand U8663 (N_8663,N_6385,N_6528);
xor U8664 (N_8664,N_5005,N_6108);
xnor U8665 (N_8665,N_5042,N_5429);
xor U8666 (N_8666,N_5433,N_5713);
or U8667 (N_8667,N_5472,N_6715);
nand U8668 (N_8668,N_6650,N_5250);
and U8669 (N_8669,N_6424,N_7120);
or U8670 (N_8670,N_6007,N_5092);
and U8671 (N_8671,N_5075,N_6841);
or U8672 (N_8672,N_6613,N_6376);
xor U8673 (N_8673,N_5046,N_6910);
nand U8674 (N_8674,N_5039,N_5167);
or U8675 (N_8675,N_6119,N_6222);
and U8676 (N_8676,N_5231,N_6165);
or U8677 (N_8677,N_5578,N_6601);
or U8678 (N_8678,N_6230,N_6129);
and U8679 (N_8679,N_6560,N_6944);
or U8680 (N_8680,N_5463,N_7446);
xnor U8681 (N_8681,N_5551,N_7024);
nor U8682 (N_8682,N_6789,N_6608);
xor U8683 (N_8683,N_5571,N_6951);
or U8684 (N_8684,N_6289,N_6185);
and U8685 (N_8685,N_5635,N_6341);
xor U8686 (N_8686,N_5942,N_5679);
and U8687 (N_8687,N_6099,N_6102);
nor U8688 (N_8688,N_6428,N_5659);
nor U8689 (N_8689,N_6711,N_5387);
or U8690 (N_8690,N_7008,N_5937);
xnor U8691 (N_8691,N_6033,N_6567);
nor U8692 (N_8692,N_5556,N_7382);
xnor U8693 (N_8693,N_7242,N_6169);
nand U8694 (N_8694,N_5424,N_5576);
nand U8695 (N_8695,N_5136,N_6614);
nand U8696 (N_8696,N_5211,N_5655);
nand U8697 (N_8697,N_5505,N_6975);
nand U8698 (N_8698,N_5111,N_7469);
nand U8699 (N_8699,N_6931,N_6675);
nor U8700 (N_8700,N_6375,N_5015);
or U8701 (N_8701,N_7365,N_7448);
nand U8702 (N_8702,N_6239,N_6485);
nand U8703 (N_8703,N_7224,N_5060);
nand U8704 (N_8704,N_5930,N_7389);
nand U8705 (N_8705,N_6483,N_6225);
xnor U8706 (N_8706,N_7465,N_6794);
xnor U8707 (N_8707,N_6612,N_7484);
xor U8708 (N_8708,N_6784,N_6678);
and U8709 (N_8709,N_6105,N_6623);
xor U8710 (N_8710,N_6638,N_6110);
nor U8711 (N_8711,N_5095,N_6297);
or U8712 (N_8712,N_7068,N_6240);
and U8713 (N_8713,N_5057,N_5237);
nor U8714 (N_8714,N_5124,N_5404);
xor U8715 (N_8715,N_5943,N_5224);
xor U8716 (N_8716,N_6591,N_6907);
nand U8717 (N_8717,N_6316,N_5432);
xnor U8718 (N_8718,N_6529,N_7357);
xor U8719 (N_8719,N_6429,N_5105);
xor U8720 (N_8720,N_5705,N_5823);
nor U8721 (N_8721,N_5891,N_5448);
or U8722 (N_8722,N_5987,N_6431);
or U8723 (N_8723,N_6582,N_6838);
and U8724 (N_8724,N_5494,N_6683);
nor U8725 (N_8725,N_6906,N_6190);
or U8726 (N_8726,N_5499,N_7349);
nor U8727 (N_8727,N_5871,N_7267);
and U8728 (N_8728,N_5471,N_6933);
nand U8729 (N_8729,N_5782,N_7063);
nand U8730 (N_8730,N_5813,N_5587);
or U8731 (N_8731,N_5315,N_5708);
nand U8732 (N_8732,N_7140,N_6198);
or U8733 (N_8733,N_6279,N_7306);
and U8734 (N_8734,N_6947,N_7212);
nor U8735 (N_8735,N_5280,N_6909);
nor U8736 (N_8736,N_5038,N_5021);
and U8737 (N_8737,N_5880,N_6839);
and U8738 (N_8738,N_7296,N_6401);
and U8739 (N_8739,N_5071,N_5970);
or U8740 (N_8740,N_5933,N_5975);
nor U8741 (N_8741,N_5350,N_6570);
nand U8742 (N_8742,N_5801,N_5008);
nand U8743 (N_8743,N_6845,N_7163);
nor U8744 (N_8744,N_6353,N_6444);
or U8745 (N_8745,N_6218,N_7211);
nor U8746 (N_8746,N_5345,N_7040);
xnor U8747 (N_8747,N_6767,N_6547);
nand U8748 (N_8748,N_7022,N_5769);
and U8749 (N_8749,N_5126,N_7408);
xor U8750 (N_8750,N_6554,N_7348);
nand U8751 (N_8751,N_6458,N_5540);
xor U8752 (N_8752,N_5363,N_6465);
and U8753 (N_8753,N_6857,N_5187);
nand U8754 (N_8754,N_5782,N_5465);
xnor U8755 (N_8755,N_5893,N_5584);
nor U8756 (N_8756,N_5114,N_7260);
or U8757 (N_8757,N_6532,N_7279);
xnor U8758 (N_8758,N_6376,N_5583);
nor U8759 (N_8759,N_6314,N_5714);
or U8760 (N_8760,N_6635,N_5874);
and U8761 (N_8761,N_5410,N_5242);
and U8762 (N_8762,N_7194,N_5738);
xnor U8763 (N_8763,N_6762,N_6206);
xor U8764 (N_8764,N_7004,N_5224);
nor U8765 (N_8765,N_5177,N_6061);
nor U8766 (N_8766,N_7485,N_5706);
and U8767 (N_8767,N_6809,N_5006);
or U8768 (N_8768,N_6990,N_5049);
nand U8769 (N_8769,N_7120,N_5748);
nor U8770 (N_8770,N_7162,N_5592);
xor U8771 (N_8771,N_7371,N_5971);
nor U8772 (N_8772,N_5287,N_7287);
xor U8773 (N_8773,N_6759,N_6523);
nand U8774 (N_8774,N_6524,N_5296);
or U8775 (N_8775,N_7057,N_7484);
nor U8776 (N_8776,N_6490,N_5165);
nor U8777 (N_8777,N_7283,N_5355);
nor U8778 (N_8778,N_6185,N_5886);
and U8779 (N_8779,N_6765,N_5976);
and U8780 (N_8780,N_5519,N_7355);
xnor U8781 (N_8781,N_5339,N_5995);
or U8782 (N_8782,N_7325,N_7293);
nand U8783 (N_8783,N_5778,N_5815);
xor U8784 (N_8784,N_6219,N_7335);
or U8785 (N_8785,N_6572,N_6922);
nor U8786 (N_8786,N_5127,N_5858);
nor U8787 (N_8787,N_6159,N_5390);
and U8788 (N_8788,N_6920,N_7042);
nand U8789 (N_8789,N_7258,N_5953);
xor U8790 (N_8790,N_6265,N_6750);
nand U8791 (N_8791,N_5870,N_6107);
and U8792 (N_8792,N_6729,N_6921);
nand U8793 (N_8793,N_5993,N_6777);
or U8794 (N_8794,N_5034,N_5167);
xor U8795 (N_8795,N_7350,N_5492);
or U8796 (N_8796,N_6384,N_5366);
and U8797 (N_8797,N_6024,N_6085);
nand U8798 (N_8798,N_5306,N_7361);
nand U8799 (N_8799,N_5188,N_6231);
xor U8800 (N_8800,N_6943,N_6051);
nor U8801 (N_8801,N_7441,N_5777);
xnor U8802 (N_8802,N_6628,N_5618);
xor U8803 (N_8803,N_7388,N_6162);
nor U8804 (N_8804,N_5987,N_6068);
nor U8805 (N_8805,N_6153,N_5375);
or U8806 (N_8806,N_5138,N_7100);
nand U8807 (N_8807,N_6386,N_5828);
xnor U8808 (N_8808,N_6798,N_6387);
and U8809 (N_8809,N_5455,N_5771);
nor U8810 (N_8810,N_6312,N_5556);
nor U8811 (N_8811,N_5000,N_6587);
xnor U8812 (N_8812,N_6901,N_5100);
nor U8813 (N_8813,N_7091,N_5825);
nand U8814 (N_8814,N_5206,N_6598);
and U8815 (N_8815,N_5056,N_6665);
and U8816 (N_8816,N_5069,N_5599);
nand U8817 (N_8817,N_5550,N_6364);
and U8818 (N_8818,N_5408,N_7233);
and U8819 (N_8819,N_6445,N_7252);
nor U8820 (N_8820,N_6359,N_6700);
xnor U8821 (N_8821,N_6884,N_6636);
nor U8822 (N_8822,N_7211,N_6919);
xnor U8823 (N_8823,N_5336,N_5041);
nor U8824 (N_8824,N_5605,N_6909);
nor U8825 (N_8825,N_6802,N_6038);
nor U8826 (N_8826,N_7173,N_7074);
nor U8827 (N_8827,N_6510,N_5761);
xor U8828 (N_8828,N_5153,N_5623);
nand U8829 (N_8829,N_5521,N_5181);
xor U8830 (N_8830,N_6056,N_6861);
and U8831 (N_8831,N_5127,N_6781);
or U8832 (N_8832,N_7065,N_7367);
xnor U8833 (N_8833,N_7001,N_6278);
or U8834 (N_8834,N_5049,N_5075);
and U8835 (N_8835,N_5095,N_6418);
nor U8836 (N_8836,N_6648,N_5291);
or U8837 (N_8837,N_7488,N_6942);
and U8838 (N_8838,N_6262,N_7424);
nand U8839 (N_8839,N_6188,N_7098);
nand U8840 (N_8840,N_6692,N_6213);
nor U8841 (N_8841,N_5879,N_5730);
or U8842 (N_8842,N_5745,N_6386);
xor U8843 (N_8843,N_6332,N_7310);
or U8844 (N_8844,N_6312,N_5665);
or U8845 (N_8845,N_6093,N_7007);
xnor U8846 (N_8846,N_6489,N_5843);
or U8847 (N_8847,N_6003,N_6738);
and U8848 (N_8848,N_5013,N_6795);
nand U8849 (N_8849,N_6686,N_6088);
nor U8850 (N_8850,N_5133,N_5989);
nor U8851 (N_8851,N_6287,N_5063);
nand U8852 (N_8852,N_5033,N_7244);
and U8853 (N_8853,N_5832,N_6835);
nor U8854 (N_8854,N_5121,N_6120);
nand U8855 (N_8855,N_6274,N_5652);
nor U8856 (N_8856,N_6928,N_6685);
nand U8857 (N_8857,N_5562,N_5011);
nor U8858 (N_8858,N_5119,N_6667);
nor U8859 (N_8859,N_6057,N_5911);
nor U8860 (N_8860,N_6134,N_6351);
nand U8861 (N_8861,N_6412,N_5012);
and U8862 (N_8862,N_6528,N_6616);
xnor U8863 (N_8863,N_5559,N_7273);
xnor U8864 (N_8864,N_6185,N_6244);
xor U8865 (N_8865,N_5624,N_6745);
xor U8866 (N_8866,N_7224,N_5326);
and U8867 (N_8867,N_6975,N_5485);
and U8868 (N_8868,N_5160,N_6705);
nand U8869 (N_8869,N_5150,N_7393);
xnor U8870 (N_8870,N_6985,N_6359);
xnor U8871 (N_8871,N_7462,N_5671);
or U8872 (N_8872,N_6877,N_5857);
and U8873 (N_8873,N_7288,N_5562);
nand U8874 (N_8874,N_5487,N_5122);
nor U8875 (N_8875,N_7431,N_5960);
or U8876 (N_8876,N_5512,N_7136);
xnor U8877 (N_8877,N_5409,N_5583);
xor U8878 (N_8878,N_6851,N_7051);
xor U8879 (N_8879,N_7157,N_6988);
nand U8880 (N_8880,N_7403,N_5645);
nor U8881 (N_8881,N_6135,N_7255);
nor U8882 (N_8882,N_5872,N_5998);
nand U8883 (N_8883,N_5419,N_6977);
nand U8884 (N_8884,N_6413,N_6263);
nand U8885 (N_8885,N_5646,N_5941);
and U8886 (N_8886,N_5498,N_7266);
nand U8887 (N_8887,N_6649,N_6124);
and U8888 (N_8888,N_6896,N_6872);
xor U8889 (N_8889,N_6282,N_7278);
xnor U8890 (N_8890,N_5072,N_7396);
nand U8891 (N_8891,N_5363,N_5758);
nand U8892 (N_8892,N_5847,N_6301);
xnor U8893 (N_8893,N_6531,N_5817);
xor U8894 (N_8894,N_6373,N_7456);
nor U8895 (N_8895,N_7336,N_7244);
xnor U8896 (N_8896,N_6766,N_7455);
nand U8897 (N_8897,N_6703,N_6552);
or U8898 (N_8898,N_5910,N_5447);
nor U8899 (N_8899,N_5943,N_5549);
nand U8900 (N_8900,N_5304,N_5188);
nand U8901 (N_8901,N_5623,N_6373);
or U8902 (N_8902,N_7077,N_6078);
and U8903 (N_8903,N_7442,N_6745);
or U8904 (N_8904,N_6633,N_5597);
xnor U8905 (N_8905,N_6528,N_6525);
xnor U8906 (N_8906,N_5622,N_6802);
or U8907 (N_8907,N_6332,N_7350);
xor U8908 (N_8908,N_6914,N_6185);
xnor U8909 (N_8909,N_5387,N_7197);
nand U8910 (N_8910,N_7485,N_7149);
xnor U8911 (N_8911,N_6872,N_7422);
and U8912 (N_8912,N_6914,N_6830);
or U8913 (N_8913,N_6679,N_6186);
and U8914 (N_8914,N_5138,N_6364);
nand U8915 (N_8915,N_5544,N_6698);
nor U8916 (N_8916,N_6000,N_7314);
nor U8917 (N_8917,N_7153,N_6715);
nand U8918 (N_8918,N_7489,N_5984);
or U8919 (N_8919,N_7343,N_5631);
or U8920 (N_8920,N_6282,N_6626);
xnor U8921 (N_8921,N_6124,N_5961);
or U8922 (N_8922,N_5605,N_5200);
nand U8923 (N_8923,N_5314,N_5507);
nand U8924 (N_8924,N_6808,N_7341);
nor U8925 (N_8925,N_7493,N_6617);
or U8926 (N_8926,N_6288,N_6592);
or U8927 (N_8927,N_6951,N_5735);
nor U8928 (N_8928,N_5462,N_6605);
xnor U8929 (N_8929,N_7495,N_5318);
nand U8930 (N_8930,N_6463,N_7245);
nand U8931 (N_8931,N_7144,N_7022);
or U8932 (N_8932,N_5864,N_6795);
nand U8933 (N_8933,N_7255,N_5128);
and U8934 (N_8934,N_5404,N_6273);
xor U8935 (N_8935,N_5191,N_6404);
nor U8936 (N_8936,N_6523,N_6476);
and U8937 (N_8937,N_5025,N_6230);
nor U8938 (N_8938,N_5591,N_7388);
nor U8939 (N_8939,N_5003,N_6291);
and U8940 (N_8940,N_7014,N_5799);
and U8941 (N_8941,N_6868,N_6440);
or U8942 (N_8942,N_7026,N_5670);
and U8943 (N_8943,N_6569,N_6095);
or U8944 (N_8944,N_6558,N_5064);
or U8945 (N_8945,N_6900,N_5917);
and U8946 (N_8946,N_6292,N_6048);
or U8947 (N_8947,N_5317,N_6201);
or U8948 (N_8948,N_5674,N_6668);
or U8949 (N_8949,N_7342,N_6321);
and U8950 (N_8950,N_5696,N_6894);
nor U8951 (N_8951,N_5259,N_5959);
nand U8952 (N_8952,N_7112,N_5509);
nor U8953 (N_8953,N_6795,N_5227);
nor U8954 (N_8954,N_6274,N_5037);
or U8955 (N_8955,N_6344,N_5060);
nand U8956 (N_8956,N_6841,N_7380);
or U8957 (N_8957,N_5034,N_6837);
and U8958 (N_8958,N_6263,N_5976);
xnor U8959 (N_8959,N_6537,N_6253);
xor U8960 (N_8960,N_7170,N_7367);
nor U8961 (N_8961,N_5652,N_6350);
and U8962 (N_8962,N_5323,N_5691);
and U8963 (N_8963,N_5049,N_6618);
or U8964 (N_8964,N_6607,N_7419);
nor U8965 (N_8965,N_5628,N_5923);
and U8966 (N_8966,N_6093,N_5510);
and U8967 (N_8967,N_5308,N_7210);
nor U8968 (N_8968,N_5574,N_5214);
nand U8969 (N_8969,N_6844,N_5911);
xor U8970 (N_8970,N_5113,N_7002);
xnor U8971 (N_8971,N_5900,N_6297);
and U8972 (N_8972,N_6833,N_6613);
and U8973 (N_8973,N_5020,N_5175);
xor U8974 (N_8974,N_5109,N_5931);
or U8975 (N_8975,N_7218,N_6732);
and U8976 (N_8976,N_5193,N_5677);
and U8977 (N_8977,N_6398,N_5273);
nand U8978 (N_8978,N_5123,N_6674);
or U8979 (N_8979,N_5757,N_6306);
or U8980 (N_8980,N_5637,N_5137);
and U8981 (N_8981,N_6604,N_5585);
or U8982 (N_8982,N_5760,N_5325);
or U8983 (N_8983,N_5846,N_6524);
and U8984 (N_8984,N_6575,N_7222);
and U8985 (N_8985,N_6270,N_6621);
xor U8986 (N_8986,N_6362,N_6952);
xnor U8987 (N_8987,N_5242,N_6114);
or U8988 (N_8988,N_5461,N_6299);
nor U8989 (N_8989,N_5950,N_6775);
nor U8990 (N_8990,N_5387,N_6207);
nand U8991 (N_8991,N_5660,N_6872);
nor U8992 (N_8992,N_6118,N_7226);
nand U8993 (N_8993,N_5493,N_6291);
or U8994 (N_8994,N_7205,N_6206);
or U8995 (N_8995,N_7143,N_7305);
or U8996 (N_8996,N_5286,N_6520);
nand U8997 (N_8997,N_5715,N_5842);
nor U8998 (N_8998,N_5494,N_6857);
nor U8999 (N_8999,N_6934,N_7190);
nor U9000 (N_9000,N_7333,N_6938);
xor U9001 (N_9001,N_6778,N_6007);
and U9002 (N_9002,N_6143,N_6638);
nand U9003 (N_9003,N_6081,N_5870);
nor U9004 (N_9004,N_6876,N_5355);
or U9005 (N_9005,N_6795,N_5315);
xor U9006 (N_9006,N_7014,N_6887);
nand U9007 (N_9007,N_7266,N_5874);
or U9008 (N_9008,N_7278,N_5393);
nor U9009 (N_9009,N_6281,N_5740);
or U9010 (N_9010,N_6297,N_6496);
or U9011 (N_9011,N_5085,N_6798);
nand U9012 (N_9012,N_5991,N_7059);
nor U9013 (N_9013,N_5379,N_6153);
xor U9014 (N_9014,N_6820,N_6628);
nor U9015 (N_9015,N_6690,N_6604);
or U9016 (N_9016,N_6690,N_6523);
nand U9017 (N_9017,N_6590,N_6507);
nor U9018 (N_9018,N_5416,N_7421);
and U9019 (N_9019,N_6141,N_6922);
xnor U9020 (N_9020,N_5704,N_5277);
or U9021 (N_9021,N_7129,N_6273);
xor U9022 (N_9022,N_7287,N_5282);
or U9023 (N_9023,N_6996,N_6200);
nor U9024 (N_9024,N_7199,N_6514);
xor U9025 (N_9025,N_5751,N_5490);
nor U9026 (N_9026,N_7041,N_5209);
nand U9027 (N_9027,N_5905,N_6274);
nor U9028 (N_9028,N_5936,N_5042);
or U9029 (N_9029,N_6310,N_5609);
nor U9030 (N_9030,N_5814,N_7034);
or U9031 (N_9031,N_5104,N_7224);
nand U9032 (N_9032,N_7404,N_5463);
xnor U9033 (N_9033,N_6313,N_6817);
and U9034 (N_9034,N_6224,N_6512);
nor U9035 (N_9035,N_7036,N_5642);
and U9036 (N_9036,N_5545,N_6000);
or U9037 (N_9037,N_5335,N_7255);
nand U9038 (N_9038,N_6626,N_5182);
or U9039 (N_9039,N_5997,N_6247);
nand U9040 (N_9040,N_5846,N_6857);
nand U9041 (N_9041,N_5493,N_7078);
nand U9042 (N_9042,N_6611,N_5031);
xor U9043 (N_9043,N_5809,N_5434);
and U9044 (N_9044,N_7268,N_5654);
nand U9045 (N_9045,N_7357,N_5105);
xor U9046 (N_9046,N_5592,N_6236);
nor U9047 (N_9047,N_6186,N_5132);
xnor U9048 (N_9048,N_6171,N_5667);
or U9049 (N_9049,N_7124,N_7270);
nor U9050 (N_9050,N_7410,N_5662);
xor U9051 (N_9051,N_6140,N_6343);
nor U9052 (N_9052,N_5757,N_5707);
nor U9053 (N_9053,N_7207,N_6169);
or U9054 (N_9054,N_6213,N_7402);
or U9055 (N_9055,N_6256,N_6404);
and U9056 (N_9056,N_6382,N_5671);
xor U9057 (N_9057,N_5438,N_6537);
and U9058 (N_9058,N_5717,N_5012);
and U9059 (N_9059,N_5522,N_6088);
xnor U9060 (N_9060,N_7361,N_5121);
or U9061 (N_9061,N_7320,N_5487);
or U9062 (N_9062,N_5750,N_5060);
nor U9063 (N_9063,N_6280,N_7213);
and U9064 (N_9064,N_7041,N_5741);
nor U9065 (N_9065,N_5049,N_5267);
or U9066 (N_9066,N_5695,N_5539);
nand U9067 (N_9067,N_6681,N_5308);
xor U9068 (N_9068,N_6564,N_5611);
and U9069 (N_9069,N_7408,N_7293);
or U9070 (N_9070,N_6893,N_5291);
and U9071 (N_9071,N_5188,N_5580);
xor U9072 (N_9072,N_7164,N_5020);
nand U9073 (N_9073,N_5201,N_6571);
and U9074 (N_9074,N_6049,N_7216);
nand U9075 (N_9075,N_6915,N_5904);
or U9076 (N_9076,N_7454,N_7025);
nand U9077 (N_9077,N_5924,N_7361);
nand U9078 (N_9078,N_6355,N_5719);
nand U9079 (N_9079,N_5263,N_5743);
nand U9080 (N_9080,N_6120,N_6362);
nand U9081 (N_9081,N_5180,N_7227);
xor U9082 (N_9082,N_6187,N_5450);
and U9083 (N_9083,N_7324,N_7010);
nand U9084 (N_9084,N_5942,N_5044);
or U9085 (N_9085,N_6918,N_6870);
nand U9086 (N_9086,N_5491,N_5290);
nand U9087 (N_9087,N_6998,N_5544);
or U9088 (N_9088,N_6591,N_5208);
xor U9089 (N_9089,N_5522,N_6993);
nor U9090 (N_9090,N_6270,N_5958);
or U9091 (N_9091,N_7280,N_7111);
xor U9092 (N_9092,N_5638,N_5913);
nand U9093 (N_9093,N_7148,N_7390);
nand U9094 (N_9094,N_6200,N_6684);
and U9095 (N_9095,N_7170,N_6725);
nand U9096 (N_9096,N_6204,N_5859);
and U9097 (N_9097,N_6121,N_6020);
xor U9098 (N_9098,N_5641,N_5091);
or U9099 (N_9099,N_5084,N_5189);
or U9100 (N_9100,N_5774,N_6705);
or U9101 (N_9101,N_7317,N_6129);
and U9102 (N_9102,N_5572,N_6626);
nand U9103 (N_9103,N_6955,N_6062);
and U9104 (N_9104,N_6437,N_6413);
and U9105 (N_9105,N_5973,N_6944);
xor U9106 (N_9106,N_5811,N_5993);
or U9107 (N_9107,N_5575,N_5441);
or U9108 (N_9108,N_6928,N_7492);
xnor U9109 (N_9109,N_7437,N_6067);
and U9110 (N_9110,N_5169,N_7449);
xnor U9111 (N_9111,N_5571,N_5221);
nor U9112 (N_9112,N_5135,N_7326);
nor U9113 (N_9113,N_5738,N_6615);
and U9114 (N_9114,N_6731,N_5969);
nand U9115 (N_9115,N_5945,N_7292);
and U9116 (N_9116,N_5391,N_5143);
and U9117 (N_9117,N_5383,N_7059);
nor U9118 (N_9118,N_5439,N_5188);
xor U9119 (N_9119,N_5941,N_7235);
xor U9120 (N_9120,N_6084,N_5028);
nand U9121 (N_9121,N_7227,N_6320);
nor U9122 (N_9122,N_5458,N_5140);
or U9123 (N_9123,N_6211,N_6400);
and U9124 (N_9124,N_6194,N_5595);
and U9125 (N_9125,N_7368,N_7240);
nand U9126 (N_9126,N_5711,N_6119);
and U9127 (N_9127,N_5391,N_6451);
nand U9128 (N_9128,N_6134,N_5231);
xnor U9129 (N_9129,N_5555,N_5209);
or U9130 (N_9130,N_7251,N_5150);
nor U9131 (N_9131,N_7362,N_5438);
xor U9132 (N_9132,N_5392,N_6872);
or U9133 (N_9133,N_7160,N_5132);
nand U9134 (N_9134,N_5319,N_5569);
or U9135 (N_9135,N_6343,N_6163);
nand U9136 (N_9136,N_5156,N_7314);
or U9137 (N_9137,N_7310,N_6813);
nor U9138 (N_9138,N_6733,N_6582);
nor U9139 (N_9139,N_6176,N_6334);
or U9140 (N_9140,N_7044,N_5871);
and U9141 (N_9141,N_7373,N_5520);
and U9142 (N_9142,N_5906,N_6687);
nor U9143 (N_9143,N_6023,N_7293);
xnor U9144 (N_9144,N_5512,N_5697);
and U9145 (N_9145,N_5828,N_7054);
nand U9146 (N_9146,N_6977,N_5703);
xnor U9147 (N_9147,N_6008,N_7297);
xnor U9148 (N_9148,N_5473,N_7272);
nor U9149 (N_9149,N_5973,N_5215);
nor U9150 (N_9150,N_5214,N_5670);
nor U9151 (N_9151,N_7155,N_6487);
xnor U9152 (N_9152,N_5012,N_5091);
or U9153 (N_9153,N_6228,N_6766);
or U9154 (N_9154,N_5968,N_5535);
nand U9155 (N_9155,N_6271,N_5490);
xor U9156 (N_9156,N_6722,N_5665);
nand U9157 (N_9157,N_5447,N_6318);
or U9158 (N_9158,N_6338,N_5122);
nor U9159 (N_9159,N_5660,N_7302);
nor U9160 (N_9160,N_5592,N_6072);
nor U9161 (N_9161,N_6224,N_7230);
and U9162 (N_9162,N_5894,N_7223);
nand U9163 (N_9163,N_7224,N_7371);
or U9164 (N_9164,N_5399,N_6323);
xor U9165 (N_9165,N_6910,N_5518);
nand U9166 (N_9166,N_6057,N_5835);
nor U9167 (N_9167,N_5526,N_5280);
and U9168 (N_9168,N_6517,N_5303);
or U9169 (N_9169,N_6622,N_6220);
or U9170 (N_9170,N_5914,N_7360);
xnor U9171 (N_9171,N_6304,N_5500);
xnor U9172 (N_9172,N_6870,N_7057);
nor U9173 (N_9173,N_6400,N_5510);
nand U9174 (N_9174,N_6373,N_7343);
or U9175 (N_9175,N_5941,N_6670);
or U9176 (N_9176,N_7024,N_7196);
and U9177 (N_9177,N_6009,N_7412);
nor U9178 (N_9178,N_6985,N_6153);
nor U9179 (N_9179,N_6372,N_6439);
or U9180 (N_9180,N_6921,N_6611);
nand U9181 (N_9181,N_7387,N_5350);
nor U9182 (N_9182,N_6233,N_6824);
or U9183 (N_9183,N_5012,N_6740);
and U9184 (N_9184,N_5546,N_5478);
nor U9185 (N_9185,N_7012,N_5055);
nand U9186 (N_9186,N_5675,N_5955);
nand U9187 (N_9187,N_5304,N_6663);
or U9188 (N_9188,N_7103,N_7476);
or U9189 (N_9189,N_6457,N_6028);
nor U9190 (N_9190,N_5188,N_6029);
nand U9191 (N_9191,N_5732,N_7368);
nor U9192 (N_9192,N_5330,N_7045);
xnor U9193 (N_9193,N_5063,N_5857);
nand U9194 (N_9194,N_6086,N_7415);
xor U9195 (N_9195,N_6057,N_7263);
nor U9196 (N_9196,N_6523,N_6586);
xor U9197 (N_9197,N_5997,N_6501);
nand U9198 (N_9198,N_5714,N_5216);
and U9199 (N_9199,N_6197,N_7219);
xor U9200 (N_9200,N_7215,N_6586);
nand U9201 (N_9201,N_7173,N_7244);
or U9202 (N_9202,N_5727,N_5662);
or U9203 (N_9203,N_6319,N_7436);
xor U9204 (N_9204,N_6066,N_6738);
nor U9205 (N_9205,N_7172,N_6787);
nor U9206 (N_9206,N_5291,N_6319);
xnor U9207 (N_9207,N_6081,N_6390);
and U9208 (N_9208,N_5423,N_7421);
xor U9209 (N_9209,N_5024,N_6899);
nand U9210 (N_9210,N_5562,N_7426);
and U9211 (N_9211,N_5163,N_6268);
and U9212 (N_9212,N_6709,N_7116);
nand U9213 (N_9213,N_5034,N_6835);
nor U9214 (N_9214,N_6723,N_7059);
nor U9215 (N_9215,N_5123,N_6419);
nor U9216 (N_9216,N_7040,N_5917);
xnor U9217 (N_9217,N_6864,N_6485);
and U9218 (N_9218,N_6501,N_6573);
and U9219 (N_9219,N_5997,N_6431);
nand U9220 (N_9220,N_5849,N_7146);
or U9221 (N_9221,N_7264,N_7013);
xor U9222 (N_9222,N_6397,N_5143);
nor U9223 (N_9223,N_6199,N_5680);
xnor U9224 (N_9224,N_6461,N_5374);
xor U9225 (N_9225,N_6066,N_6975);
or U9226 (N_9226,N_6896,N_5796);
and U9227 (N_9227,N_5057,N_7006);
xor U9228 (N_9228,N_5040,N_5000);
xnor U9229 (N_9229,N_5715,N_5259);
xnor U9230 (N_9230,N_5343,N_6226);
or U9231 (N_9231,N_5576,N_7379);
xor U9232 (N_9232,N_5330,N_5920);
nand U9233 (N_9233,N_7428,N_5421);
xnor U9234 (N_9234,N_5363,N_5342);
nand U9235 (N_9235,N_5757,N_5600);
nand U9236 (N_9236,N_7349,N_6508);
and U9237 (N_9237,N_6765,N_5249);
nor U9238 (N_9238,N_5247,N_7089);
nand U9239 (N_9239,N_5887,N_5547);
nor U9240 (N_9240,N_6603,N_6997);
and U9241 (N_9241,N_5462,N_5171);
nor U9242 (N_9242,N_6683,N_5732);
or U9243 (N_9243,N_5738,N_6891);
and U9244 (N_9244,N_6656,N_5246);
or U9245 (N_9245,N_7150,N_6792);
xnor U9246 (N_9246,N_5728,N_6970);
nand U9247 (N_9247,N_5718,N_5457);
nor U9248 (N_9248,N_5658,N_5457);
or U9249 (N_9249,N_6340,N_7056);
nand U9250 (N_9250,N_7440,N_5096);
or U9251 (N_9251,N_5447,N_5421);
or U9252 (N_9252,N_6826,N_7178);
or U9253 (N_9253,N_7418,N_7236);
or U9254 (N_9254,N_6371,N_6949);
nor U9255 (N_9255,N_6460,N_5455);
or U9256 (N_9256,N_7430,N_6717);
nor U9257 (N_9257,N_6278,N_6104);
and U9258 (N_9258,N_7474,N_5611);
and U9259 (N_9259,N_7151,N_7407);
and U9260 (N_9260,N_6529,N_6371);
and U9261 (N_9261,N_6934,N_6949);
or U9262 (N_9262,N_5541,N_6537);
nand U9263 (N_9263,N_7245,N_6226);
nand U9264 (N_9264,N_5905,N_5320);
nand U9265 (N_9265,N_5596,N_6223);
or U9266 (N_9266,N_7102,N_6900);
and U9267 (N_9267,N_6638,N_7406);
or U9268 (N_9268,N_6642,N_7117);
nor U9269 (N_9269,N_7275,N_6156);
nand U9270 (N_9270,N_6847,N_6788);
xnor U9271 (N_9271,N_5981,N_6729);
nand U9272 (N_9272,N_6483,N_7180);
and U9273 (N_9273,N_6289,N_6002);
and U9274 (N_9274,N_5239,N_7035);
nor U9275 (N_9275,N_6695,N_7391);
and U9276 (N_9276,N_7039,N_5065);
and U9277 (N_9277,N_6096,N_6303);
nand U9278 (N_9278,N_6427,N_6467);
or U9279 (N_9279,N_5232,N_5125);
nor U9280 (N_9280,N_5613,N_6505);
and U9281 (N_9281,N_5249,N_5991);
xnor U9282 (N_9282,N_5595,N_6717);
xor U9283 (N_9283,N_6705,N_5526);
and U9284 (N_9284,N_5683,N_5053);
nor U9285 (N_9285,N_7274,N_7026);
or U9286 (N_9286,N_6975,N_5341);
and U9287 (N_9287,N_7212,N_5136);
xnor U9288 (N_9288,N_7383,N_5241);
or U9289 (N_9289,N_7392,N_5258);
or U9290 (N_9290,N_5304,N_5582);
nand U9291 (N_9291,N_6274,N_5953);
or U9292 (N_9292,N_6015,N_7149);
or U9293 (N_9293,N_6388,N_7268);
nand U9294 (N_9294,N_5893,N_6209);
nand U9295 (N_9295,N_5807,N_7000);
and U9296 (N_9296,N_5392,N_6945);
or U9297 (N_9297,N_5363,N_5929);
and U9298 (N_9298,N_5164,N_6759);
nor U9299 (N_9299,N_6015,N_7206);
xnor U9300 (N_9300,N_5943,N_6961);
nor U9301 (N_9301,N_6655,N_6059);
xor U9302 (N_9302,N_6995,N_5084);
nor U9303 (N_9303,N_6897,N_5796);
or U9304 (N_9304,N_5810,N_6151);
nand U9305 (N_9305,N_5140,N_6064);
xnor U9306 (N_9306,N_6930,N_5462);
xnor U9307 (N_9307,N_7151,N_7114);
nor U9308 (N_9308,N_6648,N_7462);
nor U9309 (N_9309,N_6696,N_6371);
nand U9310 (N_9310,N_5714,N_6158);
or U9311 (N_9311,N_6205,N_6253);
and U9312 (N_9312,N_7479,N_5315);
or U9313 (N_9313,N_6872,N_7123);
or U9314 (N_9314,N_5094,N_6736);
or U9315 (N_9315,N_7409,N_7452);
or U9316 (N_9316,N_5671,N_6564);
xnor U9317 (N_9317,N_5380,N_6726);
xor U9318 (N_9318,N_7080,N_6571);
nor U9319 (N_9319,N_6968,N_6580);
nand U9320 (N_9320,N_5248,N_6678);
or U9321 (N_9321,N_6224,N_7469);
nor U9322 (N_9322,N_7353,N_6397);
nor U9323 (N_9323,N_6852,N_6844);
nand U9324 (N_9324,N_5835,N_7365);
xnor U9325 (N_9325,N_7266,N_5975);
nor U9326 (N_9326,N_7078,N_6243);
nand U9327 (N_9327,N_5754,N_7328);
xnor U9328 (N_9328,N_7431,N_6613);
or U9329 (N_9329,N_5906,N_5177);
or U9330 (N_9330,N_7243,N_7451);
xor U9331 (N_9331,N_5452,N_5861);
nand U9332 (N_9332,N_6147,N_7161);
or U9333 (N_9333,N_5275,N_6466);
nor U9334 (N_9334,N_7406,N_6129);
or U9335 (N_9335,N_7022,N_5218);
and U9336 (N_9336,N_6861,N_6110);
and U9337 (N_9337,N_5671,N_5221);
nor U9338 (N_9338,N_7068,N_6353);
nor U9339 (N_9339,N_5876,N_6015);
and U9340 (N_9340,N_7275,N_6310);
nand U9341 (N_9341,N_6769,N_5298);
xnor U9342 (N_9342,N_7287,N_6121);
nor U9343 (N_9343,N_5060,N_5645);
or U9344 (N_9344,N_6001,N_6739);
nor U9345 (N_9345,N_6023,N_6972);
and U9346 (N_9346,N_5069,N_7425);
and U9347 (N_9347,N_7031,N_7250);
nor U9348 (N_9348,N_6501,N_5687);
xnor U9349 (N_9349,N_6274,N_5429);
xor U9350 (N_9350,N_5991,N_6064);
nor U9351 (N_9351,N_5279,N_7413);
nand U9352 (N_9352,N_6639,N_6550);
nor U9353 (N_9353,N_6589,N_5677);
nand U9354 (N_9354,N_6200,N_5574);
and U9355 (N_9355,N_5593,N_7044);
xor U9356 (N_9356,N_5071,N_6427);
xor U9357 (N_9357,N_5892,N_6949);
nor U9358 (N_9358,N_5293,N_6432);
xnor U9359 (N_9359,N_6806,N_6060);
and U9360 (N_9360,N_7106,N_5139);
xor U9361 (N_9361,N_7286,N_5218);
nor U9362 (N_9362,N_6204,N_7078);
xnor U9363 (N_9363,N_5733,N_7077);
or U9364 (N_9364,N_7036,N_7237);
and U9365 (N_9365,N_6082,N_6073);
or U9366 (N_9366,N_5493,N_6401);
xor U9367 (N_9367,N_7326,N_6270);
or U9368 (N_9368,N_5641,N_7070);
nand U9369 (N_9369,N_6839,N_6410);
nor U9370 (N_9370,N_6083,N_6595);
nor U9371 (N_9371,N_7129,N_6380);
or U9372 (N_9372,N_5590,N_5228);
and U9373 (N_9373,N_6988,N_5620);
nor U9374 (N_9374,N_6977,N_5070);
and U9375 (N_9375,N_6055,N_5065);
xor U9376 (N_9376,N_5313,N_6881);
xor U9377 (N_9377,N_5050,N_6133);
nand U9378 (N_9378,N_5052,N_6861);
xor U9379 (N_9379,N_5260,N_7296);
xnor U9380 (N_9380,N_6125,N_6447);
or U9381 (N_9381,N_6593,N_5313);
nand U9382 (N_9382,N_7005,N_5990);
nand U9383 (N_9383,N_5865,N_6248);
or U9384 (N_9384,N_6272,N_5950);
xnor U9385 (N_9385,N_5442,N_5832);
or U9386 (N_9386,N_5117,N_6344);
nor U9387 (N_9387,N_5750,N_6383);
or U9388 (N_9388,N_6253,N_5465);
xnor U9389 (N_9389,N_6539,N_5418);
nor U9390 (N_9390,N_7222,N_6087);
nand U9391 (N_9391,N_7339,N_6793);
or U9392 (N_9392,N_5577,N_5022);
nand U9393 (N_9393,N_5170,N_5898);
xor U9394 (N_9394,N_5820,N_5829);
xor U9395 (N_9395,N_5107,N_6621);
or U9396 (N_9396,N_6804,N_5294);
xnor U9397 (N_9397,N_5875,N_7047);
and U9398 (N_9398,N_6245,N_5071);
nand U9399 (N_9399,N_7215,N_6157);
xnor U9400 (N_9400,N_7153,N_7174);
nor U9401 (N_9401,N_5564,N_7402);
nor U9402 (N_9402,N_7476,N_6156);
nand U9403 (N_9403,N_5875,N_7474);
nand U9404 (N_9404,N_5106,N_6792);
nor U9405 (N_9405,N_6115,N_5676);
nand U9406 (N_9406,N_6002,N_6438);
nand U9407 (N_9407,N_6795,N_7252);
nand U9408 (N_9408,N_5561,N_5169);
xor U9409 (N_9409,N_7182,N_5156);
and U9410 (N_9410,N_6181,N_5736);
xnor U9411 (N_9411,N_7339,N_6027);
nor U9412 (N_9412,N_6380,N_6253);
nand U9413 (N_9413,N_6395,N_5698);
or U9414 (N_9414,N_5501,N_6078);
xor U9415 (N_9415,N_6886,N_7304);
nor U9416 (N_9416,N_6981,N_7354);
nor U9417 (N_9417,N_6405,N_6572);
xor U9418 (N_9418,N_6721,N_6418);
or U9419 (N_9419,N_5608,N_7247);
nor U9420 (N_9420,N_6240,N_7439);
nor U9421 (N_9421,N_5403,N_5134);
nor U9422 (N_9422,N_5666,N_5238);
xor U9423 (N_9423,N_7022,N_6475);
nor U9424 (N_9424,N_5495,N_7187);
xor U9425 (N_9425,N_5630,N_7422);
or U9426 (N_9426,N_7466,N_7022);
and U9427 (N_9427,N_5186,N_6666);
and U9428 (N_9428,N_7235,N_5189);
and U9429 (N_9429,N_5363,N_6009);
or U9430 (N_9430,N_6786,N_5338);
and U9431 (N_9431,N_6970,N_7252);
or U9432 (N_9432,N_7277,N_5039);
xnor U9433 (N_9433,N_7234,N_5077);
nand U9434 (N_9434,N_5807,N_6827);
nor U9435 (N_9435,N_5844,N_6933);
nand U9436 (N_9436,N_7378,N_6028);
or U9437 (N_9437,N_7356,N_5490);
nor U9438 (N_9438,N_7324,N_5471);
and U9439 (N_9439,N_6702,N_7096);
and U9440 (N_9440,N_5685,N_6340);
or U9441 (N_9441,N_5820,N_7399);
nand U9442 (N_9442,N_5386,N_5885);
nand U9443 (N_9443,N_6216,N_6223);
nand U9444 (N_9444,N_5928,N_5736);
xor U9445 (N_9445,N_6620,N_7342);
or U9446 (N_9446,N_5988,N_7432);
xor U9447 (N_9447,N_5265,N_6156);
or U9448 (N_9448,N_6665,N_7191);
xor U9449 (N_9449,N_6688,N_5467);
or U9450 (N_9450,N_5989,N_5895);
xor U9451 (N_9451,N_6084,N_5464);
nand U9452 (N_9452,N_6525,N_6864);
or U9453 (N_9453,N_6369,N_5745);
and U9454 (N_9454,N_5704,N_6124);
xor U9455 (N_9455,N_6620,N_6091);
nor U9456 (N_9456,N_5854,N_6856);
or U9457 (N_9457,N_7138,N_5193);
nor U9458 (N_9458,N_6039,N_5086);
nand U9459 (N_9459,N_5758,N_7060);
and U9460 (N_9460,N_5245,N_7105);
nor U9461 (N_9461,N_5035,N_6680);
or U9462 (N_9462,N_5031,N_6491);
xnor U9463 (N_9463,N_6653,N_5202);
nor U9464 (N_9464,N_6763,N_5696);
nand U9465 (N_9465,N_5501,N_7436);
nand U9466 (N_9466,N_7321,N_7141);
and U9467 (N_9467,N_5547,N_6536);
and U9468 (N_9468,N_6117,N_7467);
and U9469 (N_9469,N_6486,N_7031);
or U9470 (N_9470,N_7202,N_6844);
nor U9471 (N_9471,N_5226,N_7227);
xor U9472 (N_9472,N_6945,N_5234);
and U9473 (N_9473,N_5823,N_6581);
or U9474 (N_9474,N_7137,N_6670);
xor U9475 (N_9475,N_7072,N_5069);
or U9476 (N_9476,N_7450,N_6888);
nand U9477 (N_9477,N_6620,N_5115);
nand U9478 (N_9478,N_7066,N_6523);
and U9479 (N_9479,N_6210,N_6913);
xnor U9480 (N_9480,N_6006,N_6962);
or U9481 (N_9481,N_5879,N_5926);
and U9482 (N_9482,N_6474,N_6265);
or U9483 (N_9483,N_6186,N_7186);
nor U9484 (N_9484,N_5328,N_6075);
nor U9485 (N_9485,N_6819,N_7232);
nor U9486 (N_9486,N_5111,N_6838);
nor U9487 (N_9487,N_5994,N_6289);
nor U9488 (N_9488,N_5707,N_6314);
and U9489 (N_9489,N_5272,N_6923);
or U9490 (N_9490,N_6894,N_5736);
nand U9491 (N_9491,N_7234,N_6704);
or U9492 (N_9492,N_6634,N_5408);
and U9493 (N_9493,N_7428,N_6526);
xor U9494 (N_9494,N_5435,N_6407);
nand U9495 (N_9495,N_6881,N_6739);
or U9496 (N_9496,N_6142,N_5901);
and U9497 (N_9497,N_5375,N_7201);
nand U9498 (N_9498,N_6205,N_5543);
or U9499 (N_9499,N_5382,N_5735);
and U9500 (N_9500,N_6429,N_7202);
nand U9501 (N_9501,N_5258,N_7068);
xnor U9502 (N_9502,N_6139,N_6068);
xnor U9503 (N_9503,N_5164,N_5557);
or U9504 (N_9504,N_6777,N_6474);
or U9505 (N_9505,N_6543,N_5565);
nand U9506 (N_9506,N_5908,N_7122);
nor U9507 (N_9507,N_5619,N_5000);
xor U9508 (N_9508,N_5273,N_5087);
nand U9509 (N_9509,N_7070,N_7146);
or U9510 (N_9510,N_5763,N_7268);
or U9511 (N_9511,N_5317,N_7188);
and U9512 (N_9512,N_7348,N_6859);
and U9513 (N_9513,N_6745,N_7435);
nand U9514 (N_9514,N_7385,N_6782);
nand U9515 (N_9515,N_5627,N_7100);
nor U9516 (N_9516,N_5121,N_6130);
or U9517 (N_9517,N_5180,N_7017);
xnor U9518 (N_9518,N_5012,N_6996);
nor U9519 (N_9519,N_6156,N_5478);
or U9520 (N_9520,N_6197,N_7140);
nor U9521 (N_9521,N_5029,N_5722);
or U9522 (N_9522,N_5572,N_6274);
xor U9523 (N_9523,N_6247,N_6239);
and U9524 (N_9524,N_6758,N_6824);
nor U9525 (N_9525,N_6896,N_6046);
nand U9526 (N_9526,N_5490,N_5333);
xnor U9527 (N_9527,N_6364,N_6102);
xor U9528 (N_9528,N_7233,N_5065);
and U9529 (N_9529,N_6304,N_6640);
or U9530 (N_9530,N_6275,N_6629);
xnor U9531 (N_9531,N_5210,N_6014);
nor U9532 (N_9532,N_5098,N_6830);
xnor U9533 (N_9533,N_6675,N_7266);
or U9534 (N_9534,N_7254,N_6883);
or U9535 (N_9535,N_6353,N_5112);
xor U9536 (N_9536,N_7316,N_6490);
xnor U9537 (N_9537,N_7220,N_5639);
nand U9538 (N_9538,N_5990,N_7316);
nand U9539 (N_9539,N_5196,N_6239);
nor U9540 (N_9540,N_5344,N_6506);
and U9541 (N_9541,N_5987,N_5403);
and U9542 (N_9542,N_5804,N_5542);
nand U9543 (N_9543,N_7337,N_5100);
and U9544 (N_9544,N_5035,N_5498);
nor U9545 (N_9545,N_5431,N_7206);
or U9546 (N_9546,N_5678,N_5653);
nand U9547 (N_9547,N_6300,N_6864);
nand U9548 (N_9548,N_5206,N_6431);
xor U9549 (N_9549,N_6703,N_6606);
nor U9550 (N_9550,N_6775,N_5913);
or U9551 (N_9551,N_6131,N_5932);
nand U9552 (N_9552,N_6797,N_6570);
nand U9553 (N_9553,N_6764,N_6486);
nand U9554 (N_9554,N_6120,N_5592);
or U9555 (N_9555,N_7117,N_6979);
nor U9556 (N_9556,N_5072,N_7175);
xor U9557 (N_9557,N_5018,N_7344);
or U9558 (N_9558,N_5266,N_6710);
nor U9559 (N_9559,N_6739,N_7354);
and U9560 (N_9560,N_7127,N_5527);
or U9561 (N_9561,N_5285,N_7192);
nand U9562 (N_9562,N_6373,N_6986);
or U9563 (N_9563,N_5566,N_6961);
or U9564 (N_9564,N_5119,N_6674);
or U9565 (N_9565,N_5904,N_6044);
and U9566 (N_9566,N_5802,N_5186);
nand U9567 (N_9567,N_5829,N_5929);
nand U9568 (N_9568,N_5861,N_5311);
nand U9569 (N_9569,N_5169,N_5522);
xor U9570 (N_9570,N_6777,N_6344);
nor U9571 (N_9571,N_6276,N_5066);
xor U9572 (N_9572,N_7070,N_6037);
xnor U9573 (N_9573,N_6960,N_6602);
or U9574 (N_9574,N_5472,N_6503);
nand U9575 (N_9575,N_7428,N_7471);
or U9576 (N_9576,N_7363,N_6593);
nor U9577 (N_9577,N_6032,N_6175);
nor U9578 (N_9578,N_6988,N_6583);
or U9579 (N_9579,N_5752,N_5179);
nand U9580 (N_9580,N_5013,N_5904);
nand U9581 (N_9581,N_6038,N_5794);
or U9582 (N_9582,N_5446,N_7353);
nor U9583 (N_9583,N_7419,N_6844);
and U9584 (N_9584,N_5923,N_7320);
or U9585 (N_9585,N_6944,N_6836);
xor U9586 (N_9586,N_5027,N_6066);
xnor U9587 (N_9587,N_5991,N_6866);
xnor U9588 (N_9588,N_6732,N_7410);
nand U9589 (N_9589,N_7464,N_5875);
nor U9590 (N_9590,N_5737,N_7489);
nor U9591 (N_9591,N_5260,N_5966);
nor U9592 (N_9592,N_5103,N_5106);
and U9593 (N_9593,N_5084,N_5843);
nor U9594 (N_9594,N_5618,N_5858);
xor U9595 (N_9595,N_7324,N_6041);
and U9596 (N_9596,N_6234,N_5441);
and U9597 (N_9597,N_5865,N_6609);
and U9598 (N_9598,N_7252,N_5140);
and U9599 (N_9599,N_6523,N_6538);
xor U9600 (N_9600,N_6457,N_7409);
xor U9601 (N_9601,N_6934,N_5929);
xnor U9602 (N_9602,N_5513,N_5213);
nand U9603 (N_9603,N_6288,N_5419);
xor U9604 (N_9604,N_6845,N_5810);
nor U9605 (N_9605,N_6479,N_6834);
and U9606 (N_9606,N_7102,N_5964);
nand U9607 (N_9607,N_5507,N_7364);
or U9608 (N_9608,N_5220,N_6387);
nor U9609 (N_9609,N_6055,N_6582);
or U9610 (N_9610,N_5754,N_6320);
or U9611 (N_9611,N_7453,N_6263);
xor U9612 (N_9612,N_7229,N_5766);
nor U9613 (N_9613,N_6883,N_6447);
nor U9614 (N_9614,N_5842,N_5065);
or U9615 (N_9615,N_6175,N_5642);
and U9616 (N_9616,N_5008,N_7288);
and U9617 (N_9617,N_5019,N_5949);
nand U9618 (N_9618,N_7116,N_5733);
xor U9619 (N_9619,N_6041,N_6687);
xor U9620 (N_9620,N_6668,N_7014);
nand U9621 (N_9621,N_7423,N_5544);
nand U9622 (N_9622,N_7274,N_5636);
xnor U9623 (N_9623,N_6500,N_6821);
and U9624 (N_9624,N_5690,N_5218);
and U9625 (N_9625,N_6578,N_5042);
xor U9626 (N_9626,N_5445,N_6541);
nand U9627 (N_9627,N_6914,N_6226);
xor U9628 (N_9628,N_5402,N_6223);
nand U9629 (N_9629,N_7327,N_5025);
xnor U9630 (N_9630,N_6494,N_7304);
nor U9631 (N_9631,N_6191,N_5134);
nor U9632 (N_9632,N_5500,N_5956);
nand U9633 (N_9633,N_5383,N_6108);
and U9634 (N_9634,N_7005,N_5732);
xnor U9635 (N_9635,N_5915,N_5053);
nand U9636 (N_9636,N_7256,N_6769);
nand U9637 (N_9637,N_6232,N_7196);
xor U9638 (N_9638,N_6494,N_6253);
or U9639 (N_9639,N_7352,N_7048);
nand U9640 (N_9640,N_6644,N_7237);
nand U9641 (N_9641,N_5293,N_5694);
nand U9642 (N_9642,N_5357,N_5416);
xor U9643 (N_9643,N_6137,N_6483);
nand U9644 (N_9644,N_6336,N_5426);
and U9645 (N_9645,N_5229,N_7134);
xnor U9646 (N_9646,N_5974,N_6729);
and U9647 (N_9647,N_7474,N_7195);
nor U9648 (N_9648,N_6871,N_5059);
or U9649 (N_9649,N_6897,N_5615);
nand U9650 (N_9650,N_6751,N_6621);
xor U9651 (N_9651,N_7341,N_5129);
and U9652 (N_9652,N_6866,N_7279);
or U9653 (N_9653,N_6605,N_5234);
and U9654 (N_9654,N_5448,N_5092);
or U9655 (N_9655,N_6796,N_6165);
or U9656 (N_9656,N_5464,N_6517);
or U9657 (N_9657,N_5345,N_6499);
nand U9658 (N_9658,N_6361,N_6450);
and U9659 (N_9659,N_6189,N_6484);
and U9660 (N_9660,N_5526,N_7327);
nand U9661 (N_9661,N_6718,N_5379);
or U9662 (N_9662,N_6248,N_6215);
and U9663 (N_9663,N_6290,N_5704);
and U9664 (N_9664,N_7359,N_6218);
nand U9665 (N_9665,N_6611,N_7332);
nor U9666 (N_9666,N_6079,N_7415);
nand U9667 (N_9667,N_5038,N_5599);
xnor U9668 (N_9668,N_5529,N_5580);
nand U9669 (N_9669,N_6605,N_5728);
and U9670 (N_9670,N_6543,N_5661);
nand U9671 (N_9671,N_6634,N_5070);
xor U9672 (N_9672,N_6330,N_7387);
nand U9673 (N_9673,N_6473,N_6044);
xor U9674 (N_9674,N_7144,N_6149);
or U9675 (N_9675,N_6423,N_6541);
nor U9676 (N_9676,N_5433,N_5611);
and U9677 (N_9677,N_6451,N_5169);
nand U9678 (N_9678,N_6627,N_6361);
or U9679 (N_9679,N_6778,N_5983);
xor U9680 (N_9680,N_6129,N_6039);
and U9681 (N_9681,N_6583,N_7368);
nand U9682 (N_9682,N_6684,N_7495);
or U9683 (N_9683,N_5738,N_5369);
nor U9684 (N_9684,N_6104,N_5360);
nand U9685 (N_9685,N_7208,N_6984);
and U9686 (N_9686,N_6929,N_7271);
or U9687 (N_9687,N_5773,N_5603);
xnor U9688 (N_9688,N_6911,N_5051);
nand U9689 (N_9689,N_5391,N_6719);
and U9690 (N_9690,N_5899,N_7107);
nand U9691 (N_9691,N_5278,N_6213);
nor U9692 (N_9692,N_7491,N_6860);
or U9693 (N_9693,N_6276,N_5103);
or U9694 (N_9694,N_5808,N_5084);
nand U9695 (N_9695,N_5046,N_7297);
xor U9696 (N_9696,N_5504,N_5848);
nor U9697 (N_9697,N_7385,N_7357);
or U9698 (N_9698,N_6483,N_7021);
nand U9699 (N_9699,N_5648,N_5124);
xor U9700 (N_9700,N_6260,N_6399);
xnor U9701 (N_9701,N_5427,N_5754);
nand U9702 (N_9702,N_5365,N_7284);
nand U9703 (N_9703,N_5040,N_5547);
nand U9704 (N_9704,N_6176,N_5756);
xor U9705 (N_9705,N_6568,N_6042);
nand U9706 (N_9706,N_5911,N_6730);
or U9707 (N_9707,N_5335,N_6159);
or U9708 (N_9708,N_5318,N_6316);
xnor U9709 (N_9709,N_5233,N_6950);
xor U9710 (N_9710,N_6468,N_6138);
or U9711 (N_9711,N_6963,N_6780);
nand U9712 (N_9712,N_6401,N_7204);
nand U9713 (N_9713,N_6722,N_6902);
nand U9714 (N_9714,N_7400,N_6649);
or U9715 (N_9715,N_6620,N_6572);
xor U9716 (N_9716,N_5955,N_5731);
xnor U9717 (N_9717,N_5605,N_7065);
xnor U9718 (N_9718,N_5502,N_5029);
or U9719 (N_9719,N_5848,N_5523);
xnor U9720 (N_9720,N_7385,N_5586);
or U9721 (N_9721,N_7486,N_6617);
nand U9722 (N_9722,N_5828,N_6079);
and U9723 (N_9723,N_5973,N_5837);
nand U9724 (N_9724,N_5518,N_5272);
nor U9725 (N_9725,N_6888,N_5316);
nor U9726 (N_9726,N_5921,N_6826);
xnor U9727 (N_9727,N_7174,N_5388);
and U9728 (N_9728,N_5903,N_6170);
and U9729 (N_9729,N_7117,N_7067);
nor U9730 (N_9730,N_6326,N_6674);
xnor U9731 (N_9731,N_5620,N_5646);
and U9732 (N_9732,N_7215,N_6739);
xor U9733 (N_9733,N_5037,N_5609);
or U9734 (N_9734,N_6153,N_5139);
xnor U9735 (N_9735,N_6519,N_6198);
xnor U9736 (N_9736,N_6922,N_6284);
xor U9737 (N_9737,N_5634,N_5853);
and U9738 (N_9738,N_6766,N_6018);
xnor U9739 (N_9739,N_5955,N_5068);
nor U9740 (N_9740,N_5932,N_6466);
nor U9741 (N_9741,N_7060,N_7181);
and U9742 (N_9742,N_6649,N_7214);
nand U9743 (N_9743,N_6652,N_6577);
nor U9744 (N_9744,N_6638,N_6964);
and U9745 (N_9745,N_6673,N_5694);
and U9746 (N_9746,N_6804,N_7401);
or U9747 (N_9747,N_5684,N_7481);
nand U9748 (N_9748,N_5521,N_5150);
xnor U9749 (N_9749,N_5443,N_5779);
or U9750 (N_9750,N_5813,N_7321);
and U9751 (N_9751,N_6684,N_7483);
or U9752 (N_9752,N_7339,N_5635);
nand U9753 (N_9753,N_5405,N_5095);
xor U9754 (N_9754,N_5394,N_6718);
nor U9755 (N_9755,N_6309,N_7365);
or U9756 (N_9756,N_5219,N_5825);
nor U9757 (N_9757,N_6476,N_6612);
or U9758 (N_9758,N_6730,N_6336);
xor U9759 (N_9759,N_6098,N_7343);
or U9760 (N_9760,N_5462,N_6701);
nor U9761 (N_9761,N_7078,N_7081);
nor U9762 (N_9762,N_7387,N_6442);
nor U9763 (N_9763,N_6962,N_5444);
and U9764 (N_9764,N_5864,N_7263);
xnor U9765 (N_9765,N_5078,N_5864);
nor U9766 (N_9766,N_6047,N_5079);
nand U9767 (N_9767,N_6272,N_6927);
or U9768 (N_9768,N_5154,N_5689);
or U9769 (N_9769,N_5579,N_5053);
and U9770 (N_9770,N_6422,N_6678);
or U9771 (N_9771,N_7479,N_7214);
xnor U9772 (N_9772,N_7482,N_6356);
xnor U9773 (N_9773,N_5139,N_6934);
nor U9774 (N_9774,N_5232,N_5265);
xor U9775 (N_9775,N_5549,N_5440);
and U9776 (N_9776,N_6413,N_7486);
nor U9777 (N_9777,N_7116,N_6665);
nor U9778 (N_9778,N_6651,N_6229);
nand U9779 (N_9779,N_6559,N_6125);
or U9780 (N_9780,N_5996,N_6797);
xor U9781 (N_9781,N_7481,N_5776);
or U9782 (N_9782,N_7035,N_5841);
or U9783 (N_9783,N_6996,N_7358);
or U9784 (N_9784,N_6765,N_7298);
and U9785 (N_9785,N_5258,N_5564);
nand U9786 (N_9786,N_7203,N_6738);
nand U9787 (N_9787,N_6995,N_7322);
or U9788 (N_9788,N_7423,N_6373);
or U9789 (N_9789,N_6316,N_6570);
nand U9790 (N_9790,N_6434,N_5966);
nand U9791 (N_9791,N_6049,N_7110);
nor U9792 (N_9792,N_5089,N_5305);
nor U9793 (N_9793,N_5084,N_6165);
xnor U9794 (N_9794,N_7232,N_5704);
nand U9795 (N_9795,N_7216,N_7115);
xnor U9796 (N_9796,N_5681,N_5011);
and U9797 (N_9797,N_5234,N_5939);
xnor U9798 (N_9798,N_7343,N_6585);
and U9799 (N_9799,N_7232,N_6548);
nor U9800 (N_9800,N_7364,N_5383);
and U9801 (N_9801,N_5610,N_6616);
xnor U9802 (N_9802,N_7465,N_5057);
nor U9803 (N_9803,N_7462,N_6428);
xor U9804 (N_9804,N_6945,N_7464);
xnor U9805 (N_9805,N_7215,N_7224);
nor U9806 (N_9806,N_5764,N_7374);
xnor U9807 (N_9807,N_5133,N_5434);
nor U9808 (N_9808,N_6450,N_6847);
xnor U9809 (N_9809,N_5121,N_5680);
and U9810 (N_9810,N_6553,N_6023);
and U9811 (N_9811,N_7360,N_6952);
nor U9812 (N_9812,N_5207,N_7044);
nand U9813 (N_9813,N_5554,N_5325);
or U9814 (N_9814,N_6151,N_6277);
and U9815 (N_9815,N_7404,N_6481);
xor U9816 (N_9816,N_6092,N_7404);
nor U9817 (N_9817,N_6135,N_5575);
and U9818 (N_9818,N_5012,N_5751);
nand U9819 (N_9819,N_7178,N_6010);
nand U9820 (N_9820,N_6565,N_5533);
and U9821 (N_9821,N_6755,N_6562);
xnor U9822 (N_9822,N_7474,N_6537);
and U9823 (N_9823,N_7038,N_5460);
and U9824 (N_9824,N_7343,N_6638);
nand U9825 (N_9825,N_5805,N_6225);
xnor U9826 (N_9826,N_6389,N_5631);
nand U9827 (N_9827,N_5762,N_6986);
nand U9828 (N_9828,N_5892,N_5484);
xnor U9829 (N_9829,N_5189,N_7040);
xor U9830 (N_9830,N_6933,N_6724);
nand U9831 (N_9831,N_7383,N_6622);
xor U9832 (N_9832,N_7153,N_6933);
nor U9833 (N_9833,N_6260,N_6160);
xor U9834 (N_9834,N_6085,N_5650);
nand U9835 (N_9835,N_5193,N_6731);
and U9836 (N_9836,N_5011,N_7104);
nor U9837 (N_9837,N_6839,N_7423);
and U9838 (N_9838,N_7087,N_5864);
xor U9839 (N_9839,N_6700,N_5685);
or U9840 (N_9840,N_7339,N_6594);
and U9841 (N_9841,N_5897,N_7327);
xnor U9842 (N_9842,N_5152,N_5272);
and U9843 (N_9843,N_6900,N_6998);
nand U9844 (N_9844,N_5820,N_6121);
nor U9845 (N_9845,N_7476,N_6856);
nand U9846 (N_9846,N_6063,N_5659);
nor U9847 (N_9847,N_7468,N_6337);
nand U9848 (N_9848,N_5298,N_7208);
and U9849 (N_9849,N_5814,N_6843);
xor U9850 (N_9850,N_6621,N_7482);
nor U9851 (N_9851,N_5083,N_5314);
and U9852 (N_9852,N_5515,N_5350);
nor U9853 (N_9853,N_5797,N_5923);
and U9854 (N_9854,N_6876,N_7030);
nand U9855 (N_9855,N_5758,N_7083);
nor U9856 (N_9856,N_7393,N_7087);
nand U9857 (N_9857,N_7027,N_5222);
xnor U9858 (N_9858,N_6339,N_7262);
nand U9859 (N_9859,N_6657,N_6335);
nor U9860 (N_9860,N_5154,N_6295);
or U9861 (N_9861,N_6068,N_6101);
xnor U9862 (N_9862,N_6393,N_7002);
nand U9863 (N_9863,N_6304,N_7479);
nand U9864 (N_9864,N_6916,N_5876);
nor U9865 (N_9865,N_7072,N_5724);
xor U9866 (N_9866,N_6100,N_7169);
xnor U9867 (N_9867,N_5191,N_5481);
xor U9868 (N_9868,N_5411,N_7011);
nor U9869 (N_9869,N_5885,N_5189);
nand U9870 (N_9870,N_6622,N_7217);
xor U9871 (N_9871,N_5693,N_5935);
nand U9872 (N_9872,N_6777,N_6421);
nor U9873 (N_9873,N_5630,N_7144);
and U9874 (N_9874,N_6965,N_7080);
xnor U9875 (N_9875,N_5565,N_6219);
and U9876 (N_9876,N_5871,N_5340);
xor U9877 (N_9877,N_6252,N_5373);
nand U9878 (N_9878,N_7472,N_6537);
nor U9879 (N_9879,N_5745,N_5513);
nand U9880 (N_9880,N_6285,N_5955);
or U9881 (N_9881,N_5438,N_6921);
and U9882 (N_9882,N_5389,N_5820);
xor U9883 (N_9883,N_6266,N_6702);
xnor U9884 (N_9884,N_5632,N_6213);
xnor U9885 (N_9885,N_5030,N_6742);
or U9886 (N_9886,N_7131,N_6052);
xor U9887 (N_9887,N_7202,N_7014);
xnor U9888 (N_9888,N_6260,N_6154);
nand U9889 (N_9889,N_5916,N_7445);
and U9890 (N_9890,N_6178,N_5071);
xor U9891 (N_9891,N_5030,N_5157);
nor U9892 (N_9892,N_5756,N_7198);
xnor U9893 (N_9893,N_6287,N_5828);
xor U9894 (N_9894,N_6307,N_5021);
and U9895 (N_9895,N_5226,N_7150);
and U9896 (N_9896,N_7099,N_5323);
or U9897 (N_9897,N_7410,N_5560);
xor U9898 (N_9898,N_5006,N_7256);
or U9899 (N_9899,N_5226,N_6688);
nor U9900 (N_9900,N_6373,N_6987);
and U9901 (N_9901,N_5556,N_6822);
or U9902 (N_9902,N_7172,N_6123);
nand U9903 (N_9903,N_6229,N_6041);
and U9904 (N_9904,N_7308,N_5619);
or U9905 (N_9905,N_5544,N_6570);
or U9906 (N_9906,N_5504,N_5108);
or U9907 (N_9907,N_5944,N_7100);
or U9908 (N_9908,N_6144,N_7093);
nand U9909 (N_9909,N_6922,N_6642);
and U9910 (N_9910,N_5322,N_5989);
xor U9911 (N_9911,N_6144,N_5123);
and U9912 (N_9912,N_6638,N_5493);
nand U9913 (N_9913,N_5546,N_5940);
xnor U9914 (N_9914,N_7013,N_6440);
nor U9915 (N_9915,N_7095,N_6311);
nand U9916 (N_9916,N_5160,N_6725);
nor U9917 (N_9917,N_6619,N_5529);
or U9918 (N_9918,N_5287,N_5274);
nand U9919 (N_9919,N_7353,N_6889);
or U9920 (N_9920,N_5626,N_6855);
nor U9921 (N_9921,N_6935,N_7216);
nor U9922 (N_9922,N_5254,N_7285);
nor U9923 (N_9923,N_5988,N_6366);
xor U9924 (N_9924,N_6157,N_6374);
xnor U9925 (N_9925,N_6680,N_7251);
or U9926 (N_9926,N_5232,N_6904);
xnor U9927 (N_9927,N_5669,N_6766);
nand U9928 (N_9928,N_6368,N_5083);
nand U9929 (N_9929,N_5260,N_5549);
and U9930 (N_9930,N_5556,N_7034);
and U9931 (N_9931,N_5825,N_5710);
and U9932 (N_9932,N_5099,N_6805);
nand U9933 (N_9933,N_5323,N_5696);
nor U9934 (N_9934,N_6745,N_6722);
nand U9935 (N_9935,N_5257,N_7339);
xnor U9936 (N_9936,N_6029,N_5258);
or U9937 (N_9937,N_6686,N_6406);
or U9938 (N_9938,N_6178,N_6740);
nor U9939 (N_9939,N_5971,N_6640);
and U9940 (N_9940,N_7029,N_6861);
nor U9941 (N_9941,N_6033,N_6207);
xnor U9942 (N_9942,N_6875,N_6107);
and U9943 (N_9943,N_6578,N_5549);
nor U9944 (N_9944,N_5102,N_7112);
nand U9945 (N_9945,N_5289,N_7285);
xnor U9946 (N_9946,N_6847,N_5729);
nor U9947 (N_9947,N_6340,N_5162);
and U9948 (N_9948,N_6017,N_5492);
xnor U9949 (N_9949,N_5207,N_7190);
nor U9950 (N_9950,N_7455,N_7490);
nand U9951 (N_9951,N_6053,N_5286);
and U9952 (N_9952,N_5173,N_6474);
nand U9953 (N_9953,N_5235,N_6155);
and U9954 (N_9954,N_7044,N_5063);
nand U9955 (N_9955,N_6175,N_6998);
nor U9956 (N_9956,N_5264,N_6357);
nor U9957 (N_9957,N_6838,N_5426);
xor U9958 (N_9958,N_7341,N_5976);
nor U9959 (N_9959,N_6206,N_7289);
or U9960 (N_9960,N_6910,N_5499);
or U9961 (N_9961,N_6348,N_5226);
and U9962 (N_9962,N_6245,N_7461);
and U9963 (N_9963,N_5950,N_6640);
nor U9964 (N_9964,N_6302,N_5975);
nand U9965 (N_9965,N_6528,N_6257);
and U9966 (N_9966,N_5389,N_7445);
xnor U9967 (N_9967,N_7176,N_5444);
xor U9968 (N_9968,N_5002,N_6866);
and U9969 (N_9969,N_6772,N_7124);
xor U9970 (N_9970,N_6649,N_5553);
nor U9971 (N_9971,N_5152,N_5361);
and U9972 (N_9972,N_6633,N_6764);
nand U9973 (N_9973,N_7171,N_6468);
xor U9974 (N_9974,N_6222,N_5603);
and U9975 (N_9975,N_5659,N_7197);
and U9976 (N_9976,N_5444,N_6093);
or U9977 (N_9977,N_6787,N_7075);
xor U9978 (N_9978,N_5130,N_5174);
xor U9979 (N_9979,N_6918,N_6075);
nor U9980 (N_9980,N_6283,N_5444);
nor U9981 (N_9981,N_7040,N_6834);
or U9982 (N_9982,N_5915,N_5505);
nor U9983 (N_9983,N_6689,N_5334);
or U9984 (N_9984,N_7232,N_7382);
and U9985 (N_9985,N_5277,N_5101);
or U9986 (N_9986,N_5692,N_6722);
or U9987 (N_9987,N_5810,N_6240);
nor U9988 (N_9988,N_5203,N_5955);
or U9989 (N_9989,N_5671,N_5433);
xor U9990 (N_9990,N_5393,N_6477);
nand U9991 (N_9991,N_6762,N_5028);
nor U9992 (N_9992,N_6293,N_7470);
xnor U9993 (N_9993,N_6636,N_6391);
or U9994 (N_9994,N_7125,N_6793);
xor U9995 (N_9995,N_6429,N_7409);
xnor U9996 (N_9996,N_5879,N_7473);
xnor U9997 (N_9997,N_7224,N_7193);
and U9998 (N_9998,N_6008,N_6828);
nand U9999 (N_9999,N_6759,N_6972);
xnor U10000 (N_10000,N_9912,N_8501);
nand U10001 (N_10001,N_7997,N_9109);
nor U10002 (N_10002,N_7787,N_9091);
and U10003 (N_10003,N_8897,N_8484);
nand U10004 (N_10004,N_7732,N_9512);
and U10005 (N_10005,N_8673,N_7859);
or U10006 (N_10006,N_8202,N_8298);
xnor U10007 (N_10007,N_7579,N_9907);
and U10008 (N_10008,N_9225,N_9351);
nand U10009 (N_10009,N_9662,N_8831);
nor U10010 (N_10010,N_7613,N_8913);
xor U10011 (N_10011,N_9743,N_9003);
and U10012 (N_10012,N_8013,N_8381);
nand U10013 (N_10013,N_7687,N_8768);
nand U10014 (N_10014,N_9058,N_7805);
nor U10015 (N_10015,N_7561,N_7546);
nand U10016 (N_10016,N_9827,N_9390);
nand U10017 (N_10017,N_8372,N_8490);
xor U10018 (N_10018,N_9839,N_9468);
xnor U10019 (N_10019,N_9239,N_7910);
and U10020 (N_10020,N_9127,N_9207);
or U10021 (N_10021,N_9153,N_7933);
xor U10022 (N_10022,N_7500,N_9307);
nor U10023 (N_10023,N_8564,N_7689);
nand U10024 (N_10024,N_9466,N_8903);
xnor U10025 (N_10025,N_8854,N_9000);
nor U10026 (N_10026,N_8129,N_9240);
and U10027 (N_10027,N_8241,N_9728);
and U10028 (N_10028,N_9038,N_9476);
and U10029 (N_10029,N_7651,N_7605);
nand U10030 (N_10030,N_8520,N_8819);
nand U10031 (N_10031,N_9876,N_8261);
nand U10032 (N_10032,N_8603,N_8009);
or U10033 (N_10033,N_9546,N_9253);
xnor U10034 (N_10034,N_8042,N_9009);
xor U10035 (N_10035,N_9126,N_8999);
or U10036 (N_10036,N_8223,N_7534);
nor U10037 (N_10037,N_9623,N_7768);
xnor U10038 (N_10038,N_9522,N_7939);
and U10039 (N_10039,N_9864,N_8857);
nand U10040 (N_10040,N_9167,N_7666);
or U10041 (N_10041,N_9588,N_8655);
and U10042 (N_10042,N_8405,N_9228);
nor U10043 (N_10043,N_9917,N_9227);
xnor U10044 (N_10044,N_7517,N_9120);
or U10045 (N_10045,N_9551,N_8196);
and U10046 (N_10046,N_7681,N_9834);
nor U10047 (N_10047,N_7807,N_7956);
nor U10048 (N_10048,N_8328,N_9041);
or U10049 (N_10049,N_8273,N_9299);
and U10050 (N_10050,N_8380,N_8324);
and U10051 (N_10051,N_9104,N_9659);
xor U10052 (N_10052,N_7583,N_9475);
and U10053 (N_10053,N_8580,N_7931);
or U10054 (N_10054,N_8868,N_9331);
and U10055 (N_10055,N_8001,N_9828);
xnor U10056 (N_10056,N_9704,N_7536);
nand U10057 (N_10057,N_7657,N_9204);
nor U10058 (N_10058,N_9703,N_9825);
nand U10059 (N_10059,N_8724,N_8134);
nor U10060 (N_10060,N_8537,N_9031);
nand U10061 (N_10061,N_8739,N_7801);
and U10062 (N_10062,N_9134,N_8199);
xnor U10063 (N_10063,N_9820,N_9333);
xor U10064 (N_10064,N_9628,N_8278);
xnor U10065 (N_10065,N_9050,N_7620);
and U10066 (N_10066,N_8522,N_8299);
nor U10067 (N_10067,N_7922,N_8975);
and U10068 (N_10068,N_7983,N_8974);
and U10069 (N_10069,N_8708,N_8253);
nor U10070 (N_10070,N_9328,N_7909);
and U10071 (N_10071,N_8647,N_8720);
xor U10072 (N_10072,N_8763,N_9015);
xor U10073 (N_10073,N_9151,N_8275);
nand U10074 (N_10074,N_9183,N_9283);
nand U10075 (N_10075,N_7659,N_8234);
or U10076 (N_10076,N_8876,N_9309);
nor U10077 (N_10077,N_7547,N_9192);
xor U10078 (N_10078,N_7692,N_9173);
xor U10079 (N_10079,N_9098,N_9556);
nor U10080 (N_10080,N_9918,N_9800);
nor U10081 (N_10081,N_8164,N_8075);
xnor U10082 (N_10082,N_8599,N_7593);
nor U10083 (N_10083,N_9482,N_7861);
and U10084 (N_10084,N_9814,N_8945);
or U10085 (N_10085,N_9906,N_8117);
nand U10086 (N_10086,N_7580,N_8576);
and U10087 (N_10087,N_9570,N_7758);
nor U10088 (N_10088,N_9561,N_9099);
xor U10089 (N_10089,N_7566,N_8590);
and U10090 (N_10090,N_8400,N_9181);
or U10091 (N_10091,N_7836,N_9100);
xor U10092 (N_10092,N_8296,N_8227);
xnor U10093 (N_10093,N_8753,N_7646);
xor U10094 (N_10094,N_9729,N_9089);
or U10095 (N_10095,N_8806,N_9625);
xnor U10096 (N_10096,N_9999,N_9550);
and U10097 (N_10097,N_9016,N_9544);
or U10098 (N_10098,N_9784,N_8841);
or U10099 (N_10099,N_9238,N_9245);
or U10100 (N_10100,N_7788,N_8973);
or U10101 (N_10101,N_9298,N_7835);
and U10102 (N_10102,N_9187,N_8459);
nor U10103 (N_10103,N_7540,N_8939);
nor U10104 (N_10104,N_8243,N_8587);
xor U10105 (N_10105,N_9319,N_7789);
or U10106 (N_10106,N_9140,N_9866);
and U10107 (N_10107,N_9286,N_7890);
nor U10108 (N_10108,N_8748,N_8169);
and U10109 (N_10109,N_7844,N_9036);
xnor U10110 (N_10110,N_8991,N_7893);
nor U10111 (N_10111,N_7706,N_8715);
or U10112 (N_10112,N_8718,N_7718);
xor U10113 (N_10113,N_9592,N_7809);
nand U10114 (N_10114,N_7746,N_8055);
or U10115 (N_10115,N_8048,N_9752);
xnor U10116 (N_10116,N_9944,N_9744);
and U10117 (N_10117,N_8650,N_8450);
nor U10118 (N_10118,N_8597,N_8112);
xnor U10119 (N_10119,N_9485,N_7565);
xor U10120 (N_10120,N_8823,N_8224);
or U10121 (N_10121,N_9809,N_9053);
nor U10122 (N_10122,N_8376,N_8280);
xor U10123 (N_10123,N_9255,N_8466);
nor U10124 (N_10124,N_9219,N_8835);
and U10125 (N_10125,N_7631,N_8730);
and U10126 (N_10126,N_8967,N_8014);
nand U10127 (N_10127,N_8249,N_9869);
and U10128 (N_10128,N_9765,N_9209);
nor U10129 (N_10129,N_9710,N_8270);
and U10130 (N_10130,N_8548,N_9933);
nand U10131 (N_10131,N_8060,N_8552);
nor U10132 (N_10132,N_8267,N_8526);
xnor U10133 (N_10133,N_9223,N_8363);
and U10134 (N_10134,N_9982,N_9817);
nand U10135 (N_10135,N_8547,N_8953);
and U10136 (N_10136,N_9017,N_8632);
nand U10137 (N_10137,N_8978,N_7920);
xor U10138 (N_10138,N_8961,N_8761);
xor U10139 (N_10139,N_8302,N_7812);
xor U10140 (N_10140,N_9101,N_9997);
xor U10141 (N_10141,N_7735,N_8678);
nor U10142 (N_10142,N_9273,N_8127);
or U10143 (N_10143,N_9367,N_8439);
xnor U10144 (N_10144,N_8561,N_9885);
xnor U10145 (N_10145,N_7914,N_7919);
or U10146 (N_10146,N_8078,N_8852);
and U10147 (N_10147,N_9123,N_9121);
nand U10148 (N_10148,N_7766,N_8346);
or U10149 (N_10149,N_9762,N_9521);
nand U10150 (N_10150,N_7610,N_8116);
nor U10151 (N_10151,N_8383,N_8741);
nor U10152 (N_10152,N_8263,N_7906);
nor U10153 (N_10153,N_7690,N_7796);
and U10154 (N_10154,N_8707,N_7526);
or U10155 (N_10155,N_7656,N_8932);
xor U10156 (N_10156,N_8710,N_8044);
nand U10157 (N_10157,N_8779,N_8331);
xnor U10158 (N_10158,N_9667,N_9547);
nor U10159 (N_10159,N_9614,N_8879);
nor U10160 (N_10160,N_8881,N_8122);
nand U10161 (N_10161,N_9062,N_7503);
nor U10162 (N_10162,N_8290,N_7682);
nor U10163 (N_10163,N_8456,N_9783);
or U10164 (N_10164,N_8690,N_9111);
nand U10165 (N_10165,N_9585,N_8562);
nor U10166 (N_10166,N_8107,N_8816);
and U10167 (N_10167,N_8900,N_7652);
or U10168 (N_10168,N_7717,N_8524);
nor U10169 (N_10169,N_8133,N_9177);
nand U10170 (N_10170,N_7992,N_8722);
and U10171 (N_10171,N_8410,N_8478);
xor U10172 (N_10172,N_9481,N_8142);
and U10173 (N_10173,N_8794,N_8181);
nor U10174 (N_10174,N_9088,N_8110);
or U10175 (N_10175,N_9741,N_9757);
xor U10176 (N_10176,N_8307,N_8737);
xor U10177 (N_10177,N_9108,N_9862);
nand U10178 (N_10178,N_9086,N_8336);
nand U10179 (N_10179,N_8862,N_8152);
or U10180 (N_10180,N_8361,N_9459);
nor U10181 (N_10181,N_8432,N_8856);
nor U10182 (N_10182,N_8515,N_8322);
nand U10183 (N_10183,N_8658,N_8230);
nor U10184 (N_10184,N_7609,N_8842);
and U10185 (N_10185,N_8440,N_8514);
nor U10186 (N_10186,N_9833,N_9405);
and U10187 (N_10187,N_7592,N_7637);
xnor U10188 (N_10188,N_9664,N_8265);
or U10189 (N_10189,N_7867,N_7697);
nor U10190 (N_10190,N_9158,N_7808);
xnor U10191 (N_10191,N_7753,N_8613);
xnor U10192 (N_10192,N_9665,N_8866);
xor U10193 (N_10193,N_8005,N_8283);
nand U10194 (N_10194,N_9985,N_9334);
nand U10195 (N_10195,N_9148,N_9575);
or U10196 (N_10196,N_9449,N_8742);
nand U10197 (N_10197,N_9023,N_9868);
or U10198 (N_10198,N_7994,N_9169);
or U10199 (N_10199,N_8624,N_8000);
nand U10200 (N_10200,N_9190,N_7888);
xor U10201 (N_10201,N_9622,N_7509);
or U10202 (N_10202,N_9727,N_9927);
and U10203 (N_10203,N_7964,N_9479);
and U10204 (N_10204,N_8586,N_9528);
or U10205 (N_10205,N_9454,N_8684);
nand U10206 (N_10206,N_8480,N_9430);
or U10207 (N_10207,N_8211,N_8512);
nor U10208 (N_10208,N_9066,N_8143);
nand U10209 (N_10209,N_9683,N_8915);
or U10210 (N_10210,N_9034,N_9505);
and U10211 (N_10211,N_8053,N_7870);
xor U10212 (N_10212,N_7792,N_7774);
or U10213 (N_10213,N_7771,N_9714);
and U10214 (N_10214,N_9684,N_9188);
nand U10215 (N_10215,N_8834,N_8814);
xor U10216 (N_10216,N_9007,N_8846);
nor U10217 (N_10217,N_9737,N_8538);
nand U10218 (N_10218,N_9423,N_9543);
or U10219 (N_10219,N_7621,N_7701);
or U10220 (N_10220,N_7538,N_9692);
xnor U10221 (N_10221,N_7639,N_8616);
and U10222 (N_10222,N_9358,N_8661);
nor U10223 (N_10223,N_9749,N_8717);
or U10224 (N_10224,N_9632,N_7733);
xor U10225 (N_10225,N_8565,N_7567);
xnor U10226 (N_10226,N_9144,N_8104);
nand U10227 (N_10227,N_9175,N_7991);
and U10228 (N_10228,N_8539,N_9365);
or U10229 (N_10229,N_9832,N_8061);
and U10230 (N_10230,N_7853,N_9563);
nor U10231 (N_10231,N_9558,N_9473);
nand U10232 (N_10232,N_9962,N_9750);
or U10233 (N_10233,N_8904,N_9890);
nor U10234 (N_10234,N_7935,N_8063);
nand U10235 (N_10235,N_8445,N_9940);
or U10236 (N_10236,N_9029,N_9600);
and U10237 (N_10237,N_7982,N_9527);
or U10238 (N_10238,N_8186,N_9271);
nand U10239 (N_10239,N_9152,N_7705);
nor U10240 (N_10240,N_8289,N_8451);
and U10241 (N_10241,N_7677,N_8917);
xor U10242 (N_10242,N_8385,N_7679);
nor U10243 (N_10243,N_8706,N_8443);
nand U10244 (N_10244,N_9707,N_8529);
nor U10245 (N_10245,N_9332,N_9325);
and U10246 (N_10246,N_9445,N_9576);
and U10247 (N_10247,N_8506,N_8228);
or U10248 (N_10248,N_7924,N_7751);
nand U10249 (N_10249,N_8923,N_9461);
xnor U10250 (N_10250,N_8485,N_8210);
and U10251 (N_10251,N_9656,N_8756);
or U10252 (N_10252,N_7976,N_9769);
xnor U10253 (N_10253,N_8884,N_8309);
nor U10254 (N_10254,N_8146,N_9421);
nor U10255 (N_10255,N_8402,N_9165);
and U10256 (N_10256,N_9612,N_8882);
xor U10257 (N_10257,N_8019,N_7762);
or U10258 (N_10258,N_9560,N_9191);
or U10259 (N_10259,N_8920,N_8219);
xnor U10260 (N_10260,N_8065,N_9026);
and U10261 (N_10261,N_8193,N_9577);
and U10262 (N_10262,N_8303,N_8551);
xnor U10263 (N_10263,N_7944,N_8032);
or U10264 (N_10264,N_8138,N_8209);
and U10265 (N_10265,N_9530,N_8132);
xor U10266 (N_10266,N_8339,N_7930);
nand U10267 (N_10267,N_9198,N_7529);
and U10268 (N_10268,N_7668,N_9384);
nor U10269 (N_10269,N_8969,N_9392);
xor U10270 (N_10270,N_9807,N_8621);
xnor U10271 (N_10271,N_9156,N_7996);
xnor U10272 (N_10272,N_8214,N_9269);
or U10273 (N_10273,N_7628,N_8293);
or U10274 (N_10274,N_9439,N_8928);
nand U10275 (N_10275,N_8012,N_7847);
nand U10276 (N_10276,N_8885,N_9206);
and U10277 (N_10277,N_8676,N_8271);
or U10278 (N_10278,N_8037,N_7806);
or U10279 (N_10279,N_9082,N_9128);
or U10280 (N_10280,N_8574,N_7780);
or U10281 (N_10281,N_9259,N_9263);
and U10282 (N_10282,N_9571,N_8015);
nand U10283 (N_10283,N_9617,N_7804);
nor U10284 (N_10284,N_9778,N_7672);
nand U10285 (N_10285,N_8113,N_9400);
nand U10286 (N_10286,N_7785,N_7726);
nand U10287 (N_10287,N_9730,N_9138);
nand U10288 (N_10288,N_9396,N_8509);
nand U10289 (N_10289,N_7872,N_9777);
nor U10290 (N_10290,N_8617,N_9386);
nand U10291 (N_10291,N_9624,N_8709);
nand U10292 (N_10292,N_8752,N_8062);
and U10293 (N_10293,N_8906,N_9873);
xor U10294 (N_10294,N_8926,N_9077);
nand U10295 (N_10295,N_8471,N_9201);
nand U10296 (N_10296,N_7745,N_8148);
nand U10297 (N_10297,N_9019,N_9792);
and U10298 (N_10298,N_8773,N_7654);
xnor U10299 (N_10299,N_8891,N_9257);
nand U10300 (N_10300,N_9774,N_9626);
or U10301 (N_10301,N_9135,N_7721);
and U10302 (N_10302,N_8072,N_8180);
nand U10303 (N_10303,N_7731,N_7863);
and U10304 (N_10304,N_8631,N_7527);
or U10305 (N_10305,N_9806,N_7649);
and U10306 (N_10306,N_9831,N_9302);
and U10307 (N_10307,N_7967,N_9539);
nor U10308 (N_10308,N_9432,N_8629);
nor U10309 (N_10309,N_8163,N_7819);
xor U10310 (N_10310,N_9764,N_8384);
or U10311 (N_10311,N_7747,N_9433);
nand U10312 (N_10312,N_8156,N_9160);
nand U10313 (N_10313,N_8924,N_8971);
and U10314 (N_10314,N_8908,N_7840);
and U10315 (N_10315,N_9318,N_7937);
xor U10316 (N_10316,N_9695,N_7838);
or U10317 (N_10317,N_8101,N_9984);
xor U10318 (N_10318,N_9420,N_9346);
nand U10319 (N_10319,N_8855,N_9678);
xnor U10320 (N_10320,N_9568,N_8546);
or U10321 (N_10321,N_9211,N_8927);
and U10322 (N_10322,N_7653,N_8284);
nand U10323 (N_10323,N_9602,N_8326);
and U10324 (N_10324,N_7736,N_9079);
or U10325 (N_10325,N_9686,N_8337);
or U10326 (N_10326,N_7802,N_8304);
and U10327 (N_10327,N_8568,N_7894);
nand U10328 (N_10328,N_7798,N_8236);
or U10329 (N_10329,N_9083,N_9176);
xor U10330 (N_10330,N_9105,N_9132);
and U10331 (N_10331,N_7782,N_8231);
xnor U10332 (N_10332,N_8994,N_7588);
or U10333 (N_10333,N_9797,N_8663);
xor U10334 (N_10334,N_7722,N_9642);
or U10335 (N_10335,N_9477,N_8183);
nand U10336 (N_10336,N_7643,N_9895);
and U10337 (N_10337,N_9103,N_9262);
and U10338 (N_10338,N_9295,N_8544);
or U10339 (N_10339,N_8849,N_9119);
xnor U10340 (N_10340,N_8081,N_7522);
or U10341 (N_10341,N_8525,N_8245);
nor U10342 (N_10342,N_9047,N_8308);
nand U10343 (N_10343,N_9660,N_9964);
or U10344 (N_10344,N_7683,N_8497);
nand U10345 (N_10345,N_7704,N_9141);
nor U10346 (N_10346,N_8919,N_7908);
or U10347 (N_10347,N_8644,N_9450);
nor U10348 (N_10348,N_9620,N_9993);
nand U10349 (N_10349,N_8258,N_8332);
and U10350 (N_10350,N_9587,N_9357);
or U10351 (N_10351,N_8511,N_9954);
nor U10352 (N_10352,N_9483,N_9829);
or U10353 (N_10353,N_8626,N_7978);
xor U10354 (N_10354,N_8206,N_8770);
or U10355 (N_10355,N_8046,N_7946);
nand U10356 (N_10356,N_8418,N_9013);
and U10357 (N_10357,N_7525,N_7658);
nor U10358 (N_10358,N_8345,N_8185);
nor U10359 (N_10359,N_9702,N_7663);
or U10360 (N_10360,N_9818,N_9314);
nand U10361 (N_10361,N_8195,N_8825);
nand U10362 (N_10362,N_9781,N_8725);
or U10363 (N_10363,N_8171,N_7988);
and U10364 (N_10364,N_8287,N_9166);
xnor U10365 (N_10365,N_8494,N_8909);
nand U10366 (N_10366,N_8233,N_9159);
or U10367 (N_10367,N_8672,N_9495);
xor U10368 (N_10368,N_9028,N_8373);
nand U10369 (N_10369,N_8878,N_7511);
xnor U10370 (N_10370,N_9846,N_8281);
nor U10371 (N_10371,N_8649,N_9874);
nor U10372 (N_10372,N_9478,N_8184);
and U10373 (N_10373,N_9785,N_9589);
or U10374 (N_10374,N_9130,N_8022);
xnor U10375 (N_10375,N_9672,N_7549);
and U10376 (N_10376,N_9677,N_9643);
nor U10377 (N_10377,N_9706,N_7869);
xnor U10378 (N_10378,N_8479,N_8802);
nand U10379 (N_10379,N_8396,N_8697);
xor U10380 (N_10380,N_9203,N_7505);
and U10381 (N_10381,N_9854,N_9972);
or U10382 (N_10382,N_7817,N_7737);
or U10383 (N_10383,N_9756,N_9248);
nand U10384 (N_10384,N_7767,N_7923);
nor U10385 (N_10385,N_8775,N_8795);
and U10386 (N_10386,N_9812,N_9001);
nand U10387 (N_10387,N_8205,N_8172);
nor U10388 (N_10388,N_9768,N_9621);
nor U10389 (N_10389,N_7744,N_9639);
nor U10390 (N_10390,N_8301,N_8056);
or U10391 (N_10391,N_8563,N_9075);
and U10392 (N_10392,N_9360,N_9920);
or U10393 (N_10393,N_8623,N_9627);
and U10394 (N_10394,N_8865,N_8870);
nand U10395 (N_10395,N_8108,N_8517);
nor U10396 (N_10396,N_9317,N_8203);
or U10397 (N_10397,N_7951,N_7851);
nor U10398 (N_10398,N_9233,N_7776);
nand U10399 (N_10399,N_9518,N_9913);
or U10400 (N_10400,N_9995,N_7986);
or U10401 (N_10401,N_8957,N_8811);
nand U10402 (N_10402,N_7947,N_8887);
nor U10403 (N_10403,N_9429,N_8996);
nand U10404 (N_10404,N_9929,N_8784);
nor U10405 (N_10405,N_7501,N_9287);
or U10406 (N_10406,N_9139,N_8872);
nand U10407 (N_10407,N_8793,N_9451);
nand U10408 (N_10408,N_8378,N_8235);
and U10409 (N_10409,N_9986,N_9310);
nand U10410 (N_10410,N_7596,N_9071);
nand U10411 (N_10411,N_7600,N_8064);
and U10412 (N_10412,N_9265,N_7794);
nand U10413 (N_10413,N_8011,N_9422);
and U10414 (N_10414,N_8719,N_9763);
or U10415 (N_10415,N_9112,N_9841);
and U10416 (N_10416,N_7715,N_8131);
and U10417 (N_10417,N_9282,N_8733);
nand U10418 (N_10418,N_8782,N_9060);
and U10419 (N_10419,N_8701,N_9548);
and U10420 (N_10420,N_9244,N_7950);
nand U10421 (N_10421,N_7590,N_9676);
nand U10422 (N_10422,N_9958,N_7848);
and U10423 (N_10423,N_9005,N_9393);
xor U10424 (N_10424,N_9798,N_8686);
and U10425 (N_10425,N_8740,N_8502);
nor U10426 (N_10426,N_9410,N_9935);
nand U10427 (N_10427,N_7917,N_7587);
nor U10428 (N_10428,N_9409,N_9796);
xnor U10429 (N_10429,N_7612,N_7626);
and U10430 (N_10430,N_8197,N_9535);
or U10431 (N_10431,N_7913,N_8434);
nand U10432 (N_10432,N_8902,N_7729);
nand U10433 (N_10433,N_9124,N_8914);
and U10434 (N_10434,N_8791,N_9214);
xor U10435 (N_10435,N_8455,N_7925);
nor U10436 (N_10436,N_7678,N_9754);
or U10437 (N_10437,N_7691,N_9049);
and U10438 (N_10438,N_8468,N_8716);
or U10439 (N_10439,N_8907,N_7712);
nor U10440 (N_10440,N_9960,N_8179);
and U10441 (N_10441,N_7577,N_9855);
nor U10442 (N_10442,N_8334,N_9277);
and U10443 (N_10443,N_9337,N_7942);
or U10444 (N_10444,N_9524,N_8404);
xor U10445 (N_10445,N_8160,N_9447);
nand U10446 (N_10446,N_8832,N_9251);
or U10447 (N_10447,N_8329,N_9145);
nand U10448 (N_10448,N_8333,N_9971);
and U10449 (N_10449,N_8094,N_9462);
nand U10450 (N_10450,N_8300,N_9883);
or U10451 (N_10451,N_8992,N_9306);
nor U10452 (N_10452,N_7823,N_8170);
nand U10453 (N_10453,N_8579,N_7660);
and U10454 (N_10454,N_8705,N_7734);
nand U10455 (N_10455,N_9603,N_9252);
xor U10456 (N_10456,N_8419,N_9301);
nor U10457 (N_10457,N_9849,N_8041);
nand U10458 (N_10458,N_9303,N_8150);
or U10459 (N_10459,N_7603,N_7816);
xnor U10460 (N_10460,N_8130,N_8682);
nor U10461 (N_10461,N_9553,N_8428);
or U10462 (N_10462,N_8747,N_9965);
nand U10463 (N_10463,N_8609,N_7750);
nor U10464 (N_10464,N_9994,N_9387);
xnor U10465 (N_10465,N_9107,N_7959);
nor U10466 (N_10466,N_9691,N_8662);
and U10467 (N_10467,N_8883,N_9065);
nand U10468 (N_10468,N_9407,N_8216);
and U10469 (N_10469,N_8685,N_8294);
and U10470 (N_10470,N_9669,N_9968);
nor U10471 (N_10471,N_8154,N_9200);
nand U10472 (N_10472,N_9237,N_8344);
or U10473 (N_10473,N_8038,N_9713);
nor U10474 (N_10474,N_8125,N_9315);
nor U10475 (N_10475,N_9709,N_9736);
xnor U10476 (N_10476,N_8377,N_7961);
nand U10477 (N_10477,N_8366,N_8394);
xnor U10478 (N_10478,N_9569,N_9969);
nand U10479 (N_10479,N_7968,N_7573);
nand U10480 (N_10480,N_8429,N_9196);
nand U10481 (N_10481,N_8452,N_9415);
or U10482 (N_10482,N_8764,N_8247);
xor U10483 (N_10483,N_9292,N_9385);
nor U10484 (N_10484,N_9537,N_8407);
and U10485 (N_10485,N_8826,N_9637);
nor U10486 (N_10486,N_8731,N_7829);
xnor U10487 (N_10487,N_8036,N_9352);
or U10488 (N_10488,N_7855,N_9012);
xor U10489 (N_10489,N_9094,N_8962);
or U10490 (N_10490,N_7685,N_9261);
nand U10491 (N_10491,N_9725,N_7601);
or U10492 (N_10492,N_7535,N_9919);
or U10493 (N_10493,N_8315,N_7606);
xnor U10494 (N_10494,N_8279,N_7900);
and U10495 (N_10495,N_8873,N_8353);
and U10496 (N_10496,N_9526,N_8892);
and U10497 (N_10497,N_7645,N_9411);
nor U10498 (N_10498,N_9871,N_9342);
xnor U10499 (N_10499,N_8364,N_9157);
or U10500 (N_10500,N_9296,N_7514);
nand U10501 (N_10501,N_7519,N_9035);
or U10502 (N_10502,N_9776,N_8578);
xnor U10503 (N_10503,N_9250,N_7882);
xnor U10504 (N_10504,N_9990,N_7647);
or U10505 (N_10505,N_8805,N_8476);
xor U10506 (N_10506,N_8843,N_9220);
or U10507 (N_10507,N_9989,N_9705);
nand U10508 (N_10508,N_7852,N_8734);
or U10509 (N_10509,N_7757,N_9063);
nand U10510 (N_10510,N_8910,N_9129);
nor U10511 (N_10511,N_9398,N_8467);
xnor U10512 (N_10512,N_9746,N_9117);
nor U10513 (N_10513,N_8930,N_8099);
nor U10514 (N_10514,N_8583,N_7597);
or U10515 (N_10515,N_9020,N_8571);
or U10516 (N_10516,N_8596,N_8808);
nand U10517 (N_10517,N_7568,N_9372);
xnor U10518 (N_10518,N_8584,N_8824);
and U10519 (N_10519,N_9241,N_7544);
or U10520 (N_10520,N_9195,N_8713);
and U10521 (N_10521,N_8933,N_8021);
nand U10522 (N_10522,N_8847,N_9279);
nor U10523 (N_10523,N_9782,N_9523);
nor U10524 (N_10524,N_9801,N_8598);
and U10525 (N_10525,N_8141,N_9164);
nor U10526 (N_10526,N_7634,N_8807);
nor U10527 (N_10527,N_8664,N_8341);
nor U10528 (N_10528,N_8749,N_9647);
or U10529 (N_10529,N_9330,N_7531);
nand U10530 (N_10530,N_8358,N_8213);
and U10531 (N_10531,N_9666,N_9980);
nand U10532 (N_10532,N_9480,N_9037);
and U10533 (N_10533,N_9087,N_8120);
or U10534 (N_10534,N_7885,N_8395);
nor U10535 (N_10535,N_9930,N_8040);
nor U10536 (N_10536,N_8204,N_9516);
nand U10537 (N_10537,N_7877,N_7826);
nor U10538 (N_10538,N_8155,N_9668);
nor U10539 (N_10539,N_8457,N_9453);
xnor U10540 (N_10540,N_8695,N_7604);
and U10541 (N_10541,N_8257,N_9538);
xnor U10542 (N_10542,N_8692,N_7554);
xor U10543 (N_10543,N_7858,N_8951);
xor U10544 (N_10544,N_8536,N_7553);
xor U10545 (N_10545,N_9819,N_9413);
xnor U10546 (N_10546,N_9803,N_7707);
or U10547 (N_10547,N_7739,N_7843);
nand U10548 (N_10548,N_8894,N_8943);
xnor U10549 (N_10549,N_9943,N_7781);
or U10550 (N_10550,N_7741,N_9574);
and U10551 (N_10551,N_8946,N_9114);
nand U10552 (N_10552,N_8533,N_9006);
xor U10553 (N_10553,N_9947,N_8774);
or U10554 (N_10554,N_9578,N_7875);
nor U10555 (N_10555,N_7857,N_7576);
nor U10556 (N_10556,N_8620,N_8666);
and U10557 (N_10557,N_8026,N_8277);
or U10558 (N_10558,N_9349,N_8157);
xnor U10559 (N_10559,N_8829,N_9742);
xnor U10560 (N_10560,N_9708,N_9434);
xor U10561 (N_10561,N_9904,N_7694);
or U10562 (N_10562,N_9021,N_7644);
xor U10563 (N_10563,N_9805,N_9284);
or U10564 (N_10564,N_8863,N_9324);
nor U10565 (N_10565,N_9565,N_7614);
or U10566 (N_10566,N_9716,N_9671);
or U10567 (N_10567,N_8528,N_8988);
nand U10568 (N_10568,N_7695,N_9064);
nand U10569 (N_10569,N_7578,N_7640);
or U10570 (N_10570,N_9533,N_7602);
nor U10571 (N_10571,N_9996,N_8033);
nand U10572 (N_10572,N_9366,N_9653);
xnor U10573 (N_10573,N_8771,N_9567);
nor U10574 (N_10574,N_9418,N_8374);
or U10575 (N_10575,N_9787,N_9654);
xnor U10576 (N_10576,N_9232,N_7918);
xnor U10577 (N_10577,N_8665,N_9813);
nor U10578 (N_10578,N_7599,N_9564);
nand U10579 (N_10579,N_7815,N_9168);
xor U10580 (N_10580,N_7724,N_9300);
or U10581 (N_10581,N_8595,N_9040);
nand U10582 (N_10582,N_9618,N_9278);
or U10583 (N_10583,N_9953,N_8858);
or U10584 (N_10584,N_9773,N_8413);
xor U10585 (N_10585,N_7892,N_8393);
or U10586 (N_10586,N_8637,N_8675);
xor U10587 (N_10587,N_8192,N_7676);
and U10588 (N_10588,N_7969,N_9745);
or U10589 (N_10589,N_9888,N_9507);
xor U10590 (N_10590,N_8636,N_7963);
or U10591 (N_10591,N_9657,N_8505);
nand U10592 (N_10592,N_8607,N_8618);
or U10593 (N_10593,N_7638,N_8838);
nand U10594 (N_10594,N_9597,N_7784);
nand U10595 (N_10595,N_9373,N_7770);
or U10596 (N_10596,N_7675,N_8425);
xnor U10597 (N_10597,N_7990,N_9902);
or U10598 (N_10598,N_9428,N_7849);
nor U10599 (N_10599,N_8642,N_7876);
xnor U10600 (N_10600,N_9840,N_9967);
and U10601 (N_10601,N_8898,N_7508);
and U10602 (N_10602,N_7513,N_8751);
and U10603 (N_10603,N_9815,N_9931);
xor U10604 (N_10604,N_8567,N_8610);
or U10605 (N_10605,N_9948,N_9397);
nand U10606 (N_10606,N_9679,N_9224);
or U10607 (N_10607,N_7756,N_8557);
and U10608 (N_10608,N_7545,N_9051);
or U10609 (N_10609,N_7763,N_9027);
nand U10610 (N_10610,N_7830,N_8758);
and U10611 (N_10611,N_9733,N_9802);
and U10612 (N_10612,N_8274,N_8895);
nand U10613 (N_10613,N_8194,N_9755);
nor U10614 (N_10614,N_9879,N_8177);
xnor U10615 (N_10615,N_8354,N_9504);
nand U10616 (N_10616,N_9208,N_8487);
nor U10617 (N_10617,N_8700,N_8674);
xor U10618 (N_10618,N_9808,N_9922);
or U10619 (N_10619,N_7623,N_9008);
and U10620 (N_10620,N_9681,N_9486);
xor U10621 (N_10621,N_9863,N_7995);
and U10622 (N_10622,N_7674,N_9090);
nand U10623 (N_10623,N_7510,N_8769);
nand U10624 (N_10624,N_7555,N_8365);
and U10625 (N_10625,N_8516,N_7552);
nand U10626 (N_10626,N_8698,N_9934);
or U10627 (N_10627,N_7921,N_8688);
xor U10628 (N_10628,N_7803,N_9186);
and U10629 (N_10629,N_8508,N_9881);
nand U10630 (N_10630,N_7824,N_7708);
xor U10631 (N_10631,N_8426,N_8781);
or U10632 (N_10632,N_9116,N_7749);
nor U10633 (N_10633,N_8349,N_8444);
and U10634 (N_10634,N_9857,N_8639);
and U10635 (N_10635,N_7516,N_9514);
or U10636 (N_10636,N_9059,N_8935);
or U10637 (N_10637,N_8260,N_9983);
nand U10638 (N_10638,N_7854,N_8820);
nor U10639 (N_10639,N_8783,N_7860);
and U10640 (N_10640,N_7518,N_9611);
and U10641 (N_10641,N_8059,N_9723);
nand U10642 (N_10642,N_7928,N_8523);
or U10643 (N_10643,N_7629,N_7720);
nand U10644 (N_10644,N_9363,N_9966);
or U10645 (N_10645,N_9189,N_7879);
xor U10646 (N_10646,N_9844,N_8934);
nand U10647 (N_10647,N_8392,N_9775);
or U10648 (N_10648,N_9249,N_8890);
or U10649 (N_10649,N_9594,N_8979);
nand U10650 (N_10650,N_7569,N_9424);
nor U10651 (N_10651,N_8379,N_9335);
nand U10652 (N_10652,N_8215,N_9323);
and U10653 (N_10653,N_8633,N_8232);
xor U10654 (N_10654,N_8442,N_9344);
xor U10655 (N_10655,N_9853,N_9184);
nand U10656 (N_10656,N_9106,N_9789);
xor U10657 (N_10657,N_9431,N_9979);
nor U10658 (N_10658,N_8409,N_8810);
and U10659 (N_10659,N_9915,N_8314);
nor U10660 (N_10660,N_9715,N_8093);
nor U10661 (N_10661,N_7903,N_7989);
or U10662 (N_10662,N_7667,N_9470);
nand U10663 (N_10663,N_7591,N_9963);
xnor U10664 (N_10664,N_9630,N_9345);
and U10665 (N_10665,N_9356,N_9555);
nor U10666 (N_10666,N_9143,N_9154);
xnor U10667 (N_10667,N_8068,N_8390);
nand U10668 (N_10668,N_7635,N_8711);
or U10669 (N_10669,N_9838,N_7581);
or U10670 (N_10670,N_8977,N_9354);
nand U10671 (N_10671,N_7740,N_9952);
nor U10672 (N_10672,N_8925,N_8079);
nor U10673 (N_10673,N_8787,N_9280);
or U10674 (N_10674,N_8653,N_9780);
nor U10675 (N_10675,N_9720,N_9908);
or U10676 (N_10676,N_8201,N_7938);
and U10677 (N_10677,N_9025,N_9858);
nand U10678 (N_10678,N_7632,N_8968);
xor U10679 (N_10679,N_8144,N_7680);
nor U10680 (N_10680,N_9842,N_9835);
xnor U10681 (N_10681,N_7954,N_7783);
nor U10682 (N_10682,N_7832,N_9329);
nor U10683 (N_10683,N_7671,N_8812);
xor U10684 (N_10684,N_9590,N_8929);
and U10685 (N_10685,N_9215,N_8295);
or U10686 (N_10686,N_9068,N_8652);
xor U10687 (N_10687,N_7822,N_9970);
or U10688 (N_10688,N_9740,N_7584);
and U10689 (N_10689,N_8976,N_8477);
or U10690 (N_10690,N_7710,N_9210);
or U10691 (N_10691,N_7542,N_9520);
xnor U10692 (N_10692,N_7793,N_9212);
and U10693 (N_10693,N_7866,N_7728);
or U10694 (N_10694,N_7943,N_9655);
xor U10695 (N_10695,N_7795,N_8940);
nor U10696 (N_10696,N_7563,N_9894);
xnor U10697 (N_10697,N_8051,N_8149);
xnor U10698 (N_10698,N_8375,N_8488);
or U10699 (N_10699,N_9057,N_8966);
xnor U10700 (N_10700,N_9898,N_8255);
or U10701 (N_10701,N_8189,N_9886);
nand U10702 (N_10702,N_8789,N_8408);
or U10703 (N_10703,N_9845,N_9939);
nor U10704 (N_10704,N_9137,N_8422);
xor U10705 (N_10705,N_9884,N_7559);
nor U10706 (N_10706,N_9270,N_7562);
nand U10707 (N_10707,N_9739,N_7940);
and U10708 (N_10708,N_7800,N_7955);
xor U10709 (N_10709,N_7625,N_7987);
and U10710 (N_10710,N_7974,N_9452);
nor U10711 (N_10711,N_7523,N_9753);
xor U10712 (N_10712,N_9472,N_8660);
nor U10713 (N_10713,N_8447,N_9163);
and U10714 (N_10714,N_8627,N_9338);
and U10715 (N_10715,N_8995,N_8745);
and U10716 (N_10716,N_9909,N_8899);
nor U10717 (N_10717,N_8115,N_9542);
nor U10718 (N_10718,N_8723,N_8641);
nand U10719 (N_10719,N_7878,N_8958);
nand U10720 (N_10720,N_9404,N_9457);
and U10721 (N_10721,N_9959,N_8424);
xor U10722 (N_10722,N_9402,N_9024);
or U10723 (N_10723,N_8778,N_9115);
xnor U10724 (N_10724,N_8168,N_7619);
nand U10725 (N_10725,N_9515,N_8386);
nor U10726 (N_10726,N_9772,N_8575);
nor U10727 (N_10727,N_8416,N_9002);
nor U10728 (N_10728,N_7617,N_9987);
or U10729 (N_10729,N_7582,N_7936);
and U10730 (N_10730,N_8556,N_7630);
or U10731 (N_10731,N_8980,N_9419);
or U10732 (N_10732,N_9370,N_7759);
nor U10733 (N_10733,N_8521,N_9957);
nor U10734 (N_10734,N_8712,N_8465);
or U10735 (N_10735,N_9221,N_8936);
nand U10736 (N_10736,N_8839,N_9489);
nor U10737 (N_10737,N_9193,N_8473);
or U10738 (N_10738,N_8985,N_7669);
nand U10739 (N_10739,N_8483,N_9794);
nand U10740 (N_10740,N_8188,N_7833);
xor U10741 (N_10741,N_8942,N_8355);
nand U10742 (N_10742,N_8591,N_8984);
nor U10743 (N_10743,N_8368,N_8462);
and U10744 (N_10744,N_8614,N_8669);
nand U10745 (N_10745,N_8397,N_7586);
and U10746 (N_10746,N_7641,N_8415);
xnor U10747 (N_10747,N_7786,N_7571);
nand U10748 (N_10748,N_9506,N_9880);
and U10749 (N_10749,N_7520,N_7754);
and U10750 (N_10750,N_7957,N_9811);
or U10751 (N_10751,N_8266,N_8746);
nor U10752 (N_10752,N_9950,N_9343);
or U10753 (N_10753,N_8860,N_9976);
nor U10754 (N_10754,N_8028,N_7881);
and U10755 (N_10755,N_7897,N_9872);
and U10756 (N_10756,N_9816,N_9634);
or U10757 (N_10757,N_9738,N_8801);
xor U10758 (N_10758,N_9092,N_7558);
nand U10759 (N_10759,N_8114,N_9290);
or U10760 (N_10760,N_9488,N_7834);
xnor U10761 (N_10761,N_7761,N_8137);
nand U10762 (N_10762,N_8343,N_9205);
nor U10763 (N_10763,N_9336,N_8493);
nand U10764 (N_10764,N_9998,N_9416);
nand U10765 (N_10765,N_8024,N_7831);
nand U10766 (N_10766,N_9039,N_8087);
or U10767 (N_10767,N_9793,N_9973);
nor U10768 (N_10768,N_8246,N_7560);
xor U10769 (N_10769,N_9572,N_7548);
or U10770 (N_10770,N_7865,N_8638);
or U10771 (N_10771,N_9004,N_8198);
and U10772 (N_10772,N_9734,N_9610);
nor U10773 (N_10773,N_9608,N_8084);
or U10774 (N_10774,N_8507,N_9604);
nand U10775 (N_10775,N_9717,N_9272);
and U10776 (N_10776,N_9131,N_9312);
nand U10777 (N_10777,N_9474,N_8128);
and U10778 (N_10778,N_8369,N_9629);
and U10779 (N_10779,N_9951,N_8896);
nor U10780 (N_10780,N_8844,N_9821);
and U10781 (N_10781,N_8727,N_7755);
or U10782 (N_10782,N_8092,N_7556);
nor U10783 (N_10783,N_8225,N_9110);
and U10784 (N_10784,N_7874,N_7594);
and U10785 (N_10785,N_8292,N_9502);
nand U10786 (N_10786,N_9946,N_7703);
xor U10787 (N_10787,N_9511,N_9403);
xor U10788 (N_10788,N_9374,N_8147);
xnor U10789 (N_10789,N_9146,N_9043);
nand U10790 (N_10790,N_8039,N_8702);
nand U10791 (N_10791,N_8070,N_8605);
and U10792 (N_10792,N_7585,N_8139);
nand U10793 (N_10793,N_7686,N_7730);
xor U10794 (N_10794,N_9582,N_9541);
or U10795 (N_10795,N_8683,N_8109);
xnor U10796 (N_10796,N_8628,N_7575);
nand U10797 (N_10797,N_7810,N_8091);
xnor U10798 (N_10798,N_8259,N_8123);
xor U10799 (N_10799,N_8086,N_8342);
nand U10800 (N_10800,N_8667,N_9455);
xnor U10801 (N_10801,N_9534,N_7670);
nand U10802 (N_10802,N_9136,N_7999);
xor U10803 (N_10803,N_8221,N_9905);
xor U10804 (N_10804,N_8729,N_9171);
nand U10805 (N_10805,N_9389,N_7898);
and U10806 (N_10806,N_7814,N_8360);
nor U10807 (N_10807,N_8531,N_8288);
nand U10808 (N_10808,N_9540,N_9975);
xor U10809 (N_10809,N_9417,N_9911);
and U10810 (N_10810,N_7820,N_8760);
nand U10811 (N_10811,N_8964,N_8815);
or U10812 (N_10812,N_8313,N_9735);
and U10813 (N_10813,N_9921,N_9491);
nor U10814 (N_10814,N_7512,N_8799);
nand U10815 (N_10815,N_8316,N_8750);
xnor U10816 (N_10816,N_7775,N_8671);
and U10817 (N_10817,N_9490,N_9011);
and U10818 (N_10818,N_8499,N_8027);
xnor U10819 (N_10819,N_8023,N_9033);
and U10820 (N_10820,N_9054,N_9732);
and U10821 (N_10821,N_9042,N_8401);
nor U10822 (N_10822,N_9045,N_9843);
xor U10823 (N_10823,N_7572,N_8431);
or U10824 (N_10824,N_8982,N_8010);
or U10825 (N_10825,N_7719,N_8190);
or U10826 (N_10826,N_8111,N_9889);
xnor U10827 (N_10827,N_8828,N_7608);
or U10828 (N_10828,N_9492,N_7696);
and U10829 (N_10829,N_8668,N_8535);
xnor U10830 (N_10830,N_9788,N_9799);
and U10831 (N_10831,N_7902,N_9456);
and U10832 (N_10832,N_9619,N_8986);
nor U10833 (N_10833,N_7960,N_8166);
nand U10834 (N_10834,N_9591,N_7665);
xor U10835 (N_10835,N_9362,N_9185);
nand U10836 (N_10836,N_9978,N_9412);
or U10837 (N_10837,N_7948,N_8677);
and U10838 (N_10838,N_9391,N_8420);
nand U10839 (N_10839,N_8754,N_7945);
or U10840 (N_10840,N_9401,N_7524);
xnor U10841 (N_10841,N_8357,N_9426);
xnor U10842 (N_10842,N_8833,N_7975);
xor U10843 (N_10843,N_8848,N_9046);
nand U10844 (N_10844,N_9722,N_8656);
and U10845 (N_10845,N_9649,N_8085);
xor U10846 (N_10846,N_8938,N_8635);
or U10847 (N_10847,N_9770,N_9498);
or U10848 (N_10848,N_9593,N_8474);
or U10849 (N_10849,N_7752,N_9322);
and U10850 (N_10850,N_7901,N_9595);
or U10851 (N_10851,N_9631,N_8625);
nand U10852 (N_10852,N_7607,N_8822);
nand U10853 (N_10853,N_9699,N_9275);
xor U10854 (N_10854,N_9606,N_9549);
nor U10855 (N_10855,N_9327,N_8513);
nand U10856 (N_10856,N_9583,N_9388);
nor U10857 (N_10857,N_8912,N_7624);
or U10858 (N_10858,N_9941,N_9638);
and U10859 (N_10859,N_9751,N_9698);
xor U10860 (N_10860,N_8560,N_9500);
and U10861 (N_10861,N_9875,N_9791);
and U10862 (N_10862,N_9928,N_7662);
and U10863 (N_10863,N_8461,N_7932);
nand U10864 (N_10864,N_8320,N_9438);
nand U10865 (N_10865,N_8140,N_8218);
and U10866 (N_10866,N_9501,N_8714);
nor U10867 (N_10867,N_7570,N_8018);
nor U10868 (N_10868,N_8016,N_7688);
nand U10869 (N_10869,N_7850,N_8827);
or U10870 (N_10870,N_9685,N_8993);
or U10871 (N_10871,N_8871,N_9217);
nor U10872 (N_10872,N_9562,N_9861);
and U10873 (N_10873,N_9179,N_8463);
nand U10874 (N_10874,N_9910,N_8098);
xnor U10875 (N_10875,N_9281,N_7949);
or U10876 (N_10876,N_8453,N_7981);
or U10877 (N_10877,N_9687,N_8359);
xnor U10878 (N_10878,N_8057,N_8886);
xnor U10879 (N_10879,N_8530,N_9682);
and U10880 (N_10880,N_8421,N_7598);
xnor U10881 (N_10881,N_8335,N_7557);
and U10882 (N_10882,N_8119,N_9067);
or U10883 (N_10883,N_8035,N_8990);
nor U10884 (N_10884,N_8136,N_8550);
xor U10885 (N_10885,N_9856,N_8726);
nor U10886 (N_10886,N_9748,N_7574);
or U10887 (N_10887,N_9339,N_9955);
xor U10888 (N_10888,N_9030,N_9443);
nand U10889 (N_10889,N_9870,N_8191);
and U10890 (N_10890,N_8796,N_8766);
xnor U10891 (N_10891,N_7965,N_9645);
xnor U10892 (N_10892,N_8983,N_8759);
or U10893 (N_10893,N_8319,N_9010);
xor U10894 (N_10894,N_8489,N_9635);
and U10895 (N_10895,N_8518,N_9264);
and U10896 (N_10896,N_7533,N_8600);
or U10897 (N_10897,N_8481,N_8272);
xnor U10898 (N_10898,N_8100,N_7799);
xor U10899 (N_10899,N_7713,N_9901);
nor U10900 (N_10900,N_9394,N_8162);
nand U10901 (N_10901,N_8687,N_8317);
xnor U10902 (N_10902,N_8173,N_9436);
nand U10903 (N_10903,N_8743,N_7702);
nor U10904 (N_10904,N_9616,N_8167);
and U10905 (N_10905,N_7873,N_7837);
and U10906 (N_10906,N_8417,N_8002);
and U10907 (N_10907,N_8285,N_7772);
or U10908 (N_10908,N_9326,N_7622);
nand U10909 (N_10909,N_8458,N_8460);
nor U10910 (N_10910,N_8997,N_8126);
nand U10911 (N_10911,N_9897,N_7764);
and U10912 (N_10912,N_8960,N_9949);
nor U10913 (N_10913,N_9924,N_9440);
nor U10914 (N_10914,N_9305,N_7543);
xnor U10915 (N_10915,N_9650,N_8696);
nand U10916 (N_10916,N_9194,N_7589);
nor U10917 (N_10917,N_9519,N_9170);
nor U10918 (N_10918,N_8052,N_9651);
nor U10919 (N_10919,N_9371,N_9022);
nor U10920 (N_10920,N_9230,N_7839);
nor U10921 (N_10921,N_9766,N_9347);
or U10922 (N_10922,N_7699,N_8350);
xor U10923 (N_10923,N_8269,N_8558);
nand U10924 (N_10924,N_8047,N_8765);
and U10925 (N_10925,N_9851,N_9460);
and U10926 (N_10926,N_9826,N_7714);
nor U10927 (N_10927,N_7648,N_9810);
nand U10928 (N_10928,N_9513,N_8498);
xnor U10929 (N_10929,N_9427,N_9525);
nor U10930 (N_10930,N_7769,N_8103);
or U10931 (N_10931,N_7979,N_8577);
and U10932 (N_10932,N_8555,N_8780);
and U10933 (N_10933,N_9579,N_7962);
and U10934 (N_10934,N_7642,N_9938);
and U10935 (N_10935,N_9694,N_7664);
or U10936 (N_10936,N_9256,N_9487);
xnor U10937 (N_10937,N_9945,N_9382);
xor U10938 (N_10938,N_9517,N_8464);
nor U10939 (N_10939,N_8581,N_8554);
or U10940 (N_10940,N_8800,N_8007);
or U10941 (N_10941,N_8077,N_8096);
nand U10942 (N_10942,N_8240,N_7971);
xor U10943 (N_10943,N_9133,N_9824);
xor U10944 (N_10944,N_8387,N_8403);
xnor U10945 (N_10945,N_8472,N_9222);
nor U10946 (N_10946,N_8572,N_9399);
xnor U10947 (N_10947,N_9308,N_8475);
nor U10948 (N_10948,N_9055,N_8987);
nand U10949 (N_10949,N_9675,N_8161);
nand U10950 (N_10950,N_9586,N_8956);
or U10951 (N_10951,N_8744,N_9102);
nand U10952 (N_10952,N_7551,N_9865);
nor U10953 (N_10953,N_8310,N_7765);
and U10954 (N_10954,N_9974,N_8438);
and U10955 (N_10955,N_9235,N_8970);
xnor U10956 (N_10956,N_8311,N_9601);
or U10957 (N_10957,N_7773,N_8566);
nor U10958 (N_10958,N_9790,N_9258);
and U10959 (N_10959,N_9093,N_9294);
nand U10960 (N_10960,N_9448,N_8256);
nand U10961 (N_10961,N_7864,N_8776);
xnor U10962 (N_10962,N_7537,N_9689);
or U10963 (N_10963,N_8325,N_9216);
nand U10964 (N_10964,N_7618,N_7627);
or U10965 (N_10965,N_8352,N_8151);
or U10966 (N_10966,N_9353,N_8604);
nand U10967 (N_10967,N_9747,N_9178);
nand U10968 (N_10968,N_9381,N_9471);
nor U10969 (N_10969,N_7984,N_9557);
nor U10970 (N_10970,N_9084,N_8772);
nand U10971 (N_10971,N_9276,N_8689);
nand U10972 (N_10972,N_8601,N_8135);
nand U10973 (N_10973,N_8305,N_8694);
nand U10974 (N_10974,N_8399,N_9674);
xor U10975 (N_10975,N_7748,N_9822);
nand U10976 (N_10976,N_9113,N_9361);
xor U10977 (N_10977,N_7661,N_9887);
and U10978 (N_10978,N_9321,N_8226);
and U10979 (N_10979,N_7927,N_7507);
nor U10980 (N_10980,N_9867,N_8043);
xnor U10981 (N_10981,N_8174,N_7915);
nand U10982 (N_10982,N_9688,N_8145);
or U10983 (N_10983,N_9061,N_8436);
nand U10984 (N_10984,N_9378,N_8029);
and U10985 (N_10985,N_8911,N_9718);
nor U10986 (N_10986,N_8388,N_8340);
xnor U10987 (N_10987,N_8268,N_8972);
and U10988 (N_10988,N_9376,N_9172);
and U10989 (N_10989,N_7911,N_9932);
and U10990 (N_10990,N_8510,N_8492);
or U10991 (N_10991,N_9670,N_8777);
nor U10992 (N_10992,N_8818,N_8611);
nand U10993 (N_10993,N_8542,N_7970);
and U10994 (N_10994,N_9644,N_8291);
nor U10995 (N_10995,N_8389,N_8297);
nor U10996 (N_10996,N_8798,N_8699);
nor U10997 (N_10997,N_9444,N_7725);
nor U10998 (N_10998,N_8423,N_8830);
nor U10999 (N_10999,N_8165,N_9425);
nor U11000 (N_11000,N_9368,N_8504);
or U11001 (N_11001,N_8593,N_8888);
and U11002 (N_11002,N_8159,N_9364);
nand U11003 (N_11003,N_7871,N_8963);
nor U11004 (N_11004,N_9658,N_7550);
nor U11005 (N_11005,N_7883,N_9641);
nor U11006 (N_11006,N_8500,N_9288);
nor U11007 (N_11007,N_7655,N_9266);
nor U11008 (N_11008,N_8864,N_9052);
or U11009 (N_11009,N_8351,N_9395);
or U11010 (N_11010,N_8850,N_9509);
or U11011 (N_11011,N_7539,N_9758);
and U11012 (N_11012,N_8654,N_7846);
xnor U11013 (N_11013,N_8545,N_7880);
or U11014 (N_11014,N_9070,N_9359);
or U11015 (N_11015,N_9701,N_8859);
and U11016 (N_11016,N_7899,N_8076);
nand U11017 (N_11017,N_8981,N_8901);
nor U11018 (N_11018,N_9726,N_9377);
or U11019 (N_11019,N_8680,N_7716);
or U11020 (N_11020,N_7698,N_9690);
nor U11021 (N_11021,N_7709,N_8691);
nand U11022 (N_11022,N_7564,N_8785);
xor U11023 (N_11023,N_7868,N_8347);
xnor U11024 (N_11024,N_8003,N_8851);
and U11025 (N_11025,N_9605,N_8058);
or U11026 (N_11026,N_9260,N_9213);
or U11027 (N_11027,N_8540,N_9285);
and U11028 (N_11028,N_7926,N_9464);
or U11029 (N_11029,N_8867,N_8792);
and U11030 (N_11030,N_9852,N_9926);
or U11031 (N_11031,N_8323,N_8212);
or U11032 (N_11032,N_9072,N_9771);
xnor U11033 (N_11033,N_9607,N_8238);
or U11034 (N_11034,N_9652,N_7711);
nand U11035 (N_11035,N_8220,N_8559);
and U11036 (N_11036,N_8941,N_8949);
and U11037 (N_11037,N_7886,N_9018);
xor U11038 (N_11038,N_9199,N_9056);
and U11039 (N_11039,N_8693,N_8121);
nand U11040 (N_11040,N_8435,N_8252);
nand U11041 (N_11041,N_9435,N_8937);
and U11042 (N_11042,N_8237,N_9566);
xnor U11043 (N_11043,N_8250,N_7521);
and U11044 (N_11044,N_8790,N_9599);
and U11045 (N_11045,N_8950,N_9246);
or U11046 (N_11046,N_7856,N_9267);
nor U11047 (N_11047,N_8312,N_8254);
nand U11048 (N_11048,N_9380,N_8755);
nand U11049 (N_11049,N_7912,N_9355);
xor U11050 (N_11050,N_8527,N_8837);
or U11051 (N_11051,N_8176,N_8612);
nor U11052 (N_11052,N_8809,N_7952);
nand U11053 (N_11053,N_9536,N_9916);
or U11054 (N_11054,N_9903,N_8767);
or U11055 (N_11055,N_8073,N_7828);
and U11056 (N_11056,N_7693,N_8006);
or U11057 (N_11057,N_8861,N_9823);
and U11058 (N_11058,N_7905,N_7742);
and U11059 (N_11059,N_7595,N_7700);
nor U11060 (N_11060,N_7985,N_7907);
nand U11061 (N_11061,N_7813,N_8602);
nand U11062 (N_11062,N_9613,N_9914);
nand U11063 (N_11063,N_9341,N_9596);
nor U11064 (N_11064,N_7941,N_9584);
nor U11065 (N_11065,N_8437,N_9988);
xnor U11066 (N_11066,N_9896,N_9532);
xnor U11067 (N_11067,N_8229,N_9795);
xor U11068 (N_11068,N_7916,N_8553);
nand U11069 (N_11069,N_7953,N_8588);
and U11070 (N_11070,N_9441,N_9243);
nand U11071 (N_11071,N_8853,N_8757);
xor U11072 (N_11072,N_7845,N_8398);
nor U11073 (N_11073,N_9497,N_8845);
xor U11074 (N_11074,N_8449,N_9155);
nor U11075 (N_11075,N_8430,N_9446);
or U11076 (N_11076,N_8589,N_8648);
nor U11077 (N_11077,N_8088,N_8348);
and U11078 (N_11078,N_9484,N_8083);
xor U11079 (N_11079,N_9892,N_8916);
nor U11080 (N_11080,N_8370,N_7818);
xor U11081 (N_11081,N_9531,N_7727);
nand U11082 (N_11082,N_7541,N_9182);
and U11083 (N_11083,N_8541,N_9465);
nand U11084 (N_11084,N_9711,N_9712);
nand U11085 (N_11085,N_8721,N_8008);
and U11086 (N_11086,N_8549,N_9899);
and U11087 (N_11087,N_8622,N_8582);
xor U11088 (N_11088,N_8869,N_8095);
xor U11089 (N_11089,N_7842,N_8318);
or U11090 (N_11090,N_7904,N_8640);
nor U11091 (N_11091,N_7790,N_8262);
or U11092 (N_11092,N_9226,N_8330);
and U11093 (N_11093,N_9313,N_9254);
or U11094 (N_11094,N_9554,N_8153);
or U11095 (N_11095,N_8239,N_7973);
nand U11096 (N_11096,N_9150,N_8102);
and U11097 (N_11097,N_9350,N_7506);
xor U11098 (N_11098,N_8594,N_7760);
and U11099 (N_11099,N_7884,N_8905);
nor U11100 (N_11100,N_9180,N_9236);
nor U11101 (N_11101,N_7502,N_8071);
or U11102 (N_11102,N_9859,N_8406);
nor U11103 (N_11103,N_9142,N_8634);
nor U11104 (N_11104,N_7841,N_8367);
xor U11105 (N_11105,N_9078,N_8645);
nor U11106 (N_11106,N_9469,N_9125);
nand U11107 (N_11107,N_9383,N_8877);
or U11108 (N_11108,N_7825,N_8391);
nor U11109 (N_11109,N_8248,N_8411);
and U11110 (N_11110,N_9779,N_8356);
and U11111 (N_11111,N_9936,N_9095);
nand U11112 (N_11112,N_9414,N_8952);
xnor U11113 (N_11113,N_8998,N_9991);
nand U11114 (N_11114,N_8681,N_7891);
or U11115 (N_11115,N_9615,N_8989);
and U11116 (N_11116,N_9073,N_7797);
xnor U11117 (N_11117,N_8030,N_8657);
xor U11118 (N_11118,N_7887,N_9696);
and U11119 (N_11119,N_9633,N_9406);
or U11120 (N_11120,N_8570,N_9293);
or U11121 (N_11121,N_8569,N_7743);
nand U11122 (N_11122,N_9297,N_9218);
and U11123 (N_11123,N_7791,N_7821);
nand U11124 (N_11124,N_9848,N_9508);
nand U11125 (N_11125,N_8804,N_8020);
xor U11126 (N_11126,N_7889,N_7528);
nand U11127 (N_11127,N_9648,N_8948);
nand U11128 (N_11128,N_8338,N_8158);
and U11129 (N_11129,N_9580,N_8264);
xor U11130 (N_11130,N_9923,N_9581);
nand U11131 (N_11131,N_9882,N_9080);
nand U11132 (N_11132,N_8817,N_7611);
nand U11133 (N_11133,N_8276,N_8965);
nand U11134 (N_11134,N_9850,N_9340);
nand U11135 (N_11135,N_8414,N_9096);
or U11136 (N_11136,N_8182,N_8630);
nand U11137 (N_11137,N_9069,N_7827);
and U11138 (N_11138,N_9609,N_9122);
xnor U11139 (N_11139,N_7972,N_8244);
nor U11140 (N_11140,N_9202,N_8821);
nor U11141 (N_11141,N_8503,N_8470);
and U11142 (N_11142,N_8069,N_9760);
or U11143 (N_11143,N_9992,N_7633);
and U11144 (N_11144,N_8082,N_8187);
and U11145 (N_11145,N_8944,N_9463);
and U11146 (N_11146,N_7896,N_8362);
nand U11147 (N_11147,N_8050,N_8097);
nor U11148 (N_11148,N_8242,N_8049);
or U11149 (N_11149,N_8433,N_7980);
xor U11150 (N_11150,N_9348,N_9663);
nand U11151 (N_11151,N_9956,N_8080);
xor U11152 (N_11152,N_9437,N_7778);
xnor U11153 (N_11153,N_9767,N_9229);
xnor U11154 (N_11154,N_9161,N_9847);
and U11155 (N_11155,N_9961,N_8217);
nor U11156 (N_11156,N_9320,N_9673);
xnor U11157 (N_11157,N_8797,N_9311);
xor U11158 (N_11158,N_8491,N_9268);
and U11159 (N_11159,N_9369,N_8738);
xnor U11160 (N_11160,N_9837,N_8124);
and U11161 (N_11161,N_7650,N_9719);
or U11162 (N_11162,N_9231,N_8670);
xnor U11163 (N_11163,N_9242,N_9700);
xor U11164 (N_11164,N_9458,N_8495);
xor U11165 (N_11165,N_8679,N_8954);
nand U11166 (N_11166,N_8606,N_7636);
or U11167 (N_11167,N_8017,N_9877);
or U11168 (N_11168,N_8446,N_9048);
xor U11169 (N_11169,N_7673,N_8813);
nand U11170 (N_11170,N_8592,N_9081);
nand U11171 (N_11171,N_8454,N_9893);
nor U11172 (N_11172,N_8427,N_8208);
xor U11173 (N_11173,N_7929,N_9467);
xnor U11174 (N_11174,N_8735,N_9836);
or U11175 (N_11175,N_8659,N_7895);
nand U11176 (N_11176,N_9860,N_8034);
nor U11177 (N_11177,N_9804,N_8959);
nand U11178 (N_11178,N_8880,N_8306);
nand U11179 (N_11179,N_8762,N_8004);
and U11180 (N_11180,N_7777,N_9942);
nand U11181 (N_11181,N_7504,N_8496);
xor U11182 (N_11182,N_8482,N_9640);
or U11183 (N_11183,N_8207,N_8874);
nor U11184 (N_11184,N_8067,N_8585);
xnor U11185 (N_11185,N_9759,N_8321);
nand U11186 (N_11186,N_9724,N_8728);
xnor U11187 (N_11187,N_8251,N_9247);
or U11188 (N_11188,N_9761,N_7515);
nor U11189 (N_11189,N_9496,N_8921);
nand U11190 (N_11190,N_9032,N_8788);
nor U11191 (N_11191,N_9304,N_8090);
nand U11192 (N_11192,N_8175,N_9085);
xor U11193 (N_11193,N_7998,N_9937);
or U11194 (N_11194,N_8074,N_8200);
nand U11195 (N_11195,N_8836,N_9197);
xor U11196 (N_11196,N_7615,N_9097);
and U11197 (N_11197,N_8732,N_8534);
nand U11198 (N_11198,N_8922,N_8105);
and U11199 (N_11199,N_7723,N_8918);
xnor U11200 (N_11200,N_8486,N_8893);
or U11201 (N_11201,N_9044,N_9646);
nor U11202 (N_11202,N_7977,N_7993);
nor U11203 (N_11203,N_9442,N_9147);
or U11204 (N_11204,N_9680,N_7811);
and U11205 (N_11205,N_9375,N_9174);
nor U11206 (N_11206,N_8736,N_9598);
and U11207 (N_11207,N_9234,N_8178);
nand U11208 (N_11208,N_9661,N_8382);
nor U11209 (N_11209,N_9636,N_8947);
nor U11210 (N_11210,N_9529,N_8441);
nand U11211 (N_11211,N_9510,N_8543);
nand U11212 (N_11212,N_9074,N_9149);
nor U11213 (N_11213,N_9316,N_9559);
nor U11214 (N_11214,N_8875,N_8089);
and U11215 (N_11215,N_9981,N_9721);
and U11216 (N_11216,N_9925,N_9545);
xnor U11217 (N_11217,N_9977,N_9379);
and U11218 (N_11218,N_9830,N_9878);
xor U11219 (N_11219,N_9891,N_7934);
xor U11220 (N_11220,N_8519,N_7862);
or U11221 (N_11221,N_8643,N_9076);
or U11222 (N_11222,N_8282,N_8118);
or U11223 (N_11223,N_9786,N_7966);
nor U11224 (N_11224,N_9494,N_9900);
nand U11225 (N_11225,N_9552,N_8615);
nand U11226 (N_11226,N_8327,N_8054);
and U11227 (N_11227,N_8412,N_8889);
or U11228 (N_11228,N_8066,N_9573);
nand U11229 (N_11229,N_7958,N_8532);
nor U11230 (N_11230,N_8608,N_9503);
or U11231 (N_11231,N_8106,N_8025);
nor U11232 (N_11232,N_7530,N_8448);
nor U11233 (N_11233,N_8031,N_8651);
and U11234 (N_11234,N_9162,N_9118);
nand U11235 (N_11235,N_8573,N_8931);
or U11236 (N_11236,N_7738,N_9697);
and U11237 (N_11237,N_9499,N_8286);
nor U11238 (N_11238,N_8045,N_8619);
or U11239 (N_11239,N_7532,N_9014);
nor U11240 (N_11240,N_9693,N_8840);
xnor U11241 (N_11241,N_8646,N_9289);
and U11242 (N_11242,N_8704,N_9493);
xor U11243 (N_11243,N_8703,N_9274);
or U11244 (N_11244,N_8786,N_8222);
or U11245 (N_11245,N_8955,N_7684);
xnor U11246 (N_11246,N_7779,N_9731);
or U11247 (N_11247,N_8803,N_7616);
nor U11248 (N_11248,N_8469,N_8371);
xor U11249 (N_11249,N_9408,N_9291);
and U11250 (N_11250,N_8132,N_9909);
or U11251 (N_11251,N_7658,N_8742);
nor U11252 (N_11252,N_8735,N_9025);
nand U11253 (N_11253,N_9523,N_9176);
or U11254 (N_11254,N_9570,N_8734);
nand U11255 (N_11255,N_9118,N_9751);
and U11256 (N_11256,N_8415,N_9439);
or U11257 (N_11257,N_8198,N_8229);
xor U11258 (N_11258,N_8422,N_7595);
and U11259 (N_11259,N_7734,N_8733);
nor U11260 (N_11260,N_8955,N_9030);
or U11261 (N_11261,N_9466,N_9189);
nand U11262 (N_11262,N_7534,N_8115);
or U11263 (N_11263,N_8200,N_9815);
xor U11264 (N_11264,N_8617,N_8694);
and U11265 (N_11265,N_7918,N_8031);
xor U11266 (N_11266,N_8714,N_7683);
nand U11267 (N_11267,N_9003,N_9833);
and U11268 (N_11268,N_9649,N_8210);
and U11269 (N_11269,N_7782,N_9845);
nand U11270 (N_11270,N_8978,N_9881);
and U11271 (N_11271,N_9328,N_9407);
and U11272 (N_11272,N_7962,N_8347);
nor U11273 (N_11273,N_9740,N_8452);
xor U11274 (N_11274,N_7999,N_7582);
or U11275 (N_11275,N_8901,N_9779);
and U11276 (N_11276,N_8795,N_9145);
or U11277 (N_11277,N_9824,N_8246);
or U11278 (N_11278,N_8784,N_8941);
nand U11279 (N_11279,N_8269,N_8078);
or U11280 (N_11280,N_8057,N_9321);
xnor U11281 (N_11281,N_9239,N_7667);
and U11282 (N_11282,N_7886,N_8369);
xnor U11283 (N_11283,N_9744,N_7516);
xor U11284 (N_11284,N_9329,N_8398);
or U11285 (N_11285,N_8147,N_9189);
nor U11286 (N_11286,N_9234,N_8104);
nor U11287 (N_11287,N_8708,N_7820);
xor U11288 (N_11288,N_9087,N_8515);
nor U11289 (N_11289,N_8893,N_8673);
nor U11290 (N_11290,N_9395,N_8628);
and U11291 (N_11291,N_8419,N_9641);
nor U11292 (N_11292,N_9226,N_8742);
and U11293 (N_11293,N_9210,N_8906);
nand U11294 (N_11294,N_8056,N_9696);
or U11295 (N_11295,N_7860,N_7656);
xor U11296 (N_11296,N_9532,N_7884);
nor U11297 (N_11297,N_8287,N_7953);
xor U11298 (N_11298,N_8644,N_9682);
nor U11299 (N_11299,N_8973,N_9608);
or U11300 (N_11300,N_9897,N_8940);
or U11301 (N_11301,N_9702,N_8826);
xor U11302 (N_11302,N_8882,N_7896);
or U11303 (N_11303,N_8441,N_9895);
nand U11304 (N_11304,N_9182,N_9691);
or U11305 (N_11305,N_7904,N_8764);
nand U11306 (N_11306,N_7605,N_8304);
nand U11307 (N_11307,N_9816,N_8778);
nor U11308 (N_11308,N_8330,N_7698);
and U11309 (N_11309,N_9464,N_7807);
and U11310 (N_11310,N_7964,N_8916);
nand U11311 (N_11311,N_9012,N_9050);
and U11312 (N_11312,N_8459,N_9145);
or U11313 (N_11313,N_9044,N_8125);
xor U11314 (N_11314,N_9365,N_8677);
nand U11315 (N_11315,N_7649,N_9492);
xor U11316 (N_11316,N_9873,N_7621);
or U11317 (N_11317,N_9501,N_9401);
xor U11318 (N_11318,N_8364,N_8078);
xor U11319 (N_11319,N_8651,N_8440);
or U11320 (N_11320,N_7597,N_7891);
nor U11321 (N_11321,N_9080,N_8739);
xnor U11322 (N_11322,N_9941,N_8906);
nand U11323 (N_11323,N_8214,N_8411);
and U11324 (N_11324,N_8119,N_8140);
nor U11325 (N_11325,N_8325,N_8862);
nand U11326 (N_11326,N_8655,N_8664);
nor U11327 (N_11327,N_7569,N_9964);
or U11328 (N_11328,N_8078,N_9087);
xnor U11329 (N_11329,N_8450,N_7737);
xor U11330 (N_11330,N_7817,N_9309);
and U11331 (N_11331,N_8276,N_7691);
or U11332 (N_11332,N_7923,N_9429);
nor U11333 (N_11333,N_9096,N_8662);
xor U11334 (N_11334,N_7656,N_9104);
nand U11335 (N_11335,N_8040,N_8612);
xor U11336 (N_11336,N_8859,N_9460);
or U11337 (N_11337,N_9193,N_8695);
nand U11338 (N_11338,N_7755,N_8784);
and U11339 (N_11339,N_9325,N_8605);
xnor U11340 (N_11340,N_8596,N_9301);
xor U11341 (N_11341,N_7651,N_7883);
xnor U11342 (N_11342,N_9881,N_7774);
xnor U11343 (N_11343,N_7691,N_7672);
and U11344 (N_11344,N_9151,N_8495);
and U11345 (N_11345,N_9870,N_8622);
and U11346 (N_11346,N_7997,N_8101);
xnor U11347 (N_11347,N_9696,N_7556);
xnor U11348 (N_11348,N_9066,N_8571);
or U11349 (N_11349,N_8312,N_9881);
nand U11350 (N_11350,N_7726,N_8255);
nor U11351 (N_11351,N_9098,N_9472);
and U11352 (N_11352,N_9465,N_9933);
nand U11353 (N_11353,N_9632,N_9083);
nand U11354 (N_11354,N_7831,N_9432);
xnor U11355 (N_11355,N_9488,N_9950);
nand U11356 (N_11356,N_8818,N_8062);
xor U11357 (N_11357,N_8339,N_9707);
xnor U11358 (N_11358,N_8467,N_7844);
xnor U11359 (N_11359,N_9099,N_9832);
xnor U11360 (N_11360,N_9347,N_9619);
nor U11361 (N_11361,N_9117,N_8615);
or U11362 (N_11362,N_9329,N_8672);
nor U11363 (N_11363,N_8256,N_9862);
and U11364 (N_11364,N_8159,N_8043);
or U11365 (N_11365,N_8518,N_7622);
and U11366 (N_11366,N_8995,N_8837);
or U11367 (N_11367,N_8146,N_7514);
and U11368 (N_11368,N_8708,N_9150);
nor U11369 (N_11369,N_9677,N_9641);
nor U11370 (N_11370,N_9772,N_9904);
and U11371 (N_11371,N_8894,N_8439);
xnor U11372 (N_11372,N_8153,N_7575);
nand U11373 (N_11373,N_8188,N_9169);
and U11374 (N_11374,N_7725,N_9748);
nand U11375 (N_11375,N_7982,N_8911);
xor U11376 (N_11376,N_7814,N_7684);
and U11377 (N_11377,N_8976,N_8600);
nand U11378 (N_11378,N_8765,N_8055);
and U11379 (N_11379,N_7990,N_9646);
nor U11380 (N_11380,N_9485,N_7721);
xnor U11381 (N_11381,N_9816,N_8442);
or U11382 (N_11382,N_9845,N_8229);
xor U11383 (N_11383,N_9426,N_8574);
nor U11384 (N_11384,N_8978,N_8595);
xnor U11385 (N_11385,N_9300,N_8404);
and U11386 (N_11386,N_9846,N_8906);
xor U11387 (N_11387,N_9266,N_8169);
and U11388 (N_11388,N_9739,N_9068);
xor U11389 (N_11389,N_7851,N_9590);
nand U11390 (N_11390,N_8072,N_8580);
nor U11391 (N_11391,N_9031,N_7749);
nand U11392 (N_11392,N_8772,N_7832);
or U11393 (N_11393,N_9170,N_8908);
xor U11394 (N_11394,N_9644,N_7708);
and U11395 (N_11395,N_8065,N_9899);
xnor U11396 (N_11396,N_8889,N_8190);
xnor U11397 (N_11397,N_9570,N_7879);
nand U11398 (N_11398,N_8642,N_8604);
xnor U11399 (N_11399,N_9875,N_8520);
and U11400 (N_11400,N_9383,N_8051);
or U11401 (N_11401,N_8021,N_9159);
and U11402 (N_11402,N_7694,N_9220);
nand U11403 (N_11403,N_8434,N_8632);
or U11404 (N_11404,N_7671,N_9290);
xor U11405 (N_11405,N_8627,N_7799);
nor U11406 (N_11406,N_9695,N_9597);
and U11407 (N_11407,N_9014,N_9458);
nand U11408 (N_11408,N_9888,N_8951);
or U11409 (N_11409,N_9546,N_9555);
nand U11410 (N_11410,N_8719,N_9191);
nor U11411 (N_11411,N_9785,N_9203);
and U11412 (N_11412,N_8847,N_8194);
nor U11413 (N_11413,N_8089,N_9789);
nand U11414 (N_11414,N_8363,N_9814);
nor U11415 (N_11415,N_8352,N_9016);
or U11416 (N_11416,N_9898,N_9723);
nor U11417 (N_11417,N_8405,N_8484);
xor U11418 (N_11418,N_8768,N_9807);
xor U11419 (N_11419,N_9980,N_8117);
nor U11420 (N_11420,N_9648,N_7606);
nand U11421 (N_11421,N_8388,N_7548);
xnor U11422 (N_11422,N_8000,N_9968);
nand U11423 (N_11423,N_7800,N_9697);
or U11424 (N_11424,N_8656,N_8318);
or U11425 (N_11425,N_8512,N_8013);
xor U11426 (N_11426,N_9037,N_9774);
xor U11427 (N_11427,N_9049,N_8233);
nor U11428 (N_11428,N_8330,N_9199);
nand U11429 (N_11429,N_7941,N_7903);
nor U11430 (N_11430,N_7547,N_9028);
or U11431 (N_11431,N_8662,N_7721);
or U11432 (N_11432,N_8406,N_8537);
and U11433 (N_11433,N_8955,N_9804);
nand U11434 (N_11434,N_9748,N_8422);
or U11435 (N_11435,N_8803,N_8714);
nand U11436 (N_11436,N_9758,N_9317);
and U11437 (N_11437,N_7684,N_8577);
and U11438 (N_11438,N_8179,N_8082);
and U11439 (N_11439,N_7938,N_9474);
or U11440 (N_11440,N_9236,N_8214);
or U11441 (N_11441,N_8804,N_9824);
nor U11442 (N_11442,N_9227,N_9477);
or U11443 (N_11443,N_7514,N_8075);
or U11444 (N_11444,N_8784,N_9461);
nor U11445 (N_11445,N_7622,N_9115);
and U11446 (N_11446,N_8534,N_9116);
and U11447 (N_11447,N_9293,N_8210);
or U11448 (N_11448,N_7692,N_9241);
and U11449 (N_11449,N_9502,N_8032);
nand U11450 (N_11450,N_7533,N_7844);
nor U11451 (N_11451,N_8082,N_8822);
and U11452 (N_11452,N_7758,N_7784);
nor U11453 (N_11453,N_8823,N_7888);
xor U11454 (N_11454,N_8591,N_9191);
or U11455 (N_11455,N_8601,N_8930);
or U11456 (N_11456,N_8232,N_9235);
xor U11457 (N_11457,N_8300,N_9471);
and U11458 (N_11458,N_8221,N_9584);
nand U11459 (N_11459,N_8925,N_9613);
nand U11460 (N_11460,N_8843,N_8725);
nand U11461 (N_11461,N_8782,N_7659);
and U11462 (N_11462,N_8614,N_8859);
xor U11463 (N_11463,N_8669,N_9626);
xnor U11464 (N_11464,N_9061,N_8106);
or U11465 (N_11465,N_8190,N_9093);
xor U11466 (N_11466,N_7859,N_8375);
nand U11467 (N_11467,N_8965,N_7655);
and U11468 (N_11468,N_9295,N_8942);
nor U11469 (N_11469,N_9081,N_9936);
or U11470 (N_11470,N_8749,N_7845);
xor U11471 (N_11471,N_9117,N_7766);
or U11472 (N_11472,N_8593,N_8076);
xnor U11473 (N_11473,N_8269,N_9060);
nand U11474 (N_11474,N_7660,N_9463);
nand U11475 (N_11475,N_9235,N_9440);
nor U11476 (N_11476,N_8945,N_9715);
or U11477 (N_11477,N_7708,N_9859);
xor U11478 (N_11478,N_8488,N_8024);
and U11479 (N_11479,N_9056,N_8549);
nand U11480 (N_11480,N_9303,N_8190);
or U11481 (N_11481,N_8727,N_8524);
nor U11482 (N_11482,N_8239,N_9609);
and U11483 (N_11483,N_7921,N_7978);
nand U11484 (N_11484,N_8532,N_8540);
and U11485 (N_11485,N_8753,N_8329);
or U11486 (N_11486,N_9739,N_8466);
xor U11487 (N_11487,N_9805,N_9731);
nand U11488 (N_11488,N_9427,N_9911);
nor U11489 (N_11489,N_9036,N_8448);
nand U11490 (N_11490,N_8453,N_7581);
xor U11491 (N_11491,N_9692,N_8989);
nand U11492 (N_11492,N_9455,N_9504);
and U11493 (N_11493,N_8992,N_8538);
and U11494 (N_11494,N_8241,N_8631);
nor U11495 (N_11495,N_9116,N_9531);
and U11496 (N_11496,N_8426,N_8306);
nor U11497 (N_11497,N_8147,N_8545);
nand U11498 (N_11498,N_9662,N_8907);
and U11499 (N_11499,N_8542,N_7758);
nand U11500 (N_11500,N_9843,N_9097);
or U11501 (N_11501,N_9487,N_7668);
and U11502 (N_11502,N_8106,N_8547);
or U11503 (N_11503,N_9186,N_8647);
xnor U11504 (N_11504,N_7810,N_9094);
nand U11505 (N_11505,N_8812,N_9945);
nand U11506 (N_11506,N_8055,N_8538);
and U11507 (N_11507,N_9007,N_9109);
xnor U11508 (N_11508,N_8617,N_7804);
nand U11509 (N_11509,N_7745,N_8785);
nand U11510 (N_11510,N_7740,N_8867);
nand U11511 (N_11511,N_9615,N_9731);
xor U11512 (N_11512,N_7984,N_9323);
nand U11513 (N_11513,N_9273,N_9058);
and U11514 (N_11514,N_9488,N_9865);
nor U11515 (N_11515,N_8291,N_9107);
nor U11516 (N_11516,N_9279,N_9169);
nor U11517 (N_11517,N_8393,N_8722);
and U11518 (N_11518,N_9017,N_8070);
or U11519 (N_11519,N_8696,N_9366);
and U11520 (N_11520,N_8793,N_8448);
nand U11521 (N_11521,N_8988,N_7503);
nand U11522 (N_11522,N_9957,N_9992);
xnor U11523 (N_11523,N_9987,N_9525);
nor U11524 (N_11524,N_8255,N_7685);
or U11525 (N_11525,N_8458,N_7548);
xnor U11526 (N_11526,N_8920,N_8724);
nand U11527 (N_11527,N_8984,N_9027);
xor U11528 (N_11528,N_8633,N_8550);
or U11529 (N_11529,N_9809,N_8744);
nor U11530 (N_11530,N_8218,N_8064);
xor U11531 (N_11531,N_7888,N_8261);
xor U11532 (N_11532,N_7780,N_8200);
or U11533 (N_11533,N_9377,N_7554);
nor U11534 (N_11534,N_9841,N_9445);
nor U11535 (N_11535,N_7579,N_8451);
or U11536 (N_11536,N_9195,N_8821);
and U11537 (N_11537,N_7715,N_7799);
nor U11538 (N_11538,N_8656,N_9417);
nand U11539 (N_11539,N_9131,N_8494);
and U11540 (N_11540,N_8832,N_8218);
nand U11541 (N_11541,N_9324,N_9928);
or U11542 (N_11542,N_9369,N_7682);
nand U11543 (N_11543,N_9386,N_7939);
xor U11544 (N_11544,N_8138,N_8141);
nor U11545 (N_11545,N_9011,N_7923);
nor U11546 (N_11546,N_8421,N_9662);
xnor U11547 (N_11547,N_8855,N_7963);
and U11548 (N_11548,N_9484,N_7547);
nor U11549 (N_11549,N_9737,N_8712);
nand U11550 (N_11550,N_9278,N_9027);
nor U11551 (N_11551,N_9864,N_9132);
or U11552 (N_11552,N_9085,N_9811);
nand U11553 (N_11553,N_8557,N_7835);
and U11554 (N_11554,N_9337,N_8971);
or U11555 (N_11555,N_7921,N_8931);
xor U11556 (N_11556,N_8536,N_9879);
and U11557 (N_11557,N_9292,N_8871);
nor U11558 (N_11558,N_9386,N_8823);
nor U11559 (N_11559,N_9461,N_7609);
or U11560 (N_11560,N_7532,N_7542);
xor U11561 (N_11561,N_7903,N_7532);
nor U11562 (N_11562,N_9594,N_9567);
nor U11563 (N_11563,N_9249,N_9191);
or U11564 (N_11564,N_8288,N_7684);
xnor U11565 (N_11565,N_7978,N_9975);
and U11566 (N_11566,N_8231,N_9538);
nor U11567 (N_11567,N_7807,N_8284);
and U11568 (N_11568,N_9652,N_8734);
nand U11569 (N_11569,N_8675,N_8691);
nor U11570 (N_11570,N_8467,N_9382);
nor U11571 (N_11571,N_9272,N_9666);
nand U11572 (N_11572,N_9967,N_9968);
nor U11573 (N_11573,N_8672,N_9597);
nor U11574 (N_11574,N_8037,N_9435);
nand U11575 (N_11575,N_7833,N_9875);
xor U11576 (N_11576,N_9753,N_8592);
nand U11577 (N_11577,N_7783,N_9027);
or U11578 (N_11578,N_9574,N_8994);
nor U11579 (N_11579,N_9776,N_9901);
and U11580 (N_11580,N_7569,N_8441);
nor U11581 (N_11581,N_8784,N_8284);
and U11582 (N_11582,N_7516,N_7642);
nor U11583 (N_11583,N_9643,N_9713);
nor U11584 (N_11584,N_8821,N_8132);
nor U11585 (N_11585,N_7839,N_8905);
nor U11586 (N_11586,N_8794,N_7681);
and U11587 (N_11587,N_8426,N_8513);
or U11588 (N_11588,N_7733,N_8588);
and U11589 (N_11589,N_7660,N_9117);
and U11590 (N_11590,N_9198,N_8485);
xor U11591 (N_11591,N_8870,N_8889);
and U11592 (N_11592,N_9302,N_7895);
and U11593 (N_11593,N_8624,N_8421);
nand U11594 (N_11594,N_8942,N_9152);
nand U11595 (N_11595,N_9536,N_8450);
and U11596 (N_11596,N_9374,N_9269);
and U11597 (N_11597,N_8367,N_7783);
nor U11598 (N_11598,N_8157,N_8257);
nor U11599 (N_11599,N_9219,N_7756);
nor U11600 (N_11600,N_9395,N_7660);
nand U11601 (N_11601,N_8911,N_8553);
nor U11602 (N_11602,N_9522,N_8755);
nand U11603 (N_11603,N_9682,N_8522);
xnor U11604 (N_11604,N_9053,N_8785);
and U11605 (N_11605,N_9312,N_7850);
nand U11606 (N_11606,N_8910,N_7961);
xor U11607 (N_11607,N_8937,N_9146);
or U11608 (N_11608,N_8052,N_8919);
nand U11609 (N_11609,N_8414,N_8756);
nand U11610 (N_11610,N_9812,N_9436);
nand U11611 (N_11611,N_8490,N_7866);
and U11612 (N_11612,N_9820,N_7713);
and U11613 (N_11613,N_8363,N_9285);
and U11614 (N_11614,N_9912,N_9445);
nand U11615 (N_11615,N_7652,N_7505);
nand U11616 (N_11616,N_9679,N_8447);
xor U11617 (N_11617,N_9696,N_8899);
xnor U11618 (N_11618,N_9580,N_8424);
and U11619 (N_11619,N_8966,N_9403);
or U11620 (N_11620,N_8570,N_9935);
xnor U11621 (N_11621,N_9333,N_8897);
nor U11622 (N_11622,N_8723,N_7550);
and U11623 (N_11623,N_9122,N_9749);
nand U11624 (N_11624,N_9371,N_7993);
xor U11625 (N_11625,N_9699,N_8885);
xor U11626 (N_11626,N_8717,N_8668);
and U11627 (N_11627,N_7853,N_7509);
nand U11628 (N_11628,N_8840,N_9218);
nor U11629 (N_11629,N_9813,N_9658);
and U11630 (N_11630,N_8833,N_8655);
nand U11631 (N_11631,N_9560,N_9197);
xnor U11632 (N_11632,N_9006,N_9464);
nor U11633 (N_11633,N_9951,N_9034);
and U11634 (N_11634,N_8805,N_9354);
or U11635 (N_11635,N_7789,N_8133);
nor U11636 (N_11636,N_7895,N_8356);
or U11637 (N_11637,N_8010,N_9339);
nor U11638 (N_11638,N_9396,N_9580);
and U11639 (N_11639,N_9029,N_8134);
nor U11640 (N_11640,N_9402,N_9329);
nand U11641 (N_11641,N_9395,N_9020);
xnor U11642 (N_11642,N_9542,N_9800);
and U11643 (N_11643,N_9461,N_8695);
or U11644 (N_11644,N_9289,N_8879);
and U11645 (N_11645,N_8305,N_8386);
nand U11646 (N_11646,N_9618,N_8273);
nor U11647 (N_11647,N_9968,N_8167);
or U11648 (N_11648,N_8976,N_9292);
and U11649 (N_11649,N_9146,N_7701);
and U11650 (N_11650,N_8787,N_9559);
or U11651 (N_11651,N_8811,N_9979);
xnor U11652 (N_11652,N_8386,N_9119);
nor U11653 (N_11653,N_8313,N_7591);
nor U11654 (N_11654,N_7638,N_8827);
and U11655 (N_11655,N_9920,N_9685);
nor U11656 (N_11656,N_9253,N_9054);
xor U11657 (N_11657,N_8997,N_8501);
xor U11658 (N_11658,N_8349,N_8216);
nor U11659 (N_11659,N_9788,N_9302);
nor U11660 (N_11660,N_7754,N_9432);
nor U11661 (N_11661,N_9039,N_9902);
xnor U11662 (N_11662,N_8028,N_7819);
nor U11663 (N_11663,N_7850,N_7548);
nor U11664 (N_11664,N_9815,N_7529);
xnor U11665 (N_11665,N_7630,N_8782);
and U11666 (N_11666,N_8923,N_9921);
xnor U11667 (N_11667,N_9122,N_9277);
xnor U11668 (N_11668,N_8644,N_8878);
nor U11669 (N_11669,N_9680,N_9334);
nor U11670 (N_11670,N_8869,N_9913);
xor U11671 (N_11671,N_9303,N_9483);
xor U11672 (N_11672,N_8948,N_7505);
and U11673 (N_11673,N_9305,N_8277);
or U11674 (N_11674,N_9208,N_8919);
nor U11675 (N_11675,N_7697,N_7840);
and U11676 (N_11676,N_9585,N_8769);
nand U11677 (N_11677,N_9256,N_8973);
nor U11678 (N_11678,N_9871,N_9295);
nand U11679 (N_11679,N_8646,N_8383);
xor U11680 (N_11680,N_8897,N_8340);
xor U11681 (N_11681,N_8621,N_8122);
or U11682 (N_11682,N_8224,N_8191);
and U11683 (N_11683,N_8314,N_9309);
nand U11684 (N_11684,N_9301,N_9015);
xnor U11685 (N_11685,N_9754,N_9798);
or U11686 (N_11686,N_8311,N_8526);
or U11687 (N_11687,N_9159,N_9430);
nor U11688 (N_11688,N_9223,N_8256);
or U11689 (N_11689,N_9060,N_9608);
and U11690 (N_11690,N_9326,N_7843);
nand U11691 (N_11691,N_7741,N_8798);
nor U11692 (N_11692,N_8497,N_7646);
or U11693 (N_11693,N_9558,N_9977);
or U11694 (N_11694,N_7892,N_7779);
nor U11695 (N_11695,N_7809,N_9711);
or U11696 (N_11696,N_7728,N_7768);
nand U11697 (N_11697,N_7772,N_8266);
nor U11698 (N_11698,N_7979,N_8884);
xnor U11699 (N_11699,N_8699,N_7512);
or U11700 (N_11700,N_9006,N_8145);
nor U11701 (N_11701,N_9284,N_9004);
or U11702 (N_11702,N_8850,N_9919);
nand U11703 (N_11703,N_9805,N_8045);
and U11704 (N_11704,N_7785,N_8193);
or U11705 (N_11705,N_7992,N_7649);
or U11706 (N_11706,N_9616,N_8425);
and U11707 (N_11707,N_9828,N_9927);
nand U11708 (N_11708,N_7526,N_7933);
nand U11709 (N_11709,N_8605,N_8095);
and U11710 (N_11710,N_8208,N_8242);
or U11711 (N_11711,N_7828,N_8087);
nor U11712 (N_11712,N_9462,N_8361);
and U11713 (N_11713,N_8703,N_9777);
nor U11714 (N_11714,N_7694,N_9271);
xor U11715 (N_11715,N_8742,N_8237);
nor U11716 (N_11716,N_9790,N_7969);
or U11717 (N_11717,N_7716,N_8029);
and U11718 (N_11718,N_8229,N_7767);
nor U11719 (N_11719,N_8383,N_8896);
nor U11720 (N_11720,N_8477,N_8017);
nor U11721 (N_11721,N_7665,N_9088);
nand U11722 (N_11722,N_8362,N_8534);
nand U11723 (N_11723,N_9127,N_9519);
xor U11724 (N_11724,N_9453,N_8389);
nand U11725 (N_11725,N_9663,N_8390);
nor U11726 (N_11726,N_8730,N_9988);
xnor U11727 (N_11727,N_9610,N_7540);
nor U11728 (N_11728,N_9999,N_9372);
xnor U11729 (N_11729,N_8661,N_9620);
and U11730 (N_11730,N_7671,N_9151);
and U11731 (N_11731,N_8991,N_9874);
and U11732 (N_11732,N_9470,N_9218);
or U11733 (N_11733,N_8633,N_7888);
nand U11734 (N_11734,N_9473,N_8384);
nand U11735 (N_11735,N_7614,N_7638);
and U11736 (N_11736,N_8146,N_8571);
and U11737 (N_11737,N_8525,N_7557);
nand U11738 (N_11738,N_9604,N_7598);
and U11739 (N_11739,N_8979,N_7757);
nand U11740 (N_11740,N_7761,N_9948);
and U11741 (N_11741,N_9352,N_7869);
and U11742 (N_11742,N_9368,N_8614);
xnor U11743 (N_11743,N_9699,N_9045);
and U11744 (N_11744,N_9153,N_9705);
nand U11745 (N_11745,N_7592,N_9170);
xor U11746 (N_11746,N_7950,N_9368);
nor U11747 (N_11747,N_9880,N_7533);
xnor U11748 (N_11748,N_8114,N_8575);
xor U11749 (N_11749,N_7902,N_9521);
and U11750 (N_11750,N_9689,N_9798);
or U11751 (N_11751,N_8829,N_8143);
or U11752 (N_11752,N_7830,N_7992);
nor U11753 (N_11753,N_7776,N_7832);
nand U11754 (N_11754,N_8620,N_7569);
nor U11755 (N_11755,N_9121,N_9597);
and U11756 (N_11756,N_7793,N_9576);
nand U11757 (N_11757,N_7710,N_9011);
xnor U11758 (N_11758,N_9391,N_8149);
xor U11759 (N_11759,N_9520,N_9722);
and U11760 (N_11760,N_9119,N_7756);
xor U11761 (N_11761,N_7930,N_8768);
or U11762 (N_11762,N_9139,N_8108);
or U11763 (N_11763,N_9765,N_7909);
nor U11764 (N_11764,N_8700,N_9809);
nor U11765 (N_11765,N_9566,N_7927);
nor U11766 (N_11766,N_9692,N_8231);
or U11767 (N_11767,N_9360,N_8036);
xnor U11768 (N_11768,N_7953,N_8703);
and U11769 (N_11769,N_9819,N_8992);
xnor U11770 (N_11770,N_8526,N_9635);
and U11771 (N_11771,N_9753,N_8209);
xnor U11772 (N_11772,N_9480,N_9921);
nand U11773 (N_11773,N_9782,N_9969);
nand U11774 (N_11774,N_9497,N_9306);
and U11775 (N_11775,N_9226,N_8680);
xnor U11776 (N_11776,N_8411,N_9697);
or U11777 (N_11777,N_8440,N_8307);
nand U11778 (N_11778,N_8310,N_9195);
nor U11779 (N_11779,N_7789,N_7811);
nand U11780 (N_11780,N_9858,N_8647);
and U11781 (N_11781,N_7820,N_8464);
nand U11782 (N_11782,N_7874,N_9664);
xor U11783 (N_11783,N_9860,N_7908);
nor U11784 (N_11784,N_8985,N_8118);
and U11785 (N_11785,N_8438,N_8997);
or U11786 (N_11786,N_9669,N_8641);
nand U11787 (N_11787,N_7894,N_9525);
xor U11788 (N_11788,N_8485,N_8196);
or U11789 (N_11789,N_9069,N_9983);
nand U11790 (N_11790,N_8610,N_8450);
nor U11791 (N_11791,N_8001,N_8623);
and U11792 (N_11792,N_8428,N_8007);
xor U11793 (N_11793,N_8217,N_8575);
xor U11794 (N_11794,N_9800,N_7637);
and U11795 (N_11795,N_7645,N_7770);
nand U11796 (N_11796,N_7939,N_9861);
and U11797 (N_11797,N_8295,N_8573);
xnor U11798 (N_11798,N_9701,N_9354);
nor U11799 (N_11799,N_9574,N_9516);
and U11800 (N_11800,N_9297,N_9460);
nor U11801 (N_11801,N_7867,N_8411);
or U11802 (N_11802,N_7626,N_9031);
and U11803 (N_11803,N_9419,N_8101);
xnor U11804 (N_11804,N_9831,N_8251);
nor U11805 (N_11805,N_9460,N_9547);
or U11806 (N_11806,N_7799,N_9508);
nand U11807 (N_11807,N_7670,N_8724);
xnor U11808 (N_11808,N_7849,N_7831);
or U11809 (N_11809,N_7824,N_9604);
nand U11810 (N_11810,N_9245,N_8633);
or U11811 (N_11811,N_7586,N_9248);
nand U11812 (N_11812,N_8196,N_8499);
or U11813 (N_11813,N_9571,N_7531);
or U11814 (N_11814,N_8592,N_9199);
and U11815 (N_11815,N_9921,N_9602);
or U11816 (N_11816,N_9841,N_8330);
xor U11817 (N_11817,N_8366,N_8949);
xnor U11818 (N_11818,N_8914,N_8571);
xnor U11819 (N_11819,N_8030,N_9474);
xnor U11820 (N_11820,N_8072,N_9954);
and U11821 (N_11821,N_7802,N_8568);
xnor U11822 (N_11822,N_7520,N_9944);
and U11823 (N_11823,N_9936,N_8273);
and U11824 (N_11824,N_8760,N_8825);
and U11825 (N_11825,N_9114,N_9597);
xnor U11826 (N_11826,N_9541,N_9893);
and U11827 (N_11827,N_8431,N_8408);
and U11828 (N_11828,N_8936,N_9617);
and U11829 (N_11829,N_7966,N_8365);
xnor U11830 (N_11830,N_8848,N_7916);
xor U11831 (N_11831,N_7678,N_9581);
nor U11832 (N_11832,N_8028,N_8532);
nor U11833 (N_11833,N_8655,N_9332);
nand U11834 (N_11834,N_8522,N_9709);
nor U11835 (N_11835,N_7708,N_8224);
nor U11836 (N_11836,N_8927,N_9543);
nor U11837 (N_11837,N_8012,N_8830);
or U11838 (N_11838,N_9035,N_8492);
nand U11839 (N_11839,N_8272,N_8507);
nand U11840 (N_11840,N_8661,N_8745);
and U11841 (N_11841,N_9910,N_8638);
xor U11842 (N_11842,N_8636,N_7588);
xor U11843 (N_11843,N_7692,N_7635);
and U11844 (N_11844,N_8959,N_7684);
xnor U11845 (N_11845,N_9456,N_8993);
or U11846 (N_11846,N_8327,N_9247);
nand U11847 (N_11847,N_8087,N_8134);
nor U11848 (N_11848,N_9583,N_7767);
xor U11849 (N_11849,N_9210,N_8288);
or U11850 (N_11850,N_8011,N_9498);
xor U11851 (N_11851,N_9200,N_8768);
nor U11852 (N_11852,N_9928,N_9393);
xnor U11853 (N_11853,N_9912,N_9541);
nor U11854 (N_11854,N_9070,N_9162);
nor U11855 (N_11855,N_8627,N_9811);
and U11856 (N_11856,N_8080,N_9347);
and U11857 (N_11857,N_8608,N_8279);
and U11858 (N_11858,N_7686,N_8668);
xnor U11859 (N_11859,N_9625,N_9319);
or U11860 (N_11860,N_7546,N_9052);
and U11861 (N_11861,N_9777,N_7976);
nor U11862 (N_11862,N_8880,N_8156);
xnor U11863 (N_11863,N_9851,N_7976);
nand U11864 (N_11864,N_8162,N_7625);
nor U11865 (N_11865,N_9759,N_9101);
xor U11866 (N_11866,N_8453,N_8396);
or U11867 (N_11867,N_8245,N_8454);
nor U11868 (N_11868,N_9759,N_9829);
nor U11869 (N_11869,N_8083,N_8980);
or U11870 (N_11870,N_9423,N_7933);
xor U11871 (N_11871,N_7894,N_9717);
xor U11872 (N_11872,N_9840,N_9474);
nand U11873 (N_11873,N_9585,N_7965);
and U11874 (N_11874,N_9029,N_8117);
and U11875 (N_11875,N_8906,N_9919);
nor U11876 (N_11876,N_8137,N_7544);
nand U11877 (N_11877,N_7597,N_8207);
and U11878 (N_11878,N_8006,N_9299);
and U11879 (N_11879,N_9161,N_8399);
nand U11880 (N_11880,N_9621,N_8865);
and U11881 (N_11881,N_8271,N_9815);
or U11882 (N_11882,N_7736,N_9544);
and U11883 (N_11883,N_8712,N_9034);
or U11884 (N_11884,N_8195,N_9901);
nand U11885 (N_11885,N_7552,N_8609);
xnor U11886 (N_11886,N_7967,N_9945);
and U11887 (N_11887,N_9190,N_7718);
and U11888 (N_11888,N_7921,N_8957);
nor U11889 (N_11889,N_7577,N_8879);
xor U11890 (N_11890,N_8401,N_8039);
nand U11891 (N_11891,N_7891,N_8961);
nor U11892 (N_11892,N_7527,N_8869);
nand U11893 (N_11893,N_8388,N_9599);
nand U11894 (N_11894,N_7540,N_9673);
xnor U11895 (N_11895,N_9304,N_8177);
nand U11896 (N_11896,N_7884,N_9221);
and U11897 (N_11897,N_7689,N_7881);
nor U11898 (N_11898,N_8853,N_9653);
xnor U11899 (N_11899,N_7931,N_8095);
and U11900 (N_11900,N_9562,N_8378);
or U11901 (N_11901,N_7896,N_7899);
nand U11902 (N_11902,N_9429,N_7934);
xnor U11903 (N_11903,N_9851,N_9099);
xnor U11904 (N_11904,N_7772,N_9368);
nor U11905 (N_11905,N_8371,N_8216);
and U11906 (N_11906,N_8558,N_8455);
or U11907 (N_11907,N_7590,N_9424);
nand U11908 (N_11908,N_9300,N_8888);
xor U11909 (N_11909,N_7624,N_9264);
nand U11910 (N_11910,N_7505,N_7792);
and U11911 (N_11911,N_9670,N_8586);
nand U11912 (N_11912,N_7821,N_8428);
nor U11913 (N_11913,N_8748,N_9220);
nand U11914 (N_11914,N_8903,N_9118);
nor U11915 (N_11915,N_9280,N_8770);
nand U11916 (N_11916,N_9841,N_9707);
nor U11917 (N_11917,N_8517,N_8834);
or U11918 (N_11918,N_7854,N_8311);
and U11919 (N_11919,N_9796,N_9390);
nand U11920 (N_11920,N_8421,N_9102);
nand U11921 (N_11921,N_8628,N_7880);
nor U11922 (N_11922,N_7952,N_8632);
or U11923 (N_11923,N_7807,N_8938);
xor U11924 (N_11924,N_9573,N_9308);
nand U11925 (N_11925,N_8300,N_8283);
or U11926 (N_11926,N_9420,N_9479);
nor U11927 (N_11927,N_9642,N_7667);
and U11928 (N_11928,N_7563,N_7535);
nor U11929 (N_11929,N_9237,N_8658);
nor U11930 (N_11930,N_8309,N_9156);
or U11931 (N_11931,N_8193,N_8768);
xor U11932 (N_11932,N_7580,N_8286);
and U11933 (N_11933,N_8572,N_8662);
and U11934 (N_11934,N_8084,N_8902);
nand U11935 (N_11935,N_8050,N_9409);
nor U11936 (N_11936,N_7796,N_9772);
nor U11937 (N_11937,N_8964,N_9089);
or U11938 (N_11938,N_8551,N_7539);
and U11939 (N_11939,N_8033,N_8759);
nand U11940 (N_11940,N_9036,N_9172);
and U11941 (N_11941,N_9539,N_8817);
or U11942 (N_11942,N_8771,N_7586);
or U11943 (N_11943,N_8497,N_8600);
nand U11944 (N_11944,N_7675,N_7800);
or U11945 (N_11945,N_9467,N_9868);
nand U11946 (N_11946,N_8963,N_8997);
or U11947 (N_11947,N_9279,N_8215);
nand U11948 (N_11948,N_7904,N_8669);
xor U11949 (N_11949,N_7663,N_9422);
xor U11950 (N_11950,N_9472,N_8590);
and U11951 (N_11951,N_7654,N_8357);
nand U11952 (N_11952,N_7805,N_7610);
or U11953 (N_11953,N_8550,N_9555);
and U11954 (N_11954,N_7881,N_9675);
and U11955 (N_11955,N_7554,N_7619);
and U11956 (N_11956,N_8134,N_9890);
nand U11957 (N_11957,N_7632,N_7773);
and U11958 (N_11958,N_9434,N_8406);
xor U11959 (N_11959,N_8550,N_8850);
and U11960 (N_11960,N_7732,N_8237);
xor U11961 (N_11961,N_8478,N_9595);
and U11962 (N_11962,N_8647,N_8815);
and U11963 (N_11963,N_8525,N_8341);
xnor U11964 (N_11964,N_8684,N_9522);
xnor U11965 (N_11965,N_7603,N_9078);
nor U11966 (N_11966,N_9958,N_7509);
and U11967 (N_11967,N_8600,N_9949);
xor U11968 (N_11968,N_9039,N_8505);
nand U11969 (N_11969,N_7800,N_9579);
or U11970 (N_11970,N_9353,N_8772);
or U11971 (N_11971,N_7984,N_9796);
xor U11972 (N_11972,N_9364,N_9241);
xnor U11973 (N_11973,N_9952,N_9622);
xnor U11974 (N_11974,N_7820,N_9537);
and U11975 (N_11975,N_8172,N_9517);
nand U11976 (N_11976,N_8888,N_9798);
or U11977 (N_11977,N_9818,N_8838);
nand U11978 (N_11978,N_8586,N_8804);
nand U11979 (N_11979,N_9075,N_9573);
or U11980 (N_11980,N_7992,N_9642);
xor U11981 (N_11981,N_9982,N_9755);
xnor U11982 (N_11982,N_8501,N_8339);
nor U11983 (N_11983,N_9907,N_9176);
and U11984 (N_11984,N_9417,N_9021);
nor U11985 (N_11985,N_9299,N_9924);
and U11986 (N_11986,N_7673,N_7690);
nand U11987 (N_11987,N_8534,N_8509);
nand U11988 (N_11988,N_8043,N_7634);
or U11989 (N_11989,N_8263,N_9347);
or U11990 (N_11990,N_9710,N_9716);
or U11991 (N_11991,N_9672,N_9229);
or U11992 (N_11992,N_8033,N_7936);
xnor U11993 (N_11993,N_9719,N_9468);
or U11994 (N_11994,N_7520,N_8253);
nor U11995 (N_11995,N_9840,N_8874);
nor U11996 (N_11996,N_7821,N_9617);
nor U11997 (N_11997,N_8282,N_8015);
xor U11998 (N_11998,N_7941,N_8495);
xor U11999 (N_11999,N_8324,N_8454);
nand U12000 (N_12000,N_9702,N_9895);
and U12001 (N_12001,N_8783,N_8927);
xor U12002 (N_12002,N_9525,N_9300);
nor U12003 (N_12003,N_8001,N_8988);
or U12004 (N_12004,N_9699,N_8455);
and U12005 (N_12005,N_8128,N_7695);
or U12006 (N_12006,N_7532,N_8130);
and U12007 (N_12007,N_9275,N_8987);
nand U12008 (N_12008,N_8360,N_9009);
or U12009 (N_12009,N_9608,N_7876);
xnor U12010 (N_12010,N_7765,N_9675);
xnor U12011 (N_12011,N_7612,N_9541);
or U12012 (N_12012,N_9604,N_7506);
xnor U12013 (N_12013,N_8139,N_9251);
or U12014 (N_12014,N_8871,N_8910);
and U12015 (N_12015,N_7761,N_8358);
and U12016 (N_12016,N_9696,N_9093);
nand U12017 (N_12017,N_9250,N_7704);
or U12018 (N_12018,N_9903,N_9855);
nand U12019 (N_12019,N_9094,N_8809);
nor U12020 (N_12020,N_9811,N_7740);
and U12021 (N_12021,N_8676,N_9250);
nand U12022 (N_12022,N_9166,N_8934);
nor U12023 (N_12023,N_8762,N_8368);
xnor U12024 (N_12024,N_9168,N_7629);
nand U12025 (N_12025,N_9665,N_7579);
nor U12026 (N_12026,N_7744,N_8795);
xnor U12027 (N_12027,N_9073,N_8682);
nand U12028 (N_12028,N_9427,N_9515);
nor U12029 (N_12029,N_7858,N_9928);
nor U12030 (N_12030,N_8654,N_8202);
nor U12031 (N_12031,N_9632,N_7516);
nand U12032 (N_12032,N_9688,N_9498);
xnor U12033 (N_12033,N_8339,N_7884);
xnor U12034 (N_12034,N_8319,N_7646);
and U12035 (N_12035,N_9505,N_9354);
xnor U12036 (N_12036,N_9771,N_7625);
xnor U12037 (N_12037,N_9300,N_7876);
and U12038 (N_12038,N_9024,N_9903);
xor U12039 (N_12039,N_9407,N_8401);
and U12040 (N_12040,N_7674,N_8154);
and U12041 (N_12041,N_9191,N_9152);
nor U12042 (N_12042,N_7514,N_9710);
nand U12043 (N_12043,N_8158,N_7780);
and U12044 (N_12044,N_8650,N_9247);
or U12045 (N_12045,N_8178,N_8486);
and U12046 (N_12046,N_9167,N_8115);
xnor U12047 (N_12047,N_7982,N_7890);
nand U12048 (N_12048,N_9086,N_8579);
nand U12049 (N_12049,N_9777,N_9359);
nand U12050 (N_12050,N_7783,N_9639);
nor U12051 (N_12051,N_9355,N_8311);
xnor U12052 (N_12052,N_8172,N_7755);
and U12053 (N_12053,N_8902,N_9719);
nand U12054 (N_12054,N_7556,N_8070);
nand U12055 (N_12055,N_8221,N_8156);
xor U12056 (N_12056,N_8050,N_8324);
nand U12057 (N_12057,N_9070,N_7857);
xnor U12058 (N_12058,N_8539,N_8524);
nor U12059 (N_12059,N_9288,N_7510);
and U12060 (N_12060,N_8709,N_9044);
nor U12061 (N_12061,N_9236,N_8641);
nand U12062 (N_12062,N_9340,N_8327);
nand U12063 (N_12063,N_9023,N_9708);
xnor U12064 (N_12064,N_8870,N_8669);
nor U12065 (N_12065,N_9703,N_9636);
xor U12066 (N_12066,N_9325,N_9901);
nand U12067 (N_12067,N_9295,N_9031);
nand U12068 (N_12068,N_8012,N_7548);
or U12069 (N_12069,N_7943,N_9303);
nor U12070 (N_12070,N_8656,N_7662);
nor U12071 (N_12071,N_8337,N_9386);
or U12072 (N_12072,N_7766,N_9027);
nor U12073 (N_12073,N_8209,N_8373);
xnor U12074 (N_12074,N_9598,N_9502);
xnor U12075 (N_12075,N_9334,N_8572);
nand U12076 (N_12076,N_7759,N_8727);
nor U12077 (N_12077,N_9423,N_8147);
xor U12078 (N_12078,N_9876,N_7564);
nor U12079 (N_12079,N_8103,N_9381);
or U12080 (N_12080,N_7691,N_8331);
nand U12081 (N_12081,N_9213,N_7626);
xnor U12082 (N_12082,N_7926,N_8074);
nor U12083 (N_12083,N_8492,N_8679);
or U12084 (N_12084,N_9761,N_8814);
nand U12085 (N_12085,N_7581,N_9249);
and U12086 (N_12086,N_8680,N_7853);
or U12087 (N_12087,N_9751,N_9718);
or U12088 (N_12088,N_8082,N_7969);
nand U12089 (N_12089,N_8606,N_9498);
nor U12090 (N_12090,N_9873,N_8440);
and U12091 (N_12091,N_9595,N_9587);
nand U12092 (N_12092,N_9866,N_7502);
xor U12093 (N_12093,N_9977,N_9722);
or U12094 (N_12094,N_9301,N_7532);
nor U12095 (N_12095,N_9765,N_9949);
nor U12096 (N_12096,N_8762,N_7811);
or U12097 (N_12097,N_9902,N_9806);
xnor U12098 (N_12098,N_8778,N_9928);
nor U12099 (N_12099,N_8167,N_9601);
nand U12100 (N_12100,N_8162,N_9530);
nor U12101 (N_12101,N_7708,N_8463);
nor U12102 (N_12102,N_7981,N_8903);
xor U12103 (N_12103,N_9346,N_8324);
and U12104 (N_12104,N_9311,N_8782);
nand U12105 (N_12105,N_9842,N_9754);
and U12106 (N_12106,N_9322,N_9129);
or U12107 (N_12107,N_7946,N_9012);
nor U12108 (N_12108,N_9888,N_8339);
xnor U12109 (N_12109,N_8269,N_9214);
nor U12110 (N_12110,N_8616,N_8655);
or U12111 (N_12111,N_9448,N_9720);
nor U12112 (N_12112,N_7877,N_8928);
nor U12113 (N_12113,N_9728,N_9469);
nor U12114 (N_12114,N_8139,N_9423);
nor U12115 (N_12115,N_9445,N_9501);
nand U12116 (N_12116,N_9784,N_8533);
xor U12117 (N_12117,N_8104,N_7983);
or U12118 (N_12118,N_7612,N_9631);
xor U12119 (N_12119,N_8792,N_9834);
nor U12120 (N_12120,N_9908,N_8001);
xnor U12121 (N_12121,N_9841,N_8730);
xnor U12122 (N_12122,N_9244,N_9824);
xor U12123 (N_12123,N_8598,N_9872);
or U12124 (N_12124,N_8020,N_7586);
nor U12125 (N_12125,N_7783,N_9053);
or U12126 (N_12126,N_7602,N_8978);
nor U12127 (N_12127,N_9427,N_9091);
xnor U12128 (N_12128,N_7680,N_9042);
and U12129 (N_12129,N_8271,N_9709);
nand U12130 (N_12130,N_9324,N_7919);
xnor U12131 (N_12131,N_8989,N_9178);
nor U12132 (N_12132,N_9485,N_9671);
or U12133 (N_12133,N_7627,N_8591);
and U12134 (N_12134,N_8208,N_9671);
nand U12135 (N_12135,N_8652,N_7683);
nand U12136 (N_12136,N_9594,N_7644);
nor U12137 (N_12137,N_8512,N_8701);
xnor U12138 (N_12138,N_9874,N_8128);
or U12139 (N_12139,N_9645,N_7808);
nor U12140 (N_12140,N_9330,N_9498);
xor U12141 (N_12141,N_9488,N_8729);
or U12142 (N_12142,N_8571,N_8154);
and U12143 (N_12143,N_8690,N_8283);
or U12144 (N_12144,N_9514,N_8174);
nor U12145 (N_12145,N_8140,N_8203);
or U12146 (N_12146,N_8810,N_8283);
xor U12147 (N_12147,N_9955,N_8018);
xnor U12148 (N_12148,N_9223,N_9232);
and U12149 (N_12149,N_9041,N_9310);
xnor U12150 (N_12150,N_9840,N_9763);
xor U12151 (N_12151,N_9791,N_8545);
xor U12152 (N_12152,N_8897,N_7511);
or U12153 (N_12153,N_9647,N_9250);
or U12154 (N_12154,N_8804,N_8576);
nor U12155 (N_12155,N_8329,N_8131);
nand U12156 (N_12156,N_9632,N_9855);
xor U12157 (N_12157,N_8266,N_8564);
nor U12158 (N_12158,N_8103,N_9612);
or U12159 (N_12159,N_7515,N_8182);
or U12160 (N_12160,N_8502,N_7997);
nor U12161 (N_12161,N_9633,N_8189);
and U12162 (N_12162,N_8607,N_9075);
and U12163 (N_12163,N_7507,N_9858);
or U12164 (N_12164,N_8584,N_8631);
or U12165 (N_12165,N_8564,N_9994);
xnor U12166 (N_12166,N_7792,N_9992);
or U12167 (N_12167,N_9189,N_9879);
xnor U12168 (N_12168,N_8077,N_8348);
nor U12169 (N_12169,N_8288,N_9420);
nor U12170 (N_12170,N_8785,N_7841);
nand U12171 (N_12171,N_8669,N_9123);
and U12172 (N_12172,N_7599,N_8661);
or U12173 (N_12173,N_8229,N_8969);
xor U12174 (N_12174,N_9623,N_9707);
xnor U12175 (N_12175,N_8693,N_7889);
and U12176 (N_12176,N_8245,N_8021);
and U12177 (N_12177,N_7714,N_7655);
and U12178 (N_12178,N_7896,N_8634);
xnor U12179 (N_12179,N_8571,N_9454);
xnor U12180 (N_12180,N_8553,N_9214);
and U12181 (N_12181,N_9819,N_9893);
or U12182 (N_12182,N_7697,N_7524);
xnor U12183 (N_12183,N_9316,N_9795);
and U12184 (N_12184,N_7727,N_8996);
nor U12185 (N_12185,N_7622,N_9826);
nor U12186 (N_12186,N_9506,N_7655);
and U12187 (N_12187,N_7658,N_8447);
and U12188 (N_12188,N_8227,N_9748);
nor U12189 (N_12189,N_8842,N_9059);
nor U12190 (N_12190,N_9410,N_9528);
and U12191 (N_12191,N_9183,N_8648);
xor U12192 (N_12192,N_9655,N_9200);
nor U12193 (N_12193,N_9348,N_8097);
and U12194 (N_12194,N_8231,N_9595);
xor U12195 (N_12195,N_9735,N_8852);
nand U12196 (N_12196,N_8627,N_9902);
or U12197 (N_12197,N_9889,N_7849);
nand U12198 (N_12198,N_7594,N_8061);
nand U12199 (N_12199,N_8971,N_8030);
and U12200 (N_12200,N_9235,N_8914);
nand U12201 (N_12201,N_8898,N_8042);
xnor U12202 (N_12202,N_9169,N_9999);
xnor U12203 (N_12203,N_7528,N_9582);
xor U12204 (N_12204,N_8143,N_8781);
nand U12205 (N_12205,N_9172,N_7738);
or U12206 (N_12206,N_9043,N_9072);
nand U12207 (N_12207,N_8826,N_9722);
nand U12208 (N_12208,N_8726,N_8718);
xor U12209 (N_12209,N_7678,N_9845);
nand U12210 (N_12210,N_9487,N_8416);
and U12211 (N_12211,N_9525,N_9236);
xnor U12212 (N_12212,N_8788,N_7849);
xor U12213 (N_12213,N_7746,N_8514);
nand U12214 (N_12214,N_8864,N_9858);
nand U12215 (N_12215,N_8101,N_9740);
or U12216 (N_12216,N_8530,N_9482);
or U12217 (N_12217,N_7902,N_9159);
nand U12218 (N_12218,N_9534,N_9868);
xor U12219 (N_12219,N_8896,N_9073);
nor U12220 (N_12220,N_8515,N_9703);
nand U12221 (N_12221,N_7983,N_9992);
and U12222 (N_12222,N_9526,N_8524);
or U12223 (N_12223,N_9621,N_9820);
nand U12224 (N_12224,N_7814,N_7745);
nor U12225 (N_12225,N_9333,N_7531);
nor U12226 (N_12226,N_7629,N_7881);
xnor U12227 (N_12227,N_9673,N_7837);
and U12228 (N_12228,N_9857,N_9386);
nand U12229 (N_12229,N_8463,N_8918);
xor U12230 (N_12230,N_9097,N_8946);
nor U12231 (N_12231,N_8482,N_9844);
nand U12232 (N_12232,N_8391,N_7598);
nand U12233 (N_12233,N_8875,N_8019);
nand U12234 (N_12234,N_8147,N_8010);
and U12235 (N_12235,N_9234,N_8523);
or U12236 (N_12236,N_9708,N_8128);
xnor U12237 (N_12237,N_9040,N_9138);
or U12238 (N_12238,N_8913,N_8491);
nor U12239 (N_12239,N_9974,N_7596);
or U12240 (N_12240,N_9480,N_8601);
nand U12241 (N_12241,N_9164,N_8275);
nor U12242 (N_12242,N_9091,N_9932);
xor U12243 (N_12243,N_9591,N_7767);
or U12244 (N_12244,N_7588,N_7787);
and U12245 (N_12245,N_9187,N_9823);
or U12246 (N_12246,N_8516,N_7730);
nand U12247 (N_12247,N_8483,N_9022);
nand U12248 (N_12248,N_8043,N_8193);
xnor U12249 (N_12249,N_9208,N_8522);
or U12250 (N_12250,N_7960,N_9379);
xnor U12251 (N_12251,N_7975,N_9296);
nand U12252 (N_12252,N_8996,N_7756);
xor U12253 (N_12253,N_9143,N_8717);
nand U12254 (N_12254,N_8102,N_8606);
nor U12255 (N_12255,N_8386,N_9741);
and U12256 (N_12256,N_7568,N_8172);
or U12257 (N_12257,N_9454,N_9379);
or U12258 (N_12258,N_7934,N_9609);
xor U12259 (N_12259,N_9565,N_9953);
and U12260 (N_12260,N_9123,N_8394);
nor U12261 (N_12261,N_9908,N_8559);
nand U12262 (N_12262,N_9647,N_7674);
or U12263 (N_12263,N_8492,N_8254);
xnor U12264 (N_12264,N_8957,N_8167);
nand U12265 (N_12265,N_7569,N_9909);
nor U12266 (N_12266,N_7615,N_9095);
xor U12267 (N_12267,N_9367,N_7574);
xnor U12268 (N_12268,N_8138,N_8799);
or U12269 (N_12269,N_9834,N_9581);
or U12270 (N_12270,N_7845,N_8149);
nor U12271 (N_12271,N_8416,N_9817);
and U12272 (N_12272,N_8728,N_8068);
or U12273 (N_12273,N_9907,N_7642);
xor U12274 (N_12274,N_9402,N_9067);
nor U12275 (N_12275,N_9880,N_7916);
nand U12276 (N_12276,N_9492,N_9290);
nand U12277 (N_12277,N_9815,N_8739);
xnor U12278 (N_12278,N_8535,N_9202);
nand U12279 (N_12279,N_9445,N_9274);
nand U12280 (N_12280,N_7953,N_7586);
or U12281 (N_12281,N_8152,N_8760);
nor U12282 (N_12282,N_8315,N_9992);
and U12283 (N_12283,N_8358,N_8324);
or U12284 (N_12284,N_9121,N_8056);
nand U12285 (N_12285,N_9375,N_7973);
xnor U12286 (N_12286,N_7961,N_8966);
xnor U12287 (N_12287,N_8768,N_8926);
and U12288 (N_12288,N_9897,N_8902);
nand U12289 (N_12289,N_9103,N_8233);
xor U12290 (N_12290,N_8970,N_9923);
nand U12291 (N_12291,N_8937,N_9211);
or U12292 (N_12292,N_9485,N_8992);
or U12293 (N_12293,N_9698,N_9185);
and U12294 (N_12294,N_9245,N_8002);
xor U12295 (N_12295,N_7544,N_7914);
and U12296 (N_12296,N_8447,N_9393);
xor U12297 (N_12297,N_8875,N_7924);
xor U12298 (N_12298,N_8640,N_7723);
nand U12299 (N_12299,N_7611,N_8873);
and U12300 (N_12300,N_8087,N_7594);
and U12301 (N_12301,N_7761,N_9634);
nand U12302 (N_12302,N_8555,N_8470);
nor U12303 (N_12303,N_8989,N_7592);
nand U12304 (N_12304,N_9557,N_9167);
nand U12305 (N_12305,N_7717,N_9235);
nand U12306 (N_12306,N_8649,N_7723);
nor U12307 (N_12307,N_7534,N_7642);
nor U12308 (N_12308,N_9309,N_9279);
nand U12309 (N_12309,N_8991,N_9022);
nor U12310 (N_12310,N_8065,N_7687);
xor U12311 (N_12311,N_7721,N_7573);
nand U12312 (N_12312,N_7724,N_9781);
nor U12313 (N_12313,N_7736,N_9266);
and U12314 (N_12314,N_8960,N_9443);
nor U12315 (N_12315,N_8894,N_7992);
or U12316 (N_12316,N_7785,N_9601);
xnor U12317 (N_12317,N_9035,N_8457);
and U12318 (N_12318,N_8273,N_9453);
nand U12319 (N_12319,N_8583,N_8382);
nor U12320 (N_12320,N_9321,N_9503);
or U12321 (N_12321,N_9053,N_9751);
and U12322 (N_12322,N_9544,N_9116);
nor U12323 (N_12323,N_8372,N_9449);
and U12324 (N_12324,N_8164,N_8920);
and U12325 (N_12325,N_9805,N_9446);
xnor U12326 (N_12326,N_7551,N_7634);
and U12327 (N_12327,N_8617,N_7542);
and U12328 (N_12328,N_9510,N_8123);
xor U12329 (N_12329,N_9059,N_9543);
xnor U12330 (N_12330,N_7547,N_7550);
xor U12331 (N_12331,N_7807,N_9181);
and U12332 (N_12332,N_8249,N_8051);
nand U12333 (N_12333,N_8497,N_8903);
and U12334 (N_12334,N_9647,N_7969);
or U12335 (N_12335,N_9503,N_7635);
nor U12336 (N_12336,N_9716,N_9586);
or U12337 (N_12337,N_8195,N_7873);
or U12338 (N_12338,N_9396,N_7598);
and U12339 (N_12339,N_7529,N_9110);
nand U12340 (N_12340,N_8601,N_9391);
xnor U12341 (N_12341,N_8897,N_8541);
nand U12342 (N_12342,N_8729,N_9719);
or U12343 (N_12343,N_9809,N_8971);
or U12344 (N_12344,N_9441,N_9936);
nand U12345 (N_12345,N_8441,N_8139);
or U12346 (N_12346,N_8692,N_9509);
nor U12347 (N_12347,N_8541,N_9626);
xnor U12348 (N_12348,N_9002,N_8739);
or U12349 (N_12349,N_9662,N_8385);
and U12350 (N_12350,N_7539,N_9914);
or U12351 (N_12351,N_9593,N_7688);
nand U12352 (N_12352,N_7696,N_8700);
nor U12353 (N_12353,N_7951,N_9702);
and U12354 (N_12354,N_8315,N_9677);
or U12355 (N_12355,N_9103,N_9449);
or U12356 (N_12356,N_9453,N_9719);
or U12357 (N_12357,N_8240,N_8423);
xor U12358 (N_12358,N_9325,N_8500);
nor U12359 (N_12359,N_9845,N_8306);
nand U12360 (N_12360,N_8837,N_9007);
nor U12361 (N_12361,N_9746,N_9821);
nor U12362 (N_12362,N_8958,N_8511);
nor U12363 (N_12363,N_9996,N_8024);
and U12364 (N_12364,N_9436,N_9483);
xnor U12365 (N_12365,N_9244,N_9830);
and U12366 (N_12366,N_7942,N_9520);
xnor U12367 (N_12367,N_8604,N_7798);
nand U12368 (N_12368,N_8167,N_9744);
or U12369 (N_12369,N_9114,N_9656);
nor U12370 (N_12370,N_9907,N_7817);
and U12371 (N_12371,N_9393,N_7701);
nand U12372 (N_12372,N_8058,N_8368);
or U12373 (N_12373,N_9168,N_8665);
or U12374 (N_12374,N_8972,N_9779);
xnor U12375 (N_12375,N_8650,N_8265);
nand U12376 (N_12376,N_9399,N_9946);
nor U12377 (N_12377,N_8650,N_8615);
xor U12378 (N_12378,N_9670,N_9637);
or U12379 (N_12379,N_9387,N_7850);
and U12380 (N_12380,N_9131,N_7725);
nor U12381 (N_12381,N_8473,N_9918);
nand U12382 (N_12382,N_8132,N_9114);
or U12383 (N_12383,N_9379,N_8378);
nand U12384 (N_12384,N_9483,N_8652);
nand U12385 (N_12385,N_8408,N_9816);
nand U12386 (N_12386,N_8047,N_8967);
xnor U12387 (N_12387,N_7675,N_8422);
xnor U12388 (N_12388,N_9459,N_8121);
nor U12389 (N_12389,N_8960,N_7765);
nor U12390 (N_12390,N_7668,N_7677);
or U12391 (N_12391,N_8776,N_9307);
and U12392 (N_12392,N_7571,N_8228);
or U12393 (N_12393,N_9217,N_8112);
nand U12394 (N_12394,N_8184,N_8717);
nor U12395 (N_12395,N_8355,N_8489);
nor U12396 (N_12396,N_9158,N_9392);
nor U12397 (N_12397,N_7548,N_8481);
nand U12398 (N_12398,N_9491,N_8654);
nand U12399 (N_12399,N_9599,N_9843);
nor U12400 (N_12400,N_8447,N_8095);
xnor U12401 (N_12401,N_8625,N_9845);
or U12402 (N_12402,N_8575,N_8345);
nor U12403 (N_12403,N_8624,N_8676);
or U12404 (N_12404,N_9516,N_8495);
or U12405 (N_12405,N_8912,N_9675);
or U12406 (N_12406,N_9548,N_9546);
xnor U12407 (N_12407,N_9134,N_8389);
xnor U12408 (N_12408,N_9702,N_8154);
nand U12409 (N_12409,N_8128,N_8454);
or U12410 (N_12410,N_9442,N_7642);
nand U12411 (N_12411,N_8373,N_9018);
and U12412 (N_12412,N_7502,N_8148);
nor U12413 (N_12413,N_8683,N_9316);
and U12414 (N_12414,N_7795,N_8458);
nor U12415 (N_12415,N_9390,N_7504);
nand U12416 (N_12416,N_7768,N_9894);
and U12417 (N_12417,N_8842,N_9419);
xnor U12418 (N_12418,N_8668,N_9111);
nor U12419 (N_12419,N_8264,N_9751);
nor U12420 (N_12420,N_8731,N_9612);
nor U12421 (N_12421,N_8292,N_9890);
nand U12422 (N_12422,N_8379,N_7720);
and U12423 (N_12423,N_9335,N_8805);
nor U12424 (N_12424,N_9973,N_8526);
xor U12425 (N_12425,N_9999,N_8003);
xnor U12426 (N_12426,N_9027,N_8030);
xnor U12427 (N_12427,N_9469,N_8222);
and U12428 (N_12428,N_8584,N_9188);
xnor U12429 (N_12429,N_8419,N_8275);
nand U12430 (N_12430,N_7750,N_8242);
and U12431 (N_12431,N_8929,N_9285);
or U12432 (N_12432,N_9053,N_7807);
nand U12433 (N_12433,N_8859,N_9439);
nor U12434 (N_12434,N_9741,N_9220);
or U12435 (N_12435,N_9662,N_9527);
xor U12436 (N_12436,N_7957,N_9910);
or U12437 (N_12437,N_9538,N_9162);
and U12438 (N_12438,N_8409,N_9676);
nand U12439 (N_12439,N_8491,N_9849);
or U12440 (N_12440,N_8986,N_8724);
nor U12441 (N_12441,N_8587,N_9978);
and U12442 (N_12442,N_9079,N_8548);
nor U12443 (N_12443,N_8985,N_8322);
nor U12444 (N_12444,N_9044,N_7618);
nand U12445 (N_12445,N_9813,N_8336);
xnor U12446 (N_12446,N_7661,N_8841);
or U12447 (N_12447,N_7513,N_8641);
xnor U12448 (N_12448,N_8375,N_9479);
nor U12449 (N_12449,N_9352,N_8293);
or U12450 (N_12450,N_7921,N_9117);
nand U12451 (N_12451,N_7950,N_9492);
nand U12452 (N_12452,N_8688,N_8238);
and U12453 (N_12453,N_9701,N_9745);
xnor U12454 (N_12454,N_9334,N_7831);
nor U12455 (N_12455,N_8775,N_9846);
nand U12456 (N_12456,N_8447,N_7743);
and U12457 (N_12457,N_8641,N_8767);
nor U12458 (N_12458,N_8789,N_8485);
xor U12459 (N_12459,N_9401,N_9967);
xor U12460 (N_12460,N_7548,N_8736);
or U12461 (N_12461,N_8441,N_8183);
xnor U12462 (N_12462,N_9467,N_9476);
or U12463 (N_12463,N_9924,N_9845);
nand U12464 (N_12464,N_9402,N_8115);
or U12465 (N_12465,N_8320,N_8719);
xor U12466 (N_12466,N_9550,N_8992);
xnor U12467 (N_12467,N_8714,N_7732);
xor U12468 (N_12468,N_9319,N_9690);
nand U12469 (N_12469,N_9401,N_9969);
nor U12470 (N_12470,N_9891,N_8510);
xnor U12471 (N_12471,N_9357,N_8508);
or U12472 (N_12472,N_9998,N_9195);
or U12473 (N_12473,N_8298,N_8320);
and U12474 (N_12474,N_9820,N_9062);
nand U12475 (N_12475,N_9175,N_9795);
or U12476 (N_12476,N_7832,N_7735);
nand U12477 (N_12477,N_9001,N_9918);
xnor U12478 (N_12478,N_9320,N_9487);
or U12479 (N_12479,N_7567,N_8029);
or U12480 (N_12480,N_7919,N_8321);
nor U12481 (N_12481,N_7755,N_8141);
nand U12482 (N_12482,N_9979,N_8606);
and U12483 (N_12483,N_9824,N_9192);
xor U12484 (N_12484,N_9815,N_7828);
nor U12485 (N_12485,N_8889,N_9107);
xnor U12486 (N_12486,N_9615,N_9923);
nand U12487 (N_12487,N_7656,N_7621);
nand U12488 (N_12488,N_8233,N_8290);
and U12489 (N_12489,N_9646,N_8428);
and U12490 (N_12490,N_8886,N_8140);
and U12491 (N_12491,N_8324,N_8570);
and U12492 (N_12492,N_7651,N_9231);
and U12493 (N_12493,N_7705,N_8462);
nand U12494 (N_12494,N_8186,N_9130);
xnor U12495 (N_12495,N_8058,N_9028);
or U12496 (N_12496,N_8083,N_7775);
xnor U12497 (N_12497,N_9994,N_8261);
xor U12498 (N_12498,N_7793,N_9206);
or U12499 (N_12499,N_9385,N_8151);
nand U12500 (N_12500,N_11000,N_10818);
nand U12501 (N_12501,N_12243,N_12093);
xnor U12502 (N_12502,N_11970,N_10682);
nand U12503 (N_12503,N_12405,N_10422);
or U12504 (N_12504,N_10340,N_11793);
or U12505 (N_12505,N_10401,N_10030);
and U12506 (N_12506,N_10306,N_12477);
and U12507 (N_12507,N_10949,N_11275);
nor U12508 (N_12508,N_12367,N_10527);
nand U12509 (N_12509,N_10877,N_10294);
nand U12510 (N_12510,N_10373,N_12476);
xor U12511 (N_12511,N_11966,N_12497);
and U12512 (N_12512,N_10979,N_11112);
xor U12513 (N_12513,N_10497,N_12046);
nand U12514 (N_12514,N_11483,N_11193);
xnor U12515 (N_12515,N_12107,N_12132);
or U12516 (N_12516,N_11185,N_11202);
nand U12517 (N_12517,N_10663,N_11991);
nand U12518 (N_12518,N_11233,N_10563);
nand U12519 (N_12519,N_10800,N_10515);
or U12520 (N_12520,N_11496,N_11219);
xnor U12521 (N_12521,N_10405,N_11844);
and U12522 (N_12522,N_11684,N_10413);
nand U12523 (N_12523,N_11557,N_11682);
nor U12524 (N_12524,N_11025,N_10417);
or U12525 (N_12525,N_10636,N_12258);
nand U12526 (N_12526,N_12185,N_11169);
nand U12527 (N_12527,N_10133,N_11027);
and U12528 (N_12528,N_10927,N_10074);
or U12529 (N_12529,N_11959,N_11900);
or U12530 (N_12530,N_11377,N_11479);
nor U12531 (N_12531,N_10318,N_11104);
nor U12532 (N_12532,N_11468,N_11034);
nand U12533 (N_12533,N_10247,N_11519);
or U12534 (N_12534,N_10312,N_12004);
nand U12535 (N_12535,N_12293,N_12189);
or U12536 (N_12536,N_10040,N_10073);
or U12537 (N_12537,N_11473,N_11842);
nand U12538 (N_12538,N_10214,N_10208);
and U12539 (N_12539,N_11748,N_12439);
or U12540 (N_12540,N_12340,N_12059);
nor U12541 (N_12541,N_10063,N_11457);
nand U12542 (N_12542,N_12122,N_10322);
and U12543 (N_12543,N_10084,N_10591);
nand U12544 (N_12544,N_12130,N_12074);
or U12545 (N_12545,N_10232,N_12406);
and U12546 (N_12546,N_10275,N_11786);
or U12547 (N_12547,N_10062,N_12193);
and U12548 (N_12548,N_11373,N_12385);
xnor U12549 (N_12549,N_10538,N_11419);
nand U12550 (N_12550,N_12156,N_10910);
nand U12551 (N_12551,N_10414,N_12294);
or U12552 (N_12552,N_10112,N_10940);
and U12553 (N_12553,N_11893,N_11056);
nor U12554 (N_12554,N_11642,N_11766);
xor U12555 (N_12555,N_11646,N_10688);
or U12556 (N_12556,N_11635,N_11880);
nand U12557 (N_12557,N_10824,N_11733);
nor U12558 (N_12558,N_12388,N_11184);
nand U12559 (N_12559,N_11330,N_11234);
nand U12560 (N_12560,N_10242,N_11238);
xor U12561 (N_12561,N_10190,N_12018);
or U12562 (N_12562,N_12273,N_11476);
or U12563 (N_12563,N_12414,N_12263);
and U12564 (N_12564,N_12325,N_11171);
nor U12565 (N_12565,N_10878,N_11804);
or U12566 (N_12566,N_11097,N_10530);
nand U12567 (N_12567,N_11788,N_11870);
or U12568 (N_12568,N_11322,N_10193);
nand U12569 (N_12569,N_10267,N_11658);
nand U12570 (N_12570,N_10119,N_11006);
nor U12571 (N_12571,N_11347,N_10540);
xnor U12572 (N_12572,N_11992,N_11738);
or U12573 (N_12573,N_11720,N_11161);
nor U12574 (N_12574,N_11877,N_10658);
nor U12575 (N_12575,N_11997,N_12037);
xnor U12576 (N_12576,N_11785,N_10633);
nor U12577 (N_12577,N_10158,N_11266);
and U12578 (N_12578,N_10635,N_11407);
nand U12579 (N_12579,N_12011,N_12464);
or U12580 (N_12580,N_11432,N_10192);
nor U12581 (N_12581,N_11976,N_10015);
xnor U12582 (N_12582,N_10713,N_10529);
or U12583 (N_12583,N_11953,N_11618);
nand U12584 (N_12584,N_10196,N_11146);
nor U12585 (N_12585,N_11872,N_10987);
or U12586 (N_12586,N_10123,N_10472);
and U12587 (N_12587,N_12346,N_12114);
nand U12588 (N_12588,N_10924,N_10553);
and U12589 (N_12589,N_11022,N_11349);
or U12590 (N_12590,N_10408,N_10561);
or U12591 (N_12591,N_10539,N_11863);
nor U12592 (N_12592,N_10328,N_10447);
and U12593 (N_12593,N_12136,N_10980);
xnor U12594 (N_12594,N_11704,N_11076);
xor U12595 (N_12595,N_10742,N_10816);
or U12596 (N_12596,N_10227,N_10953);
nand U12597 (N_12597,N_12213,N_10241);
nor U12598 (N_12598,N_10933,N_11866);
xor U12599 (N_12599,N_11497,N_10420);
and U12600 (N_12600,N_10215,N_12111);
or U12601 (N_12601,N_11297,N_11879);
xor U12602 (N_12602,N_11464,N_12327);
xnor U12603 (N_12603,N_11084,N_11606);
or U12604 (N_12604,N_12396,N_12473);
or U12605 (N_12605,N_10850,N_11727);
and U12606 (N_12606,N_11481,N_10695);
xnor U12607 (N_12607,N_11851,N_11749);
or U12608 (N_12608,N_11527,N_11260);
xor U12609 (N_12609,N_12051,N_12053);
nand U12610 (N_12610,N_11320,N_10674);
nand U12611 (N_12611,N_10727,N_10046);
nand U12612 (N_12612,N_11399,N_12375);
or U12613 (N_12613,N_12373,N_11003);
or U12614 (N_12614,N_10519,N_10024);
and U12615 (N_12615,N_10342,N_12479);
or U12616 (N_12616,N_10025,N_10085);
nor U12617 (N_12617,N_10991,N_11968);
nand U12618 (N_12618,N_10929,N_10363);
and U12619 (N_12619,N_12308,N_12088);
or U12620 (N_12620,N_11021,N_10345);
xnor U12621 (N_12621,N_11382,N_11281);
or U12622 (N_12622,N_11050,N_11102);
xnor U12623 (N_12623,N_10205,N_11080);
and U12624 (N_12624,N_11012,N_10153);
nand U12625 (N_12625,N_10070,N_10412);
xor U12626 (N_12626,N_10610,N_10185);
nand U12627 (N_12627,N_10848,N_10533);
or U12628 (N_12628,N_11280,N_11378);
nand U12629 (N_12629,N_10442,N_11036);
nand U12630 (N_12630,N_11743,N_11467);
and U12631 (N_12631,N_10130,N_12007);
and U12632 (N_12632,N_10182,N_12319);
nand U12633 (N_12633,N_11708,N_12324);
and U12634 (N_12634,N_10143,N_12448);
and U12635 (N_12635,N_12409,N_11869);
nand U12636 (N_12636,N_12474,N_11449);
nand U12637 (N_12637,N_10096,N_12389);
and U12638 (N_12638,N_10941,N_10165);
xor U12639 (N_12639,N_12211,N_12177);
nand U12640 (N_12640,N_10840,N_10043);
or U12641 (N_12641,N_11327,N_10579);
nand U12642 (N_12642,N_10932,N_11137);
nor U12643 (N_12643,N_11882,N_12309);
or U12644 (N_12644,N_10194,N_10601);
xnor U12645 (N_12645,N_11676,N_12126);
xor U12646 (N_12646,N_10741,N_11125);
xnor U12647 (N_12647,N_11074,N_11086);
nand U12648 (N_12648,N_12280,N_12371);
and U12649 (N_12649,N_10285,N_12103);
nor U12650 (N_12650,N_12026,N_11532);
nor U12651 (N_12651,N_10726,N_12424);
xor U12652 (N_12652,N_11858,N_10005);
xor U12653 (N_12653,N_11261,N_10917);
or U12654 (N_12654,N_10588,N_10951);
nor U12655 (N_12655,N_10467,N_10817);
nor U12656 (N_12656,N_10260,N_10327);
or U12657 (N_12657,N_12207,N_11552);
xor U12658 (N_12658,N_10673,N_10645);
nor U12659 (N_12659,N_12256,N_11665);
nor U12660 (N_12660,N_12456,N_12174);
and U12661 (N_12661,N_11741,N_10339);
nor U12662 (N_12662,N_10384,N_12173);
nor U12663 (N_12663,N_10534,N_10221);
nand U12664 (N_12664,N_10464,N_10201);
xnor U12665 (N_12665,N_12457,N_11069);
and U12666 (N_12666,N_10549,N_11540);
and U12667 (N_12667,N_11865,N_10289);
nand U12668 (N_12668,N_10487,N_12247);
and U12669 (N_12669,N_11899,N_12119);
and U12670 (N_12670,N_10052,N_11641);
xnor U12671 (N_12671,N_11216,N_12386);
and U12672 (N_12672,N_10048,N_10370);
or U12673 (N_12673,N_10458,N_11747);
nand U12674 (N_12674,N_10469,N_11818);
or U12675 (N_12675,N_11591,N_12246);
xnor U12676 (N_12676,N_11750,N_11368);
xor U12677 (N_12677,N_10268,N_11017);
or U12678 (N_12678,N_12090,N_12337);
or U12679 (N_12679,N_11114,N_10386);
xor U12680 (N_12680,N_11896,N_10081);
and U12681 (N_12681,N_11394,N_10646);
or U12682 (N_12682,N_11987,N_11414);
or U12683 (N_12683,N_11744,N_10863);
xnor U12684 (N_12684,N_10416,N_10775);
nand U12685 (N_12685,N_10685,N_11445);
xnor U12686 (N_12686,N_11052,N_10297);
nor U12687 (N_12687,N_11190,N_10456);
xor U12688 (N_12688,N_12355,N_11242);
nand U12689 (N_12689,N_11290,N_10066);
nand U12690 (N_12690,N_11745,N_11762);
and U12691 (N_12691,N_11311,N_12144);
nand U12692 (N_12692,N_11506,N_11888);
and U12693 (N_12693,N_11580,N_11087);
and U12694 (N_12694,N_10399,N_10429);
xor U12695 (N_12695,N_10856,N_11376);
and U12696 (N_12696,N_11430,N_11400);
nor U12697 (N_12697,N_12267,N_12498);
or U12698 (N_12698,N_11612,N_11735);
nand U12699 (N_12699,N_11918,N_12184);
or U12700 (N_12700,N_11324,N_10441);
xor U12701 (N_12701,N_11107,N_11910);
nand U12702 (N_12702,N_12468,N_12075);
xor U12703 (N_12703,N_11181,N_11650);
or U12704 (N_12704,N_10307,N_12281);
xnor U12705 (N_12705,N_11256,N_11384);
nand U12706 (N_12706,N_10167,N_11323);
and U12707 (N_12707,N_10337,N_10955);
xnor U12708 (N_12708,N_12219,N_10224);
nor U12709 (N_12709,N_11436,N_12290);
or U12710 (N_12710,N_10016,N_11406);
or U12711 (N_12711,N_11862,N_11329);
or U12712 (N_12712,N_10266,N_11636);
and U12713 (N_12713,N_11815,N_10555);
xor U12714 (N_12714,N_12358,N_12086);
nand U12715 (N_12715,N_11699,N_11709);
and U12716 (N_12716,N_10783,N_11828);
xnor U12717 (N_12717,N_11152,N_12368);
nor U12718 (N_12718,N_11032,N_12353);
nand U12719 (N_12719,N_12301,N_10578);
and U12720 (N_12720,N_10630,N_10263);
nand U12721 (N_12721,N_12370,N_11604);
nand U12722 (N_12722,N_10730,N_10317);
xor U12723 (N_12723,N_10526,N_12445);
nand U12724 (N_12724,N_10476,N_12264);
and U12725 (N_12725,N_10675,N_11803);
or U12726 (N_12726,N_10738,N_12049);
nor U12727 (N_12727,N_11802,N_11182);
nor U12728 (N_12728,N_10693,N_10943);
or U12729 (N_12729,N_11537,N_10501);
or U12730 (N_12730,N_11318,N_11031);
nand U12731 (N_12731,N_11974,N_12151);
nor U12732 (N_12732,N_10956,N_11405);
nand U12733 (N_12733,N_11660,N_11617);
xor U12734 (N_12734,N_11939,N_11934);
nand U12735 (N_12735,N_11048,N_10841);
xnor U12736 (N_12736,N_10828,N_10827);
and U12737 (N_12737,N_10159,N_10865);
and U12738 (N_12738,N_10602,N_12435);
or U12739 (N_12739,N_12104,N_11447);
and U12740 (N_12740,N_11028,N_12099);
or U12741 (N_12741,N_10651,N_12228);
and U12742 (N_12742,N_11516,N_11408);
xor U12743 (N_12743,N_11071,N_11353);
xor U12744 (N_12744,N_10976,N_10152);
nand U12745 (N_12745,N_11463,N_11705);
nor U12746 (N_12746,N_10452,N_11060);
nand U12747 (N_12747,N_11906,N_12372);
nor U12748 (N_12748,N_10258,N_12187);
xnor U12749 (N_12749,N_10388,N_11556);
or U12750 (N_12750,N_10985,N_11120);
xor U12751 (N_12751,N_11312,N_11549);
nand U12752 (N_12752,N_10321,N_10057);
or U12753 (N_12753,N_11545,N_10203);
xor U12754 (N_12754,N_11131,N_12205);
or U12755 (N_12755,N_11901,N_11252);
nor U12756 (N_12756,N_10032,N_12029);
and U12757 (N_12757,N_10964,N_11822);
xor U12758 (N_12758,N_10517,N_10836);
nand U12759 (N_12759,N_10436,N_11397);
xor U12760 (N_12760,N_10128,N_11515);
and U12761 (N_12761,N_11587,N_10614);
and U12762 (N_12762,N_11616,N_12128);
nand U12763 (N_12763,N_12387,N_11930);
and U12764 (N_12764,N_10587,N_11841);
or U12765 (N_12765,N_11840,N_12282);
xnor U12766 (N_12766,N_10029,N_10148);
nand U12767 (N_12767,N_11466,N_10483);
or U12768 (N_12768,N_10886,N_12040);
or U12769 (N_12769,N_12223,N_11946);
nor U12770 (N_12770,N_12197,N_12490);
and U12771 (N_12771,N_12050,N_10377);
or U12772 (N_12772,N_10749,N_11799);
or U12773 (N_12773,N_11683,N_11962);
or U12774 (N_12774,N_11791,N_12335);
nor U12775 (N_12775,N_11334,N_11692);
or U12776 (N_12776,N_11434,N_11439);
or U12777 (N_12777,N_10525,N_10724);
or U12778 (N_12778,N_10560,N_10712);
nor U12779 (N_12779,N_12001,N_11885);
xnor U12780 (N_12780,N_10644,N_11702);
xnor U12781 (N_12781,N_10564,N_10831);
and U12782 (N_12782,N_11106,N_11912);
and U12783 (N_12783,N_10522,N_12461);
xnor U12784 (N_12784,N_12254,N_11534);
and U12785 (N_12785,N_10499,N_10619);
and U12786 (N_12786,N_10438,N_10795);
nor U12787 (N_12787,N_10656,N_11800);
or U12788 (N_12788,N_10790,N_11530);
or U12789 (N_12789,N_12240,N_10333);
and U12790 (N_12790,N_10814,N_10315);
and U12791 (N_12791,N_12305,N_11833);
or U12792 (N_12792,N_12449,N_10557);
xor U12793 (N_12793,N_10905,N_10845);
and U12794 (N_12794,N_10049,N_12020);
nand U12795 (N_12795,N_10216,N_11110);
or U12796 (N_12796,N_12291,N_11177);
nand U12797 (N_12797,N_11148,N_10968);
nor U12798 (N_12798,N_11053,N_11894);
xnor U12799 (N_12799,N_11203,N_11095);
or U12800 (N_12800,N_10879,N_10027);
nor U12801 (N_12801,N_11680,N_12403);
nand U12802 (N_12802,N_10565,N_12005);
nand U12803 (N_12803,N_11282,N_11092);
nor U12804 (N_12804,N_11725,N_12338);
and U12805 (N_12805,N_10475,N_12257);
xor U12806 (N_12806,N_12478,N_11949);
nor U12807 (N_12807,N_11528,N_10813);
or U12808 (N_12808,N_11484,N_11787);
nor U12809 (N_12809,N_12454,N_10351);
nand U12810 (N_12810,N_11550,N_11628);
or U12811 (N_12811,N_10625,N_12098);
xnor U12812 (N_12812,N_10038,N_12393);
and U12813 (N_12813,N_11967,N_10142);
nand U12814 (N_12814,N_11622,N_10002);
or U12815 (N_12815,N_11420,N_10972);
nand U12816 (N_12816,N_10240,N_12418);
nor U12817 (N_12817,N_11435,N_10047);
or U12818 (N_12818,N_12462,N_11227);
and U12819 (N_12819,N_10760,N_10776);
and U12820 (N_12820,N_11296,N_12069);
xnor U12821 (N_12821,N_11624,N_12296);
xor U12822 (N_12822,N_10524,N_11990);
or U12823 (N_12823,N_11035,N_10191);
nor U12824 (N_12824,N_12416,N_11569);
or U12825 (N_12825,N_11627,N_11637);
xor U12826 (N_12826,N_11632,N_12276);
and U12827 (N_12827,N_10183,N_12038);
nand U12828 (N_12828,N_11574,N_11663);
xnor U12829 (N_12829,N_11013,N_10108);
and U12830 (N_12830,N_10572,N_10714);
or U12831 (N_12831,N_11147,N_10718);
xor U12832 (N_12832,N_11480,N_12342);
nor U12833 (N_12833,N_10493,N_10786);
nor U12834 (N_12834,N_11426,N_12450);
nand U12835 (N_12835,N_11914,N_12164);
xnor U12836 (N_12836,N_10075,N_11066);
nor U12837 (N_12837,N_12183,N_11994);
or U12838 (N_12838,N_12143,N_12180);
and U12839 (N_12839,N_11208,N_10900);
nor U12840 (N_12840,N_10041,N_11359);
nand U12841 (N_12841,N_11350,N_10236);
nor U12842 (N_12842,N_11999,N_11740);
or U12843 (N_12843,N_11172,N_10514);
xor U12844 (N_12844,N_10734,N_10132);
nor U12845 (N_12845,N_10450,N_10948);
or U12846 (N_12846,N_10906,N_11941);
or U12847 (N_12847,N_11272,N_11546);
nor U12848 (N_12848,N_11456,N_11771);
nor U12849 (N_12849,N_10308,N_11836);
and U12850 (N_12850,N_12350,N_11498);
nor U12851 (N_12851,N_10304,N_11175);
and U12852 (N_12852,N_12226,N_12003);
and U12853 (N_12853,N_11731,N_11767);
nor U12854 (N_12854,N_12106,N_11383);
xnor U12855 (N_12855,N_12420,N_11475);
and U12856 (N_12856,N_11115,N_11387);
or U12857 (N_12857,N_11333,N_12123);
and U12858 (N_12858,N_12313,N_11716);
nand U12859 (N_12859,N_11697,N_10562);
nand U12860 (N_12860,N_12165,N_12369);
nor U12861 (N_12861,N_10107,N_11176);
and U12862 (N_12862,N_11345,N_10789);
or U12863 (N_12863,N_10551,N_10605);
xor U12864 (N_12864,N_11278,N_12494);
or U12865 (N_12865,N_11551,N_11313);
nor U12866 (N_12866,N_10222,N_10832);
nand U12867 (N_12867,N_10282,N_10757);
xor U12868 (N_12868,N_12407,N_10309);
and U12869 (N_12869,N_11908,N_10821);
or U12870 (N_12870,N_10083,N_10770);
and U12871 (N_12871,N_12014,N_12295);
xnor U12872 (N_12872,N_10995,N_11501);
xnor U12873 (N_12873,N_10810,N_11118);
and U12874 (N_12874,N_10058,N_10245);
xor U12875 (N_12875,N_11935,N_11805);
and U12876 (N_12876,N_10690,N_12215);
or U12877 (N_12877,N_10060,N_10931);
or U12878 (N_12878,N_10791,N_12292);
and U12879 (N_12879,N_10782,N_10150);
nand U12880 (N_12880,N_11821,N_10861);
xor U12881 (N_12881,N_10448,N_12285);
or U12882 (N_12882,N_12101,N_10668);
nand U12883 (N_12883,N_12057,N_10833);
nand U12884 (N_12884,N_10647,N_11897);
xnor U12885 (N_12885,N_12070,N_12289);
nor U12886 (N_12886,N_10253,N_11890);
and U12887 (N_12887,N_12467,N_12200);
and U12888 (N_12888,N_10366,N_10763);
or U12889 (N_12889,N_10305,N_11687);
nand U12890 (N_12890,N_12314,N_11562);
or U12891 (N_12891,N_11911,N_10707);
nor U12892 (N_12892,N_10103,N_11427);
nor U12893 (N_12893,N_11082,N_10360);
and U12894 (N_12894,N_12384,N_10854);
or U12895 (N_12895,N_11392,N_12044);
xor U12896 (N_12896,N_11482,N_10488);
nand U12897 (N_12897,N_10138,N_11507);
or U12898 (N_12898,N_10080,N_10589);
or U12899 (N_12899,N_12162,N_10099);
or U12900 (N_12900,N_10396,N_12008);
and U12901 (N_12901,N_10455,N_12283);
or U12902 (N_12902,N_11213,N_11656);
nand U12903 (N_12903,N_10076,N_10485);
nor U12904 (N_12904,N_10952,N_11487);
or U12905 (N_12905,N_12465,N_10039);
nand U12906 (N_12906,N_10755,N_10912);
xnor U12907 (N_12907,N_12013,N_10104);
xor U12908 (N_12908,N_10535,N_10166);
and U12909 (N_12909,N_10957,N_11153);
nand U12910 (N_12910,N_11638,N_10667);
and U12911 (N_12911,N_11640,N_10238);
xnor U12912 (N_12912,N_12031,N_10457);
nor U12913 (N_12913,N_10271,N_10989);
and U12914 (N_12914,N_10117,N_11722);
or U12915 (N_12915,N_11761,N_10352);
xnor U12916 (N_12916,N_11411,N_12469);
and U12917 (N_12917,N_10355,N_11868);
or U12918 (N_12918,N_11211,N_12058);
xor U12919 (N_12919,N_10385,N_11180);
nor U12920 (N_12920,N_12419,N_11343);
nand U12921 (N_12921,N_10872,N_11251);
or U12922 (N_12922,N_10802,N_11288);
nor U12923 (N_12923,N_11763,N_11443);
nand U12924 (N_12924,N_11416,N_10509);
xor U12925 (N_12925,N_12459,N_11909);
xor U12926 (N_12926,N_10744,N_10283);
or U12927 (N_12927,N_11755,N_11143);
nor U12928 (N_12928,N_10178,N_10748);
or U12929 (N_12929,N_11303,N_11919);
or U12930 (N_12930,N_11187,N_10697);
nor U12931 (N_12931,N_12095,N_10965);
or U12932 (N_12932,N_10855,N_11116);
nor U12933 (N_12933,N_12488,N_10761);
and U12934 (N_12934,N_10944,N_12487);
nand U12935 (N_12935,N_10531,N_12146);
or U12936 (N_12936,N_11326,N_10975);
xnor U12937 (N_12937,N_12251,N_10028);
xor U12938 (N_12938,N_10722,N_11905);
and U12939 (N_12939,N_10959,N_10808);
or U12940 (N_12940,N_11239,N_12019);
xnor U12941 (N_12941,N_11404,N_11486);
and U12942 (N_12942,N_11571,N_11752);
and U12943 (N_12943,N_11240,N_10478);
nand U12944 (N_12944,N_10151,N_11328);
and U12945 (N_12945,N_11732,N_10978);
or U12946 (N_12946,N_10508,N_10569);
nand U12947 (N_12947,N_11594,N_11300);
and U12948 (N_12948,N_10197,N_10252);
xnor U12949 (N_12949,N_12427,N_10451);
or U12950 (N_12950,N_10583,N_12030);
or U12951 (N_12951,N_11079,N_12178);
xor U12952 (N_12952,N_11668,N_12400);
and U12953 (N_12953,N_11267,N_11834);
or U12954 (N_12954,N_10437,N_10157);
nand U12955 (N_12955,N_11790,N_10160);
xor U12956 (N_12956,N_10616,N_12115);
xor U12957 (N_12957,N_10703,N_10313);
nor U12958 (N_12958,N_12138,N_11958);
nand U12959 (N_12959,N_10392,N_12209);
nand U12960 (N_12960,N_10585,N_11796);
or U12961 (N_12961,N_11988,N_12304);
xnor U12962 (N_12962,N_12377,N_11491);
nor U12963 (N_12963,N_10402,N_12110);
nand U12964 (N_12964,N_10219,N_11593);
xor U12965 (N_12965,N_10629,N_11871);
nor U12966 (N_12966,N_10461,N_10034);
nor U12967 (N_12967,N_10484,N_10498);
nor U12968 (N_12968,N_11241,N_11521);
xnor U12969 (N_12969,N_12429,N_10421);
or U12970 (N_12970,N_11402,N_10586);
nand U12971 (N_12971,N_10849,N_11985);
nand U12972 (N_12972,N_11932,N_12081);
nand U12973 (N_12973,N_10676,N_11157);
nand U12974 (N_12974,N_11724,N_11448);
nand U12975 (N_12975,N_11465,N_11883);
nand U12976 (N_12976,N_12045,N_10210);
xor U12977 (N_12977,N_12380,N_10834);
nand U12978 (N_12978,N_12278,N_11596);
nand U12979 (N_12979,N_11813,N_11460);
and U12980 (N_12980,N_10835,N_12482);
nor U12981 (N_12981,N_11829,N_12381);
nor U12982 (N_12982,N_12475,N_10390);
or U12983 (N_12983,N_11586,N_10885);
nand U12984 (N_12984,N_11681,N_10554);
or U12985 (N_12985,N_12411,N_10639);
or U12986 (N_12986,N_11209,N_11611);
nand U12987 (N_12987,N_11235,N_12204);
nand U12988 (N_12988,N_11287,N_10725);
and U12989 (N_12989,N_10136,N_10403);
nor U12990 (N_12990,N_10504,N_10938);
and U12991 (N_12991,N_10794,N_11830);
nor U12992 (N_12992,N_11409,N_11986);
nand U12993 (N_12993,N_11943,N_10740);
xnor U12994 (N_12994,N_12000,N_10575);
or U12995 (N_12995,N_12191,N_10882);
and U12996 (N_12996,N_12382,N_11956);
and U12997 (N_12997,N_12425,N_11271);
nand U12998 (N_12998,N_10146,N_12043);
or U12999 (N_12999,N_10164,N_10883);
nand U13000 (N_13000,N_10298,N_12284);
nor U13001 (N_13001,N_12194,N_10110);
and U13002 (N_13002,N_11955,N_10996);
or U13003 (N_13003,N_11924,N_10778);
nor U13004 (N_13004,N_10611,N_10387);
xor U13005 (N_13005,N_11163,N_11533);
nand U13006 (N_13006,N_10866,N_11304);
or U13007 (N_13007,N_10694,N_12230);
xor U13008 (N_13008,N_11695,N_10642);
or U13009 (N_13009,N_10568,N_12176);
nand U13010 (N_13010,N_11352,N_10687);
xor U13011 (N_13011,N_10280,N_10163);
nor U13012 (N_13012,N_12334,N_10513);
and U13013 (N_13013,N_12272,N_11221);
xnor U13014 (N_13014,N_11849,N_12172);
nand U13015 (N_13015,N_12442,N_11938);
and U13016 (N_13016,N_10660,N_12443);
xor U13017 (N_13017,N_11688,N_11217);
and U13018 (N_13018,N_11250,N_11993);
nand U13019 (N_13019,N_10983,N_12299);
nand U13020 (N_13020,N_10440,N_10407);
and U13021 (N_13021,N_10295,N_11773);
or U13022 (N_13022,N_10577,N_12065);
nand U13023 (N_13023,N_11718,N_12078);
or U13024 (N_13024,N_10095,N_11075);
or U13025 (N_13025,N_10358,N_10918);
nor U13026 (N_13026,N_10463,N_11155);
nor U13027 (N_13027,N_11293,N_11584);
or U13028 (N_13028,N_11451,N_10753);
nor U13029 (N_13029,N_11164,N_11054);
xnor U13030 (N_13030,N_12306,N_10705);
or U13031 (N_13031,N_11602,N_12072);
xor U13032 (N_13032,N_11945,N_11831);
nand U13033 (N_13033,N_11362,N_11192);
xnor U13034 (N_13034,N_11122,N_12035);
and U13035 (N_13035,N_10830,N_11237);
xor U13036 (N_13036,N_12436,N_10180);
or U13037 (N_13037,N_10928,N_12440);
or U13038 (N_13038,N_12428,N_11753);
xnor U13039 (N_13039,N_11807,N_11614);
and U13040 (N_13040,N_12466,N_10068);
or U13041 (N_13041,N_10664,N_10632);
and U13042 (N_13042,N_10141,N_10430);
or U13043 (N_13043,N_11096,N_12190);
nor U13044 (N_13044,N_12460,N_11717);
nor U13045 (N_13045,N_10842,N_10762);
xor U13046 (N_13046,N_10823,N_11619);
or U13047 (N_13047,N_11291,N_12259);
nand U13048 (N_13048,N_12232,N_12458);
or U13049 (N_13049,N_10376,N_11369);
nand U13050 (N_13050,N_10100,N_11124);
and U13051 (N_13051,N_11388,N_11620);
xor U13052 (N_13052,N_11666,N_12236);
or U13053 (N_13053,N_12034,N_11294);
and U13054 (N_13054,N_10121,N_10265);
and U13055 (N_13055,N_10011,N_10925);
nand U13056 (N_13056,N_11101,N_12202);
and U13057 (N_13057,N_10186,N_12157);
and U13058 (N_13058,N_10088,N_10672);
nand U13059 (N_13059,N_12109,N_10359);
nand U13060 (N_13060,N_10600,N_10127);
xor U13061 (N_13061,N_11492,N_12198);
and U13062 (N_13062,N_10709,N_11065);
nand U13063 (N_13063,N_10615,N_11895);
xnor U13064 (N_13064,N_11279,N_11931);
xor U13065 (N_13065,N_10570,N_10433);
nor U13066 (N_13066,N_11459,N_10973);
nand U13067 (N_13067,N_12168,N_11979);
and U13068 (N_13068,N_10281,N_10346);
nor U13069 (N_13069,N_10173,N_11564);
or U13070 (N_13070,N_10223,N_11130);
or U13071 (N_13071,N_10168,N_11995);
and U13072 (N_13072,N_11358,N_12056);
xor U13073 (N_13073,N_11262,N_10506);
and U13074 (N_13074,N_11255,N_12201);
xnor U13075 (N_13075,N_10607,N_11973);
and U13076 (N_13076,N_10310,N_10594);
nand U13077 (N_13077,N_11212,N_11810);
nand U13078 (N_13078,N_11670,N_11525);
and U13079 (N_13079,N_11774,N_10348);
xor U13080 (N_13080,N_11707,N_12079);
xnor U13081 (N_13081,N_10174,N_11057);
nand U13082 (N_13082,N_11607,N_11671);
nor U13083 (N_13083,N_10922,N_12066);
nand U13084 (N_13084,N_11264,N_11133);
nand U13085 (N_13085,N_12307,N_11058);
or U13086 (N_13086,N_12260,N_11059);
and U13087 (N_13087,N_12241,N_10907);
nor U13088 (N_13088,N_11928,N_10573);
and U13089 (N_13089,N_10460,N_12329);
nand U13090 (N_13090,N_12485,N_10666);
nor U13091 (N_13091,N_11390,N_12087);
xnor U13092 (N_13092,N_12270,N_10172);
xor U13093 (N_13093,N_11338,N_10206);
xor U13094 (N_13094,N_12404,N_11247);
or U13095 (N_13095,N_12410,N_12206);
and U13096 (N_13096,N_10654,N_11566);
nand U13097 (N_13097,N_11690,N_11371);
or U13098 (N_13098,N_12333,N_11559);
xor U13099 (N_13099,N_11020,N_11218);
xnor U13100 (N_13100,N_11043,N_11644);
nand U13101 (N_13101,N_11342,N_11062);
xor U13102 (N_13102,N_12063,N_11204);
xor U13103 (N_13103,N_10233,N_10244);
xor U13104 (N_13104,N_10091,N_11915);
xnor U13105 (N_13105,N_12084,N_10930);
or U13106 (N_13106,N_10873,N_12235);
xor U13107 (N_13107,N_10393,N_12231);
xor U13108 (N_13108,N_10708,N_10584);
and U13109 (N_13109,N_10053,N_11696);
and U13110 (N_13110,N_10536,N_10768);
or U13111 (N_13111,N_11188,N_11816);
and U13112 (N_13112,N_11088,N_12413);
nor U13113 (N_13113,N_10093,N_12100);
nor U13114 (N_13114,N_10259,N_12366);
nor U13115 (N_13115,N_11957,N_11412);
or U13116 (N_13116,N_10617,N_11067);
or U13117 (N_13117,N_12339,N_10637);
xnor U13118 (N_13118,N_11008,N_10286);
nor U13119 (N_13119,N_11488,N_10913);
xor U13120 (N_13120,N_11270,N_12117);
nand U13121 (N_13121,N_11274,N_10809);
nand U13122 (N_13122,N_10874,N_10251);
nand U13123 (N_13123,N_12395,N_11795);
nand U13124 (N_13124,N_11814,N_10657);
nand U13125 (N_13125,N_11167,N_10179);
nor U13126 (N_13126,N_11710,N_11440);
and U13127 (N_13127,N_11038,N_11356);
and U13128 (N_13128,N_11839,N_10606);
xor U13129 (N_13129,N_10735,N_11140);
and U13130 (N_13130,N_10065,N_11061);
nand U13131 (N_13131,N_10552,N_12356);
and U13132 (N_13132,N_11567,N_10634);
xnor U13133 (N_13133,N_11712,N_10291);
or U13134 (N_13134,N_11070,N_11049);
or U13135 (N_13135,N_10316,N_11554);
and U13136 (N_13136,N_11860,N_11511);
nand U13137 (N_13137,N_10229,N_11573);
nand U13138 (N_13138,N_11100,N_11243);
xor U13139 (N_13139,N_10711,N_11183);
or U13140 (N_13140,N_10510,N_12105);
xor U13141 (N_13141,N_11174,N_11922);
and U13142 (N_13142,N_10037,N_12451);
xor U13143 (N_13143,N_10652,N_11726);
and U13144 (N_13144,N_10087,N_11570);
xnor U13145 (N_13145,N_11662,N_10988);
xnor U13146 (N_13146,N_11113,N_12312);
xor U13147 (N_13147,N_11780,N_10819);
nand U13148 (N_13148,N_10097,N_11981);
xnor U13149 (N_13149,N_10489,N_12227);
and U13150 (N_13150,N_11673,N_10805);
nand U13151 (N_13151,N_10217,N_10875);
and U13152 (N_13152,N_11832,N_10124);
nand U13153 (N_13153,N_11158,N_11433);
xnor U13154 (N_13154,N_11903,N_11429);
nand U13155 (N_13155,N_11454,N_10019);
nand U13156 (N_13156,N_10012,N_11307);
nand U13157 (N_13157,N_10364,N_11269);
and U13158 (N_13158,N_11127,N_11513);
or U13159 (N_13159,N_10631,N_11314);
nand U13160 (N_13160,N_11168,N_10496);
xnor U13161 (N_13161,N_11232,N_10686);
xnor U13162 (N_13162,N_11063,N_12166);
nand U13163 (N_13163,N_10375,N_11357);
nor U13164 (N_13164,N_10623,N_11856);
or U13165 (N_13165,N_11565,N_10332);
and U13166 (N_13166,N_11077,N_10008);
or U13167 (N_13167,N_10077,N_11236);
and U13168 (N_13168,N_12472,N_10902);
xor U13169 (N_13169,N_11595,N_10071);
and U13170 (N_13170,N_11667,N_11625);
nand U13171 (N_13171,N_11889,N_11355);
xnor U13172 (N_13172,N_10374,N_11042);
nor U13173 (N_13173,N_12052,N_10729);
or U13174 (N_13174,N_10279,N_11083);
nor U13175 (N_13175,N_12480,N_11904);
nor U13176 (N_13176,N_11305,N_10443);
xnor U13177 (N_13177,N_10171,N_12447);
xor U13178 (N_13178,N_10916,N_12310);
nand U13179 (N_13179,N_11819,N_12392);
nand U13180 (N_13180,N_11055,N_10270);
and U13181 (N_13181,N_12083,N_11415);
nor U13182 (N_13182,N_11907,N_11878);
nand U13183 (N_13183,N_10147,N_10486);
or U13184 (N_13184,N_10198,N_10580);
or U13185 (N_13185,N_12234,N_12220);
xnor U13186 (N_13186,N_11820,N_12269);
nand U13187 (N_13187,N_11823,N_10170);
or U13188 (N_13188,N_10628,N_12068);
and U13189 (N_13189,N_11228,N_12470);
nand U13190 (N_13190,N_10559,N_11972);
nor U13191 (N_13191,N_11339,N_10303);
and U13192 (N_13192,N_10406,N_12175);
or U13193 (N_13193,N_11916,N_10888);
nor U13194 (N_13194,N_11630,N_10009);
nand U13195 (N_13195,N_11524,N_11129);
nand U13196 (N_13196,N_11782,N_12208);
xor U13197 (N_13197,N_11301,N_12431);
or U13198 (N_13198,N_11536,N_11073);
and U13199 (N_13199,N_11737,N_12318);
nor U13200 (N_13200,N_11853,N_11478);
xor U13201 (N_13201,N_11942,N_11892);
nor U13202 (N_13202,N_10990,N_10765);
nand U13203 (N_13203,N_11577,N_10548);
and U13204 (N_13204,N_10710,N_11039);
and U13205 (N_13205,N_10131,N_12145);
nor U13206 (N_13206,N_11698,N_12222);
nor U13207 (N_13207,N_10626,N_11944);
nand U13208 (N_13208,N_11634,N_11446);
xor U13209 (N_13209,N_11675,N_11452);
xnor U13210 (N_13210,N_10432,N_11655);
and U13211 (N_13211,N_11045,N_11568);
nand U13212 (N_13212,N_10649,N_11186);
or U13213 (N_13213,N_12237,N_12359);
nand U13214 (N_13214,N_10926,N_11876);
nand U13215 (N_13215,N_10934,N_11801);
nand U13216 (N_13216,N_11734,N_11886);
and U13217 (N_13217,N_10301,N_12491);
and U13218 (N_13218,N_11351,N_10444);
xor U13219 (N_13219,N_10671,N_12398);
nor U13220 (N_13220,N_12023,N_12361);
nand U13221 (N_13221,N_10331,N_10700);
nor U13222 (N_13222,N_11678,N_10596);
xor U13223 (N_13223,N_12493,N_10135);
xor U13224 (N_13224,N_10200,N_10184);
xnor U13225 (N_13225,N_11374,N_11162);
nor U13226 (N_13226,N_12321,N_10759);
and U13227 (N_13227,N_11677,N_10792);
xnor U13228 (N_13228,N_10249,N_12134);
and U13229 (N_13229,N_11723,N_10500);
xor U13230 (N_13230,N_11348,N_10323);
and U13231 (N_13231,N_10923,N_11850);
and U13232 (N_13232,N_10064,N_10092);
nor U13233 (N_13233,N_10939,N_12002);
and U13234 (N_13234,N_11441,N_11657);
or U13235 (N_13235,N_11952,N_10825);
xor U13236 (N_13236,N_11651,N_10445);
nand U13237 (N_13237,N_10169,N_10669);
or U13238 (N_13238,N_10395,N_12032);
nand U13239 (N_13239,N_10982,N_10434);
and U13240 (N_13240,N_10627,N_12415);
nor U13241 (N_13241,N_10653,N_12323);
or U13242 (N_13242,N_12154,N_10449);
xor U13243 (N_13243,N_11579,N_11714);
and U13244 (N_13244,N_11123,N_12330);
and U13245 (N_13245,N_12077,N_11845);
or U13246 (N_13246,N_11253,N_10896);
and U13247 (N_13247,N_11341,N_10947);
and U13248 (N_13248,N_11971,N_10994);
or U13249 (N_13249,N_11824,N_12121);
and U13250 (N_13250,N_11510,N_11041);
or U13251 (N_13251,N_10706,N_12492);
xor U13252 (N_13252,N_11393,N_11555);
and U13253 (N_13253,N_11245,N_10428);
or U13254 (N_13254,N_10262,N_11458);
xor U13255 (N_13255,N_12010,N_12374);
nand U13256 (N_13256,N_11703,N_11613);
nand U13257 (N_13257,N_10881,N_10966);
or U13258 (N_13258,N_11259,N_12016);
nand U13259 (N_13259,N_11715,N_11553);
or U13260 (N_13260,N_12390,N_11442);
nor U13261 (N_13261,N_11664,N_12147);
nand U13262 (N_13262,N_12150,N_12006);
and U13263 (N_13263,N_10118,N_10621);
xnor U13264 (N_13264,N_11589,N_11867);
nand U13265 (N_13265,N_12244,N_10851);
and U13266 (N_13266,N_11363,N_10638);
nor U13267 (N_13267,N_12328,N_10004);
or U13268 (N_13268,N_10921,N_11543);
xor U13269 (N_13269,N_10302,N_10784);
and U13270 (N_13270,N_10477,N_10545);
and U13271 (N_13271,N_11609,N_11847);
xnor U13272 (N_13272,N_10264,N_10140);
xnor U13273 (N_13273,N_10471,N_11843);
or U13274 (N_13274,N_10411,N_11170);
nand U13275 (N_13275,N_11044,N_11284);
and U13276 (N_13276,N_11902,N_11588);
and U13277 (N_13277,N_10869,N_12277);
xor U13278 (N_13278,N_10006,N_10807);
nor U13279 (N_13279,N_10347,N_11418);
or U13280 (N_13280,N_11585,N_10176);
nand U13281 (N_13281,N_11535,N_12097);
nand U13282 (N_13282,N_11539,N_11825);
or U13283 (N_13283,N_11423,N_10162);
xnor U13284 (N_13284,N_11948,N_10404);
xnor U13285 (N_13285,N_12089,N_10532);
xor U13286 (N_13286,N_12376,N_10777);
nand U13287 (N_13287,N_11425,N_11495);
nor U13288 (N_13288,N_11653,N_10780);
xnor U13289 (N_13289,N_11265,N_11838);
and U13290 (N_13290,N_12024,N_10255);
or U13291 (N_13291,N_10681,N_11248);
nand U13292 (N_13292,N_10891,N_10520);
and U13293 (N_13293,N_10898,N_10769);
xor U13294 (N_13294,N_12054,N_10593);
xnor U13295 (N_13295,N_11729,N_10299);
or U13296 (N_13296,N_10296,N_10114);
or U13297 (N_13297,N_10511,N_11998);
nand U13298 (N_13298,N_11764,N_11340);
and U13299 (N_13299,N_10622,N_10423);
xnor U13300 (N_13300,N_12199,N_11461);
nand U13301 (N_13301,N_12192,N_11386);
nor U13302 (N_13302,N_10523,N_12484);
xnor U13303 (N_13303,N_11195,N_10661);
xor U13304 (N_13304,N_10752,N_10126);
nand U13305 (N_13305,N_12218,N_12076);
nor U13306 (N_13306,N_12345,N_11751);
and U13307 (N_13307,N_12118,N_10969);
xor U13308 (N_13308,N_10595,N_10018);
xnor U13309 (N_13309,N_12085,N_10723);
nor U13310 (N_13310,N_10779,N_12160);
xnor U13311 (N_13311,N_12463,N_11694);
and U13312 (N_13312,N_10904,N_11030);
and U13313 (N_13313,N_12249,N_11015);
xnor U13314 (N_13314,N_12242,N_11779);
nor U13315 (N_13315,N_11672,N_11354);
nand U13316 (N_13316,N_10847,N_10254);
nand U13317 (N_13317,N_12135,N_10919);
and U13318 (N_13318,N_11933,N_10482);
nor U13319 (N_13319,N_11610,N_10276);
or U13320 (N_13320,N_11179,N_10454);
or U13321 (N_13321,N_11346,N_10620);
xnor U13322 (N_13322,N_11693,N_10597);
or U13323 (N_13323,N_10567,N_12315);
or U13324 (N_13324,N_11002,N_12499);
xor U13325 (N_13325,N_10102,N_10574);
xnor U13326 (N_13326,N_11826,N_12155);
and U13327 (N_13327,N_11700,N_11285);
and U13328 (N_13328,N_11982,N_11547);
xor U13329 (N_13329,N_12379,N_11674);
or U13330 (N_13330,N_11523,N_12159);
or U13331 (N_13331,N_10893,N_12496);
or U13332 (N_13332,N_10803,N_10870);
nand U13333 (N_13333,N_12022,N_10993);
and U13334 (N_13334,N_12274,N_10187);
nor U13335 (N_13335,N_11295,N_11230);
nand U13336 (N_13336,N_10122,N_10698);
xor U13337 (N_13337,N_11531,N_12096);
nand U13338 (N_13338,N_10400,N_10609);
xnor U13339 (N_13339,N_11652,N_10231);
or U13340 (N_13340,N_11605,N_11037);
nand U13341 (N_13341,N_10889,N_10903);
or U13342 (N_13342,N_11951,N_12225);
xor U13343 (N_13343,N_11317,N_11739);
and U13344 (N_13344,N_10678,N_11151);
nor U13345 (N_13345,N_12113,N_11370);
xnor U13346 (N_13346,N_11144,N_10045);
and U13347 (N_13347,N_10970,N_10998);
and U13348 (N_13348,N_10211,N_10648);
nor U13349 (N_13349,N_12248,N_12186);
and U13350 (N_13350,N_10679,N_11648);
nand U13351 (N_13351,N_10890,N_10801);
nor U13352 (N_13352,N_11254,N_10235);
nor U13353 (N_13353,N_10446,N_10007);
nand U13354 (N_13354,N_10894,N_10367);
nor U13355 (N_13355,N_10365,N_11561);
xor U13356 (N_13356,N_11224,N_10079);
nor U13357 (N_13357,N_10202,N_11395);
and U13358 (N_13358,N_11210,N_10608);
nand U13359 (N_13359,N_10897,N_10439);
and U13360 (N_13360,N_10468,N_10257);
xor U13361 (N_13361,N_12326,N_10115);
and U13362 (N_13362,N_12133,N_11462);
nand U13363 (N_13363,N_10737,N_11331);
nor U13364 (N_13364,N_12365,N_10576);
xnor U13365 (N_13365,N_10937,N_10023);
nor U13366 (N_13366,N_11756,N_11875);
nand U13367 (N_13367,N_12179,N_10599);
or U13368 (N_13368,N_10733,N_12255);
nand U13369 (N_13369,N_11921,N_10550);
and U13370 (N_13370,N_11026,N_11051);
nand U13371 (N_13371,N_11582,N_12120);
nand U13372 (N_13372,N_12252,N_12348);
or U13373 (N_13373,N_11139,N_11961);
nand U13374 (N_13374,N_11706,N_10967);
and U13375 (N_13375,N_10341,N_11827);
xnor U13376 (N_13376,N_11367,N_11508);
nand U13377 (N_13377,N_11989,N_10962);
or U13378 (N_13378,N_11887,N_11389);
or U13379 (N_13379,N_12082,N_11940);
xnor U13380 (N_13380,N_11598,N_10228);
and U13381 (N_13381,N_10680,N_10746);
or U13382 (N_13382,N_10431,N_12061);
and U13383 (N_13383,N_12261,N_10188);
and U13384 (N_13384,N_10225,N_10844);
nand U13385 (N_13385,N_11023,N_11608);
nand U13386 (N_13386,N_10492,N_11159);
xnor U13387 (N_13387,N_12444,N_10113);
or U13388 (N_13388,N_11200,N_10382);
or U13389 (N_13389,N_12239,N_12317);
nand U13390 (N_13390,N_11686,N_12336);
nand U13391 (N_13391,N_10691,N_10380);
nor U13392 (N_13392,N_12233,N_10072);
or U13393 (N_13393,N_11196,N_11538);
xor U13394 (N_13394,N_12357,N_11776);
or U13395 (N_13395,N_10721,N_11286);
and U13396 (N_13396,N_11754,N_10343);
xnor U13397 (N_13397,N_12182,N_11214);
nand U13398 (N_13398,N_12412,N_10349);
xor U13399 (N_13399,N_10212,N_11365);
nor U13400 (N_13400,N_10129,N_10839);
and U13401 (N_13401,N_10812,N_12286);
or U13402 (N_13402,N_12402,N_11019);
or U13403 (N_13403,N_11661,N_10003);
nand U13404 (N_13404,N_11713,N_11310);
and U13405 (N_13405,N_10546,N_10799);
nor U13406 (N_13406,N_11806,N_10022);
xor U13407 (N_13407,N_12300,N_11765);
xnor U13408 (N_13408,N_11917,N_10862);
nand U13409 (N_13409,N_11149,N_10204);
and U13410 (N_13410,N_12048,N_10059);
nand U13411 (N_13411,N_11794,N_11855);
nor U13412 (N_13412,N_12495,N_11811);
xor U13413 (N_13413,N_12344,N_11578);
or U13414 (N_13414,N_10785,N_11659);
xnor U13415 (N_13415,N_10837,N_11499);
nand U13416 (N_13416,N_10677,N_11529);
nand U13417 (N_13417,N_10942,N_12455);
nand U13418 (N_13418,N_11009,N_10798);
or U13419 (N_13419,N_10189,N_10479);
or U13420 (N_13420,N_12297,N_12161);
xnor U13421 (N_13421,N_11319,N_10541);
xor U13422 (N_13422,N_12483,N_11789);
nor U13423 (N_13423,N_12210,N_12341);
nand U13424 (N_13424,N_11360,N_10581);
nor U13425 (N_13425,N_10717,N_11859);
nand U13426 (N_13426,N_10415,N_11485);
nand U13427 (N_13427,N_11315,N_11431);
nor U13428 (N_13428,N_11522,N_10427);
nor U13429 (N_13429,N_10269,N_12360);
or U13430 (N_13430,N_10031,N_11450);
nor U13431 (N_13431,N_11257,N_11273);
nor U13432 (N_13432,N_11581,N_12129);
or U13433 (N_13433,N_11583,N_10319);
and U13434 (N_13434,N_10418,N_10507);
or U13435 (N_13435,N_11090,N_10261);
xor U13436 (N_13436,N_10699,N_11004);
xnor U13437 (N_13437,N_12214,N_11518);
nor U13438 (N_13438,N_10256,N_10105);
nor U13439 (N_13439,N_11633,N_10272);
xor U13440 (N_13440,N_10017,N_11719);
or U13441 (N_13441,N_10021,N_12080);
or U13442 (N_13442,N_11222,N_11775);
and U13443 (N_13443,N_10820,N_12217);
or U13444 (N_13444,N_10683,N_12073);
xnor U13445 (N_13445,N_11597,N_11783);
xnor U13446 (N_13446,N_11469,N_10843);
or U13447 (N_13447,N_12212,N_10424);
xnor U13448 (N_13448,N_10234,N_10470);
or U13449 (N_13449,N_10689,N_12288);
xor U13450 (N_13450,N_11244,N_12221);
and U13451 (N_13451,N_10329,N_11385);
nand U13452 (N_13452,N_11316,N_12438);
nand U13453 (N_13453,N_11965,N_12149);
nor U13454 (N_13454,N_10852,N_11424);
nand U13455 (N_13455,N_12195,N_10624);
nor U13456 (N_13456,N_10750,N_11742);
xnor U13457 (N_13457,N_12229,N_11852);
nand U13458 (N_13458,N_10728,N_10116);
and U13459 (N_13459,N_11770,N_10314);
xnor U13460 (N_13460,N_11306,N_10641);
and U13461 (N_13461,N_11344,N_11846);
xor U13462 (N_13462,N_11141,N_10701);
xor U13463 (N_13463,N_11575,N_12092);
xor U13464 (N_13464,N_11422,N_12401);
xnor U13465 (N_13465,N_10859,N_12430);
or U13466 (N_13466,N_11453,N_10901);
xnor U13467 (N_13467,N_11258,N_11592);
nand U13468 (N_13468,N_11493,N_10887);
nor U13469 (N_13469,N_10491,N_10936);
or U13470 (N_13470,N_12015,N_10494);
nand U13471 (N_13471,N_11470,N_10521);
or U13472 (N_13472,N_11505,N_11477);
or U13473 (N_13473,N_12140,N_10981);
and U13474 (N_13474,N_10250,N_10354);
nor U13475 (N_13475,N_11154,N_12152);
nor U13476 (N_13476,N_11558,N_11728);
or U13477 (N_13477,N_11490,N_10590);
and U13478 (N_13478,N_10963,N_11500);
xor U13479 (N_13479,N_11150,N_10111);
and U13480 (N_13480,N_11016,N_12060);
or U13481 (N_13481,N_12108,N_11215);
and U13482 (N_13482,N_11927,N_11757);
or U13483 (N_13483,N_10243,N_10876);
or U13484 (N_13484,N_12298,N_10603);
xor U13485 (N_13485,N_10582,N_12131);
xnor U13486 (N_13486,N_11623,N_11848);
nor U13487 (N_13487,N_12354,N_10013);
xnor U13488 (N_13488,N_12397,N_11117);
and U13489 (N_13489,N_12322,N_11173);
or U13490 (N_13490,N_10665,N_11277);
and U13491 (N_13491,N_12047,N_11165);
nand U13492 (N_13492,N_10324,N_11758);
nor U13493 (N_13493,N_12422,N_11444);
xnor U13494 (N_13494,N_11544,N_10325);
nand U13495 (N_13495,N_11308,N_11298);
or U13496 (N_13496,N_11960,N_11001);
nand U13497 (N_13497,N_10139,N_11891);
or U13498 (N_13498,N_11639,N_12399);
or U13499 (N_13499,N_11132,N_10719);
nand U13500 (N_13500,N_12394,N_10288);
xor U13501 (N_13501,N_10702,N_11166);
nand U13502 (N_13502,N_12017,N_10078);
xnor U13503 (N_13503,N_10378,N_12203);
or U13504 (N_13504,N_10094,N_10481);
xnor U13505 (N_13505,N_10287,N_11380);
xor U13506 (N_13506,N_11679,N_11977);
nor U13507 (N_13507,N_11014,N_10082);
nand U13508 (N_13508,N_11950,N_10815);
or U13509 (N_13509,N_11401,N_10716);
and U13510 (N_13510,N_11223,N_11576);
or U13511 (N_13511,N_10435,N_10984);
nor U13512 (N_13512,N_11768,N_11781);
xnor U13513 (N_13513,N_10273,N_11160);
nand U13514 (N_13514,N_10000,N_10764);
and U13515 (N_13515,N_12347,N_10826);
xnor U13516 (N_13516,N_10774,N_11809);
and U13517 (N_13517,N_10155,N_12127);
or U13518 (N_13518,N_10868,N_11156);
and U13519 (N_13519,N_11375,N_11881);
nor U13520 (N_13520,N_12169,N_10274);
nor U13521 (N_13521,N_11455,N_12094);
xnor U13522 (N_13522,N_11206,N_11379);
nand U13523 (N_13523,N_10860,N_11542);
nand U13524 (N_13524,N_11226,N_10544);
or U13525 (N_13525,N_11134,N_11197);
and U13526 (N_13526,N_10383,N_12158);
xor U13527 (N_13527,N_11548,N_12265);
xor U13528 (N_13528,N_12446,N_10684);
or U13529 (N_13529,N_12139,N_11111);
xnor U13530 (N_13530,N_10935,N_10462);
nor U13531 (N_13531,N_12349,N_10109);
nand U13532 (N_13532,N_10035,N_11064);
xor U13533 (N_13533,N_10731,N_10154);
nand U13534 (N_13534,N_12039,N_10618);
and U13535 (N_13535,N_11601,N_11309);
nor U13536 (N_13536,N_10220,N_12224);
nor U13537 (N_13537,N_11621,N_11873);
and U13538 (N_13538,N_12071,N_10670);
nor U13539 (N_13539,N_11517,N_11837);
nor U13540 (N_13540,N_10954,N_11502);
and U13541 (N_13541,N_10290,N_11520);
xor U13542 (N_13542,N_11207,N_10946);
or U13543 (N_13543,N_10368,N_10495);
and U13544 (N_13544,N_10300,N_10858);
xnor U13545 (N_13545,N_10571,N_12437);
nor U13546 (N_13546,N_11920,N_10914);
nor U13547 (N_13547,N_10822,N_10177);
or U13548 (N_13548,N_12062,N_10207);
xnor U13549 (N_13549,N_10050,N_11085);
xnor U13550 (N_13550,N_10537,N_11108);
nor U13551 (N_13551,N_10106,N_12421);
nor U13552 (N_13552,N_11325,N_11417);
nand U13553 (N_13553,N_10459,N_10089);
xnor U13554 (N_13554,N_11996,N_11471);
nor U13555 (N_13555,N_10001,N_12153);
or U13556 (N_13556,N_10137,N_10864);
and U13557 (N_13557,N_10643,N_10743);
nor U13558 (N_13558,N_11937,N_10311);
nand U13559 (N_13559,N_11136,N_12027);
and U13560 (N_13560,N_10389,N_10992);
or U13561 (N_13561,N_11494,N_11189);
and U13562 (N_13562,N_10067,N_11413);
xor U13563 (N_13563,N_10846,N_10756);
nand U13564 (N_13564,N_11109,N_10248);
xnor U13565 (N_13565,N_12170,N_10604);
nand U13566 (N_13566,N_10381,N_10226);
nand U13567 (N_13567,N_12279,N_11094);
nand U13568 (N_13568,N_10044,N_11010);
nor U13569 (N_13569,N_10758,N_11936);
nand U13570 (N_13570,N_10650,N_11645);
nand U13571 (N_13571,N_10284,N_11590);
and U13572 (N_13572,N_11138,N_11861);
and U13573 (N_13573,N_12250,N_11730);
nand U13574 (N_13574,N_12378,N_11923);
nand U13575 (N_13575,N_10696,N_11337);
or U13576 (N_13576,N_12391,N_10958);
nor U13577 (N_13577,N_12262,N_11194);
nand U13578 (N_13578,N_11798,N_11276);
nor U13579 (N_13579,N_11366,N_10293);
xor U13580 (N_13580,N_10920,N_11145);
nor U13581 (N_13581,N_11603,N_12042);
or U13582 (N_13582,N_10014,N_10426);
or U13583 (N_13583,N_12036,N_10326);
nand U13584 (N_13584,N_12408,N_12188);
nor U13585 (N_13585,N_11336,N_11563);
and U13586 (N_13586,N_10199,N_10356);
nand U13587 (N_13587,N_10556,N_11817);
xor U13588 (N_13588,N_11760,N_11103);
nand U13589 (N_13589,N_10410,N_10098);
or U13590 (N_13590,N_11615,N_10425);
or U13591 (N_13591,N_10503,N_10010);
nand U13592 (N_13592,N_11268,N_12275);
or U13593 (N_13593,N_11526,N_11093);
nand U13594 (N_13594,N_12181,N_12271);
nor U13595 (N_13595,N_11777,N_11778);
nor U13596 (N_13596,N_11135,N_10335);
xor U13597 (N_13597,N_10175,N_12441);
or U13598 (N_13598,N_10277,N_11835);
or U13599 (N_13599,N_10338,N_11142);
or U13600 (N_13600,N_11403,N_11249);
or U13601 (N_13601,N_11797,N_12351);
xnor U13602 (N_13602,N_11007,N_11599);
xor U13603 (N_13603,N_10543,N_10371);
and U13604 (N_13604,N_12171,N_10156);
xnor U13605 (N_13605,N_10394,N_11178);
nand U13606 (N_13606,N_10950,N_11769);
nor U13607 (N_13607,N_11504,N_10986);
and U13608 (N_13608,N_11649,N_10278);
nor U13609 (N_13609,N_11046,N_10033);
nor U13610 (N_13610,N_10061,N_10911);
nor U13611 (N_13611,N_11759,N_12332);
xnor U13612 (N_13612,N_10796,N_12033);
and U13613 (N_13613,N_10884,N_10369);
and U13614 (N_13614,N_11784,N_10945);
nor U13615 (N_13615,N_12481,N_11225);
xnor U13616 (N_13616,N_12041,N_12426);
or U13617 (N_13617,N_11381,N_11398);
and U13618 (N_13618,N_10120,N_12433);
and U13619 (N_13619,N_10806,N_11980);
nand U13620 (N_13620,N_10195,N_11396);
and U13621 (N_13621,N_10542,N_11808);
nand U13622 (N_13622,N_10772,N_11302);
nor U13623 (N_13623,N_10566,N_10218);
xnor U13624 (N_13624,N_10398,N_10787);
and U13625 (N_13625,N_11081,N_10419);
nor U13626 (N_13626,N_12320,N_11654);
or U13627 (N_13627,N_10054,N_10598);
and U13628 (N_13628,N_12364,N_11299);
or U13629 (N_13629,N_10149,N_12352);
or U13630 (N_13630,N_12012,N_11631);
and U13631 (N_13631,N_10101,N_10974);
or U13632 (N_13632,N_11126,N_11541);
nor U13633 (N_13633,N_11018,N_10909);
nand U13634 (N_13634,N_10391,N_10161);
or U13635 (N_13635,N_12112,N_10051);
nor U13636 (N_13636,N_12489,N_10747);
nand U13637 (N_13637,N_10528,N_10320);
xnor U13638 (N_13638,N_11929,N_11954);
xor U13639 (N_13639,N_11229,N_10899);
nor U13640 (N_13640,N_11024,N_10336);
nor U13641 (N_13641,N_12116,N_12142);
and U13642 (N_13642,N_10871,N_10361);
xnor U13643 (N_13643,N_11040,N_11600);
or U13644 (N_13644,N_12028,N_11864);
or U13645 (N_13645,N_10409,N_10915);
or U13646 (N_13646,N_11321,N_11489);
or U13647 (N_13647,N_12303,N_10732);
nor U13648 (N_13648,N_11438,N_10020);
nand U13649 (N_13649,N_10971,N_11978);
or U13650 (N_13650,N_11428,N_11410);
nor U13651 (N_13651,N_12025,N_12021);
xnor U13652 (N_13652,N_10857,N_10739);
nand U13653 (N_13653,N_11068,N_10518);
nor U13654 (N_13654,N_12302,N_12268);
nor U13655 (N_13655,N_10480,N_10895);
or U13656 (N_13656,N_11199,N_10771);
nor U13657 (N_13657,N_10069,N_11263);
xnor U13658 (N_13658,N_10793,N_11246);
xor U13659 (N_13659,N_11033,N_11047);
and U13660 (N_13660,N_10292,N_11746);
or U13661 (N_13661,N_10042,N_10502);
or U13662 (N_13662,N_11098,N_12148);
xnor U13663 (N_13663,N_12434,N_10592);
or U13664 (N_13664,N_11421,N_10811);
xor U13665 (N_13665,N_12363,N_10838);
nand U13666 (N_13666,N_11701,N_11198);
nand U13667 (N_13667,N_10960,N_11089);
xnor U13668 (N_13668,N_11512,N_11560);
nand U13669 (N_13669,N_10999,N_11964);
nor U13670 (N_13670,N_11105,N_11685);
nor U13671 (N_13671,N_11283,N_11857);
nand U13672 (N_13672,N_10330,N_11874);
nand U13673 (N_13673,N_11372,N_11091);
and U13674 (N_13674,N_12137,N_10754);
nor U13675 (N_13675,N_11926,N_10036);
nor U13676 (N_13676,N_10788,N_10613);
nor U13677 (N_13677,N_10829,N_10473);
and U13678 (N_13678,N_12067,N_10908);
xor U13679 (N_13679,N_12266,N_11289);
xnor U13680 (N_13680,N_10892,N_10490);
nor U13681 (N_13681,N_10767,N_11711);
nor U13682 (N_13682,N_10715,N_12064);
nor U13683 (N_13683,N_11884,N_10961);
and U13684 (N_13684,N_10350,N_10751);
xnor U13685 (N_13685,N_11898,N_10655);
and U13686 (N_13686,N_11332,N_12055);
and U13687 (N_13687,N_10362,N_10773);
nand U13688 (N_13688,N_11231,N_10465);
xnor U13689 (N_13689,N_10134,N_12102);
and U13690 (N_13690,N_11514,N_10474);
and U13691 (N_13691,N_12167,N_11643);
nor U13692 (N_13692,N_11335,N_10766);
xnor U13693 (N_13693,N_10246,N_10086);
nor U13694 (N_13694,N_12432,N_10209);
xor U13695 (N_13695,N_10505,N_12287);
nand U13696 (N_13696,N_11119,N_12316);
nor U13697 (N_13697,N_11975,N_10704);
xor U13698 (N_13698,N_12141,N_10453);
nor U13699 (N_13699,N_10213,N_10026);
nor U13700 (N_13700,N_10781,N_11078);
nand U13701 (N_13701,N_12423,N_11913);
nand U13702 (N_13702,N_12238,N_11736);
nand U13703 (N_13703,N_11361,N_12362);
xor U13704 (N_13704,N_11947,N_11201);
and U13705 (N_13705,N_10662,N_11792);
and U13706 (N_13706,N_10344,N_11029);
and U13707 (N_13707,N_10547,N_12163);
or U13708 (N_13708,N_11011,N_11292);
xnor U13709 (N_13709,N_11364,N_11812);
and U13710 (N_13710,N_10055,N_11472);
xor U13711 (N_13711,N_11220,N_11963);
or U13712 (N_13712,N_10612,N_11121);
or U13713 (N_13713,N_10237,N_10145);
or U13714 (N_13714,N_10144,N_11969);
or U13715 (N_13715,N_10880,N_10466);
xnor U13716 (N_13716,N_10125,N_10379);
or U13717 (N_13717,N_11626,N_11647);
nand U13718 (N_13718,N_10090,N_11474);
nand U13719 (N_13719,N_10797,N_12453);
xor U13720 (N_13720,N_11772,N_12343);
xnor U13721 (N_13721,N_11691,N_10372);
and U13722 (N_13722,N_11984,N_10181);
and U13723 (N_13723,N_11391,N_11925);
or U13724 (N_13724,N_10558,N_10512);
nor U13725 (N_13725,N_11854,N_10804);
or U13726 (N_13726,N_11509,N_10239);
or U13727 (N_13727,N_12245,N_10357);
nor U13728 (N_13728,N_11437,N_11689);
and U13729 (N_13729,N_10353,N_10853);
nor U13730 (N_13730,N_10659,N_12009);
xor U13731 (N_13731,N_10056,N_11721);
xnor U13732 (N_13732,N_12311,N_10230);
xnor U13733 (N_13733,N_12124,N_10997);
or U13734 (N_13734,N_11983,N_12417);
nand U13735 (N_13735,N_11072,N_11099);
nor U13736 (N_13736,N_11669,N_10516);
nor U13737 (N_13737,N_11629,N_10720);
nor U13738 (N_13738,N_11503,N_12125);
and U13739 (N_13739,N_11205,N_10977);
nand U13740 (N_13740,N_10692,N_12216);
nor U13741 (N_13741,N_12452,N_11005);
xnor U13742 (N_13742,N_12196,N_12486);
xnor U13743 (N_13743,N_10867,N_11128);
and U13744 (N_13744,N_12331,N_10334);
or U13745 (N_13745,N_10640,N_10397);
nor U13746 (N_13746,N_12091,N_10736);
or U13747 (N_13747,N_11191,N_12253);
nand U13748 (N_13748,N_10745,N_12471);
xor U13749 (N_13749,N_11572,N_12383);
xnor U13750 (N_13750,N_10538,N_11569);
nand U13751 (N_13751,N_10518,N_11173);
or U13752 (N_13752,N_10934,N_11000);
and U13753 (N_13753,N_10025,N_10037);
nor U13754 (N_13754,N_10027,N_11007);
xor U13755 (N_13755,N_11346,N_10476);
or U13756 (N_13756,N_11339,N_11134);
or U13757 (N_13757,N_12236,N_11787);
or U13758 (N_13758,N_12196,N_10872);
nor U13759 (N_13759,N_11885,N_11697);
nand U13760 (N_13760,N_10223,N_10652);
or U13761 (N_13761,N_12028,N_11365);
nor U13762 (N_13762,N_10664,N_11803);
or U13763 (N_13763,N_11543,N_11985);
nor U13764 (N_13764,N_10338,N_10668);
xor U13765 (N_13765,N_10536,N_10858);
and U13766 (N_13766,N_11774,N_11362);
and U13767 (N_13767,N_10651,N_10452);
xor U13768 (N_13768,N_10445,N_10755);
or U13769 (N_13769,N_12302,N_11394);
or U13770 (N_13770,N_11377,N_12362);
xnor U13771 (N_13771,N_10314,N_10666);
xnor U13772 (N_13772,N_11193,N_10820);
nand U13773 (N_13773,N_10641,N_10213);
or U13774 (N_13774,N_10725,N_11459);
nand U13775 (N_13775,N_10520,N_12048);
nor U13776 (N_13776,N_11196,N_11803);
nand U13777 (N_13777,N_12257,N_10887);
or U13778 (N_13778,N_11115,N_10095);
or U13779 (N_13779,N_11241,N_12109);
xor U13780 (N_13780,N_10822,N_10406);
or U13781 (N_13781,N_11575,N_11115);
or U13782 (N_13782,N_12251,N_11233);
nand U13783 (N_13783,N_12150,N_11354);
nand U13784 (N_13784,N_12486,N_12388);
nand U13785 (N_13785,N_12209,N_11067);
nor U13786 (N_13786,N_10471,N_10313);
nand U13787 (N_13787,N_10908,N_11981);
nor U13788 (N_13788,N_10604,N_12432);
and U13789 (N_13789,N_10977,N_10121);
nor U13790 (N_13790,N_10516,N_11963);
nand U13791 (N_13791,N_10501,N_12426);
or U13792 (N_13792,N_11933,N_10591);
nor U13793 (N_13793,N_12342,N_10092);
xnor U13794 (N_13794,N_10087,N_12264);
or U13795 (N_13795,N_11991,N_10586);
xnor U13796 (N_13796,N_10432,N_12062);
nor U13797 (N_13797,N_10911,N_10816);
nor U13798 (N_13798,N_10940,N_11031);
xor U13799 (N_13799,N_12435,N_10524);
xor U13800 (N_13800,N_10853,N_11115);
or U13801 (N_13801,N_11491,N_10158);
or U13802 (N_13802,N_12454,N_11842);
and U13803 (N_13803,N_11587,N_11206);
nand U13804 (N_13804,N_11595,N_11491);
or U13805 (N_13805,N_10044,N_10212);
nand U13806 (N_13806,N_12497,N_10673);
and U13807 (N_13807,N_11385,N_10093);
nand U13808 (N_13808,N_10611,N_12443);
or U13809 (N_13809,N_10576,N_11140);
and U13810 (N_13810,N_11951,N_12059);
nand U13811 (N_13811,N_10135,N_10491);
xnor U13812 (N_13812,N_10281,N_11083);
nand U13813 (N_13813,N_11537,N_10017);
xnor U13814 (N_13814,N_10227,N_10725);
nand U13815 (N_13815,N_10753,N_10132);
xor U13816 (N_13816,N_10400,N_10183);
xor U13817 (N_13817,N_12083,N_10908);
or U13818 (N_13818,N_10536,N_10526);
xnor U13819 (N_13819,N_11499,N_11234);
or U13820 (N_13820,N_11405,N_11095);
or U13821 (N_13821,N_10741,N_10188);
xnor U13822 (N_13822,N_12468,N_10723);
or U13823 (N_13823,N_10660,N_12281);
nor U13824 (N_13824,N_10619,N_10225);
nor U13825 (N_13825,N_11625,N_10501);
nand U13826 (N_13826,N_11989,N_10374);
xor U13827 (N_13827,N_10656,N_12229);
nand U13828 (N_13828,N_10974,N_10548);
and U13829 (N_13829,N_11009,N_10609);
nand U13830 (N_13830,N_10025,N_10537);
or U13831 (N_13831,N_10161,N_12256);
xnor U13832 (N_13832,N_12491,N_10449);
and U13833 (N_13833,N_12343,N_10702);
or U13834 (N_13834,N_11500,N_11529);
nor U13835 (N_13835,N_10303,N_11772);
nand U13836 (N_13836,N_12432,N_11281);
and U13837 (N_13837,N_11619,N_10574);
or U13838 (N_13838,N_11758,N_12460);
and U13839 (N_13839,N_12025,N_10849);
nand U13840 (N_13840,N_12110,N_10835);
nand U13841 (N_13841,N_10943,N_11946);
nor U13842 (N_13842,N_11688,N_11744);
xor U13843 (N_13843,N_11311,N_11758);
nor U13844 (N_13844,N_11218,N_10513);
xnor U13845 (N_13845,N_10409,N_12395);
and U13846 (N_13846,N_11477,N_12057);
xor U13847 (N_13847,N_10256,N_11805);
nand U13848 (N_13848,N_11557,N_11241);
xor U13849 (N_13849,N_12213,N_10846);
nor U13850 (N_13850,N_11346,N_10077);
and U13851 (N_13851,N_11655,N_10002);
or U13852 (N_13852,N_11059,N_10533);
nand U13853 (N_13853,N_11712,N_10407);
xor U13854 (N_13854,N_12421,N_12431);
or U13855 (N_13855,N_11024,N_10490);
or U13856 (N_13856,N_11068,N_11920);
and U13857 (N_13857,N_11549,N_12236);
xnor U13858 (N_13858,N_11693,N_11770);
nor U13859 (N_13859,N_10946,N_12393);
nor U13860 (N_13860,N_10957,N_11757);
nor U13861 (N_13861,N_12342,N_10064);
or U13862 (N_13862,N_12228,N_10033);
nor U13863 (N_13863,N_11656,N_10562);
nor U13864 (N_13864,N_11100,N_10269);
nand U13865 (N_13865,N_11944,N_10425);
or U13866 (N_13866,N_12497,N_11877);
nor U13867 (N_13867,N_11477,N_10245);
nor U13868 (N_13868,N_11868,N_10904);
xor U13869 (N_13869,N_10228,N_10167);
nand U13870 (N_13870,N_11609,N_12359);
or U13871 (N_13871,N_11498,N_11541);
nand U13872 (N_13872,N_10451,N_12102);
nor U13873 (N_13873,N_12299,N_12162);
or U13874 (N_13874,N_12190,N_10223);
xnor U13875 (N_13875,N_11443,N_10902);
or U13876 (N_13876,N_11932,N_10582);
nand U13877 (N_13877,N_12160,N_10989);
and U13878 (N_13878,N_10529,N_10913);
or U13879 (N_13879,N_11841,N_12141);
nand U13880 (N_13880,N_11136,N_10862);
and U13881 (N_13881,N_11450,N_11707);
and U13882 (N_13882,N_11577,N_12106);
xor U13883 (N_13883,N_11396,N_11772);
nor U13884 (N_13884,N_10550,N_11734);
or U13885 (N_13885,N_11528,N_11415);
and U13886 (N_13886,N_10245,N_12331);
or U13887 (N_13887,N_12266,N_11437);
or U13888 (N_13888,N_12331,N_11694);
nor U13889 (N_13889,N_10301,N_10555);
nand U13890 (N_13890,N_10696,N_11737);
nand U13891 (N_13891,N_10087,N_10483);
nor U13892 (N_13892,N_10428,N_11391);
xor U13893 (N_13893,N_10733,N_12281);
nor U13894 (N_13894,N_10565,N_12050);
nor U13895 (N_13895,N_10630,N_10496);
and U13896 (N_13896,N_10733,N_10259);
nor U13897 (N_13897,N_11770,N_12172);
and U13898 (N_13898,N_11910,N_10340);
nand U13899 (N_13899,N_10263,N_12135);
nand U13900 (N_13900,N_12205,N_10484);
xor U13901 (N_13901,N_10803,N_10809);
and U13902 (N_13902,N_10530,N_11292);
or U13903 (N_13903,N_12359,N_11891);
and U13904 (N_13904,N_10332,N_12260);
nand U13905 (N_13905,N_10979,N_11029);
or U13906 (N_13906,N_12467,N_11223);
or U13907 (N_13907,N_11952,N_12471);
xor U13908 (N_13908,N_11729,N_11404);
nor U13909 (N_13909,N_10615,N_12345);
and U13910 (N_13910,N_12361,N_10652);
nor U13911 (N_13911,N_11896,N_11354);
or U13912 (N_13912,N_11464,N_11723);
or U13913 (N_13913,N_11183,N_10146);
or U13914 (N_13914,N_11818,N_10292);
and U13915 (N_13915,N_11175,N_12025);
nand U13916 (N_13916,N_10638,N_11306);
nand U13917 (N_13917,N_10410,N_10226);
or U13918 (N_13918,N_11093,N_10353);
or U13919 (N_13919,N_10768,N_10553);
and U13920 (N_13920,N_11395,N_10637);
nand U13921 (N_13921,N_12103,N_10172);
xor U13922 (N_13922,N_10023,N_10447);
and U13923 (N_13923,N_10304,N_10207);
and U13924 (N_13924,N_10910,N_10469);
xnor U13925 (N_13925,N_11525,N_12394);
nor U13926 (N_13926,N_11784,N_11360);
or U13927 (N_13927,N_11248,N_11957);
nor U13928 (N_13928,N_11613,N_11367);
nand U13929 (N_13929,N_11249,N_12463);
xnor U13930 (N_13930,N_10819,N_10787);
nand U13931 (N_13931,N_10156,N_12429);
nor U13932 (N_13932,N_10471,N_12285);
xnor U13933 (N_13933,N_12178,N_10055);
and U13934 (N_13934,N_11289,N_11373);
or U13935 (N_13935,N_11549,N_10296);
xor U13936 (N_13936,N_10427,N_10631);
and U13937 (N_13937,N_10251,N_10618);
nor U13938 (N_13938,N_12127,N_11279);
xnor U13939 (N_13939,N_11978,N_10772);
nand U13940 (N_13940,N_10386,N_11547);
and U13941 (N_13941,N_10519,N_11529);
nand U13942 (N_13942,N_12195,N_10016);
or U13943 (N_13943,N_10928,N_11049);
nor U13944 (N_13944,N_10118,N_10741);
and U13945 (N_13945,N_10554,N_11577);
and U13946 (N_13946,N_12349,N_10815);
nand U13947 (N_13947,N_10270,N_11714);
nor U13948 (N_13948,N_10861,N_12184);
nor U13949 (N_13949,N_10284,N_10541);
and U13950 (N_13950,N_11396,N_11456);
and U13951 (N_13951,N_11683,N_10695);
and U13952 (N_13952,N_12317,N_11752);
xnor U13953 (N_13953,N_10302,N_11222);
and U13954 (N_13954,N_11313,N_11023);
xnor U13955 (N_13955,N_10290,N_10679);
or U13956 (N_13956,N_11690,N_12179);
nor U13957 (N_13957,N_11438,N_11493);
or U13958 (N_13958,N_11118,N_11329);
or U13959 (N_13959,N_11758,N_12476);
nor U13960 (N_13960,N_11247,N_10532);
nor U13961 (N_13961,N_12365,N_12083);
or U13962 (N_13962,N_11169,N_10114);
nand U13963 (N_13963,N_11434,N_10851);
or U13964 (N_13964,N_10661,N_12353);
nor U13965 (N_13965,N_12187,N_10178);
xor U13966 (N_13966,N_12127,N_10774);
or U13967 (N_13967,N_10425,N_10684);
nand U13968 (N_13968,N_11237,N_10471);
nand U13969 (N_13969,N_11072,N_10175);
nor U13970 (N_13970,N_12483,N_10524);
nor U13971 (N_13971,N_12090,N_11660);
or U13972 (N_13972,N_11060,N_12321);
and U13973 (N_13973,N_10210,N_10628);
and U13974 (N_13974,N_10648,N_10698);
or U13975 (N_13975,N_12345,N_10114);
or U13976 (N_13976,N_10852,N_11874);
xor U13977 (N_13977,N_11021,N_10587);
xor U13978 (N_13978,N_10450,N_10123);
nand U13979 (N_13979,N_12379,N_10701);
and U13980 (N_13980,N_10347,N_12342);
and U13981 (N_13981,N_10783,N_10676);
and U13982 (N_13982,N_10873,N_11984);
and U13983 (N_13983,N_10108,N_11856);
nand U13984 (N_13984,N_10780,N_11819);
xnor U13985 (N_13985,N_11334,N_12214);
xnor U13986 (N_13986,N_12027,N_10273);
or U13987 (N_13987,N_11567,N_12387);
and U13988 (N_13988,N_11824,N_11672);
nand U13989 (N_13989,N_11010,N_10242);
nand U13990 (N_13990,N_10616,N_10338);
nand U13991 (N_13991,N_10541,N_10008);
or U13992 (N_13992,N_11877,N_10669);
nor U13993 (N_13993,N_10751,N_11456);
nor U13994 (N_13994,N_11729,N_10841);
and U13995 (N_13995,N_11707,N_10649);
nor U13996 (N_13996,N_11300,N_10817);
nor U13997 (N_13997,N_11997,N_11181);
and U13998 (N_13998,N_11886,N_11295);
or U13999 (N_13999,N_11327,N_10990);
nand U14000 (N_14000,N_11741,N_12365);
nand U14001 (N_14001,N_10138,N_12356);
nand U14002 (N_14002,N_11961,N_11429);
or U14003 (N_14003,N_11027,N_12439);
nor U14004 (N_14004,N_10712,N_12418);
nand U14005 (N_14005,N_12139,N_10325);
and U14006 (N_14006,N_12223,N_11586);
nand U14007 (N_14007,N_11452,N_10749);
xnor U14008 (N_14008,N_12047,N_10199);
nand U14009 (N_14009,N_10651,N_10546);
and U14010 (N_14010,N_10895,N_12444);
nor U14011 (N_14011,N_10745,N_10655);
xor U14012 (N_14012,N_10966,N_12059);
xnor U14013 (N_14013,N_10360,N_10274);
and U14014 (N_14014,N_11409,N_12304);
nor U14015 (N_14015,N_12084,N_11757);
nand U14016 (N_14016,N_12439,N_10187);
and U14017 (N_14017,N_10229,N_10609);
and U14018 (N_14018,N_11288,N_10176);
nand U14019 (N_14019,N_12135,N_12242);
nand U14020 (N_14020,N_11697,N_11410);
xor U14021 (N_14021,N_10790,N_11749);
or U14022 (N_14022,N_11222,N_11968);
or U14023 (N_14023,N_10074,N_10731);
nor U14024 (N_14024,N_12441,N_11294);
and U14025 (N_14025,N_11797,N_11560);
xor U14026 (N_14026,N_11879,N_11049);
xor U14027 (N_14027,N_11404,N_12217);
and U14028 (N_14028,N_12404,N_11540);
nor U14029 (N_14029,N_10466,N_10853);
nor U14030 (N_14030,N_11556,N_10026);
or U14031 (N_14031,N_10886,N_12069);
and U14032 (N_14032,N_10340,N_11014);
nand U14033 (N_14033,N_11111,N_11498);
or U14034 (N_14034,N_11452,N_12109);
nor U14035 (N_14035,N_10165,N_12127);
nor U14036 (N_14036,N_11047,N_10257);
nand U14037 (N_14037,N_12398,N_11212);
or U14038 (N_14038,N_11150,N_10701);
xnor U14039 (N_14039,N_10653,N_11430);
xnor U14040 (N_14040,N_11534,N_11416);
or U14041 (N_14041,N_10141,N_10288);
or U14042 (N_14042,N_12130,N_12011);
or U14043 (N_14043,N_10092,N_10300);
nor U14044 (N_14044,N_11170,N_11589);
xor U14045 (N_14045,N_12046,N_11989);
nor U14046 (N_14046,N_10096,N_11003);
nor U14047 (N_14047,N_12421,N_11574);
and U14048 (N_14048,N_10135,N_11489);
and U14049 (N_14049,N_11161,N_11559);
or U14050 (N_14050,N_10924,N_10170);
or U14051 (N_14051,N_11197,N_11398);
xor U14052 (N_14052,N_11344,N_11807);
xnor U14053 (N_14053,N_10648,N_10794);
or U14054 (N_14054,N_10460,N_10197);
or U14055 (N_14055,N_10244,N_10811);
and U14056 (N_14056,N_10055,N_10981);
nand U14057 (N_14057,N_11165,N_10323);
and U14058 (N_14058,N_11119,N_11789);
and U14059 (N_14059,N_11211,N_10253);
nand U14060 (N_14060,N_11281,N_10514);
or U14061 (N_14061,N_11094,N_11841);
nor U14062 (N_14062,N_12258,N_12074);
nor U14063 (N_14063,N_11970,N_10317);
nand U14064 (N_14064,N_11801,N_11550);
or U14065 (N_14065,N_11235,N_11869);
xor U14066 (N_14066,N_10786,N_10781);
nor U14067 (N_14067,N_11034,N_10552);
nor U14068 (N_14068,N_12183,N_11027);
or U14069 (N_14069,N_10387,N_12049);
or U14070 (N_14070,N_10264,N_10060);
nand U14071 (N_14071,N_10550,N_10962);
xor U14072 (N_14072,N_10758,N_11473);
nand U14073 (N_14073,N_10080,N_11481);
nor U14074 (N_14074,N_11411,N_12078);
xor U14075 (N_14075,N_10528,N_10612);
or U14076 (N_14076,N_10973,N_11649);
or U14077 (N_14077,N_11071,N_11201);
or U14078 (N_14078,N_11472,N_11228);
or U14079 (N_14079,N_10286,N_11563);
and U14080 (N_14080,N_10686,N_10770);
nand U14081 (N_14081,N_10272,N_11145);
nor U14082 (N_14082,N_11342,N_11216);
nor U14083 (N_14083,N_11867,N_12012);
and U14084 (N_14084,N_11765,N_10453);
nor U14085 (N_14085,N_10219,N_10788);
nor U14086 (N_14086,N_11160,N_11432);
and U14087 (N_14087,N_12029,N_11904);
and U14088 (N_14088,N_12392,N_11786);
nor U14089 (N_14089,N_10009,N_11951);
and U14090 (N_14090,N_10859,N_12273);
and U14091 (N_14091,N_10383,N_12361);
and U14092 (N_14092,N_10292,N_10835);
xnor U14093 (N_14093,N_10756,N_12240);
or U14094 (N_14094,N_10120,N_11819);
xor U14095 (N_14095,N_10099,N_10161);
nand U14096 (N_14096,N_11694,N_12381);
or U14097 (N_14097,N_11234,N_11781);
nand U14098 (N_14098,N_11369,N_12037);
nor U14099 (N_14099,N_11130,N_12286);
nand U14100 (N_14100,N_12257,N_11122);
nand U14101 (N_14101,N_12201,N_12035);
nand U14102 (N_14102,N_10059,N_11003);
nor U14103 (N_14103,N_10008,N_12225);
xnor U14104 (N_14104,N_10411,N_10947);
nor U14105 (N_14105,N_11744,N_10686);
and U14106 (N_14106,N_12376,N_11113);
nor U14107 (N_14107,N_10240,N_11369);
nand U14108 (N_14108,N_10036,N_11035);
nor U14109 (N_14109,N_11481,N_11962);
nand U14110 (N_14110,N_10024,N_10509);
nand U14111 (N_14111,N_12196,N_10397);
and U14112 (N_14112,N_11031,N_10447);
nand U14113 (N_14113,N_12461,N_10471);
xnor U14114 (N_14114,N_12090,N_10699);
nand U14115 (N_14115,N_10736,N_11480);
or U14116 (N_14116,N_11134,N_10738);
and U14117 (N_14117,N_11873,N_11295);
xnor U14118 (N_14118,N_10211,N_10359);
nand U14119 (N_14119,N_10934,N_11977);
xor U14120 (N_14120,N_11177,N_12367);
xnor U14121 (N_14121,N_12399,N_10345);
xnor U14122 (N_14122,N_11696,N_10456);
and U14123 (N_14123,N_10755,N_10827);
and U14124 (N_14124,N_12097,N_11141);
nand U14125 (N_14125,N_10204,N_12316);
or U14126 (N_14126,N_11237,N_11414);
or U14127 (N_14127,N_11676,N_10041);
xor U14128 (N_14128,N_11877,N_10441);
xnor U14129 (N_14129,N_10929,N_10336);
nand U14130 (N_14130,N_12002,N_10807);
xor U14131 (N_14131,N_12047,N_12356);
xor U14132 (N_14132,N_10558,N_10419);
nor U14133 (N_14133,N_11763,N_12081);
and U14134 (N_14134,N_10365,N_10362);
nand U14135 (N_14135,N_11599,N_11210);
and U14136 (N_14136,N_10276,N_11454);
nand U14137 (N_14137,N_11583,N_10737);
nand U14138 (N_14138,N_10743,N_12021);
and U14139 (N_14139,N_11248,N_10313);
nand U14140 (N_14140,N_10913,N_10879);
nor U14141 (N_14141,N_11488,N_11270);
and U14142 (N_14142,N_10953,N_11805);
nand U14143 (N_14143,N_11532,N_10876);
nand U14144 (N_14144,N_11330,N_10743);
xor U14145 (N_14145,N_11566,N_10881);
and U14146 (N_14146,N_10964,N_12067);
nand U14147 (N_14147,N_11083,N_11797);
and U14148 (N_14148,N_11248,N_10345);
or U14149 (N_14149,N_11624,N_11564);
xnor U14150 (N_14150,N_11047,N_10571);
or U14151 (N_14151,N_10662,N_12486);
or U14152 (N_14152,N_12127,N_10773);
nand U14153 (N_14153,N_10102,N_11473);
and U14154 (N_14154,N_10042,N_11460);
xor U14155 (N_14155,N_10747,N_11553);
nor U14156 (N_14156,N_11109,N_10995);
and U14157 (N_14157,N_12164,N_12371);
nand U14158 (N_14158,N_10784,N_12322);
xnor U14159 (N_14159,N_11719,N_11357);
or U14160 (N_14160,N_11777,N_10762);
and U14161 (N_14161,N_10899,N_10810);
nor U14162 (N_14162,N_10025,N_11431);
xnor U14163 (N_14163,N_10591,N_12262);
and U14164 (N_14164,N_11090,N_10643);
or U14165 (N_14165,N_11754,N_11373);
or U14166 (N_14166,N_10178,N_11578);
or U14167 (N_14167,N_11938,N_11185);
nand U14168 (N_14168,N_11188,N_11448);
xor U14169 (N_14169,N_11589,N_10876);
xor U14170 (N_14170,N_10893,N_11043);
nor U14171 (N_14171,N_11672,N_11667);
or U14172 (N_14172,N_10210,N_10911);
and U14173 (N_14173,N_11043,N_11650);
nor U14174 (N_14174,N_12130,N_12019);
and U14175 (N_14175,N_12260,N_10130);
and U14176 (N_14176,N_12000,N_10440);
and U14177 (N_14177,N_10523,N_11761);
nand U14178 (N_14178,N_11239,N_11220);
and U14179 (N_14179,N_10912,N_11641);
and U14180 (N_14180,N_11805,N_10690);
xnor U14181 (N_14181,N_10956,N_11425);
and U14182 (N_14182,N_10495,N_10024);
and U14183 (N_14183,N_11431,N_12093);
and U14184 (N_14184,N_11577,N_11586);
nor U14185 (N_14185,N_10335,N_10461);
and U14186 (N_14186,N_10527,N_11151);
and U14187 (N_14187,N_10914,N_10771);
nand U14188 (N_14188,N_11356,N_11303);
nor U14189 (N_14189,N_12252,N_10018);
and U14190 (N_14190,N_12234,N_11945);
xnor U14191 (N_14191,N_11585,N_10495);
nand U14192 (N_14192,N_12395,N_10331);
xor U14193 (N_14193,N_11836,N_10773);
xor U14194 (N_14194,N_10593,N_11698);
nand U14195 (N_14195,N_11244,N_10739);
nand U14196 (N_14196,N_11122,N_12409);
xnor U14197 (N_14197,N_11506,N_10624);
or U14198 (N_14198,N_10577,N_11374);
xnor U14199 (N_14199,N_11162,N_10750);
nand U14200 (N_14200,N_11672,N_10161);
or U14201 (N_14201,N_10993,N_10966);
nor U14202 (N_14202,N_11906,N_11593);
nand U14203 (N_14203,N_11644,N_12424);
and U14204 (N_14204,N_11482,N_10076);
and U14205 (N_14205,N_12491,N_10576);
nand U14206 (N_14206,N_11189,N_12280);
and U14207 (N_14207,N_10878,N_10963);
nor U14208 (N_14208,N_10200,N_11221);
and U14209 (N_14209,N_12322,N_10377);
and U14210 (N_14210,N_10555,N_12037);
xnor U14211 (N_14211,N_11574,N_11878);
nor U14212 (N_14212,N_12302,N_10313);
nor U14213 (N_14213,N_10367,N_11417);
xnor U14214 (N_14214,N_12402,N_10673);
or U14215 (N_14215,N_10684,N_11260);
and U14216 (N_14216,N_10584,N_12236);
nand U14217 (N_14217,N_10202,N_11083);
xnor U14218 (N_14218,N_11167,N_11024);
or U14219 (N_14219,N_11423,N_10319);
or U14220 (N_14220,N_11810,N_10082);
nand U14221 (N_14221,N_11631,N_11054);
xor U14222 (N_14222,N_11964,N_10325);
nor U14223 (N_14223,N_11450,N_10884);
nor U14224 (N_14224,N_11656,N_11785);
nor U14225 (N_14225,N_12463,N_10800);
nand U14226 (N_14226,N_12470,N_12057);
nor U14227 (N_14227,N_10086,N_11254);
xnor U14228 (N_14228,N_10520,N_10339);
nor U14229 (N_14229,N_10143,N_11649);
nor U14230 (N_14230,N_11186,N_10727);
or U14231 (N_14231,N_11559,N_10286);
and U14232 (N_14232,N_11137,N_12058);
and U14233 (N_14233,N_11127,N_10022);
and U14234 (N_14234,N_12091,N_10898);
or U14235 (N_14235,N_11056,N_11835);
and U14236 (N_14236,N_11367,N_10312);
and U14237 (N_14237,N_12069,N_12355);
and U14238 (N_14238,N_10509,N_10697);
xor U14239 (N_14239,N_11476,N_10128);
or U14240 (N_14240,N_10895,N_11386);
nand U14241 (N_14241,N_10603,N_11107);
xor U14242 (N_14242,N_11643,N_12257);
xor U14243 (N_14243,N_12496,N_10038);
xor U14244 (N_14244,N_12468,N_10369);
nor U14245 (N_14245,N_12013,N_10681);
nand U14246 (N_14246,N_10177,N_10902);
or U14247 (N_14247,N_10360,N_11627);
or U14248 (N_14248,N_11485,N_10075);
nand U14249 (N_14249,N_12094,N_10545);
and U14250 (N_14250,N_10769,N_11835);
nor U14251 (N_14251,N_11840,N_11138);
nand U14252 (N_14252,N_12367,N_11250);
nor U14253 (N_14253,N_10135,N_11385);
nand U14254 (N_14254,N_11674,N_11747);
xor U14255 (N_14255,N_11175,N_11494);
xnor U14256 (N_14256,N_10375,N_10049);
xnor U14257 (N_14257,N_11810,N_11141);
or U14258 (N_14258,N_10250,N_10491);
nand U14259 (N_14259,N_10186,N_12284);
nand U14260 (N_14260,N_10261,N_12363);
or U14261 (N_14261,N_10179,N_11417);
and U14262 (N_14262,N_11742,N_10375);
nand U14263 (N_14263,N_10701,N_10769);
or U14264 (N_14264,N_12338,N_12443);
xnor U14265 (N_14265,N_11744,N_12123);
or U14266 (N_14266,N_11169,N_10337);
or U14267 (N_14267,N_11022,N_11476);
xor U14268 (N_14268,N_10927,N_11812);
nand U14269 (N_14269,N_11174,N_10721);
or U14270 (N_14270,N_11789,N_12219);
nand U14271 (N_14271,N_10886,N_10145);
and U14272 (N_14272,N_11373,N_10002);
xnor U14273 (N_14273,N_12447,N_11806);
xnor U14274 (N_14274,N_10005,N_11810);
nand U14275 (N_14275,N_10151,N_11443);
or U14276 (N_14276,N_11492,N_10100);
or U14277 (N_14277,N_10405,N_10415);
or U14278 (N_14278,N_12024,N_10524);
xnor U14279 (N_14279,N_11880,N_11037);
nor U14280 (N_14280,N_12074,N_12141);
nand U14281 (N_14281,N_10326,N_10053);
or U14282 (N_14282,N_11765,N_11450);
xnor U14283 (N_14283,N_10824,N_12308);
nand U14284 (N_14284,N_10513,N_12041);
and U14285 (N_14285,N_11981,N_11235);
xor U14286 (N_14286,N_11877,N_11871);
nand U14287 (N_14287,N_10384,N_10390);
nand U14288 (N_14288,N_10765,N_12155);
xnor U14289 (N_14289,N_10314,N_10327);
xnor U14290 (N_14290,N_10225,N_12238);
and U14291 (N_14291,N_10072,N_10512);
and U14292 (N_14292,N_11708,N_10533);
and U14293 (N_14293,N_11778,N_10502);
nor U14294 (N_14294,N_10992,N_10907);
xor U14295 (N_14295,N_10312,N_10358);
nand U14296 (N_14296,N_10459,N_11307);
nor U14297 (N_14297,N_10184,N_11630);
xor U14298 (N_14298,N_11792,N_10891);
nor U14299 (N_14299,N_11906,N_10188);
nand U14300 (N_14300,N_12399,N_11844);
xor U14301 (N_14301,N_12416,N_10882);
nand U14302 (N_14302,N_12128,N_11987);
nor U14303 (N_14303,N_10881,N_10688);
xnor U14304 (N_14304,N_10912,N_11604);
nor U14305 (N_14305,N_11832,N_10858);
xnor U14306 (N_14306,N_10963,N_11960);
and U14307 (N_14307,N_11314,N_12107);
xnor U14308 (N_14308,N_10582,N_12324);
and U14309 (N_14309,N_10043,N_11376);
and U14310 (N_14310,N_11041,N_11420);
nor U14311 (N_14311,N_11278,N_10621);
or U14312 (N_14312,N_12108,N_10775);
or U14313 (N_14313,N_12162,N_12314);
nor U14314 (N_14314,N_10985,N_11381);
nand U14315 (N_14315,N_10624,N_11187);
nand U14316 (N_14316,N_10696,N_11834);
nand U14317 (N_14317,N_10700,N_12066);
and U14318 (N_14318,N_11424,N_10509);
nand U14319 (N_14319,N_10306,N_11218);
xnor U14320 (N_14320,N_11772,N_12269);
nand U14321 (N_14321,N_12141,N_10395);
or U14322 (N_14322,N_11104,N_11112);
xnor U14323 (N_14323,N_10983,N_10865);
nand U14324 (N_14324,N_11326,N_11494);
or U14325 (N_14325,N_12486,N_10323);
xnor U14326 (N_14326,N_10756,N_10664);
xor U14327 (N_14327,N_10250,N_10881);
nor U14328 (N_14328,N_11401,N_11155);
and U14329 (N_14329,N_11828,N_10267);
or U14330 (N_14330,N_10758,N_11513);
nor U14331 (N_14331,N_10614,N_12314);
and U14332 (N_14332,N_10294,N_12073);
xor U14333 (N_14333,N_12149,N_11252);
nor U14334 (N_14334,N_12169,N_10493);
or U14335 (N_14335,N_10779,N_11275);
or U14336 (N_14336,N_11807,N_12211);
xnor U14337 (N_14337,N_11438,N_11343);
nand U14338 (N_14338,N_10328,N_11046);
xor U14339 (N_14339,N_10907,N_10765);
xor U14340 (N_14340,N_11657,N_12123);
nor U14341 (N_14341,N_10052,N_10633);
nor U14342 (N_14342,N_11066,N_11501);
nor U14343 (N_14343,N_12124,N_10621);
nor U14344 (N_14344,N_12006,N_11919);
nand U14345 (N_14345,N_10937,N_12170);
nand U14346 (N_14346,N_12341,N_11958);
and U14347 (N_14347,N_10948,N_10497);
nor U14348 (N_14348,N_10105,N_11585);
nand U14349 (N_14349,N_11568,N_11784);
and U14350 (N_14350,N_10731,N_10156);
or U14351 (N_14351,N_12237,N_10052);
xnor U14352 (N_14352,N_11667,N_12268);
xnor U14353 (N_14353,N_11071,N_12094);
or U14354 (N_14354,N_11349,N_11046);
nand U14355 (N_14355,N_12000,N_10209);
nor U14356 (N_14356,N_12216,N_10267);
and U14357 (N_14357,N_10958,N_10876);
and U14358 (N_14358,N_11175,N_11279);
and U14359 (N_14359,N_11964,N_10082);
and U14360 (N_14360,N_10629,N_10706);
or U14361 (N_14361,N_12371,N_10107);
xor U14362 (N_14362,N_12090,N_11163);
nor U14363 (N_14363,N_12005,N_11344);
nand U14364 (N_14364,N_11152,N_10078);
and U14365 (N_14365,N_10655,N_10513);
and U14366 (N_14366,N_11863,N_10428);
and U14367 (N_14367,N_11156,N_11480);
nor U14368 (N_14368,N_11772,N_10613);
or U14369 (N_14369,N_11943,N_10743);
nand U14370 (N_14370,N_10662,N_11610);
and U14371 (N_14371,N_11141,N_10226);
nand U14372 (N_14372,N_10116,N_10197);
nand U14373 (N_14373,N_10578,N_11786);
and U14374 (N_14374,N_10741,N_10969);
nand U14375 (N_14375,N_12310,N_10323);
xor U14376 (N_14376,N_11846,N_12220);
xor U14377 (N_14377,N_11937,N_11557);
nand U14378 (N_14378,N_11265,N_11379);
nand U14379 (N_14379,N_12290,N_10194);
or U14380 (N_14380,N_10850,N_10688);
nor U14381 (N_14381,N_10273,N_10493);
nor U14382 (N_14382,N_11727,N_12292);
and U14383 (N_14383,N_12208,N_11645);
nand U14384 (N_14384,N_10943,N_10094);
and U14385 (N_14385,N_12135,N_11515);
and U14386 (N_14386,N_11988,N_11372);
nand U14387 (N_14387,N_11473,N_10182);
nand U14388 (N_14388,N_10760,N_11064);
xnor U14389 (N_14389,N_12460,N_11464);
and U14390 (N_14390,N_10897,N_11824);
and U14391 (N_14391,N_11777,N_11039);
or U14392 (N_14392,N_10603,N_11586);
nand U14393 (N_14393,N_11239,N_11292);
nand U14394 (N_14394,N_11483,N_12138);
nand U14395 (N_14395,N_11553,N_12068);
nor U14396 (N_14396,N_11155,N_12139);
and U14397 (N_14397,N_12004,N_11524);
nor U14398 (N_14398,N_10904,N_12068);
and U14399 (N_14399,N_12101,N_11165);
or U14400 (N_14400,N_11564,N_11491);
and U14401 (N_14401,N_11622,N_10860);
nor U14402 (N_14402,N_11424,N_10686);
or U14403 (N_14403,N_12106,N_12068);
nor U14404 (N_14404,N_11267,N_11600);
and U14405 (N_14405,N_11125,N_11079);
and U14406 (N_14406,N_11688,N_10770);
xor U14407 (N_14407,N_11243,N_12325);
xnor U14408 (N_14408,N_10374,N_11054);
and U14409 (N_14409,N_11853,N_11364);
xnor U14410 (N_14410,N_10900,N_11639);
nor U14411 (N_14411,N_10390,N_11950);
xor U14412 (N_14412,N_11518,N_11944);
and U14413 (N_14413,N_12489,N_10021);
or U14414 (N_14414,N_10093,N_10336);
and U14415 (N_14415,N_11791,N_11759);
nor U14416 (N_14416,N_11840,N_10872);
nor U14417 (N_14417,N_12129,N_11323);
xnor U14418 (N_14418,N_12185,N_12240);
nor U14419 (N_14419,N_11817,N_11189);
or U14420 (N_14420,N_10682,N_11522);
nor U14421 (N_14421,N_11373,N_11965);
nor U14422 (N_14422,N_11593,N_10045);
nand U14423 (N_14423,N_10662,N_12156);
xnor U14424 (N_14424,N_10471,N_11353);
xnor U14425 (N_14425,N_11557,N_11849);
nor U14426 (N_14426,N_11051,N_11534);
nor U14427 (N_14427,N_10317,N_12480);
nor U14428 (N_14428,N_11788,N_10999);
nand U14429 (N_14429,N_11704,N_12365);
nor U14430 (N_14430,N_11254,N_10627);
or U14431 (N_14431,N_11608,N_10407);
nand U14432 (N_14432,N_12097,N_10962);
nor U14433 (N_14433,N_10392,N_11923);
nand U14434 (N_14434,N_12196,N_11381);
nand U14435 (N_14435,N_10862,N_10109);
nor U14436 (N_14436,N_10407,N_10322);
nand U14437 (N_14437,N_10074,N_10344);
xnor U14438 (N_14438,N_10696,N_12335);
xor U14439 (N_14439,N_11683,N_12027);
or U14440 (N_14440,N_10248,N_10855);
nand U14441 (N_14441,N_12031,N_10051);
or U14442 (N_14442,N_10438,N_10422);
nor U14443 (N_14443,N_11775,N_12091);
xnor U14444 (N_14444,N_10634,N_11658);
nor U14445 (N_14445,N_10774,N_12046);
or U14446 (N_14446,N_10123,N_11503);
nand U14447 (N_14447,N_11627,N_10927);
xor U14448 (N_14448,N_10183,N_12042);
nand U14449 (N_14449,N_10909,N_12058);
nand U14450 (N_14450,N_11301,N_11327);
or U14451 (N_14451,N_10474,N_11823);
xnor U14452 (N_14452,N_11388,N_11937);
or U14453 (N_14453,N_12322,N_10903);
and U14454 (N_14454,N_11696,N_12443);
xor U14455 (N_14455,N_11307,N_12493);
nand U14456 (N_14456,N_11866,N_11714);
or U14457 (N_14457,N_11774,N_11214);
xor U14458 (N_14458,N_11652,N_10120);
and U14459 (N_14459,N_10276,N_11292);
nand U14460 (N_14460,N_12304,N_11084);
or U14461 (N_14461,N_11948,N_12267);
and U14462 (N_14462,N_10988,N_11987);
xor U14463 (N_14463,N_12157,N_10436);
or U14464 (N_14464,N_11811,N_12296);
nor U14465 (N_14465,N_11742,N_11781);
xor U14466 (N_14466,N_11025,N_10594);
and U14467 (N_14467,N_11797,N_11337);
nor U14468 (N_14468,N_10059,N_11532);
nor U14469 (N_14469,N_11726,N_10349);
or U14470 (N_14470,N_10771,N_11914);
and U14471 (N_14471,N_10775,N_11743);
xnor U14472 (N_14472,N_10638,N_12039);
nand U14473 (N_14473,N_11237,N_10566);
or U14474 (N_14474,N_11165,N_12412);
nor U14475 (N_14475,N_10116,N_10297);
or U14476 (N_14476,N_10241,N_10892);
and U14477 (N_14477,N_12043,N_10309);
and U14478 (N_14478,N_12114,N_11067);
or U14479 (N_14479,N_12477,N_10418);
nand U14480 (N_14480,N_12017,N_11099);
nand U14481 (N_14481,N_10734,N_11960);
and U14482 (N_14482,N_11024,N_10501);
nor U14483 (N_14483,N_10447,N_12051);
xnor U14484 (N_14484,N_12027,N_10199);
nor U14485 (N_14485,N_12129,N_10371);
or U14486 (N_14486,N_10385,N_10438);
nor U14487 (N_14487,N_12031,N_11882);
and U14488 (N_14488,N_11842,N_10234);
or U14489 (N_14489,N_12215,N_11759);
xor U14490 (N_14490,N_11396,N_10218);
nand U14491 (N_14491,N_12000,N_11358);
or U14492 (N_14492,N_10838,N_10606);
nor U14493 (N_14493,N_11385,N_12348);
xor U14494 (N_14494,N_11790,N_11216);
and U14495 (N_14495,N_12086,N_12229);
nor U14496 (N_14496,N_11011,N_10741);
nor U14497 (N_14497,N_10465,N_10809);
nand U14498 (N_14498,N_10186,N_11713);
and U14499 (N_14499,N_10327,N_12346);
nor U14500 (N_14500,N_10675,N_10293);
nand U14501 (N_14501,N_11379,N_12382);
and U14502 (N_14502,N_11646,N_10438);
nor U14503 (N_14503,N_11648,N_11484);
nand U14504 (N_14504,N_11169,N_10827);
xnor U14505 (N_14505,N_10804,N_11231);
nand U14506 (N_14506,N_10823,N_11325);
nand U14507 (N_14507,N_11235,N_11758);
and U14508 (N_14508,N_12174,N_10866);
nor U14509 (N_14509,N_12329,N_11669);
nor U14510 (N_14510,N_11409,N_12442);
or U14511 (N_14511,N_11135,N_10683);
xnor U14512 (N_14512,N_10915,N_11601);
nand U14513 (N_14513,N_11873,N_10220);
or U14514 (N_14514,N_10609,N_12435);
and U14515 (N_14515,N_12005,N_10934);
and U14516 (N_14516,N_10059,N_11047);
xnor U14517 (N_14517,N_10866,N_12413);
nor U14518 (N_14518,N_12261,N_11142);
nor U14519 (N_14519,N_12089,N_10378);
and U14520 (N_14520,N_10161,N_10209);
and U14521 (N_14521,N_12199,N_10067);
or U14522 (N_14522,N_10800,N_11683);
nor U14523 (N_14523,N_12255,N_10228);
nor U14524 (N_14524,N_11863,N_11358);
nand U14525 (N_14525,N_12215,N_12232);
nand U14526 (N_14526,N_12191,N_11260);
nand U14527 (N_14527,N_10173,N_12269);
xnor U14528 (N_14528,N_12312,N_12347);
and U14529 (N_14529,N_12218,N_10438);
or U14530 (N_14530,N_10097,N_11858);
xnor U14531 (N_14531,N_10352,N_11844);
or U14532 (N_14532,N_11987,N_10520);
or U14533 (N_14533,N_10689,N_10822);
nand U14534 (N_14534,N_10286,N_12255);
nand U14535 (N_14535,N_12044,N_10059);
or U14536 (N_14536,N_12302,N_10198);
and U14537 (N_14537,N_11263,N_10280);
nand U14538 (N_14538,N_10919,N_10243);
nand U14539 (N_14539,N_10882,N_10092);
xor U14540 (N_14540,N_12292,N_11134);
nor U14541 (N_14541,N_11430,N_12243);
nor U14542 (N_14542,N_12457,N_10333);
and U14543 (N_14543,N_10331,N_11310);
and U14544 (N_14544,N_11133,N_10328);
xor U14545 (N_14545,N_12488,N_10965);
nand U14546 (N_14546,N_12160,N_10346);
xnor U14547 (N_14547,N_11850,N_12041);
nor U14548 (N_14548,N_10794,N_10197);
xnor U14549 (N_14549,N_10559,N_10881);
xor U14550 (N_14550,N_12462,N_11474);
xor U14551 (N_14551,N_10904,N_12228);
and U14552 (N_14552,N_10736,N_12495);
or U14553 (N_14553,N_12472,N_12413);
nand U14554 (N_14554,N_11172,N_12200);
nor U14555 (N_14555,N_11831,N_11547);
xnor U14556 (N_14556,N_11247,N_11577);
and U14557 (N_14557,N_12012,N_11923);
nand U14558 (N_14558,N_12362,N_10020);
nand U14559 (N_14559,N_11475,N_10560);
nor U14560 (N_14560,N_11444,N_12176);
or U14561 (N_14561,N_10506,N_11697);
nand U14562 (N_14562,N_11514,N_10776);
or U14563 (N_14563,N_11616,N_11568);
xnor U14564 (N_14564,N_10279,N_10152);
nor U14565 (N_14565,N_11355,N_11816);
xnor U14566 (N_14566,N_10671,N_11263);
or U14567 (N_14567,N_10183,N_12345);
and U14568 (N_14568,N_10513,N_10158);
or U14569 (N_14569,N_11674,N_11791);
nor U14570 (N_14570,N_10607,N_12041);
and U14571 (N_14571,N_12023,N_11605);
nand U14572 (N_14572,N_12332,N_11408);
and U14573 (N_14573,N_12105,N_12002);
nor U14574 (N_14574,N_10563,N_11748);
or U14575 (N_14575,N_10637,N_11072);
or U14576 (N_14576,N_10226,N_11812);
nand U14577 (N_14577,N_11531,N_11320);
xnor U14578 (N_14578,N_12471,N_10180);
nand U14579 (N_14579,N_10997,N_10372);
nor U14580 (N_14580,N_11207,N_10584);
or U14581 (N_14581,N_10364,N_11022);
and U14582 (N_14582,N_12013,N_10082);
nor U14583 (N_14583,N_11727,N_11448);
and U14584 (N_14584,N_11010,N_10397);
xnor U14585 (N_14585,N_10254,N_10672);
nor U14586 (N_14586,N_12325,N_11571);
nor U14587 (N_14587,N_11804,N_11467);
or U14588 (N_14588,N_11863,N_11872);
nor U14589 (N_14589,N_11756,N_10942);
xor U14590 (N_14590,N_12370,N_10963);
xor U14591 (N_14591,N_10830,N_10581);
or U14592 (N_14592,N_10225,N_11889);
nand U14593 (N_14593,N_10846,N_12238);
xnor U14594 (N_14594,N_10447,N_11862);
or U14595 (N_14595,N_10633,N_11295);
and U14596 (N_14596,N_10019,N_11795);
nor U14597 (N_14597,N_11011,N_12059);
nand U14598 (N_14598,N_10175,N_11817);
nand U14599 (N_14599,N_10952,N_12353);
nand U14600 (N_14600,N_11323,N_12019);
nand U14601 (N_14601,N_10007,N_10849);
and U14602 (N_14602,N_12431,N_12168);
or U14603 (N_14603,N_11311,N_11318);
nand U14604 (N_14604,N_12304,N_12294);
xnor U14605 (N_14605,N_11849,N_10408);
and U14606 (N_14606,N_12102,N_10868);
xor U14607 (N_14607,N_10123,N_10198);
and U14608 (N_14608,N_10075,N_10408);
nor U14609 (N_14609,N_11792,N_10301);
or U14610 (N_14610,N_12376,N_10300);
xnor U14611 (N_14611,N_11430,N_12258);
nand U14612 (N_14612,N_11055,N_12132);
or U14613 (N_14613,N_10996,N_10010);
and U14614 (N_14614,N_10433,N_11166);
xor U14615 (N_14615,N_12175,N_12494);
or U14616 (N_14616,N_12316,N_10558);
nand U14617 (N_14617,N_10653,N_10612);
xnor U14618 (N_14618,N_12190,N_12098);
nor U14619 (N_14619,N_12106,N_10929);
or U14620 (N_14620,N_10956,N_12193);
nor U14621 (N_14621,N_11978,N_11981);
nand U14622 (N_14622,N_11231,N_10728);
nand U14623 (N_14623,N_11259,N_12328);
and U14624 (N_14624,N_12216,N_10407);
nand U14625 (N_14625,N_10088,N_11508);
or U14626 (N_14626,N_10218,N_12191);
xnor U14627 (N_14627,N_11391,N_10907);
nor U14628 (N_14628,N_10265,N_10236);
and U14629 (N_14629,N_12231,N_11355);
or U14630 (N_14630,N_11572,N_11411);
nand U14631 (N_14631,N_11596,N_11390);
xnor U14632 (N_14632,N_12352,N_11325);
xor U14633 (N_14633,N_10009,N_11892);
nand U14634 (N_14634,N_11786,N_10930);
and U14635 (N_14635,N_10153,N_12386);
nand U14636 (N_14636,N_11360,N_11163);
xor U14637 (N_14637,N_10992,N_11429);
xnor U14638 (N_14638,N_11470,N_10143);
or U14639 (N_14639,N_12456,N_10475);
nor U14640 (N_14640,N_10598,N_12322);
nand U14641 (N_14641,N_12090,N_11740);
or U14642 (N_14642,N_11973,N_11263);
xnor U14643 (N_14643,N_10309,N_10572);
xnor U14644 (N_14644,N_11282,N_11450);
or U14645 (N_14645,N_12222,N_11864);
nor U14646 (N_14646,N_12239,N_11136);
xnor U14647 (N_14647,N_11725,N_11632);
nand U14648 (N_14648,N_10393,N_12362);
xnor U14649 (N_14649,N_11358,N_11634);
nor U14650 (N_14650,N_12333,N_12155);
and U14651 (N_14651,N_12042,N_11723);
nand U14652 (N_14652,N_12013,N_11975);
and U14653 (N_14653,N_11505,N_12311);
nor U14654 (N_14654,N_11708,N_11005);
nand U14655 (N_14655,N_10452,N_12053);
and U14656 (N_14656,N_11402,N_11888);
and U14657 (N_14657,N_10289,N_10014);
or U14658 (N_14658,N_10687,N_11795);
nor U14659 (N_14659,N_10892,N_11743);
nor U14660 (N_14660,N_10798,N_10439);
and U14661 (N_14661,N_10720,N_11320);
and U14662 (N_14662,N_10703,N_11606);
xor U14663 (N_14663,N_10675,N_11318);
nor U14664 (N_14664,N_11587,N_10256);
or U14665 (N_14665,N_10583,N_11692);
or U14666 (N_14666,N_10465,N_11151);
xnor U14667 (N_14667,N_10269,N_11317);
nor U14668 (N_14668,N_11750,N_10800);
nor U14669 (N_14669,N_10791,N_12083);
xnor U14670 (N_14670,N_10442,N_10776);
or U14671 (N_14671,N_11239,N_11982);
nor U14672 (N_14672,N_10590,N_10327);
or U14673 (N_14673,N_11210,N_10317);
nand U14674 (N_14674,N_11348,N_10158);
or U14675 (N_14675,N_10470,N_10559);
and U14676 (N_14676,N_10407,N_11007);
xor U14677 (N_14677,N_10913,N_11530);
nand U14678 (N_14678,N_10953,N_10964);
nand U14679 (N_14679,N_11443,N_10596);
xnor U14680 (N_14680,N_11332,N_10938);
xor U14681 (N_14681,N_11206,N_12421);
nor U14682 (N_14682,N_11503,N_11770);
nand U14683 (N_14683,N_10740,N_11592);
nor U14684 (N_14684,N_10375,N_10900);
nor U14685 (N_14685,N_11220,N_10435);
or U14686 (N_14686,N_12441,N_11126);
nand U14687 (N_14687,N_10204,N_11034);
or U14688 (N_14688,N_11893,N_12241);
or U14689 (N_14689,N_12461,N_10409);
and U14690 (N_14690,N_11089,N_11358);
and U14691 (N_14691,N_10747,N_12193);
nor U14692 (N_14692,N_11261,N_12212);
and U14693 (N_14693,N_11417,N_12341);
and U14694 (N_14694,N_11656,N_10047);
and U14695 (N_14695,N_11241,N_10268);
nand U14696 (N_14696,N_11734,N_11440);
or U14697 (N_14697,N_12191,N_12257);
and U14698 (N_14698,N_10799,N_12493);
xor U14699 (N_14699,N_11643,N_10291);
or U14700 (N_14700,N_12117,N_11591);
xnor U14701 (N_14701,N_10548,N_11694);
xor U14702 (N_14702,N_10654,N_11618);
nor U14703 (N_14703,N_11237,N_11798);
xnor U14704 (N_14704,N_12085,N_10161);
xnor U14705 (N_14705,N_11028,N_11935);
xor U14706 (N_14706,N_11014,N_11975);
xnor U14707 (N_14707,N_11569,N_10106);
nand U14708 (N_14708,N_12341,N_11590);
nand U14709 (N_14709,N_10547,N_12107);
nor U14710 (N_14710,N_11180,N_10666);
nand U14711 (N_14711,N_12182,N_11045);
nor U14712 (N_14712,N_12402,N_12119);
xor U14713 (N_14713,N_10449,N_12053);
nand U14714 (N_14714,N_12167,N_11855);
nor U14715 (N_14715,N_11445,N_12254);
nand U14716 (N_14716,N_11279,N_10755);
nand U14717 (N_14717,N_11899,N_11290);
and U14718 (N_14718,N_12140,N_11129);
xor U14719 (N_14719,N_11149,N_11250);
xnor U14720 (N_14720,N_11380,N_10609);
nor U14721 (N_14721,N_10791,N_10079);
nand U14722 (N_14722,N_10064,N_11851);
nor U14723 (N_14723,N_11574,N_10515);
nor U14724 (N_14724,N_10220,N_11982);
or U14725 (N_14725,N_11804,N_10120);
nand U14726 (N_14726,N_10875,N_10569);
or U14727 (N_14727,N_12241,N_11642);
nand U14728 (N_14728,N_10255,N_11325);
or U14729 (N_14729,N_11876,N_11705);
and U14730 (N_14730,N_11346,N_12296);
and U14731 (N_14731,N_11329,N_12499);
or U14732 (N_14732,N_11549,N_10378);
nand U14733 (N_14733,N_11472,N_11202);
nand U14734 (N_14734,N_10234,N_11538);
nor U14735 (N_14735,N_12281,N_10661);
nor U14736 (N_14736,N_12217,N_11258);
nand U14737 (N_14737,N_11586,N_10299);
or U14738 (N_14738,N_11872,N_10122);
xnor U14739 (N_14739,N_11140,N_12437);
nand U14740 (N_14740,N_10642,N_11657);
xor U14741 (N_14741,N_10725,N_12470);
nor U14742 (N_14742,N_12361,N_12155);
xnor U14743 (N_14743,N_11355,N_11800);
and U14744 (N_14744,N_11678,N_10865);
nor U14745 (N_14745,N_10717,N_11978);
nand U14746 (N_14746,N_12033,N_11937);
or U14747 (N_14747,N_10109,N_12429);
nor U14748 (N_14748,N_12041,N_10551);
nor U14749 (N_14749,N_10109,N_12159);
or U14750 (N_14750,N_11530,N_10116);
nand U14751 (N_14751,N_11921,N_11694);
or U14752 (N_14752,N_11783,N_11256);
xor U14753 (N_14753,N_10249,N_10236);
and U14754 (N_14754,N_10394,N_10083);
xnor U14755 (N_14755,N_11472,N_12334);
nand U14756 (N_14756,N_10589,N_12251);
and U14757 (N_14757,N_10291,N_11928);
nand U14758 (N_14758,N_11030,N_12013);
nand U14759 (N_14759,N_11561,N_11741);
and U14760 (N_14760,N_11425,N_10544);
nand U14761 (N_14761,N_10093,N_12215);
nor U14762 (N_14762,N_12140,N_12214);
xor U14763 (N_14763,N_10782,N_11244);
nand U14764 (N_14764,N_11314,N_11217);
or U14765 (N_14765,N_12483,N_10556);
nor U14766 (N_14766,N_12413,N_12054);
or U14767 (N_14767,N_11015,N_11167);
nor U14768 (N_14768,N_10769,N_11889);
and U14769 (N_14769,N_10925,N_10616);
nand U14770 (N_14770,N_12073,N_10149);
xnor U14771 (N_14771,N_11010,N_10339);
nor U14772 (N_14772,N_10812,N_11861);
and U14773 (N_14773,N_12205,N_10464);
or U14774 (N_14774,N_11811,N_11604);
nor U14775 (N_14775,N_11333,N_10390);
xor U14776 (N_14776,N_11726,N_12470);
and U14777 (N_14777,N_10252,N_11536);
nor U14778 (N_14778,N_11013,N_11238);
nand U14779 (N_14779,N_11402,N_12014);
nand U14780 (N_14780,N_10212,N_11151);
nor U14781 (N_14781,N_11579,N_12021);
xnor U14782 (N_14782,N_10745,N_10690);
nand U14783 (N_14783,N_11758,N_12241);
and U14784 (N_14784,N_11575,N_10489);
and U14785 (N_14785,N_11611,N_10638);
nor U14786 (N_14786,N_11988,N_10382);
xnor U14787 (N_14787,N_10624,N_11782);
or U14788 (N_14788,N_10976,N_11056);
and U14789 (N_14789,N_11637,N_11106);
xor U14790 (N_14790,N_11078,N_11160);
nor U14791 (N_14791,N_11894,N_10285);
or U14792 (N_14792,N_11184,N_10075);
or U14793 (N_14793,N_11083,N_11727);
nor U14794 (N_14794,N_11900,N_11280);
or U14795 (N_14795,N_11722,N_10485);
nand U14796 (N_14796,N_10300,N_11331);
or U14797 (N_14797,N_10871,N_11717);
and U14798 (N_14798,N_10565,N_11910);
or U14799 (N_14799,N_11788,N_10433);
nor U14800 (N_14800,N_10274,N_10182);
or U14801 (N_14801,N_10083,N_11238);
nor U14802 (N_14802,N_12104,N_11105);
or U14803 (N_14803,N_10741,N_10897);
or U14804 (N_14804,N_10347,N_11341);
xor U14805 (N_14805,N_10648,N_11117);
xnor U14806 (N_14806,N_10581,N_10082);
and U14807 (N_14807,N_11653,N_10083);
and U14808 (N_14808,N_12250,N_11844);
and U14809 (N_14809,N_11343,N_11346);
nand U14810 (N_14810,N_10770,N_10813);
xor U14811 (N_14811,N_10581,N_12206);
nand U14812 (N_14812,N_10828,N_11160);
nor U14813 (N_14813,N_10424,N_11962);
nand U14814 (N_14814,N_12153,N_11075);
and U14815 (N_14815,N_11315,N_11113);
nor U14816 (N_14816,N_12187,N_10238);
or U14817 (N_14817,N_12070,N_10774);
xor U14818 (N_14818,N_11100,N_10453);
nor U14819 (N_14819,N_11961,N_10968);
or U14820 (N_14820,N_11711,N_10291);
or U14821 (N_14821,N_11040,N_11341);
and U14822 (N_14822,N_11699,N_11510);
nor U14823 (N_14823,N_12469,N_11044);
or U14824 (N_14824,N_10921,N_12150);
and U14825 (N_14825,N_12378,N_12463);
xor U14826 (N_14826,N_11648,N_10299);
and U14827 (N_14827,N_10490,N_12289);
or U14828 (N_14828,N_11149,N_11154);
or U14829 (N_14829,N_10145,N_11591);
or U14830 (N_14830,N_11120,N_11871);
and U14831 (N_14831,N_10835,N_10914);
and U14832 (N_14832,N_11327,N_10199);
xor U14833 (N_14833,N_11166,N_12247);
and U14834 (N_14834,N_12146,N_12426);
or U14835 (N_14835,N_10047,N_10048);
or U14836 (N_14836,N_12062,N_10849);
and U14837 (N_14837,N_12112,N_10554);
xnor U14838 (N_14838,N_10748,N_11445);
and U14839 (N_14839,N_11877,N_11795);
nor U14840 (N_14840,N_11670,N_12468);
or U14841 (N_14841,N_12179,N_11950);
nand U14842 (N_14842,N_11179,N_12259);
or U14843 (N_14843,N_10861,N_10507);
nand U14844 (N_14844,N_11046,N_10638);
or U14845 (N_14845,N_10120,N_11704);
xnor U14846 (N_14846,N_10166,N_10904);
or U14847 (N_14847,N_10962,N_10936);
nand U14848 (N_14848,N_10945,N_12142);
and U14849 (N_14849,N_10245,N_12075);
nand U14850 (N_14850,N_10309,N_10557);
or U14851 (N_14851,N_11710,N_10368);
or U14852 (N_14852,N_11506,N_11395);
xor U14853 (N_14853,N_11437,N_10654);
and U14854 (N_14854,N_12303,N_11568);
nor U14855 (N_14855,N_10385,N_11951);
xor U14856 (N_14856,N_12419,N_11075);
nor U14857 (N_14857,N_11571,N_12347);
or U14858 (N_14858,N_10720,N_12110);
xor U14859 (N_14859,N_11098,N_11748);
nand U14860 (N_14860,N_11668,N_11077);
and U14861 (N_14861,N_11233,N_11543);
xor U14862 (N_14862,N_11898,N_11431);
or U14863 (N_14863,N_10709,N_10691);
or U14864 (N_14864,N_10978,N_11323);
and U14865 (N_14865,N_11978,N_12097);
nand U14866 (N_14866,N_10031,N_11701);
nor U14867 (N_14867,N_12488,N_12049);
and U14868 (N_14868,N_10580,N_10637);
nor U14869 (N_14869,N_10864,N_10985);
or U14870 (N_14870,N_10270,N_11211);
nand U14871 (N_14871,N_11450,N_10027);
or U14872 (N_14872,N_10091,N_10039);
xor U14873 (N_14873,N_11135,N_10273);
nand U14874 (N_14874,N_10807,N_10576);
xor U14875 (N_14875,N_12365,N_11269);
or U14876 (N_14876,N_10115,N_10231);
nor U14877 (N_14877,N_11556,N_11624);
or U14878 (N_14878,N_10768,N_10430);
xnor U14879 (N_14879,N_10945,N_10670);
xnor U14880 (N_14880,N_12257,N_11634);
nand U14881 (N_14881,N_12207,N_12219);
and U14882 (N_14882,N_10358,N_10236);
or U14883 (N_14883,N_12400,N_10525);
nand U14884 (N_14884,N_11041,N_11881);
nand U14885 (N_14885,N_12483,N_12382);
or U14886 (N_14886,N_12385,N_11716);
xor U14887 (N_14887,N_11435,N_11808);
xnor U14888 (N_14888,N_10844,N_11454);
nor U14889 (N_14889,N_11740,N_12204);
and U14890 (N_14890,N_10205,N_10694);
and U14891 (N_14891,N_12366,N_11003);
nor U14892 (N_14892,N_10619,N_11649);
and U14893 (N_14893,N_11091,N_10289);
xor U14894 (N_14894,N_11234,N_10727);
and U14895 (N_14895,N_11534,N_10814);
and U14896 (N_14896,N_11248,N_10661);
nor U14897 (N_14897,N_10925,N_11213);
nor U14898 (N_14898,N_11100,N_10778);
nor U14899 (N_14899,N_11037,N_11074);
nand U14900 (N_14900,N_12082,N_11834);
and U14901 (N_14901,N_12424,N_10511);
or U14902 (N_14902,N_12419,N_10805);
or U14903 (N_14903,N_11509,N_11177);
xnor U14904 (N_14904,N_11568,N_12474);
nand U14905 (N_14905,N_10762,N_10310);
xor U14906 (N_14906,N_10651,N_12224);
nand U14907 (N_14907,N_11982,N_11856);
nand U14908 (N_14908,N_10418,N_11646);
and U14909 (N_14909,N_12430,N_10441);
and U14910 (N_14910,N_10606,N_10104);
or U14911 (N_14911,N_10740,N_12048);
nand U14912 (N_14912,N_11839,N_11589);
nor U14913 (N_14913,N_11942,N_12389);
or U14914 (N_14914,N_11300,N_10133);
and U14915 (N_14915,N_12269,N_10527);
or U14916 (N_14916,N_10543,N_11665);
nand U14917 (N_14917,N_11269,N_11750);
xor U14918 (N_14918,N_10873,N_10623);
and U14919 (N_14919,N_11263,N_10683);
nor U14920 (N_14920,N_11071,N_12339);
xnor U14921 (N_14921,N_11980,N_11082);
nor U14922 (N_14922,N_11106,N_11981);
xnor U14923 (N_14923,N_10469,N_10938);
nand U14924 (N_14924,N_11104,N_11522);
nand U14925 (N_14925,N_11497,N_11009);
or U14926 (N_14926,N_12455,N_11342);
nor U14927 (N_14927,N_12224,N_10466);
nand U14928 (N_14928,N_10374,N_11831);
nand U14929 (N_14929,N_11916,N_12167);
nand U14930 (N_14930,N_11468,N_10671);
and U14931 (N_14931,N_11466,N_11124);
or U14932 (N_14932,N_11761,N_10765);
nand U14933 (N_14933,N_11820,N_11779);
nor U14934 (N_14934,N_11221,N_10486);
xnor U14935 (N_14935,N_11362,N_10860);
xnor U14936 (N_14936,N_12111,N_11152);
xor U14937 (N_14937,N_10571,N_10298);
nand U14938 (N_14938,N_11383,N_11669);
or U14939 (N_14939,N_10273,N_11499);
nand U14940 (N_14940,N_12096,N_12088);
and U14941 (N_14941,N_11901,N_12266);
nor U14942 (N_14942,N_12220,N_10370);
or U14943 (N_14943,N_11842,N_11797);
and U14944 (N_14944,N_11221,N_10581);
or U14945 (N_14945,N_10134,N_10423);
or U14946 (N_14946,N_11600,N_10082);
xor U14947 (N_14947,N_11481,N_11802);
and U14948 (N_14948,N_11313,N_11540);
xor U14949 (N_14949,N_10989,N_11097);
or U14950 (N_14950,N_10695,N_10173);
nor U14951 (N_14951,N_11743,N_10582);
or U14952 (N_14952,N_10018,N_10178);
or U14953 (N_14953,N_10739,N_10480);
nand U14954 (N_14954,N_11777,N_11226);
and U14955 (N_14955,N_10305,N_12433);
nand U14956 (N_14956,N_11345,N_10773);
nand U14957 (N_14957,N_10143,N_11593);
nor U14958 (N_14958,N_10832,N_12297);
or U14959 (N_14959,N_11935,N_11753);
nand U14960 (N_14960,N_10538,N_11660);
and U14961 (N_14961,N_12040,N_12327);
or U14962 (N_14962,N_10923,N_11149);
nor U14963 (N_14963,N_12035,N_11331);
nand U14964 (N_14964,N_12194,N_10680);
and U14965 (N_14965,N_11062,N_10855);
and U14966 (N_14966,N_10537,N_10186);
nand U14967 (N_14967,N_10296,N_10810);
or U14968 (N_14968,N_10244,N_11972);
nand U14969 (N_14969,N_11410,N_10444);
or U14970 (N_14970,N_11842,N_10576);
nor U14971 (N_14971,N_11001,N_11531);
and U14972 (N_14972,N_10088,N_10588);
or U14973 (N_14973,N_10474,N_11549);
or U14974 (N_14974,N_10049,N_11833);
nor U14975 (N_14975,N_10507,N_10323);
nor U14976 (N_14976,N_10368,N_10438);
or U14977 (N_14977,N_11232,N_12086);
or U14978 (N_14978,N_11273,N_10897);
nor U14979 (N_14979,N_12351,N_10956);
xnor U14980 (N_14980,N_11518,N_10430);
or U14981 (N_14981,N_10421,N_11318);
nor U14982 (N_14982,N_10513,N_11525);
nand U14983 (N_14983,N_11815,N_10410);
nand U14984 (N_14984,N_12081,N_10517);
nand U14985 (N_14985,N_11885,N_10361);
and U14986 (N_14986,N_10392,N_10588);
nor U14987 (N_14987,N_10971,N_11290);
or U14988 (N_14988,N_11459,N_11006);
xnor U14989 (N_14989,N_10341,N_10908);
nor U14990 (N_14990,N_11172,N_10245);
xnor U14991 (N_14991,N_12074,N_10970);
xor U14992 (N_14992,N_10010,N_10651);
nor U14993 (N_14993,N_10405,N_11857);
nand U14994 (N_14994,N_11602,N_10825);
xnor U14995 (N_14995,N_12117,N_12300);
xor U14996 (N_14996,N_11970,N_10753);
and U14997 (N_14997,N_10540,N_10863);
nor U14998 (N_14998,N_12301,N_10157);
nand U14999 (N_14999,N_12475,N_10513);
nor U15000 (N_15000,N_13125,N_12763);
nand U15001 (N_15001,N_14383,N_13187);
nand U15002 (N_15002,N_12613,N_14849);
nor U15003 (N_15003,N_13114,N_12894);
or U15004 (N_15004,N_13315,N_13810);
nor U15005 (N_15005,N_13213,N_14059);
xor U15006 (N_15006,N_14810,N_14174);
and U15007 (N_15007,N_13185,N_13794);
xor U15008 (N_15008,N_14424,N_14209);
or U15009 (N_15009,N_14392,N_14558);
and U15010 (N_15010,N_13874,N_14274);
or U15011 (N_15011,N_13010,N_14702);
and U15012 (N_15012,N_13283,N_14560);
or U15013 (N_15013,N_14811,N_14917);
nand U15014 (N_15014,N_13799,N_13851);
xnor U15015 (N_15015,N_14304,N_13872);
and U15016 (N_15016,N_13764,N_13102);
and U15017 (N_15017,N_14318,N_12594);
xnor U15018 (N_15018,N_12671,N_13113);
or U15019 (N_15019,N_12754,N_14454);
nor U15020 (N_15020,N_12903,N_13277);
nor U15021 (N_15021,N_14226,N_13757);
nor U15022 (N_15022,N_12838,N_13622);
nand U15023 (N_15023,N_13739,N_14524);
xnor U15024 (N_15024,N_13494,N_12726);
xnor U15025 (N_15025,N_12652,N_13716);
or U15026 (N_15026,N_14580,N_13720);
xor U15027 (N_15027,N_14007,N_14643);
and U15028 (N_15028,N_12541,N_12574);
nand U15029 (N_15029,N_14427,N_12720);
nor U15030 (N_15030,N_14111,N_13147);
or U15031 (N_15031,N_13328,N_14404);
or U15032 (N_15032,N_14141,N_12665);
xor U15033 (N_15033,N_14614,N_14017);
nand U15034 (N_15034,N_14447,N_13983);
xnor U15035 (N_15035,N_13308,N_12576);
nor U15036 (N_15036,N_12623,N_12622);
nand U15037 (N_15037,N_14449,N_13921);
and U15038 (N_15038,N_12690,N_14704);
or U15039 (N_15039,N_14587,N_13355);
xor U15040 (N_15040,N_13914,N_14589);
xor U15041 (N_15041,N_12591,N_14605);
or U15042 (N_15042,N_14024,N_14649);
xor U15043 (N_15043,N_12633,N_14296);
xor U15044 (N_15044,N_12802,N_14433);
or U15045 (N_15045,N_13659,N_12519);
nor U15046 (N_15046,N_14489,N_14106);
or U15047 (N_15047,N_14933,N_12571);
or U15048 (N_15048,N_12952,N_12626);
or U15049 (N_15049,N_13203,N_12874);
nand U15050 (N_15050,N_13364,N_14420);
and U15051 (N_15051,N_13427,N_12771);
nand U15052 (N_15052,N_13870,N_14464);
and U15053 (N_15053,N_13955,N_13060);
xor U15054 (N_15054,N_13404,N_12785);
nand U15055 (N_15055,N_12801,N_13719);
and U15056 (N_15056,N_13141,N_14157);
and U15057 (N_15057,N_12592,N_14981);
and U15058 (N_15058,N_13941,N_14134);
nand U15059 (N_15059,N_12538,N_14081);
nand U15060 (N_15060,N_13423,N_13030);
nand U15061 (N_15061,N_14579,N_14323);
nor U15062 (N_15062,N_13433,N_14232);
nand U15063 (N_15063,N_13497,N_14572);
xnor U15064 (N_15064,N_12523,N_13304);
nor U15065 (N_15065,N_12542,N_14343);
and U15066 (N_15066,N_12799,N_13119);
or U15067 (N_15067,N_13037,N_13812);
nor U15068 (N_15068,N_14995,N_14241);
xor U15069 (N_15069,N_14066,N_14993);
and U15070 (N_15070,N_13070,N_13844);
nor U15071 (N_15071,N_13432,N_12647);
nand U15072 (N_15072,N_12746,N_14475);
nand U15073 (N_15073,N_12853,N_14728);
and U15074 (N_15074,N_12867,N_13396);
nand U15075 (N_15075,N_14508,N_12779);
and U15076 (N_15076,N_13149,N_12937);
and U15077 (N_15077,N_13986,N_14992);
nand U15078 (N_15078,N_12527,N_14294);
nor U15079 (N_15079,N_14611,N_14990);
xor U15080 (N_15080,N_13057,N_13649);
and U15081 (N_15081,N_13855,N_13292);
and U15082 (N_15082,N_14921,N_13152);
xor U15083 (N_15083,N_14836,N_14909);
or U15084 (N_15084,N_12605,N_13223);
nand U15085 (N_15085,N_13353,N_14506);
nor U15086 (N_15086,N_12843,N_13498);
xnor U15087 (N_15087,N_13643,N_12960);
and U15088 (N_15088,N_13572,N_13031);
nand U15089 (N_15089,N_14786,N_13603);
and U15090 (N_15090,N_13545,N_14263);
and U15091 (N_15091,N_13687,N_14575);
nand U15092 (N_15092,N_13845,N_14636);
or U15093 (N_15093,N_13880,N_13461);
and U15094 (N_15094,N_12927,N_13318);
xor U15095 (N_15095,N_13202,N_14253);
nor U15096 (N_15096,N_12641,N_13631);
and U15097 (N_15097,N_14503,N_14275);
xor U15098 (N_15098,N_14431,N_14395);
nor U15099 (N_15099,N_14281,N_14391);
or U15100 (N_15100,N_13701,N_14255);
xor U15101 (N_15101,N_12819,N_12938);
nand U15102 (N_15102,N_12756,N_13281);
xor U15103 (N_15103,N_14735,N_12558);
and U15104 (N_15104,N_13744,N_12737);
and U15105 (N_15105,N_13510,N_14718);
and U15106 (N_15106,N_14051,N_13549);
or U15107 (N_15107,N_12856,N_12944);
or U15108 (N_15108,N_14827,N_13121);
nor U15109 (N_15109,N_13592,N_13373);
or U15110 (N_15110,N_12738,N_14135);
or U15111 (N_15111,N_13873,N_13877);
or U15112 (N_15112,N_14912,N_14320);
and U15113 (N_15113,N_14600,N_14003);
nor U15114 (N_15114,N_12818,N_14831);
or U15115 (N_15115,N_13201,N_13234);
or U15116 (N_15116,N_13309,N_14989);
and U15117 (N_15117,N_14128,N_12981);
and U15118 (N_15118,N_13481,N_14271);
and U15119 (N_15119,N_13783,N_14915);
or U15120 (N_15120,N_13733,N_13050);
nor U15121 (N_15121,N_13382,N_14940);
xor U15122 (N_15122,N_13492,N_14664);
and U15123 (N_15123,N_13018,N_13412);
nor U15124 (N_15124,N_14257,N_13204);
xnor U15125 (N_15125,N_12932,N_14821);
nand U15126 (N_15126,N_12503,N_14741);
or U15127 (N_15127,N_12520,N_14440);
and U15128 (N_15128,N_12986,N_12793);
xor U15129 (N_15129,N_14476,N_12947);
and U15130 (N_15130,N_13178,N_13192);
and U15131 (N_15131,N_13157,N_14259);
nand U15132 (N_15132,N_13953,N_13507);
xnor U15133 (N_15133,N_14100,N_12828);
nand U15134 (N_15134,N_14149,N_13245);
or U15135 (N_15135,N_12621,N_14366);
nor U15136 (N_15136,N_14617,N_14722);
nor U15137 (N_15137,N_14077,N_14799);
nand U15138 (N_15138,N_14947,N_13418);
or U15139 (N_15139,N_13891,N_13957);
xor U15140 (N_15140,N_12524,N_12717);
nand U15141 (N_15141,N_12729,N_13605);
nor U15142 (N_15142,N_12922,N_13906);
or U15143 (N_15143,N_13322,N_13860);
nor U15144 (N_15144,N_12718,N_14672);
xor U15145 (N_15145,N_14734,N_13271);
and U15146 (N_15146,N_12862,N_13841);
nand U15147 (N_15147,N_14897,N_12996);
or U15148 (N_15148,N_14914,N_12943);
nor U15149 (N_15149,N_14711,N_14759);
xor U15150 (N_15150,N_14610,N_12772);
and U15151 (N_15151,N_14820,N_14481);
xnor U15152 (N_15152,N_14109,N_13680);
nor U15153 (N_15153,N_13750,N_14886);
nor U15154 (N_15154,N_14783,N_12757);
nor U15155 (N_15155,N_13616,N_12615);
xnor U15156 (N_15156,N_13473,N_14154);
xnor U15157 (N_15157,N_14049,N_13391);
or U15158 (N_15158,N_13881,N_12821);
and U15159 (N_15159,N_13039,N_13337);
and U15160 (N_15160,N_12871,N_13021);
nand U15161 (N_15161,N_13267,N_13142);
nand U15162 (N_15162,N_13761,N_12666);
xor U15163 (N_15163,N_12941,N_14311);
and U15164 (N_15164,N_13032,N_13711);
nor U15165 (N_15165,N_14014,N_12566);
nand U15166 (N_15166,N_12685,N_12739);
or U15167 (N_15167,N_14858,N_14022);
or U15168 (N_15168,N_13968,N_14844);
xnor U15169 (N_15169,N_13013,N_12640);
xor U15170 (N_15170,N_14678,N_14548);
nor U15171 (N_15171,N_12815,N_13746);
nand U15172 (N_15172,N_14772,N_12733);
and U15173 (N_15173,N_13671,N_13995);
nand U15174 (N_15174,N_12829,N_13782);
or U15175 (N_15175,N_12533,N_13883);
nand U15176 (N_15176,N_12510,N_13969);
or U15177 (N_15177,N_14179,N_13313);
or U15178 (N_15178,N_13814,N_14574);
xnor U15179 (N_15179,N_12724,N_13697);
or U15180 (N_15180,N_13707,N_13573);
and U15181 (N_15181,N_14302,N_13601);
nand U15182 (N_15182,N_12910,N_14126);
nor U15183 (N_15183,N_13096,N_13205);
nand U15184 (N_15184,N_13491,N_13749);
and U15185 (N_15185,N_14339,N_13227);
or U15186 (N_15186,N_13862,N_14593);
nand U15187 (N_15187,N_13100,N_13407);
and U15188 (N_15188,N_13604,N_13439);
or U15189 (N_15189,N_14554,N_12681);
nor U15190 (N_15190,N_13048,N_13496);
nor U15191 (N_15191,N_14763,N_13665);
or U15192 (N_15192,N_13903,N_14334);
or U15193 (N_15193,N_12808,N_13256);
or U15194 (N_15194,N_12939,N_12777);
and U15195 (N_15195,N_13935,N_14971);
or U15196 (N_15196,N_14522,N_12830);
and U15197 (N_15197,N_14514,N_14078);
xnor U15198 (N_15198,N_13965,N_13093);
or U15199 (N_15199,N_12512,N_14237);
xnor U15200 (N_15200,N_13135,N_13893);
and U15201 (N_15201,N_14752,N_13884);
and U15202 (N_15202,N_13811,N_14069);
nand U15203 (N_15203,N_13335,N_14616);
and U15204 (N_15204,N_14796,N_13779);
and U15205 (N_15205,N_13158,N_13217);
and U15206 (N_15206,N_13194,N_14098);
and U15207 (N_15207,N_13791,N_12762);
nor U15208 (N_15208,N_13774,N_13876);
xor U15209 (N_15209,N_12766,N_12860);
and U15210 (N_15210,N_14520,N_14452);
and U15211 (N_15211,N_14129,N_14932);
or U15212 (N_15212,N_12865,N_13395);
nand U15213 (N_15213,N_13105,N_12839);
and U15214 (N_15214,N_13648,N_12926);
or U15215 (N_15215,N_12847,N_13082);
nor U15216 (N_15216,N_13366,N_14155);
and U15217 (N_15217,N_14876,N_14270);
and U15218 (N_15218,N_14695,N_14056);
xnor U15219 (N_15219,N_14723,N_12611);
xor U15220 (N_15220,N_12677,N_13793);
nor U15221 (N_15221,N_14467,N_12700);
nand U15222 (N_15222,N_12961,N_14252);
nand U15223 (N_15223,N_14784,N_14743);
xnor U15224 (N_15224,N_14519,N_14905);
or U15225 (N_15225,N_14544,N_12689);
and U15226 (N_15226,N_14653,N_14386);
xor U15227 (N_15227,N_13111,N_13897);
nand U15228 (N_15228,N_13686,N_13555);
nand U15229 (N_15229,N_14691,N_13288);
xor U15230 (N_15230,N_13773,N_12883);
xor U15231 (N_15231,N_14895,N_13843);
or U15232 (N_15232,N_13300,N_13700);
nand U15233 (N_15233,N_14585,N_13011);
xnor U15234 (N_15234,N_14987,N_13343);
or U15235 (N_15235,N_13087,N_13517);
and U15236 (N_15236,N_13869,N_13836);
and U15237 (N_15237,N_14652,N_12565);
and U15238 (N_15238,N_12563,N_13816);
nor U15239 (N_15239,N_13219,N_13156);
and U15240 (N_15240,N_14730,N_14461);
nor U15241 (N_15241,N_13828,N_14607);
and U15242 (N_15242,N_14016,N_14234);
or U15243 (N_15243,N_14350,N_14436);
nand U15244 (N_15244,N_14325,N_14555);
nor U15245 (N_15245,N_12971,N_14708);
nor U15246 (N_15246,N_14770,N_14118);
and U15247 (N_15247,N_14701,N_12603);
nor U15248 (N_15248,N_14124,N_12678);
nand U15249 (N_15249,N_13095,N_14629);
xnor U15250 (N_15250,N_13973,N_13994);
nor U15251 (N_15251,N_13354,N_13826);
and U15252 (N_15252,N_14742,N_14358);
and U15253 (N_15253,N_12673,N_13940);
and U15254 (N_15254,N_14842,N_13465);
or U15255 (N_15255,N_13637,N_13381);
nand U15256 (N_15256,N_14974,N_14890);
nor U15257 (N_15257,N_12516,N_12743);
nor U15258 (N_15258,N_12716,N_13636);
nand U15259 (N_15259,N_13402,N_14689);
and U15260 (N_15260,N_13489,N_13210);
xnor U15261 (N_15261,N_12982,N_13691);
or U15262 (N_15262,N_13608,N_14755);
and U15263 (N_15263,N_13977,N_13476);
nor U15264 (N_15264,N_13260,N_14687);
nor U15265 (N_15265,N_13005,N_13682);
xor U15266 (N_15266,N_13307,N_14005);
nor U15267 (N_15267,N_14512,N_14855);
nand U15268 (N_15268,N_13434,N_14997);
and U15269 (N_15269,N_14818,N_12625);
nand U15270 (N_15270,N_14804,N_14189);
or U15271 (N_15271,N_14457,N_13228);
xor U15272 (N_15272,N_14597,N_12866);
and U15273 (N_15273,N_14031,N_14891);
or U15274 (N_15274,N_12977,N_13741);
and U15275 (N_15275,N_13211,N_14806);
nor U15276 (N_15276,N_14582,N_13695);
nor U15277 (N_15277,N_12974,N_12696);
nand U15278 (N_15278,N_14462,N_14307);
nor U15279 (N_15279,N_12786,N_12901);
nand U15280 (N_15280,N_14470,N_13471);
or U15281 (N_15281,N_14483,N_12547);
or U15282 (N_15282,N_13323,N_14058);
or U15283 (N_15283,N_14385,N_14023);
xnor U15284 (N_15284,N_13472,N_14020);
nor U15285 (N_15285,N_14047,N_13180);
or U15286 (N_15286,N_12564,N_14071);
and U15287 (N_15287,N_13618,N_14874);
nor U15288 (N_15288,N_14191,N_14352);
and U15289 (N_15289,N_13430,N_14920);
or U15290 (N_15290,N_13028,N_13825);
nor U15291 (N_15291,N_13003,N_12973);
and U15292 (N_15292,N_13676,N_14513);
or U15293 (N_15293,N_13675,N_13438);
nor U15294 (N_15294,N_13270,N_12789);
xor U15295 (N_15295,N_14500,N_13350);
xnor U15296 (N_15296,N_13019,N_14502);
nor U15297 (N_15297,N_12848,N_14907);
nand U15298 (N_15298,N_13085,N_12787);
or U15299 (N_15299,N_13196,N_14731);
xnor U15300 (N_15300,N_14869,N_14324);
nand U15301 (N_15301,N_14301,N_14110);
nor U15302 (N_15302,N_13878,N_13462);
and U15303 (N_15303,N_13520,N_14238);
and U15304 (N_15304,N_12526,N_13822);
xor U15305 (N_15305,N_12561,N_14724);
xor U15306 (N_15306,N_12768,N_13321);
xor U15307 (N_15307,N_14843,N_14446);
and U15308 (N_15308,N_14173,N_13242);
nand U15309 (N_15309,N_14305,N_12784);
and U15310 (N_15310,N_14036,N_14828);
xor U15311 (N_15311,N_13305,N_12727);
nand U15312 (N_15312,N_12836,N_14389);
nand U15313 (N_15313,N_14299,N_14026);
xnor U15314 (N_15314,N_14822,N_14390);
nor U15315 (N_15315,N_13590,N_14762);
xnor U15316 (N_15316,N_13866,N_12505);
or U15317 (N_15317,N_14144,N_13046);
xnor U15318 (N_15318,N_13992,N_13817);
xor U15319 (N_15319,N_12940,N_13926);
nor U15320 (N_15320,N_13535,N_14659);
nand U15321 (N_15321,N_14057,N_12674);
and U15322 (N_15322,N_12885,N_13124);
or U15323 (N_15323,N_14674,N_14774);
and U15324 (N_15324,N_14277,N_13751);
and U15325 (N_15325,N_14073,N_14557);
and U15326 (N_15326,N_14581,N_13301);
nand U15327 (N_15327,N_12638,N_13996);
nor U15328 (N_15328,N_14090,N_14428);
or U15329 (N_15329,N_14983,N_12736);
nor U15330 (N_15330,N_12525,N_12698);
nor U15331 (N_15331,N_12988,N_12804);
or U15332 (N_15332,N_13143,N_12909);
nand U15333 (N_15333,N_13222,N_14248);
nand U15334 (N_15334,N_12595,N_13987);
nand U15335 (N_15335,N_12854,N_13611);
nand U15336 (N_15336,N_13886,N_12904);
nand U15337 (N_15337,N_13829,N_13101);
xor U15338 (N_15338,N_13106,N_14480);
and U15339 (N_15339,N_14562,N_13128);
and U15340 (N_15340,N_14205,N_13181);
and U15341 (N_15341,N_13650,N_13079);
and U15342 (N_15342,N_14959,N_14683);
and U15343 (N_15343,N_14777,N_14121);
and U15344 (N_15344,N_13394,N_13594);
nand U15345 (N_15345,N_14875,N_13597);
nor U15346 (N_15346,N_14421,N_13875);
nor U15347 (N_15347,N_13853,N_13654);
or U15348 (N_15348,N_13635,N_13154);
and U15349 (N_15349,N_13718,N_13740);
nand U15350 (N_15350,N_14130,N_14794);
or U15351 (N_15351,N_13902,N_13329);
nand U15352 (N_15352,N_14948,N_14625);
xor U15353 (N_15353,N_14781,N_13752);
and U15354 (N_15354,N_12851,N_12978);
or U15355 (N_15355,N_14713,N_12508);
xor U15356 (N_15356,N_13306,N_14928);
nand U15357 (N_15357,N_14779,N_13130);
and U15358 (N_15358,N_13077,N_12604);
or U15359 (N_15359,N_13966,N_14244);
nor U15360 (N_15360,N_14079,N_13979);
nand U15361 (N_15361,N_14387,N_14904);
or U15362 (N_15362,N_14185,N_13689);
or U15363 (N_15363,N_12795,N_12539);
nor U15364 (N_15364,N_13571,N_12893);
or U15365 (N_15365,N_13705,N_14679);
xnor U15366 (N_15366,N_14196,N_14628);
and U15367 (N_15367,N_14571,N_13537);
or U15368 (N_15368,N_14814,N_13839);
xnor U15369 (N_15369,N_13909,N_13344);
xor U15370 (N_15370,N_12959,N_13723);
xor U15371 (N_15371,N_13647,N_13577);
and U15372 (N_15372,N_13352,N_14878);
and U15373 (N_15373,N_13199,N_13446);
nand U15374 (N_15374,N_14166,N_12859);
or U15375 (N_15375,N_14095,N_12907);
or U15376 (N_15376,N_13400,N_12597);
nor U15377 (N_15377,N_12749,N_13324);
and U15378 (N_15378,N_13464,N_14943);
nor U15379 (N_15379,N_12543,N_14685);
nor U15380 (N_15380,N_14097,N_13652);
or U15381 (N_15381,N_14105,N_14559);
nand U15382 (N_15382,N_13161,N_13712);
and U15383 (N_15383,N_14091,N_14086);
nor U15384 (N_15384,N_14509,N_14567);
and U15385 (N_15385,N_13393,N_14087);
xor U15386 (N_15386,N_13892,N_12887);
nor U15387 (N_15387,N_13683,N_13195);
and U15388 (N_15388,N_14805,N_13122);
nand U15389 (N_15389,N_14761,N_14293);
nor U15390 (N_15390,N_14478,N_14926);
or U15391 (N_15391,N_14337,N_14034);
and U15392 (N_15392,N_13399,N_13770);
and U15393 (N_15393,N_12740,N_13052);
xnor U15394 (N_15394,N_14613,N_13858);
xor U15395 (N_15395,N_13454,N_14316);
or U15396 (N_15396,N_14941,N_13327);
nor U15397 (N_15397,N_12536,N_14848);
xnor U15398 (N_15398,N_14249,N_13236);
and U15399 (N_15399,N_14199,N_14092);
and U15400 (N_15400,N_13484,N_14202);
and U15401 (N_15401,N_14028,N_13123);
and U15402 (N_15402,N_14361,N_12925);
nand U15403 (N_15403,N_13930,N_13591);
or U15404 (N_15404,N_14319,N_12598);
nor U15405 (N_15405,N_13997,N_14737);
nor U15406 (N_15406,N_13061,N_12572);
nand U15407 (N_15407,N_12534,N_12989);
xor U15408 (N_15408,N_13976,N_14491);
or U15409 (N_15409,N_12741,N_14621);
or U15410 (N_15410,N_12984,N_13392);
nand U15411 (N_15411,N_13868,N_14326);
nor U15412 (N_15412,N_13753,N_14936);
and U15413 (N_15413,N_12834,N_12687);
nand U15414 (N_15414,N_14107,N_13661);
or U15415 (N_15415,N_12794,N_12844);
nand U15416 (N_15416,N_13600,N_13109);
nand U15417 (N_15417,N_14030,N_13041);
nand U15418 (N_15418,N_12511,N_12770);
xnor U15419 (N_15419,N_12600,N_13413);
xnor U15420 (N_15420,N_13795,N_12898);
and U15421 (N_15421,N_14927,N_12661);
nand U15422 (N_15422,N_13499,N_14055);
and U15423 (N_15423,N_14220,N_12998);
or U15424 (N_15424,N_14807,N_12655);
nand U15425 (N_15425,N_13703,N_12560);
nand U15426 (N_15426,N_13004,N_13530);
or U15427 (N_15427,N_13850,N_14171);
or U15428 (N_15428,N_13049,N_14450);
xor U15429 (N_15429,N_14847,N_13907);
xor U15430 (N_15430,N_14542,N_13110);
nor U15431 (N_15431,N_14523,N_13229);
or U15432 (N_15432,N_14052,N_13512);
and U15433 (N_15433,N_12897,N_14009);
and U15434 (N_15434,N_14789,N_14364);
and U15435 (N_15435,N_12972,N_13849);
or U15436 (N_15436,N_14321,N_14860);
or U15437 (N_15437,N_13728,N_13627);
nor U15438 (N_15438,N_13312,N_14744);
nand U15439 (N_15439,N_13602,N_14538);
nor U15440 (N_15440,N_14340,N_13506);
nor U15441 (N_15441,N_14733,N_13628);
nor U15442 (N_15442,N_14403,N_14570);
xor U15443 (N_15443,N_13371,N_13083);
nand U15444 (N_15444,N_14314,N_14823);
xnor U15445 (N_15445,N_13065,N_13375);
nand U15446 (N_15446,N_13377,N_13388);
xor U15447 (N_15447,N_14965,N_14988);
or U15448 (N_15448,N_13027,N_12521);
or U15449 (N_15449,N_13831,N_12509);
and U15450 (N_15450,N_12500,N_13521);
nor U15451 (N_15451,N_12535,N_14042);
nor U15452 (N_15452,N_12966,N_13326);
or U15453 (N_15453,N_14206,N_12990);
and U15454 (N_15454,N_13495,N_14114);
nor U15455 (N_15455,N_13846,N_13086);
nor U15456 (N_15456,N_13081,N_13129);
nand U15457 (N_15457,N_13452,N_12748);
nand U15458 (N_15458,N_13074,N_13330);
nand U15459 (N_15459,N_14850,N_13363);
and U15460 (N_15460,N_14750,N_13579);
and U15461 (N_15461,N_13848,N_13084);
and U15462 (N_15462,N_13238,N_12896);
nor U15463 (N_15463,N_14910,N_13911);
and U15464 (N_15464,N_13539,N_14788);
nand U15465 (N_15465,N_12826,N_13043);
nor U15466 (N_15466,N_14363,N_12899);
and U15467 (N_15467,N_13112,N_12976);
xor U15468 (N_15468,N_14896,N_12889);
or U15469 (N_15469,N_13664,N_14156);
or U15470 (N_15470,N_14113,N_13899);
nand U15471 (N_15471,N_14360,N_12506);
and U15472 (N_15472,N_13405,N_14726);
xor U15473 (N_15473,N_13020,N_14335);
and U15474 (N_15474,N_14525,N_14516);
xor U15475 (N_15475,N_14064,N_13674);
and U15476 (N_15476,N_14336,N_12750);
xnor U15477 (N_15477,N_13493,N_13999);
and U15478 (N_15478,N_13437,N_14647);
nor U15479 (N_15479,N_13239,N_14758);
nand U15480 (N_15480,N_13387,N_14884);
nand U15481 (N_15481,N_14388,N_14153);
nor U15482 (N_15482,N_12568,N_14594);
or U15483 (N_15483,N_14535,N_12882);
xnor U15484 (N_15484,N_12570,N_12759);
or U15485 (N_15485,N_12823,N_14435);
and U15486 (N_15486,N_13206,N_12608);
nor U15487 (N_15487,N_13240,N_13480);
nor U15488 (N_15488,N_13882,N_12513);
or U15489 (N_15489,N_12587,N_12814);
nand U15490 (N_15490,N_13153,N_14211);
and U15491 (N_15491,N_13459,N_13617);
nand U15492 (N_15492,N_14309,N_12664);
or U15493 (N_15493,N_13666,N_12765);
and U15494 (N_15494,N_12965,N_13500);
nor U15495 (N_15495,N_13336,N_14150);
nor U15496 (N_15496,N_12744,N_13927);
and U15497 (N_15497,N_13541,N_14231);
and U15498 (N_15498,N_14682,N_14159);
and U15499 (N_15499,N_13466,N_14423);
nor U15500 (N_15500,N_12902,N_13508);
and U15501 (N_15501,N_13470,N_14598);
nand U15502 (N_15502,N_14528,N_14808);
nor U15503 (N_15503,N_14116,N_13155);
or U15504 (N_15504,N_12954,N_14344);
nand U15505 (N_15505,N_14485,N_14379);
nand U15506 (N_15506,N_13726,N_14254);
nor U15507 (N_15507,N_13598,N_13022);
and U15508 (N_15508,N_14929,N_12934);
nand U15509 (N_15509,N_13790,N_14402);
xor U15510 (N_15510,N_12644,N_14357);
xor U15511 (N_15511,N_14456,N_13837);
nor U15512 (N_15512,N_14666,N_12725);
and U15513 (N_15513,N_13818,N_13696);
nand U15514 (N_15514,N_14676,N_13543);
nor U15515 (N_15515,N_13174,N_12663);
and U15516 (N_15516,N_13528,N_13006);
and U15517 (N_15517,N_12588,N_13754);
xnor U15518 (N_15518,N_12955,N_13588);
nor U15519 (N_15519,N_13068,N_12583);
nor U15520 (N_15520,N_14645,N_14550);
and U15521 (N_15521,N_12628,N_12964);
or U15522 (N_15522,N_12712,N_14637);
and U15523 (N_15523,N_13939,N_14673);
nand U15524 (N_15524,N_14925,N_14412);
nand U15525 (N_15525,N_14841,N_14887);
xnor U15526 (N_15526,N_14510,N_14760);
nor U15527 (N_15527,N_14720,N_12549);
and U15528 (N_15528,N_13072,N_13133);
and U15529 (N_15529,N_14082,N_13678);
nor U15530 (N_15530,N_13088,N_14496);
and U15531 (N_15531,N_14000,N_13044);
xor U15532 (N_15532,N_12713,N_13765);
or U15533 (N_15533,N_14184,N_12694);
or U15534 (N_15534,N_14957,N_14696);
and U15535 (N_15535,N_13990,N_13777);
nor U15536 (N_15536,N_14815,N_13144);
nor U15537 (N_15537,N_12669,N_13801);
nand U15538 (N_15538,N_14686,N_13212);
and U15539 (N_15539,N_13861,N_14566);
or U15540 (N_15540,N_14656,N_13599);
and U15541 (N_15541,N_14778,N_14362);
nand U15542 (N_15542,N_13424,N_13356);
nand U15543 (N_15543,N_13633,N_14380);
nand U15544 (N_15544,N_13835,N_14706);
and U15545 (N_15545,N_12639,N_14719);
nor U15546 (N_15546,N_13929,N_14472);
or U15547 (N_15547,N_13175,N_13980);
nor U15548 (N_15548,N_13257,N_13706);
nor U15549 (N_15549,N_14800,N_12711);
nor U15550 (N_15550,N_14715,N_14738);
and U15551 (N_15551,N_14650,N_14864);
nor U15552 (N_15552,N_14349,N_13538);
xor U15553 (N_15553,N_13947,N_14330);
xnor U15554 (N_15554,N_14757,N_13655);
xnor U15555 (N_15555,N_13220,N_14161);
xor U15556 (N_15556,N_13436,N_14374);
nand U15557 (N_15557,N_13249,N_14622);
nor U15558 (N_15558,N_12637,N_12888);
and U15559 (N_15559,N_14651,N_14705);
and U15560 (N_15560,N_13607,N_13169);
and U15561 (N_15561,N_12532,N_12654);
xor U15562 (N_15562,N_13584,N_14280);
and U15563 (N_15563,N_13191,N_14215);
nand U15564 (N_15564,N_14225,N_13285);
nand U15565 (N_15565,N_12811,N_14675);
nand U15566 (N_15566,N_13457,N_14230);
and U15567 (N_15567,N_13710,N_14329);
nor U15568 (N_15568,N_13988,N_14076);
xor U15569 (N_15569,N_14192,N_14444);
nor U15570 (N_15570,N_13445,N_14817);
nand U15571 (N_15571,N_13362,N_13291);
and U15572 (N_15572,N_13815,N_13578);
xnor U15573 (N_15573,N_14868,N_12708);
or U15574 (N_15574,N_13293,N_14998);
xor U15575 (N_15575,N_14505,N_14445);
and U15576 (N_15576,N_13524,N_13559);
nand U15577 (N_15577,N_12858,N_12810);
xnor U15578 (N_15578,N_12994,N_14729);
xor U15579 (N_15579,N_14590,N_14494);
nand U15580 (N_15580,N_13040,N_13132);
or U15581 (N_15581,N_12697,N_13485);
nand U15582 (N_15582,N_12747,N_12933);
and U15583 (N_15583,N_13745,N_13583);
and U15584 (N_15584,N_14029,N_13348);
and U15585 (N_15585,N_13298,N_14977);
nand U15586 (N_15586,N_13208,N_12841);
nand U15587 (N_15587,N_14551,N_13732);
nand U15588 (N_15588,N_13280,N_13029);
xor U15589 (N_15589,N_14881,N_14966);
and U15590 (N_15590,N_12918,N_13570);
nand U15591 (N_15591,N_12703,N_13821);
nor U15592 (N_15592,N_13807,N_13898);
xor U15593 (N_15593,N_14749,N_12905);
and U15594 (N_15594,N_14348,N_13663);
xnor U15595 (N_15595,N_14276,N_12731);
and U15596 (N_15596,N_14300,N_14094);
or U15597 (N_15597,N_12775,N_12518);
and U15598 (N_15598,N_13150,N_13094);
xor U15599 (N_15599,N_14183,N_14490);
nor U15600 (N_15600,N_13341,N_14187);
nor U15601 (N_15601,N_14955,N_12569);
or U15602 (N_15602,N_13698,N_14775);
or U15603 (N_15603,N_14488,N_14394);
or U15604 (N_15604,N_14398,N_12788);
nand U15605 (N_15605,N_14534,N_13231);
or U15606 (N_15606,N_14477,N_14203);
or U15607 (N_15607,N_14657,N_13214);
and U15608 (N_15608,N_12531,N_13842);
and U15609 (N_15609,N_13871,N_13615);
nor U15610 (N_15610,N_13529,N_14934);
and U15611 (N_15611,N_12931,N_13184);
xor U15612 (N_15612,N_13808,N_13425);
xnor U15613 (N_15613,N_14101,N_13717);
xnor U15614 (N_15614,N_13246,N_14400);
nand U15615 (N_15615,N_14859,N_13759);
xor U15616 (N_15616,N_13854,N_14958);
and U15617 (N_15617,N_12546,N_14169);
nor U15618 (N_15618,N_14332,N_13045);
nand U15619 (N_15619,N_14846,N_13702);
or U15620 (N_15620,N_13959,N_12886);
nor U15621 (N_15621,N_12662,N_14592);
and U15622 (N_15622,N_13667,N_14367);
nand U15623 (N_15623,N_12812,N_12796);
xnor U15624 (N_15624,N_14530,N_14290);
or U15625 (N_15625,N_13035,N_14635);
nand U15626 (N_15626,N_12620,N_12970);
nor U15627 (N_15627,N_14982,N_13340);
nand U15628 (N_15628,N_14583,N_13254);
xor U15629 (N_15629,N_13098,N_13550);
and U15630 (N_15630,N_13295,N_14046);
or U15631 (N_15631,N_14062,N_14857);
and U15632 (N_15632,N_14830,N_13230);
nand U15633 (N_15633,N_14260,N_13653);
or U15634 (N_15634,N_13642,N_13544);
or U15635 (N_15635,N_14168,N_14136);
or U15636 (N_15636,N_13755,N_14194);
xor U15637 (N_15637,N_13075,N_14083);
xor U15638 (N_15638,N_14233,N_14644);
xor U15639 (N_15639,N_14527,N_13444);
or U15640 (N_15640,N_12979,N_12672);
nor U15641 (N_15641,N_13748,N_12791);
nand U15642 (N_15642,N_14175,N_13786);
and U15643 (N_15643,N_14602,N_13406);
or U15644 (N_15644,N_14663,N_14727);
nand U15645 (N_15645,N_13378,N_14167);
nand U15646 (N_15646,N_12833,N_13054);
and U15647 (N_15647,N_14816,N_13137);
nand U15648 (N_15648,N_14041,N_13949);
and U15649 (N_15649,N_12692,N_12630);
xor U15650 (N_15650,N_14198,N_14954);
nor U15651 (N_15651,N_13501,N_14006);
and U15652 (N_15652,N_13261,N_14903);
or U15653 (N_15653,N_12869,N_13804);
nor U15654 (N_15654,N_14067,N_13551);
or U15655 (N_15655,N_14413,N_13679);
nand U15656 (N_15656,N_12714,N_14414);
and U15657 (N_15657,N_14463,N_12806);
xnor U15658 (N_15658,N_13511,N_14065);
and U15659 (N_15659,N_14697,N_13609);
nand U15660 (N_15660,N_14122,N_14576);
and U15661 (N_15661,N_14960,N_14837);
nor U15662 (N_15662,N_14952,N_14038);
xnor U15663 (N_15663,N_13064,N_13107);
xnor U15664 (N_15664,N_14019,N_12634);
nor U15665 (N_15665,N_13796,N_13923);
nor U15666 (N_15666,N_14208,N_12624);
nand U15667 (N_15667,N_14972,N_13273);
or U15668 (N_15668,N_13542,N_13369);
nand U15669 (N_15669,N_14840,N_13218);
nand U15670 (N_15670,N_14951,N_13938);
nand U15671 (N_15671,N_12660,N_13630);
or U15672 (N_15672,N_14239,N_13563);
or U15673 (N_15673,N_12951,N_14979);
nand U15674 (N_15674,N_14978,N_12653);
nand U15675 (N_15675,N_14563,N_14356);
or U15676 (N_15676,N_13165,N_12803);
or U15677 (N_15677,N_14267,N_12863);
or U15678 (N_15678,N_13398,N_14924);
or U15679 (N_15679,N_12648,N_14393);
and U15680 (N_15680,N_13365,N_13047);
and U15681 (N_15681,N_14370,N_14545);
or U15682 (N_15682,N_14351,N_14468);
or U15683 (N_15683,N_14085,N_13115);
and U15684 (N_15684,N_12593,N_13108);
xor U15685 (N_15685,N_12917,N_14201);
nor U15686 (N_15686,N_14944,N_14217);
nor U15687 (N_15687,N_12502,N_13482);
and U15688 (N_15688,N_12877,N_12913);
xnor U15689 (N_15689,N_14410,N_13463);
nor U15690 (N_15690,N_14540,N_14443);
nor U15691 (N_15691,N_14375,N_14265);
and U15692 (N_15692,N_13547,N_12705);
and U15693 (N_15693,N_14753,N_14584);
and U15694 (N_15694,N_13251,N_14798);
and U15695 (N_15695,N_13690,N_12868);
or U15696 (N_15696,N_12643,N_14591);
and U15697 (N_15697,N_14791,N_12824);
and U15698 (N_15698,N_12682,N_13830);
or U15699 (N_15699,N_12552,N_13163);
nand U15700 (N_15700,N_14406,N_12602);
or U15701 (N_15701,N_13431,N_14870);
nand U15702 (N_15702,N_14039,N_13606);
and U15703 (N_15703,N_12849,N_14214);
or U15704 (N_15704,N_14451,N_12945);
xnor U15705 (N_15705,N_13160,N_14900);
and U15706 (N_15706,N_14417,N_13776);
nor U15707 (N_15707,N_12761,N_13922);
and U15708 (N_15708,N_14834,N_13978);
nor U15709 (N_15709,N_13441,N_14289);
nor U15710 (N_15710,N_13915,N_13713);
nor U15711 (N_15711,N_13769,N_14303);
and U15712 (N_15712,N_12728,N_13736);
xnor U15713 (N_15713,N_14787,N_12857);
nor U15714 (N_15714,N_14397,N_13558);
or U15715 (N_15715,N_14405,N_14586);
nand U15716 (N_15716,N_13116,N_14096);
nor U15717 (N_15717,N_13714,N_13069);
and U15718 (N_15718,N_12840,N_13126);
or U15719 (N_15719,N_14852,N_14632);
nand U15720 (N_15720,N_13809,N_13342);
nand U15721 (N_15721,N_13345,N_14004);
xor U15722 (N_15722,N_14002,N_13800);
and U15723 (N_15723,N_13189,N_14286);
or U15724 (N_15724,N_13933,N_14240);
or U15725 (N_15725,N_14913,N_12517);
nand U15726 (N_15726,N_13610,N_14382);
xnor U15727 (N_15727,N_13863,N_13596);
nor U15728 (N_15728,N_14670,N_13533);
nor U15729 (N_15729,N_12845,N_14213);
nor U15730 (N_15730,N_12715,N_12778);
nor U15731 (N_15731,N_14127,N_14495);
nand U15732 (N_15732,N_14297,N_13932);
xnor U15733 (N_15733,N_14888,N_12658);
nor U15734 (N_15734,N_13946,N_14768);
or U15735 (N_15735,N_13595,N_13286);
and U15736 (N_15736,N_13333,N_13566);
and U15737 (N_15737,N_13747,N_14164);
nand U15738 (N_15738,N_13198,N_12911);
and U15739 (N_15739,N_13403,N_13426);
and U15740 (N_15740,N_12559,N_13614);
and U15741 (N_15741,N_14790,N_14448);
nand U15742 (N_15742,N_12629,N_13490);
nand U15743 (N_15743,N_14152,N_12953);
or U15744 (N_15744,N_13120,N_12688);
nor U15745 (N_15745,N_13958,N_13621);
xor U15746 (N_15746,N_14552,N_14273);
nand U15747 (N_15747,N_13827,N_14725);
nand U15748 (N_15748,N_14518,N_12504);
or U15749 (N_15749,N_13009,N_13934);
nand U15750 (N_15750,N_14032,N_14283);
nand U15751 (N_15751,N_14070,N_12730);
and U15752 (N_15752,N_13780,N_13408);
and U15753 (N_15753,N_14908,N_14547);
or U15754 (N_15754,N_14812,N_12567);
nor U15755 (N_15755,N_13447,N_14801);
or U15756 (N_15756,N_14245,N_12753);
nor U15757 (N_15757,N_13767,N_13415);
xnor U15758 (N_15758,N_14766,N_14246);
and U15759 (N_15759,N_13346,N_14053);
nand U15760 (N_15760,N_13974,N_14803);
nand U15761 (N_15761,N_13944,N_13787);
nand U15762 (N_15762,N_12636,N_14313);
or U15763 (N_15763,N_13272,N_13073);
xor U15764 (N_15764,N_14655,N_13738);
xor U15765 (N_15765,N_13991,N_13813);
nor U15766 (N_15766,N_14968,N_14795);
nand U15767 (N_15767,N_14408,N_13936);
and U15768 (N_15768,N_13838,N_13982);
nand U15769 (N_15769,N_14885,N_14994);
nor U15770 (N_15770,N_14521,N_13505);
and U15771 (N_15771,N_14080,N_13263);
nor U15772 (N_15772,N_12837,N_13657);
nand U15773 (N_15773,N_14633,N_13458);
nor U15774 (N_15774,N_14631,N_13644);
and U15775 (N_15775,N_14515,N_13186);
and U15776 (N_15776,N_13067,N_13134);
nor U15777 (N_15777,N_14862,N_14825);
or U15778 (N_15778,N_13895,N_13139);
nor U15779 (N_15779,N_14942,N_14608);
xor U15780 (N_15780,N_13367,N_13956);
and U15781 (N_15781,N_13612,N_13673);
nor U15782 (N_15782,N_13477,N_14170);
nor U15783 (N_15783,N_13641,N_14498);
xor U15784 (N_15784,N_14204,N_13297);
nand U15785 (N_15785,N_12890,N_14568);
and U15786 (N_15786,N_14050,N_13562);
nand U15787 (N_15787,N_14640,N_12557);
or U15788 (N_15788,N_14284,N_13970);
nor U15789 (N_15789,N_13390,N_13925);
nand U15790 (N_15790,N_14937,N_14872);
or U15791 (N_15791,N_12670,N_13449);
and U15792 (N_15792,N_14368,N_13146);
nand U15793 (N_15793,N_14377,N_12820);
nor U15794 (N_15794,N_14132,N_13190);
xor U15795 (N_15795,N_14210,N_14147);
xnor U15796 (N_15796,N_14764,N_13226);
and U15797 (N_15797,N_12916,N_14354);
nor U15798 (N_15798,N_14378,N_12782);
xor U15799 (N_15799,N_12707,N_12948);
xor U15800 (N_15800,N_13320,N_12522);
xor U15801 (N_15801,N_13172,N_13151);
nor U15802 (N_15802,N_13681,N_14353);
xnor U15803 (N_15803,N_13901,N_13904);
and U15804 (N_15804,N_13613,N_13890);
or U15805 (N_15805,N_12679,N_12649);
xor U15806 (N_15806,N_12967,N_12704);
xor U15807 (N_15807,N_13693,N_13428);
or U15808 (N_15808,N_14985,N_13414);
or U15809 (N_15809,N_13296,N_14624);
and U15810 (N_15810,N_14278,N_14251);
xor U15811 (N_15811,N_13766,N_14961);
and U15812 (N_15812,N_13639,N_12957);
or U15813 (N_15813,N_12798,N_13168);
nand U15814 (N_15814,N_12805,N_14061);
and U15815 (N_15815,N_13176,N_14182);
xor U15816 (N_15816,N_12991,N_14854);
xnor U15817 (N_15817,N_14641,N_13440);
and U15818 (N_15818,N_14606,N_13948);
and U15819 (N_15819,N_14707,N_14785);
nor U15820 (N_15820,N_13797,N_13536);
nand U15821 (N_15821,N_12864,N_14342);
or U15822 (N_15822,N_12831,N_12734);
or U15823 (N_15823,N_13889,N_13159);
and U15824 (N_15824,N_12949,N_13266);
or U15825 (N_15825,N_14373,N_13715);
xor U15826 (N_15826,N_13359,N_13023);
nor U15827 (N_15827,N_13984,N_13104);
and U15828 (N_15828,N_14549,N_12920);
or U15829 (N_15829,N_13699,N_12908);
nor U15830 (N_15830,N_14626,N_13001);
or U15831 (N_15831,N_14074,N_13177);
nor U15832 (N_15832,N_13200,N_13170);
nand U15833 (N_15833,N_13962,N_14499);
nand U15834 (N_15834,N_12683,N_12767);
or U15835 (N_15835,N_12581,N_12659);
and U15836 (N_15836,N_14419,N_14507);
or U15837 (N_15837,N_13725,N_13708);
nor U15838 (N_15838,N_14824,N_13971);
and U15839 (N_15839,N_14693,N_13859);
or U15840 (N_15840,N_13103,N_12680);
or U15841 (N_15841,N_12935,N_14474);
nor U15842 (N_15842,N_13952,N_14556);
xnor U15843 (N_15843,N_12585,N_13007);
nand U15844 (N_15844,N_13347,N_13314);
nor U15845 (N_15845,N_13488,N_13376);
and U15846 (N_15846,N_12813,N_14291);
nor U15847 (N_15847,N_13287,N_14949);
nor U15848 (N_15848,N_14612,N_12645);
nor U15849 (N_15849,N_13401,N_12919);
nor U15850 (N_15850,N_14853,N_12781);
nor U15851 (N_15851,N_14541,N_12872);
nand U15852 (N_15852,N_13805,N_14021);
nor U15853 (N_15853,N_13532,N_14037);
nand U15854 (N_15854,N_13803,N_13216);
or U15855 (N_15855,N_14553,N_13015);
or U15856 (N_15856,N_12554,N_14748);
and U15857 (N_15857,N_13138,N_13097);
nor U15858 (N_15858,N_14322,N_12545);
and U15859 (N_15859,N_14662,N_13456);
nor U15860 (N_15860,N_13221,N_14176);
nor U15861 (N_15861,N_14714,N_13919);
nor U15862 (N_15862,N_13225,N_14117);
nand U15863 (N_15863,N_13760,N_13503);
nor U15864 (N_15864,N_12514,N_13053);
or U15865 (N_15865,N_14359,N_14991);
or U15866 (N_15866,N_14430,N_13385);
nor U15867 (N_15867,N_12835,N_14867);
nand U15868 (N_15868,N_14543,N_12556);
nand U15869 (N_15869,N_13164,N_13182);
or U15870 (N_15870,N_14181,N_14648);
xnor U15871 (N_15871,N_13090,N_13756);
xnor U15872 (N_15872,N_14880,N_14422);
or U15873 (N_15873,N_13487,N_13568);
nor U15874 (N_15874,N_13688,N_14894);
and U15875 (N_15875,N_12721,N_14001);
xor U15876 (N_15876,N_12956,N_14346);
nand U15877 (N_15877,N_13416,N_14901);
and U15878 (N_15878,N_14138,N_13179);
or U15879 (N_15879,N_13062,N_14381);
nor U15880 (N_15880,N_13410,N_12596);
nor U15881 (N_15881,N_14599,N_12958);
nand U15882 (N_15882,N_14690,N_14177);
or U15883 (N_15883,N_14102,N_13332);
xnor U15884 (N_15884,N_14218,N_13924);
or U15885 (N_15885,N_12881,N_12895);
and U15886 (N_15886,N_14145,N_14967);
nand U15887 (N_15887,N_13145,N_13730);
nor U15888 (N_15888,N_14243,N_13008);
nand U15889 (N_15889,N_14120,N_13646);
nor U15890 (N_15890,N_14809,N_14899);
nor U15891 (N_15891,N_13758,N_13224);
and U15892 (N_15892,N_13672,N_14709);
nor U15893 (N_15893,N_14438,N_14877);
and U15894 (N_15894,N_13248,N_14865);
nor U15895 (N_15895,N_14546,N_12969);
or U15896 (N_15896,N_13626,N_12722);
nor U15897 (N_15897,N_14425,N_13942);
and U15898 (N_15898,N_14418,N_13634);
nor U15899 (N_15899,N_14160,N_13089);
nor U15900 (N_15900,N_13370,N_14700);
xor U15901 (N_15901,N_12609,N_13832);
and U15902 (N_15902,N_14638,N_14115);
xor U15903 (N_15903,N_14434,N_13419);
nor U15904 (N_15904,N_14588,N_13455);
nand U15905 (N_15905,N_12992,N_14531);
and U15906 (N_15906,N_14222,N_12575);
and U15907 (N_15907,N_13900,N_13091);
and U15908 (N_15908,N_12879,N_14533);
xnor U15909 (N_15909,N_12723,N_13879);
nand U15910 (N_15910,N_13311,N_13737);
nor U15911 (N_15911,N_14469,N_12695);
nor U15912 (N_15912,N_13722,N_14615);
xor U15913 (N_15913,N_13548,N_12975);
and U15914 (N_15914,N_14484,N_13960);
nand U15915 (N_15915,N_14459,N_13275);
or U15916 (N_15916,N_14819,N_13469);
xor U15917 (N_15917,N_14756,N_14200);
nor U15918 (N_15918,N_12635,N_13840);
xnor U15919 (N_15919,N_12884,N_13660);
and U15920 (N_15920,N_14879,N_14893);
nand U15921 (N_15921,N_14473,N_13580);
and U15922 (N_15922,N_14112,N_13569);
nand U15923 (N_15923,N_12900,N_14573);
xnor U15924 (N_15924,N_14411,N_13864);
or U15925 (N_15925,N_13197,N_14782);
nand U15926 (N_15926,N_13357,N_14455);
or U15927 (N_15927,N_14376,N_14680);
xor U15928 (N_15928,N_12914,N_12607);
nor U15929 (N_15929,N_13762,N_13625);
and U15930 (N_15930,N_14699,N_14838);
nor U15931 (N_15931,N_13443,N_13554);
and U15932 (N_15932,N_14282,N_14285);
xor U15933 (N_15933,N_14119,N_14654);
or U15934 (N_15934,N_13279,N_13945);
nand U15935 (N_15935,N_13931,N_12825);
and U15936 (N_15936,N_13268,N_13785);
nor U15937 (N_15937,N_14732,N_14609);
or U15938 (N_15938,N_14980,N_14916);
nor U15939 (N_15939,N_13834,N_13778);
nor U15940 (N_15940,N_12827,N_14658);
nand U15941 (N_15941,N_13917,N_14178);
or U15942 (N_15942,N_13709,N_13802);
and U15943 (N_15943,N_14010,N_13981);
or U15944 (N_15944,N_14015,N_13379);
nand U15945 (N_15945,N_14578,N_12709);
nor U15946 (N_15946,N_13575,N_14235);
and U15947 (N_15947,N_13574,N_12528);
and U15948 (N_15948,N_14956,N_12529);
or U15949 (N_15949,N_13002,N_12946);
xnor U15950 (N_15950,N_14970,N_12880);
and U15951 (N_15951,N_13148,N_12555);
or U15952 (N_15952,N_13534,N_12735);
nor U15953 (N_15953,N_13166,N_12816);
nor U15954 (N_15954,N_14620,N_14486);
and U15955 (N_15955,N_14453,N_13789);
and U15956 (N_15956,N_14288,N_14008);
nand U15957 (N_15957,N_14619,N_13993);
xor U15958 (N_15958,N_12619,N_12997);
or U15959 (N_15959,N_14946,N_14151);
xor U15960 (N_15960,N_14736,N_13885);
xnor U15961 (N_15961,N_12632,N_13284);
or U15962 (N_15962,N_13908,N_13516);
nand U15963 (N_15963,N_13916,N_14104);
xnor U15964 (N_15964,N_13038,N_13972);
and U15965 (N_15965,N_13451,N_14873);
xor U15966 (N_15966,N_13265,N_14108);
and U15967 (N_15967,N_14228,N_13080);
nand U15968 (N_15968,N_14517,N_12573);
xor U15969 (N_15969,N_14532,N_13623);
or U15970 (N_15970,N_12507,N_14902);
nand U15971 (N_15971,N_13775,N_12760);
xor U15972 (N_15972,N_14054,N_14180);
and U15973 (N_15973,N_13442,N_14973);
or U15974 (N_15974,N_14793,N_14439);
nor U15975 (N_15975,N_14308,N_12650);
and U15976 (N_15976,N_14048,N_12562);
or U15977 (N_15977,N_12942,N_13847);
xnor U15978 (N_15978,N_13274,N_14739);
nor U15979 (N_15979,N_12783,N_14999);
and U15980 (N_15980,N_13651,N_12993);
nand U15981 (N_15981,N_14315,N_12870);
or U15982 (N_15982,N_13066,N_13078);
xnor U15983 (N_15983,N_13784,N_13276);
nor U15984 (N_15984,N_13063,N_14317);
nand U15985 (N_15985,N_13386,N_13731);
xor U15986 (N_15986,N_13684,N_13963);
nor U15987 (N_15987,N_13820,N_14684);
or U15988 (N_15988,N_13303,N_14465);
nor U15989 (N_15989,N_14529,N_14197);
xnor U15990 (N_15990,N_13513,N_14964);
or U15991 (N_15991,N_12686,N_12968);
nor U15992 (N_15992,N_12774,N_12995);
and U15993 (N_15993,N_13867,N_13024);
nand U15994 (N_15994,N_14935,N_13632);
or U15995 (N_15995,N_14660,N_14011);
or U15996 (N_15996,N_13526,N_14148);
nor U15997 (N_15997,N_12691,N_12980);
nand U15998 (N_15998,N_13788,N_13264);
nor U15999 (N_15999,N_14401,N_13351);
nand U16000 (N_16000,N_14216,N_14258);
nor U16001 (N_16001,N_14272,N_14984);
xor U16002 (N_16002,N_14331,N_12699);
or U16003 (N_16003,N_13299,N_14163);
nor U16004 (N_16004,N_14025,N_12963);
nand U16005 (N_16005,N_12614,N_12878);
or U16006 (N_16006,N_12667,N_13581);
and U16007 (N_16007,N_12809,N_12668);
nor U16008 (N_16008,N_13912,N_13033);
xnor U16009 (N_16009,N_13127,N_12915);
nand U16010 (N_16010,N_12745,N_14409);
xnor U16011 (N_16011,N_13215,N_14845);
xnor U16012 (N_16012,N_14962,N_13058);
nor U16013 (N_16013,N_13207,N_12599);
nor U16014 (N_16014,N_13525,N_14242);
nor U16015 (N_16015,N_13319,N_12676);
nor U16016 (N_16016,N_14043,N_14372);
or U16017 (N_16017,N_12550,N_14458);
xor U16018 (N_16018,N_12548,N_12751);
and U16019 (N_16019,N_12861,N_13014);
or U16020 (N_16020,N_13975,N_12928);
nand U16021 (N_16021,N_13928,N_13417);
or U16022 (N_16022,N_13282,N_14856);
or U16023 (N_16023,N_12842,N_13025);
nor U16024 (N_16024,N_14256,N_14623);
nor U16025 (N_16025,N_14661,N_12983);
and U16026 (N_16026,N_14634,N_13193);
and U16027 (N_16027,N_12675,N_14040);
or U16028 (N_16028,N_13012,N_13694);
nand U16029 (N_16029,N_14539,N_14345);
and U16030 (N_16030,N_12929,N_14416);
and U16031 (N_16031,N_14537,N_14306);
nor U16032 (N_16032,N_13640,N_13453);
nor U16033 (N_16033,N_14093,N_13527);
or U16034 (N_16034,N_13704,N_14347);
or U16035 (N_16035,N_12719,N_14829);
and U16036 (N_16036,N_14668,N_14133);
nand U16037 (N_16037,N_13593,N_12616);
and U16038 (N_16038,N_12646,N_13358);
nand U16039 (N_16039,N_13620,N_13824);
nor U16040 (N_16040,N_14338,N_12924);
and U16041 (N_16041,N_13317,N_14898);
or U16042 (N_16042,N_14072,N_14027);
xnor U16043 (N_16043,N_14190,N_13244);
nand U16044 (N_16044,N_13763,N_14746);
or U16045 (N_16045,N_12651,N_13662);
nor U16046 (N_16046,N_13468,N_13950);
and U16047 (N_16047,N_14207,N_12589);
nor U16048 (N_16048,N_14432,N_12617);
xor U16049 (N_16049,N_14931,N_14771);
xor U16050 (N_16050,N_14221,N_13383);
nand U16051 (N_16051,N_14497,N_13967);
or U16052 (N_16052,N_13557,N_14922);
xor U16053 (N_16053,N_14075,N_13183);
nand U16054 (N_16054,N_13173,N_14963);
or U16055 (N_16055,N_14143,N_13743);
or U16056 (N_16056,N_14487,N_13658);
and U16057 (N_16057,N_14813,N_14833);
and U16058 (N_16058,N_13518,N_12742);
or U16059 (N_16059,N_13071,N_14396);
xor U16060 (N_16060,N_14236,N_14437);
nor U16061 (N_16061,N_12776,N_13823);
and U16062 (N_16062,N_14123,N_14751);
nor U16063 (N_16063,N_12936,N_13059);
or U16064 (N_16064,N_14826,N_14269);
xnor U16065 (N_16065,N_13361,N_12764);
or U16066 (N_16066,N_13397,N_13771);
and U16067 (N_16067,N_14223,N_12530);
nand U16068 (N_16068,N_14012,N_13685);
xnor U16069 (N_16069,N_12822,N_13561);
or U16070 (N_16070,N_14694,N_14327);
or U16071 (N_16071,N_13985,N_13232);
or U16072 (N_16072,N_13380,N_13638);
nor U16073 (N_16073,N_13806,N_13421);
xor U16074 (N_16074,N_14627,N_13255);
or U16075 (N_16075,N_13467,N_14765);
nand U16076 (N_16076,N_12850,N_14717);
and U16077 (N_16077,N_14618,N_13951);
or U16078 (N_16078,N_14482,N_12612);
nor U16079 (N_16079,N_14287,N_14369);
and U16080 (N_16080,N_13798,N_13857);
xor U16081 (N_16081,N_12930,N_13034);
nor U16082 (N_16082,N_14939,N_12578);
nor U16083 (N_16083,N_14227,N_14429);
nor U16084 (N_16084,N_14142,N_14851);
or U16085 (N_16085,N_12601,N_12987);
nand U16086 (N_16086,N_13000,N_14224);
or U16087 (N_16087,N_13360,N_14692);
nand U16088 (N_16088,N_14341,N_13209);
xnor U16089 (N_16089,N_13565,N_13734);
nand U16090 (N_16090,N_12832,N_14193);
xnor U16091 (N_16091,N_14460,N_14033);
nand U16092 (N_16092,N_13964,N_14247);
nand U16093 (N_16093,N_13629,N_14767);
or U16094 (N_16094,N_13056,N_12618);
nand U16095 (N_16095,N_12610,N_12817);
and U16096 (N_16096,N_12710,N_12846);
and U16097 (N_16097,N_14747,N_14745);
nor U16098 (N_16098,N_13131,N_13233);
nand U16099 (N_16099,N_14892,N_12892);
xnor U16100 (N_16100,N_13237,N_14595);
nor U16101 (N_16101,N_14835,N_14365);
or U16102 (N_16102,N_13450,N_14195);
nor U16103 (N_16103,N_12590,N_14780);
or U16104 (N_16104,N_14035,N_14630);
and U16105 (N_16105,N_13429,N_13349);
xor U16106 (N_16106,N_14219,N_13515);
and U16107 (N_16107,N_13241,N_13913);
nor U16108 (N_16108,N_14310,N_12923);
nor U16109 (N_16109,N_12656,N_13819);
nor U16110 (N_16110,N_14754,N_14861);
nor U16111 (N_16111,N_12642,N_14137);
nand U16112 (N_16112,N_13026,N_14125);
xnor U16113 (N_16113,N_14415,N_14279);
nor U16114 (N_16114,N_12580,N_13905);
or U16115 (N_16115,N_13894,N_12631);
xnor U16116 (N_16116,N_13768,N_14565);
or U16117 (N_16117,N_14013,N_12732);
and U16118 (N_16118,N_14504,N_13910);
nand U16119 (N_16119,N_14871,N_14044);
xnor U16120 (N_16120,N_12606,N_13781);
nand U16121 (N_16121,N_14792,N_13668);
or U16122 (N_16122,N_14603,N_13852);
nand U16123 (N_16123,N_13519,N_13721);
xor U16124 (N_16124,N_13865,N_14172);
nor U16125 (N_16125,N_14262,N_14511);
and U16126 (N_16126,N_13099,N_14088);
nand U16127 (N_16127,N_14131,N_14564);
xor U16128 (N_16128,N_14212,N_13331);
and U16129 (N_16129,N_13514,N_13502);
or U16130 (N_16130,N_13372,N_13334);
nand U16131 (N_16131,N_12515,N_13669);
and U16132 (N_16132,N_13460,N_14188);
xnor U16133 (N_16133,N_13316,N_13692);
nor U16134 (N_16134,N_14646,N_14399);
nand U16135 (N_16135,N_13076,N_14716);
and U16136 (N_16136,N_14969,N_14721);
and U16137 (N_16137,N_13937,N_12701);
nor U16138 (N_16138,N_12921,N_13582);
xor U16139 (N_16139,N_12912,N_13483);
nand U16140 (N_16140,N_12755,N_14671);
or U16141 (N_16141,N_14802,N_13253);
or U16142 (N_16142,N_13435,N_13325);
xor U16143 (N_16143,N_12875,N_14975);
and U16144 (N_16144,N_14268,N_13531);
nor U16145 (N_16145,N_13587,N_12579);
and U16146 (N_16146,N_13051,N_14384);
or U16147 (N_16147,N_14561,N_13294);
and U16148 (N_16148,N_14103,N_12577);
or U16149 (N_16149,N_14976,N_12540);
and U16150 (N_16150,N_13833,N_13888);
nand U16151 (N_16151,N_13586,N_13724);
nor U16152 (N_16152,N_14938,N_14604);
nor U16153 (N_16153,N_14953,N_13504);
nor U16154 (N_16154,N_13670,N_13289);
and U16155 (N_16155,N_13118,N_13016);
nor U16156 (N_16156,N_13117,N_12553);
or U16157 (N_16157,N_13136,N_12999);
xor U16158 (N_16158,N_14165,N_12807);
xor U16159 (N_16159,N_13262,N_13887);
and U16160 (N_16160,N_13645,N_12950);
nor U16161 (N_16161,N_14355,N_14407);
xnor U16162 (N_16162,N_13188,N_14839);
xnor U16163 (N_16163,N_14426,N_13409);
xnor U16164 (N_16164,N_13742,N_14045);
nor U16165 (N_16165,N_12769,N_13339);
nand U16166 (N_16166,N_13055,N_14911);
or U16167 (N_16167,N_13589,N_13422);
xor U16168 (N_16168,N_13677,N_13729);
nor U16169 (N_16169,N_13247,N_13235);
and U16170 (N_16170,N_14139,N_12752);
nor U16171 (N_16171,N_13540,N_12852);
xor U16172 (N_16172,N_14493,N_14923);
and U16173 (N_16173,N_12962,N_14089);
nor U16174 (N_16174,N_14371,N_13656);
nor U16175 (N_16175,N_14084,N_13856);
or U16176 (N_16176,N_13252,N_12797);
and U16177 (N_16177,N_14442,N_14986);
nor U16178 (N_16178,N_12544,N_14292);
nand U16179 (N_16179,N_14882,N_14492);
or U16180 (N_16180,N_13624,N_13092);
or U16181 (N_16181,N_12758,N_14832);
and U16182 (N_16182,N_14471,N_13162);
xnor U16183 (N_16183,N_14298,N_14665);
and U16184 (N_16184,N_14601,N_12985);
nor U16185 (N_16185,N_14950,N_14295);
or U16186 (N_16186,N_13918,N_13619);
or U16187 (N_16187,N_12706,N_13302);
xnor U16188 (N_16188,N_12501,N_14162);
nor U16189 (N_16189,N_13556,N_14712);
or U16190 (N_16190,N_13474,N_13167);
nor U16191 (N_16191,N_13310,N_14710);
nor U16192 (N_16192,N_14328,N_13243);
nor U16193 (N_16193,N_14889,N_13250);
or U16194 (N_16194,N_12800,N_13564);
nand U16195 (N_16195,N_13585,N_14018);
or U16196 (N_16196,N_12855,N_14186);
and U16197 (N_16197,N_14479,N_13523);
xor U16198 (N_16198,N_14996,N_13961);
nand U16199 (N_16199,N_13509,N_13017);
or U16200 (N_16200,N_12627,N_14919);
and U16201 (N_16201,N_13896,N_12582);
nand U16202 (N_16202,N_14866,N_12702);
and U16203 (N_16203,N_13278,N_13954);
xor U16204 (N_16204,N_14146,N_14536);
nand U16205 (N_16205,N_14797,N_13338);
nor U16206 (N_16206,N_13735,N_13546);
xor U16207 (N_16207,N_14681,N_14441);
nand U16208 (N_16208,N_14312,N_14703);
nand U16209 (N_16209,N_13368,N_13448);
or U16210 (N_16210,N_14698,N_14906);
xor U16211 (N_16211,N_14229,N_14945);
nand U16212 (N_16212,N_14677,N_13943);
and U16213 (N_16213,N_14526,N_12773);
xor U16214 (N_16214,N_14596,N_12551);
and U16215 (N_16215,N_14060,N_13269);
or U16216 (N_16216,N_13792,N_14158);
xnor U16217 (N_16217,N_13478,N_14773);
nor U16218 (N_16218,N_13989,N_12684);
nor U16219 (N_16219,N_13553,N_12876);
xor U16220 (N_16220,N_12891,N_12780);
xor U16221 (N_16221,N_14769,N_14266);
xnor U16222 (N_16222,N_14639,N_13374);
nand U16223 (N_16223,N_14642,N_14930);
and U16224 (N_16224,N_12693,N_14068);
or U16225 (N_16225,N_13920,N_14667);
or U16226 (N_16226,N_13258,N_13042);
xor U16227 (N_16227,N_13479,N_13290);
nand U16228 (N_16228,N_13384,N_12790);
xor U16229 (N_16229,N_14883,N_12873);
xnor U16230 (N_16230,N_13560,N_14140);
and U16231 (N_16231,N_14264,N_14261);
or U16232 (N_16232,N_13576,N_13727);
nor U16233 (N_16233,N_13998,N_12586);
nand U16234 (N_16234,N_13411,N_14918);
nor U16235 (N_16235,N_14501,N_13389);
nor U16236 (N_16236,N_14466,N_12537);
nor U16237 (N_16237,N_13772,N_13259);
nand U16238 (N_16238,N_12792,N_13475);
nor U16239 (N_16239,N_14099,N_13522);
nor U16240 (N_16240,N_13552,N_14863);
nor U16241 (N_16241,N_14063,N_13420);
or U16242 (N_16242,N_14333,N_13171);
and U16243 (N_16243,N_14577,N_13486);
nor U16244 (N_16244,N_13140,N_13036);
and U16245 (N_16245,N_14688,N_13567);
xor U16246 (N_16246,N_12584,N_14740);
nand U16247 (N_16247,N_14776,N_14669);
or U16248 (N_16248,N_12906,N_12657);
nand U16249 (N_16249,N_14250,N_14569);
nor U16250 (N_16250,N_12865,N_14651);
and U16251 (N_16251,N_14592,N_13060);
nor U16252 (N_16252,N_14165,N_14479);
nand U16253 (N_16253,N_13739,N_12809);
or U16254 (N_16254,N_13378,N_13414);
or U16255 (N_16255,N_13818,N_14761);
or U16256 (N_16256,N_14593,N_14591);
and U16257 (N_16257,N_13917,N_12671);
nor U16258 (N_16258,N_14193,N_14340);
nand U16259 (N_16259,N_14981,N_12857);
nand U16260 (N_16260,N_12576,N_13261);
or U16261 (N_16261,N_13643,N_14666);
xor U16262 (N_16262,N_13715,N_13990);
or U16263 (N_16263,N_13055,N_14216);
nand U16264 (N_16264,N_13429,N_12839);
and U16265 (N_16265,N_14054,N_14420);
xnor U16266 (N_16266,N_13499,N_14754);
xnor U16267 (N_16267,N_14811,N_12859);
and U16268 (N_16268,N_13405,N_14359);
and U16269 (N_16269,N_13216,N_14750);
xor U16270 (N_16270,N_13163,N_13932);
and U16271 (N_16271,N_14485,N_13529);
and U16272 (N_16272,N_14055,N_12909);
xor U16273 (N_16273,N_13158,N_13621);
nand U16274 (N_16274,N_14561,N_14134);
nor U16275 (N_16275,N_14460,N_14834);
and U16276 (N_16276,N_13935,N_13326);
xnor U16277 (N_16277,N_13728,N_13983);
and U16278 (N_16278,N_13254,N_13770);
or U16279 (N_16279,N_12561,N_13554);
or U16280 (N_16280,N_12655,N_13494);
or U16281 (N_16281,N_13090,N_12943);
nor U16282 (N_16282,N_14855,N_14546);
or U16283 (N_16283,N_13268,N_13094);
nand U16284 (N_16284,N_13033,N_13010);
nand U16285 (N_16285,N_13995,N_13110);
nand U16286 (N_16286,N_12882,N_13467);
xnor U16287 (N_16287,N_14247,N_13813);
nand U16288 (N_16288,N_12536,N_13652);
or U16289 (N_16289,N_14510,N_13970);
nor U16290 (N_16290,N_14023,N_13941);
and U16291 (N_16291,N_14338,N_12732);
xor U16292 (N_16292,N_13206,N_14925);
nor U16293 (N_16293,N_12613,N_12876);
or U16294 (N_16294,N_13177,N_14473);
and U16295 (N_16295,N_13688,N_14634);
and U16296 (N_16296,N_14442,N_14180);
nand U16297 (N_16297,N_12970,N_14039);
nand U16298 (N_16298,N_13303,N_14690);
nor U16299 (N_16299,N_12879,N_12909);
xnor U16300 (N_16300,N_14162,N_12812);
nand U16301 (N_16301,N_14449,N_13815);
nand U16302 (N_16302,N_14059,N_14935);
nor U16303 (N_16303,N_13015,N_12559);
xor U16304 (N_16304,N_13539,N_14587);
nor U16305 (N_16305,N_12817,N_14668);
xor U16306 (N_16306,N_14111,N_13577);
or U16307 (N_16307,N_14176,N_12511);
and U16308 (N_16308,N_13513,N_13156);
and U16309 (N_16309,N_12738,N_14053);
xor U16310 (N_16310,N_12678,N_12684);
xnor U16311 (N_16311,N_14098,N_14400);
xor U16312 (N_16312,N_14003,N_13657);
nor U16313 (N_16313,N_14572,N_14180);
or U16314 (N_16314,N_14172,N_14438);
nand U16315 (N_16315,N_13512,N_13174);
or U16316 (N_16316,N_14742,N_12778);
xor U16317 (N_16317,N_14018,N_13939);
or U16318 (N_16318,N_14577,N_12531);
nor U16319 (N_16319,N_14744,N_12887);
and U16320 (N_16320,N_13219,N_14647);
nor U16321 (N_16321,N_14869,N_14859);
nand U16322 (N_16322,N_13104,N_14401);
and U16323 (N_16323,N_14865,N_13150);
xnor U16324 (N_16324,N_13803,N_14977);
and U16325 (N_16325,N_13659,N_14724);
nor U16326 (N_16326,N_13729,N_14831);
nand U16327 (N_16327,N_14110,N_13140);
or U16328 (N_16328,N_12818,N_13690);
nand U16329 (N_16329,N_12945,N_13602);
or U16330 (N_16330,N_13495,N_13013);
nand U16331 (N_16331,N_14134,N_13555);
xnor U16332 (N_16332,N_14464,N_14579);
and U16333 (N_16333,N_13503,N_13622);
and U16334 (N_16334,N_13272,N_12984);
nand U16335 (N_16335,N_14130,N_14233);
or U16336 (N_16336,N_12706,N_14848);
or U16337 (N_16337,N_14523,N_13550);
and U16338 (N_16338,N_13447,N_12874);
xor U16339 (N_16339,N_12675,N_12687);
nand U16340 (N_16340,N_14893,N_14102);
nand U16341 (N_16341,N_14404,N_13796);
xor U16342 (N_16342,N_13932,N_13784);
and U16343 (N_16343,N_12640,N_14118);
nand U16344 (N_16344,N_13285,N_14366);
or U16345 (N_16345,N_13237,N_13410);
nand U16346 (N_16346,N_12734,N_13885);
or U16347 (N_16347,N_12754,N_14332);
and U16348 (N_16348,N_12663,N_13957);
or U16349 (N_16349,N_12912,N_12940);
nand U16350 (N_16350,N_14858,N_12749);
and U16351 (N_16351,N_12907,N_14296);
xnor U16352 (N_16352,N_13266,N_13486);
xor U16353 (N_16353,N_14084,N_12938);
nor U16354 (N_16354,N_12653,N_13550);
or U16355 (N_16355,N_12632,N_14093);
xor U16356 (N_16356,N_13044,N_14777);
xor U16357 (N_16357,N_14671,N_14547);
or U16358 (N_16358,N_14682,N_14152);
xor U16359 (N_16359,N_14310,N_13296);
nor U16360 (N_16360,N_12841,N_13733);
and U16361 (N_16361,N_14116,N_14823);
nand U16362 (N_16362,N_12712,N_14152);
and U16363 (N_16363,N_14125,N_14025);
and U16364 (N_16364,N_12805,N_14110);
xor U16365 (N_16365,N_13969,N_14149);
and U16366 (N_16366,N_14172,N_14836);
or U16367 (N_16367,N_13391,N_14341);
and U16368 (N_16368,N_14894,N_14156);
or U16369 (N_16369,N_13904,N_13147);
nand U16370 (N_16370,N_13274,N_13259);
xnor U16371 (N_16371,N_14884,N_13077);
nand U16372 (N_16372,N_14371,N_14783);
or U16373 (N_16373,N_14423,N_13599);
xor U16374 (N_16374,N_12807,N_13122);
xor U16375 (N_16375,N_12821,N_13139);
nand U16376 (N_16376,N_13199,N_13195);
xnor U16377 (N_16377,N_14924,N_13552);
or U16378 (N_16378,N_13322,N_12856);
or U16379 (N_16379,N_13532,N_13289);
and U16380 (N_16380,N_14472,N_12980);
nand U16381 (N_16381,N_14385,N_14633);
xnor U16382 (N_16382,N_12915,N_13758);
xor U16383 (N_16383,N_12509,N_14244);
xor U16384 (N_16384,N_14703,N_12723);
xnor U16385 (N_16385,N_14834,N_13826);
nor U16386 (N_16386,N_14681,N_12560);
nand U16387 (N_16387,N_12767,N_14768);
or U16388 (N_16388,N_13775,N_13385);
and U16389 (N_16389,N_14970,N_13137);
and U16390 (N_16390,N_14844,N_14007);
and U16391 (N_16391,N_13228,N_14522);
nand U16392 (N_16392,N_12500,N_14376);
nand U16393 (N_16393,N_14445,N_14632);
or U16394 (N_16394,N_14631,N_13077);
xor U16395 (N_16395,N_12829,N_13006);
nand U16396 (N_16396,N_13631,N_14691);
xor U16397 (N_16397,N_13390,N_14602);
nand U16398 (N_16398,N_12619,N_14739);
xnor U16399 (N_16399,N_13054,N_14220);
and U16400 (N_16400,N_14830,N_13932);
nor U16401 (N_16401,N_12836,N_14827);
and U16402 (N_16402,N_12642,N_14932);
xnor U16403 (N_16403,N_14555,N_13025);
or U16404 (N_16404,N_13164,N_13377);
and U16405 (N_16405,N_14468,N_14362);
nor U16406 (N_16406,N_14208,N_13177);
nand U16407 (N_16407,N_13110,N_14976);
and U16408 (N_16408,N_13939,N_13567);
xor U16409 (N_16409,N_14558,N_14804);
nand U16410 (N_16410,N_12794,N_14706);
xnor U16411 (N_16411,N_12667,N_14174);
and U16412 (N_16412,N_13201,N_13620);
nor U16413 (N_16413,N_13191,N_14594);
and U16414 (N_16414,N_14984,N_14631);
and U16415 (N_16415,N_13504,N_13335);
xnor U16416 (N_16416,N_13263,N_14751);
and U16417 (N_16417,N_13653,N_13722);
xnor U16418 (N_16418,N_12699,N_13485);
or U16419 (N_16419,N_13817,N_13758);
or U16420 (N_16420,N_13019,N_12763);
nand U16421 (N_16421,N_13384,N_14464);
or U16422 (N_16422,N_14787,N_12877);
xor U16423 (N_16423,N_12702,N_14121);
nor U16424 (N_16424,N_14443,N_14683);
and U16425 (N_16425,N_14301,N_12500);
and U16426 (N_16426,N_13911,N_12618);
and U16427 (N_16427,N_14301,N_13699);
and U16428 (N_16428,N_14607,N_14552);
nor U16429 (N_16429,N_14644,N_14207);
nor U16430 (N_16430,N_12680,N_14457);
or U16431 (N_16431,N_14020,N_12952);
and U16432 (N_16432,N_13213,N_13281);
nor U16433 (N_16433,N_13552,N_14714);
xnor U16434 (N_16434,N_13464,N_13970);
nor U16435 (N_16435,N_12991,N_12621);
nand U16436 (N_16436,N_14204,N_14454);
nor U16437 (N_16437,N_14642,N_13252);
nand U16438 (N_16438,N_14350,N_14194);
xnor U16439 (N_16439,N_14858,N_14814);
xor U16440 (N_16440,N_13117,N_12748);
xnor U16441 (N_16441,N_14219,N_14714);
nand U16442 (N_16442,N_13701,N_14042);
or U16443 (N_16443,N_14844,N_12526);
nor U16444 (N_16444,N_14481,N_14327);
nor U16445 (N_16445,N_13926,N_14444);
xnor U16446 (N_16446,N_13142,N_13299);
nand U16447 (N_16447,N_14635,N_13642);
and U16448 (N_16448,N_14271,N_14061);
xor U16449 (N_16449,N_14461,N_12629);
and U16450 (N_16450,N_14872,N_13213);
and U16451 (N_16451,N_13242,N_14585);
and U16452 (N_16452,N_14933,N_14396);
and U16453 (N_16453,N_14550,N_13262);
nand U16454 (N_16454,N_13724,N_13190);
nor U16455 (N_16455,N_14205,N_13015);
nand U16456 (N_16456,N_13188,N_14295);
or U16457 (N_16457,N_12698,N_12509);
and U16458 (N_16458,N_12860,N_13693);
nor U16459 (N_16459,N_14639,N_12832);
xor U16460 (N_16460,N_14754,N_12580);
xnor U16461 (N_16461,N_14517,N_13356);
nand U16462 (N_16462,N_14325,N_14621);
xnor U16463 (N_16463,N_12689,N_13195);
and U16464 (N_16464,N_13217,N_14657);
nand U16465 (N_16465,N_13846,N_14947);
or U16466 (N_16466,N_14268,N_13189);
and U16467 (N_16467,N_13186,N_13624);
and U16468 (N_16468,N_14914,N_14103);
xor U16469 (N_16469,N_13858,N_14373);
or U16470 (N_16470,N_13958,N_13503);
and U16471 (N_16471,N_13448,N_13943);
xor U16472 (N_16472,N_14357,N_14020);
nor U16473 (N_16473,N_13039,N_14854);
nor U16474 (N_16474,N_12731,N_14596);
nand U16475 (N_16475,N_14530,N_14468);
xnor U16476 (N_16476,N_13905,N_14023);
nand U16477 (N_16477,N_13306,N_14956);
and U16478 (N_16478,N_14363,N_13141);
nand U16479 (N_16479,N_12629,N_12604);
and U16480 (N_16480,N_14184,N_13926);
and U16481 (N_16481,N_14937,N_13523);
or U16482 (N_16482,N_12832,N_14764);
nand U16483 (N_16483,N_12728,N_14269);
xnor U16484 (N_16484,N_13222,N_14783);
nor U16485 (N_16485,N_14857,N_14569);
and U16486 (N_16486,N_12704,N_12840);
nor U16487 (N_16487,N_14806,N_13805);
xnor U16488 (N_16488,N_14563,N_12535);
nand U16489 (N_16489,N_13418,N_13294);
or U16490 (N_16490,N_14327,N_13303);
xnor U16491 (N_16491,N_13409,N_14169);
or U16492 (N_16492,N_13144,N_13930);
or U16493 (N_16493,N_14735,N_13607);
and U16494 (N_16494,N_12849,N_14805);
nor U16495 (N_16495,N_13485,N_14989);
nor U16496 (N_16496,N_12575,N_12607);
nor U16497 (N_16497,N_13142,N_14402);
and U16498 (N_16498,N_13886,N_13707);
nor U16499 (N_16499,N_13898,N_14366);
xnor U16500 (N_16500,N_13525,N_13672);
nor U16501 (N_16501,N_12971,N_14110);
or U16502 (N_16502,N_13481,N_14280);
and U16503 (N_16503,N_13053,N_12670);
or U16504 (N_16504,N_14573,N_14408);
nand U16505 (N_16505,N_13487,N_12966);
xnor U16506 (N_16506,N_14754,N_14412);
nor U16507 (N_16507,N_12892,N_13087);
nor U16508 (N_16508,N_14290,N_14229);
nand U16509 (N_16509,N_12639,N_14371);
and U16510 (N_16510,N_13995,N_13407);
nand U16511 (N_16511,N_12990,N_13396);
or U16512 (N_16512,N_14581,N_13227);
or U16513 (N_16513,N_13720,N_14434);
and U16514 (N_16514,N_14405,N_13802);
or U16515 (N_16515,N_12699,N_13927);
nand U16516 (N_16516,N_14357,N_14893);
or U16517 (N_16517,N_13008,N_13885);
nand U16518 (N_16518,N_14336,N_12806);
nor U16519 (N_16519,N_14686,N_13480);
nor U16520 (N_16520,N_13034,N_14154);
nand U16521 (N_16521,N_13460,N_13255);
nor U16522 (N_16522,N_13296,N_13051);
nor U16523 (N_16523,N_14706,N_14718);
xnor U16524 (N_16524,N_14318,N_14569);
nor U16525 (N_16525,N_13963,N_12626);
xor U16526 (N_16526,N_13823,N_12908);
xor U16527 (N_16527,N_14747,N_12764);
or U16528 (N_16528,N_14026,N_13445);
nand U16529 (N_16529,N_13726,N_14926);
or U16530 (N_16530,N_13091,N_13787);
or U16531 (N_16531,N_14137,N_12971);
or U16532 (N_16532,N_13967,N_14261);
or U16533 (N_16533,N_12504,N_14800);
and U16534 (N_16534,N_13107,N_12749);
and U16535 (N_16535,N_14675,N_13317);
and U16536 (N_16536,N_13973,N_14049);
xor U16537 (N_16537,N_14941,N_12676);
nor U16538 (N_16538,N_13562,N_14258);
xnor U16539 (N_16539,N_13622,N_14632);
nor U16540 (N_16540,N_14713,N_14870);
nor U16541 (N_16541,N_13259,N_13578);
xor U16542 (N_16542,N_12835,N_13432);
or U16543 (N_16543,N_14261,N_13387);
or U16544 (N_16544,N_13408,N_12840);
nand U16545 (N_16545,N_14772,N_13993);
xor U16546 (N_16546,N_14404,N_14065);
nor U16547 (N_16547,N_13590,N_12566);
or U16548 (N_16548,N_14785,N_13937);
nand U16549 (N_16549,N_13124,N_13638);
xor U16550 (N_16550,N_14734,N_13398);
nor U16551 (N_16551,N_13371,N_13134);
nand U16552 (N_16552,N_12818,N_14306);
xor U16553 (N_16553,N_13569,N_14681);
and U16554 (N_16554,N_13368,N_12710);
nand U16555 (N_16555,N_13559,N_14032);
nand U16556 (N_16556,N_14477,N_14242);
or U16557 (N_16557,N_12984,N_14491);
or U16558 (N_16558,N_13957,N_13547);
nor U16559 (N_16559,N_13012,N_14582);
nand U16560 (N_16560,N_14569,N_13883);
nor U16561 (N_16561,N_12729,N_13496);
or U16562 (N_16562,N_14603,N_14086);
nand U16563 (N_16563,N_13786,N_13619);
xnor U16564 (N_16564,N_13828,N_14072);
and U16565 (N_16565,N_14613,N_14391);
and U16566 (N_16566,N_13479,N_14569);
or U16567 (N_16567,N_14605,N_13118);
nor U16568 (N_16568,N_13877,N_13213);
nor U16569 (N_16569,N_12507,N_14588);
nor U16570 (N_16570,N_13468,N_14013);
and U16571 (N_16571,N_13403,N_12505);
nor U16572 (N_16572,N_14380,N_14168);
and U16573 (N_16573,N_14734,N_14434);
nand U16574 (N_16574,N_14687,N_14522);
or U16575 (N_16575,N_14107,N_14945);
nand U16576 (N_16576,N_14921,N_12802);
and U16577 (N_16577,N_13966,N_14274);
or U16578 (N_16578,N_13525,N_14975);
xor U16579 (N_16579,N_14238,N_13428);
nand U16580 (N_16580,N_14125,N_12786);
nor U16581 (N_16581,N_14583,N_12895);
nor U16582 (N_16582,N_12513,N_12644);
or U16583 (N_16583,N_14669,N_13673);
nand U16584 (N_16584,N_14410,N_13933);
and U16585 (N_16585,N_13084,N_14519);
and U16586 (N_16586,N_13858,N_14394);
and U16587 (N_16587,N_12874,N_13873);
and U16588 (N_16588,N_13060,N_13406);
and U16589 (N_16589,N_13271,N_14433);
or U16590 (N_16590,N_14763,N_13204);
nor U16591 (N_16591,N_14524,N_14447);
and U16592 (N_16592,N_14346,N_12767);
nand U16593 (N_16593,N_14522,N_14021);
xor U16594 (N_16594,N_14914,N_13304);
nand U16595 (N_16595,N_13511,N_14122);
nor U16596 (N_16596,N_13030,N_13958);
and U16597 (N_16597,N_13058,N_14797);
xor U16598 (N_16598,N_14015,N_14936);
nand U16599 (N_16599,N_12547,N_14854);
nand U16600 (N_16600,N_13280,N_14661);
and U16601 (N_16601,N_13523,N_13636);
xnor U16602 (N_16602,N_14548,N_14883);
xor U16603 (N_16603,N_14819,N_12595);
nand U16604 (N_16604,N_13099,N_12978);
and U16605 (N_16605,N_13852,N_13274);
and U16606 (N_16606,N_14877,N_13079);
xor U16607 (N_16607,N_12995,N_12763);
nor U16608 (N_16608,N_14754,N_13741);
nor U16609 (N_16609,N_13341,N_13169);
xor U16610 (N_16610,N_14891,N_14569);
nand U16611 (N_16611,N_13145,N_12644);
or U16612 (N_16612,N_13438,N_14394);
xnor U16613 (N_16613,N_14305,N_13807);
or U16614 (N_16614,N_14405,N_12937);
and U16615 (N_16615,N_14410,N_14290);
or U16616 (N_16616,N_12913,N_14563);
nand U16617 (N_16617,N_13689,N_14541);
nor U16618 (N_16618,N_13634,N_13281);
nor U16619 (N_16619,N_14526,N_14672);
nand U16620 (N_16620,N_12506,N_13130);
or U16621 (N_16621,N_13224,N_14886);
xor U16622 (N_16622,N_13998,N_13450);
xor U16623 (N_16623,N_13201,N_13005);
xor U16624 (N_16624,N_14132,N_14909);
xor U16625 (N_16625,N_14454,N_14245);
nor U16626 (N_16626,N_13922,N_13789);
nor U16627 (N_16627,N_12673,N_13980);
or U16628 (N_16628,N_13679,N_12895);
xnor U16629 (N_16629,N_13956,N_13351);
nand U16630 (N_16630,N_13701,N_14701);
and U16631 (N_16631,N_12852,N_13127);
xnor U16632 (N_16632,N_12764,N_13568);
or U16633 (N_16633,N_13802,N_13315);
xor U16634 (N_16634,N_14181,N_12945);
xor U16635 (N_16635,N_12502,N_12717);
or U16636 (N_16636,N_14074,N_14814);
nand U16637 (N_16637,N_13275,N_13956);
xor U16638 (N_16638,N_13038,N_14501);
xor U16639 (N_16639,N_13458,N_13990);
and U16640 (N_16640,N_14849,N_13855);
or U16641 (N_16641,N_13396,N_14919);
nand U16642 (N_16642,N_14190,N_13699);
or U16643 (N_16643,N_13615,N_14416);
or U16644 (N_16644,N_13124,N_12886);
and U16645 (N_16645,N_14293,N_12848);
nor U16646 (N_16646,N_13000,N_12928);
nand U16647 (N_16647,N_12677,N_12647);
and U16648 (N_16648,N_13892,N_13715);
xor U16649 (N_16649,N_14566,N_12579);
nand U16650 (N_16650,N_13028,N_13160);
and U16651 (N_16651,N_14451,N_14470);
xor U16652 (N_16652,N_13391,N_13558);
xor U16653 (N_16653,N_12797,N_13796);
or U16654 (N_16654,N_13451,N_13109);
nand U16655 (N_16655,N_14435,N_13071);
and U16656 (N_16656,N_13184,N_12564);
xnor U16657 (N_16657,N_13188,N_13140);
and U16658 (N_16658,N_13261,N_13231);
nor U16659 (N_16659,N_13683,N_14719);
xnor U16660 (N_16660,N_13516,N_13394);
and U16661 (N_16661,N_12794,N_13144);
and U16662 (N_16662,N_14920,N_14331);
nand U16663 (N_16663,N_13832,N_12509);
and U16664 (N_16664,N_13941,N_14764);
nand U16665 (N_16665,N_14471,N_12933);
nand U16666 (N_16666,N_14282,N_14240);
and U16667 (N_16667,N_12604,N_13462);
and U16668 (N_16668,N_13963,N_12646);
nor U16669 (N_16669,N_14314,N_14662);
or U16670 (N_16670,N_13182,N_12938);
xnor U16671 (N_16671,N_14468,N_13859);
nor U16672 (N_16672,N_14086,N_13912);
nor U16673 (N_16673,N_13400,N_13748);
nor U16674 (N_16674,N_14481,N_14495);
nor U16675 (N_16675,N_13601,N_13890);
or U16676 (N_16676,N_12742,N_12828);
xor U16677 (N_16677,N_12821,N_13812);
or U16678 (N_16678,N_13366,N_13500);
xnor U16679 (N_16679,N_13229,N_13587);
nand U16680 (N_16680,N_14462,N_13324);
nand U16681 (N_16681,N_13493,N_13844);
and U16682 (N_16682,N_14955,N_14578);
nand U16683 (N_16683,N_14769,N_13069);
and U16684 (N_16684,N_13193,N_13060);
xnor U16685 (N_16685,N_13303,N_13347);
or U16686 (N_16686,N_12526,N_12922);
nor U16687 (N_16687,N_14392,N_14336);
or U16688 (N_16688,N_14156,N_12929);
nand U16689 (N_16689,N_14561,N_13022);
or U16690 (N_16690,N_13950,N_13816);
or U16691 (N_16691,N_13704,N_14593);
and U16692 (N_16692,N_12737,N_13937);
nand U16693 (N_16693,N_12502,N_14267);
nand U16694 (N_16694,N_12553,N_12599);
nor U16695 (N_16695,N_14072,N_14243);
xnor U16696 (N_16696,N_13544,N_14045);
or U16697 (N_16697,N_12814,N_12528);
nand U16698 (N_16698,N_14733,N_13224);
nand U16699 (N_16699,N_13827,N_13141);
xnor U16700 (N_16700,N_12873,N_14847);
nor U16701 (N_16701,N_12768,N_13987);
or U16702 (N_16702,N_12683,N_12763);
or U16703 (N_16703,N_13525,N_14537);
nor U16704 (N_16704,N_13116,N_12582);
and U16705 (N_16705,N_14945,N_13843);
and U16706 (N_16706,N_14518,N_14980);
and U16707 (N_16707,N_13244,N_13524);
and U16708 (N_16708,N_14752,N_13212);
nand U16709 (N_16709,N_14766,N_14209);
xor U16710 (N_16710,N_12774,N_13465);
and U16711 (N_16711,N_12970,N_14234);
xnor U16712 (N_16712,N_12857,N_13316);
xnor U16713 (N_16713,N_13623,N_14692);
nand U16714 (N_16714,N_14755,N_14052);
nand U16715 (N_16715,N_14688,N_13107);
and U16716 (N_16716,N_13496,N_14191);
or U16717 (N_16717,N_13908,N_13962);
xnor U16718 (N_16718,N_12866,N_13797);
nand U16719 (N_16719,N_13525,N_13548);
nor U16720 (N_16720,N_14213,N_13063);
xor U16721 (N_16721,N_13054,N_13275);
nand U16722 (N_16722,N_14733,N_12805);
nor U16723 (N_16723,N_14571,N_13062);
or U16724 (N_16724,N_14220,N_14601);
nor U16725 (N_16725,N_14755,N_13188);
nand U16726 (N_16726,N_12808,N_13858);
or U16727 (N_16727,N_13608,N_13264);
xnor U16728 (N_16728,N_14649,N_13917);
nor U16729 (N_16729,N_13570,N_14803);
nor U16730 (N_16730,N_13754,N_13789);
and U16731 (N_16731,N_13157,N_14982);
xnor U16732 (N_16732,N_13035,N_14917);
or U16733 (N_16733,N_12663,N_12947);
nand U16734 (N_16734,N_13210,N_13246);
xor U16735 (N_16735,N_14026,N_14569);
nor U16736 (N_16736,N_14107,N_12560);
xor U16737 (N_16737,N_12516,N_13973);
nor U16738 (N_16738,N_12752,N_14042);
xor U16739 (N_16739,N_14069,N_13941);
xor U16740 (N_16740,N_14555,N_12999);
or U16741 (N_16741,N_14354,N_13900);
nor U16742 (N_16742,N_14059,N_14758);
or U16743 (N_16743,N_14815,N_14312);
or U16744 (N_16744,N_14083,N_14602);
xor U16745 (N_16745,N_13854,N_14850);
or U16746 (N_16746,N_13780,N_12525);
or U16747 (N_16747,N_14653,N_12996);
nand U16748 (N_16748,N_14280,N_13831);
nand U16749 (N_16749,N_14719,N_14464);
and U16750 (N_16750,N_14297,N_14986);
nor U16751 (N_16751,N_13270,N_12976);
and U16752 (N_16752,N_13552,N_14026);
and U16753 (N_16753,N_14009,N_14364);
nor U16754 (N_16754,N_14028,N_13433);
nand U16755 (N_16755,N_12838,N_13027);
or U16756 (N_16756,N_13022,N_13835);
xor U16757 (N_16757,N_14193,N_12937);
nand U16758 (N_16758,N_14361,N_14188);
nor U16759 (N_16759,N_14265,N_12654);
or U16760 (N_16760,N_12774,N_12714);
and U16761 (N_16761,N_13823,N_13861);
and U16762 (N_16762,N_13179,N_14186);
xnor U16763 (N_16763,N_13566,N_14722);
nor U16764 (N_16764,N_14282,N_12790);
xor U16765 (N_16765,N_13341,N_14921);
nor U16766 (N_16766,N_14381,N_14242);
nand U16767 (N_16767,N_13064,N_12946);
or U16768 (N_16768,N_14863,N_13359);
or U16769 (N_16769,N_14584,N_13197);
nor U16770 (N_16770,N_14273,N_12848);
xnor U16771 (N_16771,N_13814,N_13653);
or U16772 (N_16772,N_13260,N_13429);
or U16773 (N_16773,N_13868,N_12524);
nand U16774 (N_16774,N_14360,N_13018);
nor U16775 (N_16775,N_12681,N_13814);
or U16776 (N_16776,N_13002,N_12869);
nor U16777 (N_16777,N_13502,N_13577);
nand U16778 (N_16778,N_13599,N_13046);
nor U16779 (N_16779,N_13958,N_14603);
xnor U16780 (N_16780,N_13197,N_14432);
nor U16781 (N_16781,N_12945,N_12555);
xnor U16782 (N_16782,N_14606,N_13902);
nand U16783 (N_16783,N_13481,N_14224);
xor U16784 (N_16784,N_14626,N_13375);
or U16785 (N_16785,N_14387,N_12710);
nor U16786 (N_16786,N_14020,N_13706);
xor U16787 (N_16787,N_13255,N_14711);
and U16788 (N_16788,N_13491,N_12907);
or U16789 (N_16789,N_13203,N_14699);
and U16790 (N_16790,N_12938,N_13624);
nor U16791 (N_16791,N_12811,N_13525);
and U16792 (N_16792,N_13860,N_14956);
xor U16793 (N_16793,N_14525,N_12641);
nor U16794 (N_16794,N_14837,N_14565);
nor U16795 (N_16795,N_14203,N_13679);
nand U16796 (N_16796,N_14240,N_14921);
or U16797 (N_16797,N_13062,N_14154);
or U16798 (N_16798,N_14103,N_12857);
or U16799 (N_16799,N_13553,N_12760);
and U16800 (N_16800,N_13064,N_14808);
and U16801 (N_16801,N_14203,N_14437);
or U16802 (N_16802,N_13215,N_12668);
and U16803 (N_16803,N_14915,N_13908);
xnor U16804 (N_16804,N_14526,N_13771);
and U16805 (N_16805,N_14733,N_14112);
and U16806 (N_16806,N_13405,N_13501);
and U16807 (N_16807,N_13092,N_12545);
nand U16808 (N_16808,N_12803,N_13491);
xnor U16809 (N_16809,N_14038,N_14492);
xor U16810 (N_16810,N_14648,N_13355);
and U16811 (N_16811,N_13702,N_12608);
xor U16812 (N_16812,N_13371,N_14811);
nor U16813 (N_16813,N_14192,N_13750);
nand U16814 (N_16814,N_14331,N_13354);
and U16815 (N_16815,N_14538,N_12840);
and U16816 (N_16816,N_13328,N_14483);
xor U16817 (N_16817,N_13893,N_12970);
nand U16818 (N_16818,N_13810,N_14736);
nor U16819 (N_16819,N_14846,N_14775);
and U16820 (N_16820,N_13111,N_14077);
or U16821 (N_16821,N_13450,N_13218);
or U16822 (N_16822,N_13396,N_13250);
and U16823 (N_16823,N_13689,N_12542);
xor U16824 (N_16824,N_12527,N_14695);
xnor U16825 (N_16825,N_13133,N_13839);
nor U16826 (N_16826,N_12770,N_12861);
nand U16827 (N_16827,N_14903,N_13164);
nand U16828 (N_16828,N_14277,N_14687);
or U16829 (N_16829,N_13313,N_14124);
and U16830 (N_16830,N_12792,N_13918);
or U16831 (N_16831,N_13154,N_13167);
or U16832 (N_16832,N_14424,N_14578);
nor U16833 (N_16833,N_14834,N_13677);
or U16834 (N_16834,N_13278,N_13669);
and U16835 (N_16835,N_13659,N_12873);
xnor U16836 (N_16836,N_12890,N_14992);
nor U16837 (N_16837,N_14731,N_14047);
xnor U16838 (N_16838,N_13846,N_13956);
xnor U16839 (N_16839,N_12715,N_13429);
and U16840 (N_16840,N_12772,N_13024);
nand U16841 (N_16841,N_13008,N_12905);
xnor U16842 (N_16842,N_14786,N_13632);
nor U16843 (N_16843,N_13349,N_13556);
or U16844 (N_16844,N_13029,N_13450);
and U16845 (N_16845,N_13798,N_13027);
and U16846 (N_16846,N_13250,N_14287);
or U16847 (N_16847,N_13602,N_14642);
or U16848 (N_16848,N_14483,N_14881);
nor U16849 (N_16849,N_12513,N_13125);
or U16850 (N_16850,N_14968,N_14990);
xor U16851 (N_16851,N_14780,N_12867);
and U16852 (N_16852,N_12686,N_13634);
xnor U16853 (N_16853,N_14066,N_13595);
xnor U16854 (N_16854,N_13186,N_14006);
nand U16855 (N_16855,N_14855,N_13660);
or U16856 (N_16856,N_13511,N_13340);
nand U16857 (N_16857,N_14985,N_12967);
xnor U16858 (N_16858,N_13462,N_14320);
xnor U16859 (N_16859,N_13604,N_12597);
or U16860 (N_16860,N_14907,N_14105);
nor U16861 (N_16861,N_14689,N_13784);
and U16862 (N_16862,N_14188,N_12763);
or U16863 (N_16863,N_14770,N_14360);
xor U16864 (N_16864,N_14459,N_13390);
and U16865 (N_16865,N_12965,N_12788);
nor U16866 (N_16866,N_14270,N_12846);
nand U16867 (N_16867,N_13802,N_13478);
xnor U16868 (N_16868,N_14364,N_14281);
or U16869 (N_16869,N_13030,N_13752);
and U16870 (N_16870,N_13175,N_14561);
nand U16871 (N_16871,N_14700,N_14732);
and U16872 (N_16872,N_13583,N_12587);
or U16873 (N_16873,N_13176,N_14353);
nand U16874 (N_16874,N_13556,N_13539);
nand U16875 (N_16875,N_12805,N_14351);
xnor U16876 (N_16876,N_13993,N_14368);
nand U16877 (N_16877,N_14507,N_14844);
or U16878 (N_16878,N_14117,N_13055);
and U16879 (N_16879,N_13329,N_14958);
xor U16880 (N_16880,N_14129,N_13353);
or U16881 (N_16881,N_14580,N_14763);
xor U16882 (N_16882,N_13042,N_14850);
xor U16883 (N_16883,N_12757,N_14684);
xnor U16884 (N_16884,N_14131,N_14106);
xor U16885 (N_16885,N_12834,N_14766);
nor U16886 (N_16886,N_12571,N_14284);
xnor U16887 (N_16887,N_14559,N_13798);
or U16888 (N_16888,N_13326,N_12500);
and U16889 (N_16889,N_14608,N_14877);
and U16890 (N_16890,N_13214,N_14278);
or U16891 (N_16891,N_14329,N_14890);
xnor U16892 (N_16892,N_14586,N_14295);
and U16893 (N_16893,N_14201,N_12961);
nand U16894 (N_16894,N_14410,N_12859);
or U16895 (N_16895,N_14293,N_13506);
or U16896 (N_16896,N_13506,N_13309);
nor U16897 (N_16897,N_13503,N_12759);
and U16898 (N_16898,N_13629,N_12805);
xnor U16899 (N_16899,N_14548,N_14976);
or U16900 (N_16900,N_14788,N_14878);
nand U16901 (N_16901,N_13136,N_13377);
nor U16902 (N_16902,N_14637,N_13757);
and U16903 (N_16903,N_13600,N_12531);
xnor U16904 (N_16904,N_12863,N_13399);
or U16905 (N_16905,N_14261,N_14047);
xnor U16906 (N_16906,N_12760,N_14192);
xnor U16907 (N_16907,N_13510,N_13250);
nor U16908 (N_16908,N_12956,N_12554);
nand U16909 (N_16909,N_13914,N_13897);
nand U16910 (N_16910,N_12672,N_13732);
or U16911 (N_16911,N_14760,N_13239);
nor U16912 (N_16912,N_12563,N_14171);
or U16913 (N_16913,N_13073,N_14065);
or U16914 (N_16914,N_13924,N_13721);
xnor U16915 (N_16915,N_14103,N_12902);
nand U16916 (N_16916,N_14680,N_13632);
nand U16917 (N_16917,N_14928,N_14205);
nand U16918 (N_16918,N_13307,N_13698);
nor U16919 (N_16919,N_13351,N_14759);
nor U16920 (N_16920,N_12960,N_13868);
xnor U16921 (N_16921,N_14147,N_14079);
and U16922 (N_16922,N_12618,N_13932);
and U16923 (N_16923,N_12678,N_13155);
or U16924 (N_16924,N_12838,N_14113);
nand U16925 (N_16925,N_14402,N_14655);
xor U16926 (N_16926,N_13180,N_13775);
nor U16927 (N_16927,N_12758,N_14895);
or U16928 (N_16928,N_12967,N_13350);
xor U16929 (N_16929,N_12940,N_14071);
nand U16930 (N_16930,N_14116,N_13027);
and U16931 (N_16931,N_14260,N_14700);
nand U16932 (N_16932,N_14466,N_13740);
xor U16933 (N_16933,N_13783,N_14055);
and U16934 (N_16934,N_14098,N_14905);
or U16935 (N_16935,N_13316,N_13329);
xor U16936 (N_16936,N_13006,N_14697);
and U16937 (N_16937,N_14623,N_12837);
xor U16938 (N_16938,N_13981,N_13648);
and U16939 (N_16939,N_14190,N_12921);
nor U16940 (N_16940,N_14831,N_13584);
nor U16941 (N_16941,N_13090,N_14833);
and U16942 (N_16942,N_14471,N_12579);
xnor U16943 (N_16943,N_14942,N_13903);
nand U16944 (N_16944,N_14743,N_14913);
nor U16945 (N_16945,N_12879,N_13144);
and U16946 (N_16946,N_14054,N_14310);
nor U16947 (N_16947,N_13254,N_12923);
xnor U16948 (N_16948,N_12964,N_14182);
and U16949 (N_16949,N_13817,N_13787);
or U16950 (N_16950,N_12976,N_14692);
nand U16951 (N_16951,N_12505,N_14785);
nand U16952 (N_16952,N_13807,N_14763);
nand U16953 (N_16953,N_13093,N_13828);
or U16954 (N_16954,N_12858,N_12518);
nand U16955 (N_16955,N_14476,N_14990);
or U16956 (N_16956,N_14255,N_13357);
and U16957 (N_16957,N_13457,N_13026);
and U16958 (N_16958,N_14386,N_14748);
xor U16959 (N_16959,N_14420,N_14887);
and U16960 (N_16960,N_12916,N_13497);
xor U16961 (N_16961,N_13084,N_14218);
nor U16962 (N_16962,N_12927,N_14140);
and U16963 (N_16963,N_12761,N_14121);
nand U16964 (N_16964,N_13273,N_13322);
xnor U16965 (N_16965,N_14035,N_13506);
nor U16966 (N_16966,N_14517,N_13111);
nand U16967 (N_16967,N_14201,N_12677);
nor U16968 (N_16968,N_13172,N_14522);
nand U16969 (N_16969,N_13105,N_13757);
xnor U16970 (N_16970,N_14785,N_13254);
nor U16971 (N_16971,N_13536,N_14466);
xor U16972 (N_16972,N_14558,N_13100);
nand U16973 (N_16973,N_14262,N_13572);
xor U16974 (N_16974,N_14459,N_14772);
or U16975 (N_16975,N_14140,N_14205);
xnor U16976 (N_16976,N_14932,N_14786);
xor U16977 (N_16977,N_12661,N_12504);
xor U16978 (N_16978,N_14331,N_13356);
and U16979 (N_16979,N_12528,N_12704);
or U16980 (N_16980,N_12805,N_13745);
nand U16981 (N_16981,N_13962,N_14909);
or U16982 (N_16982,N_14904,N_14276);
nor U16983 (N_16983,N_12975,N_14787);
or U16984 (N_16984,N_12560,N_14131);
and U16985 (N_16985,N_13234,N_14985);
and U16986 (N_16986,N_13671,N_12944);
or U16987 (N_16987,N_12946,N_14556);
nor U16988 (N_16988,N_14662,N_14456);
nor U16989 (N_16989,N_12779,N_13367);
and U16990 (N_16990,N_13126,N_13550);
xnor U16991 (N_16991,N_13110,N_12947);
nand U16992 (N_16992,N_13890,N_13487);
xnor U16993 (N_16993,N_14810,N_13185);
nor U16994 (N_16994,N_14734,N_13830);
nand U16995 (N_16995,N_13698,N_14115);
nor U16996 (N_16996,N_12606,N_12730);
and U16997 (N_16997,N_14630,N_12527);
and U16998 (N_16998,N_13693,N_14173);
nor U16999 (N_16999,N_14544,N_14135);
nor U17000 (N_17000,N_14573,N_13213);
and U17001 (N_17001,N_13121,N_13033);
nor U17002 (N_17002,N_12904,N_14522);
or U17003 (N_17003,N_14166,N_12613);
nand U17004 (N_17004,N_13589,N_13738);
nor U17005 (N_17005,N_14146,N_13301);
nor U17006 (N_17006,N_12636,N_14723);
nand U17007 (N_17007,N_13354,N_14338);
or U17008 (N_17008,N_14021,N_14960);
nand U17009 (N_17009,N_13953,N_13892);
or U17010 (N_17010,N_13353,N_14475);
and U17011 (N_17011,N_13819,N_12812);
xnor U17012 (N_17012,N_13674,N_12737);
or U17013 (N_17013,N_14261,N_12794);
nand U17014 (N_17014,N_14048,N_13408);
nor U17015 (N_17015,N_14337,N_14817);
nand U17016 (N_17016,N_13721,N_13911);
and U17017 (N_17017,N_14000,N_12971);
nand U17018 (N_17018,N_13213,N_14246);
nand U17019 (N_17019,N_14910,N_14057);
or U17020 (N_17020,N_12592,N_14919);
and U17021 (N_17021,N_14006,N_14123);
nand U17022 (N_17022,N_14527,N_14114);
nand U17023 (N_17023,N_13958,N_13780);
nand U17024 (N_17024,N_13324,N_14459);
xnor U17025 (N_17025,N_14341,N_13981);
nor U17026 (N_17026,N_13055,N_13208);
nor U17027 (N_17027,N_13374,N_13967);
nand U17028 (N_17028,N_14016,N_14202);
and U17029 (N_17029,N_12838,N_14785);
nand U17030 (N_17030,N_13317,N_14543);
nand U17031 (N_17031,N_13265,N_14299);
nand U17032 (N_17032,N_14915,N_12569);
nor U17033 (N_17033,N_13602,N_13403);
nor U17034 (N_17034,N_12574,N_13867);
or U17035 (N_17035,N_13250,N_12675);
or U17036 (N_17036,N_13378,N_14457);
nand U17037 (N_17037,N_12571,N_13224);
nor U17038 (N_17038,N_13803,N_14998);
or U17039 (N_17039,N_13908,N_12821);
nand U17040 (N_17040,N_12848,N_13257);
xnor U17041 (N_17041,N_12872,N_13220);
and U17042 (N_17042,N_14198,N_12841);
xnor U17043 (N_17043,N_14925,N_13888);
or U17044 (N_17044,N_12640,N_13186);
or U17045 (N_17045,N_14534,N_13405);
or U17046 (N_17046,N_13371,N_13092);
xnor U17047 (N_17047,N_13638,N_12624);
xnor U17048 (N_17048,N_14847,N_14106);
or U17049 (N_17049,N_13676,N_12862);
xnor U17050 (N_17050,N_12714,N_13042);
and U17051 (N_17051,N_13214,N_13553);
and U17052 (N_17052,N_14721,N_14281);
nor U17053 (N_17053,N_13030,N_12727);
and U17054 (N_17054,N_13574,N_14213);
and U17055 (N_17055,N_14718,N_12965);
or U17056 (N_17056,N_14436,N_13784);
and U17057 (N_17057,N_13995,N_13336);
xnor U17058 (N_17058,N_13590,N_14292);
nand U17059 (N_17059,N_14725,N_13214);
and U17060 (N_17060,N_12789,N_13933);
xnor U17061 (N_17061,N_12970,N_14370);
nor U17062 (N_17062,N_13249,N_13194);
nand U17063 (N_17063,N_14859,N_12640);
nor U17064 (N_17064,N_14251,N_12982);
nor U17065 (N_17065,N_14615,N_13322);
xor U17066 (N_17066,N_13457,N_13480);
xnor U17067 (N_17067,N_13950,N_14704);
nor U17068 (N_17068,N_13868,N_14982);
xnor U17069 (N_17069,N_13022,N_12727);
nand U17070 (N_17070,N_14035,N_14794);
nand U17071 (N_17071,N_13481,N_14216);
and U17072 (N_17072,N_13928,N_14359);
nor U17073 (N_17073,N_13622,N_13872);
or U17074 (N_17074,N_14001,N_13994);
and U17075 (N_17075,N_14858,N_14512);
nand U17076 (N_17076,N_14945,N_13221);
or U17077 (N_17077,N_13848,N_12868);
xor U17078 (N_17078,N_14198,N_14123);
nand U17079 (N_17079,N_13528,N_13838);
xor U17080 (N_17080,N_14155,N_12946);
and U17081 (N_17081,N_13669,N_14845);
nand U17082 (N_17082,N_14097,N_13358);
and U17083 (N_17083,N_13597,N_14454);
nand U17084 (N_17084,N_13184,N_12664);
nor U17085 (N_17085,N_14700,N_13324);
nand U17086 (N_17086,N_13119,N_13650);
xor U17087 (N_17087,N_13793,N_12902);
and U17088 (N_17088,N_14220,N_14454);
xor U17089 (N_17089,N_14827,N_13801);
or U17090 (N_17090,N_14949,N_13329);
xnor U17091 (N_17091,N_14473,N_12818);
xor U17092 (N_17092,N_13050,N_12765);
and U17093 (N_17093,N_13968,N_13791);
nor U17094 (N_17094,N_12627,N_12818);
and U17095 (N_17095,N_14871,N_13544);
or U17096 (N_17096,N_13841,N_13737);
or U17097 (N_17097,N_13503,N_13376);
nand U17098 (N_17098,N_13914,N_13868);
xor U17099 (N_17099,N_14719,N_14834);
xnor U17100 (N_17100,N_13094,N_14455);
and U17101 (N_17101,N_13349,N_12784);
xnor U17102 (N_17102,N_13479,N_12745);
nor U17103 (N_17103,N_14425,N_14053);
and U17104 (N_17104,N_14490,N_13676);
nor U17105 (N_17105,N_12578,N_14784);
and U17106 (N_17106,N_13518,N_12891);
and U17107 (N_17107,N_13487,N_13684);
nand U17108 (N_17108,N_13487,N_13212);
nor U17109 (N_17109,N_14586,N_13416);
and U17110 (N_17110,N_13112,N_14165);
xnor U17111 (N_17111,N_13670,N_13131);
xor U17112 (N_17112,N_13684,N_13526);
nor U17113 (N_17113,N_14837,N_12514);
xnor U17114 (N_17114,N_13021,N_14982);
nor U17115 (N_17115,N_13675,N_12537);
nor U17116 (N_17116,N_13731,N_13687);
xnor U17117 (N_17117,N_14833,N_14964);
xor U17118 (N_17118,N_13207,N_14986);
or U17119 (N_17119,N_12625,N_14414);
nand U17120 (N_17120,N_14371,N_13387);
or U17121 (N_17121,N_13109,N_13750);
and U17122 (N_17122,N_14038,N_14130);
xnor U17123 (N_17123,N_13816,N_14593);
and U17124 (N_17124,N_14833,N_14163);
xor U17125 (N_17125,N_14511,N_14547);
and U17126 (N_17126,N_13387,N_14429);
and U17127 (N_17127,N_12788,N_12840);
or U17128 (N_17128,N_13854,N_12532);
and U17129 (N_17129,N_12791,N_13933);
or U17130 (N_17130,N_14063,N_14688);
nor U17131 (N_17131,N_12987,N_12595);
nor U17132 (N_17132,N_14181,N_13606);
or U17133 (N_17133,N_13688,N_12905);
nand U17134 (N_17134,N_14918,N_12585);
or U17135 (N_17135,N_12703,N_14689);
nor U17136 (N_17136,N_14957,N_13430);
nand U17137 (N_17137,N_13615,N_12794);
or U17138 (N_17138,N_12920,N_13625);
and U17139 (N_17139,N_12520,N_12629);
nand U17140 (N_17140,N_12947,N_13334);
or U17141 (N_17141,N_14314,N_14879);
nand U17142 (N_17142,N_13700,N_13124);
or U17143 (N_17143,N_14109,N_14438);
and U17144 (N_17144,N_13876,N_13279);
nand U17145 (N_17145,N_14797,N_13497);
nor U17146 (N_17146,N_14632,N_13900);
xnor U17147 (N_17147,N_14661,N_14166);
or U17148 (N_17148,N_13532,N_13723);
nor U17149 (N_17149,N_14837,N_14125);
nor U17150 (N_17150,N_14201,N_13819);
xnor U17151 (N_17151,N_14893,N_14859);
or U17152 (N_17152,N_13041,N_14226);
xor U17153 (N_17153,N_13290,N_13595);
or U17154 (N_17154,N_14012,N_13735);
or U17155 (N_17155,N_12827,N_14030);
and U17156 (N_17156,N_14554,N_13838);
xor U17157 (N_17157,N_14149,N_14505);
xnor U17158 (N_17158,N_13222,N_14491);
or U17159 (N_17159,N_14876,N_14890);
nand U17160 (N_17160,N_13446,N_14114);
or U17161 (N_17161,N_12593,N_12568);
or U17162 (N_17162,N_12856,N_14121);
xnor U17163 (N_17163,N_12663,N_14973);
nand U17164 (N_17164,N_12964,N_13447);
and U17165 (N_17165,N_13103,N_14960);
nor U17166 (N_17166,N_14049,N_13865);
nor U17167 (N_17167,N_14431,N_12992);
nand U17168 (N_17168,N_14211,N_14267);
nor U17169 (N_17169,N_13797,N_14823);
xor U17170 (N_17170,N_13370,N_14066);
or U17171 (N_17171,N_12919,N_12858);
and U17172 (N_17172,N_12704,N_12883);
xor U17173 (N_17173,N_14260,N_14946);
nand U17174 (N_17174,N_12738,N_14384);
and U17175 (N_17175,N_13142,N_14803);
and U17176 (N_17176,N_14847,N_13850);
or U17177 (N_17177,N_13018,N_13742);
nand U17178 (N_17178,N_13225,N_13337);
nand U17179 (N_17179,N_13889,N_13045);
nor U17180 (N_17180,N_12942,N_13652);
or U17181 (N_17181,N_13906,N_12598);
nand U17182 (N_17182,N_13452,N_13455);
or U17183 (N_17183,N_14773,N_14880);
xor U17184 (N_17184,N_13338,N_14207);
nor U17185 (N_17185,N_14640,N_12838);
nor U17186 (N_17186,N_14866,N_13726);
nor U17187 (N_17187,N_12967,N_13732);
nand U17188 (N_17188,N_13385,N_12937);
nor U17189 (N_17189,N_12737,N_14872);
nor U17190 (N_17190,N_13494,N_14537);
or U17191 (N_17191,N_14941,N_14189);
and U17192 (N_17192,N_12966,N_14692);
xnor U17193 (N_17193,N_14340,N_13052);
nor U17194 (N_17194,N_12512,N_13730);
and U17195 (N_17195,N_12732,N_14415);
or U17196 (N_17196,N_13643,N_14351);
or U17197 (N_17197,N_14945,N_12918);
nand U17198 (N_17198,N_13003,N_13566);
xor U17199 (N_17199,N_12687,N_14921);
nor U17200 (N_17200,N_13066,N_14685);
nor U17201 (N_17201,N_12744,N_13462);
or U17202 (N_17202,N_14570,N_14316);
and U17203 (N_17203,N_14568,N_13649);
nor U17204 (N_17204,N_14460,N_12594);
nor U17205 (N_17205,N_13342,N_13838);
or U17206 (N_17206,N_13363,N_12725);
nor U17207 (N_17207,N_13714,N_14097);
and U17208 (N_17208,N_13163,N_13482);
nand U17209 (N_17209,N_13275,N_14520);
nor U17210 (N_17210,N_12558,N_13520);
or U17211 (N_17211,N_13045,N_12945);
nor U17212 (N_17212,N_14767,N_14409);
and U17213 (N_17213,N_13710,N_14268);
xnor U17214 (N_17214,N_14622,N_12872);
or U17215 (N_17215,N_13324,N_12774);
xor U17216 (N_17216,N_14454,N_12998);
nand U17217 (N_17217,N_14704,N_13857);
or U17218 (N_17218,N_14735,N_12778);
or U17219 (N_17219,N_12714,N_13441);
nor U17220 (N_17220,N_13315,N_12597);
nand U17221 (N_17221,N_14436,N_13800);
nand U17222 (N_17222,N_14186,N_12582);
or U17223 (N_17223,N_13331,N_12780);
or U17224 (N_17224,N_13619,N_12664);
nor U17225 (N_17225,N_14742,N_12832);
and U17226 (N_17226,N_14319,N_14524);
xnor U17227 (N_17227,N_14244,N_12819);
xor U17228 (N_17228,N_13961,N_13585);
nor U17229 (N_17229,N_14380,N_14387);
and U17230 (N_17230,N_12643,N_14834);
xnor U17231 (N_17231,N_14794,N_13735);
xnor U17232 (N_17232,N_14001,N_13552);
or U17233 (N_17233,N_13309,N_12873);
or U17234 (N_17234,N_12546,N_14069);
and U17235 (N_17235,N_12545,N_13122);
and U17236 (N_17236,N_13662,N_12852);
nor U17237 (N_17237,N_12530,N_14732);
nor U17238 (N_17238,N_12600,N_14029);
nor U17239 (N_17239,N_13836,N_14091);
nand U17240 (N_17240,N_13082,N_12758);
nand U17241 (N_17241,N_13914,N_14051);
or U17242 (N_17242,N_14397,N_13706);
nor U17243 (N_17243,N_12799,N_13826);
nand U17244 (N_17244,N_12533,N_14862);
or U17245 (N_17245,N_13427,N_14672);
or U17246 (N_17246,N_12679,N_13983);
or U17247 (N_17247,N_12664,N_13987);
and U17248 (N_17248,N_13449,N_14455);
and U17249 (N_17249,N_13606,N_14946);
or U17250 (N_17250,N_14441,N_13432);
and U17251 (N_17251,N_13690,N_14247);
xnor U17252 (N_17252,N_13131,N_14383);
or U17253 (N_17253,N_13116,N_13516);
nand U17254 (N_17254,N_12674,N_13706);
nor U17255 (N_17255,N_14279,N_13930);
nand U17256 (N_17256,N_13412,N_12908);
nor U17257 (N_17257,N_14306,N_13233);
or U17258 (N_17258,N_12551,N_14621);
and U17259 (N_17259,N_14425,N_13895);
xor U17260 (N_17260,N_13208,N_13353);
nand U17261 (N_17261,N_12868,N_14254);
nor U17262 (N_17262,N_14850,N_12661);
and U17263 (N_17263,N_14337,N_13281);
xor U17264 (N_17264,N_14836,N_13609);
nor U17265 (N_17265,N_13565,N_14359);
or U17266 (N_17266,N_12824,N_14063);
or U17267 (N_17267,N_13556,N_13536);
or U17268 (N_17268,N_12817,N_13614);
or U17269 (N_17269,N_13279,N_14058);
nand U17270 (N_17270,N_13261,N_12818);
nor U17271 (N_17271,N_14916,N_14758);
nand U17272 (N_17272,N_13121,N_13321);
nor U17273 (N_17273,N_14628,N_13101);
nand U17274 (N_17274,N_13174,N_13417);
xnor U17275 (N_17275,N_14522,N_12902);
nand U17276 (N_17276,N_12866,N_13955);
nor U17277 (N_17277,N_13391,N_13576);
and U17278 (N_17278,N_13426,N_14920);
xor U17279 (N_17279,N_14734,N_14395);
xnor U17280 (N_17280,N_14902,N_14152);
nand U17281 (N_17281,N_14886,N_14484);
or U17282 (N_17282,N_14818,N_14384);
nand U17283 (N_17283,N_13055,N_14142);
nand U17284 (N_17284,N_14752,N_13628);
and U17285 (N_17285,N_13558,N_13062);
or U17286 (N_17286,N_14333,N_12750);
nor U17287 (N_17287,N_12528,N_14404);
nand U17288 (N_17288,N_12525,N_13290);
and U17289 (N_17289,N_12939,N_13704);
xnor U17290 (N_17290,N_12511,N_14846);
nor U17291 (N_17291,N_14512,N_14463);
nor U17292 (N_17292,N_13660,N_13252);
nand U17293 (N_17293,N_13824,N_13852);
nand U17294 (N_17294,N_14422,N_12835);
and U17295 (N_17295,N_12768,N_13446);
nor U17296 (N_17296,N_12877,N_13572);
nor U17297 (N_17297,N_12922,N_12670);
or U17298 (N_17298,N_14274,N_14649);
or U17299 (N_17299,N_13347,N_13365);
or U17300 (N_17300,N_12973,N_14458);
xnor U17301 (N_17301,N_13666,N_13188);
nor U17302 (N_17302,N_13683,N_14676);
and U17303 (N_17303,N_13223,N_13471);
or U17304 (N_17304,N_13281,N_14690);
or U17305 (N_17305,N_12899,N_13957);
nand U17306 (N_17306,N_13831,N_14029);
xnor U17307 (N_17307,N_13391,N_14253);
xnor U17308 (N_17308,N_14794,N_14885);
xor U17309 (N_17309,N_12564,N_12500);
and U17310 (N_17310,N_14127,N_13427);
nor U17311 (N_17311,N_13216,N_13807);
nand U17312 (N_17312,N_14182,N_12535);
xor U17313 (N_17313,N_13114,N_13081);
or U17314 (N_17314,N_13902,N_12860);
and U17315 (N_17315,N_13709,N_14211);
and U17316 (N_17316,N_14377,N_13858);
or U17317 (N_17317,N_14116,N_13691);
nor U17318 (N_17318,N_13776,N_13390);
and U17319 (N_17319,N_14641,N_12594);
nor U17320 (N_17320,N_13973,N_13145);
or U17321 (N_17321,N_13981,N_13569);
xnor U17322 (N_17322,N_14786,N_14105);
or U17323 (N_17323,N_14941,N_14324);
nand U17324 (N_17324,N_13672,N_12926);
nor U17325 (N_17325,N_14803,N_14456);
nor U17326 (N_17326,N_14781,N_14777);
nand U17327 (N_17327,N_14043,N_13135);
nand U17328 (N_17328,N_12736,N_14142);
nand U17329 (N_17329,N_12941,N_13572);
nor U17330 (N_17330,N_13269,N_12734);
nand U17331 (N_17331,N_14291,N_14234);
nand U17332 (N_17332,N_14745,N_13122);
nor U17333 (N_17333,N_14666,N_13976);
nand U17334 (N_17334,N_12711,N_14732);
and U17335 (N_17335,N_14108,N_14070);
nand U17336 (N_17336,N_13704,N_13176);
and U17337 (N_17337,N_13551,N_14273);
nand U17338 (N_17338,N_12779,N_12572);
xnor U17339 (N_17339,N_12931,N_14272);
and U17340 (N_17340,N_13061,N_14870);
xor U17341 (N_17341,N_13315,N_12575);
and U17342 (N_17342,N_14913,N_13617);
nor U17343 (N_17343,N_14047,N_14519);
nand U17344 (N_17344,N_14246,N_13720);
nor U17345 (N_17345,N_14730,N_12944);
nand U17346 (N_17346,N_12540,N_14795);
xnor U17347 (N_17347,N_12869,N_14664);
xor U17348 (N_17348,N_13917,N_13388);
and U17349 (N_17349,N_14153,N_14446);
and U17350 (N_17350,N_14067,N_12816);
nand U17351 (N_17351,N_13121,N_12665);
and U17352 (N_17352,N_12971,N_14870);
xor U17353 (N_17353,N_13850,N_12681);
nor U17354 (N_17354,N_12941,N_14942);
or U17355 (N_17355,N_13542,N_13021);
or U17356 (N_17356,N_13581,N_14905);
nand U17357 (N_17357,N_12923,N_14840);
and U17358 (N_17358,N_13159,N_14171);
or U17359 (N_17359,N_13598,N_14672);
or U17360 (N_17360,N_13568,N_14718);
nor U17361 (N_17361,N_12751,N_13850);
and U17362 (N_17362,N_12633,N_14530);
or U17363 (N_17363,N_13826,N_13173);
nor U17364 (N_17364,N_14676,N_13091);
nor U17365 (N_17365,N_13203,N_12804);
and U17366 (N_17366,N_14789,N_12576);
nor U17367 (N_17367,N_14895,N_14515);
xnor U17368 (N_17368,N_13812,N_13808);
xor U17369 (N_17369,N_13820,N_14734);
nand U17370 (N_17370,N_14068,N_13804);
xnor U17371 (N_17371,N_14289,N_12747);
nand U17372 (N_17372,N_14685,N_12649);
or U17373 (N_17373,N_13325,N_13910);
nand U17374 (N_17374,N_13576,N_12785);
nand U17375 (N_17375,N_13971,N_13403);
and U17376 (N_17376,N_13416,N_13528);
xor U17377 (N_17377,N_13149,N_13649);
xnor U17378 (N_17378,N_14908,N_14208);
xor U17379 (N_17379,N_14923,N_13241);
nand U17380 (N_17380,N_13687,N_14615);
nand U17381 (N_17381,N_13759,N_14851);
nor U17382 (N_17382,N_14492,N_12710);
or U17383 (N_17383,N_12766,N_12609);
or U17384 (N_17384,N_13862,N_13970);
nor U17385 (N_17385,N_14874,N_12892);
and U17386 (N_17386,N_14382,N_14155);
or U17387 (N_17387,N_12945,N_14493);
and U17388 (N_17388,N_12827,N_14151);
nand U17389 (N_17389,N_12835,N_13232);
nand U17390 (N_17390,N_12655,N_12584);
nor U17391 (N_17391,N_13305,N_14138);
nor U17392 (N_17392,N_13598,N_14320);
nand U17393 (N_17393,N_13622,N_13854);
and U17394 (N_17394,N_14081,N_14638);
nor U17395 (N_17395,N_14478,N_12945);
nand U17396 (N_17396,N_14805,N_13630);
and U17397 (N_17397,N_13108,N_12600);
nor U17398 (N_17398,N_13472,N_13688);
and U17399 (N_17399,N_13054,N_13673);
and U17400 (N_17400,N_12948,N_13629);
or U17401 (N_17401,N_14643,N_14862);
nand U17402 (N_17402,N_14097,N_14950);
xnor U17403 (N_17403,N_13459,N_12737);
xnor U17404 (N_17404,N_13119,N_14833);
nor U17405 (N_17405,N_14546,N_14673);
xnor U17406 (N_17406,N_13632,N_13388);
xnor U17407 (N_17407,N_14105,N_14352);
nand U17408 (N_17408,N_14833,N_13725);
and U17409 (N_17409,N_13138,N_14849);
xnor U17410 (N_17410,N_13087,N_12816);
nor U17411 (N_17411,N_14107,N_14110);
and U17412 (N_17412,N_14432,N_14624);
nand U17413 (N_17413,N_14458,N_12980);
nand U17414 (N_17414,N_12537,N_14262);
and U17415 (N_17415,N_13295,N_13778);
and U17416 (N_17416,N_13117,N_12728);
nand U17417 (N_17417,N_12909,N_14459);
or U17418 (N_17418,N_12569,N_14671);
nand U17419 (N_17419,N_13653,N_13695);
or U17420 (N_17420,N_14472,N_14441);
nand U17421 (N_17421,N_14508,N_14566);
nand U17422 (N_17422,N_14180,N_12816);
nand U17423 (N_17423,N_13489,N_13214);
nor U17424 (N_17424,N_13299,N_14006);
xnor U17425 (N_17425,N_13084,N_14295);
or U17426 (N_17426,N_13207,N_13540);
nand U17427 (N_17427,N_12676,N_13011);
or U17428 (N_17428,N_12731,N_12621);
xor U17429 (N_17429,N_13696,N_14842);
xnor U17430 (N_17430,N_13181,N_13183);
nor U17431 (N_17431,N_12751,N_14760);
xnor U17432 (N_17432,N_14761,N_13257);
nor U17433 (N_17433,N_13871,N_14381);
and U17434 (N_17434,N_12597,N_14511);
xnor U17435 (N_17435,N_12726,N_14760);
xnor U17436 (N_17436,N_13453,N_14480);
and U17437 (N_17437,N_12711,N_14807);
nor U17438 (N_17438,N_13939,N_14627);
nand U17439 (N_17439,N_12600,N_13457);
nor U17440 (N_17440,N_13954,N_12850);
and U17441 (N_17441,N_13907,N_14589);
xor U17442 (N_17442,N_13124,N_13625);
nand U17443 (N_17443,N_14563,N_14250);
or U17444 (N_17444,N_14028,N_14715);
nand U17445 (N_17445,N_13117,N_13992);
and U17446 (N_17446,N_14891,N_13810);
or U17447 (N_17447,N_14085,N_12834);
or U17448 (N_17448,N_14316,N_14874);
nor U17449 (N_17449,N_13733,N_13194);
nand U17450 (N_17450,N_14474,N_14144);
and U17451 (N_17451,N_13411,N_14564);
and U17452 (N_17452,N_14960,N_13817);
and U17453 (N_17453,N_13818,N_13687);
nand U17454 (N_17454,N_14515,N_14227);
nand U17455 (N_17455,N_13625,N_13574);
nand U17456 (N_17456,N_12860,N_12520);
nand U17457 (N_17457,N_13709,N_12915);
nand U17458 (N_17458,N_14053,N_13981);
or U17459 (N_17459,N_13867,N_13298);
xnor U17460 (N_17460,N_13191,N_14956);
xor U17461 (N_17461,N_14038,N_14079);
xor U17462 (N_17462,N_14720,N_13198);
and U17463 (N_17463,N_14828,N_13097);
and U17464 (N_17464,N_12703,N_14296);
xor U17465 (N_17465,N_12766,N_12696);
xnor U17466 (N_17466,N_14429,N_12777);
or U17467 (N_17467,N_13826,N_14477);
nand U17468 (N_17468,N_13062,N_14597);
and U17469 (N_17469,N_14703,N_14984);
nor U17470 (N_17470,N_13734,N_13454);
nand U17471 (N_17471,N_13730,N_14857);
and U17472 (N_17472,N_14775,N_12882);
nor U17473 (N_17473,N_12779,N_14419);
or U17474 (N_17474,N_13528,N_13213);
nand U17475 (N_17475,N_12955,N_14789);
or U17476 (N_17476,N_14949,N_12952);
nand U17477 (N_17477,N_14682,N_13258);
and U17478 (N_17478,N_12616,N_12809);
or U17479 (N_17479,N_14116,N_13610);
or U17480 (N_17480,N_14209,N_13075);
xor U17481 (N_17481,N_13780,N_13322);
nand U17482 (N_17482,N_13956,N_12854);
nor U17483 (N_17483,N_14762,N_13086);
or U17484 (N_17484,N_13666,N_12716);
nor U17485 (N_17485,N_13253,N_12587);
or U17486 (N_17486,N_13819,N_14881);
xor U17487 (N_17487,N_13318,N_13591);
and U17488 (N_17488,N_13264,N_14289);
xor U17489 (N_17489,N_14048,N_12872);
or U17490 (N_17490,N_13150,N_14197);
and U17491 (N_17491,N_12862,N_13154);
and U17492 (N_17492,N_14605,N_12810);
nand U17493 (N_17493,N_12503,N_12563);
or U17494 (N_17494,N_14590,N_13916);
and U17495 (N_17495,N_13607,N_14143);
xor U17496 (N_17496,N_14199,N_13407);
nor U17497 (N_17497,N_13038,N_12984);
or U17498 (N_17498,N_13275,N_12786);
nor U17499 (N_17499,N_14889,N_12809);
nor U17500 (N_17500,N_16753,N_15414);
xor U17501 (N_17501,N_16598,N_17217);
xor U17502 (N_17502,N_16431,N_15969);
xnor U17503 (N_17503,N_15380,N_15312);
xnor U17504 (N_17504,N_16810,N_15474);
or U17505 (N_17505,N_16470,N_15041);
or U17506 (N_17506,N_16168,N_16434);
nor U17507 (N_17507,N_16841,N_15092);
or U17508 (N_17508,N_15272,N_15655);
nand U17509 (N_17509,N_16881,N_15755);
nand U17510 (N_17510,N_17146,N_16048);
xnor U17511 (N_17511,N_15129,N_16556);
nor U17512 (N_17512,N_15706,N_16619);
or U17513 (N_17513,N_15248,N_15680);
or U17514 (N_17514,N_16047,N_15276);
nand U17515 (N_17515,N_16240,N_16550);
nand U17516 (N_17516,N_16879,N_16129);
xor U17517 (N_17517,N_17058,N_16067);
nor U17518 (N_17518,N_17265,N_15395);
nor U17519 (N_17519,N_16906,N_16307);
or U17520 (N_17520,N_15374,N_16063);
xnor U17521 (N_17521,N_15244,N_16682);
and U17522 (N_17522,N_15641,N_16575);
xnor U17523 (N_17523,N_15271,N_16544);
nor U17524 (N_17524,N_15894,N_16033);
and U17525 (N_17525,N_15348,N_16337);
nor U17526 (N_17526,N_17356,N_15064);
nand U17527 (N_17527,N_15168,N_17466);
nor U17528 (N_17528,N_15143,N_15379);
nor U17529 (N_17529,N_15038,N_16280);
or U17530 (N_17530,N_17410,N_15559);
nor U17531 (N_17531,N_16911,N_15998);
nand U17532 (N_17532,N_16354,N_15565);
or U17533 (N_17533,N_16254,N_15552);
nor U17534 (N_17534,N_15128,N_15822);
nand U17535 (N_17535,N_15554,N_16954);
xnor U17536 (N_17536,N_16940,N_17176);
and U17537 (N_17537,N_16673,N_16386);
xor U17538 (N_17538,N_16430,N_15991);
nand U17539 (N_17539,N_15192,N_16840);
or U17540 (N_17540,N_16790,N_16667);
and U17541 (N_17541,N_15615,N_17330);
nor U17542 (N_17542,N_15116,N_15166);
nand U17543 (N_17543,N_16686,N_16321);
xnor U17544 (N_17544,N_16006,N_16065);
xor U17545 (N_17545,N_17203,N_17370);
or U17546 (N_17546,N_17354,N_16757);
nand U17547 (N_17547,N_15747,N_16620);
or U17548 (N_17548,N_15634,N_16477);
nand U17549 (N_17549,N_15120,N_15697);
xnor U17550 (N_17550,N_17383,N_15810);
and U17551 (N_17551,N_17469,N_16356);
and U17552 (N_17552,N_15289,N_16745);
nor U17553 (N_17553,N_15577,N_15441);
xor U17554 (N_17554,N_16946,N_17348);
nand U17555 (N_17555,N_15051,N_16573);
and U17556 (N_17556,N_16135,N_15376);
or U17557 (N_17557,N_15781,N_15639);
nor U17558 (N_17558,N_15338,N_17406);
xnor U17559 (N_17559,N_16057,N_15324);
or U17560 (N_17560,N_15873,N_17191);
nor U17561 (N_17561,N_15936,N_16595);
xor U17562 (N_17562,N_16521,N_15131);
and U17563 (N_17563,N_15902,N_17188);
xnor U17564 (N_17564,N_16983,N_15540);
or U17565 (N_17565,N_16499,N_16678);
and U17566 (N_17566,N_16623,N_17210);
nor U17567 (N_17567,N_16484,N_16238);
nor U17568 (N_17568,N_17281,N_16461);
or U17569 (N_17569,N_17396,N_15549);
nand U17570 (N_17570,N_16059,N_16085);
nor U17571 (N_17571,N_15506,N_16567);
xnor U17572 (N_17572,N_15420,N_15068);
and U17573 (N_17573,N_17213,N_15584);
xnor U17574 (N_17574,N_15892,N_15572);
nor U17575 (N_17575,N_16510,N_17016);
or U17576 (N_17576,N_17273,N_16471);
nand U17577 (N_17577,N_15180,N_16007);
nand U17578 (N_17578,N_15357,N_15973);
nor U17579 (N_17579,N_17425,N_16476);
or U17580 (N_17580,N_15976,N_15996);
nor U17581 (N_17581,N_17082,N_15378);
and U17582 (N_17582,N_15161,N_15606);
nor U17583 (N_17583,N_16456,N_15829);
and U17584 (N_17584,N_15553,N_16995);
and U17585 (N_17585,N_15528,N_15284);
or U17586 (N_17586,N_15297,N_15929);
nor U17587 (N_17587,N_16074,N_17399);
nand U17588 (N_17588,N_15462,N_17483);
xor U17589 (N_17589,N_16396,N_16817);
xor U17590 (N_17590,N_16541,N_15313);
nand U17591 (N_17591,N_16522,N_15764);
or U17592 (N_17592,N_15621,N_17229);
nand U17593 (N_17593,N_15483,N_17166);
xnor U17594 (N_17594,N_17103,N_17024);
xor U17595 (N_17595,N_17062,N_16202);
or U17596 (N_17596,N_15725,N_17253);
xor U17597 (N_17597,N_16261,N_16764);
xnor U17598 (N_17598,N_15359,N_15874);
or U17599 (N_17599,N_16593,N_15020);
and U17600 (N_17600,N_15292,N_17398);
or U17601 (N_17601,N_16459,N_15527);
xor U17602 (N_17602,N_15144,N_16791);
and U17603 (N_17603,N_16862,N_17363);
and U17604 (N_17604,N_17460,N_17079);
and U17605 (N_17605,N_16565,N_16773);
or U17606 (N_17606,N_17038,N_15358);
nand U17607 (N_17607,N_15921,N_17012);
or U17608 (N_17608,N_16338,N_16821);
nand U17609 (N_17609,N_16045,N_15971);
and U17610 (N_17610,N_15728,N_15118);
and U17611 (N_17611,N_15405,N_15072);
nor U17612 (N_17612,N_16318,N_16144);
nor U17613 (N_17613,N_17431,N_17340);
nor U17614 (N_17614,N_15027,N_17452);
and U17615 (N_17615,N_16467,N_15173);
and U17616 (N_17616,N_16752,N_17465);
xor U17617 (N_17617,N_15486,N_15582);
or U17618 (N_17618,N_16640,N_15899);
nor U17619 (N_17619,N_15596,N_16343);
xnor U17620 (N_17620,N_15211,N_15365);
nand U17621 (N_17621,N_15788,N_15049);
nor U17622 (N_17622,N_16709,N_15001);
xor U17623 (N_17623,N_15366,N_16674);
and U17624 (N_17624,N_16634,N_17083);
and U17625 (N_17625,N_15856,N_16637);
xnor U17626 (N_17626,N_16600,N_16805);
nand U17627 (N_17627,N_16704,N_16286);
xor U17628 (N_17628,N_17163,N_15141);
or U17629 (N_17629,N_15022,N_15419);
nand U17630 (N_17630,N_15053,N_17366);
xor U17631 (N_17631,N_15826,N_16487);
xnor U17632 (N_17632,N_17059,N_15838);
or U17633 (N_17633,N_15662,N_17490);
xnor U17634 (N_17634,N_17400,N_16270);
or U17635 (N_17635,N_15912,N_15467);
or U17636 (N_17636,N_15784,N_16207);
nor U17637 (N_17637,N_17480,N_15354);
nor U17638 (N_17638,N_15150,N_16225);
xor U17639 (N_17639,N_16861,N_17385);
xor U17640 (N_17640,N_16108,N_15266);
xnor U17641 (N_17641,N_16251,N_15627);
and U17642 (N_17642,N_15351,N_16690);
or U17643 (N_17643,N_17044,N_16643);
or U17644 (N_17644,N_15253,N_16912);
and U17645 (N_17645,N_15385,N_17201);
nor U17646 (N_17646,N_15672,N_15981);
xor U17647 (N_17647,N_16176,N_17264);
nor U17648 (N_17648,N_17262,N_16857);
and U17649 (N_17649,N_16003,N_16241);
nor U17650 (N_17650,N_16145,N_16333);
or U17651 (N_17651,N_16425,N_15147);
or U17652 (N_17652,N_15372,N_16796);
or U17653 (N_17653,N_15602,N_15461);
nand U17654 (N_17654,N_15095,N_15328);
nand U17655 (N_17655,N_15670,N_16198);
and U17656 (N_17656,N_16093,N_17078);
xor U17657 (N_17657,N_16053,N_15862);
nand U17658 (N_17658,N_17156,N_16922);
xor U17659 (N_17659,N_15194,N_17296);
nand U17660 (N_17660,N_16956,N_16214);
and U17661 (N_17661,N_15175,N_15302);
nor U17662 (N_17662,N_16441,N_15932);
and U17663 (N_17663,N_15952,N_16485);
nor U17664 (N_17664,N_15629,N_15609);
xnor U17665 (N_17665,N_15203,N_15526);
xor U17666 (N_17666,N_17393,N_17301);
or U17667 (N_17667,N_15371,N_17242);
nor U17668 (N_17668,N_16661,N_17190);
or U17669 (N_17669,N_15361,N_16894);
or U17670 (N_17670,N_15098,N_15668);
nor U17671 (N_17671,N_17472,N_17484);
and U17672 (N_17672,N_15722,N_17423);
and U17673 (N_17673,N_15958,N_17372);
or U17674 (N_17674,N_16031,N_16827);
nor U17675 (N_17675,N_15032,N_15162);
xor U17676 (N_17676,N_17358,N_17321);
xor U17677 (N_17677,N_16604,N_16414);
nand U17678 (N_17678,N_17489,N_15455);
nor U17679 (N_17679,N_16320,N_15114);
nand U17680 (N_17680,N_17057,N_15164);
nand U17681 (N_17681,N_16304,N_16529);
xnor U17682 (N_17682,N_15630,N_15654);
or U17683 (N_17683,N_17280,N_16277);
or U17684 (N_17684,N_15108,N_16646);
xor U17685 (N_17685,N_15314,N_16961);
xor U17686 (N_17686,N_16801,N_16483);
and U17687 (N_17687,N_15469,N_17300);
and U17688 (N_17688,N_16187,N_16437);
or U17689 (N_17689,N_16591,N_16888);
nor U17690 (N_17690,N_16860,N_15881);
nor U17691 (N_17691,N_15174,N_16473);
nor U17692 (N_17692,N_16504,N_17179);
and U17693 (N_17693,N_15623,N_17223);
or U17694 (N_17694,N_16099,N_15692);
nor U17695 (N_17695,N_16271,N_17445);
xor U17696 (N_17696,N_15993,N_16289);
and U17697 (N_17697,N_17310,N_16018);
nand U17698 (N_17698,N_16957,N_17014);
and U17699 (N_17699,N_16754,N_16855);
nor U17700 (N_17700,N_15094,N_16147);
nand U17701 (N_17701,N_15088,N_16783);
nand U17702 (N_17702,N_16402,N_16442);
nor U17703 (N_17703,N_17339,N_17107);
nand U17704 (N_17704,N_16815,N_16878);
nand U17705 (N_17705,N_15423,N_16014);
or U17706 (N_17706,N_15003,N_15752);
xnor U17707 (N_17707,N_16568,N_17468);
nand U17708 (N_17708,N_15868,N_17361);
and U17709 (N_17709,N_16535,N_15063);
or U17710 (N_17710,N_15270,N_16342);
or U17711 (N_17711,N_15057,N_16421);
xnor U17712 (N_17712,N_15226,N_15675);
nand U17713 (N_17713,N_16279,N_15055);
or U17714 (N_17714,N_16518,N_16103);
or U17715 (N_17715,N_16087,N_16844);
or U17716 (N_17716,N_16895,N_17063);
or U17717 (N_17717,N_16475,N_15957);
nor U17718 (N_17718,N_16204,N_15500);
nor U17719 (N_17719,N_17180,N_17316);
nand U17720 (N_17720,N_15221,N_16589);
xnor U17721 (N_17721,N_15659,N_15727);
nand U17722 (N_17722,N_17199,N_17420);
xor U17723 (N_17723,N_15511,N_16968);
and U17724 (N_17724,N_16050,N_15513);
and U17725 (N_17725,N_17276,N_15193);
nand U17726 (N_17726,N_15917,N_16334);
nor U17727 (N_17727,N_15877,N_16724);
xor U17728 (N_17728,N_15994,N_16073);
nand U17729 (N_17729,N_15139,N_16364);
and U17730 (N_17730,N_15529,N_15903);
and U17731 (N_17731,N_15442,N_17471);
or U17732 (N_17732,N_17042,N_16676);
nand U17733 (N_17733,N_15340,N_15595);
xor U17734 (N_17734,N_16260,N_15652);
or U17735 (N_17735,N_15763,N_15674);
or U17736 (N_17736,N_16479,N_16360);
and U17737 (N_17737,N_16692,N_16398);
nor U17738 (N_17738,N_17432,N_17033);
nor U17739 (N_17739,N_15718,N_15508);
nor U17740 (N_17740,N_16186,N_16875);
and U17741 (N_17741,N_17308,N_15538);
xnor U17742 (N_17742,N_16263,N_16019);
xnor U17743 (N_17743,N_17053,N_16451);
nor U17744 (N_17744,N_15233,N_15399);
and U17745 (N_17745,N_16419,N_17257);
or U17746 (N_17746,N_16828,N_16068);
or U17747 (N_17747,N_15254,N_15574);
nand U17748 (N_17748,N_16071,N_16100);
xnor U17749 (N_17749,N_17113,N_17030);
nand U17750 (N_17750,N_15897,N_16769);
or U17751 (N_17751,N_16030,N_15050);
nor U17752 (N_17752,N_15077,N_16554);
xnor U17753 (N_17753,N_15645,N_15940);
nor U17754 (N_17754,N_15883,N_16220);
nand U17755 (N_17755,N_15824,N_16378);
and U17756 (N_17756,N_16949,N_15724);
xor U17757 (N_17757,N_16196,N_15514);
or U17758 (N_17758,N_16493,N_16997);
nor U17759 (N_17759,N_16835,N_16699);
nor U17760 (N_17760,N_15269,N_15882);
nor U17761 (N_17761,N_17164,N_15377);
nor U17762 (N_17762,N_16438,N_16596);
nand U17763 (N_17763,N_16613,N_15495);
or U17764 (N_17764,N_15091,N_16998);
nand U17765 (N_17765,N_17475,N_15096);
and U17766 (N_17766,N_17121,N_16223);
or U17767 (N_17767,N_16944,N_17120);
or U17768 (N_17768,N_17022,N_15242);
and U17769 (N_17769,N_15772,N_16269);
nor U17770 (N_17770,N_15310,N_17206);
nor U17771 (N_17771,N_15657,N_16352);
nand U17772 (N_17772,N_15210,N_16344);
or U17773 (N_17773,N_15214,N_16802);
or U17774 (N_17774,N_17129,N_17287);
or U17775 (N_17775,N_15158,N_15866);
xnor U17776 (N_17776,N_16727,N_15341);
or U17777 (N_17777,N_16300,N_15171);
and U17778 (N_17778,N_15541,N_16715);
or U17779 (N_17779,N_17158,N_15900);
nand U17780 (N_17780,N_15915,N_15619);
and U17781 (N_17781,N_16545,N_16730);
nand U17782 (N_17782,N_16055,N_17499);
nor U17783 (N_17783,N_17110,N_15044);
nor U17784 (N_17784,N_15922,N_15263);
nor U17785 (N_17785,N_15945,N_15804);
xor U17786 (N_17786,N_15575,N_15036);
or U17787 (N_17787,N_16500,N_17411);
xnor U17788 (N_17788,N_17274,N_16776);
or U17789 (N_17789,N_16605,N_15750);
nor U17790 (N_17790,N_17114,N_16088);
nand U17791 (N_17791,N_16884,N_16813);
nor U17792 (N_17792,N_15524,N_15847);
nand U17793 (N_17793,N_15653,N_15632);
nand U17794 (N_17794,N_17167,N_16206);
and U17795 (N_17795,N_15961,N_15533);
and U17796 (N_17796,N_16788,N_15539);
and U17797 (N_17797,N_15133,N_15291);
and U17798 (N_17798,N_15696,N_15382);
and U17799 (N_17799,N_16418,N_16644);
xor U17800 (N_17800,N_15317,N_17359);
and U17801 (N_17801,N_15821,N_16762);
nand U17802 (N_17802,N_16371,N_15798);
or U17803 (N_17803,N_16948,N_15779);
nor U17804 (N_17804,N_17408,N_15978);
xor U17805 (N_17805,N_16635,N_15891);
nand U17806 (N_17806,N_17171,N_16151);
nor U17807 (N_17807,N_16649,N_16517);
xor U17808 (N_17808,N_17076,N_17195);
nor U17809 (N_17809,N_17336,N_15026);
nor U17810 (N_17810,N_16236,N_16959);
nor U17811 (N_17811,N_16851,N_16587);
nand U17812 (N_17812,N_15245,N_16958);
xnor U17813 (N_17813,N_17093,N_16987);
or U17814 (N_17814,N_16527,N_15274);
or U17815 (N_17815,N_15307,N_15867);
xor U17816 (N_17816,N_17261,N_15176);
and U17817 (N_17817,N_16316,N_15217);
xnor U17818 (N_17818,N_16481,N_15628);
nand U17819 (N_17819,N_16512,N_16327);
or U17820 (N_17820,N_15910,N_16576);
and U17821 (N_17821,N_15099,N_17143);
nand U17822 (N_17822,N_15195,N_16765);
or U17823 (N_17823,N_16919,N_16152);
nor U17824 (N_17824,N_16787,N_16774);
xnor U17825 (N_17825,N_15531,N_15404);
nand U17826 (N_17826,N_15806,N_16106);
nor U17827 (N_17827,N_16384,N_17119);
nand U17828 (N_17828,N_15059,N_17297);
xor U17829 (N_17829,N_17285,N_16924);
nand U17830 (N_17830,N_16750,N_15446);
or U17831 (N_17831,N_15710,N_16420);
or U17832 (N_17832,N_15587,N_15601);
nor U17833 (N_17833,N_16651,N_16558);
and U17834 (N_17834,N_15303,N_16938);
nand U17835 (N_17835,N_16423,N_15853);
nor U17836 (N_17836,N_17258,N_15663);
or U17837 (N_17837,N_16120,N_17089);
xnor U17838 (N_17838,N_16373,N_16250);
and U17839 (N_17839,N_16910,N_15898);
nand U17840 (N_17840,N_15151,N_17311);
or U17841 (N_17841,N_15013,N_16193);
xor U17842 (N_17842,N_15428,N_15849);
nor U17843 (N_17843,N_16173,N_16592);
and U17844 (N_17844,N_16761,N_15833);
and U17845 (N_17845,N_15624,N_15391);
or U17846 (N_17846,N_15169,N_16814);
nor U17847 (N_17847,N_17312,N_17270);
and U17848 (N_17848,N_15842,N_16285);
nor U17849 (N_17849,N_16222,N_15209);
xor U17850 (N_17850,N_16149,N_15669);
nor U17851 (N_17851,N_16642,N_16991);
xnor U17852 (N_17852,N_15797,N_15614);
or U17853 (N_17853,N_15509,N_15556);
xor U17854 (N_17854,N_16266,N_16472);
nand U17855 (N_17855,N_15557,N_17160);
xor U17856 (N_17856,N_15010,N_17192);
nand U17857 (N_17857,N_16188,N_16976);
nor U17858 (N_17858,N_15626,N_16917);
or U17859 (N_17859,N_17417,N_16234);
xnor U17860 (N_17860,N_17004,N_16199);
xor U17861 (N_17861,N_15109,N_16101);
nand U17862 (N_17862,N_15618,N_15255);
nand U17863 (N_17863,N_16291,N_16697);
nand U17864 (N_17864,N_16233,N_16252);
or U17865 (N_17865,N_16812,N_16448);
or U17866 (N_17866,N_16366,N_16084);
nand U17867 (N_17867,N_15002,N_17194);
or U17868 (N_17868,N_16117,N_17225);
and U17869 (N_17869,N_15799,N_15542);
nor U17870 (N_17870,N_15861,N_15426);
and U17871 (N_17871,N_16109,N_15989);
and U17872 (N_17872,N_15362,N_15017);
nand U17873 (N_17873,N_15590,N_17478);
and U17874 (N_17874,N_16993,N_15705);
xor U17875 (N_17875,N_16929,N_16706);
xnor U17876 (N_17876,N_15406,N_16215);
nor U17877 (N_17877,N_15852,N_17134);
xnor U17878 (N_17878,N_17127,N_16695);
nor U17879 (N_17879,N_17485,N_16163);
nand U17880 (N_17880,N_16648,N_16411);
and U17881 (N_17881,N_15914,N_15383);
and U17882 (N_17882,N_16666,N_15658);
xor U17883 (N_17883,N_17350,N_15878);
nor U17884 (N_17884,N_15283,N_15074);
and U17885 (N_17885,N_15855,N_17198);
and U17886 (N_17886,N_15190,N_15103);
nand U17887 (N_17887,N_15440,N_15241);
nor U17888 (N_17888,N_16131,N_15941);
xnor U17889 (N_17889,N_16226,N_16052);
xor U17890 (N_17890,N_15097,N_16733);
nand U17891 (N_17891,N_15594,N_15968);
nor U17892 (N_17892,N_16909,N_16209);
and U17893 (N_17893,N_16182,N_15012);
xnor U17894 (N_17894,N_17045,N_15712);
or U17895 (N_17895,N_16639,N_15485);
nand U17896 (N_17896,N_15392,N_17052);
nand U17897 (N_17897,N_17434,N_16696);
nand U17898 (N_17898,N_16701,N_16989);
xor U17899 (N_17899,N_15334,N_16584);
nor U17900 (N_17900,N_15153,N_15137);
nand U17901 (N_17901,N_17453,N_15931);
and U17902 (N_17902,N_17401,N_17235);
xor U17903 (N_17903,N_16845,N_15530);
nand U17904 (N_17904,N_15223,N_15667);
nor U17905 (N_17905,N_17418,N_17096);
nand U17906 (N_17906,N_16323,N_15367);
and U17907 (N_17907,N_16161,N_16992);
and U17908 (N_17908,N_17027,N_16463);
nor U17909 (N_17909,N_15212,N_16244);
or U17910 (N_17910,N_17088,N_16941);
xor U17911 (N_17911,N_16066,N_16115);
xnor U17912 (N_17912,N_15938,N_16302);
nor U17913 (N_17913,N_16520,N_16148);
and U17914 (N_17914,N_16276,N_16039);
nand U17915 (N_17915,N_17267,N_16726);
and U17916 (N_17916,N_16986,N_15992);
nand U17917 (N_17917,N_15793,N_17123);
nor U17918 (N_17918,N_17496,N_15650);
and U17919 (N_17919,N_15316,N_16749);
or U17920 (N_17920,N_16893,N_16468);
and U17921 (N_17921,N_15684,N_15454);
nor U17922 (N_17922,N_15184,N_15682);
or U17923 (N_17923,N_15293,N_15573);
nand U17924 (N_17924,N_16886,N_16089);
nand U17925 (N_17925,N_16979,N_15548);
nor U17926 (N_17926,N_15858,N_17133);
or U17927 (N_17927,N_16332,N_17072);
nor U17928 (N_17928,N_17246,N_16408);
nor U17929 (N_17929,N_15746,N_15890);
and U17930 (N_17930,N_15389,N_16716);
or U17931 (N_17931,N_17462,N_15319);
xnor U17932 (N_17932,N_15984,N_16150);
nor U17933 (N_17933,N_17086,N_16982);
nand U17934 (N_17934,N_15815,N_15492);
and U17935 (N_17935,N_15807,N_15895);
xnor U17936 (N_17936,N_15146,N_17046);
or U17937 (N_17937,N_15988,N_17071);
or U17938 (N_17938,N_15646,N_15543);
nor U17939 (N_17939,N_15149,N_15522);
and U17940 (N_17940,N_15677,N_16114);
nand U17941 (N_17941,N_15840,N_16628);
or U17942 (N_17942,N_17305,N_15235);
or U17943 (N_17943,N_17395,N_17221);
or U17944 (N_17944,N_17112,N_17327);
nand U17945 (N_17945,N_16759,N_17433);
xnor U17946 (N_17946,N_16780,N_16656);
nor U17947 (N_17947,N_16027,N_16578);
and U17948 (N_17948,N_17230,N_16559);
xnor U17949 (N_17949,N_15709,N_15083);
nor U17950 (N_17950,N_15040,N_16617);
nor U17951 (N_17951,N_16612,N_16478);
or U17952 (N_17952,N_16610,N_17404);
or U17953 (N_17953,N_17299,N_17322);
nand U17954 (N_17954,N_16768,N_17141);
nor U17955 (N_17955,N_15222,N_15643);
and U17956 (N_17956,N_17154,N_15578);
and U17957 (N_17957,N_16928,N_16966);
or U17958 (N_17958,N_16061,N_16908);
xnor U17959 (N_17959,N_16357,N_15970);
or U17960 (N_17960,N_15859,N_16963);
and U17961 (N_17961,N_16183,N_17477);
xor U17962 (N_17962,N_15716,N_15299);
and U17963 (N_17963,N_16760,N_17003);
nand U17964 (N_17964,N_16890,N_16111);
nor U17965 (N_17965,N_16097,N_17337);
and U17966 (N_17966,N_16970,N_15258);
and U17967 (N_17967,N_15927,N_15476);
xnor U17968 (N_17968,N_16892,N_15676);
xor U17969 (N_17969,N_17272,N_15124);
xnor U17970 (N_17970,N_16837,N_17384);
or U17971 (N_17971,N_16819,N_16076);
or U17972 (N_17972,N_15751,N_16002);
and U17973 (N_17973,N_15948,N_15439);
or U17974 (N_17974,N_15787,N_17001);
nand U17975 (N_17975,N_15691,N_16169);
or U17976 (N_17976,N_16525,N_16116);
nor U17977 (N_17977,N_16918,N_16090);
or U17978 (N_17978,N_17151,N_17260);
nor U17979 (N_17979,N_17303,N_16804);
or U17980 (N_17980,N_16662,N_15637);
nor U17981 (N_17981,N_15951,N_16348);
xnor U17982 (N_17982,N_17087,N_17011);
nor U17983 (N_17983,N_16849,N_15320);
nand U17984 (N_17984,N_16950,N_15736);
xnor U17985 (N_17985,N_16735,N_17439);
nand U17986 (N_17986,N_16913,N_17211);
nor U17987 (N_17987,N_15481,N_17279);
or U17988 (N_17988,N_15130,N_15950);
or U17989 (N_17989,N_15498,N_16008);
nand U17990 (N_17990,N_16741,N_16210);
and U17991 (N_17991,N_17357,N_15197);
or U17992 (N_17992,N_17255,N_17302);
xor U17993 (N_17993,N_16417,N_16876);
nand U17994 (N_17994,N_16839,N_15305);
or U17995 (N_17995,N_15579,N_15326);
xor U17996 (N_17996,N_16079,N_17320);
or U17997 (N_17997,N_15850,N_15835);
and U17998 (N_17998,N_16519,N_16502);
xnor U17999 (N_17999,N_16679,N_16060);
nand U18000 (N_18000,N_15586,N_15488);
or U18001 (N_18001,N_15448,N_15410);
nand U18002 (N_18002,N_16809,N_16664);
nor U18003 (N_18003,N_15039,N_17189);
nand U18004 (N_18004,N_16772,N_16064);
xnor U18005 (N_18005,N_16738,N_15015);
and U18006 (N_18006,N_15105,N_16377);
nor U18007 (N_18007,N_16985,N_16655);
or U18008 (N_18008,N_16503,N_15452);
nand U18009 (N_18009,N_15142,N_15430);
and U18010 (N_18010,N_15790,N_16681);
nor U18011 (N_18011,N_16684,N_15393);
or U18012 (N_18012,N_15134,N_17147);
xnor U18013 (N_18013,N_16345,N_16947);
nand U18014 (N_18014,N_15331,N_16870);
or U18015 (N_18015,N_17185,N_15384);
xor U18016 (N_18016,N_16112,N_16823);
nand U18017 (N_18017,N_15648,N_16789);
or U18018 (N_18018,N_15318,N_15546);
xnor U18019 (N_18019,N_15823,N_16228);
xor U18020 (N_18020,N_16856,N_17268);
nand U18021 (N_18021,N_16363,N_16864);
and U18022 (N_18022,N_15880,N_16509);
and U18023 (N_18023,N_15783,N_16197);
xnor U18024 (N_18024,N_15934,N_15946);
xor U18025 (N_18025,N_16133,N_16482);
xnor U18026 (N_18026,N_15545,N_16040);
xor U18027 (N_18027,N_16630,N_15550);
or U18028 (N_18028,N_16208,N_17150);
and U18029 (N_18029,N_15631,N_15477);
nor U18030 (N_18030,N_16218,N_15995);
and U18031 (N_18031,N_17454,N_16491);
nand U18032 (N_18032,N_15346,N_17288);
nor U18033 (N_18033,N_15465,N_16191);
or U18034 (N_18034,N_15671,N_15434);
and U18035 (N_18035,N_16863,N_17440);
xnor U18036 (N_18036,N_15585,N_15535);
or U18037 (N_18037,N_15959,N_15178);
or U18038 (N_18038,N_15997,N_16967);
and U18039 (N_18039,N_15347,N_16224);
nand U18040 (N_18040,N_16091,N_15246);
and U18041 (N_18041,N_15104,N_17334);
nand U18042 (N_18042,N_16278,N_15762);
nor U18043 (N_18043,N_16355,N_15791);
or U18044 (N_18044,N_16555,N_16092);
or U18045 (N_18045,N_15851,N_16779);
or U18046 (N_18046,N_16194,N_15256);
and U18047 (N_18047,N_15794,N_17067);
xnor U18048 (N_18048,N_17216,N_16376);
nand U18049 (N_18049,N_16652,N_16290);
nor U18050 (N_18050,N_15980,N_15748);
nor U18051 (N_18051,N_15857,N_16387);
nand U18052 (N_18052,N_16590,N_15416);
nor U18053 (N_18053,N_16708,N_17218);
nor U18054 (N_18054,N_15181,N_16009);
nand U18055 (N_18055,N_16723,N_15715);
nor U18056 (N_18056,N_15126,N_17442);
nand U18057 (N_18057,N_15031,N_17013);
nand U18058 (N_18058,N_15863,N_17259);
or U18059 (N_18059,N_16582,N_15484);
and U18060 (N_18060,N_15928,N_16349);
nor U18061 (N_18061,N_17323,N_17309);
nor U18062 (N_18062,N_15381,N_15247);
or U18063 (N_18063,N_15534,N_15512);
and U18064 (N_18064,N_17144,N_17286);
and U18065 (N_18065,N_17168,N_15888);
nand U18066 (N_18066,N_15743,N_16426);
nand U18067 (N_18067,N_17345,N_17331);
nor U18068 (N_18068,N_16734,N_16155);
nand U18069 (N_18069,N_15062,N_16325);
xnor U18070 (N_18070,N_15167,N_16179);
or U18071 (N_18071,N_17173,N_15812);
xnor U18072 (N_18072,N_15033,N_16866);
or U18073 (N_18073,N_17498,N_15259);
or U18074 (N_18074,N_15695,N_16615);
and U18075 (N_18075,N_16180,N_15785);
nand U18076 (N_18076,N_16981,N_15576);
nand U18077 (N_18077,N_17208,N_16042);
and U18078 (N_18078,N_16539,N_16514);
nor U18079 (N_18079,N_16415,N_15457);
nand U18080 (N_18080,N_16372,N_15045);
or U18081 (N_18081,N_16248,N_16685);
nor U18082 (N_18082,N_17493,N_16051);
nor U18083 (N_18083,N_15975,N_17436);
xor U18084 (N_18084,N_17470,N_15123);
nor U18085 (N_18085,N_15425,N_15547);
nand U18086 (N_18086,N_15449,N_15753);
and U18087 (N_18087,N_16852,N_15982);
and U18088 (N_18088,N_15067,N_15561);
nor U18089 (N_18089,N_15865,N_16309);
and U18090 (N_18090,N_16588,N_15019);
or U18091 (N_18091,N_16854,N_15438);
and U18092 (N_18092,N_16859,N_15742);
xor U18093 (N_18093,N_16633,N_15435);
nand U18094 (N_18094,N_16795,N_15368);
and U18095 (N_18095,N_16375,N_17456);
nand U18096 (N_18096,N_15335,N_16023);
nand U18097 (N_18097,N_15085,N_15344);
and U18098 (N_18098,N_15795,N_17318);
and U18099 (N_18099,N_16873,N_16936);
xnor U18100 (N_18100,N_15121,N_17040);
nand U18101 (N_18101,N_15232,N_17152);
xor U18102 (N_18102,N_15830,N_16887);
xnor U18103 (N_18103,N_15433,N_16654);
nand U18104 (N_18104,N_15458,N_15215);
or U18105 (N_18105,N_17250,N_17497);
nor U18106 (N_18106,N_16025,N_16160);
or U18107 (N_18107,N_16897,N_15544);
nor U18108 (N_18108,N_16004,N_16232);
nor U18109 (N_18109,N_17157,N_16939);
or U18110 (N_18110,N_15160,N_16832);
nor U18111 (N_18111,N_17325,N_16346);
nor U18112 (N_18112,N_16369,N_16058);
and U18113 (N_18113,N_15239,N_15827);
and U18114 (N_18114,N_16794,N_17204);
or U18115 (N_18115,N_15520,N_15521);
or U18116 (N_18116,N_15909,N_16036);
nor U18117 (N_18117,N_16718,N_15219);
nor U18118 (N_18118,N_16742,N_16022);
nand U18119 (N_18119,N_16454,N_17051);
or U18120 (N_18120,N_15635,N_15225);
xnor U18121 (N_18121,N_17077,N_15711);
or U18122 (N_18122,N_16677,N_16636);
nand U18123 (N_18123,N_16937,N_16381);
and U18124 (N_18124,N_16283,N_16172);
nand U18125 (N_18125,N_15375,N_15583);
xor U18126 (N_18126,N_16113,N_16404);
nand U18127 (N_18127,N_15649,N_17283);
or U18128 (N_18128,N_17313,N_16563);
nor U18129 (N_18129,N_17373,N_17021);
or U18130 (N_18130,N_16212,N_15636);
nor U18131 (N_18131,N_17414,N_16942);
nand U18132 (N_18132,N_15260,N_15268);
or U18133 (N_18133,N_15218,N_16146);
and U18134 (N_18134,N_17379,N_16299);
nor U18135 (N_18135,N_15599,N_15523);
nor U18136 (N_18136,N_17200,N_16931);
nor U18137 (N_18137,N_15445,N_16329);
nor U18138 (N_18138,N_15777,N_16698);
nand U18139 (N_18139,N_16907,N_16842);
or U18140 (N_18140,N_15930,N_17403);
nand U18141 (N_18141,N_15122,N_16392);
or U18142 (N_18142,N_15157,N_16847);
or U18143 (N_18143,N_17066,N_16178);
nor U18144 (N_18144,N_15421,N_16326);
nand U18145 (N_18145,N_15007,N_15417);
or U18146 (N_18146,N_17377,N_15593);
nor U18147 (N_18147,N_15819,N_15363);
xnor U18148 (N_18148,N_17232,N_17131);
xor U18149 (N_18149,N_16308,N_16551);
nor U18150 (N_18150,N_17324,N_16751);
or U18151 (N_18151,N_15870,N_16916);
xor U18152 (N_18152,N_15700,N_16157);
nand U18153 (N_18153,N_15845,N_15478);
or U18154 (N_18154,N_15415,N_15854);
xor U18155 (N_18155,N_15154,N_16663);
nand U18156 (N_18156,N_15499,N_16341);
xor U18157 (N_18157,N_17364,N_17054);
and U18158 (N_18158,N_16490,N_17343);
or U18159 (N_18159,N_17142,N_17205);
nand U18160 (N_18160,N_15678,N_16331);
xor U18161 (N_18161,N_16062,N_16268);
and U18162 (N_18162,N_15688,N_16086);
or U18163 (N_18163,N_17175,N_15687);
nand U18164 (N_18164,N_15983,N_16755);
nand U18165 (N_18165,N_15413,N_16399);
xor U18166 (N_18166,N_15825,N_16505);
and U18167 (N_18167,N_16528,N_17026);
and U18168 (N_18168,N_16707,N_15885);
nor U18169 (N_18169,N_15089,N_16166);
and U18170 (N_18170,N_16833,N_15884);
xor U18171 (N_18171,N_16711,N_16903);
nand U18172 (N_18172,N_15820,N_16035);
nand U18173 (N_18173,N_15183,N_16243);
and U18174 (N_18174,N_17020,N_15516);
and U18175 (N_18175,N_17237,N_16850);
and U18176 (N_18176,N_15186,N_16822);
and U18177 (N_18177,N_15112,N_16523);
and U18178 (N_18178,N_16336,N_17226);
and U18179 (N_18179,N_15911,N_15875);
xnor U18180 (N_18180,N_16132,N_15836);
xnor U18181 (N_18181,N_17252,N_16351);
and U18182 (N_18182,N_15679,N_15739);
and U18183 (N_18183,N_17349,N_17090);
nand U18184 (N_18184,N_16219,N_15396);
and U18185 (N_18185,N_17031,N_15612);
nand U18186 (N_18186,N_16943,N_17064);
and U18187 (N_18187,N_17092,N_15555);
xor U18188 (N_18188,N_15407,N_15065);
or U18189 (N_18189,N_17032,N_16952);
nor U18190 (N_18190,N_15280,N_15960);
nand U18191 (N_18191,N_15402,N_15749);
xor U18192 (N_18192,N_17174,N_15016);
or U18193 (N_18193,N_15411,N_16536);
nand U18194 (N_18194,N_15605,N_16046);
nand U18195 (N_18195,N_15412,N_15087);
xor U18196 (N_18196,N_15592,N_15343);
xnor U18197 (N_18197,N_17391,N_16553);
nand U18198 (N_18198,N_16581,N_17037);
or U18199 (N_18199,N_17249,N_16028);
xnor U18200 (N_18200,N_16195,N_16353);
or U18201 (N_18201,N_15400,N_16675);
nor U18202 (N_18202,N_16400,N_15397);
or U18203 (N_18203,N_17155,N_16306);
nor U18204 (N_18204,N_16669,N_15464);
or U18205 (N_18205,N_17117,N_16339);
or U18206 (N_18206,N_16192,N_16720);
nor U18207 (N_18207,N_16239,N_15110);
nor U18208 (N_18208,N_15262,N_15604);
nor U18209 (N_18209,N_17298,N_16122);
xnor U18210 (N_18210,N_16139,N_16609);
nand U18211 (N_18211,N_16165,N_17438);
and U18212 (N_18212,N_15665,N_15443);
nor U18213 (N_18213,N_16811,N_16935);
nand U18214 (N_18214,N_16303,N_16782);
and U18215 (N_18215,N_15352,N_16631);
xnor U18216 (N_18216,N_16549,N_15904);
nor U18217 (N_18217,N_15234,N_16955);
or U18218 (N_18218,N_17389,N_16393);
or U18219 (N_18219,N_15999,N_15182);
xor U18220 (N_18220,N_16439,N_16200);
xor U18221 (N_18221,N_16577,N_15745);
and U18222 (N_18222,N_15600,N_16310);
nor U18223 (N_18223,N_16102,N_17458);
xor U18224 (N_18224,N_15610,N_17109);
or U18225 (N_18225,N_17319,N_16242);
and U18226 (N_18226,N_15954,N_15388);
nor U18227 (N_18227,N_15403,N_16818);
or U18228 (N_18228,N_17202,N_16170);
xor U18229 (N_18229,N_16719,N_17457);
and U18230 (N_18230,N_16158,N_17227);
and U18231 (N_18231,N_16580,N_17376);
nand U18232 (N_18232,N_16846,N_15236);
or U18233 (N_18233,N_15776,N_15698);
xnor U18234 (N_18234,N_17284,N_17314);
xnor U18235 (N_18235,N_15907,N_16319);
nor U18236 (N_18236,N_16401,N_16853);
or U18237 (N_18237,N_16466,N_15207);
xor U18238 (N_18238,N_17132,N_16245);
xnor U18239 (N_18239,N_16389,N_15102);
or U18240 (N_18240,N_16496,N_15315);
nand U18241 (N_18241,N_16960,N_17122);
xnor U18242 (N_18242,N_17165,N_16777);
nor U18243 (N_18243,N_16365,N_16725);
and U18244 (N_18244,N_17028,N_17068);
nor U18245 (N_18245,N_16140,N_15767);
and U18246 (N_18246,N_15598,N_17482);
and U18247 (N_18247,N_15809,N_17292);
nand U18248 (N_18248,N_15702,N_15202);
nor U18249 (N_18249,N_16262,N_16702);
or U18250 (N_18250,N_16181,N_17412);
and U18251 (N_18251,N_17104,N_16249);
xnor U18252 (N_18252,N_16574,N_16650);
nor U18253 (N_18253,N_15090,N_16246);
or U18254 (N_18254,N_15803,N_16340);
or U18255 (N_18255,N_16237,N_15796);
nand U18256 (N_18256,N_15198,N_15093);
or U18257 (N_18257,N_15265,N_17214);
nor U18258 (N_18258,N_15906,N_16190);
or U18259 (N_18259,N_15733,N_15350);
or U18260 (N_18260,N_16534,N_15075);
nor U18261 (N_18261,N_16572,N_15864);
and U18262 (N_18262,N_15277,N_15170);
and U18263 (N_18263,N_15778,N_15768);
and U18264 (N_18264,N_16978,N_16601);
xnor U18265 (N_18265,N_15000,N_15972);
nand U18266 (N_18266,N_16533,N_16721);
and U18267 (N_18267,N_16930,N_16474);
nand U18268 (N_18268,N_16034,N_15480);
and U18269 (N_18269,N_15977,N_17084);
nand U18270 (N_18270,N_15496,N_15287);
nand U18271 (N_18271,N_15082,N_16898);
and U18272 (N_18272,N_15304,N_16570);
nand U18273 (N_18273,N_17241,N_16824);
nand U18274 (N_18274,N_16831,N_15035);
xnor U18275 (N_18275,N_15052,N_15213);
nor U18276 (N_18276,N_16830,N_16501);
nand U18277 (N_18277,N_17234,N_17491);
nand U18278 (N_18278,N_17135,N_17486);
and U18279 (N_18279,N_16041,N_17035);
nand U18280 (N_18280,N_16710,N_15782);
or U18281 (N_18281,N_17422,N_16990);
nand U18282 (N_18282,N_16971,N_16107);
nand U18283 (N_18283,N_16792,N_16566);
nor U18284 (N_18284,N_15633,N_16142);
nand U18285 (N_18285,N_15336,N_16359);
or U18286 (N_18286,N_17271,N_16530);
and U18287 (N_18287,N_15566,N_16994);
xor U18288 (N_18288,N_15966,N_15437);
or U18289 (N_18289,N_15730,N_15588);
or U18290 (N_18290,N_16380,N_16693);
xnor U18291 (N_18291,N_15505,N_16513);
and U18292 (N_18292,N_15084,N_15756);
or U18293 (N_18293,N_17474,N_17282);
xor U18294 (N_18294,N_15282,N_16744);
or U18295 (N_18295,N_15519,N_15311);
and U18296 (N_18296,N_16105,N_16096);
and U18297 (N_18297,N_15551,N_16923);
nand U18298 (N_18298,N_16433,N_16800);
or U18299 (N_18299,N_16315,N_16546);
nand U18300 (N_18300,N_15869,N_16292);
xnor U18301 (N_18301,N_16080,N_15229);
nand U18302 (N_18302,N_16552,N_17463);
nor U18303 (N_18303,N_17041,N_16743);
or U18304 (N_18304,N_15689,N_17008);
and U18305 (N_18305,N_15949,N_15786);
nand U18306 (N_18306,N_16784,N_15196);
nand U18307 (N_18307,N_16413,N_17055);
or U18308 (N_18308,N_15054,N_15436);
xnor U18309 (N_18309,N_17183,N_15373);
or U18310 (N_18310,N_15515,N_15138);
and U18311 (N_18311,N_17007,N_16597);
or U18312 (N_18312,N_16618,N_16446);
and U18313 (N_18313,N_15200,N_17006);
nand U18314 (N_18314,N_15939,N_16128);
nand U18315 (N_18315,N_15243,N_15460);
xor U18316 (N_18316,N_16868,N_17448);
and U18317 (N_18317,N_16629,N_15386);
and U18318 (N_18318,N_15811,N_15805);
or U18319 (N_18319,N_15332,N_16799);
nand U18320 (N_18320,N_17351,N_15444);
and U18321 (N_18321,N_17182,N_16221);
xor U18322 (N_18322,N_16436,N_15876);
nand U18323 (N_18323,N_15908,N_15647);
xor U18324 (N_18324,N_15281,N_17464);
nand U18325 (N_18325,N_17451,N_17098);
nor U18326 (N_18326,N_15721,N_15451);
or U18327 (N_18327,N_15401,N_16611);
xnor U18328 (N_18328,N_15148,N_15069);
nor U18329 (N_18329,N_16255,N_16069);
nor U18330 (N_18330,N_15353,N_16072);
and U18331 (N_18331,N_15325,N_16660);
and U18332 (N_18332,N_17074,N_16259);
and U18333 (N_18333,N_15740,N_16098);
xor U18334 (N_18334,N_17115,N_15708);
xnor U18335 (N_18335,N_16497,N_17080);
nand U18336 (N_18336,N_16189,N_15597);
nor U18337 (N_18337,N_16156,N_15567);
xor U18338 (N_18338,N_17140,N_15701);
xnor U18339 (N_18339,N_16808,N_15923);
xnor U18340 (N_18340,N_15046,N_15076);
xnor U18341 (N_18341,N_16427,N_16460);
nor U18342 (N_18342,N_15155,N_16138);
xnor U18343 (N_18343,N_15887,N_16999);
nand U18344 (N_18344,N_17447,N_16767);
nand U18345 (N_18345,N_17029,N_15296);
nor U18346 (N_18346,N_16313,N_16880);
or U18347 (N_18347,N_17170,N_16301);
nand U18348 (N_18348,N_17329,N_17009);
and U18349 (N_18349,N_17137,N_15078);
xnor U18350 (N_18350,N_15510,N_17224);
or U18351 (N_18351,N_17149,N_17219);
nor U18352 (N_18352,N_17317,N_16267);
and U18353 (N_18353,N_16740,N_17069);
nand U18354 (N_18354,N_17307,N_16462);
xor U18355 (N_18355,N_17461,N_17421);
and U18356 (N_18356,N_16095,N_16953);
nand U18357 (N_18357,N_16024,N_16739);
nor U18358 (N_18358,N_16049,N_16691);
or U18359 (N_18359,N_17415,N_16756);
nor U18360 (N_18360,N_17481,N_15962);
nor U18361 (N_18361,N_16077,N_16763);
nor U18362 (N_18362,N_15843,N_16450);
and U18363 (N_18363,N_16770,N_17378);
nor U18364 (N_18364,N_16798,N_17102);
nor U18365 (N_18365,N_15127,N_15119);
nand U18366 (N_18366,N_15872,N_17392);
and U18367 (N_18367,N_17402,N_15471);
or U18368 (N_18368,N_16217,N_15345);
or U18369 (N_18369,N_16368,N_16561);
and U18370 (N_18370,N_16626,N_16227);
nand U18371 (N_18371,N_17315,N_16647);
and U18372 (N_18372,N_16524,N_16312);
nand U18373 (N_18373,N_17073,N_16374);
or U18374 (N_18374,N_16511,N_16902);
xnor U18375 (N_18375,N_17333,N_15490);
nor U18376 (N_18376,N_17369,N_15986);
or U18377 (N_18377,N_17139,N_16858);
and U18378 (N_18378,N_16562,N_16607);
xor U18379 (N_18379,N_17172,N_16167);
and U18380 (N_18380,N_17124,N_15501);
nor U18381 (N_18381,N_15642,N_15935);
nand U18382 (N_18382,N_15238,N_15489);
or U18383 (N_18383,N_16492,N_16516);
and U18384 (N_18384,N_17446,N_17197);
and U18385 (N_18385,N_15479,N_16044);
xor U18386 (N_18386,N_15106,N_16032);
nand U18387 (N_18387,N_17335,N_15023);
nor U18388 (N_18388,N_15249,N_16540);
xnor U18389 (N_18389,N_15942,N_16786);
nand U18390 (N_18390,N_16543,N_16975);
and U18391 (N_18391,N_15330,N_16901);
and U18392 (N_18392,N_15517,N_16201);
and U18393 (N_18393,N_16383,N_17081);
or U18394 (N_18394,N_16037,N_16429);
xor U18395 (N_18395,N_16391,N_15985);
or U18396 (N_18396,N_16125,N_15879);
and U18397 (N_18397,N_16579,N_15955);
nor U18398 (N_18398,N_16964,N_15589);
or U18399 (N_18399,N_17061,N_16011);
xor U18400 (N_18400,N_15525,N_16185);
nor U18401 (N_18401,N_15737,N_16825);
nand U18402 (N_18402,N_16457,N_16489);
nand U18403 (N_18403,N_16896,N_17236);
nor U18404 (N_18404,N_15447,N_17049);
xor U18405 (N_18405,N_15279,N_15660);
xnor U18406 (N_18406,N_15937,N_16515);
and U18407 (N_18407,N_15224,N_16614);
and U18408 (N_18408,N_15569,N_17294);
or U18409 (N_18409,N_15409,N_16700);
nand U18410 (N_18410,N_15159,N_16328);
nand U18411 (N_18411,N_15030,N_17347);
nand U18412 (N_18412,N_17390,N_15603);
nor U18413 (N_18413,N_15278,N_16211);
nor U18414 (N_18414,N_15327,N_15177);
or U18415 (N_18415,N_16412,N_15113);
nor U18416 (N_18416,N_16385,N_17130);
or U18417 (N_18417,N_16867,N_15140);
xnor U18418 (N_18418,N_16432,N_15285);
or U18419 (N_18419,N_15841,N_15694);
xor U18420 (N_18420,N_17075,N_15086);
nand U18421 (N_18421,N_16311,N_15732);
or U18422 (N_18422,N_16882,N_15661);
and U18423 (N_18423,N_17413,N_15780);
and U18424 (N_18424,N_16820,N_16671);
nand U18425 (N_18425,N_16110,N_16653);
or U18426 (N_18426,N_16465,N_16972);
or U18427 (N_18427,N_15638,N_16921);
nor U18428 (N_18428,N_16732,N_15580);
and U18429 (N_18429,N_15275,N_15848);
and U18430 (N_18430,N_16508,N_15494);
and U18431 (N_18431,N_17374,N_16174);
nand U18432 (N_18432,N_17444,N_15066);
and U18433 (N_18433,N_15532,N_15886);
or U18434 (N_18434,N_17266,N_15228);
nor U18435 (N_18435,N_17495,N_17449);
xor U18436 (N_18436,N_16367,N_15611);
and U18437 (N_18437,N_17346,N_15360);
or U18438 (N_18438,N_16729,N_16548);
xnor U18439 (N_18439,N_16542,N_15644);
and U18440 (N_18440,N_17161,N_16606);
nand U18441 (N_18441,N_16872,N_17025);
xor U18442 (N_18442,N_15704,N_17492);
nand U18443 (N_18443,N_16962,N_16594);
or U18444 (N_18444,N_15920,N_17435);
or U18445 (N_18445,N_16627,N_15432);
and U18446 (N_18446,N_16253,N_16026);
nand U18447 (N_18447,N_16689,N_17240);
nand U18448 (N_18448,N_15301,N_16075);
nor U18449 (N_18449,N_15172,N_15683);
nor U18450 (N_18450,N_16899,N_15714);
nor U18451 (N_18451,N_16771,N_16670);
and U18452 (N_18452,N_15286,N_16883);
nand U18453 (N_18453,N_17397,N_17125);
nand U18454 (N_18454,N_16256,N_15355);
xor U18455 (N_18455,N_15773,N_16748);
xnor U18456 (N_18456,N_17409,N_16758);
or U18457 (N_18457,N_16532,N_16622);
nand U18458 (N_18458,N_16265,N_15468);
nand U18459 (N_18459,N_15979,N_15924);
or U18460 (N_18460,N_15625,N_15398);
xnor U18461 (N_18461,N_16284,N_15227);
nand U18462 (N_18462,N_16632,N_15792);
nand U18463 (N_18463,N_17278,N_16118);
nand U18464 (N_18464,N_16127,N_16797);
nor U18465 (N_18465,N_16370,N_17269);
and U18466 (N_18466,N_17018,N_16714);
nor U18467 (N_18467,N_17091,N_15298);
xor U18468 (N_18468,N_15450,N_17162);
xnor U18469 (N_18469,N_15204,N_15713);
or U18470 (N_18470,N_17382,N_15422);
xor U18471 (N_18471,N_15518,N_17019);
nand U18472 (N_18472,N_16296,N_16969);
nand U18473 (N_18473,N_16445,N_16571);
nor U18474 (N_18474,N_15006,N_17036);
or U18475 (N_18475,N_17184,N_17494);
xnor U18476 (N_18476,N_16164,N_17169);
nor U18477 (N_18477,N_15775,N_16016);
nor U18478 (N_18478,N_16205,N_17332);
nand U18479 (N_18479,N_15800,N_15189);
nand U18480 (N_18480,N_16362,N_16104);
xnor U18481 (N_18481,N_15808,N_16264);
nand U18482 (N_18482,N_16793,N_15766);
nand U18483 (N_18483,N_15613,N_15967);
nand U18484 (N_18484,N_17186,N_16231);
and U18485 (N_18485,N_16247,N_15844);
nor U18486 (N_18486,N_16130,N_15493);
or U18487 (N_18487,N_16469,N_15250);
and U18488 (N_18488,N_16945,N_16537);
nor U18489 (N_18489,N_17341,N_15919);
or U18490 (N_18490,N_17215,N_17352);
nor U18491 (N_18491,N_15329,N_15342);
nand U18492 (N_18492,N_15738,N_15107);
or U18493 (N_18493,N_15568,N_15216);
xnor U18494 (N_18494,N_16317,N_16659);
and U18495 (N_18495,N_15789,N_16136);
and U18496 (N_18496,N_15475,N_15944);
or U18497 (N_18497,N_15571,N_15562);
and U18498 (N_18498,N_16177,N_15056);
xnor U18499 (N_18499,N_16586,N_15060);
or U18500 (N_18500,N_16781,N_17430);
or U18501 (N_18501,N_17371,N_15987);
and U18502 (N_18502,N_17100,N_16121);
nand U18503 (N_18503,N_15502,N_15364);
or U18504 (N_18504,N_16672,N_16203);
or U18505 (N_18505,N_16885,N_15681);
nor U18506 (N_18506,N_15179,N_15860);
nor U18507 (N_18507,N_17289,N_16694);
nor U18508 (N_18508,N_17047,N_17050);
xnor U18509 (N_18509,N_16775,N_16834);
nand U18510 (N_18510,N_16171,N_15754);
and U18511 (N_18511,N_15008,N_15163);
nor U18512 (N_18512,N_15080,N_17256);
xor U18513 (N_18513,N_16616,N_17002);
and U18514 (N_18514,N_15037,N_16891);
and U18515 (N_18515,N_15707,N_16602);
xor U18516 (N_18516,N_16645,N_16394);
xor U18517 (N_18517,N_17459,N_16440);
and U18518 (N_18518,N_17473,N_16070);
or U18519 (N_18519,N_15759,N_16703);
nor U18520 (N_18520,N_16424,N_15918);
xor U18521 (N_18521,N_16920,N_15760);
or U18522 (N_18522,N_17043,N_16984);
or U18523 (N_18523,N_17116,N_15136);
nand U18524 (N_18524,N_15048,N_17212);
nor U18525 (N_18525,N_17326,N_15071);
nand U18526 (N_18526,N_15021,N_15025);
or U18527 (N_18527,N_17118,N_17441);
or U18528 (N_18528,N_16322,N_15507);
or U18529 (N_18529,N_16980,N_17017);
xnor U18530 (N_18530,N_15816,N_15761);
xnor U18531 (N_18531,N_17178,N_15974);
nand U18532 (N_18532,N_16829,N_17136);
nand U18533 (N_18533,N_15473,N_16314);
nand U18534 (N_18534,N_16282,N_16082);
or U18535 (N_18535,N_15264,N_16915);
or U18536 (N_18536,N_17181,N_15817);
and U18537 (N_18537,N_17338,N_16488);
xnor U18538 (N_18538,N_15294,N_15774);
nor U18539 (N_18539,N_16010,N_16747);
xor U18540 (N_18540,N_15504,N_16925);
nor U18541 (N_18541,N_16235,N_15308);
nor U18542 (N_18542,N_15956,N_15288);
xnor U18543 (N_18543,N_17248,N_15252);
xor U18544 (N_18544,N_15156,N_16162);
xnor U18545 (N_18545,N_17138,N_15191);
nand U18546 (N_18546,N_15871,N_15491);
nor U18547 (N_18547,N_16974,N_15240);
or U18548 (N_18548,N_15230,N_16153);
nor U18549 (N_18549,N_15005,N_15424);
and U18550 (N_18550,N_16137,N_17426);
nand U18551 (N_18551,N_17375,N_16583);
and U18552 (N_18552,N_16410,N_17177);
or U18553 (N_18553,N_16012,N_15014);
and U18554 (N_18554,N_17238,N_15472);
nor U18555 (N_18555,N_17424,N_17380);
nor U18556 (N_18556,N_15206,N_17467);
xnor U18557 (N_18557,N_16625,N_16877);
or U18558 (N_18558,N_16350,N_15261);
nor U18559 (N_18559,N_16494,N_16230);
or U18560 (N_18560,N_16480,N_15666);
and U18561 (N_18561,N_17010,N_16889);
nor U18562 (N_18562,N_15560,N_16021);
nand U18563 (N_18563,N_17222,N_15018);
nor U18564 (N_18564,N_17228,N_16298);
or U18565 (N_18565,N_16013,N_17106);
xnor U18566 (N_18566,N_16486,N_16932);
xnor U18567 (N_18567,N_16293,N_17239);
or U18568 (N_18568,N_16599,N_16458);
and U18569 (N_18569,N_16435,N_15734);
nand U18570 (N_18570,N_16531,N_15965);
or U18571 (N_18571,N_17488,N_17291);
nor U18572 (N_18572,N_16657,N_17039);
xor U18573 (N_18573,N_17251,N_16056);
or U18574 (N_18574,N_15889,N_17476);
nand U18575 (N_18575,N_16507,N_15834);
or U18576 (N_18576,N_16848,N_15640);
or U18577 (N_18577,N_17386,N_15802);
and U18578 (N_18578,N_17381,N_16816);
xnor U18579 (N_18579,N_16403,N_17455);
nor U18580 (N_18580,N_15690,N_15251);
nand U18581 (N_18581,N_15004,N_16015);
nor U18582 (N_18582,N_16665,N_15100);
and U18583 (N_18583,N_15616,N_16766);
nor U18584 (N_18584,N_16836,N_17097);
or U18585 (N_18585,N_15029,N_16865);
and U18586 (N_18586,N_16495,N_16449);
or U18587 (N_18587,N_16216,N_17070);
nand U18588 (N_18588,N_16621,N_15470);
xnor U18589 (N_18589,N_16281,N_16965);
and U18590 (N_18590,N_15720,N_15893);
nand U18591 (N_18591,N_15188,N_17405);
xnor U18592 (N_18592,N_16560,N_16506);
nor U18593 (N_18593,N_17407,N_15073);
xnor U18594 (N_18594,N_17085,N_16933);
or U18595 (N_18595,N_15418,N_16297);
nand U18596 (N_18596,N_17126,N_15564);
or U18597 (N_18597,N_15145,N_15322);
and U18598 (N_18598,N_16705,N_16409);
or U18599 (N_18599,N_15152,N_16641);
nor U18600 (N_18600,N_15656,N_17193);
and U18601 (N_18601,N_16874,N_16294);
xor U18602 (N_18602,N_16288,N_16330);
nand U18603 (N_18603,N_16807,N_15744);
xor U18604 (N_18604,N_15769,N_15741);
xor U18605 (N_18605,N_15536,N_16806);
or U18606 (N_18606,N_15456,N_16143);
and U18607 (N_18607,N_17342,N_17328);
nor U18608 (N_18608,N_16347,N_16422);
or U18609 (N_18609,N_17108,N_16843);
nor U18610 (N_18610,N_15132,N_15042);
and U18611 (N_18611,N_15607,N_16305);
and U18612 (N_18612,N_16871,N_17209);
and U18613 (N_18613,N_15591,N_15356);
and U18614 (N_18614,N_15237,N_15231);
or U18615 (N_18615,N_17101,N_16668);
or U18616 (N_18616,N_15390,N_15832);
xor U18617 (N_18617,N_15814,N_15664);
nand U18618 (N_18618,N_16295,N_16464);
nor U18619 (N_18619,N_16078,N_15337);
nand U18620 (N_18620,N_15273,N_15011);
or U18621 (N_18621,N_15699,N_17263);
and U18622 (N_18622,N_16838,N_15201);
and U18623 (N_18623,N_16728,N_16526);
nand U18624 (N_18624,N_17344,N_16977);
and U18625 (N_18625,N_17387,N_17231);
or U18626 (N_18626,N_17487,N_15719);
nor U18627 (N_18627,N_16397,N_15497);
xor U18628 (N_18628,N_16900,N_17290);
or U18629 (N_18629,N_15453,N_16658);
nand U18630 (N_18630,N_16175,N_17368);
nor U18631 (N_18631,N_15620,N_16904);
xnor U18632 (N_18632,N_16416,N_15309);
or U18633 (N_18633,N_16585,N_15839);
nor U18634 (N_18634,N_15333,N_17275);
xnor U18635 (N_18635,N_15896,N_17428);
and U18636 (N_18636,N_16498,N_16081);
nand U18637 (N_18637,N_16083,N_15925);
xor U18638 (N_18638,N_16683,N_17416);
nor U18639 (N_18639,N_17244,N_15081);
and U18640 (N_18640,N_16029,N_17220);
or U18641 (N_18641,N_15135,N_17233);
and U18642 (N_18642,N_17005,N_16275);
or U18643 (N_18643,N_15916,N_15686);
nand U18644 (N_18644,N_17095,N_15061);
or U18645 (N_18645,N_16869,N_15926);
nor U18646 (N_18646,N_16443,N_16785);
and U18647 (N_18647,N_17034,N_15731);
and U18648 (N_18648,N_15570,N_16184);
and U18649 (N_18649,N_17207,N_15723);
nand U18650 (N_18650,N_15185,N_17394);
nand U18651 (N_18651,N_16390,N_16731);
xor U18652 (N_18652,N_15370,N_16043);
nor U18653 (N_18653,N_15617,N_16538);
nand U18654 (N_18654,N_15257,N_16407);
xnor U18655 (N_18655,N_15117,N_15463);
and U18656 (N_18656,N_17247,N_16229);
and U18657 (N_18657,N_17293,N_15058);
nor U18658 (N_18658,N_16453,N_15369);
and U18659 (N_18659,N_17023,N_16608);
nor U18660 (N_18660,N_17056,N_15125);
nand U18661 (N_18661,N_15765,N_15187);
nand U18662 (N_18662,N_15963,N_15408);
xor U18663 (N_18663,N_15043,N_15208);
nand U18664 (N_18664,N_16569,N_15729);
and U18665 (N_18665,N_15339,N_16951);
nor U18666 (N_18666,N_16124,N_16017);
or U18667 (N_18667,N_17388,N_15828);
or U18668 (N_18668,N_16126,N_15953);
nor U18669 (N_18669,N_15622,N_15427);
nand U18670 (N_18670,N_16257,N_15651);
and U18671 (N_18671,N_16154,N_17000);
or U18672 (N_18672,N_16712,N_16736);
nor U18673 (N_18673,N_16379,N_16624);
xor U18674 (N_18674,N_15321,N_16934);
nand U18675 (N_18675,N_17443,N_17015);
xor U18676 (N_18676,N_16826,N_16746);
or U18677 (N_18677,N_16778,N_15101);
nor U18678 (N_18678,N_15024,N_17105);
nor U18679 (N_18679,N_16361,N_17295);
or U18680 (N_18680,N_15034,N_17148);
nor U18681 (N_18681,N_15466,N_16803);
xor U18682 (N_18682,N_17128,N_16020);
nand U18683 (N_18683,N_15028,N_17367);
nand U18684 (N_18684,N_16094,N_15673);
nand U18685 (N_18685,N_15482,N_16119);
nor U18686 (N_18686,N_17159,N_17065);
and U18687 (N_18687,N_15990,N_16638);
nor U18688 (N_18688,N_15703,N_15165);
or U18689 (N_18689,N_15487,N_15306);
nor U18690 (N_18690,N_17243,N_15685);
nor U18691 (N_18691,N_16996,N_16557);
nor U18692 (N_18692,N_16914,N_17355);
xnor U18693 (N_18693,N_15758,N_17254);
and U18694 (N_18694,N_17450,N_15813);
or U18695 (N_18695,N_16680,N_17111);
nor U18696 (N_18696,N_16273,N_17304);
nor U18697 (N_18697,N_15220,N_15717);
nand U18698 (N_18698,N_15079,N_15199);
xor U18699 (N_18699,N_16447,N_15429);
nand U18700 (N_18700,N_17360,N_16713);
nor U18701 (N_18701,N_16324,N_16388);
nor U18702 (N_18702,N_15537,N_15771);
or U18703 (N_18703,N_15431,N_16926);
or U18704 (N_18704,N_15459,N_16274);
or U18705 (N_18705,N_15563,N_15503);
or U18706 (N_18706,N_17153,N_15964);
nor U18707 (N_18707,N_17145,N_17479);
nand U18708 (N_18708,N_15387,N_15394);
and U18709 (N_18709,N_15290,N_15801);
xor U18710 (N_18710,N_15267,N_15933);
nor U18711 (N_18711,N_15757,N_15295);
nor U18712 (N_18712,N_15735,N_16737);
xor U18713 (N_18713,N_15901,N_15837);
xor U18714 (N_18714,N_16717,N_15323);
nor U18715 (N_18715,N_16688,N_15558);
or U18716 (N_18716,N_16988,N_15846);
nor U18717 (N_18717,N_16395,N_16687);
or U18718 (N_18718,N_17427,N_16973);
or U18719 (N_18719,N_15770,N_15009);
and U18720 (N_18720,N_16428,N_16123);
or U18721 (N_18721,N_15726,N_16000);
xnor U18722 (N_18722,N_17353,N_16406);
xor U18723 (N_18723,N_16722,N_16005);
xnor U18724 (N_18724,N_17277,N_16272);
nor U18725 (N_18725,N_15581,N_16159);
or U18726 (N_18726,N_17048,N_16603);
nand U18727 (N_18727,N_17060,N_17187);
nand U18728 (N_18728,N_16452,N_16564);
xor U18729 (N_18729,N_15905,N_15047);
xor U18730 (N_18730,N_16287,N_15608);
or U18731 (N_18731,N_17437,N_16444);
nor U18732 (N_18732,N_17099,N_16258);
and U18733 (N_18733,N_17306,N_16335);
and U18734 (N_18734,N_17429,N_17362);
and U18735 (N_18735,N_15300,N_15205);
nor U18736 (N_18736,N_16905,N_15818);
nor U18737 (N_18737,N_16358,N_15943);
nand U18738 (N_18738,N_17094,N_16054);
nand U18739 (N_18739,N_16213,N_16038);
and U18740 (N_18740,N_15913,N_16455);
and U18741 (N_18741,N_16001,N_15070);
xor U18742 (N_18742,N_16141,N_16382);
xnor U18743 (N_18743,N_15115,N_17419);
and U18744 (N_18744,N_16927,N_16405);
or U18745 (N_18745,N_15831,N_17245);
and U18746 (N_18746,N_17196,N_16547);
or U18747 (N_18747,N_15111,N_16134);
and U18748 (N_18748,N_15349,N_15947);
or U18749 (N_18749,N_17365,N_15693);
nor U18750 (N_18750,N_16821,N_17147);
or U18751 (N_18751,N_17026,N_17227);
xor U18752 (N_18752,N_15531,N_17288);
and U18753 (N_18753,N_17332,N_15404);
or U18754 (N_18754,N_16411,N_17469);
nand U18755 (N_18755,N_17242,N_15039);
or U18756 (N_18756,N_16670,N_15813);
and U18757 (N_18757,N_16635,N_15176);
xor U18758 (N_18758,N_16273,N_15041);
and U18759 (N_18759,N_16600,N_16413);
and U18760 (N_18760,N_15340,N_15573);
xnor U18761 (N_18761,N_16287,N_17470);
and U18762 (N_18762,N_16686,N_15252);
nand U18763 (N_18763,N_16836,N_15432);
or U18764 (N_18764,N_15077,N_17060);
nor U18765 (N_18765,N_16330,N_16946);
nor U18766 (N_18766,N_15736,N_15890);
nor U18767 (N_18767,N_16941,N_16395);
nor U18768 (N_18768,N_16572,N_17204);
nand U18769 (N_18769,N_16233,N_17317);
nand U18770 (N_18770,N_16736,N_15751);
xnor U18771 (N_18771,N_17032,N_16730);
and U18772 (N_18772,N_16871,N_16348);
or U18773 (N_18773,N_16771,N_16278);
nand U18774 (N_18774,N_15930,N_15631);
and U18775 (N_18775,N_16059,N_17364);
nor U18776 (N_18776,N_16391,N_16661);
or U18777 (N_18777,N_15860,N_15938);
nor U18778 (N_18778,N_16332,N_17091);
nand U18779 (N_18779,N_16410,N_15111);
nand U18780 (N_18780,N_17297,N_15838);
nand U18781 (N_18781,N_16978,N_15824);
nand U18782 (N_18782,N_17444,N_16005);
and U18783 (N_18783,N_16903,N_16862);
and U18784 (N_18784,N_16675,N_15471);
or U18785 (N_18785,N_16379,N_17358);
nand U18786 (N_18786,N_15521,N_15460);
and U18787 (N_18787,N_17067,N_15120);
nand U18788 (N_18788,N_16532,N_15436);
xnor U18789 (N_18789,N_15137,N_15645);
nor U18790 (N_18790,N_16577,N_15179);
and U18791 (N_18791,N_16904,N_16001);
nand U18792 (N_18792,N_17002,N_15362);
nand U18793 (N_18793,N_17271,N_16612);
xor U18794 (N_18794,N_15091,N_16167);
nor U18795 (N_18795,N_15355,N_15331);
nand U18796 (N_18796,N_17159,N_15971);
and U18797 (N_18797,N_17057,N_15764);
nand U18798 (N_18798,N_17226,N_15593);
and U18799 (N_18799,N_15464,N_17285);
and U18800 (N_18800,N_16792,N_15905);
nand U18801 (N_18801,N_15567,N_15520);
nor U18802 (N_18802,N_17233,N_15740);
and U18803 (N_18803,N_15787,N_15805);
nand U18804 (N_18804,N_15331,N_17092);
or U18805 (N_18805,N_16350,N_16767);
and U18806 (N_18806,N_16639,N_15407);
or U18807 (N_18807,N_15360,N_16010);
and U18808 (N_18808,N_17209,N_15954);
xor U18809 (N_18809,N_17266,N_16502);
nand U18810 (N_18810,N_17468,N_17405);
and U18811 (N_18811,N_15648,N_15747);
or U18812 (N_18812,N_15864,N_16716);
nor U18813 (N_18813,N_15305,N_17405);
nand U18814 (N_18814,N_15676,N_16962);
nor U18815 (N_18815,N_16309,N_16797);
nand U18816 (N_18816,N_16753,N_15429);
nand U18817 (N_18817,N_17105,N_16842);
xor U18818 (N_18818,N_15759,N_16674);
or U18819 (N_18819,N_15822,N_15431);
nor U18820 (N_18820,N_15352,N_17292);
and U18821 (N_18821,N_16196,N_17373);
nor U18822 (N_18822,N_17406,N_15133);
nor U18823 (N_18823,N_15423,N_15915);
nand U18824 (N_18824,N_16123,N_17348);
and U18825 (N_18825,N_15272,N_16963);
or U18826 (N_18826,N_16285,N_16076);
and U18827 (N_18827,N_17479,N_15839);
nor U18828 (N_18828,N_15307,N_17380);
and U18829 (N_18829,N_17456,N_16364);
nand U18830 (N_18830,N_15197,N_16802);
or U18831 (N_18831,N_17198,N_15239);
and U18832 (N_18832,N_15398,N_16923);
nand U18833 (N_18833,N_15411,N_16515);
nand U18834 (N_18834,N_15125,N_17003);
nand U18835 (N_18835,N_15871,N_15684);
nand U18836 (N_18836,N_15740,N_17028);
or U18837 (N_18837,N_15149,N_15726);
xor U18838 (N_18838,N_16642,N_15202);
xor U18839 (N_18839,N_15744,N_15923);
xor U18840 (N_18840,N_16666,N_15651);
and U18841 (N_18841,N_16077,N_15515);
or U18842 (N_18842,N_16190,N_16501);
and U18843 (N_18843,N_16129,N_16282);
and U18844 (N_18844,N_16537,N_15061);
nor U18845 (N_18845,N_16245,N_17004);
xnor U18846 (N_18846,N_15008,N_15065);
and U18847 (N_18847,N_16663,N_16135);
nand U18848 (N_18848,N_16563,N_17168);
and U18849 (N_18849,N_16515,N_17172);
nor U18850 (N_18850,N_15937,N_17301);
nand U18851 (N_18851,N_16464,N_17490);
nand U18852 (N_18852,N_15574,N_16858);
nor U18853 (N_18853,N_15269,N_16631);
and U18854 (N_18854,N_15760,N_15703);
xnor U18855 (N_18855,N_15222,N_16033);
nand U18856 (N_18856,N_15241,N_17197);
xor U18857 (N_18857,N_15465,N_15469);
nand U18858 (N_18858,N_15032,N_17454);
xor U18859 (N_18859,N_15686,N_17288);
and U18860 (N_18860,N_15625,N_16583);
or U18861 (N_18861,N_16717,N_16033);
nand U18862 (N_18862,N_16993,N_16070);
xor U18863 (N_18863,N_15075,N_15216);
or U18864 (N_18864,N_16361,N_17401);
and U18865 (N_18865,N_15097,N_15143);
and U18866 (N_18866,N_16809,N_15557);
and U18867 (N_18867,N_15042,N_16823);
nand U18868 (N_18868,N_15524,N_15143);
and U18869 (N_18869,N_16068,N_16214);
nand U18870 (N_18870,N_17351,N_16381);
or U18871 (N_18871,N_17110,N_16870);
and U18872 (N_18872,N_17399,N_15514);
or U18873 (N_18873,N_17284,N_15336);
and U18874 (N_18874,N_15588,N_17414);
or U18875 (N_18875,N_15141,N_15456);
nor U18876 (N_18876,N_15796,N_16145);
nand U18877 (N_18877,N_17046,N_17195);
nor U18878 (N_18878,N_16974,N_16065);
nor U18879 (N_18879,N_17071,N_17423);
and U18880 (N_18880,N_15841,N_15366);
and U18881 (N_18881,N_16936,N_15135);
and U18882 (N_18882,N_15899,N_16386);
nor U18883 (N_18883,N_16083,N_17424);
nand U18884 (N_18884,N_15572,N_17467);
xor U18885 (N_18885,N_17088,N_15118);
or U18886 (N_18886,N_16554,N_16824);
xor U18887 (N_18887,N_15370,N_16543);
and U18888 (N_18888,N_16537,N_15847);
xor U18889 (N_18889,N_16226,N_16890);
nand U18890 (N_18890,N_15667,N_17238);
xnor U18891 (N_18891,N_16753,N_17173);
nand U18892 (N_18892,N_17145,N_16287);
nand U18893 (N_18893,N_16406,N_17368);
or U18894 (N_18894,N_17459,N_16485);
and U18895 (N_18895,N_17308,N_15446);
nand U18896 (N_18896,N_16373,N_16838);
nand U18897 (N_18897,N_17343,N_16028);
nor U18898 (N_18898,N_15017,N_15824);
xor U18899 (N_18899,N_17229,N_15134);
xor U18900 (N_18900,N_17184,N_16091);
nand U18901 (N_18901,N_17030,N_15464);
nor U18902 (N_18902,N_17446,N_15470);
nand U18903 (N_18903,N_17309,N_16660);
nand U18904 (N_18904,N_16816,N_17225);
nor U18905 (N_18905,N_15422,N_16977);
xor U18906 (N_18906,N_16660,N_15062);
nand U18907 (N_18907,N_17135,N_16965);
or U18908 (N_18908,N_15284,N_15261);
nand U18909 (N_18909,N_15866,N_15736);
and U18910 (N_18910,N_15662,N_16218);
or U18911 (N_18911,N_16921,N_16539);
xor U18912 (N_18912,N_16894,N_17100);
and U18913 (N_18913,N_17390,N_17067);
or U18914 (N_18914,N_15746,N_15018);
nor U18915 (N_18915,N_15889,N_17197);
xor U18916 (N_18916,N_15819,N_15953);
xor U18917 (N_18917,N_17033,N_16717);
xor U18918 (N_18918,N_16195,N_16043);
and U18919 (N_18919,N_16990,N_16280);
nor U18920 (N_18920,N_16024,N_15338);
or U18921 (N_18921,N_16064,N_15240);
nand U18922 (N_18922,N_15085,N_16686);
xor U18923 (N_18923,N_17094,N_17200);
or U18924 (N_18924,N_15529,N_16912);
and U18925 (N_18925,N_15064,N_15348);
nand U18926 (N_18926,N_15130,N_16489);
nor U18927 (N_18927,N_15976,N_16772);
or U18928 (N_18928,N_17344,N_15888);
or U18929 (N_18929,N_16133,N_16641);
and U18930 (N_18930,N_16620,N_15207);
xor U18931 (N_18931,N_15939,N_15121);
xnor U18932 (N_18932,N_16155,N_17231);
nor U18933 (N_18933,N_15872,N_17221);
nor U18934 (N_18934,N_15787,N_15587);
nor U18935 (N_18935,N_17358,N_16358);
and U18936 (N_18936,N_15640,N_15686);
and U18937 (N_18937,N_16288,N_17269);
or U18938 (N_18938,N_15828,N_16537);
or U18939 (N_18939,N_17488,N_15769);
nand U18940 (N_18940,N_17229,N_16248);
nor U18941 (N_18941,N_17427,N_17040);
xor U18942 (N_18942,N_16893,N_15736);
xor U18943 (N_18943,N_15848,N_15269);
nor U18944 (N_18944,N_16132,N_17155);
or U18945 (N_18945,N_16420,N_17341);
and U18946 (N_18946,N_16181,N_15642);
or U18947 (N_18947,N_15054,N_15872);
nand U18948 (N_18948,N_16402,N_16024);
xor U18949 (N_18949,N_16548,N_17495);
xor U18950 (N_18950,N_16395,N_16728);
and U18951 (N_18951,N_17331,N_15472);
or U18952 (N_18952,N_15053,N_17265);
and U18953 (N_18953,N_15672,N_16831);
nand U18954 (N_18954,N_15069,N_17008);
or U18955 (N_18955,N_17345,N_16539);
xor U18956 (N_18956,N_16255,N_15064);
xnor U18957 (N_18957,N_16293,N_15123);
xor U18958 (N_18958,N_16576,N_16462);
nor U18959 (N_18959,N_15987,N_16496);
and U18960 (N_18960,N_16125,N_17108);
xor U18961 (N_18961,N_16019,N_15108);
nor U18962 (N_18962,N_17223,N_16705);
or U18963 (N_18963,N_17169,N_16907);
nand U18964 (N_18964,N_15123,N_16556);
or U18965 (N_18965,N_15265,N_16286);
nand U18966 (N_18966,N_15747,N_16508);
and U18967 (N_18967,N_17357,N_16135);
xnor U18968 (N_18968,N_16053,N_17108);
and U18969 (N_18969,N_15773,N_16416);
and U18970 (N_18970,N_15305,N_15145);
xnor U18971 (N_18971,N_15173,N_16907);
nor U18972 (N_18972,N_16737,N_17205);
nand U18973 (N_18973,N_15988,N_15396);
nor U18974 (N_18974,N_17330,N_17464);
or U18975 (N_18975,N_15164,N_17309);
and U18976 (N_18976,N_15473,N_15922);
nor U18977 (N_18977,N_17450,N_15673);
and U18978 (N_18978,N_15077,N_16290);
xnor U18979 (N_18979,N_16069,N_17462);
or U18980 (N_18980,N_16651,N_16878);
or U18981 (N_18981,N_15529,N_15347);
and U18982 (N_18982,N_16632,N_15324);
and U18983 (N_18983,N_15823,N_16608);
and U18984 (N_18984,N_17463,N_15050);
nor U18985 (N_18985,N_16166,N_15554);
and U18986 (N_18986,N_16106,N_15661);
nand U18987 (N_18987,N_16609,N_16156);
nand U18988 (N_18988,N_15795,N_15453);
and U18989 (N_18989,N_16497,N_16113);
and U18990 (N_18990,N_16957,N_16249);
and U18991 (N_18991,N_15897,N_15943);
and U18992 (N_18992,N_17266,N_16518);
or U18993 (N_18993,N_16319,N_16410);
and U18994 (N_18994,N_15449,N_16359);
xnor U18995 (N_18995,N_15922,N_16756);
nand U18996 (N_18996,N_17172,N_15674);
xnor U18997 (N_18997,N_15853,N_16907);
or U18998 (N_18998,N_17230,N_16106);
xor U18999 (N_18999,N_15464,N_15637);
xor U19000 (N_19000,N_15661,N_17178);
and U19001 (N_19001,N_16257,N_15761);
xnor U19002 (N_19002,N_15979,N_15499);
xnor U19003 (N_19003,N_15772,N_16155);
nand U19004 (N_19004,N_15961,N_17141);
xnor U19005 (N_19005,N_16828,N_15574);
or U19006 (N_19006,N_17312,N_15543);
and U19007 (N_19007,N_15486,N_16779);
and U19008 (N_19008,N_16635,N_16655);
or U19009 (N_19009,N_16314,N_17091);
or U19010 (N_19010,N_15689,N_15985);
and U19011 (N_19011,N_16878,N_16650);
nor U19012 (N_19012,N_16691,N_16879);
nor U19013 (N_19013,N_16969,N_15801);
nand U19014 (N_19014,N_16015,N_17273);
nor U19015 (N_19015,N_17403,N_15951);
nand U19016 (N_19016,N_16821,N_16126);
nand U19017 (N_19017,N_17474,N_17219);
nand U19018 (N_19018,N_15608,N_15491);
xor U19019 (N_19019,N_17008,N_15848);
and U19020 (N_19020,N_17169,N_16526);
xor U19021 (N_19021,N_16601,N_16029);
xor U19022 (N_19022,N_15853,N_17454);
nand U19023 (N_19023,N_15431,N_15771);
nor U19024 (N_19024,N_15405,N_15733);
nand U19025 (N_19025,N_15202,N_15523);
xnor U19026 (N_19026,N_16168,N_15235);
nand U19027 (N_19027,N_15318,N_16445);
nor U19028 (N_19028,N_16284,N_15199);
and U19029 (N_19029,N_16969,N_15519);
and U19030 (N_19030,N_16017,N_16294);
and U19031 (N_19031,N_17422,N_16849);
xnor U19032 (N_19032,N_15952,N_15942);
xor U19033 (N_19033,N_17274,N_16089);
xor U19034 (N_19034,N_17436,N_16883);
nor U19035 (N_19035,N_15043,N_17423);
xor U19036 (N_19036,N_17346,N_17285);
nor U19037 (N_19037,N_15992,N_16267);
and U19038 (N_19038,N_15364,N_17124);
xnor U19039 (N_19039,N_16455,N_15465);
nor U19040 (N_19040,N_16781,N_17250);
or U19041 (N_19041,N_16468,N_17186);
and U19042 (N_19042,N_15793,N_17223);
and U19043 (N_19043,N_17381,N_15909);
nand U19044 (N_19044,N_15210,N_17324);
or U19045 (N_19045,N_16359,N_17369);
nand U19046 (N_19046,N_16246,N_16338);
nor U19047 (N_19047,N_16109,N_16387);
nor U19048 (N_19048,N_16963,N_16388);
xnor U19049 (N_19049,N_17437,N_15558);
and U19050 (N_19050,N_15819,N_15751);
xnor U19051 (N_19051,N_16847,N_17215);
xor U19052 (N_19052,N_16588,N_15443);
or U19053 (N_19053,N_16158,N_16495);
nor U19054 (N_19054,N_15565,N_16373);
and U19055 (N_19055,N_15724,N_17302);
xnor U19056 (N_19056,N_17178,N_17459);
or U19057 (N_19057,N_16260,N_15457);
and U19058 (N_19058,N_16829,N_16852);
nor U19059 (N_19059,N_17244,N_17329);
nor U19060 (N_19060,N_15401,N_16997);
nor U19061 (N_19061,N_16732,N_15753);
nand U19062 (N_19062,N_17454,N_16976);
and U19063 (N_19063,N_15834,N_17227);
and U19064 (N_19064,N_16001,N_16568);
nor U19065 (N_19065,N_16156,N_16010);
and U19066 (N_19066,N_15063,N_16644);
nand U19067 (N_19067,N_16933,N_16230);
xor U19068 (N_19068,N_16061,N_15665);
and U19069 (N_19069,N_16895,N_16432);
and U19070 (N_19070,N_16306,N_15637);
nor U19071 (N_19071,N_16452,N_15023);
nor U19072 (N_19072,N_16677,N_17034);
nand U19073 (N_19073,N_17072,N_17057);
and U19074 (N_19074,N_17305,N_16490);
xnor U19075 (N_19075,N_16824,N_17298);
nand U19076 (N_19076,N_17403,N_16610);
or U19077 (N_19077,N_15243,N_16442);
nor U19078 (N_19078,N_16373,N_16875);
and U19079 (N_19079,N_15093,N_16708);
xnor U19080 (N_19080,N_16908,N_15269);
nand U19081 (N_19081,N_15895,N_16607);
and U19082 (N_19082,N_16887,N_15885);
or U19083 (N_19083,N_17025,N_17235);
or U19084 (N_19084,N_15685,N_15948);
or U19085 (N_19085,N_17090,N_16645);
nand U19086 (N_19086,N_16212,N_17175);
nand U19087 (N_19087,N_16534,N_15739);
nor U19088 (N_19088,N_16369,N_15709);
xor U19089 (N_19089,N_15127,N_17379);
and U19090 (N_19090,N_15647,N_15642);
nor U19091 (N_19091,N_16162,N_16092);
xor U19092 (N_19092,N_15641,N_15169);
xor U19093 (N_19093,N_17313,N_15349);
and U19094 (N_19094,N_15661,N_15796);
nand U19095 (N_19095,N_15075,N_16488);
xnor U19096 (N_19096,N_17116,N_17307);
and U19097 (N_19097,N_17420,N_17397);
xnor U19098 (N_19098,N_16944,N_15512);
or U19099 (N_19099,N_15548,N_16564);
xnor U19100 (N_19100,N_16442,N_15360);
nor U19101 (N_19101,N_16693,N_15451);
nor U19102 (N_19102,N_15829,N_15140);
xor U19103 (N_19103,N_17083,N_17160);
xnor U19104 (N_19104,N_16232,N_16462);
xnor U19105 (N_19105,N_16072,N_15680);
and U19106 (N_19106,N_16236,N_15492);
or U19107 (N_19107,N_15422,N_17124);
nand U19108 (N_19108,N_15897,N_15759);
or U19109 (N_19109,N_16323,N_17277);
nand U19110 (N_19110,N_15150,N_16378);
xor U19111 (N_19111,N_17288,N_16199);
xor U19112 (N_19112,N_16765,N_17275);
and U19113 (N_19113,N_16856,N_17071);
or U19114 (N_19114,N_15063,N_15413);
nand U19115 (N_19115,N_15202,N_15409);
nand U19116 (N_19116,N_15737,N_17484);
nor U19117 (N_19117,N_16174,N_15247);
nand U19118 (N_19118,N_17246,N_16536);
nand U19119 (N_19119,N_15114,N_15169);
and U19120 (N_19120,N_17434,N_16581);
nand U19121 (N_19121,N_15530,N_15127);
or U19122 (N_19122,N_15404,N_15265);
and U19123 (N_19123,N_15012,N_17116);
nand U19124 (N_19124,N_16887,N_15177);
nand U19125 (N_19125,N_16613,N_15018);
and U19126 (N_19126,N_15375,N_17297);
xnor U19127 (N_19127,N_17419,N_16533);
xor U19128 (N_19128,N_16803,N_15016);
or U19129 (N_19129,N_15829,N_16949);
nor U19130 (N_19130,N_16121,N_16194);
nand U19131 (N_19131,N_16411,N_17324);
nand U19132 (N_19132,N_15405,N_16337);
or U19133 (N_19133,N_16877,N_15052);
xnor U19134 (N_19134,N_16554,N_15255);
nor U19135 (N_19135,N_16165,N_16632);
xnor U19136 (N_19136,N_15211,N_17178);
nand U19137 (N_19137,N_17430,N_15469);
nand U19138 (N_19138,N_15940,N_16290);
nand U19139 (N_19139,N_15096,N_16264);
nor U19140 (N_19140,N_17473,N_17114);
or U19141 (N_19141,N_17329,N_16701);
xor U19142 (N_19142,N_16048,N_16973);
or U19143 (N_19143,N_15470,N_16994);
nor U19144 (N_19144,N_15106,N_15112);
and U19145 (N_19145,N_16773,N_16069);
xor U19146 (N_19146,N_15133,N_16221);
and U19147 (N_19147,N_16801,N_16898);
nand U19148 (N_19148,N_16500,N_15630);
or U19149 (N_19149,N_16709,N_16234);
nand U19150 (N_19150,N_16949,N_17412);
nor U19151 (N_19151,N_15472,N_16284);
nand U19152 (N_19152,N_15489,N_16562);
or U19153 (N_19153,N_15582,N_15373);
nor U19154 (N_19154,N_17064,N_16601);
nand U19155 (N_19155,N_16710,N_16668);
or U19156 (N_19156,N_15215,N_15660);
nor U19157 (N_19157,N_15644,N_16406);
and U19158 (N_19158,N_16313,N_15630);
and U19159 (N_19159,N_16245,N_16201);
xor U19160 (N_19160,N_17062,N_16641);
nor U19161 (N_19161,N_16833,N_16306);
xnor U19162 (N_19162,N_15785,N_16071);
nand U19163 (N_19163,N_16181,N_15019);
or U19164 (N_19164,N_15415,N_16353);
xnor U19165 (N_19165,N_15876,N_16851);
and U19166 (N_19166,N_17129,N_16001);
nand U19167 (N_19167,N_15307,N_17395);
nand U19168 (N_19168,N_16713,N_15119);
and U19169 (N_19169,N_15053,N_15860);
xnor U19170 (N_19170,N_15543,N_17319);
nor U19171 (N_19171,N_15002,N_17468);
and U19172 (N_19172,N_16491,N_16962);
xnor U19173 (N_19173,N_15699,N_15408);
nor U19174 (N_19174,N_16125,N_17004);
nor U19175 (N_19175,N_17201,N_16018);
nand U19176 (N_19176,N_15598,N_16652);
nor U19177 (N_19177,N_15939,N_15492);
or U19178 (N_19178,N_15831,N_17493);
nand U19179 (N_19179,N_17392,N_16203);
nand U19180 (N_19180,N_17034,N_16239);
or U19181 (N_19181,N_17039,N_17334);
nor U19182 (N_19182,N_15168,N_17085);
and U19183 (N_19183,N_16353,N_17170);
and U19184 (N_19184,N_15105,N_15452);
xor U19185 (N_19185,N_15414,N_16387);
or U19186 (N_19186,N_15571,N_15087);
nand U19187 (N_19187,N_15974,N_15624);
and U19188 (N_19188,N_15386,N_17363);
nor U19189 (N_19189,N_15308,N_15405);
nand U19190 (N_19190,N_15860,N_16525);
nor U19191 (N_19191,N_15043,N_16994);
nor U19192 (N_19192,N_15868,N_16882);
or U19193 (N_19193,N_16505,N_16138);
and U19194 (N_19194,N_16801,N_15061);
nand U19195 (N_19195,N_17425,N_15838);
xor U19196 (N_19196,N_15350,N_16233);
nand U19197 (N_19197,N_16725,N_17466);
and U19198 (N_19198,N_15643,N_15690);
nor U19199 (N_19199,N_15725,N_15647);
nand U19200 (N_19200,N_16535,N_16140);
xnor U19201 (N_19201,N_17058,N_17192);
and U19202 (N_19202,N_16249,N_15862);
or U19203 (N_19203,N_17111,N_17279);
xnor U19204 (N_19204,N_15509,N_17060);
xnor U19205 (N_19205,N_16057,N_16232);
nor U19206 (N_19206,N_17283,N_17250);
and U19207 (N_19207,N_15121,N_15777);
nor U19208 (N_19208,N_15694,N_16907);
or U19209 (N_19209,N_15339,N_15220);
nor U19210 (N_19210,N_17197,N_16149);
xor U19211 (N_19211,N_16326,N_16697);
nand U19212 (N_19212,N_15501,N_16782);
nor U19213 (N_19213,N_17071,N_15416);
and U19214 (N_19214,N_16344,N_15034);
xor U19215 (N_19215,N_15148,N_16678);
nor U19216 (N_19216,N_16130,N_17213);
and U19217 (N_19217,N_16195,N_15211);
nor U19218 (N_19218,N_15704,N_15255);
or U19219 (N_19219,N_15498,N_15844);
nor U19220 (N_19220,N_15339,N_16895);
nor U19221 (N_19221,N_15035,N_16325);
and U19222 (N_19222,N_16894,N_15710);
nand U19223 (N_19223,N_15016,N_17472);
or U19224 (N_19224,N_15361,N_15778);
nand U19225 (N_19225,N_15501,N_16948);
and U19226 (N_19226,N_16371,N_16511);
and U19227 (N_19227,N_15027,N_17346);
nand U19228 (N_19228,N_17005,N_15372);
xnor U19229 (N_19229,N_16280,N_16023);
or U19230 (N_19230,N_16730,N_16921);
xnor U19231 (N_19231,N_16413,N_15753);
nor U19232 (N_19232,N_16020,N_15840);
nand U19233 (N_19233,N_15784,N_17316);
or U19234 (N_19234,N_16562,N_15220);
or U19235 (N_19235,N_15732,N_16381);
nand U19236 (N_19236,N_17151,N_15983);
and U19237 (N_19237,N_15708,N_15894);
and U19238 (N_19238,N_17247,N_16034);
xor U19239 (N_19239,N_17478,N_16985);
and U19240 (N_19240,N_16411,N_15705);
nor U19241 (N_19241,N_15808,N_17026);
or U19242 (N_19242,N_15353,N_16075);
nand U19243 (N_19243,N_15283,N_17116);
and U19244 (N_19244,N_17291,N_15744);
or U19245 (N_19245,N_15017,N_15292);
nand U19246 (N_19246,N_16707,N_15231);
and U19247 (N_19247,N_17271,N_17337);
and U19248 (N_19248,N_17229,N_16907);
nor U19249 (N_19249,N_16783,N_15000);
and U19250 (N_19250,N_17353,N_16522);
nor U19251 (N_19251,N_15416,N_15484);
or U19252 (N_19252,N_17264,N_15601);
or U19253 (N_19253,N_17177,N_16889);
xnor U19254 (N_19254,N_15082,N_16476);
nand U19255 (N_19255,N_15736,N_16934);
xor U19256 (N_19256,N_17351,N_17476);
and U19257 (N_19257,N_15489,N_16840);
or U19258 (N_19258,N_15813,N_15387);
nor U19259 (N_19259,N_16130,N_17357);
and U19260 (N_19260,N_16192,N_17429);
nor U19261 (N_19261,N_15510,N_16680);
xor U19262 (N_19262,N_15774,N_16518);
nand U19263 (N_19263,N_15365,N_17289);
or U19264 (N_19264,N_16115,N_16711);
nand U19265 (N_19265,N_15197,N_17367);
xor U19266 (N_19266,N_15384,N_17101);
xnor U19267 (N_19267,N_16067,N_16421);
or U19268 (N_19268,N_15342,N_17079);
or U19269 (N_19269,N_15953,N_15214);
and U19270 (N_19270,N_17304,N_17128);
and U19271 (N_19271,N_15635,N_16472);
nor U19272 (N_19272,N_15251,N_17458);
or U19273 (N_19273,N_16255,N_15859);
nor U19274 (N_19274,N_15393,N_16209);
and U19275 (N_19275,N_16290,N_16432);
or U19276 (N_19276,N_15783,N_16095);
nand U19277 (N_19277,N_16616,N_15667);
or U19278 (N_19278,N_16013,N_17468);
xor U19279 (N_19279,N_16094,N_15487);
nor U19280 (N_19280,N_15254,N_16267);
or U19281 (N_19281,N_16899,N_16125);
nand U19282 (N_19282,N_17001,N_15494);
xor U19283 (N_19283,N_16132,N_16553);
xor U19284 (N_19284,N_17273,N_15416);
and U19285 (N_19285,N_16933,N_16326);
nand U19286 (N_19286,N_17471,N_15898);
and U19287 (N_19287,N_16875,N_15019);
and U19288 (N_19288,N_16498,N_17019);
nor U19289 (N_19289,N_17251,N_17344);
nand U19290 (N_19290,N_16758,N_15258);
nor U19291 (N_19291,N_17154,N_15952);
xor U19292 (N_19292,N_17275,N_17370);
and U19293 (N_19293,N_17378,N_16816);
and U19294 (N_19294,N_17363,N_15374);
xnor U19295 (N_19295,N_16865,N_15963);
or U19296 (N_19296,N_16208,N_15479);
nor U19297 (N_19297,N_16935,N_17171);
nand U19298 (N_19298,N_15781,N_17189);
nor U19299 (N_19299,N_17127,N_16696);
nand U19300 (N_19300,N_17242,N_16508);
nand U19301 (N_19301,N_15878,N_15080);
nand U19302 (N_19302,N_15958,N_16125);
nand U19303 (N_19303,N_15391,N_17153);
nor U19304 (N_19304,N_16696,N_16551);
and U19305 (N_19305,N_15869,N_16821);
or U19306 (N_19306,N_17369,N_17015);
nand U19307 (N_19307,N_17180,N_16260);
and U19308 (N_19308,N_16921,N_15821);
or U19309 (N_19309,N_16500,N_17024);
nor U19310 (N_19310,N_17185,N_15306);
nor U19311 (N_19311,N_17368,N_15417);
nand U19312 (N_19312,N_15470,N_15532);
and U19313 (N_19313,N_16728,N_16767);
and U19314 (N_19314,N_15216,N_15806);
nand U19315 (N_19315,N_16913,N_15926);
and U19316 (N_19316,N_17143,N_15844);
xor U19317 (N_19317,N_16758,N_15791);
nor U19318 (N_19318,N_16732,N_17483);
and U19319 (N_19319,N_16034,N_15442);
and U19320 (N_19320,N_15469,N_15139);
xnor U19321 (N_19321,N_16994,N_15244);
nand U19322 (N_19322,N_15040,N_17159);
and U19323 (N_19323,N_17263,N_17410);
or U19324 (N_19324,N_16107,N_17411);
xnor U19325 (N_19325,N_16051,N_16020);
or U19326 (N_19326,N_15878,N_15926);
and U19327 (N_19327,N_17403,N_16261);
and U19328 (N_19328,N_16626,N_15525);
nand U19329 (N_19329,N_17490,N_15191);
nand U19330 (N_19330,N_17467,N_16910);
nand U19331 (N_19331,N_16284,N_15825);
and U19332 (N_19332,N_16992,N_15393);
nor U19333 (N_19333,N_16204,N_15537);
nand U19334 (N_19334,N_16225,N_16152);
xnor U19335 (N_19335,N_15870,N_16124);
nor U19336 (N_19336,N_16332,N_15651);
nor U19337 (N_19337,N_16660,N_16562);
or U19338 (N_19338,N_16819,N_17004);
or U19339 (N_19339,N_15327,N_15981);
nor U19340 (N_19340,N_16230,N_15755);
and U19341 (N_19341,N_15594,N_16236);
nand U19342 (N_19342,N_15482,N_16133);
or U19343 (N_19343,N_15776,N_17191);
xor U19344 (N_19344,N_15360,N_17315);
nor U19345 (N_19345,N_15103,N_15204);
and U19346 (N_19346,N_15523,N_16147);
and U19347 (N_19347,N_15038,N_16698);
nand U19348 (N_19348,N_17026,N_17261);
nand U19349 (N_19349,N_16333,N_17303);
xnor U19350 (N_19350,N_16325,N_17464);
xnor U19351 (N_19351,N_17020,N_16399);
nand U19352 (N_19352,N_16718,N_15709);
nand U19353 (N_19353,N_16379,N_17281);
and U19354 (N_19354,N_15524,N_15777);
and U19355 (N_19355,N_16425,N_16546);
and U19356 (N_19356,N_17366,N_16366);
xor U19357 (N_19357,N_15358,N_16778);
xor U19358 (N_19358,N_16003,N_15987);
xor U19359 (N_19359,N_15871,N_16509);
xor U19360 (N_19360,N_15326,N_15886);
or U19361 (N_19361,N_17170,N_16890);
and U19362 (N_19362,N_15211,N_15297);
xor U19363 (N_19363,N_16980,N_16048);
xor U19364 (N_19364,N_15763,N_17193);
xnor U19365 (N_19365,N_16758,N_16461);
and U19366 (N_19366,N_15503,N_16789);
and U19367 (N_19367,N_15724,N_16723);
or U19368 (N_19368,N_17006,N_17218);
and U19369 (N_19369,N_15164,N_15542);
nand U19370 (N_19370,N_15625,N_17250);
nor U19371 (N_19371,N_17365,N_15663);
and U19372 (N_19372,N_16674,N_15821);
xor U19373 (N_19373,N_17218,N_16619);
or U19374 (N_19374,N_16631,N_16752);
nand U19375 (N_19375,N_15253,N_15357);
nand U19376 (N_19376,N_17346,N_16705);
nand U19377 (N_19377,N_15906,N_17276);
nand U19378 (N_19378,N_17467,N_17024);
xor U19379 (N_19379,N_16019,N_15975);
nor U19380 (N_19380,N_15862,N_15564);
or U19381 (N_19381,N_16620,N_16334);
xor U19382 (N_19382,N_17210,N_15719);
xnor U19383 (N_19383,N_17051,N_16477);
nand U19384 (N_19384,N_15489,N_15055);
nand U19385 (N_19385,N_16439,N_15355);
nor U19386 (N_19386,N_17319,N_15621);
nor U19387 (N_19387,N_15142,N_16469);
xnor U19388 (N_19388,N_15802,N_15069);
nor U19389 (N_19389,N_15699,N_15213);
and U19390 (N_19390,N_15303,N_16985);
nand U19391 (N_19391,N_15897,N_17431);
or U19392 (N_19392,N_17171,N_17200);
nor U19393 (N_19393,N_15755,N_17101);
or U19394 (N_19394,N_15319,N_15180);
and U19395 (N_19395,N_16719,N_17451);
or U19396 (N_19396,N_15464,N_15531);
and U19397 (N_19397,N_16045,N_15208);
nor U19398 (N_19398,N_15576,N_15093);
or U19399 (N_19399,N_16742,N_16068);
or U19400 (N_19400,N_16725,N_16747);
nand U19401 (N_19401,N_16924,N_16249);
xnor U19402 (N_19402,N_15003,N_16266);
nor U19403 (N_19403,N_16383,N_15798);
nand U19404 (N_19404,N_15084,N_15181);
nand U19405 (N_19405,N_15229,N_16342);
xnor U19406 (N_19406,N_15104,N_16242);
nand U19407 (N_19407,N_15726,N_15326);
or U19408 (N_19408,N_15516,N_15081);
nor U19409 (N_19409,N_17459,N_15013);
or U19410 (N_19410,N_15364,N_17156);
xor U19411 (N_19411,N_17415,N_15043);
and U19412 (N_19412,N_17085,N_16593);
nor U19413 (N_19413,N_17193,N_15734);
nand U19414 (N_19414,N_17235,N_17385);
or U19415 (N_19415,N_15314,N_17336);
or U19416 (N_19416,N_15133,N_16597);
nor U19417 (N_19417,N_16131,N_15392);
xor U19418 (N_19418,N_17366,N_16669);
nand U19419 (N_19419,N_15244,N_17325);
nor U19420 (N_19420,N_16562,N_16684);
and U19421 (N_19421,N_15928,N_15665);
and U19422 (N_19422,N_17104,N_16664);
xnor U19423 (N_19423,N_16391,N_15258);
xor U19424 (N_19424,N_15856,N_17013);
or U19425 (N_19425,N_16547,N_16798);
and U19426 (N_19426,N_16412,N_15604);
or U19427 (N_19427,N_15322,N_17317);
and U19428 (N_19428,N_16931,N_15682);
nor U19429 (N_19429,N_15905,N_16837);
nor U19430 (N_19430,N_15790,N_15147);
xnor U19431 (N_19431,N_15951,N_16390);
xor U19432 (N_19432,N_16578,N_15724);
nand U19433 (N_19433,N_15124,N_15848);
nor U19434 (N_19434,N_17058,N_16930);
nand U19435 (N_19435,N_16717,N_16268);
nand U19436 (N_19436,N_15228,N_16093);
and U19437 (N_19437,N_15748,N_16286);
or U19438 (N_19438,N_16606,N_16164);
nor U19439 (N_19439,N_16136,N_15293);
xnor U19440 (N_19440,N_17252,N_15385);
xnor U19441 (N_19441,N_15684,N_15420);
nand U19442 (N_19442,N_16415,N_16549);
nor U19443 (N_19443,N_17056,N_16979);
or U19444 (N_19444,N_16532,N_15332);
nor U19445 (N_19445,N_16573,N_16176);
xnor U19446 (N_19446,N_15196,N_16739);
or U19447 (N_19447,N_15104,N_17445);
nand U19448 (N_19448,N_16463,N_17444);
xnor U19449 (N_19449,N_16869,N_15318);
and U19450 (N_19450,N_16379,N_17301);
or U19451 (N_19451,N_16542,N_15215);
nor U19452 (N_19452,N_15164,N_16948);
and U19453 (N_19453,N_16153,N_16080);
xor U19454 (N_19454,N_16563,N_16655);
nor U19455 (N_19455,N_15837,N_15377);
nand U19456 (N_19456,N_16869,N_17281);
or U19457 (N_19457,N_17151,N_16619);
and U19458 (N_19458,N_15038,N_16339);
nor U19459 (N_19459,N_15113,N_17132);
or U19460 (N_19460,N_16811,N_16704);
xor U19461 (N_19461,N_16187,N_15213);
nor U19462 (N_19462,N_15677,N_15234);
nand U19463 (N_19463,N_17111,N_15837);
or U19464 (N_19464,N_17469,N_15856);
and U19465 (N_19465,N_17295,N_16616);
xor U19466 (N_19466,N_17385,N_16627);
nor U19467 (N_19467,N_15005,N_16600);
nand U19468 (N_19468,N_16986,N_17288);
nor U19469 (N_19469,N_16183,N_15265);
nand U19470 (N_19470,N_17488,N_16656);
and U19471 (N_19471,N_17480,N_15582);
and U19472 (N_19472,N_15427,N_17073);
nand U19473 (N_19473,N_16207,N_16371);
xnor U19474 (N_19474,N_15883,N_15561);
or U19475 (N_19475,N_16957,N_16544);
nand U19476 (N_19476,N_16045,N_16186);
or U19477 (N_19477,N_17248,N_16838);
xor U19478 (N_19478,N_17300,N_17253);
nand U19479 (N_19479,N_17093,N_16114);
and U19480 (N_19480,N_16959,N_17048);
xor U19481 (N_19481,N_15991,N_16248);
and U19482 (N_19482,N_15938,N_16590);
nand U19483 (N_19483,N_15535,N_17450);
xnor U19484 (N_19484,N_15568,N_16229);
and U19485 (N_19485,N_16529,N_15708);
nor U19486 (N_19486,N_15292,N_15010);
and U19487 (N_19487,N_16521,N_15499);
xor U19488 (N_19488,N_15500,N_15822);
xnor U19489 (N_19489,N_16758,N_17374);
nor U19490 (N_19490,N_15960,N_17212);
xor U19491 (N_19491,N_17186,N_16024);
nand U19492 (N_19492,N_16426,N_15563);
or U19493 (N_19493,N_17339,N_17398);
xnor U19494 (N_19494,N_15271,N_15047);
or U19495 (N_19495,N_15085,N_15277);
xor U19496 (N_19496,N_15573,N_16879);
nor U19497 (N_19497,N_16343,N_15909);
nor U19498 (N_19498,N_17226,N_15872);
or U19499 (N_19499,N_16825,N_15394);
nor U19500 (N_19500,N_15615,N_15750);
xnor U19501 (N_19501,N_15925,N_17309);
and U19502 (N_19502,N_17336,N_17029);
xnor U19503 (N_19503,N_16746,N_16068);
or U19504 (N_19504,N_15583,N_17000);
nand U19505 (N_19505,N_16965,N_16497);
nand U19506 (N_19506,N_16855,N_15079);
nand U19507 (N_19507,N_15303,N_15378);
or U19508 (N_19508,N_16166,N_16500);
nor U19509 (N_19509,N_15090,N_16150);
nand U19510 (N_19510,N_15501,N_17284);
nand U19511 (N_19511,N_15486,N_15688);
and U19512 (N_19512,N_15658,N_15778);
xor U19513 (N_19513,N_17353,N_16365);
xor U19514 (N_19514,N_15749,N_17477);
and U19515 (N_19515,N_15855,N_15255);
nand U19516 (N_19516,N_16556,N_16438);
and U19517 (N_19517,N_15896,N_15510);
xor U19518 (N_19518,N_16785,N_15557);
nand U19519 (N_19519,N_15201,N_15783);
and U19520 (N_19520,N_17217,N_15580);
nand U19521 (N_19521,N_16923,N_16581);
nand U19522 (N_19522,N_16038,N_15272);
or U19523 (N_19523,N_16609,N_15168);
and U19524 (N_19524,N_16682,N_15972);
nand U19525 (N_19525,N_15642,N_15333);
or U19526 (N_19526,N_15027,N_15982);
and U19527 (N_19527,N_15472,N_16535);
or U19528 (N_19528,N_16464,N_17498);
and U19529 (N_19529,N_16799,N_17273);
and U19530 (N_19530,N_15069,N_17410);
nor U19531 (N_19531,N_17032,N_17196);
xor U19532 (N_19532,N_15788,N_15715);
nor U19533 (N_19533,N_17071,N_16278);
nor U19534 (N_19534,N_16256,N_15379);
nor U19535 (N_19535,N_17487,N_15259);
nor U19536 (N_19536,N_15468,N_15240);
xor U19537 (N_19537,N_17149,N_16189);
xor U19538 (N_19538,N_15823,N_15491);
and U19539 (N_19539,N_15584,N_17274);
xnor U19540 (N_19540,N_15404,N_16985);
nor U19541 (N_19541,N_15348,N_16073);
nand U19542 (N_19542,N_17121,N_15345);
xor U19543 (N_19543,N_15436,N_15348);
nor U19544 (N_19544,N_15803,N_15391);
and U19545 (N_19545,N_17346,N_15514);
xor U19546 (N_19546,N_16456,N_15941);
or U19547 (N_19547,N_16794,N_15812);
nand U19548 (N_19548,N_17183,N_15303);
or U19549 (N_19549,N_15354,N_15733);
and U19550 (N_19550,N_15452,N_15309);
or U19551 (N_19551,N_16758,N_15000);
and U19552 (N_19552,N_16310,N_17110);
or U19553 (N_19553,N_16747,N_17372);
nor U19554 (N_19554,N_16483,N_16927);
or U19555 (N_19555,N_15015,N_17471);
nor U19556 (N_19556,N_15904,N_16440);
or U19557 (N_19557,N_16427,N_15628);
or U19558 (N_19558,N_15319,N_17103);
nand U19559 (N_19559,N_17229,N_15126);
nor U19560 (N_19560,N_15351,N_15056);
xor U19561 (N_19561,N_17145,N_17046);
and U19562 (N_19562,N_17255,N_17421);
nor U19563 (N_19563,N_16340,N_17176);
or U19564 (N_19564,N_15120,N_15897);
nor U19565 (N_19565,N_15188,N_15670);
nand U19566 (N_19566,N_15047,N_17158);
nor U19567 (N_19567,N_16009,N_15407);
nor U19568 (N_19568,N_15380,N_16778);
and U19569 (N_19569,N_15322,N_16555);
or U19570 (N_19570,N_16332,N_16323);
nor U19571 (N_19571,N_15662,N_17425);
nor U19572 (N_19572,N_15461,N_15152);
nor U19573 (N_19573,N_16424,N_16619);
or U19574 (N_19574,N_15761,N_15577);
xnor U19575 (N_19575,N_16017,N_16106);
xor U19576 (N_19576,N_16883,N_15571);
nor U19577 (N_19577,N_17142,N_15923);
xor U19578 (N_19578,N_17038,N_16678);
or U19579 (N_19579,N_15784,N_17034);
nor U19580 (N_19580,N_17108,N_16270);
xor U19581 (N_19581,N_15016,N_16740);
nand U19582 (N_19582,N_17476,N_15473);
or U19583 (N_19583,N_17097,N_16128);
and U19584 (N_19584,N_15510,N_16960);
or U19585 (N_19585,N_15878,N_15460);
nor U19586 (N_19586,N_15171,N_16941);
and U19587 (N_19587,N_15302,N_17174);
and U19588 (N_19588,N_17027,N_16567);
and U19589 (N_19589,N_15064,N_16312);
and U19590 (N_19590,N_15835,N_17208);
and U19591 (N_19591,N_15305,N_15998);
or U19592 (N_19592,N_15507,N_16111);
and U19593 (N_19593,N_15135,N_15005);
xnor U19594 (N_19594,N_16026,N_16127);
nand U19595 (N_19595,N_16484,N_16324);
xor U19596 (N_19596,N_15551,N_16810);
xor U19597 (N_19597,N_15338,N_17130);
or U19598 (N_19598,N_16843,N_17157);
nand U19599 (N_19599,N_15884,N_16504);
or U19600 (N_19600,N_16762,N_15366);
and U19601 (N_19601,N_16098,N_17457);
or U19602 (N_19602,N_16374,N_15659);
or U19603 (N_19603,N_15379,N_15489);
xor U19604 (N_19604,N_15943,N_15864);
nor U19605 (N_19605,N_16468,N_16705);
or U19606 (N_19606,N_15618,N_17148);
or U19607 (N_19607,N_17082,N_17378);
nor U19608 (N_19608,N_17234,N_17411);
or U19609 (N_19609,N_15370,N_15911);
nand U19610 (N_19610,N_16583,N_17162);
nor U19611 (N_19611,N_16962,N_16421);
or U19612 (N_19612,N_16784,N_15549);
nand U19613 (N_19613,N_16716,N_15027);
nor U19614 (N_19614,N_16446,N_15192);
nor U19615 (N_19615,N_16908,N_15169);
and U19616 (N_19616,N_15947,N_15564);
or U19617 (N_19617,N_17472,N_15343);
and U19618 (N_19618,N_16982,N_16968);
nor U19619 (N_19619,N_17315,N_16940);
xor U19620 (N_19620,N_16587,N_16719);
xnor U19621 (N_19621,N_15109,N_17395);
nand U19622 (N_19622,N_16371,N_16841);
xnor U19623 (N_19623,N_16525,N_16195);
nand U19624 (N_19624,N_16819,N_17345);
nand U19625 (N_19625,N_16943,N_17115);
xnor U19626 (N_19626,N_16200,N_17048);
and U19627 (N_19627,N_15487,N_15917);
and U19628 (N_19628,N_16199,N_17127);
or U19629 (N_19629,N_16001,N_16378);
nand U19630 (N_19630,N_16932,N_15267);
or U19631 (N_19631,N_15758,N_16196);
or U19632 (N_19632,N_17315,N_16263);
nand U19633 (N_19633,N_17310,N_16618);
xor U19634 (N_19634,N_16965,N_17427);
nor U19635 (N_19635,N_16544,N_15891);
nand U19636 (N_19636,N_17488,N_16440);
nor U19637 (N_19637,N_16970,N_17389);
nand U19638 (N_19638,N_16957,N_16936);
nor U19639 (N_19639,N_17453,N_16170);
xor U19640 (N_19640,N_17207,N_16711);
nor U19641 (N_19641,N_16067,N_17208);
nor U19642 (N_19642,N_15396,N_17108);
nor U19643 (N_19643,N_16091,N_16195);
nand U19644 (N_19644,N_15976,N_16054);
nand U19645 (N_19645,N_15624,N_17363);
or U19646 (N_19646,N_16184,N_15093);
or U19647 (N_19647,N_15475,N_15287);
nand U19648 (N_19648,N_15894,N_15400);
or U19649 (N_19649,N_15532,N_16626);
or U19650 (N_19650,N_17200,N_15845);
and U19651 (N_19651,N_17197,N_17423);
nor U19652 (N_19652,N_16512,N_16010);
or U19653 (N_19653,N_15619,N_16059);
nor U19654 (N_19654,N_17221,N_16099);
nand U19655 (N_19655,N_16585,N_16641);
and U19656 (N_19656,N_16107,N_16941);
xnor U19657 (N_19657,N_16624,N_15264);
nand U19658 (N_19658,N_17243,N_16499);
xnor U19659 (N_19659,N_15722,N_16690);
and U19660 (N_19660,N_16643,N_17118);
and U19661 (N_19661,N_16759,N_17231);
or U19662 (N_19662,N_16212,N_15576);
nand U19663 (N_19663,N_15778,N_17410);
xor U19664 (N_19664,N_17300,N_15294);
nand U19665 (N_19665,N_15610,N_16760);
xnor U19666 (N_19666,N_16208,N_15156);
nor U19667 (N_19667,N_16848,N_16279);
or U19668 (N_19668,N_16732,N_16222);
nor U19669 (N_19669,N_15282,N_16761);
and U19670 (N_19670,N_15781,N_16313);
or U19671 (N_19671,N_15133,N_16070);
nand U19672 (N_19672,N_15436,N_17025);
or U19673 (N_19673,N_17468,N_17203);
or U19674 (N_19674,N_16918,N_15469);
nor U19675 (N_19675,N_17218,N_16553);
and U19676 (N_19676,N_15233,N_17424);
or U19677 (N_19677,N_16073,N_16460);
nand U19678 (N_19678,N_15038,N_15264);
xor U19679 (N_19679,N_16351,N_15478);
nor U19680 (N_19680,N_16834,N_15565);
nand U19681 (N_19681,N_15896,N_15868);
or U19682 (N_19682,N_16856,N_15294);
or U19683 (N_19683,N_15830,N_16283);
or U19684 (N_19684,N_15945,N_16273);
and U19685 (N_19685,N_17044,N_15242);
nand U19686 (N_19686,N_15448,N_16836);
or U19687 (N_19687,N_17000,N_15125);
or U19688 (N_19688,N_15299,N_15202);
nor U19689 (N_19689,N_16958,N_15640);
or U19690 (N_19690,N_15532,N_16598);
nor U19691 (N_19691,N_15751,N_15662);
and U19692 (N_19692,N_15806,N_16131);
nor U19693 (N_19693,N_16596,N_15604);
and U19694 (N_19694,N_15126,N_16994);
and U19695 (N_19695,N_15556,N_16853);
and U19696 (N_19696,N_17381,N_15221);
nand U19697 (N_19697,N_16492,N_16690);
or U19698 (N_19698,N_17479,N_15516);
or U19699 (N_19699,N_16256,N_15970);
nand U19700 (N_19700,N_16500,N_16892);
and U19701 (N_19701,N_17418,N_15916);
xor U19702 (N_19702,N_15095,N_15308);
xor U19703 (N_19703,N_17044,N_15905);
xor U19704 (N_19704,N_15946,N_15809);
xnor U19705 (N_19705,N_17235,N_16171);
nor U19706 (N_19706,N_15569,N_17163);
or U19707 (N_19707,N_16793,N_15878);
or U19708 (N_19708,N_16601,N_15183);
or U19709 (N_19709,N_16151,N_16660);
or U19710 (N_19710,N_16406,N_15248);
and U19711 (N_19711,N_16790,N_16156);
and U19712 (N_19712,N_15334,N_15075);
nor U19713 (N_19713,N_15435,N_17407);
nor U19714 (N_19714,N_15178,N_16560);
nor U19715 (N_19715,N_17350,N_17005);
xnor U19716 (N_19716,N_15045,N_16568);
and U19717 (N_19717,N_15078,N_15298);
xnor U19718 (N_19718,N_15060,N_17335);
nor U19719 (N_19719,N_17195,N_15885);
nand U19720 (N_19720,N_15791,N_17157);
nor U19721 (N_19721,N_16920,N_16446);
xor U19722 (N_19722,N_15336,N_17389);
or U19723 (N_19723,N_15282,N_15021);
nand U19724 (N_19724,N_16178,N_15980);
xor U19725 (N_19725,N_16945,N_17001);
nor U19726 (N_19726,N_17061,N_15493);
or U19727 (N_19727,N_15166,N_16695);
nand U19728 (N_19728,N_16093,N_15225);
and U19729 (N_19729,N_16728,N_17211);
and U19730 (N_19730,N_17145,N_15142);
nor U19731 (N_19731,N_16196,N_16691);
xnor U19732 (N_19732,N_17397,N_15055);
nand U19733 (N_19733,N_16305,N_16985);
or U19734 (N_19734,N_17429,N_17132);
nand U19735 (N_19735,N_17164,N_15378);
and U19736 (N_19736,N_16660,N_15705);
xor U19737 (N_19737,N_17164,N_15898);
xnor U19738 (N_19738,N_15438,N_15393);
nand U19739 (N_19739,N_15729,N_16365);
or U19740 (N_19740,N_16451,N_16316);
or U19741 (N_19741,N_15599,N_15151);
nor U19742 (N_19742,N_15976,N_15844);
and U19743 (N_19743,N_15524,N_16681);
xnor U19744 (N_19744,N_15720,N_16604);
and U19745 (N_19745,N_15153,N_15969);
and U19746 (N_19746,N_15358,N_15801);
or U19747 (N_19747,N_17401,N_15463);
or U19748 (N_19748,N_16107,N_15215);
nor U19749 (N_19749,N_17094,N_15277);
xnor U19750 (N_19750,N_15846,N_15463);
and U19751 (N_19751,N_15780,N_17158);
nor U19752 (N_19752,N_15763,N_15010);
nand U19753 (N_19753,N_16488,N_16227);
xor U19754 (N_19754,N_16302,N_15760);
or U19755 (N_19755,N_16694,N_16539);
or U19756 (N_19756,N_16827,N_15373);
nor U19757 (N_19757,N_15243,N_15438);
nand U19758 (N_19758,N_16914,N_16674);
xor U19759 (N_19759,N_16589,N_15840);
and U19760 (N_19760,N_15223,N_16493);
nand U19761 (N_19761,N_15321,N_17206);
nor U19762 (N_19762,N_16723,N_15123);
nor U19763 (N_19763,N_17124,N_15945);
nor U19764 (N_19764,N_16666,N_16000);
nand U19765 (N_19765,N_15718,N_16351);
xor U19766 (N_19766,N_15274,N_15488);
nand U19767 (N_19767,N_17202,N_15668);
nor U19768 (N_19768,N_17485,N_16568);
and U19769 (N_19769,N_17010,N_17322);
and U19770 (N_19770,N_17026,N_16746);
xnor U19771 (N_19771,N_15990,N_17317);
nor U19772 (N_19772,N_15791,N_15178);
xor U19773 (N_19773,N_17317,N_16263);
nor U19774 (N_19774,N_16165,N_16119);
xnor U19775 (N_19775,N_16439,N_16965);
and U19776 (N_19776,N_16659,N_16621);
and U19777 (N_19777,N_15694,N_17198);
or U19778 (N_19778,N_15537,N_16997);
and U19779 (N_19779,N_15929,N_15078);
xor U19780 (N_19780,N_16850,N_16286);
and U19781 (N_19781,N_16289,N_17425);
or U19782 (N_19782,N_15590,N_15850);
nor U19783 (N_19783,N_15499,N_15312);
nor U19784 (N_19784,N_16453,N_16547);
nand U19785 (N_19785,N_15340,N_15982);
xnor U19786 (N_19786,N_15929,N_16403);
or U19787 (N_19787,N_15861,N_15451);
or U19788 (N_19788,N_17257,N_17332);
xor U19789 (N_19789,N_15622,N_15470);
nand U19790 (N_19790,N_15032,N_16430);
nand U19791 (N_19791,N_16816,N_15312);
nor U19792 (N_19792,N_15639,N_17417);
nand U19793 (N_19793,N_15569,N_15127);
or U19794 (N_19794,N_17379,N_15755);
and U19795 (N_19795,N_16019,N_17329);
nor U19796 (N_19796,N_16526,N_17474);
or U19797 (N_19797,N_15838,N_15280);
nor U19798 (N_19798,N_16514,N_15827);
or U19799 (N_19799,N_16405,N_16937);
xor U19800 (N_19800,N_17078,N_15215);
and U19801 (N_19801,N_16018,N_16540);
or U19802 (N_19802,N_16482,N_17136);
nand U19803 (N_19803,N_16089,N_16080);
xor U19804 (N_19804,N_16092,N_16258);
or U19805 (N_19805,N_16059,N_16395);
and U19806 (N_19806,N_15327,N_15164);
nor U19807 (N_19807,N_16554,N_15249);
or U19808 (N_19808,N_15901,N_17239);
nand U19809 (N_19809,N_15023,N_15147);
or U19810 (N_19810,N_15175,N_16618);
and U19811 (N_19811,N_17316,N_15531);
xor U19812 (N_19812,N_17308,N_16507);
nor U19813 (N_19813,N_16203,N_15930);
xnor U19814 (N_19814,N_15074,N_17207);
xnor U19815 (N_19815,N_16938,N_17399);
and U19816 (N_19816,N_15684,N_16110);
nor U19817 (N_19817,N_16658,N_16072);
nor U19818 (N_19818,N_16463,N_16413);
xnor U19819 (N_19819,N_16683,N_15428);
nor U19820 (N_19820,N_15290,N_16558);
nor U19821 (N_19821,N_17408,N_17297);
or U19822 (N_19822,N_15460,N_17349);
xnor U19823 (N_19823,N_15410,N_15557);
nand U19824 (N_19824,N_16714,N_16925);
nor U19825 (N_19825,N_16099,N_15224);
and U19826 (N_19826,N_16554,N_16590);
and U19827 (N_19827,N_16763,N_16360);
or U19828 (N_19828,N_16234,N_15672);
nand U19829 (N_19829,N_16438,N_16512);
nor U19830 (N_19830,N_16461,N_15392);
and U19831 (N_19831,N_15672,N_17219);
nand U19832 (N_19832,N_16190,N_16397);
xor U19833 (N_19833,N_15649,N_17440);
or U19834 (N_19834,N_15973,N_17451);
nor U19835 (N_19835,N_15456,N_16672);
nor U19836 (N_19836,N_17034,N_15201);
and U19837 (N_19837,N_17003,N_17125);
and U19838 (N_19838,N_16426,N_15593);
nor U19839 (N_19839,N_16830,N_16666);
xor U19840 (N_19840,N_15017,N_17153);
or U19841 (N_19841,N_15967,N_16717);
or U19842 (N_19842,N_16151,N_16424);
or U19843 (N_19843,N_16203,N_16392);
nor U19844 (N_19844,N_15209,N_17040);
and U19845 (N_19845,N_15170,N_15558);
nor U19846 (N_19846,N_16667,N_16022);
xor U19847 (N_19847,N_16249,N_15849);
xnor U19848 (N_19848,N_16904,N_15685);
and U19849 (N_19849,N_15472,N_15768);
nor U19850 (N_19850,N_16075,N_15119);
and U19851 (N_19851,N_17013,N_15238);
xor U19852 (N_19852,N_16167,N_15965);
nand U19853 (N_19853,N_15336,N_16231);
nor U19854 (N_19854,N_15229,N_15165);
nor U19855 (N_19855,N_16190,N_16484);
or U19856 (N_19856,N_15661,N_16108);
nor U19857 (N_19857,N_16436,N_16673);
nor U19858 (N_19858,N_15992,N_15374);
nand U19859 (N_19859,N_15926,N_16926);
nor U19860 (N_19860,N_16897,N_15155);
nor U19861 (N_19861,N_16282,N_15942);
or U19862 (N_19862,N_16269,N_15014);
and U19863 (N_19863,N_15149,N_15961);
or U19864 (N_19864,N_16027,N_15491);
nor U19865 (N_19865,N_15397,N_16941);
xor U19866 (N_19866,N_17038,N_15643);
and U19867 (N_19867,N_16369,N_16607);
nand U19868 (N_19868,N_15385,N_15853);
nand U19869 (N_19869,N_16833,N_17318);
and U19870 (N_19870,N_16579,N_15232);
nor U19871 (N_19871,N_16200,N_15316);
or U19872 (N_19872,N_15491,N_16199);
or U19873 (N_19873,N_17346,N_16059);
or U19874 (N_19874,N_16627,N_15961);
nor U19875 (N_19875,N_15676,N_15851);
and U19876 (N_19876,N_15457,N_15428);
xor U19877 (N_19877,N_16170,N_17494);
xnor U19878 (N_19878,N_15467,N_15753);
nand U19879 (N_19879,N_15230,N_16603);
and U19880 (N_19880,N_15006,N_17353);
or U19881 (N_19881,N_15035,N_16921);
nand U19882 (N_19882,N_17392,N_15686);
nor U19883 (N_19883,N_15423,N_15933);
nor U19884 (N_19884,N_15630,N_15140);
or U19885 (N_19885,N_17039,N_16842);
nor U19886 (N_19886,N_17463,N_15522);
or U19887 (N_19887,N_15661,N_17189);
nand U19888 (N_19888,N_15805,N_15484);
or U19889 (N_19889,N_16749,N_15327);
or U19890 (N_19890,N_17195,N_15735);
xnor U19891 (N_19891,N_16335,N_17030);
nor U19892 (N_19892,N_17389,N_15000);
nor U19893 (N_19893,N_16453,N_16694);
nand U19894 (N_19894,N_15939,N_16248);
xor U19895 (N_19895,N_15088,N_16050);
nand U19896 (N_19896,N_16622,N_15134);
nor U19897 (N_19897,N_16548,N_17367);
or U19898 (N_19898,N_16469,N_15932);
and U19899 (N_19899,N_16355,N_15427);
and U19900 (N_19900,N_16808,N_15659);
xnor U19901 (N_19901,N_15810,N_17441);
and U19902 (N_19902,N_16940,N_16494);
nor U19903 (N_19903,N_16688,N_15098);
xor U19904 (N_19904,N_15161,N_16575);
nor U19905 (N_19905,N_17371,N_15988);
or U19906 (N_19906,N_15020,N_15576);
nor U19907 (N_19907,N_16645,N_17288);
nor U19908 (N_19908,N_16519,N_17466);
and U19909 (N_19909,N_16694,N_16057);
and U19910 (N_19910,N_16019,N_15923);
xor U19911 (N_19911,N_15683,N_15912);
or U19912 (N_19912,N_16239,N_16470);
nand U19913 (N_19913,N_15048,N_16071);
and U19914 (N_19914,N_15453,N_16925);
nand U19915 (N_19915,N_16650,N_15332);
or U19916 (N_19916,N_15730,N_17410);
or U19917 (N_19917,N_17041,N_15054);
nand U19918 (N_19918,N_15539,N_15434);
nand U19919 (N_19919,N_15668,N_16119);
and U19920 (N_19920,N_15532,N_16508);
xnor U19921 (N_19921,N_15078,N_15824);
or U19922 (N_19922,N_16767,N_16366);
or U19923 (N_19923,N_15151,N_16563);
or U19924 (N_19924,N_15931,N_16273);
and U19925 (N_19925,N_16231,N_17021);
nand U19926 (N_19926,N_16123,N_15311);
xor U19927 (N_19927,N_16601,N_16453);
or U19928 (N_19928,N_15213,N_16727);
xnor U19929 (N_19929,N_16598,N_15551);
nor U19930 (N_19930,N_15471,N_17467);
nor U19931 (N_19931,N_17184,N_17187);
nand U19932 (N_19932,N_15736,N_16052);
xnor U19933 (N_19933,N_17400,N_15180);
and U19934 (N_19934,N_16098,N_16481);
and U19935 (N_19935,N_17307,N_16799);
nor U19936 (N_19936,N_16449,N_16363);
or U19937 (N_19937,N_17100,N_16434);
and U19938 (N_19938,N_16564,N_15093);
nand U19939 (N_19939,N_16222,N_17173);
xor U19940 (N_19940,N_15913,N_17354);
nor U19941 (N_19941,N_17005,N_16191);
nand U19942 (N_19942,N_15171,N_16742);
nand U19943 (N_19943,N_15907,N_17329);
nand U19944 (N_19944,N_17098,N_16056);
nor U19945 (N_19945,N_16388,N_15502);
nor U19946 (N_19946,N_17275,N_16182);
nand U19947 (N_19947,N_17336,N_15380);
nor U19948 (N_19948,N_16498,N_15320);
or U19949 (N_19949,N_16000,N_16152);
nor U19950 (N_19950,N_15822,N_16666);
nor U19951 (N_19951,N_17242,N_15731);
xor U19952 (N_19952,N_17163,N_17319);
nor U19953 (N_19953,N_17485,N_15884);
xnor U19954 (N_19954,N_17415,N_17072);
and U19955 (N_19955,N_15805,N_15598);
and U19956 (N_19956,N_16990,N_17146);
and U19957 (N_19957,N_17491,N_15206);
and U19958 (N_19958,N_17075,N_17438);
nand U19959 (N_19959,N_15887,N_17202);
xnor U19960 (N_19960,N_15481,N_17079);
nand U19961 (N_19961,N_15188,N_15680);
nand U19962 (N_19962,N_17244,N_15039);
and U19963 (N_19963,N_16607,N_17282);
nor U19964 (N_19964,N_16549,N_15291);
xor U19965 (N_19965,N_16213,N_16103);
and U19966 (N_19966,N_15569,N_17410);
nand U19967 (N_19967,N_16362,N_17417);
nand U19968 (N_19968,N_15573,N_15330);
nor U19969 (N_19969,N_15515,N_17337);
and U19970 (N_19970,N_16376,N_15817);
nor U19971 (N_19971,N_15843,N_15741);
nor U19972 (N_19972,N_16477,N_17490);
and U19973 (N_19973,N_16930,N_16845);
nand U19974 (N_19974,N_15459,N_16962);
xor U19975 (N_19975,N_15511,N_17012);
or U19976 (N_19976,N_17006,N_17448);
and U19977 (N_19977,N_17477,N_16024);
xnor U19978 (N_19978,N_15018,N_16013);
nor U19979 (N_19979,N_15857,N_15593);
xor U19980 (N_19980,N_15795,N_17458);
or U19981 (N_19981,N_15570,N_16510);
nand U19982 (N_19982,N_15638,N_15930);
xnor U19983 (N_19983,N_15526,N_15591);
xor U19984 (N_19984,N_16987,N_15162);
and U19985 (N_19985,N_15573,N_16243);
nor U19986 (N_19986,N_16639,N_15292);
or U19987 (N_19987,N_16891,N_15298);
xnor U19988 (N_19988,N_15920,N_16488);
and U19989 (N_19989,N_17306,N_15322);
nand U19990 (N_19990,N_15212,N_16591);
and U19991 (N_19991,N_16223,N_17149);
or U19992 (N_19992,N_15506,N_17467);
xnor U19993 (N_19993,N_16478,N_16080);
xor U19994 (N_19994,N_15047,N_15500);
nor U19995 (N_19995,N_16392,N_17469);
and U19996 (N_19996,N_15830,N_17450);
nor U19997 (N_19997,N_17389,N_17275);
nor U19998 (N_19998,N_17437,N_15881);
and U19999 (N_19999,N_16193,N_15032);
and U20000 (N_20000,N_18285,N_19908);
nor U20001 (N_20001,N_18754,N_18486);
xnor U20002 (N_20002,N_19018,N_18212);
xor U20003 (N_20003,N_18210,N_17650);
or U20004 (N_20004,N_18637,N_19541);
xor U20005 (N_20005,N_17748,N_18480);
nand U20006 (N_20006,N_19848,N_18275);
nor U20007 (N_20007,N_17539,N_19963);
nor U20008 (N_20008,N_18825,N_17556);
nand U20009 (N_20009,N_18393,N_18297);
and U20010 (N_20010,N_17899,N_18026);
nand U20011 (N_20011,N_18282,N_19966);
and U20012 (N_20012,N_19225,N_19166);
nand U20013 (N_20013,N_18472,N_19352);
nor U20014 (N_20014,N_19329,N_19962);
nor U20015 (N_20015,N_19955,N_19637);
or U20016 (N_20016,N_19453,N_17549);
or U20017 (N_20017,N_19892,N_18778);
or U20018 (N_20018,N_18673,N_17775);
nor U20019 (N_20019,N_18197,N_18135);
nand U20020 (N_20020,N_19192,N_17860);
xor U20021 (N_20021,N_19200,N_19891);
nor U20022 (N_20022,N_18864,N_17636);
and U20023 (N_20023,N_18281,N_18007);
xor U20024 (N_20024,N_19996,N_18676);
nor U20025 (N_20025,N_17851,N_19814);
nor U20026 (N_20026,N_18389,N_19792);
or U20027 (N_20027,N_19958,N_18974);
and U20028 (N_20028,N_17713,N_19954);
nor U20029 (N_20029,N_18614,N_18479);
nand U20030 (N_20030,N_19427,N_18196);
nand U20031 (N_20031,N_18292,N_19496);
and U20032 (N_20032,N_19097,N_19842);
or U20033 (N_20033,N_18990,N_18538);
nand U20034 (N_20034,N_18846,N_18330);
nor U20035 (N_20035,N_19417,N_19900);
xnor U20036 (N_20036,N_19838,N_17550);
nor U20037 (N_20037,N_19174,N_19970);
or U20038 (N_20038,N_19101,N_18645);
xnor U20039 (N_20039,N_17856,N_19687);
and U20040 (N_20040,N_18862,N_18712);
nor U20041 (N_20041,N_18312,N_17938);
nand U20042 (N_20042,N_18811,N_18772);
nor U20043 (N_20043,N_19939,N_19650);
or U20044 (N_20044,N_18856,N_18554);
xor U20045 (N_20045,N_17753,N_17947);
nand U20046 (N_20046,N_19447,N_19491);
or U20047 (N_20047,N_18871,N_19198);
or U20048 (N_20048,N_19671,N_18437);
nand U20049 (N_20049,N_19221,N_19064);
and U20050 (N_20050,N_19045,N_18761);
nor U20051 (N_20051,N_17566,N_19202);
nor U20052 (N_20052,N_19736,N_18505);
or U20053 (N_20053,N_18355,N_18127);
xor U20054 (N_20054,N_18626,N_18648);
and U20055 (N_20055,N_17507,N_18009);
or U20056 (N_20056,N_19394,N_18839);
nor U20057 (N_20057,N_19946,N_18488);
nor U20058 (N_20058,N_19616,N_19381);
or U20059 (N_20059,N_19607,N_19817);
and U20060 (N_20060,N_19796,N_19245);
xnor U20061 (N_20061,N_17502,N_19367);
or U20062 (N_20062,N_17803,N_18113);
and U20063 (N_20063,N_18843,N_19811);
xor U20064 (N_20064,N_18891,N_18384);
xnor U20065 (N_20065,N_17784,N_19091);
and U20066 (N_20066,N_18179,N_18216);
xnor U20067 (N_20067,N_19730,N_19191);
or U20068 (N_20068,N_18930,N_18248);
or U20069 (N_20069,N_18701,N_18077);
nor U20070 (N_20070,N_19078,N_18391);
and U20071 (N_20071,N_19278,N_18064);
or U20072 (N_20072,N_19507,N_19333);
xor U20073 (N_20073,N_19022,N_19806);
xor U20074 (N_20074,N_17805,N_19139);
nor U20075 (N_20075,N_19533,N_19921);
nor U20076 (N_20076,N_19277,N_19925);
and U20077 (N_20077,N_18332,N_17850);
xor U20078 (N_20078,N_17513,N_19033);
xnor U20079 (N_20079,N_17921,N_19084);
nand U20080 (N_20080,N_18895,N_19889);
or U20081 (N_20081,N_19463,N_17546);
xor U20082 (N_20082,N_18674,N_19873);
and U20083 (N_20083,N_19280,N_19458);
nor U20084 (N_20084,N_17822,N_18143);
and U20085 (N_20085,N_18522,N_19821);
and U20086 (N_20086,N_19731,N_19297);
nand U20087 (N_20087,N_17754,N_18193);
nand U20088 (N_20088,N_18059,N_18624);
nor U20089 (N_20089,N_17571,N_18455);
nand U20090 (N_20090,N_18867,N_18922);
or U20091 (N_20091,N_18289,N_19393);
or U20092 (N_20092,N_18691,N_18090);
xor U20093 (N_20093,N_17970,N_18129);
and U20094 (N_20094,N_17862,N_19475);
and U20095 (N_20095,N_17857,N_19069);
xor U20096 (N_20096,N_17519,N_18906);
xnor U20097 (N_20097,N_17742,N_18926);
nor U20098 (N_20098,N_19083,N_19454);
xor U20099 (N_20099,N_18866,N_18374);
nand U20100 (N_20100,N_18719,N_17501);
or U20101 (N_20101,N_19542,N_19476);
or U20102 (N_20102,N_17879,N_17757);
nand U20103 (N_20103,N_19721,N_17760);
nor U20104 (N_20104,N_19082,N_18787);
or U20105 (N_20105,N_19895,N_19754);
and U20106 (N_20106,N_18434,N_18299);
nor U20107 (N_20107,N_18447,N_18158);
nor U20108 (N_20108,N_17536,N_18329);
nand U20109 (N_20109,N_19711,N_18341);
or U20110 (N_20110,N_18547,N_17737);
xor U20111 (N_20111,N_17796,N_19852);
nor U20112 (N_20112,N_19956,N_17594);
and U20113 (N_20113,N_17816,N_18633);
and U20114 (N_20114,N_17680,N_19779);
nor U20115 (N_20115,N_17649,N_18133);
or U20116 (N_20116,N_17666,N_18584);
nor U20117 (N_20117,N_17942,N_17893);
xor U20118 (N_20118,N_19851,N_18487);
xnor U20119 (N_20119,N_18516,N_18756);
or U20120 (N_20120,N_18310,N_19087);
xnor U20121 (N_20121,N_19461,N_18670);
nor U20122 (N_20122,N_19307,N_18470);
nand U20123 (N_20123,N_18445,N_19723);
and U20124 (N_20124,N_19778,N_17962);
and U20125 (N_20125,N_19922,N_19421);
or U20126 (N_20126,N_18741,N_17696);
and U20127 (N_20127,N_19456,N_18550);
or U20128 (N_20128,N_18944,N_18927);
and U20129 (N_20129,N_19459,N_19378);
or U20130 (N_20130,N_17577,N_18313);
or U20131 (N_20131,N_19414,N_18591);
nor U20132 (N_20132,N_17526,N_19782);
and U20133 (N_20133,N_17853,N_17665);
nand U20134 (N_20134,N_19290,N_19302);
xor U20135 (N_20135,N_19219,N_19562);
and U20136 (N_20136,N_19442,N_18656);
or U20137 (N_20137,N_18072,N_18755);
xnor U20138 (N_20138,N_17761,N_19745);
nor U20139 (N_20139,N_19951,N_18677);
and U20140 (N_20140,N_17592,N_19357);
nand U20141 (N_20141,N_18597,N_17887);
nand U20142 (N_20142,N_18467,N_19250);
nand U20143 (N_20143,N_18457,N_18991);
or U20144 (N_20144,N_17533,N_17833);
nand U20145 (N_20145,N_18635,N_19434);
and U20146 (N_20146,N_18841,N_18224);
nor U20147 (N_20147,N_17509,N_18810);
and U20148 (N_20148,N_18022,N_19594);
xor U20149 (N_20149,N_19089,N_17747);
xnor U20150 (N_20150,N_17770,N_18308);
nand U20151 (N_20151,N_18442,N_19617);
nand U20152 (N_20152,N_17609,N_19478);
and U20153 (N_20153,N_18105,N_17741);
or U20154 (N_20154,N_17598,N_17905);
nor U20155 (N_20155,N_19490,N_19010);
and U20156 (N_20156,N_19989,N_19327);
and U20157 (N_20157,N_19627,N_18180);
nor U20158 (N_20158,N_19474,N_17832);
nor U20159 (N_20159,N_19488,N_18565);
or U20160 (N_20160,N_19655,N_18764);
nor U20161 (N_20161,N_17607,N_17817);
and U20162 (N_20162,N_19808,N_18784);
xor U20163 (N_20163,N_18613,N_18937);
or U20164 (N_20164,N_18278,N_18604);
and U20165 (N_20165,N_19030,N_19866);
nand U20166 (N_20166,N_18309,N_17614);
and U20167 (N_20167,N_18217,N_19812);
or U20168 (N_20168,N_17734,N_18460);
nand U20169 (N_20169,N_17984,N_17505);
or U20170 (N_20170,N_17884,N_19880);
nor U20171 (N_20171,N_18474,N_19431);
nor U20172 (N_20172,N_19677,N_17520);
and U20173 (N_20173,N_18478,N_18087);
and U20174 (N_20174,N_19398,N_19580);
nand U20175 (N_20175,N_19154,N_18094);
and U20176 (N_20176,N_19395,N_19810);
and U20177 (N_20177,N_19338,N_18435);
and U20178 (N_20178,N_18439,N_18979);
and U20179 (N_20179,N_18184,N_19377);
xor U20180 (N_20180,N_18177,N_19647);
nand U20181 (N_20181,N_18917,N_18792);
nand U20182 (N_20182,N_19971,N_17578);
and U20183 (N_20183,N_19618,N_18743);
nor U20184 (N_20184,N_19003,N_19901);
and U20185 (N_20185,N_17956,N_17957);
xor U20186 (N_20186,N_19856,N_19651);
and U20187 (N_20187,N_19011,N_17854);
or U20188 (N_20188,N_18735,N_17504);
nor U20189 (N_20189,N_17656,N_18779);
and U20190 (N_20190,N_19790,N_18786);
nand U20191 (N_20191,N_17937,N_18476);
xor U20192 (N_20192,N_19700,N_19199);
and U20193 (N_20193,N_19585,N_18629);
nand U20194 (N_20194,N_18245,N_18270);
or U20195 (N_20195,N_19017,N_18672);
and U20196 (N_20196,N_19554,N_18050);
or U20197 (N_20197,N_19320,N_19841);
or U20198 (N_20198,N_18973,N_18412);
or U20199 (N_20199,N_18508,N_19645);
and U20200 (N_20200,N_17848,N_18305);
xnor U20201 (N_20201,N_18578,N_18834);
nor U20202 (N_20202,N_19146,N_18942);
nand U20203 (N_20203,N_18288,N_19027);
nand U20204 (N_20204,N_19781,N_19959);
and U20205 (N_20205,N_18018,N_17898);
nor U20206 (N_20206,N_18823,N_18485);
nor U20207 (N_20207,N_18527,N_18581);
nor U20208 (N_20208,N_19780,N_19614);
nand U20209 (N_20209,N_19228,N_19215);
and U20210 (N_20210,N_18882,N_19141);
nor U20211 (N_20211,N_19886,N_18532);
or U20212 (N_20212,N_18892,N_17993);
nand U20213 (N_20213,N_19525,N_18176);
nor U20214 (N_20214,N_18189,N_17808);
nand U20215 (N_20215,N_19828,N_18720);
xor U20216 (N_20216,N_19203,N_19813);
xor U20217 (N_20217,N_19638,N_19117);
and U20218 (N_20218,N_17944,N_18780);
and U20219 (N_20219,N_19578,N_19771);
nand U20220 (N_20220,N_19443,N_17844);
xnor U20221 (N_20221,N_19573,N_18767);
nor U20222 (N_20222,N_18185,N_18958);
or U20223 (N_20223,N_17785,N_18397);
or U20224 (N_20224,N_18988,N_18315);
and U20225 (N_20225,N_18379,N_19094);
nand U20226 (N_20226,N_19267,N_19244);
or U20227 (N_20227,N_19483,N_18829);
or U20228 (N_20228,N_19349,N_19864);
nand U20229 (N_20229,N_18413,N_18820);
or U20230 (N_20230,N_19881,N_18259);
xor U20231 (N_20231,N_17708,N_19997);
nor U20232 (N_20232,N_18378,N_19471);
or U20233 (N_20233,N_19994,N_19513);
or U20234 (N_20234,N_17771,N_19888);
nor U20235 (N_20235,N_19360,N_19693);
or U20236 (N_20236,N_18647,N_19998);
and U20237 (N_20237,N_19912,N_19060);
xor U20238 (N_20238,N_19540,N_17729);
and U20239 (N_20239,N_18414,N_19967);
xnor U20240 (N_20240,N_18943,N_18541);
xnor U20241 (N_20241,N_19473,N_18365);
nor U20242 (N_20242,N_18542,N_18237);
or U20243 (N_20243,N_19760,N_19430);
nand U20244 (N_20244,N_18172,N_19086);
xor U20245 (N_20245,N_17903,N_19911);
and U20246 (N_20246,N_17839,N_19846);
nand U20247 (N_20247,N_17830,N_19752);
or U20248 (N_20248,N_19735,N_18835);
nor U20249 (N_20249,N_17672,N_19691);
nand U20250 (N_20250,N_19249,N_18395);
nand U20251 (N_20251,N_17620,N_18998);
nand U20252 (N_20252,N_19397,N_19505);
or U20253 (N_20253,N_19685,N_17568);
and U20254 (N_20254,N_19331,N_19095);
and U20255 (N_20255,N_17906,N_19220);
nor U20256 (N_20256,N_19213,N_17826);
or U20257 (N_20257,N_19014,N_17915);
nor U20258 (N_20258,N_19621,N_19118);
nand U20259 (N_20259,N_18428,N_18427);
nor U20260 (N_20260,N_17930,N_19798);
nand U20261 (N_20261,N_18955,N_18348);
or U20262 (N_20262,N_18001,N_19706);
xnor U20263 (N_20263,N_19226,N_18777);
and U20264 (N_20264,N_19521,N_17829);
xor U20265 (N_20265,N_18593,N_18115);
nor U20266 (N_20266,N_19999,N_18223);
nand U20267 (N_20267,N_19452,N_18514);
and U20268 (N_20268,N_17807,N_18168);
and U20269 (N_20269,N_18661,N_18244);
and U20270 (N_20270,N_19719,N_18911);
nor U20271 (N_20271,N_18410,N_17617);
xnor U20272 (N_20272,N_18536,N_18665);
and U20273 (N_20273,N_19270,N_18325);
nand U20274 (N_20274,N_18752,N_19558);
and U20275 (N_20275,N_19107,N_18298);
or U20276 (N_20276,N_19231,N_19259);
and U20277 (N_20277,N_17518,N_19072);
or U20278 (N_20278,N_19328,N_17897);
xor U20279 (N_20279,N_19389,N_18011);
xor U20280 (N_20280,N_18795,N_19919);
xor U20281 (N_20281,N_18008,N_18383);
and U20282 (N_20282,N_19597,N_18600);
or U20283 (N_20283,N_18746,N_19609);
nand U20284 (N_20284,N_18709,N_19067);
xor U20285 (N_20285,N_19859,N_18082);
and U20286 (N_20286,N_17939,N_19340);
or U20287 (N_20287,N_18257,N_18704);
nor U20288 (N_20288,N_18632,N_17963);
xor U20289 (N_20289,N_19724,N_17874);
xnor U20290 (N_20290,N_19776,N_17663);
nor U20291 (N_20291,N_18065,N_17587);
and U20292 (N_20292,N_17869,N_19283);
and U20293 (N_20293,N_17500,N_18900);
nand U20294 (N_20294,N_17685,N_18119);
nand U20295 (N_20295,N_17809,N_18664);
or U20296 (N_20296,N_18443,N_18114);
or U20297 (N_20297,N_17995,N_18889);
nor U20298 (N_20298,N_18401,N_19242);
nor U20299 (N_20299,N_19953,N_19608);
nand U20300 (N_20300,N_19756,N_17994);
nor U20301 (N_20301,N_17688,N_18546);
nand U20302 (N_20302,N_19695,N_19112);
nand U20303 (N_20303,N_18240,N_19524);
or U20304 (N_20304,N_19182,N_18070);
or U20305 (N_20305,N_18452,N_19142);
and U20306 (N_20306,N_18468,N_17767);
or U20307 (N_20307,N_18576,N_18420);
or U20308 (N_20308,N_19335,N_18710);
or U20309 (N_20309,N_19034,N_18641);
and U20310 (N_20310,N_19624,N_17732);
or U20311 (N_20311,N_17928,N_17916);
or U20312 (N_20312,N_18969,N_17628);
nor U20313 (N_20313,N_18684,N_18347);
xnor U20314 (N_20314,N_18067,N_18729);
or U20315 (N_20315,N_19289,N_17693);
and U20316 (N_20316,N_18699,N_18489);
and U20317 (N_20317,N_18254,N_17543);
and U20318 (N_20318,N_19844,N_18870);
xnor U20319 (N_20319,N_18590,N_17954);
nand U20320 (N_20320,N_18517,N_19031);
nor U20321 (N_20321,N_17981,N_18459);
nand U20322 (N_20322,N_18218,N_18350);
or U20323 (N_20323,N_17837,N_18441);
xnor U20324 (N_20324,N_19899,N_19240);
and U20325 (N_20325,N_18147,N_19871);
and U20326 (N_20326,N_19547,N_19682);
nand U20327 (N_20327,N_17682,N_17907);
or U20328 (N_20328,N_17866,N_19666);
or U20329 (N_20329,N_17553,N_19184);
and U20330 (N_20330,N_17600,N_17987);
xnor U20331 (N_20331,N_18186,N_17618);
and U20332 (N_20332,N_17831,N_19628);
nand U20333 (N_20333,N_18235,N_19744);
xnor U20334 (N_20334,N_17644,N_19630);
or U20335 (N_20335,N_19725,N_19080);
nor U20336 (N_20336,N_17664,N_18782);
or U20337 (N_20337,N_18970,N_19122);
nand U20338 (N_20338,N_19163,N_18923);
nand U20339 (N_20339,N_18725,N_19980);
and U20340 (N_20340,N_18205,N_19243);
nor U20341 (N_20341,N_17958,N_19081);
xnor U20342 (N_20342,N_18731,N_19282);
nand U20343 (N_20343,N_18530,N_19276);
nor U20344 (N_20344,N_17799,N_19559);
xor U20345 (N_20345,N_19254,N_18074);
xor U20346 (N_20346,N_18596,N_17700);
nand U20347 (N_20347,N_17782,N_19622);
or U20348 (N_20348,N_19110,N_18436);
nor U20349 (N_20349,N_19363,N_18417);
or U20350 (N_20350,N_17911,N_18750);
or U20351 (N_20351,N_18992,N_18890);
nand U20352 (N_20352,N_19286,N_17818);
nand U20353 (N_20353,N_18826,N_19920);
nand U20354 (N_20354,N_18797,N_19129);
and U20355 (N_20355,N_17750,N_19294);
nor U20356 (N_20356,N_18838,N_17972);
xnor U20357 (N_20357,N_18881,N_18372);
or U20358 (N_20358,N_17941,N_17904);
xnor U20359 (N_20359,N_19455,N_17622);
xor U20360 (N_20360,N_17586,N_18017);
nor U20361 (N_20361,N_17864,N_19990);
nor U20362 (N_20362,N_19661,N_18836);
xnor U20363 (N_20363,N_19680,N_17601);
and U20364 (N_20364,N_19001,N_17593);
and U20365 (N_20365,N_18461,N_17631);
nor U20366 (N_20366,N_19576,N_18692);
nor U20367 (N_20367,N_19937,N_19789);
or U20368 (N_20368,N_18099,N_19992);
xnor U20369 (N_20369,N_18213,N_19986);
nor U20370 (N_20370,N_17986,N_18016);
nand U20371 (N_20371,N_18802,N_18644);
xnor U20372 (N_20372,N_17707,N_18469);
nand U20373 (N_20373,N_17919,N_19879);
or U20374 (N_20374,N_18086,N_17858);
nand U20375 (N_20375,N_17670,N_19212);
and U20376 (N_20376,N_17780,N_18221);
xor U20377 (N_20377,N_19061,N_19615);
nor U20378 (N_20378,N_18095,N_17629);
or U20379 (N_20379,N_19935,N_19613);
and U20380 (N_20380,N_19484,N_17875);
nand U20381 (N_20381,N_19298,N_19234);
and U20382 (N_20382,N_17605,N_18708);
xnor U20383 (N_20383,N_18175,N_19799);
and U20384 (N_20384,N_19587,N_18872);
and U20385 (N_20385,N_18139,N_17812);
xnor U20386 (N_20386,N_18323,N_18760);
and U20387 (N_20387,N_18047,N_18242);
or U20388 (N_20388,N_18230,N_18142);
nand U20389 (N_20389,N_18561,N_19108);
nand U20390 (N_20390,N_17745,N_18322);
and U20391 (N_20391,N_18239,N_19514);
xnor U20392 (N_20392,N_18306,N_17611);
or U20393 (N_20393,N_19281,N_19652);
and U20394 (N_20394,N_19102,N_17562);
nand U20395 (N_20395,N_17959,N_18751);
nor U20396 (N_20396,N_17574,N_18769);
nor U20397 (N_20397,N_18736,N_18080);
nand U20398 (N_20398,N_17590,N_18199);
xnor U20399 (N_20399,N_18314,N_19271);
and U20400 (N_20400,N_19450,N_18660);
nand U20401 (N_20401,N_19529,N_19639);
nor U20402 (N_20402,N_18933,N_19116);
and U20403 (N_20403,N_19858,N_19460);
or U20404 (N_20404,N_18575,N_17804);
xor U20405 (N_20405,N_19365,N_18331);
and U20406 (N_20406,N_17648,N_17651);
xnor U20407 (N_20407,N_17730,N_19186);
nand U20408 (N_20408,N_18643,N_19492);
xnor U20409 (N_20409,N_18494,N_18939);
nand U20410 (N_20410,N_18302,N_18954);
xnor U20411 (N_20411,N_19293,N_19803);
xor U20412 (N_20412,N_19390,N_18931);
nor U20413 (N_20413,N_18907,N_17668);
nor U20414 (N_20414,N_19611,N_18261);
nand U20415 (N_20415,N_18078,N_17744);
xor U20416 (N_20416,N_17765,N_18421);
nand U20417 (N_20417,N_19697,N_17949);
or U20418 (N_20418,N_19111,N_18963);
and U20419 (N_20419,N_17978,N_19256);
xor U20420 (N_20420,N_18097,N_18390);
or U20421 (N_20421,N_18869,N_18985);
nor U20422 (N_20422,N_18873,N_18606);
xnor U20423 (N_20423,N_19362,N_19028);
nor U20424 (N_20424,N_19173,N_19984);
nor U20425 (N_20425,N_18765,N_19763);
xor U20426 (N_20426,N_19550,N_19712);
nor U20427 (N_20427,N_19464,N_18291);
and U20428 (N_20428,N_18818,N_18117);
nand U20429 (N_20429,N_19620,N_18631);
xor U20430 (N_20430,N_19123,N_19926);
xor U20431 (N_20431,N_19694,N_18827);
and U20432 (N_20432,N_18500,N_19209);
or U20433 (N_20433,N_19138,N_17671);
or U20434 (N_20434,N_18879,N_18776);
nand U20435 (N_20435,N_19732,N_19285);
or U20436 (N_20436,N_19995,N_18967);
nand U20437 (N_20437,N_19654,N_19158);
nor U20438 (N_20438,N_19251,N_18137);
nand U20439 (N_20439,N_19160,N_19274);
nand U20440 (N_20440,N_18983,N_19029);
xnor U20441 (N_20441,N_17652,N_17635);
nand U20442 (N_20442,N_19287,N_18646);
and U20443 (N_20443,N_17576,N_19020);
and U20444 (N_20444,N_18373,N_19235);
nand U20445 (N_20445,N_18563,N_17966);
nand U20446 (N_20446,N_17992,N_18411);
xnor U20447 (N_20447,N_19161,N_17902);
or U20448 (N_20448,N_19193,N_19016);
or U20449 (N_20449,N_17591,N_18222);
nand U20450 (N_20450,N_17841,N_17722);
nand U20451 (N_20451,N_19927,N_17813);
xor U20452 (N_20452,N_18148,N_18852);
and U20453 (N_20453,N_19265,N_19291);
or U20454 (N_20454,N_19835,N_18617);
nor U20455 (N_20455,N_17991,N_19409);
nor U20456 (N_20456,N_19435,N_19596);
nand U20457 (N_20457,N_19316,N_18418);
or U20458 (N_20458,N_18689,N_18706);
xor U20459 (N_20459,N_18821,N_19303);
and U20460 (N_20460,N_19120,N_19132);
or U20461 (N_20461,N_18948,N_19556);
or U20462 (N_20462,N_17695,N_17662);
or U20463 (N_20463,N_17878,N_19626);
or U20464 (N_20464,N_19757,N_19000);
nor U20465 (N_20465,N_18568,N_17728);
xnor U20466 (N_20466,N_18499,N_19537);
nor U20467 (N_20467,N_18110,N_18675);
or U20468 (N_20468,N_19878,N_18543);
xnor U20469 (N_20469,N_19487,N_19536);
xnor U20470 (N_20470,N_18131,N_19439);
xor U20471 (N_20471,N_17529,N_18652);
or U20472 (N_20472,N_19619,N_17752);
nor U20473 (N_20473,N_17801,N_17823);
nand U20474 (N_20474,N_18817,N_19788);
nor U20475 (N_20475,N_18620,N_18627);
nor U20476 (N_20476,N_18506,N_18667);
and U20477 (N_20477,N_18855,N_18715);
xor U20478 (N_20478,N_19188,N_19136);
nor U20479 (N_20479,N_18814,N_19632);
nand U20480 (N_20480,N_19216,N_18368);
nand U20481 (N_20481,N_19151,N_19772);
xnor U20482 (N_20482,N_19509,N_17917);
nand U20483 (N_20483,N_18858,N_18703);
or U20484 (N_20484,N_19205,N_17673);
and U20485 (N_20485,N_18512,N_19561);
nor U20486 (N_20486,N_18800,N_19148);
or U20487 (N_20487,N_18653,N_18984);
xor U20488 (N_20488,N_19702,N_19384);
or U20489 (N_20489,N_18762,N_19162);
and U20490 (N_20490,N_18697,N_18909);
nor U20491 (N_20491,N_18775,N_18369);
nor U20492 (N_20492,N_17583,N_19194);
xor U20493 (N_20493,N_19599,N_18066);
and U20494 (N_20494,N_19180,N_19893);
and U20495 (N_20495,N_19500,N_18560);
nor U20496 (N_20496,N_18128,N_19130);
nor U20497 (N_20497,N_19257,N_19009);
nand U20498 (N_20498,N_19832,N_18616);
and U20499 (N_20499,N_18111,N_19534);
or U20500 (N_20500,N_19392,N_19581);
nand U20501 (N_20501,N_19300,N_19304);
and U20502 (N_20502,N_19924,N_18136);
nor U20503 (N_20503,N_18021,N_18649);
nand U20504 (N_20504,N_18899,N_19336);
nor U20505 (N_20505,N_19058,N_19268);
and U20506 (N_20506,N_19317,N_19600);
nand U20507 (N_20507,N_19055,N_17623);
or U20508 (N_20508,N_18513,N_18049);
xnor U20509 (N_20509,N_17731,N_19560);
nor U20510 (N_20510,N_18249,N_18038);
nor U20511 (N_20511,N_19266,N_18477);
xor U20512 (N_20512,N_18409,N_19036);
xor U20513 (N_20513,N_17913,N_18075);
and U20514 (N_20514,N_17873,N_18144);
nand U20515 (N_20515,N_19241,N_19006);
or U20516 (N_20516,N_19263,N_18521);
xor U20517 (N_20517,N_19805,N_19382);
or U20518 (N_20518,N_18191,N_19531);
or U20519 (N_20519,N_17595,N_18085);
or U20520 (N_20520,N_18945,N_17868);
nand U20521 (N_20521,N_19217,N_18962);
and U20522 (N_20522,N_18200,N_17527);
or U20523 (N_20523,N_19947,N_19098);
or U20524 (N_20524,N_18051,N_18956);
xor U20525 (N_20525,N_18844,N_17781);
nand U20526 (N_20526,N_18345,N_19314);
nor U20527 (N_20527,N_19854,N_19047);
nand U20528 (N_20528,N_17867,N_18807);
and U20529 (N_20529,N_19689,N_19839);
nand U20530 (N_20530,N_18682,N_19517);
xor U20531 (N_20531,N_19444,N_18294);
or U20532 (N_20532,N_19568,N_17783);
nand U20533 (N_20533,N_19884,N_17891);
xor U20534 (N_20534,N_17900,N_19707);
nor U20535 (N_20535,N_19952,N_18096);
xor U20536 (N_20536,N_17997,N_19977);
nor U20537 (N_20537,N_18450,N_17825);
and U20538 (N_20538,N_18642,N_17777);
nor U20539 (N_20539,N_19750,N_17849);
nor U20540 (N_20540,N_17798,N_18999);
and U20541 (N_20541,N_19042,N_18759);
nor U20542 (N_20542,N_18102,N_18636);
and U20543 (N_20543,N_17739,N_19869);
and U20544 (N_20544,N_18902,N_19311);
nand U20545 (N_20545,N_19979,N_17896);
nor U20546 (N_20546,N_19761,N_19820);
and U20547 (N_20547,N_19602,N_18023);
xnor U20548 (N_20548,N_19477,N_17793);
nand U20549 (N_20549,N_19933,N_19853);
nand U20550 (N_20550,N_17872,N_18745);
xnor U20551 (N_20551,N_17934,N_18573);
xor U20552 (N_20552,N_18548,N_18953);
xnor U20553 (N_20553,N_17975,N_18303);
and U20554 (N_20554,N_18354,N_19044);
nor U20555 (N_20555,N_18630,N_18226);
and U20556 (N_20556,N_18603,N_18574);
nor U20557 (N_20557,N_18181,N_19675);
nand U20558 (N_20558,N_19169,N_18155);
nor U20559 (N_20559,N_18246,N_19785);
and U20560 (N_20560,N_18915,N_18976);
nand U20561 (N_20561,N_17691,N_19991);
nand U20562 (N_20562,N_19591,N_18952);
nor U20563 (N_20563,N_19867,N_18231);
xor U20564 (N_20564,N_18639,N_19555);
nor U20565 (N_20565,N_19155,N_18491);
or U20566 (N_20566,N_17892,N_18279);
and U20567 (N_20567,N_17755,N_19641);
or U20568 (N_20568,N_17524,N_19334);
xor U20569 (N_20569,N_18214,N_19942);
nand U20570 (N_20570,N_19318,N_19025);
nor U20571 (N_20571,N_17791,N_18093);
nand U20572 (N_20572,N_19545,N_19502);
xnor U20573 (N_20573,N_19742,N_18252);
nand U20574 (N_20574,N_18123,N_18101);
nor U20575 (N_20575,N_17889,N_18659);
xnor U20576 (N_20576,N_18885,N_19863);
nand U20577 (N_20577,N_17773,N_18535);
xor U20578 (N_20578,N_18556,N_18124);
nand U20579 (N_20579,N_18569,N_18161);
and U20580 (N_20580,N_19104,N_19601);
xor U20581 (N_20581,N_18612,N_18234);
nor U20582 (N_20582,N_18920,N_18456);
nand U20583 (N_20583,N_17909,N_17538);
nand U20584 (N_20584,N_19481,N_18605);
nor U20585 (N_20585,N_19862,N_19649);
nor U20586 (N_20586,N_18696,N_19479);
xor U20587 (N_20587,N_18243,N_18966);
or U20588 (N_20588,N_17880,N_18608);
nor U20589 (N_20589,N_17706,N_17936);
nand U20590 (N_20590,N_19100,N_19717);
and U20591 (N_20591,N_19969,N_19669);
and U20592 (N_20592,N_18531,N_18166);
or U20593 (N_20593,N_18333,N_18300);
nand U20594 (N_20594,N_19965,N_18062);
nand U20595 (N_20595,N_18274,N_19683);
nor U20596 (N_20596,N_19077,N_17694);
xnor U20597 (N_20597,N_18198,N_17689);
xor U20598 (N_20598,N_19416,N_19741);
and U20599 (N_20599,N_19634,N_17572);
and U20600 (N_20600,N_18813,N_19872);
and U20601 (N_20601,N_19743,N_18964);
and U20602 (N_20602,N_17523,N_19876);
xor U20603 (N_20603,N_19800,N_18815);
nor U20604 (N_20604,N_19520,N_18266);
or U20605 (N_20605,N_18908,N_19103);
nor U20606 (N_20606,N_18562,N_18351);
xnor U20607 (N_20607,N_17555,N_17716);
nand U20608 (N_20608,N_18429,N_19519);
nor U20609 (N_20609,N_18830,N_17554);
nor U20610 (N_20610,N_18585,N_18424);
xor U20611 (N_20611,N_18076,N_19914);
and U20612 (N_20612,N_19451,N_18526);
and U20613 (N_20613,N_18840,N_19343);
or U20614 (N_20614,N_18987,N_17885);
or U20615 (N_20615,N_18700,N_19931);
or U20616 (N_20616,N_18799,N_18680);
or U20617 (N_20617,N_18473,N_19664);
nand U20618 (N_20618,N_19310,N_19791);
xor U20619 (N_20619,N_17715,N_19323);
nor U20620 (N_20620,N_19662,N_17989);
or U20621 (N_20621,N_18029,N_18865);
nor U20622 (N_20622,N_19171,N_19433);
nor U20623 (N_20623,N_17953,N_17820);
and U20624 (N_20624,N_17772,N_18236);
nor U20625 (N_20625,N_18788,N_18707);
xnor U20626 (N_20626,N_19324,N_19686);
and U20627 (N_20627,N_18375,N_19466);
xor U20628 (N_20628,N_19167,N_18851);
nor U20629 (N_20629,N_18112,N_18326);
xnor U20630 (N_20630,N_18894,N_18657);
and U20631 (N_20631,N_17751,N_17883);
nand U20632 (N_20632,N_19945,N_19185);
nor U20633 (N_20633,N_19909,N_19713);
or U20634 (N_20634,N_19208,N_19827);
nor U20635 (N_20635,N_19391,N_19383);
xor U20636 (N_20636,N_18262,N_17955);
xnor U20637 (N_20637,N_19913,N_17508);
xnor U20638 (N_20638,N_18121,N_19569);
or U20639 (N_20639,N_18806,N_17692);
nor U20640 (N_20640,N_17675,N_19043);
nor U20641 (N_20641,N_18206,N_17687);
xnor U20642 (N_20642,N_19012,N_19402);
or U20643 (N_20643,N_18356,N_18982);
xnor U20644 (N_20644,N_18079,N_18003);
nor U20645 (N_20645,N_18496,N_18687);
or U20646 (N_20646,N_18831,N_19368);
and U20647 (N_20647,N_18621,N_19985);
or U20648 (N_20648,N_18903,N_19981);
xnor U20649 (N_20649,N_19749,N_18727);
nor U20650 (N_20650,N_19134,N_19143);
nor U20651 (N_20651,N_18732,N_17769);
nor U20652 (N_20652,N_18833,N_19948);
and U20653 (N_20653,N_19668,N_17940);
and U20654 (N_20654,N_17603,N_18433);
and U20655 (N_20655,N_19774,N_17746);
or U20656 (N_20656,N_17669,N_17821);
and U20657 (N_20657,N_19127,N_18726);
nand U20658 (N_20658,N_18733,N_19096);
nor U20659 (N_20659,N_19178,N_18408);
nand U20660 (N_20660,N_18484,N_17584);
or U20661 (N_20661,N_19960,N_19589);
xnor U20662 (N_20662,N_18949,N_17778);
nor U20663 (N_20663,N_19631,N_19236);
or U20664 (N_20664,N_18010,N_19472);
and U20665 (N_20665,N_17645,N_19370);
nand U20666 (N_20666,N_17998,N_17935);
nand U20667 (N_20667,N_18502,N_18154);
xnor U20668 (N_20668,N_18619,N_17525);
and U20669 (N_20669,N_19358,N_18748);
nand U20670 (N_20670,N_19667,N_18686);
and U20671 (N_20671,N_17701,N_19769);
and U20672 (N_20672,N_19826,N_19172);
and U20673 (N_20673,N_18924,N_18043);
and U20674 (N_20674,N_19004,N_18993);
nand U20675 (N_20675,N_18921,N_18426);
nand U20676 (N_20676,N_18448,N_19426);
or U20677 (N_20677,N_19703,N_18091);
and U20678 (N_20678,N_19164,N_19898);
nand U20679 (N_20679,N_19258,N_17723);
nand U20680 (N_20680,N_18738,N_18015);
nor U20681 (N_20681,N_19056,N_18812);
nand U20682 (N_20682,N_17828,N_18256);
or U20683 (N_20683,N_17545,N_17776);
or U20684 (N_20684,N_18173,N_19714);
and U20685 (N_20685,N_19396,N_17971);
and U20686 (N_20686,N_18723,N_18916);
xnor U20687 (N_20687,N_19566,N_18716);
and U20688 (N_20688,N_17589,N_18407);
nor U20689 (N_20689,N_18848,N_19415);
nor U20690 (N_20690,N_18804,N_18853);
nand U20691 (N_20691,N_19406,N_19237);
nor U20692 (N_20692,N_19740,N_18404);
or U20693 (N_20693,N_18625,N_17774);
nand U20694 (N_20694,N_19716,N_19915);
nand U20695 (N_20695,N_17847,N_17510);
or U20696 (N_20696,N_18758,N_18020);
nor U20697 (N_20697,N_17802,N_18069);
xor U20698 (N_20698,N_17602,N_19976);
nor U20699 (N_20699,N_17541,N_18611);
and U20700 (N_20700,N_19564,N_18232);
nor U20701 (N_20701,N_19354,N_19319);
nor U20702 (N_20702,N_19734,N_17659);
nand U20703 (N_20703,N_19253,N_19606);
nor U20704 (N_20704,N_18599,N_17678);
xnor U20705 (N_20705,N_18978,N_18571);
or U20706 (N_20706,N_17686,N_19301);
xor U20707 (N_20707,N_18971,N_18349);
or U20708 (N_20708,N_18740,N_17552);
nor U20709 (N_20709,N_18533,N_18957);
xnor U20710 (N_20710,N_19246,N_18688);
nand U20711 (N_20711,N_17945,N_18528);
and U20712 (N_20712,N_19227,N_19709);
nor U20713 (N_20713,N_19557,N_18572);
xor U20714 (N_20714,N_19309,N_19705);
nor U20715 (N_20715,N_19751,N_19470);
or U20716 (N_20716,N_18724,N_18027);
nor U20717 (N_20717,N_19106,N_17615);
xor U20718 (N_20718,N_18702,N_18422);
nand U20719 (N_20719,N_19346,N_17794);
or U20720 (N_20720,N_18598,N_18053);
nand U20721 (N_20721,N_19145,N_17625);
nand U20722 (N_20722,N_19544,N_17965);
nand U20723 (N_20723,N_19748,N_19305);
nor U20724 (N_20724,N_19699,N_19261);
nor U20725 (N_20725,N_17863,N_17547);
and U20726 (N_20726,N_18286,N_19295);
nand U20727 (N_20727,N_19570,N_17557);
and U20728 (N_20728,N_19489,N_19623);
and U20729 (N_20729,N_17990,N_18103);
or U20730 (N_20730,N_19292,N_19063);
nor U20731 (N_20731,N_18118,N_19035);
xor U20732 (N_20732,N_18033,N_17581);
and U20733 (N_20733,N_19684,N_19179);
xor U20734 (N_20734,N_19339,N_18052);
and U20735 (N_20735,N_17677,N_19206);
nand U20736 (N_20736,N_18540,N_18679);
nor U20737 (N_20737,N_19156,N_17976);
or U20738 (N_20738,N_18304,N_19902);
or U20739 (N_20739,N_19332,N_19729);
or U20740 (N_20740,N_17702,N_19910);
or U20741 (N_20741,N_19372,N_19527);
or U20742 (N_20742,N_19359,N_19648);
and U20743 (N_20743,N_18073,N_18994);
nand U20744 (N_20744,N_18228,N_19770);
nand U20745 (N_20745,N_17655,N_18698);
xor U20746 (N_20746,N_19793,N_17514);
nand U20747 (N_20747,N_17925,N_19325);
and U20748 (N_20748,N_19404,N_18919);
or U20749 (N_20749,N_17548,N_17950);
or U20750 (N_20750,N_18588,N_18941);
xor U20751 (N_20751,N_19147,N_17980);
xor U20752 (N_20752,N_17871,N_19113);
and U20753 (N_20753,N_19896,N_19883);
and U20754 (N_20754,N_17933,N_18564);
xor U20755 (N_20755,N_18293,N_18215);
nor U20756 (N_20756,N_19002,N_19592);
or U20757 (N_20757,N_19157,N_19345);
or U20758 (N_20758,N_19936,N_17727);
and U20759 (N_20759,N_17718,N_18068);
nand U20760 (N_20760,N_17642,N_19657);
and U20761 (N_20761,N_19321,N_19690);
nor U20762 (N_20762,N_19874,N_19773);
xnor U20763 (N_20763,N_19861,N_19326);
and U20764 (N_20764,N_19497,N_17918);
and U20765 (N_20765,N_19401,N_19949);
nor U20766 (N_20766,N_19204,N_17516);
xnor U20767 (N_20767,N_18190,N_19313);
and U20768 (N_20768,N_19065,N_19350);
or U20769 (N_20769,N_18269,N_18182);
nand U20770 (N_20770,N_19865,N_18327);
and U20771 (N_20771,N_18860,N_19875);
xor U20772 (N_20772,N_18162,N_17768);
nor U20773 (N_20773,N_17890,N_19093);
nand U20774 (N_20774,N_19646,N_19530);
xnor U20775 (N_20775,N_17537,N_18545);
nor U20776 (N_20776,N_17719,N_18125);
and U20777 (N_20777,N_19786,N_19023);
xor U20778 (N_20778,N_18170,N_19041);
nand U20779 (N_20779,N_19121,N_18174);
or U20780 (N_20780,N_17535,N_18747);
xnor U20781 (N_20781,N_19526,N_18423);
xor U20782 (N_20782,N_18912,N_17569);
nor U20783 (N_20783,N_19210,N_17779);
and U20784 (N_20784,N_17736,N_18381);
xnor U20785 (N_20785,N_19660,N_18845);
and U20786 (N_20786,N_19284,N_19522);
nor U20787 (N_20787,N_18006,N_19822);
or U20788 (N_20788,N_19232,N_18361);
and U20789 (N_20789,N_18146,N_19516);
xnor U20790 (N_20790,N_19057,N_17960);
or U20791 (N_20791,N_18034,N_19438);
xnor U20792 (N_20792,N_17788,N_18088);
xnor U20793 (N_20793,N_19428,N_17534);
xor U20794 (N_20794,N_18403,N_17764);
and U20795 (N_20795,N_19715,N_18938);
xnor U20796 (N_20796,N_18265,N_19109);
and U20797 (N_20797,N_19840,N_18878);
nand U20798 (N_20798,N_18024,N_18156);
and U20799 (N_20799,N_17630,N_18346);
nor U20800 (N_20800,N_18208,N_19075);
or U20801 (N_20801,N_17643,N_19794);
nand U20802 (N_20802,N_18061,N_17588);
xor U20803 (N_20803,N_18586,N_18277);
xnor U20804 (N_20804,N_19133,N_17924);
xnor U20805 (N_20805,N_17544,N_19653);
xnor U20806 (N_20806,N_17712,N_17877);
and U20807 (N_20807,N_17521,N_18046);
or U20808 (N_20808,N_19374,N_18570);
or U20809 (N_20809,N_19753,N_18370);
and U20810 (N_20810,N_17506,N_18165);
xnor U20811 (N_20811,N_18058,N_18904);
nor U20812 (N_20812,N_18685,N_18150);
xnor U20813 (N_20813,N_19816,N_19765);
nand U20814 (N_20814,N_17565,N_18824);
or U20815 (N_20815,N_19355,N_18031);
xor U20816 (N_20816,N_19125,N_19679);
nor U20817 (N_20817,N_17888,N_18524);
and U20818 (N_20818,N_19168,N_19722);
xor U20819 (N_20819,N_19904,N_17721);
nor U20820 (N_20820,N_19099,N_19975);
and U20821 (N_20821,N_18287,N_18194);
nor U20822 (N_20822,N_18463,N_19944);
and U20823 (N_20823,N_19068,N_19640);
nor U20824 (N_20824,N_18209,N_18905);
xnor U20825 (N_20825,N_17540,N_19583);
nand U20826 (N_20826,N_18877,N_19726);
or U20827 (N_20827,N_18057,N_17653);
xor U20828 (N_20828,N_19066,N_17561);
xnor U20829 (N_20829,N_18501,N_17690);
or U20830 (N_20830,N_18651,N_18283);
xnor U20831 (N_20831,N_18936,N_17724);
and U20832 (N_20832,N_19230,N_17948);
nor U20833 (N_20833,N_17758,N_19659);
nand U20834 (N_20834,N_19845,N_18048);
xor U20835 (N_20835,N_19644,N_17926);
and U20836 (N_20836,N_18549,N_17973);
and U20837 (N_20837,N_18107,N_17932);
xor U20838 (N_20838,N_18188,N_17608);
xor U20839 (N_20839,N_19747,N_18263);
nor U20840 (N_20840,N_19187,N_18658);
xnor U20841 (N_20841,N_18972,N_18711);
nand U20842 (N_20842,N_19165,N_17743);
nor U20843 (N_20843,N_17756,N_19356);
or U20844 (N_20844,N_18868,N_19021);
or U20845 (N_20845,N_19386,N_19440);
xor U20846 (N_20846,N_19777,N_19177);
and U20847 (N_20847,N_17703,N_19670);
nand U20848 (N_20848,N_19218,N_19233);
xor U20849 (N_20849,N_18415,N_19894);
xnor U20850 (N_20850,N_19499,N_17810);
or U20851 (N_20851,N_18138,N_19882);
and U20852 (N_20852,N_18201,N_18717);
nand U20853 (N_20853,N_18328,N_17979);
xnor U20854 (N_20854,N_17679,N_19252);
or U20855 (N_20855,N_19635,N_18268);
or U20856 (N_20856,N_18875,N_19364);
nand U20857 (N_20857,N_19128,N_17551);
or U20858 (N_20858,N_19807,N_18272);
nor U20859 (N_20859,N_19071,N_17792);
nand U20860 (N_20860,N_19673,N_18037);
nand U20861 (N_20861,N_18960,N_19262);
nor U20862 (N_20862,N_19153,N_19934);
nor U20863 (N_20863,N_18728,N_19115);
and U20864 (N_20864,N_19196,N_18722);
nand U20865 (N_20865,N_19906,N_19494);
nand U20866 (N_20866,N_19928,N_19818);
and U20867 (N_20867,N_19868,N_19565);
and U20868 (N_20868,N_18041,N_18126);
and U20869 (N_20869,N_18451,N_18537);
or U20870 (N_20870,N_18850,N_19337);
xor U20871 (N_20871,N_19272,N_19506);
nor U20872 (N_20872,N_18662,N_18482);
xnor U20873 (N_20873,N_17661,N_18602);
or U20874 (N_20874,N_18290,N_18464);
or U20875 (N_20875,N_19446,N_18343);
xor U20876 (N_20876,N_19603,N_19918);
nor U20877 (N_20877,N_18663,N_19486);
and U20878 (N_20878,N_17912,N_19543);
nand U20879 (N_20879,N_18071,N_17567);
xnor U20880 (N_20880,N_19930,N_18295);
xnor U20881 (N_20881,N_19462,N_19353);
nor U20882 (N_20882,N_19938,N_19643);
xnor U20883 (N_20883,N_18444,N_18580);
and U20884 (N_20884,N_19571,N_17835);
or U20885 (N_20885,N_18589,N_18618);
xor U20886 (N_20886,N_18084,N_18195);
or U20887 (N_20887,N_17914,N_17709);
nand U20888 (N_20888,N_18405,N_18440);
nor U20889 (N_20889,N_19518,N_17573);
nand U20890 (N_20890,N_19197,N_18406);
nor U20891 (N_20891,N_18392,N_17726);
and U20892 (N_20892,N_18796,N_19229);
nand U20893 (N_20893,N_19424,N_18609);
nand U20894 (N_20894,N_18898,N_19380);
or U20895 (N_20895,N_18884,N_19195);
and U20896 (N_20896,N_19943,N_19105);
nor U20897 (N_20897,N_18267,N_18783);
and U20898 (N_20898,N_17683,N_19418);
nor U20899 (N_20899,N_19836,N_19598);
or U20900 (N_20900,N_19344,N_17996);
and U20901 (N_20901,N_18036,N_19762);
or U20902 (N_20902,N_17558,N_19223);
xnor U20903 (N_20903,N_18518,N_18592);
or U20904 (N_20904,N_18163,N_19448);
or U20905 (N_20905,N_19688,N_19308);
and U20906 (N_20906,N_19552,N_19968);
nor U20907 (N_20907,N_17634,N_17604);
nor U20908 (N_20908,N_18975,N_19804);
xor U20909 (N_20909,N_19090,N_18360);
nor U20910 (N_20910,N_19877,N_18781);
nor U20911 (N_20911,N_19092,N_19342);
or U20912 (N_20912,N_17846,N_17660);
and U20913 (N_20913,N_18012,N_18104);
nand U20914 (N_20914,N_18587,N_17717);
nor U20915 (N_20915,N_18164,N_19079);
nor U20916 (N_20916,N_17646,N_17895);
xnor U20917 (N_20917,N_19152,N_17824);
nor U20918 (N_20918,N_17612,N_18035);
and U20919 (N_20919,N_18387,N_17952);
or U20920 (N_20920,N_18693,N_19351);
or U20921 (N_20921,N_18932,N_17532);
nand U20922 (N_20922,N_19797,N_19288);
and U20923 (N_20923,N_19429,N_18386);
and U20924 (N_20924,N_18739,N_18019);
nand U20925 (N_20925,N_17923,N_19511);
nand U20926 (N_20926,N_19037,N_19070);
xor U20927 (N_20927,N_18416,N_19371);
nand U20928 (N_20928,N_17740,N_19366);
nor U20929 (N_20929,N_19738,N_18650);
nand U20930 (N_20930,N_19843,N_18940);
nor U20931 (N_20931,N_19523,N_19432);
and U20932 (N_20932,N_19678,N_18100);
nand U20933 (N_20933,N_18109,N_18520);
nor U20934 (N_20934,N_18363,N_19973);
nand U20935 (N_20935,N_18774,N_18400);
xor U20936 (N_20936,N_19672,N_18997);
xor U20937 (N_20937,N_17531,N_19932);
nand U20938 (N_20938,N_17759,N_19419);
nor U20939 (N_20939,N_18790,N_18874);
or U20940 (N_20940,N_18914,N_17836);
nand U20941 (N_20941,N_17922,N_18122);
nor U20942 (N_20942,N_18690,N_17674);
or U20943 (N_20943,N_19341,N_18044);
nor U20944 (N_20944,N_19532,N_19445);
or U20945 (N_20945,N_18398,N_18171);
and U20946 (N_20946,N_19907,N_19801);
xnor U20947 (N_20947,N_19549,N_18544);
nand U20948 (N_20948,N_18628,N_18534);
and U20949 (N_20949,N_19306,N_19629);
nor U20950 (N_20950,N_18721,N_19728);
or U20951 (N_20951,N_18950,N_19347);
or U20952 (N_20952,N_18951,N_18042);
nand U20953 (N_20953,N_19595,N_19149);
xnor U20954 (N_20954,N_19214,N_18842);
xnor U20955 (N_20955,N_18357,N_19993);
nor U20956 (N_20956,N_19062,N_18340);
nand U20957 (N_20957,N_17910,N_17861);
xor U20958 (N_20958,N_18669,N_18947);
nor U20959 (N_20959,N_18187,N_19704);
nand U20960 (N_20960,N_18678,N_18465);
nand U20961 (N_20961,N_18483,N_18655);
xnor U20962 (N_20962,N_18965,N_18132);
and U20963 (N_20963,N_18334,N_18060);
xnor U20964 (N_20964,N_18929,N_18816);
xor U20965 (N_20965,N_19658,N_18462);
nor U20966 (N_20966,N_17575,N_19764);
xnor U20967 (N_20967,N_19983,N_18579);
and U20968 (N_20968,N_17882,N_18352);
nand U20969 (N_20969,N_19495,N_18771);
or U20970 (N_20970,N_19315,N_18227);
and U20971 (N_20971,N_19676,N_18431);
and U20972 (N_20972,N_17843,N_18055);
xor U20973 (N_20973,N_17503,N_19897);
nor U20974 (N_20974,N_18863,N_18399);
nor U20975 (N_20975,N_18977,N_19150);
nor U20976 (N_20976,N_17795,N_18594);
xnor U20977 (N_20977,N_18557,N_19508);
nand U20978 (N_20978,N_18837,N_19586);
nand U20979 (N_20979,N_19860,N_18229);
and U20980 (N_20980,N_19369,N_19656);
xor U20981 (N_20981,N_17964,N_19449);
xnor U20982 (N_20982,N_19767,N_19211);
nor U20983 (N_20983,N_19758,N_18737);
nand U20984 (N_20984,N_19538,N_19501);
and U20985 (N_20985,N_18385,N_18946);
and U20986 (N_20986,N_18359,N_17626);
xnor U20987 (N_20987,N_18219,N_19410);
or U20988 (N_20988,N_19929,N_18081);
nor U20989 (N_20989,N_18339,N_19815);
or U20990 (N_20990,N_17640,N_19710);
and U20991 (N_20991,N_19373,N_19510);
nand U20992 (N_20992,N_18149,N_18301);
and U20993 (N_20993,N_19361,N_19923);
and U20994 (N_20994,N_17633,N_19207);
nor U20995 (N_20995,N_19579,N_18910);
xnor U20996 (N_20996,N_18789,N_17763);
xnor U20997 (N_20997,N_19831,N_17606);
and U20998 (N_20998,N_18005,N_19890);
nor U20999 (N_20999,N_17811,N_18968);
nor U21000 (N_21000,N_18793,N_19681);
and U21001 (N_21001,N_19375,N_19755);
and U21002 (N_21002,N_17838,N_18250);
xnor U21003 (N_21003,N_18888,N_18961);
xnor U21004 (N_21004,N_19503,N_18819);
xor U21005 (N_21005,N_18886,N_19847);
xor U21006 (N_21006,N_17974,N_19809);
and U21007 (N_21007,N_19733,N_19692);
nor U21008 (N_21008,N_17647,N_17580);
xnor U21009 (N_21009,N_18089,N_17766);
nand U21010 (N_21010,N_18734,N_19074);
nand U21011 (N_21011,N_19612,N_19005);
or U21012 (N_21012,N_19420,N_17530);
nand U21013 (N_21013,N_18634,N_17982);
nand U21014 (N_21014,N_19768,N_18106);
or U21015 (N_21015,N_18358,N_17517);
nand U21016 (N_21016,N_19248,N_18438);
or U21017 (N_21017,N_17619,N_19957);
nand U21018 (N_21018,N_18504,N_18083);
nor U21019 (N_21019,N_17681,N_19411);
nand U21020 (N_21020,N_18056,N_18225);
and U21021 (N_21021,N_18466,N_19553);
nor U21022 (N_21022,N_19076,N_18311);
or U21023 (N_21023,N_18367,N_19759);
nand U21024 (N_21024,N_19170,N_18551);
and U21025 (N_21025,N_18394,N_19665);
nand U21026 (N_21026,N_19739,N_18388);
and U21027 (N_21027,N_17512,N_18523);
xnor U21028 (N_21028,N_19855,N_19437);
xor U21029 (N_21029,N_17814,N_18847);
or U21030 (N_21030,N_18430,N_19480);
nor U21031 (N_21031,N_18490,N_18481);
xnor U21032 (N_21032,N_18986,N_18493);
nand U21033 (N_21033,N_18192,N_18766);
or U21034 (N_21034,N_17886,N_18338);
nor U21035 (N_21035,N_17621,N_19405);
nand U21036 (N_21036,N_19403,N_17908);
nand U21037 (N_21037,N_19468,N_19019);
nand U21038 (N_21038,N_19720,N_19049);
nand U21039 (N_21039,N_18801,N_19126);
nand U21040 (N_21040,N_18832,N_18638);
or U21041 (N_21041,N_19698,N_17667);
and U21042 (N_21042,N_18054,N_19059);
xnor U21043 (N_21043,N_19636,N_19264);
nand U21044 (N_21044,N_18233,N_19467);
and U21045 (N_21045,N_19546,N_18419);
xnor U21046 (N_21046,N_18959,N_19642);
and U21047 (N_21047,N_19802,N_17951);
nand U21048 (N_21048,N_18317,N_18178);
or U21049 (N_21049,N_18382,N_19972);
nand U21050 (N_21050,N_17613,N_17637);
xnor U21051 (N_21051,N_19584,N_18151);
or U21052 (N_21052,N_17870,N_17632);
xor U21053 (N_21053,N_18183,N_19422);
nor U21054 (N_21054,N_18260,N_17943);
nand U21055 (N_21055,N_19032,N_19746);
or U21056 (N_21056,N_19073,N_17704);
or U21057 (N_21057,N_19834,N_17697);
and U21058 (N_21058,N_18808,N_17599);
nor U21059 (N_21059,N_18883,N_18785);
xnor U21060 (N_21060,N_19269,N_19593);
or U21061 (N_21061,N_18475,N_18610);
nand U21062 (N_21062,N_18896,N_17657);
nor U21063 (N_21063,N_18749,N_18039);
xnor U21064 (N_21064,N_17711,N_17579);
and U21065 (N_21065,N_17946,N_17563);
nand U21066 (N_21066,N_17735,N_18032);
nand U21067 (N_21067,N_18859,N_17542);
nor U21068 (N_21068,N_17815,N_18601);
nor U21069 (N_21069,N_18622,N_18380);
and U21070 (N_21070,N_19610,N_19829);
xnor U21071 (N_21071,N_19961,N_18995);
xor U21072 (N_21072,N_18695,N_19916);
xor U21073 (N_21073,N_17749,N_19940);
nor U21074 (N_21074,N_19190,N_18000);
xnor U21075 (N_21075,N_18654,N_17515);
and U21076 (N_21076,N_18040,N_18169);
and U21077 (N_21077,N_18996,N_19917);
nor U21078 (N_21078,N_17842,N_18607);
xor U21079 (N_21079,N_18157,N_18241);
xnor U21080 (N_21080,N_19412,N_18280);
and U21081 (N_21081,N_18582,N_17845);
nor U21082 (N_21082,N_19485,N_19413);
xor U21083 (N_21083,N_19238,N_19987);
or U21084 (N_21084,N_18013,N_18559);
nor U21085 (N_21085,N_19247,N_17797);
and U21086 (N_21086,N_18063,N_17852);
nand U21087 (N_21087,N_17698,N_18141);
and U21088 (N_21088,N_19183,N_18134);
and U21089 (N_21089,N_18342,N_19135);
and U21090 (N_21090,N_19039,N_17920);
nand U21091 (N_21091,N_18928,N_17999);
or U21092 (N_21092,N_19441,N_17559);
nor U21093 (N_21093,N_19941,N_18432);
xnor U21094 (N_21094,N_19050,N_17881);
or U21095 (N_21095,N_18319,N_19140);
nand U21096 (N_21096,N_17806,N_18511);
or U21097 (N_21097,N_19275,N_18773);
and U21098 (N_21098,N_17582,N_17800);
xnor U21099 (N_21099,N_18713,N_17585);
or U21100 (N_21100,N_19830,N_18396);
nand U21101 (N_21101,N_17931,N_19551);
nand U21102 (N_21102,N_18454,N_17522);
nand U21103 (N_21103,N_17714,N_19119);
xnor U21104 (N_21104,N_17725,N_19498);
nand U21105 (N_21105,N_19870,N_18770);
xnor U21106 (N_21106,N_18207,N_18828);
nor U21107 (N_21107,N_19387,N_19013);
or U21108 (N_21108,N_17988,N_17560);
and U21109 (N_21109,N_19015,N_17968);
or U21110 (N_21110,N_19457,N_19964);
or U21111 (N_21111,N_17787,N_17786);
nand U21112 (N_21112,N_18763,N_18211);
xor U21113 (N_21113,N_17827,N_18507);
xor U21114 (N_21114,N_17699,N_18714);
and U21115 (N_21115,N_17901,N_18446);
nor U21116 (N_21116,N_17654,N_18324);
or U21117 (N_21117,N_19124,N_19436);
or U21118 (N_21118,N_18503,N_19849);
nand U21119 (N_21119,N_19040,N_19787);
xor U21120 (N_21120,N_18028,N_18981);
nand U21121 (N_21121,N_17710,N_19201);
and U21122 (N_21122,N_18276,N_19048);
xor U21123 (N_21123,N_19385,N_19024);
xor U21124 (N_21124,N_19539,N_17789);
nand U21125 (N_21125,N_18264,N_18402);
or U21126 (N_21126,N_18449,N_18238);
xor U21127 (N_21127,N_18495,N_18989);
nand U21128 (N_21128,N_17840,N_18498);
nand U21129 (N_21129,N_19988,N_17738);
nor U21130 (N_21130,N_19633,N_19903);
and U21131 (N_21131,N_19783,N_19052);
and U21132 (N_21132,N_18336,N_17720);
xor U21133 (N_21133,N_18337,N_18555);
nor U21134 (N_21134,N_18202,N_18167);
and U21135 (N_21135,N_19588,N_19322);
and U21136 (N_21136,N_18335,N_17705);
nand U21137 (N_21137,N_18251,N_17676);
or U21138 (N_21138,N_17638,N_19535);
and U21139 (N_21139,N_18822,N_18362);
and U21140 (N_21140,N_19046,N_17511);
or U21141 (N_21141,N_18255,N_18284);
nand U21142 (N_21142,N_18768,N_18120);
and U21143 (N_21143,N_19330,N_19260);
nand U21144 (N_21144,N_18344,N_19469);
nand U21145 (N_21145,N_19982,N_18130);
nand U21146 (N_21146,N_17564,N_17929);
and U21147 (N_21147,N_17658,N_19504);
and U21148 (N_21148,N_19407,N_18453);
nand U21149 (N_21149,N_17865,N_19400);
nand U21150 (N_21150,N_18092,N_18320);
xnor U21151 (N_21151,N_18004,N_19175);
or U21152 (N_21152,N_17639,N_19737);
nand U21153 (N_21153,N_19465,N_18893);
nor U21154 (N_21154,N_19819,N_18376);
nor U21155 (N_21155,N_18247,N_19701);
xnor U21156 (N_21156,N_18805,N_19950);
nand U21157 (N_21157,N_19425,N_18876);
xnor U21158 (N_21158,N_18901,N_18258);
xor U21159 (N_21159,N_19563,N_18566);
xnor U21160 (N_21160,N_17570,N_18615);
nor U21161 (N_21161,N_19572,N_19974);
or U21162 (N_21162,N_19574,N_18271);
xnor U21163 (N_21163,N_17961,N_19708);
and U21164 (N_21164,N_18744,N_18425);
and U21165 (N_21165,N_17610,N_19775);
xor U21166 (N_21166,N_19887,N_17855);
xnor U21167 (N_21167,N_18742,N_19625);
xor U21168 (N_21168,N_17733,N_17819);
and U21169 (N_21169,N_17967,N_19582);
xor U21170 (N_21170,N_19053,N_18203);
or U21171 (N_21171,N_19296,N_19312);
and U21172 (N_21172,N_19590,N_18220);
and U21173 (N_21173,N_17641,N_19823);
or U21174 (N_21174,N_18857,N_18887);
nor U21175 (N_21175,N_18925,N_17969);
or U21176 (N_21176,N_17834,N_18525);
nand U21177 (N_21177,N_18510,N_18159);
xor U21178 (N_21178,N_17977,N_17927);
nand U21179 (N_21179,N_19493,N_19575);
xnor U21180 (N_21180,N_19379,N_19784);
nor U21181 (N_21181,N_19766,N_18321);
or U21182 (N_21182,N_18145,N_19727);
nand U21183 (N_21183,N_18666,N_17528);
and U21184 (N_21184,N_19279,N_18757);
or U21185 (N_21185,N_18002,N_17762);
or U21186 (N_21186,N_18861,N_19026);
nand U21187 (N_21187,N_18458,N_19222);
xor U21188 (N_21188,N_18366,N_19604);
and U21189 (N_21189,N_18492,N_18980);
nand U21190 (N_21190,N_19144,N_19824);
and U21191 (N_21191,N_19837,N_18471);
nand U21192 (N_21192,N_18371,N_19054);
nand U21193 (N_21193,N_19663,N_19905);
or U21194 (N_21194,N_18353,N_18577);
nand U21195 (N_21195,N_18803,N_18497);
nor U21196 (N_21196,N_18153,N_18558);
or U21197 (N_21197,N_18791,N_19482);
xor U21198 (N_21198,N_17684,N_17894);
and U21199 (N_21199,N_17985,N_19255);
and U21200 (N_21200,N_19825,N_19408);
nor U21201 (N_21201,N_19388,N_17876);
or U21202 (N_21202,N_19833,N_18671);
nor U21203 (N_21203,N_18160,N_18623);
and U21204 (N_21204,N_19159,N_19674);
and U21205 (N_21205,N_18567,N_18364);
xor U21206 (N_21206,N_18553,N_18377);
and U21207 (N_21207,N_19189,N_18668);
xor U21208 (N_21208,N_19885,N_19850);
nand U21209 (N_21209,N_18913,N_18030);
nand U21210 (N_21210,N_17790,N_18307);
or U21211 (N_21211,N_18253,N_17983);
xor U21212 (N_21212,N_18753,N_19008);
and U21213 (N_21213,N_18640,N_18296);
xor U21214 (N_21214,N_18854,N_18918);
xor U21215 (N_21215,N_18025,N_19007);
and U21216 (N_21216,N_19423,N_19051);
nor U21217 (N_21217,N_18583,N_18204);
nand U21218 (N_21218,N_17859,N_18595);
and U21219 (N_21219,N_18273,N_19114);
nor U21220 (N_21220,N_19567,N_18809);
nand U21221 (N_21221,N_18108,N_18509);
nor U21222 (N_21222,N_19515,N_17597);
nand U21223 (N_21223,N_18519,N_17627);
nand U21224 (N_21224,N_18539,N_18897);
or U21225 (N_21225,N_19605,N_19696);
xor U21226 (N_21226,N_17624,N_18140);
nand U21227 (N_21227,N_19399,N_18880);
nand U21228 (N_21228,N_19176,N_19131);
or U21229 (N_21229,N_18798,N_19038);
and U21230 (N_21230,N_18683,N_19299);
nor U21231 (N_21231,N_18045,N_18935);
or U21232 (N_21232,N_19273,N_17596);
or U21233 (N_21233,N_18116,N_18152);
nand U21234 (N_21234,N_19577,N_18794);
and U21235 (N_21235,N_17616,N_18705);
or U21236 (N_21236,N_19088,N_19376);
nand U21237 (N_21237,N_19137,N_19224);
nand U21238 (N_21238,N_19978,N_19795);
or U21239 (N_21239,N_18552,N_18316);
nand U21240 (N_21240,N_19857,N_18529);
xor U21241 (N_21241,N_19512,N_18730);
and U21242 (N_21242,N_18318,N_19239);
nor U21243 (N_21243,N_19528,N_19548);
nand U21244 (N_21244,N_18849,N_19085);
or U21245 (N_21245,N_18098,N_18681);
or U21246 (N_21246,N_18718,N_18934);
xnor U21247 (N_21247,N_18694,N_19718);
or U21248 (N_21248,N_18515,N_18014);
or U21249 (N_21249,N_19348,N_19181);
xnor U21250 (N_21250,N_18163,N_17950);
nand U21251 (N_21251,N_19971,N_18068);
or U21252 (N_21252,N_19801,N_17788);
nand U21253 (N_21253,N_17516,N_18899);
nand U21254 (N_21254,N_17875,N_17579);
and U21255 (N_21255,N_19203,N_17750);
nand U21256 (N_21256,N_18028,N_19099);
nor U21257 (N_21257,N_18748,N_18349);
or U21258 (N_21258,N_17727,N_17759);
nor U21259 (N_21259,N_17661,N_19827);
or U21260 (N_21260,N_18268,N_18311);
xnor U21261 (N_21261,N_19503,N_19561);
xnor U21262 (N_21262,N_17942,N_19091);
or U21263 (N_21263,N_18281,N_19586);
and U21264 (N_21264,N_18922,N_18264);
or U21265 (N_21265,N_17894,N_19660);
nor U21266 (N_21266,N_19740,N_19884);
or U21267 (N_21267,N_19163,N_17828);
and U21268 (N_21268,N_19754,N_19960);
nor U21269 (N_21269,N_17678,N_19801);
nor U21270 (N_21270,N_18486,N_18061);
and U21271 (N_21271,N_19307,N_18321);
nor U21272 (N_21272,N_18624,N_17882);
and U21273 (N_21273,N_18503,N_18339);
and U21274 (N_21274,N_18803,N_17763);
nor U21275 (N_21275,N_18702,N_18175);
and U21276 (N_21276,N_18700,N_19586);
xnor U21277 (N_21277,N_17819,N_18989);
nand U21278 (N_21278,N_19341,N_19395);
xnor U21279 (N_21279,N_17830,N_19848);
nand U21280 (N_21280,N_19779,N_18693);
xnor U21281 (N_21281,N_19688,N_19665);
nor U21282 (N_21282,N_17993,N_19378);
or U21283 (N_21283,N_19614,N_19542);
or U21284 (N_21284,N_17607,N_19001);
xnor U21285 (N_21285,N_19769,N_19286);
nor U21286 (N_21286,N_19361,N_17992);
and U21287 (N_21287,N_17839,N_17644);
or U21288 (N_21288,N_18628,N_19195);
or U21289 (N_21289,N_19608,N_18491);
xor U21290 (N_21290,N_18029,N_17842);
nor U21291 (N_21291,N_19901,N_19018);
nand U21292 (N_21292,N_19393,N_19258);
nor U21293 (N_21293,N_19476,N_19024);
xnor U21294 (N_21294,N_19221,N_19840);
nand U21295 (N_21295,N_18329,N_19432);
xnor U21296 (N_21296,N_19645,N_19206);
nor U21297 (N_21297,N_18951,N_17983);
xnor U21298 (N_21298,N_18257,N_18048);
or U21299 (N_21299,N_19178,N_17906);
or U21300 (N_21300,N_19065,N_17907);
and U21301 (N_21301,N_17947,N_19007);
nor U21302 (N_21302,N_18311,N_17943);
nand U21303 (N_21303,N_18118,N_17775);
nor U21304 (N_21304,N_18279,N_19351);
or U21305 (N_21305,N_17955,N_19222);
and U21306 (N_21306,N_19224,N_17735);
xor U21307 (N_21307,N_17795,N_19873);
or U21308 (N_21308,N_19743,N_18696);
nand U21309 (N_21309,N_18072,N_17968);
nand U21310 (N_21310,N_17512,N_19149);
xor U21311 (N_21311,N_17570,N_18556);
and U21312 (N_21312,N_19619,N_17510);
or U21313 (N_21313,N_18465,N_19794);
and U21314 (N_21314,N_19025,N_19794);
nand U21315 (N_21315,N_18883,N_18212);
and U21316 (N_21316,N_19058,N_18705);
and U21317 (N_21317,N_17656,N_18139);
and U21318 (N_21318,N_17852,N_18665);
nand U21319 (N_21319,N_19235,N_19496);
nor U21320 (N_21320,N_18115,N_17629);
and U21321 (N_21321,N_19975,N_17770);
or U21322 (N_21322,N_19873,N_18641);
or U21323 (N_21323,N_19768,N_19556);
or U21324 (N_21324,N_18015,N_18652);
and U21325 (N_21325,N_19471,N_18312);
xnor U21326 (N_21326,N_18604,N_17627);
and U21327 (N_21327,N_19847,N_18630);
and U21328 (N_21328,N_17858,N_18526);
nand U21329 (N_21329,N_19890,N_18786);
or U21330 (N_21330,N_18922,N_18533);
and U21331 (N_21331,N_19118,N_19928);
nor U21332 (N_21332,N_18561,N_18792);
nand U21333 (N_21333,N_18702,N_18253);
nor U21334 (N_21334,N_18532,N_19677);
xnor U21335 (N_21335,N_19449,N_19076);
and U21336 (N_21336,N_18966,N_19000);
and U21337 (N_21337,N_17709,N_18596);
and U21338 (N_21338,N_18579,N_18528);
nand U21339 (N_21339,N_18293,N_17548);
nand U21340 (N_21340,N_19947,N_18058);
or U21341 (N_21341,N_18034,N_18853);
nand U21342 (N_21342,N_18138,N_17850);
nand U21343 (N_21343,N_19236,N_19054);
nor U21344 (N_21344,N_17689,N_17937);
nand U21345 (N_21345,N_19969,N_18821);
and U21346 (N_21346,N_17883,N_19676);
nor U21347 (N_21347,N_19534,N_17886);
nor U21348 (N_21348,N_17806,N_18758);
nor U21349 (N_21349,N_17964,N_18034);
nor U21350 (N_21350,N_17830,N_18770);
xor U21351 (N_21351,N_19097,N_18358);
or U21352 (N_21352,N_19002,N_19601);
and U21353 (N_21353,N_19732,N_17502);
and U21354 (N_21354,N_18710,N_18838);
or U21355 (N_21355,N_17890,N_19770);
xor U21356 (N_21356,N_18226,N_19218);
nor U21357 (N_21357,N_17643,N_18758);
xnor U21358 (N_21358,N_19017,N_19988);
xor U21359 (N_21359,N_19136,N_18074);
or U21360 (N_21360,N_17609,N_19959);
nand U21361 (N_21361,N_19592,N_17776);
and U21362 (N_21362,N_19420,N_19522);
nand U21363 (N_21363,N_18134,N_18903);
nand U21364 (N_21364,N_18683,N_19792);
nand U21365 (N_21365,N_17855,N_19956);
xnor U21366 (N_21366,N_18388,N_18943);
or U21367 (N_21367,N_17932,N_19735);
xor U21368 (N_21368,N_18094,N_19014);
nor U21369 (N_21369,N_18298,N_19234);
and U21370 (N_21370,N_17856,N_19672);
or U21371 (N_21371,N_19560,N_17609);
or U21372 (N_21372,N_19905,N_19490);
and U21373 (N_21373,N_17933,N_18121);
nand U21374 (N_21374,N_18898,N_19448);
or U21375 (N_21375,N_19642,N_17909);
or U21376 (N_21376,N_19526,N_19336);
and U21377 (N_21377,N_19691,N_19332);
xnor U21378 (N_21378,N_19538,N_18249);
xor U21379 (N_21379,N_18391,N_17552);
or U21380 (N_21380,N_17648,N_18062);
or U21381 (N_21381,N_17583,N_17685);
or U21382 (N_21382,N_17943,N_19924);
and U21383 (N_21383,N_19174,N_18328);
nand U21384 (N_21384,N_19144,N_17527);
xor U21385 (N_21385,N_18283,N_18257);
or U21386 (N_21386,N_19874,N_17939);
xor U21387 (N_21387,N_18262,N_19016);
nand U21388 (N_21388,N_19656,N_18248);
and U21389 (N_21389,N_18473,N_19757);
nor U21390 (N_21390,N_19556,N_19791);
nand U21391 (N_21391,N_19734,N_19306);
or U21392 (N_21392,N_19804,N_19242);
or U21393 (N_21393,N_17685,N_19024);
nor U21394 (N_21394,N_18589,N_17972);
or U21395 (N_21395,N_18016,N_18039);
nor U21396 (N_21396,N_19132,N_19594);
xor U21397 (N_21397,N_19549,N_17707);
or U21398 (N_21398,N_18274,N_19294);
and U21399 (N_21399,N_18255,N_18219);
nor U21400 (N_21400,N_18609,N_17958);
or U21401 (N_21401,N_19322,N_19143);
xnor U21402 (N_21402,N_18405,N_19314);
nor U21403 (N_21403,N_17543,N_19165);
nand U21404 (N_21404,N_19282,N_18518);
and U21405 (N_21405,N_19340,N_19898);
and U21406 (N_21406,N_19461,N_18895);
or U21407 (N_21407,N_17503,N_18725);
or U21408 (N_21408,N_18273,N_17607);
xnor U21409 (N_21409,N_18076,N_19368);
nand U21410 (N_21410,N_19065,N_18031);
and U21411 (N_21411,N_17896,N_18146);
nand U21412 (N_21412,N_19188,N_17772);
nand U21413 (N_21413,N_19679,N_18238);
or U21414 (N_21414,N_17532,N_18360);
nand U21415 (N_21415,N_18249,N_19313);
and U21416 (N_21416,N_18123,N_18625);
xnor U21417 (N_21417,N_18402,N_18168);
nor U21418 (N_21418,N_19581,N_19650);
nor U21419 (N_21419,N_17982,N_17575);
nor U21420 (N_21420,N_19888,N_18508);
nor U21421 (N_21421,N_17997,N_19218);
nand U21422 (N_21422,N_17763,N_19312);
or U21423 (N_21423,N_18269,N_18825);
or U21424 (N_21424,N_17956,N_19436);
or U21425 (N_21425,N_18059,N_17512);
or U21426 (N_21426,N_17569,N_17802);
nor U21427 (N_21427,N_18456,N_19418);
nand U21428 (N_21428,N_17545,N_19823);
or U21429 (N_21429,N_18913,N_19245);
nand U21430 (N_21430,N_18810,N_19208);
or U21431 (N_21431,N_18452,N_19856);
nor U21432 (N_21432,N_17718,N_19513);
xnor U21433 (N_21433,N_18293,N_18617);
or U21434 (N_21434,N_18305,N_18761);
xnor U21435 (N_21435,N_18312,N_18587);
xor U21436 (N_21436,N_18849,N_18503);
nor U21437 (N_21437,N_19541,N_19725);
nand U21438 (N_21438,N_17933,N_19236);
nor U21439 (N_21439,N_19582,N_18152);
xnor U21440 (N_21440,N_17709,N_18713);
and U21441 (N_21441,N_18840,N_19915);
xnor U21442 (N_21442,N_18147,N_19192);
nand U21443 (N_21443,N_18242,N_19524);
nor U21444 (N_21444,N_19817,N_18998);
nand U21445 (N_21445,N_17994,N_17901);
nand U21446 (N_21446,N_19882,N_17820);
or U21447 (N_21447,N_19354,N_19309);
and U21448 (N_21448,N_17510,N_18422);
nand U21449 (N_21449,N_17789,N_19603);
nor U21450 (N_21450,N_18434,N_17947);
nor U21451 (N_21451,N_18702,N_18212);
xor U21452 (N_21452,N_19984,N_18096);
nand U21453 (N_21453,N_18094,N_19605);
nand U21454 (N_21454,N_17597,N_17847);
nand U21455 (N_21455,N_19095,N_18430);
xnor U21456 (N_21456,N_19305,N_19921);
and U21457 (N_21457,N_17942,N_19135);
or U21458 (N_21458,N_17500,N_19074);
nand U21459 (N_21459,N_17947,N_17604);
nor U21460 (N_21460,N_18719,N_19257);
or U21461 (N_21461,N_18259,N_18320);
nor U21462 (N_21462,N_18101,N_18321);
nor U21463 (N_21463,N_18136,N_18952);
nand U21464 (N_21464,N_19557,N_18300);
xor U21465 (N_21465,N_18873,N_19797);
nor U21466 (N_21466,N_19924,N_19990);
xor U21467 (N_21467,N_18727,N_19410);
or U21468 (N_21468,N_19211,N_18297);
or U21469 (N_21469,N_18562,N_17800);
xnor U21470 (N_21470,N_18111,N_19438);
or U21471 (N_21471,N_19709,N_19922);
and U21472 (N_21472,N_18043,N_18939);
and U21473 (N_21473,N_17793,N_19711);
and U21474 (N_21474,N_19117,N_18910);
and U21475 (N_21475,N_18922,N_18342);
or U21476 (N_21476,N_18968,N_19641);
nor U21477 (N_21477,N_18796,N_19971);
xor U21478 (N_21478,N_17515,N_18422);
and U21479 (N_21479,N_19705,N_17938);
or U21480 (N_21480,N_17655,N_18023);
or U21481 (N_21481,N_18787,N_17554);
or U21482 (N_21482,N_19758,N_19202);
nor U21483 (N_21483,N_18515,N_19143);
xnor U21484 (N_21484,N_19516,N_18499);
nand U21485 (N_21485,N_17545,N_19717);
or U21486 (N_21486,N_19223,N_18189);
nand U21487 (N_21487,N_19912,N_17552);
nand U21488 (N_21488,N_19938,N_18096);
and U21489 (N_21489,N_19807,N_18790);
nor U21490 (N_21490,N_19005,N_19968);
nor U21491 (N_21491,N_19886,N_18414);
nor U21492 (N_21492,N_18714,N_17814);
nand U21493 (N_21493,N_18344,N_19868);
nor U21494 (N_21494,N_17799,N_18360);
xnor U21495 (N_21495,N_18493,N_19289);
nand U21496 (N_21496,N_18815,N_19601);
xnor U21497 (N_21497,N_19158,N_19673);
nor U21498 (N_21498,N_18715,N_18675);
xor U21499 (N_21499,N_18869,N_19165);
xnor U21500 (N_21500,N_18808,N_18114);
nor U21501 (N_21501,N_18010,N_18997);
or U21502 (N_21502,N_18971,N_19740);
or U21503 (N_21503,N_17692,N_17662);
xor U21504 (N_21504,N_18157,N_18297);
or U21505 (N_21505,N_19772,N_17947);
xor U21506 (N_21506,N_18657,N_19372);
or U21507 (N_21507,N_18191,N_18880);
or U21508 (N_21508,N_18354,N_18923);
nor U21509 (N_21509,N_17658,N_19474);
or U21510 (N_21510,N_18028,N_18933);
nor U21511 (N_21511,N_17571,N_18642);
nor U21512 (N_21512,N_18527,N_18793);
or U21513 (N_21513,N_19612,N_18874);
or U21514 (N_21514,N_18563,N_19531);
xnor U21515 (N_21515,N_18476,N_17844);
nor U21516 (N_21516,N_18467,N_19070);
nand U21517 (N_21517,N_18471,N_18280);
nand U21518 (N_21518,N_18187,N_19051);
nor U21519 (N_21519,N_18342,N_18939);
nor U21520 (N_21520,N_19864,N_18771);
xnor U21521 (N_21521,N_19171,N_19317);
nand U21522 (N_21522,N_17952,N_18785);
nand U21523 (N_21523,N_19057,N_17509);
nor U21524 (N_21524,N_18774,N_17550);
and U21525 (N_21525,N_17862,N_18427);
nand U21526 (N_21526,N_17867,N_19806);
and U21527 (N_21527,N_17699,N_18608);
or U21528 (N_21528,N_19950,N_19594);
and U21529 (N_21529,N_19585,N_19114);
or U21530 (N_21530,N_17852,N_18808);
and U21531 (N_21531,N_18844,N_19871);
or U21532 (N_21532,N_17877,N_18963);
xor U21533 (N_21533,N_19160,N_18857);
or U21534 (N_21534,N_18117,N_19051);
and U21535 (N_21535,N_19780,N_18918);
nand U21536 (N_21536,N_18696,N_18814);
xnor U21537 (N_21537,N_19383,N_17838);
nor U21538 (N_21538,N_18415,N_19380);
nor U21539 (N_21539,N_19135,N_18493);
and U21540 (N_21540,N_17916,N_18943);
nor U21541 (N_21541,N_18652,N_18351);
nand U21542 (N_21542,N_19386,N_19206);
and U21543 (N_21543,N_17727,N_18839);
nor U21544 (N_21544,N_19787,N_18357);
or U21545 (N_21545,N_19839,N_18416);
and U21546 (N_21546,N_18502,N_17636);
and U21547 (N_21547,N_19816,N_19826);
nand U21548 (N_21548,N_17652,N_18508);
nand U21549 (N_21549,N_19622,N_17972);
nor U21550 (N_21550,N_19620,N_18991);
nand U21551 (N_21551,N_19509,N_18464);
or U21552 (N_21552,N_18729,N_18620);
xnor U21553 (N_21553,N_18503,N_18809);
nand U21554 (N_21554,N_19858,N_19272);
and U21555 (N_21555,N_17943,N_18375);
xnor U21556 (N_21556,N_17550,N_18954);
and U21557 (N_21557,N_18360,N_19380);
or U21558 (N_21558,N_18639,N_19743);
and U21559 (N_21559,N_19927,N_19547);
nand U21560 (N_21560,N_19558,N_18859);
and U21561 (N_21561,N_19954,N_18769);
nor U21562 (N_21562,N_18473,N_17619);
xor U21563 (N_21563,N_17920,N_19805);
and U21564 (N_21564,N_17881,N_18288);
nor U21565 (N_21565,N_19187,N_17635);
or U21566 (N_21566,N_18408,N_19036);
nand U21567 (N_21567,N_19791,N_19104);
and U21568 (N_21568,N_18833,N_19570);
nor U21569 (N_21569,N_19192,N_19232);
and U21570 (N_21570,N_19878,N_18557);
and U21571 (N_21571,N_18467,N_18147);
nor U21572 (N_21572,N_19144,N_19372);
or U21573 (N_21573,N_17504,N_18113);
nor U21574 (N_21574,N_17898,N_18764);
xor U21575 (N_21575,N_19111,N_19882);
nand U21576 (N_21576,N_19841,N_18243);
xnor U21577 (N_21577,N_19436,N_17949);
or U21578 (N_21578,N_19555,N_19305);
nor U21579 (N_21579,N_19693,N_18150);
and U21580 (N_21580,N_18444,N_19202);
or U21581 (N_21581,N_18253,N_17709);
xnor U21582 (N_21582,N_19417,N_17692);
or U21583 (N_21583,N_17669,N_18072);
xnor U21584 (N_21584,N_18198,N_18213);
or U21585 (N_21585,N_18926,N_18779);
and U21586 (N_21586,N_19075,N_19186);
and U21587 (N_21587,N_18967,N_19062);
nand U21588 (N_21588,N_18006,N_18321);
xnor U21589 (N_21589,N_19017,N_19046);
nand U21590 (N_21590,N_18880,N_19215);
or U21591 (N_21591,N_19760,N_19951);
and U21592 (N_21592,N_18289,N_17652);
nand U21593 (N_21593,N_17509,N_18036);
xor U21594 (N_21594,N_19739,N_18195);
and U21595 (N_21595,N_19193,N_19941);
and U21596 (N_21596,N_19684,N_18893);
nor U21597 (N_21597,N_17670,N_19719);
nand U21598 (N_21598,N_18272,N_18285);
xnor U21599 (N_21599,N_19799,N_17901);
or U21600 (N_21600,N_19370,N_19638);
xor U21601 (N_21601,N_18434,N_19893);
and U21602 (N_21602,N_18103,N_19775);
xnor U21603 (N_21603,N_19936,N_18714);
and U21604 (N_21604,N_18146,N_19481);
nor U21605 (N_21605,N_18570,N_17648);
and U21606 (N_21606,N_18268,N_19943);
nand U21607 (N_21607,N_19164,N_18405);
or U21608 (N_21608,N_18606,N_18593);
xor U21609 (N_21609,N_17934,N_18555);
and U21610 (N_21610,N_19244,N_19605);
nand U21611 (N_21611,N_19030,N_18623);
nor U21612 (N_21612,N_19159,N_17624);
or U21613 (N_21613,N_18331,N_19566);
or U21614 (N_21614,N_18948,N_18127);
nand U21615 (N_21615,N_19065,N_17962);
nor U21616 (N_21616,N_18056,N_18998);
nand U21617 (N_21617,N_18000,N_19522);
xor U21618 (N_21618,N_18210,N_18078);
or U21619 (N_21619,N_17960,N_17841);
xnor U21620 (N_21620,N_18838,N_17821);
and U21621 (N_21621,N_19211,N_18160);
xnor U21622 (N_21622,N_18689,N_18761);
nand U21623 (N_21623,N_17707,N_19459);
nand U21624 (N_21624,N_17658,N_19238);
nand U21625 (N_21625,N_18464,N_19047);
xnor U21626 (N_21626,N_19934,N_19009);
nand U21627 (N_21627,N_19592,N_19905);
or U21628 (N_21628,N_18511,N_18383);
nor U21629 (N_21629,N_19871,N_19463);
nor U21630 (N_21630,N_18407,N_17918);
or U21631 (N_21631,N_19746,N_17684);
nor U21632 (N_21632,N_17550,N_17831);
or U21633 (N_21633,N_19670,N_17505);
nand U21634 (N_21634,N_19013,N_17727);
xnor U21635 (N_21635,N_18302,N_18385);
nand U21636 (N_21636,N_18914,N_17996);
or U21637 (N_21637,N_17881,N_18295);
xor U21638 (N_21638,N_17734,N_18515);
nand U21639 (N_21639,N_19170,N_17809);
nor U21640 (N_21640,N_17526,N_18989);
or U21641 (N_21641,N_17712,N_18326);
or U21642 (N_21642,N_19274,N_19788);
nand U21643 (N_21643,N_18286,N_19104);
nor U21644 (N_21644,N_19374,N_18006);
and U21645 (N_21645,N_17559,N_19048);
or U21646 (N_21646,N_18866,N_19055);
or U21647 (N_21647,N_17592,N_18493);
or U21648 (N_21648,N_19728,N_19640);
nor U21649 (N_21649,N_19223,N_18920);
nand U21650 (N_21650,N_17917,N_18581);
nor U21651 (N_21651,N_17896,N_19788);
or U21652 (N_21652,N_19274,N_19548);
nand U21653 (N_21653,N_18488,N_17669);
or U21654 (N_21654,N_19135,N_18431);
xor U21655 (N_21655,N_17655,N_18464);
nand U21656 (N_21656,N_19208,N_18466);
and U21657 (N_21657,N_19013,N_18700);
nand U21658 (N_21658,N_18725,N_17757);
and U21659 (N_21659,N_19399,N_17712);
and U21660 (N_21660,N_19505,N_19823);
or U21661 (N_21661,N_19300,N_17586);
nor U21662 (N_21662,N_18005,N_18310);
nand U21663 (N_21663,N_18703,N_18441);
xnor U21664 (N_21664,N_18517,N_17876);
nor U21665 (N_21665,N_18926,N_18906);
nor U21666 (N_21666,N_18706,N_19277);
xor U21667 (N_21667,N_17735,N_19480);
and U21668 (N_21668,N_18961,N_19141);
xnor U21669 (N_21669,N_18611,N_19813);
nand U21670 (N_21670,N_19771,N_18129);
nand U21671 (N_21671,N_19162,N_18939);
or U21672 (N_21672,N_18098,N_18056);
nor U21673 (N_21673,N_17703,N_18332);
nand U21674 (N_21674,N_17963,N_17744);
nor U21675 (N_21675,N_18132,N_18800);
nor U21676 (N_21676,N_18784,N_19842);
nor U21677 (N_21677,N_19412,N_19884);
or U21678 (N_21678,N_19554,N_18780);
nand U21679 (N_21679,N_18535,N_18953);
and U21680 (N_21680,N_19316,N_19408);
xnor U21681 (N_21681,N_17928,N_18594);
nor U21682 (N_21682,N_18257,N_19054);
nand U21683 (N_21683,N_18435,N_18577);
nor U21684 (N_21684,N_19501,N_19287);
nand U21685 (N_21685,N_18269,N_19606);
xor U21686 (N_21686,N_19094,N_18662);
nor U21687 (N_21687,N_19580,N_19052);
or U21688 (N_21688,N_18566,N_18845);
and U21689 (N_21689,N_19667,N_18548);
or U21690 (N_21690,N_19647,N_17880);
xor U21691 (N_21691,N_18582,N_18377);
nor U21692 (N_21692,N_17894,N_17579);
nand U21693 (N_21693,N_19694,N_19718);
xnor U21694 (N_21694,N_19720,N_18106);
or U21695 (N_21695,N_17671,N_19910);
nand U21696 (N_21696,N_18720,N_18244);
and U21697 (N_21697,N_18175,N_19701);
nand U21698 (N_21698,N_19982,N_19214);
and U21699 (N_21699,N_19433,N_19043);
or U21700 (N_21700,N_19333,N_18257);
nand U21701 (N_21701,N_18693,N_19077);
or U21702 (N_21702,N_18166,N_18136);
and U21703 (N_21703,N_18013,N_19594);
or U21704 (N_21704,N_19236,N_18048);
or U21705 (N_21705,N_18351,N_17954);
nor U21706 (N_21706,N_18995,N_19922);
xor U21707 (N_21707,N_19106,N_18872);
nor U21708 (N_21708,N_18366,N_18805);
and U21709 (N_21709,N_17935,N_18191);
xor U21710 (N_21710,N_18906,N_18568);
and U21711 (N_21711,N_18389,N_19525);
nor U21712 (N_21712,N_17704,N_17619);
or U21713 (N_21713,N_17687,N_19518);
xnor U21714 (N_21714,N_19166,N_19049);
or U21715 (N_21715,N_17620,N_19014);
xnor U21716 (N_21716,N_19606,N_18163);
nand U21717 (N_21717,N_18252,N_18173);
or U21718 (N_21718,N_18407,N_18765);
xnor U21719 (N_21719,N_19528,N_19139);
nand U21720 (N_21720,N_18071,N_19016);
nor U21721 (N_21721,N_17912,N_19946);
and U21722 (N_21722,N_19703,N_18866);
xnor U21723 (N_21723,N_18824,N_19911);
nor U21724 (N_21724,N_18696,N_19863);
nand U21725 (N_21725,N_18967,N_19525);
nand U21726 (N_21726,N_19813,N_18299);
or U21727 (N_21727,N_18486,N_18545);
nand U21728 (N_21728,N_19267,N_17705);
nor U21729 (N_21729,N_17845,N_17738);
or U21730 (N_21730,N_19537,N_18164);
or U21731 (N_21731,N_17559,N_19832);
nand U21732 (N_21732,N_18792,N_18040);
nor U21733 (N_21733,N_18555,N_19975);
xor U21734 (N_21734,N_18112,N_19810);
xor U21735 (N_21735,N_18073,N_17542);
xor U21736 (N_21736,N_19584,N_18455);
and U21737 (N_21737,N_19336,N_17945);
nand U21738 (N_21738,N_18586,N_17995);
nor U21739 (N_21739,N_18772,N_18029);
and U21740 (N_21740,N_17565,N_17558);
and U21741 (N_21741,N_19690,N_17750);
nor U21742 (N_21742,N_17969,N_18012);
nor U21743 (N_21743,N_18047,N_19081);
nor U21744 (N_21744,N_18337,N_19407);
or U21745 (N_21745,N_19651,N_19648);
xor U21746 (N_21746,N_18105,N_19293);
nand U21747 (N_21747,N_18783,N_17716);
or U21748 (N_21748,N_19262,N_17808);
and U21749 (N_21749,N_18128,N_17859);
xor U21750 (N_21750,N_17943,N_18163);
and U21751 (N_21751,N_18060,N_18680);
or U21752 (N_21752,N_18705,N_18229);
nor U21753 (N_21753,N_19173,N_19143);
and U21754 (N_21754,N_19221,N_17888);
xnor U21755 (N_21755,N_19921,N_18400);
and U21756 (N_21756,N_19153,N_17665);
or U21757 (N_21757,N_19608,N_19461);
and U21758 (N_21758,N_17937,N_17931);
and U21759 (N_21759,N_18190,N_18164);
xnor U21760 (N_21760,N_19691,N_19484);
nor U21761 (N_21761,N_17992,N_19649);
nand U21762 (N_21762,N_18163,N_18535);
nand U21763 (N_21763,N_18828,N_19451);
or U21764 (N_21764,N_19375,N_19443);
xnor U21765 (N_21765,N_18689,N_19316);
nand U21766 (N_21766,N_18351,N_19099);
xor U21767 (N_21767,N_19996,N_19755);
nand U21768 (N_21768,N_19909,N_17982);
or U21769 (N_21769,N_19489,N_17585);
nand U21770 (N_21770,N_18057,N_19908);
nand U21771 (N_21771,N_18626,N_18587);
nor U21772 (N_21772,N_19563,N_17950);
nor U21773 (N_21773,N_18881,N_17503);
xnor U21774 (N_21774,N_19214,N_18044);
xnor U21775 (N_21775,N_18091,N_18259);
or U21776 (N_21776,N_19473,N_19595);
xor U21777 (N_21777,N_18658,N_19814);
or U21778 (N_21778,N_17550,N_19930);
or U21779 (N_21779,N_18442,N_19481);
nand U21780 (N_21780,N_19313,N_17916);
nand U21781 (N_21781,N_19286,N_18515);
nand U21782 (N_21782,N_19675,N_17832);
and U21783 (N_21783,N_19713,N_18059);
and U21784 (N_21784,N_18470,N_18935);
and U21785 (N_21785,N_19076,N_18058);
nand U21786 (N_21786,N_17682,N_19937);
xnor U21787 (N_21787,N_17637,N_18972);
nand U21788 (N_21788,N_18581,N_18632);
xor U21789 (N_21789,N_19792,N_19198);
or U21790 (N_21790,N_18714,N_17625);
xnor U21791 (N_21791,N_18965,N_17833);
nor U21792 (N_21792,N_19289,N_19027);
xnor U21793 (N_21793,N_19984,N_18356);
nand U21794 (N_21794,N_19003,N_19573);
xor U21795 (N_21795,N_18818,N_18107);
xor U21796 (N_21796,N_18123,N_19709);
or U21797 (N_21797,N_18962,N_19246);
xor U21798 (N_21798,N_19551,N_18586);
xor U21799 (N_21799,N_17704,N_18530);
or U21800 (N_21800,N_18396,N_18582);
or U21801 (N_21801,N_19585,N_18470);
and U21802 (N_21802,N_19118,N_18705);
or U21803 (N_21803,N_19676,N_18692);
nand U21804 (N_21804,N_19760,N_18214);
and U21805 (N_21805,N_18614,N_18161);
nand U21806 (N_21806,N_17597,N_19786);
or U21807 (N_21807,N_19032,N_18527);
xnor U21808 (N_21808,N_18704,N_18033);
xor U21809 (N_21809,N_17741,N_17897);
xor U21810 (N_21810,N_19793,N_17796);
nand U21811 (N_21811,N_18882,N_19080);
and U21812 (N_21812,N_19859,N_18671);
xor U21813 (N_21813,N_18723,N_18278);
xnor U21814 (N_21814,N_19467,N_18650);
and U21815 (N_21815,N_18598,N_17604);
nor U21816 (N_21816,N_18761,N_19617);
nand U21817 (N_21817,N_18963,N_19629);
or U21818 (N_21818,N_17685,N_18551);
xor U21819 (N_21819,N_19196,N_18483);
and U21820 (N_21820,N_17855,N_17925);
nand U21821 (N_21821,N_18701,N_19402);
or U21822 (N_21822,N_18671,N_17563);
nor U21823 (N_21823,N_17707,N_17717);
or U21824 (N_21824,N_17941,N_18162);
and U21825 (N_21825,N_18319,N_18975);
xnor U21826 (N_21826,N_19893,N_17553);
and U21827 (N_21827,N_18558,N_19142);
or U21828 (N_21828,N_17818,N_17867);
nand U21829 (N_21829,N_18686,N_17939);
nand U21830 (N_21830,N_19989,N_19465);
or U21831 (N_21831,N_18878,N_17939);
and U21832 (N_21832,N_18143,N_18696);
nor U21833 (N_21833,N_18301,N_18857);
nand U21834 (N_21834,N_17740,N_18854);
xor U21835 (N_21835,N_19025,N_19838);
nand U21836 (N_21836,N_19929,N_19850);
and U21837 (N_21837,N_18402,N_19477);
nor U21838 (N_21838,N_19368,N_17652);
or U21839 (N_21839,N_18699,N_18291);
and U21840 (N_21840,N_19135,N_17630);
xnor U21841 (N_21841,N_18642,N_17672);
nand U21842 (N_21842,N_18805,N_19907);
nand U21843 (N_21843,N_19066,N_17699);
nor U21844 (N_21844,N_18308,N_19212);
or U21845 (N_21845,N_18495,N_17677);
nand U21846 (N_21846,N_19153,N_17535);
nand U21847 (N_21847,N_18558,N_19381);
nor U21848 (N_21848,N_18958,N_19453);
and U21849 (N_21849,N_17639,N_19005);
and U21850 (N_21850,N_19155,N_18394);
nor U21851 (N_21851,N_19288,N_18101);
and U21852 (N_21852,N_18657,N_19051);
and U21853 (N_21853,N_18896,N_18735);
nand U21854 (N_21854,N_18821,N_18532);
and U21855 (N_21855,N_18802,N_18225);
xor U21856 (N_21856,N_18361,N_18566);
nand U21857 (N_21857,N_19546,N_19188);
and U21858 (N_21858,N_18462,N_19422);
or U21859 (N_21859,N_18850,N_17513);
or U21860 (N_21860,N_18174,N_19134);
nor U21861 (N_21861,N_17927,N_18234);
nand U21862 (N_21862,N_18762,N_18116);
and U21863 (N_21863,N_19699,N_19914);
nor U21864 (N_21864,N_18703,N_17967);
nor U21865 (N_21865,N_18029,N_19921);
xnor U21866 (N_21866,N_19403,N_18139);
xor U21867 (N_21867,N_19769,N_18185);
and U21868 (N_21868,N_19507,N_18788);
xor U21869 (N_21869,N_19416,N_18972);
nor U21870 (N_21870,N_18929,N_19358);
xnor U21871 (N_21871,N_19209,N_19442);
xor U21872 (N_21872,N_19598,N_17773);
and U21873 (N_21873,N_19345,N_17537);
nor U21874 (N_21874,N_18449,N_18202);
and U21875 (N_21875,N_18753,N_17685);
or U21876 (N_21876,N_19698,N_19907);
xor U21877 (N_21877,N_17665,N_18469);
xor U21878 (N_21878,N_19793,N_18534);
nand U21879 (N_21879,N_18248,N_18206);
nand U21880 (N_21880,N_19355,N_19691);
or U21881 (N_21881,N_17990,N_18666);
or U21882 (N_21882,N_18466,N_19778);
and U21883 (N_21883,N_18715,N_17705);
and U21884 (N_21884,N_18672,N_17661);
and U21885 (N_21885,N_17992,N_19416);
nor U21886 (N_21886,N_18452,N_19413);
or U21887 (N_21887,N_18539,N_19962);
or U21888 (N_21888,N_19010,N_18303);
xnor U21889 (N_21889,N_18525,N_17552);
or U21890 (N_21890,N_17840,N_18698);
or U21891 (N_21891,N_19662,N_18684);
or U21892 (N_21892,N_18030,N_18104);
nand U21893 (N_21893,N_18347,N_19443);
nand U21894 (N_21894,N_18243,N_17713);
or U21895 (N_21895,N_19505,N_19605);
xnor U21896 (N_21896,N_19858,N_17668);
and U21897 (N_21897,N_18883,N_18967);
nand U21898 (N_21898,N_19781,N_19044);
xnor U21899 (N_21899,N_18024,N_19340);
and U21900 (N_21900,N_18689,N_18554);
nor U21901 (N_21901,N_18657,N_19751);
nand U21902 (N_21902,N_19923,N_18497);
or U21903 (N_21903,N_17671,N_19274);
and U21904 (N_21904,N_18133,N_18729);
nor U21905 (N_21905,N_19255,N_19132);
and U21906 (N_21906,N_18330,N_18613);
nand U21907 (N_21907,N_18321,N_18377);
or U21908 (N_21908,N_18313,N_18876);
or U21909 (N_21909,N_18336,N_19135);
and U21910 (N_21910,N_17728,N_17636);
xor U21911 (N_21911,N_19126,N_19330);
nor U21912 (N_21912,N_18645,N_18543);
nand U21913 (N_21913,N_18074,N_18000);
nor U21914 (N_21914,N_17839,N_18512);
nand U21915 (N_21915,N_18604,N_19763);
nand U21916 (N_21916,N_19852,N_19962);
or U21917 (N_21917,N_18318,N_19433);
nor U21918 (N_21918,N_19833,N_19215);
nand U21919 (N_21919,N_17677,N_19011);
nor U21920 (N_21920,N_19155,N_18174);
nor U21921 (N_21921,N_18729,N_17960);
xnor U21922 (N_21922,N_18416,N_19392);
or U21923 (N_21923,N_18765,N_19054);
xor U21924 (N_21924,N_19738,N_18726);
and U21925 (N_21925,N_19863,N_18990);
or U21926 (N_21926,N_18315,N_18412);
nand U21927 (N_21927,N_17698,N_19538);
nor U21928 (N_21928,N_19703,N_18001);
and U21929 (N_21929,N_17554,N_18145);
and U21930 (N_21930,N_17766,N_19886);
xor U21931 (N_21931,N_19837,N_18793);
nor U21932 (N_21932,N_17997,N_18924);
xor U21933 (N_21933,N_18231,N_19422);
nor U21934 (N_21934,N_19156,N_18727);
nor U21935 (N_21935,N_19580,N_17838);
nor U21936 (N_21936,N_19640,N_19660);
and U21937 (N_21937,N_19282,N_18075);
nor U21938 (N_21938,N_19687,N_18445);
or U21939 (N_21939,N_17659,N_19704);
nor U21940 (N_21940,N_19757,N_17508);
nor U21941 (N_21941,N_18541,N_19736);
xor U21942 (N_21942,N_18702,N_18899);
and U21943 (N_21943,N_19744,N_18503);
or U21944 (N_21944,N_19511,N_18713);
xor U21945 (N_21945,N_17612,N_19964);
xor U21946 (N_21946,N_19050,N_18005);
nor U21947 (N_21947,N_19025,N_18962);
nand U21948 (N_21948,N_17795,N_18780);
xnor U21949 (N_21949,N_18470,N_17664);
nand U21950 (N_21950,N_18385,N_17901);
nor U21951 (N_21951,N_18519,N_17836);
and U21952 (N_21952,N_19851,N_18544);
nor U21953 (N_21953,N_19787,N_19333);
xor U21954 (N_21954,N_18239,N_18928);
or U21955 (N_21955,N_19968,N_17776);
and U21956 (N_21956,N_19850,N_19474);
nor U21957 (N_21957,N_19232,N_19146);
nand U21958 (N_21958,N_18388,N_18573);
and U21959 (N_21959,N_19047,N_18510);
or U21960 (N_21960,N_18613,N_18995);
or U21961 (N_21961,N_18580,N_19350);
and U21962 (N_21962,N_18398,N_19359);
and U21963 (N_21963,N_17502,N_18753);
or U21964 (N_21964,N_17627,N_19802);
nand U21965 (N_21965,N_19199,N_19419);
nor U21966 (N_21966,N_17990,N_18820);
or U21967 (N_21967,N_19775,N_19115);
or U21968 (N_21968,N_19636,N_18591);
nand U21969 (N_21969,N_18409,N_18130);
nand U21970 (N_21970,N_19896,N_19615);
nor U21971 (N_21971,N_19452,N_19468);
nand U21972 (N_21972,N_19658,N_19828);
or U21973 (N_21973,N_18478,N_18247);
nor U21974 (N_21974,N_19372,N_18719);
and U21975 (N_21975,N_18691,N_18877);
or U21976 (N_21976,N_19408,N_19089);
and U21977 (N_21977,N_18953,N_17547);
or U21978 (N_21978,N_18189,N_19755);
and U21979 (N_21979,N_17514,N_19782);
or U21980 (N_21980,N_19515,N_19110);
or U21981 (N_21981,N_17798,N_19402);
nor U21982 (N_21982,N_18376,N_19884);
or U21983 (N_21983,N_18854,N_19849);
nand U21984 (N_21984,N_19984,N_17588);
nand U21985 (N_21985,N_18504,N_17783);
xnor U21986 (N_21986,N_17762,N_19634);
or U21987 (N_21987,N_19029,N_17611);
or U21988 (N_21988,N_19528,N_17748);
nand U21989 (N_21989,N_18154,N_19447);
nand U21990 (N_21990,N_17763,N_19013);
and U21991 (N_21991,N_17685,N_18881);
xor U21992 (N_21992,N_17848,N_19620);
and U21993 (N_21993,N_19605,N_19329);
xnor U21994 (N_21994,N_19574,N_18395);
or U21995 (N_21995,N_18052,N_19942);
nand U21996 (N_21996,N_19155,N_17798);
or U21997 (N_21997,N_19196,N_19233);
nor U21998 (N_21998,N_17525,N_17564);
nand U21999 (N_21999,N_17672,N_17608);
or U22000 (N_22000,N_19635,N_19019);
or U22001 (N_22001,N_18102,N_19137);
and U22002 (N_22002,N_19847,N_18699);
xor U22003 (N_22003,N_19418,N_19149);
and U22004 (N_22004,N_19606,N_17848);
and U22005 (N_22005,N_19157,N_19396);
and U22006 (N_22006,N_17628,N_19845);
or U22007 (N_22007,N_18291,N_17676);
nor U22008 (N_22008,N_19642,N_19688);
nand U22009 (N_22009,N_18626,N_19779);
or U22010 (N_22010,N_18520,N_18658);
and U22011 (N_22011,N_19484,N_19357);
and U22012 (N_22012,N_19649,N_19591);
nand U22013 (N_22013,N_19098,N_18154);
xor U22014 (N_22014,N_19485,N_18832);
nand U22015 (N_22015,N_18875,N_18747);
or U22016 (N_22016,N_18194,N_18247);
nor U22017 (N_22017,N_19887,N_19345);
or U22018 (N_22018,N_17818,N_19054);
xor U22019 (N_22019,N_18232,N_17607);
nor U22020 (N_22020,N_19062,N_17603);
nand U22021 (N_22021,N_17817,N_18550);
xnor U22022 (N_22022,N_19732,N_18134);
nor U22023 (N_22023,N_17829,N_19894);
nor U22024 (N_22024,N_19219,N_19821);
and U22025 (N_22025,N_17605,N_18891);
or U22026 (N_22026,N_19907,N_19864);
or U22027 (N_22027,N_18003,N_18576);
and U22028 (N_22028,N_19577,N_17726);
nor U22029 (N_22029,N_18809,N_17865);
or U22030 (N_22030,N_19498,N_19207);
and U22031 (N_22031,N_17916,N_18026);
xor U22032 (N_22032,N_19223,N_17670);
nor U22033 (N_22033,N_17815,N_18149);
nand U22034 (N_22034,N_18685,N_18106);
nor U22035 (N_22035,N_19290,N_19588);
nor U22036 (N_22036,N_17984,N_18037);
or U22037 (N_22037,N_19922,N_19556);
xor U22038 (N_22038,N_19173,N_18887);
nand U22039 (N_22039,N_18828,N_19377);
or U22040 (N_22040,N_18870,N_19646);
or U22041 (N_22041,N_17862,N_19943);
nor U22042 (N_22042,N_18680,N_18761);
xnor U22043 (N_22043,N_17619,N_18330);
or U22044 (N_22044,N_19496,N_19077);
and U22045 (N_22045,N_19878,N_19877);
xor U22046 (N_22046,N_17696,N_19289);
nor U22047 (N_22047,N_19439,N_18814);
nand U22048 (N_22048,N_19454,N_17597);
and U22049 (N_22049,N_17514,N_19623);
and U22050 (N_22050,N_19240,N_17510);
or U22051 (N_22051,N_17974,N_19211);
or U22052 (N_22052,N_19923,N_17738);
nor U22053 (N_22053,N_19663,N_19022);
and U22054 (N_22054,N_19592,N_18081);
or U22055 (N_22055,N_19955,N_18856);
nor U22056 (N_22056,N_18396,N_17747);
and U22057 (N_22057,N_18965,N_17800);
and U22058 (N_22058,N_17775,N_18643);
and U22059 (N_22059,N_18112,N_18885);
or U22060 (N_22060,N_18614,N_19895);
and U22061 (N_22061,N_17679,N_19641);
or U22062 (N_22062,N_18524,N_18227);
and U22063 (N_22063,N_19562,N_17980);
or U22064 (N_22064,N_19810,N_19411);
and U22065 (N_22065,N_18517,N_17734);
nor U22066 (N_22066,N_19236,N_17739);
xor U22067 (N_22067,N_17925,N_18697);
xor U22068 (N_22068,N_18227,N_18974);
nor U22069 (N_22069,N_18018,N_19608);
or U22070 (N_22070,N_19711,N_19610);
or U22071 (N_22071,N_18358,N_17592);
and U22072 (N_22072,N_19744,N_18191);
and U22073 (N_22073,N_19721,N_17716);
and U22074 (N_22074,N_18097,N_17835);
or U22075 (N_22075,N_18011,N_19610);
nor U22076 (N_22076,N_19055,N_19640);
and U22077 (N_22077,N_19311,N_18680);
xnor U22078 (N_22078,N_19645,N_19821);
xor U22079 (N_22079,N_18722,N_18048);
nor U22080 (N_22080,N_18420,N_19480);
xor U22081 (N_22081,N_17900,N_19898);
nand U22082 (N_22082,N_17991,N_19837);
and U22083 (N_22083,N_19671,N_19348);
nand U22084 (N_22084,N_19479,N_18473);
or U22085 (N_22085,N_18247,N_18079);
nor U22086 (N_22086,N_18568,N_19211);
xnor U22087 (N_22087,N_19220,N_19153);
nor U22088 (N_22088,N_17592,N_18427);
nand U22089 (N_22089,N_19681,N_18251);
xnor U22090 (N_22090,N_19648,N_18325);
nor U22091 (N_22091,N_18284,N_19824);
xor U22092 (N_22092,N_17939,N_17551);
or U22093 (N_22093,N_18413,N_17745);
or U22094 (N_22094,N_19276,N_18814);
xor U22095 (N_22095,N_19608,N_18185);
or U22096 (N_22096,N_18933,N_17967);
and U22097 (N_22097,N_18168,N_19521);
xor U22098 (N_22098,N_17640,N_18808);
or U22099 (N_22099,N_18622,N_19796);
nand U22100 (N_22100,N_18978,N_19148);
nor U22101 (N_22101,N_18149,N_18374);
or U22102 (N_22102,N_17685,N_19058);
or U22103 (N_22103,N_19076,N_17896);
nand U22104 (N_22104,N_18750,N_17670);
nor U22105 (N_22105,N_19204,N_18734);
nor U22106 (N_22106,N_19920,N_19300);
nand U22107 (N_22107,N_19240,N_19675);
and U22108 (N_22108,N_17911,N_17711);
xor U22109 (N_22109,N_18326,N_19131);
nor U22110 (N_22110,N_17823,N_19896);
xnor U22111 (N_22111,N_17629,N_17936);
nand U22112 (N_22112,N_17595,N_19867);
xor U22113 (N_22113,N_18529,N_18400);
xor U22114 (N_22114,N_18819,N_19591);
nand U22115 (N_22115,N_18784,N_18922);
xnor U22116 (N_22116,N_19102,N_19469);
or U22117 (N_22117,N_17561,N_19506);
nand U22118 (N_22118,N_18229,N_18970);
and U22119 (N_22119,N_17886,N_19875);
xnor U22120 (N_22120,N_18572,N_19591);
and U22121 (N_22121,N_17943,N_17947);
nor U22122 (N_22122,N_19787,N_17604);
and U22123 (N_22123,N_18594,N_19296);
nand U22124 (N_22124,N_17794,N_18026);
and U22125 (N_22125,N_19256,N_18392);
nor U22126 (N_22126,N_19233,N_18111);
nand U22127 (N_22127,N_19994,N_18407);
nor U22128 (N_22128,N_18043,N_18369);
nor U22129 (N_22129,N_19212,N_18352);
xor U22130 (N_22130,N_17730,N_17987);
xor U22131 (N_22131,N_19812,N_19766);
and U22132 (N_22132,N_17622,N_18796);
xor U22133 (N_22133,N_19330,N_18716);
nand U22134 (N_22134,N_18157,N_19057);
nor U22135 (N_22135,N_19802,N_18658);
nand U22136 (N_22136,N_19333,N_19703);
and U22137 (N_22137,N_19028,N_19793);
nand U22138 (N_22138,N_19918,N_19393);
nor U22139 (N_22139,N_18241,N_17674);
or U22140 (N_22140,N_17675,N_19646);
nand U22141 (N_22141,N_19956,N_19973);
nor U22142 (N_22142,N_18483,N_17990);
xor U22143 (N_22143,N_19736,N_19142);
xor U22144 (N_22144,N_19391,N_18044);
xnor U22145 (N_22145,N_17958,N_18459);
xnor U22146 (N_22146,N_19221,N_19097);
and U22147 (N_22147,N_18082,N_17525);
nand U22148 (N_22148,N_18302,N_18639);
or U22149 (N_22149,N_18936,N_18257);
and U22150 (N_22150,N_18128,N_18601);
nand U22151 (N_22151,N_18610,N_18593);
or U22152 (N_22152,N_18723,N_17761);
or U22153 (N_22153,N_18873,N_19987);
and U22154 (N_22154,N_18242,N_18434);
xor U22155 (N_22155,N_18980,N_18463);
and U22156 (N_22156,N_19496,N_17615);
nor U22157 (N_22157,N_19360,N_18862);
nand U22158 (N_22158,N_18276,N_18810);
or U22159 (N_22159,N_18918,N_17888);
or U22160 (N_22160,N_18268,N_18487);
nor U22161 (N_22161,N_19569,N_19696);
nand U22162 (N_22162,N_19699,N_17552);
nand U22163 (N_22163,N_18183,N_17785);
and U22164 (N_22164,N_17552,N_18249);
and U22165 (N_22165,N_17716,N_18430);
nor U22166 (N_22166,N_19324,N_18103);
xnor U22167 (N_22167,N_18786,N_17810);
or U22168 (N_22168,N_18939,N_18293);
xnor U22169 (N_22169,N_19530,N_17699);
nand U22170 (N_22170,N_19856,N_19273);
and U22171 (N_22171,N_17806,N_18499);
xnor U22172 (N_22172,N_17921,N_19935);
and U22173 (N_22173,N_18356,N_18574);
or U22174 (N_22174,N_18340,N_18405);
and U22175 (N_22175,N_17655,N_18384);
xnor U22176 (N_22176,N_18380,N_18353);
nor U22177 (N_22177,N_18506,N_19979);
or U22178 (N_22178,N_18964,N_18429);
or U22179 (N_22179,N_19106,N_17933);
nor U22180 (N_22180,N_17515,N_18630);
xnor U22181 (N_22181,N_18647,N_18661);
xor U22182 (N_22182,N_18907,N_18309);
nor U22183 (N_22183,N_19185,N_18100);
or U22184 (N_22184,N_18549,N_18532);
nor U22185 (N_22185,N_18614,N_19098);
or U22186 (N_22186,N_19066,N_17547);
nand U22187 (N_22187,N_18264,N_19420);
nand U22188 (N_22188,N_17596,N_18723);
and U22189 (N_22189,N_18992,N_18072);
and U22190 (N_22190,N_17889,N_18001);
and U22191 (N_22191,N_19378,N_18429);
nor U22192 (N_22192,N_17743,N_17744);
xor U22193 (N_22193,N_18115,N_18015);
and U22194 (N_22194,N_18627,N_17681);
xor U22195 (N_22195,N_17685,N_18135);
nor U22196 (N_22196,N_19999,N_19934);
or U22197 (N_22197,N_18633,N_19754);
or U22198 (N_22198,N_17844,N_19921);
xor U22199 (N_22199,N_18067,N_17625);
nor U22200 (N_22200,N_17599,N_18290);
and U22201 (N_22201,N_18328,N_19575);
or U22202 (N_22202,N_19175,N_17946);
or U22203 (N_22203,N_18176,N_19262);
and U22204 (N_22204,N_18700,N_17527);
and U22205 (N_22205,N_18058,N_17641);
nor U22206 (N_22206,N_18282,N_18483);
nor U22207 (N_22207,N_19939,N_17840);
nor U22208 (N_22208,N_18522,N_19256);
and U22209 (N_22209,N_19780,N_19754);
nand U22210 (N_22210,N_19627,N_19940);
nor U22211 (N_22211,N_19531,N_19095);
nor U22212 (N_22212,N_19530,N_19993);
and U22213 (N_22213,N_18968,N_18266);
nor U22214 (N_22214,N_19978,N_18961);
and U22215 (N_22215,N_18195,N_18745);
or U22216 (N_22216,N_17799,N_18585);
nor U22217 (N_22217,N_17646,N_19722);
or U22218 (N_22218,N_19700,N_19014);
and U22219 (N_22219,N_18728,N_19717);
and U22220 (N_22220,N_19011,N_18639);
nor U22221 (N_22221,N_19342,N_18538);
nand U22222 (N_22222,N_18259,N_19338);
nor U22223 (N_22223,N_18685,N_18296);
nand U22224 (N_22224,N_19146,N_19538);
and U22225 (N_22225,N_19176,N_19849);
nand U22226 (N_22226,N_19127,N_19121);
nor U22227 (N_22227,N_18066,N_19348);
or U22228 (N_22228,N_17616,N_18081);
xnor U22229 (N_22229,N_17765,N_18984);
and U22230 (N_22230,N_19519,N_18078);
nor U22231 (N_22231,N_18636,N_17586);
nand U22232 (N_22232,N_18972,N_18420);
nor U22233 (N_22233,N_18422,N_18825);
and U22234 (N_22234,N_19850,N_18524);
xor U22235 (N_22235,N_17569,N_19502);
nand U22236 (N_22236,N_17865,N_18018);
and U22237 (N_22237,N_18203,N_19805);
xor U22238 (N_22238,N_18089,N_18020);
nor U22239 (N_22239,N_18742,N_18887);
and U22240 (N_22240,N_19010,N_19346);
nand U22241 (N_22241,N_18687,N_18099);
and U22242 (N_22242,N_19087,N_18443);
nand U22243 (N_22243,N_18934,N_19054);
nor U22244 (N_22244,N_18865,N_18545);
or U22245 (N_22245,N_18197,N_19776);
or U22246 (N_22246,N_19965,N_19790);
nand U22247 (N_22247,N_18518,N_17768);
or U22248 (N_22248,N_19868,N_18918);
xnor U22249 (N_22249,N_19317,N_19470);
or U22250 (N_22250,N_19501,N_19242);
nor U22251 (N_22251,N_19081,N_18194);
nor U22252 (N_22252,N_17553,N_17651);
and U22253 (N_22253,N_17715,N_19239);
nand U22254 (N_22254,N_19826,N_18852);
nor U22255 (N_22255,N_19654,N_19794);
xnor U22256 (N_22256,N_19876,N_19199);
or U22257 (N_22257,N_19993,N_18157);
xor U22258 (N_22258,N_19202,N_18084);
nor U22259 (N_22259,N_17767,N_19006);
and U22260 (N_22260,N_18016,N_19828);
nor U22261 (N_22261,N_18513,N_18365);
and U22262 (N_22262,N_18629,N_19506);
nand U22263 (N_22263,N_19796,N_17988);
nand U22264 (N_22264,N_18099,N_19154);
xnor U22265 (N_22265,N_18563,N_18099);
and U22266 (N_22266,N_19734,N_18701);
xnor U22267 (N_22267,N_18205,N_18084);
nand U22268 (N_22268,N_17703,N_19748);
nand U22269 (N_22269,N_19818,N_19291);
or U22270 (N_22270,N_19285,N_18993);
or U22271 (N_22271,N_18094,N_18315);
and U22272 (N_22272,N_18551,N_19830);
and U22273 (N_22273,N_17617,N_19468);
or U22274 (N_22274,N_19435,N_19847);
and U22275 (N_22275,N_18254,N_18654);
and U22276 (N_22276,N_18752,N_17680);
and U22277 (N_22277,N_18950,N_18915);
or U22278 (N_22278,N_17702,N_19465);
nor U22279 (N_22279,N_19154,N_19999);
nor U22280 (N_22280,N_18766,N_17651);
nor U22281 (N_22281,N_17666,N_19944);
or U22282 (N_22282,N_19720,N_19918);
and U22283 (N_22283,N_19174,N_17923);
and U22284 (N_22284,N_18848,N_18267);
and U22285 (N_22285,N_19311,N_19083);
or U22286 (N_22286,N_18697,N_18270);
xnor U22287 (N_22287,N_18069,N_18620);
nand U22288 (N_22288,N_17590,N_18767);
and U22289 (N_22289,N_17971,N_18146);
and U22290 (N_22290,N_19500,N_18975);
and U22291 (N_22291,N_17572,N_18840);
or U22292 (N_22292,N_18572,N_18544);
or U22293 (N_22293,N_19033,N_19192);
nor U22294 (N_22294,N_18323,N_17568);
and U22295 (N_22295,N_18051,N_19488);
nand U22296 (N_22296,N_18521,N_17680);
nor U22297 (N_22297,N_17666,N_19151);
xor U22298 (N_22298,N_18332,N_18829);
or U22299 (N_22299,N_19291,N_19508);
or U22300 (N_22300,N_17731,N_19567);
nor U22301 (N_22301,N_19512,N_19228);
or U22302 (N_22302,N_18295,N_18355);
and U22303 (N_22303,N_18592,N_18580);
nor U22304 (N_22304,N_19496,N_18155);
nand U22305 (N_22305,N_18995,N_18987);
xnor U22306 (N_22306,N_19200,N_19965);
nor U22307 (N_22307,N_19123,N_18150);
nand U22308 (N_22308,N_18923,N_19902);
or U22309 (N_22309,N_19632,N_18708);
or U22310 (N_22310,N_19286,N_18275);
or U22311 (N_22311,N_18770,N_18089);
nor U22312 (N_22312,N_19257,N_19260);
xor U22313 (N_22313,N_18617,N_17983);
xor U22314 (N_22314,N_17607,N_19018);
nand U22315 (N_22315,N_18188,N_18555);
or U22316 (N_22316,N_19159,N_19158);
nor U22317 (N_22317,N_18532,N_19988);
xnor U22318 (N_22318,N_19928,N_18885);
nand U22319 (N_22319,N_17652,N_18906);
and U22320 (N_22320,N_19402,N_18441);
nor U22321 (N_22321,N_18810,N_19290);
and U22322 (N_22322,N_17803,N_19461);
nor U22323 (N_22323,N_18233,N_19524);
nor U22324 (N_22324,N_19636,N_18961);
nand U22325 (N_22325,N_17898,N_18456);
and U22326 (N_22326,N_17632,N_17906);
or U22327 (N_22327,N_19104,N_18252);
nand U22328 (N_22328,N_17655,N_18472);
or U22329 (N_22329,N_19100,N_17561);
or U22330 (N_22330,N_18720,N_17783);
and U22331 (N_22331,N_19172,N_18522);
nor U22332 (N_22332,N_19640,N_18804);
or U22333 (N_22333,N_18894,N_19721);
xor U22334 (N_22334,N_18379,N_17660);
nor U22335 (N_22335,N_19183,N_18657);
nand U22336 (N_22336,N_17917,N_19637);
nand U22337 (N_22337,N_18951,N_19485);
xor U22338 (N_22338,N_17936,N_19069);
nand U22339 (N_22339,N_19303,N_18093);
nand U22340 (N_22340,N_18319,N_17636);
and U22341 (N_22341,N_19673,N_18245);
nor U22342 (N_22342,N_19860,N_18415);
and U22343 (N_22343,N_19208,N_19689);
xnor U22344 (N_22344,N_19893,N_18247);
nor U22345 (N_22345,N_18826,N_19269);
and U22346 (N_22346,N_18268,N_19892);
nand U22347 (N_22347,N_18474,N_18324);
xnor U22348 (N_22348,N_19385,N_18380);
xnor U22349 (N_22349,N_19857,N_19877);
xor U22350 (N_22350,N_18250,N_17556);
nand U22351 (N_22351,N_18782,N_18304);
nor U22352 (N_22352,N_19178,N_19489);
or U22353 (N_22353,N_18000,N_18804);
nor U22354 (N_22354,N_19781,N_18682);
and U22355 (N_22355,N_18521,N_18967);
xor U22356 (N_22356,N_17978,N_19132);
and U22357 (N_22357,N_19754,N_17693);
nand U22358 (N_22358,N_17839,N_19215);
nand U22359 (N_22359,N_19550,N_17947);
or U22360 (N_22360,N_19706,N_19933);
or U22361 (N_22361,N_17787,N_17769);
nor U22362 (N_22362,N_19298,N_18586);
or U22363 (N_22363,N_18237,N_18178);
nand U22364 (N_22364,N_18366,N_17532);
or U22365 (N_22365,N_18607,N_18466);
and U22366 (N_22366,N_19961,N_18271);
nand U22367 (N_22367,N_19474,N_19319);
or U22368 (N_22368,N_19585,N_19239);
and U22369 (N_22369,N_18878,N_18947);
nor U22370 (N_22370,N_19985,N_19995);
and U22371 (N_22371,N_17844,N_18515);
or U22372 (N_22372,N_18055,N_18474);
xnor U22373 (N_22373,N_18521,N_19783);
or U22374 (N_22374,N_18539,N_18514);
and U22375 (N_22375,N_18371,N_19197);
and U22376 (N_22376,N_18001,N_19104);
nor U22377 (N_22377,N_19075,N_19067);
and U22378 (N_22378,N_19147,N_19099);
nand U22379 (N_22379,N_19109,N_18391);
nand U22380 (N_22380,N_18440,N_17571);
xnor U22381 (N_22381,N_19134,N_18866);
and U22382 (N_22382,N_18696,N_17517);
or U22383 (N_22383,N_17809,N_17558);
nor U22384 (N_22384,N_17927,N_17978);
or U22385 (N_22385,N_19367,N_17591);
and U22386 (N_22386,N_18952,N_19054);
nand U22387 (N_22387,N_18743,N_17800);
xnor U22388 (N_22388,N_17804,N_17657);
nor U22389 (N_22389,N_19350,N_19524);
and U22390 (N_22390,N_19072,N_18370);
xor U22391 (N_22391,N_18550,N_19797);
nor U22392 (N_22392,N_18593,N_18731);
and U22393 (N_22393,N_18234,N_19447);
or U22394 (N_22394,N_17964,N_19207);
nand U22395 (N_22395,N_19439,N_19929);
xnor U22396 (N_22396,N_19766,N_18797);
nor U22397 (N_22397,N_17778,N_18506);
xor U22398 (N_22398,N_18637,N_17667);
nor U22399 (N_22399,N_19788,N_18438);
or U22400 (N_22400,N_19038,N_18795);
and U22401 (N_22401,N_19995,N_19703);
xor U22402 (N_22402,N_19912,N_17716);
xor U22403 (N_22403,N_19789,N_19317);
nor U22404 (N_22404,N_17909,N_19729);
nor U22405 (N_22405,N_17571,N_19630);
and U22406 (N_22406,N_19771,N_18851);
xnor U22407 (N_22407,N_17558,N_17507);
nor U22408 (N_22408,N_17531,N_19249);
xnor U22409 (N_22409,N_18718,N_17997);
nand U22410 (N_22410,N_19651,N_17904);
nor U22411 (N_22411,N_19324,N_19155);
xnor U22412 (N_22412,N_18649,N_19139);
nand U22413 (N_22413,N_18773,N_18716);
or U22414 (N_22414,N_19569,N_18323);
xnor U22415 (N_22415,N_19470,N_19882);
nand U22416 (N_22416,N_17632,N_17766);
or U22417 (N_22417,N_18268,N_17576);
nor U22418 (N_22418,N_19418,N_19844);
xnor U22419 (N_22419,N_19479,N_18561);
nor U22420 (N_22420,N_19342,N_19065);
nand U22421 (N_22421,N_19721,N_18160);
nand U22422 (N_22422,N_18607,N_18287);
nand U22423 (N_22423,N_19758,N_17742);
or U22424 (N_22424,N_18764,N_18226);
or U22425 (N_22425,N_17615,N_18189);
nand U22426 (N_22426,N_17640,N_18682);
and U22427 (N_22427,N_19160,N_17910);
and U22428 (N_22428,N_19176,N_19289);
nand U22429 (N_22429,N_19696,N_17573);
and U22430 (N_22430,N_19430,N_19132);
nor U22431 (N_22431,N_18747,N_19223);
nor U22432 (N_22432,N_18450,N_19510);
xnor U22433 (N_22433,N_18714,N_19808);
nor U22434 (N_22434,N_19209,N_17905);
or U22435 (N_22435,N_17998,N_18946);
nand U22436 (N_22436,N_19054,N_19585);
and U22437 (N_22437,N_17603,N_18529);
xor U22438 (N_22438,N_19446,N_19528);
nand U22439 (N_22439,N_18648,N_19829);
and U22440 (N_22440,N_19018,N_18002);
or U22441 (N_22441,N_17745,N_18303);
nand U22442 (N_22442,N_19650,N_18210);
nor U22443 (N_22443,N_19131,N_17774);
and U22444 (N_22444,N_18911,N_19989);
xor U22445 (N_22445,N_17615,N_19354);
and U22446 (N_22446,N_17567,N_18972);
xor U22447 (N_22447,N_19398,N_17945);
or U22448 (N_22448,N_18652,N_18883);
or U22449 (N_22449,N_17927,N_19753);
nand U22450 (N_22450,N_18617,N_17825);
nor U22451 (N_22451,N_19618,N_19205);
nand U22452 (N_22452,N_18774,N_17658);
and U22453 (N_22453,N_18230,N_17901);
xor U22454 (N_22454,N_18406,N_17576);
and U22455 (N_22455,N_19358,N_19416);
nor U22456 (N_22456,N_18292,N_19293);
or U22457 (N_22457,N_17924,N_19292);
nand U22458 (N_22458,N_17938,N_18839);
xor U22459 (N_22459,N_18080,N_17845);
nor U22460 (N_22460,N_19544,N_18605);
xor U22461 (N_22461,N_19904,N_19670);
xor U22462 (N_22462,N_19538,N_19014);
nand U22463 (N_22463,N_18244,N_19726);
nor U22464 (N_22464,N_19418,N_18059);
nand U22465 (N_22465,N_18561,N_18020);
nor U22466 (N_22466,N_18371,N_18570);
nand U22467 (N_22467,N_18728,N_19537);
or U22468 (N_22468,N_18841,N_17527);
xnor U22469 (N_22469,N_18570,N_18906);
nand U22470 (N_22470,N_17768,N_18838);
or U22471 (N_22471,N_19606,N_18801);
xor U22472 (N_22472,N_19376,N_18585);
and U22473 (N_22473,N_17766,N_17579);
nand U22474 (N_22474,N_19410,N_18473);
and U22475 (N_22475,N_19812,N_17576);
nand U22476 (N_22476,N_18805,N_18835);
and U22477 (N_22477,N_19157,N_18917);
nor U22478 (N_22478,N_17622,N_17812);
or U22479 (N_22479,N_19892,N_19134);
xor U22480 (N_22480,N_19442,N_18062);
nor U22481 (N_22481,N_17638,N_18534);
nand U22482 (N_22482,N_18915,N_19347);
nor U22483 (N_22483,N_17693,N_18591);
or U22484 (N_22484,N_18211,N_17641);
xnor U22485 (N_22485,N_18111,N_18159);
nor U22486 (N_22486,N_18107,N_19436);
and U22487 (N_22487,N_18573,N_18277);
nand U22488 (N_22488,N_18823,N_19423);
nand U22489 (N_22489,N_17677,N_18268);
or U22490 (N_22490,N_18274,N_19898);
nand U22491 (N_22491,N_19646,N_19877);
and U22492 (N_22492,N_19474,N_18092);
nor U22493 (N_22493,N_18416,N_18968);
nor U22494 (N_22494,N_18512,N_19193);
nand U22495 (N_22495,N_17837,N_19308);
nor U22496 (N_22496,N_19173,N_18738);
xor U22497 (N_22497,N_18431,N_19371);
nor U22498 (N_22498,N_17832,N_18170);
nor U22499 (N_22499,N_18220,N_18708);
xnor U22500 (N_22500,N_20312,N_22150);
xnor U22501 (N_22501,N_20417,N_20812);
nand U22502 (N_22502,N_22048,N_21134);
nand U22503 (N_22503,N_20227,N_21821);
or U22504 (N_22504,N_20068,N_20166);
xor U22505 (N_22505,N_21641,N_22092);
or U22506 (N_22506,N_21802,N_20803);
or U22507 (N_22507,N_21005,N_21506);
xnor U22508 (N_22508,N_20444,N_20741);
nand U22509 (N_22509,N_21168,N_20486);
or U22510 (N_22510,N_21805,N_21563);
or U22511 (N_22511,N_21696,N_21468);
nand U22512 (N_22512,N_20045,N_22071);
nor U22513 (N_22513,N_21717,N_22024);
or U22514 (N_22514,N_21020,N_20944);
or U22515 (N_22515,N_21992,N_21941);
nand U22516 (N_22516,N_21372,N_21116);
or U22517 (N_22517,N_21849,N_20351);
nand U22518 (N_22518,N_20397,N_21816);
nand U22519 (N_22519,N_21107,N_21889);
or U22520 (N_22520,N_21387,N_20214);
nor U22521 (N_22521,N_21776,N_21709);
xor U22522 (N_22522,N_21879,N_20002);
nor U22523 (N_22523,N_21469,N_21220);
xor U22524 (N_22524,N_21826,N_21775);
nor U22525 (N_22525,N_21182,N_21517);
xor U22526 (N_22526,N_20709,N_22323);
nor U22527 (N_22527,N_21571,N_21628);
and U22528 (N_22528,N_21919,N_20061);
and U22529 (N_22529,N_21969,N_21945);
nand U22530 (N_22530,N_20830,N_20906);
xnor U22531 (N_22531,N_21631,N_20152);
nand U22532 (N_22532,N_21984,N_21386);
nor U22533 (N_22533,N_20731,N_22359);
nand U22534 (N_22534,N_20996,N_20590);
xnor U22535 (N_22535,N_20897,N_20368);
and U22536 (N_22536,N_22053,N_21327);
and U22537 (N_22537,N_22171,N_20625);
nor U22538 (N_22538,N_21158,N_20951);
xnor U22539 (N_22539,N_21413,N_21659);
or U22540 (N_22540,N_20828,N_20952);
nand U22541 (N_22541,N_21562,N_20147);
and U22542 (N_22542,N_20220,N_21948);
and U22543 (N_22543,N_21519,N_22486);
xor U22544 (N_22544,N_22131,N_21378);
and U22545 (N_22545,N_20096,N_21216);
and U22546 (N_22546,N_20679,N_21783);
nand U22547 (N_22547,N_21914,N_20860);
or U22548 (N_22548,N_21973,N_21325);
nor U22549 (N_22549,N_22107,N_20307);
nor U22550 (N_22550,N_20501,N_21685);
nand U22551 (N_22551,N_20910,N_20256);
xor U22552 (N_22552,N_22253,N_20885);
or U22553 (N_22553,N_21249,N_21708);
nand U22554 (N_22554,N_20446,N_20587);
xnor U22555 (N_22555,N_21938,N_20248);
or U22556 (N_22556,N_22122,N_21532);
or U22557 (N_22557,N_22305,N_20950);
and U22558 (N_22558,N_20500,N_21366);
nand U22559 (N_22559,N_20413,N_21104);
nand U22560 (N_22560,N_20841,N_20375);
nor U22561 (N_22561,N_20322,N_20280);
and U22562 (N_22562,N_20270,N_22006);
nor U22563 (N_22563,N_20102,N_20879);
and U22564 (N_22564,N_21354,N_22363);
xnor U22565 (N_22565,N_21014,N_20311);
xnor U22566 (N_22566,N_20561,N_21291);
and U22567 (N_22567,N_21585,N_21037);
nor U22568 (N_22568,N_20518,N_20580);
or U22569 (N_22569,N_20053,N_22416);
or U22570 (N_22570,N_21435,N_20161);
nor U22571 (N_22571,N_21731,N_22090);
nor U22572 (N_22572,N_20328,N_20407);
and U22573 (N_22573,N_20752,N_20081);
or U22574 (N_22574,N_21120,N_20491);
or U22575 (N_22575,N_21953,N_22436);
xor U22576 (N_22576,N_21494,N_21219);
xnor U22577 (N_22577,N_22472,N_20034);
xnor U22578 (N_22578,N_21877,N_21210);
and U22579 (N_22579,N_20484,N_20243);
xnor U22580 (N_22580,N_20620,N_22476);
or U22581 (N_22581,N_22298,N_22213);
xor U22582 (N_22582,N_20338,N_21382);
nand U22583 (N_22583,N_21287,N_21432);
or U22584 (N_22584,N_21780,N_21925);
nor U22585 (N_22585,N_22244,N_22342);
nor U22586 (N_22586,N_21977,N_20246);
nand U22587 (N_22587,N_22258,N_20215);
nor U22588 (N_22588,N_20320,N_20678);
or U22589 (N_22589,N_21465,N_21215);
xor U22590 (N_22590,N_22319,N_20048);
nor U22591 (N_22591,N_21292,N_20915);
xor U22592 (N_22592,N_20864,N_20517);
xor U22593 (N_22593,N_20558,N_21208);
or U22594 (N_22594,N_21309,N_21408);
xor U22595 (N_22595,N_21103,N_20472);
or U22596 (N_22596,N_22477,N_22438);
nand U22597 (N_22597,N_21957,N_20768);
nor U22598 (N_22598,N_20403,N_21461);
xor U22599 (N_22599,N_21772,N_22007);
nor U22600 (N_22600,N_20800,N_22205);
or U22601 (N_22601,N_22260,N_21724);
xor U22602 (N_22602,N_20595,N_20569);
xnor U22603 (N_22603,N_22354,N_20749);
and U22604 (N_22604,N_22154,N_20074);
and U22605 (N_22605,N_20681,N_21740);
nand U22606 (N_22606,N_20998,N_21561);
xor U22607 (N_22607,N_21293,N_20576);
or U22608 (N_22608,N_20976,N_22032);
nand U22609 (N_22609,N_21131,N_22325);
or U22610 (N_22610,N_22093,N_22474);
xnor U22611 (N_22611,N_20156,N_20865);
xnor U22612 (N_22612,N_21323,N_20689);
nor U22613 (N_22613,N_21541,N_21706);
xnor U22614 (N_22614,N_21167,N_21034);
nand U22615 (N_22615,N_22182,N_20541);
xnor U22616 (N_22616,N_22062,N_21508);
nand U22617 (N_22617,N_21012,N_20715);
or U22618 (N_22618,N_21620,N_20130);
xnor U22619 (N_22619,N_20783,N_22261);
and U22620 (N_22620,N_22497,N_20792);
nor U22621 (N_22621,N_21023,N_20361);
nand U22622 (N_22622,N_20271,N_20009);
nand U22623 (N_22623,N_21243,N_20474);
or U22624 (N_22624,N_22118,N_20943);
nor U22625 (N_22625,N_21610,N_20939);
nor U22626 (N_22626,N_21252,N_22185);
nor U22627 (N_22627,N_21692,N_20921);
nor U22628 (N_22628,N_21027,N_21225);
and U22629 (N_22629,N_22398,N_20775);
nand U22630 (N_22630,N_20711,N_20259);
or U22631 (N_22631,N_20699,N_20022);
and U22632 (N_22632,N_22215,N_21085);
nand U22633 (N_22633,N_21820,N_21007);
nand U22634 (N_22634,N_21779,N_21736);
or U22635 (N_22635,N_21883,N_21240);
xor U22636 (N_22636,N_20324,N_22119);
nor U22637 (N_22637,N_21575,N_20412);
nand U22638 (N_22638,N_22255,N_21503);
nor U22639 (N_22639,N_20736,N_20958);
or U22640 (N_22640,N_20478,N_20080);
nand U22641 (N_22641,N_21431,N_21700);
nand U22642 (N_22642,N_21411,N_20172);
xor U22643 (N_22643,N_20723,N_22491);
and U22644 (N_22644,N_21666,N_22345);
nor U22645 (N_22645,N_21611,N_21434);
or U22646 (N_22646,N_21398,N_22218);
nand U22647 (N_22647,N_22029,N_20824);
nor U22648 (N_22648,N_21381,N_21365);
nor U22649 (N_22649,N_21766,N_20928);
xnor U22650 (N_22650,N_20925,N_20884);
and U22651 (N_22651,N_21464,N_20268);
and U22652 (N_22652,N_20370,N_21392);
or U22653 (N_22653,N_21466,N_20528);
or U22654 (N_22654,N_20379,N_21202);
nor U22655 (N_22655,N_20532,N_21908);
xor U22656 (N_22656,N_20377,N_20737);
xnor U22657 (N_22657,N_20111,N_21657);
nand U22658 (N_22658,N_20390,N_22113);
and U22659 (N_22659,N_21993,N_21892);
nor U22660 (N_22660,N_21792,N_21499);
and U22661 (N_22661,N_21197,N_20714);
nor U22662 (N_22662,N_22371,N_20041);
nand U22663 (N_22663,N_21830,N_20748);
or U22664 (N_22664,N_22198,N_20940);
and U22665 (N_22665,N_21172,N_21001);
nor U22666 (N_22666,N_20618,N_21545);
or U22667 (N_22667,N_21051,N_21337);
or U22668 (N_22668,N_20738,N_22186);
and U22669 (N_22669,N_21454,N_20447);
or U22670 (N_22670,N_21042,N_20688);
nand U22671 (N_22671,N_21446,N_22480);
xor U22672 (N_22672,N_21145,N_20896);
or U22673 (N_22673,N_21328,N_22036);
xor U22674 (N_22674,N_20055,N_22179);
nor U22675 (N_22675,N_22475,N_20893);
xnor U22676 (N_22676,N_21880,N_20599);
xor U22677 (N_22677,N_21095,N_20471);
and U22678 (N_22678,N_21785,N_20623);
and U22679 (N_22679,N_21974,N_21478);
xor U22680 (N_22680,N_21759,N_21937);
and U22681 (N_22681,N_20926,N_21618);
and U22682 (N_22682,N_20973,N_21595);
nor U22683 (N_22683,N_20203,N_20666);
nor U22684 (N_22684,N_21568,N_21960);
or U22685 (N_22685,N_21841,N_20790);
nor U22686 (N_22686,N_20815,N_20601);
nand U22687 (N_22687,N_20033,N_21244);
and U22688 (N_22688,N_20186,N_20570);
xnor U22689 (N_22689,N_22242,N_21604);
or U22690 (N_22690,N_22214,N_21927);
xnor U22691 (N_22691,N_20133,N_21053);
or U22692 (N_22692,N_21286,N_21749);
nand U22693 (N_22693,N_21601,N_21681);
nor U22694 (N_22694,N_20529,N_22203);
xnor U22695 (N_22695,N_20160,N_20088);
xor U22696 (N_22696,N_21033,N_20350);
nand U22697 (N_22697,N_21306,N_20739);
nor U22698 (N_22698,N_20914,N_21647);
nand U22699 (N_22699,N_21522,N_22227);
nor U22700 (N_22700,N_21317,N_20704);
nand U22701 (N_22701,N_22020,N_22259);
and U22702 (N_22702,N_20924,N_22152);
nor U22703 (N_22703,N_21019,N_21560);
nor U22704 (N_22704,N_22166,N_20682);
nor U22705 (N_22705,N_22392,N_21196);
nand U22706 (N_22706,N_20707,N_21041);
nand U22707 (N_22707,N_20276,N_21092);
and U22708 (N_22708,N_20453,N_20165);
and U22709 (N_22709,N_21718,N_20189);
nor U22710 (N_22710,N_21224,N_21473);
xnor U22711 (N_22711,N_20909,N_20706);
xnor U22712 (N_22712,N_21739,N_22478);
or U22713 (N_22713,N_21111,N_20226);
nand U22714 (N_22714,N_20605,N_20459);
or U22715 (N_22715,N_20753,N_21296);
nand U22716 (N_22716,N_20432,N_21000);
xnor U22717 (N_22717,N_22338,N_20542);
or U22718 (N_22718,N_20365,N_22043);
and U22719 (N_22719,N_21460,N_21728);
and U22720 (N_22720,N_20037,N_20819);
nor U22721 (N_22721,N_21985,N_20005);
nand U22722 (N_22722,N_21227,N_22173);
and U22723 (N_22723,N_22456,N_21295);
nor U22724 (N_22724,N_21529,N_22279);
nor U22725 (N_22725,N_21748,N_20596);
xnor U22726 (N_22726,N_21357,N_20911);
nand U22727 (N_22727,N_20347,N_20606);
and U22728 (N_22728,N_21899,N_22235);
or U22729 (N_22729,N_22415,N_21036);
nor U22730 (N_22730,N_22120,N_22278);
nand U22731 (N_22731,N_22196,N_20835);
nor U22732 (N_22732,N_20662,N_20899);
and U22733 (N_22733,N_20730,N_21358);
nor U22734 (N_22734,N_20429,N_21926);
nand U22735 (N_22735,N_22189,N_20902);
xnor U22736 (N_22736,N_22318,N_22164);
nand U22737 (N_22737,N_20573,N_21274);
and U22738 (N_22738,N_21207,N_21789);
or U22739 (N_22739,N_20180,N_20965);
or U22740 (N_22740,N_22452,N_21716);
nand U22741 (N_22741,N_21472,N_20335);
xor U22742 (N_22742,N_20981,N_20231);
xor U22743 (N_22743,N_22228,N_21376);
nand U22744 (N_22744,N_20438,N_21516);
nand U22745 (N_22745,N_21135,N_20264);
nor U22746 (N_22746,N_22422,N_20810);
or U22747 (N_22747,N_20527,N_22219);
xnor U22748 (N_22748,N_21079,N_21970);
nor U22749 (N_22749,N_21113,N_22023);
nor U22750 (N_22750,N_22421,N_21316);
xnor U22751 (N_22751,N_21598,N_20579);
or U22752 (N_22752,N_21194,N_21299);
or U22753 (N_22753,N_21046,N_20084);
or U22754 (N_22754,N_20157,N_21626);
xnor U22755 (N_22755,N_21915,N_21471);
nor U22756 (N_22756,N_20418,N_21982);
or U22757 (N_22757,N_20190,N_21363);
nor U22758 (N_22758,N_22287,N_21087);
nand U22759 (N_22759,N_20852,N_22285);
xor U22760 (N_22760,N_20986,N_21035);
xnor U22761 (N_22761,N_20535,N_20983);
nor U22762 (N_22762,N_21800,N_21263);
xnor U22763 (N_22763,N_20060,N_21646);
and U22764 (N_22764,N_20913,N_20713);
nand U22765 (N_22765,N_20170,N_21479);
xnor U22766 (N_22766,N_20954,N_21186);
nor U22767 (N_22767,N_21226,N_21679);
or U22768 (N_22768,N_21594,N_22418);
nand U22769 (N_22769,N_21272,N_20428);
xnor U22770 (N_22770,N_20992,N_22002);
or U22771 (N_22771,N_21727,N_21608);
or U22772 (N_22772,N_20063,N_20521);
nor U22773 (N_22773,N_21796,N_21771);
nand U22774 (N_22774,N_21393,N_20078);
nand U22775 (N_22775,N_22405,N_21417);
xor U22776 (N_22776,N_20254,N_21253);
and U22777 (N_22777,N_21911,N_21638);
nand U22778 (N_22778,N_20075,N_20199);
nand U22779 (N_22779,N_20871,N_20565);
and U22780 (N_22780,N_21615,N_20895);
xor U22781 (N_22781,N_20089,N_22420);
and U22782 (N_22782,N_20461,N_20331);
nand U22783 (N_22783,N_20691,N_22358);
xnor U22784 (N_22784,N_21900,N_20993);
nor U22785 (N_22785,N_20806,N_21201);
xnor U22786 (N_22786,N_21632,N_21710);
and U22787 (N_22787,N_22124,N_20833);
or U22788 (N_22788,N_21535,N_21031);
and U22789 (N_22789,N_22063,N_22499);
nand U22790 (N_22790,N_22381,N_21123);
xor U22791 (N_22791,N_21640,N_20843);
or U22792 (N_22792,N_20304,N_22394);
nand U22793 (N_22793,N_20589,N_21887);
and U22794 (N_22794,N_20877,N_21543);
nand U22795 (N_22795,N_21438,N_22324);
xnor U22796 (N_22796,N_22075,N_21581);
nand U22797 (N_22797,N_22018,N_21096);
nor U22798 (N_22798,N_21795,N_20837);
and U22799 (N_22799,N_20607,N_20740);
xor U22800 (N_22800,N_20433,N_20975);
and U22801 (N_22801,N_22362,N_20540);
or U22802 (N_22802,N_22050,N_22174);
and U22803 (N_22803,N_21038,N_21371);
or U22804 (N_22804,N_22294,N_20144);
xnor U22805 (N_22805,N_21190,N_22369);
nand U22806 (N_22806,N_21863,N_20367);
and U22807 (N_22807,N_21898,N_20148);
nand U22808 (N_22808,N_21807,N_20946);
nor U22809 (N_22809,N_21374,N_21341);
nor U22810 (N_22810,N_21838,N_20795);
nand U22811 (N_22811,N_20457,N_21798);
nor U22812 (N_22812,N_20001,N_21039);
and U22813 (N_22813,N_21961,N_21856);
and U22814 (N_22814,N_21280,N_22303);
or U22815 (N_22815,N_20138,N_21797);
or U22816 (N_22816,N_20772,N_22482);
nor U22817 (N_22817,N_21399,N_22295);
or U22818 (N_22818,N_20562,N_21199);
nand U22819 (N_22819,N_21457,N_21271);
or U22820 (N_22820,N_21267,N_22106);
nand U22821 (N_22821,N_20948,N_20255);
and U22822 (N_22822,N_21459,N_22112);
nor U22823 (N_22823,N_20647,N_22317);
nand U22824 (N_22824,N_21963,N_20901);
nand U22825 (N_22825,N_20725,N_20187);
or U22826 (N_22826,N_22217,N_21282);
and U22827 (N_22827,N_21688,N_20373);
or U22828 (N_22828,N_21068,N_21331);
or U22829 (N_22829,N_21674,N_21612);
nor U22830 (N_22830,N_21524,N_21008);
or U22831 (N_22831,N_21580,N_21858);
and U22832 (N_22832,N_20313,N_22073);
nand U22833 (N_22833,N_20593,N_20029);
nor U22834 (N_22834,N_20670,N_20564);
xnor U22835 (N_22835,N_22069,N_20099);
nor U22836 (N_22836,N_22332,N_21125);
and U22837 (N_22837,N_20757,N_20460);
and U22838 (N_22838,N_22473,N_21265);
nand U22839 (N_22839,N_20776,N_22005);
xor U22840 (N_22840,N_21232,N_20020);
and U22841 (N_22841,N_21380,N_21793);
nor U22842 (N_22842,N_20450,N_20393);
nand U22843 (N_22843,N_21990,N_22137);
or U22844 (N_22844,N_20853,N_21918);
or U22845 (N_22845,N_21475,N_20419);
nand U22846 (N_22846,N_21360,N_22437);
nand U22847 (N_22847,N_21662,N_22177);
and U22848 (N_22848,N_22460,N_21419);
or U22849 (N_22849,N_21320,N_21540);
and U22850 (N_22850,N_20690,N_22116);
nor U22851 (N_22851,N_21389,N_22494);
or U22852 (N_22852,N_20507,N_22039);
nand U22853 (N_22853,N_20880,N_22222);
or U22854 (N_22854,N_22220,N_21569);
and U22855 (N_22855,N_22289,N_22468);
nor U22856 (N_22856,N_21894,N_22229);
and U22857 (N_22857,N_21490,N_22291);
or U22858 (N_22858,N_21812,N_20401);
nand U22859 (N_22859,N_20550,N_20947);
and U22860 (N_22860,N_20094,N_22311);
or U22861 (N_22861,N_21621,N_21988);
and U22862 (N_22862,N_20057,N_22267);
nor U22863 (N_22863,N_20631,N_22254);
or U22864 (N_22864,N_21895,N_22240);
nor U22865 (N_22865,N_20277,N_21844);
xor U22866 (N_22866,N_21153,N_21021);
nand U22867 (N_22867,N_20621,N_21763);
nor U22868 (N_22868,N_22147,N_22429);
nand U22869 (N_22869,N_20137,N_21542);
xor U22870 (N_22870,N_21682,N_21995);
nor U22871 (N_22871,N_21493,N_20683);
nor U22872 (N_22872,N_20604,N_22172);
xnor U22873 (N_22873,N_22143,N_21649);
or U22874 (N_22874,N_21952,N_21209);
or U22875 (N_22875,N_20555,N_20729);
or U22876 (N_22876,N_22008,N_21003);
nor U22877 (N_22877,N_21996,N_21426);
xnor U22878 (N_22878,N_21109,N_22140);
and U22879 (N_22879,N_22492,N_21002);
nand U22880 (N_22880,N_20265,N_22331);
and U22881 (N_22881,N_20408,N_20326);
and U22882 (N_22882,N_20960,N_21301);
or U22883 (N_22883,N_21436,N_21482);
or U22884 (N_22884,N_20551,N_20437);
nand U22885 (N_22885,N_20184,N_20867);
nor U22886 (N_22886,N_20797,N_21214);
nand U22887 (N_22887,N_21070,N_21861);
nor U22888 (N_22888,N_20205,N_20435);
nand U22889 (N_22889,N_21847,N_20167);
nand U22890 (N_22890,N_21853,N_21881);
nor U22891 (N_22891,N_22212,N_21705);
nor U22892 (N_22892,N_22336,N_21213);
or U22893 (N_22893,N_22224,N_22395);
nor U22894 (N_22894,N_20364,N_21801);
nand U22895 (N_22895,N_20466,N_22268);
nor U22896 (N_22896,N_22408,N_21905);
and U22897 (N_22897,N_20387,N_21140);
or U22898 (N_22898,N_20140,N_21762);
or U22899 (N_22899,N_22386,N_20767);
or U22900 (N_22900,N_21955,N_22277);
and U22901 (N_22901,N_21848,N_21605);
or U22902 (N_22902,N_20887,N_20319);
or U22903 (N_22903,N_22489,N_21391);
or U22904 (N_22904,N_20480,N_20727);
or U22905 (N_22905,N_20352,N_22031);
nor U22906 (N_22906,N_20494,N_21016);
and U22907 (N_22907,N_21528,N_20559);
and U22908 (N_22908,N_22479,N_21527);
nor U22909 (N_22909,N_21137,N_20071);
and U22910 (N_22910,N_22009,N_21697);
nor U22911 (N_22911,N_20719,N_21311);
nor U22912 (N_22912,N_20937,N_20963);
or U22913 (N_22913,N_20876,N_21834);
or U22914 (N_22914,N_22435,N_20545);
or U22915 (N_22915,N_20207,N_22340);
and U22916 (N_22916,N_20781,N_22427);
xor U22917 (N_22917,N_22432,N_20193);
xor U22918 (N_22918,N_20610,N_21089);
and U22919 (N_22919,N_21663,N_21929);
nand U22920 (N_22920,N_21370,N_20787);
or U22921 (N_22921,N_20439,N_20892);
or U22922 (N_22922,N_20374,N_20842);
and U22923 (N_22923,N_20649,N_21344);
or U22924 (N_22924,N_21704,N_20355);
and U22925 (N_22925,N_22151,N_22077);
or U22926 (N_22926,N_20216,N_21044);
and U22927 (N_22927,N_21439,N_20445);
or U22928 (N_22928,N_20120,N_21714);
or U22929 (N_22929,N_20789,N_21015);
or U22930 (N_22930,N_20462,N_20420);
xnor U22931 (N_22931,N_22313,N_21369);
or U22932 (N_22932,N_20273,N_20321);
and U22933 (N_22933,N_21782,N_20511);
nor U22934 (N_22934,N_21256,N_22047);
and U22935 (N_22935,N_20554,N_21588);
or U22936 (N_22936,N_21453,N_21112);
or U22937 (N_22937,N_22273,N_20107);
and U22938 (N_22938,N_20238,N_20425);
xor U22939 (N_22939,N_20024,N_20332);
nand U22940 (N_22940,N_20820,N_20179);
and U22941 (N_22941,N_21388,N_21584);
nand U22942 (N_22942,N_20701,N_22180);
and U22943 (N_22943,N_20985,N_20085);
or U22944 (N_22944,N_22026,N_21578);
or U22945 (N_22945,N_20657,N_21349);
nor U22946 (N_22946,N_21707,N_20747);
nor U22947 (N_22947,N_21390,N_20955);
and U22948 (N_22948,N_20308,N_20318);
nor U22949 (N_22949,N_20746,N_21917);
nand U22950 (N_22950,N_20069,N_20376);
or U22951 (N_22951,N_21596,N_20497);
or U22952 (N_22952,N_20777,N_20919);
nand U22953 (N_22953,N_22095,N_20716);
nand U22954 (N_22954,N_20839,N_21174);
nor U22955 (N_22955,N_20223,N_21497);
nand U22956 (N_22956,N_22269,N_21088);
and U22957 (N_22957,N_22123,N_21127);
or U22958 (N_22958,N_21698,N_20040);
nand U22959 (N_22959,N_21276,N_22057);
nand U22960 (N_22960,N_20353,N_20337);
and U22961 (N_22961,N_20414,N_20643);
nor U22962 (N_22962,N_20964,N_20766);
nand U22963 (N_22963,N_20675,N_21959);
nor U22964 (N_22964,N_20143,N_21322);
or U22965 (N_22965,N_21967,N_20671);
xor U22966 (N_22966,N_20991,N_21579);
xor U22967 (N_22967,N_21218,N_20356);
or U22968 (N_22968,N_20582,N_20224);
xor U22969 (N_22969,N_20430,N_21837);
nand U22970 (N_22970,N_20941,N_22406);
nor U22971 (N_22971,N_20744,N_22379);
or U22972 (N_22972,N_21998,N_21514);
nor U22973 (N_22973,N_22250,N_22459);
xor U22974 (N_22974,N_22121,N_20953);
and U22975 (N_22975,N_21840,N_22141);
nor U22976 (N_22976,N_21069,N_21298);
or U22977 (N_22977,N_20546,N_21339);
nand U22978 (N_22978,N_22328,N_21262);
xor U22979 (N_22979,N_20987,N_20995);
xor U22980 (N_22980,N_22275,N_21356);
and U22981 (N_22981,N_22329,N_20237);
or U22982 (N_22982,N_20968,N_20646);
xnor U22983 (N_22983,N_21851,N_22074);
or U22984 (N_22984,N_20469,N_20505);
and U22985 (N_22985,N_21330,N_21484);
or U22986 (N_22986,N_21032,N_20384);
and U22987 (N_22987,N_21428,N_22356);
and U22988 (N_22988,N_20759,N_21597);
and U22989 (N_22989,N_21548,N_22388);
and U22990 (N_22990,N_20266,N_21980);
nor U22991 (N_22991,N_20536,N_20209);
nand U22992 (N_22992,N_22360,N_21162);
and U22993 (N_22993,N_20495,N_21896);
or U22994 (N_22994,N_22084,N_20552);
or U22995 (N_22995,N_21239,N_22365);
nand U22996 (N_22996,N_20176,N_21627);
nand U22997 (N_22997,N_20863,N_21081);
or U22998 (N_22998,N_20630,N_22446);
nor U22999 (N_22999,N_20856,N_20385);
xnor U23000 (N_23000,N_22207,N_20836);
nand U23001 (N_23001,N_20660,N_20769);
or U23002 (N_23002,N_20870,N_20047);
xnor U23003 (N_23003,N_22357,N_21665);
or U23004 (N_23004,N_21616,N_22129);
and U23005 (N_23005,N_22197,N_21939);
and U23006 (N_23006,N_20651,N_22467);
xnor U23007 (N_23007,N_20693,N_21396);
xor U23008 (N_23008,N_21169,N_21166);
nand U23009 (N_23009,N_20296,N_20097);
nor U23010 (N_23010,N_22284,N_21554);
and U23011 (N_23011,N_20218,N_21875);
xnor U23012 (N_23012,N_21504,N_20848);
and U23013 (N_23013,N_21891,N_21462);
and U23014 (N_23014,N_21564,N_21928);
nand U23015 (N_23015,N_20302,N_20522);
or U23016 (N_23016,N_20451,N_22445);
nand U23017 (N_23017,N_20997,N_21619);
or U23018 (N_23018,N_21126,N_20807);
xor U23019 (N_23019,N_22128,N_21159);
xor U23020 (N_23020,N_22099,N_21932);
or U23021 (N_23021,N_22041,N_22423);
nor U23022 (N_23022,N_20907,N_20282);
nand U23023 (N_23023,N_20360,N_22037);
or U23024 (N_23024,N_20929,N_21971);
nand U23025 (N_23025,N_22370,N_22447);
nor U23026 (N_23026,N_20182,N_22263);
xnor U23027 (N_23027,N_22321,N_20169);
nand U23028 (N_23028,N_22155,N_21481);
nand U23029 (N_23029,N_21950,N_21355);
xnor U23030 (N_23030,N_21994,N_21102);
nand U23031 (N_23031,N_20363,N_20105);
and U23032 (N_23032,N_20845,N_20015);
nand U23033 (N_23033,N_21195,N_20637);
xor U23034 (N_23034,N_21983,N_21683);
nand U23035 (N_23035,N_21178,N_22307);
or U23036 (N_23036,N_20966,N_20636);
and U23037 (N_23037,N_22450,N_21117);
or U23038 (N_23038,N_20653,N_20164);
xor U23039 (N_23039,N_20239,N_21273);
xor U23040 (N_23040,N_21968,N_20584);
or U23041 (N_23041,N_20510,N_21882);
or U23042 (N_23042,N_21483,N_20378);
and U23043 (N_23043,N_20912,N_20838);
or U23044 (N_23044,N_20720,N_22081);
nand U23045 (N_23045,N_22082,N_22044);
or U23046 (N_23046,N_21818,N_20113);
and U23047 (N_23047,N_20454,N_20052);
nand U23048 (N_23048,N_20090,N_20696);
nand U23049 (N_23049,N_22440,N_20917);
nor U23050 (N_23050,N_20348,N_21026);
xnor U23051 (N_23051,N_21492,N_20294);
and U23052 (N_23052,N_20597,N_21083);
and U23053 (N_23053,N_21521,N_21223);
xnor U23054 (N_23054,N_21047,N_20805);
and U23055 (N_23055,N_20724,N_21447);
and U23056 (N_23056,N_22425,N_21940);
and U23057 (N_23057,N_21814,N_22401);
and U23058 (N_23058,N_21440,N_22251);
nor U23059 (N_23059,N_21842,N_21277);
nor U23060 (N_23060,N_20006,N_20635);
xnor U23061 (N_23061,N_20116,N_20504);
or U23062 (N_23062,N_21586,N_20788);
xnor U23063 (N_23063,N_20149,N_21237);
or U23064 (N_23064,N_20027,N_21976);
nor U23065 (N_23065,N_21949,N_21733);
nor U23066 (N_23066,N_20676,N_20898);
and U23067 (N_23067,N_20410,N_21760);
xnor U23068 (N_23068,N_21054,N_20016);
xor U23069 (N_23069,N_21407,N_20627);
nand U23070 (N_23070,N_21204,N_20935);
nand U23071 (N_23071,N_21884,N_20340);
and U23072 (N_23072,N_20394,N_20530);
xnor U23073 (N_23073,N_21305,N_20121);
nand U23074 (N_23074,N_20990,N_22015);
and U23075 (N_23075,N_20000,N_21056);
nor U23076 (N_23076,N_20703,N_21200);
xnor U23077 (N_23077,N_22296,N_21222);
nor U23078 (N_23078,N_21245,N_20674);
nand U23079 (N_23079,N_21429,N_22078);
nand U23080 (N_23080,N_20624,N_21829);
and U23081 (N_23081,N_21737,N_22300);
and U23082 (N_23082,N_21852,N_20503);
and U23083 (N_23083,N_20303,N_20722);
nand U23084 (N_23084,N_21414,N_20581);
or U23085 (N_23085,N_20195,N_21839);
nand U23086 (N_23086,N_20477,N_21664);
nor U23087 (N_23087,N_21592,N_20188);
nor U23088 (N_23088,N_22402,N_21902);
and U23089 (N_23089,N_22157,N_20159);
nor U23090 (N_23090,N_22308,N_20305);
xor U23091 (N_23091,N_21769,N_20298);
or U23092 (N_23092,N_20984,N_21424);
nor U23093 (N_23093,N_21599,N_22274);
xnor U23094 (N_23094,N_21409,N_21346);
nor U23095 (N_23095,N_21835,N_22021);
nor U23096 (N_23096,N_20345,N_22153);
nand U23097 (N_23097,N_21650,N_22016);
and U23098 (N_23098,N_21176,N_21114);
xnor U23099 (N_23099,N_21750,N_21270);
nand U23100 (N_23100,N_21791,N_21525);
and U23101 (N_23101,N_22159,N_20310);
and U23102 (N_23102,N_21082,N_20289);
nand U23103 (N_23103,N_21318,N_20487);
or U23104 (N_23104,N_22352,N_21474);
nand U23105 (N_23105,N_20750,N_22210);
nand U23106 (N_23106,N_20652,N_21383);
nor U23107 (N_23107,N_21397,N_21713);
and U23108 (N_23108,N_21146,N_21086);
and U23109 (N_23109,N_21211,N_20988);
or U23110 (N_23110,N_20514,N_21746);
nand U23111 (N_23111,N_20881,N_21154);
nor U23112 (N_23112,N_20026,N_22337);
xnor U23113 (N_23113,N_21966,N_20755);
or U23114 (N_23114,N_20283,N_20846);
nor U23115 (N_23115,N_21156,N_21947);
or U23116 (N_23116,N_20272,N_21558);
nor U23117 (N_23117,N_20110,N_20575);
and U23118 (N_23118,N_21430,N_22327);
or U23119 (N_23119,N_21777,N_20537);
nor U23120 (N_23120,N_21922,N_21846);
and U23121 (N_23121,N_22366,N_21094);
or U23122 (N_23122,N_22072,N_20547);
and U23123 (N_23123,N_20012,N_22442);
xnor U23124 (N_23124,N_20531,N_22126);
and U23125 (N_23125,N_20244,N_20151);
nor U23126 (N_23126,N_20680,N_22490);
and U23127 (N_23127,N_22237,N_20809);
nand U23128 (N_23128,N_21057,N_21060);
and U23129 (N_23129,N_21052,N_20232);
xor U23130 (N_23130,N_20017,N_20967);
nand U23131 (N_23131,N_21394,N_22097);
and U23132 (N_23132,N_20252,N_20458);
or U23133 (N_23133,N_20634,N_21603);
and U23134 (N_23134,N_22264,N_21652);
and U23135 (N_23135,N_21651,N_20762);
or U23136 (N_23136,N_20103,N_20594);
and U23137 (N_23137,N_21913,N_20844);
xor U23138 (N_23138,N_21890,N_22087);
xor U23139 (N_23139,N_20771,N_21648);
xor U23140 (N_23140,N_22019,N_20577);
nor U23141 (N_23141,N_20508,N_20661);
nand U23142 (N_23142,N_21090,N_22270);
xor U23143 (N_23143,N_20468,N_21544);
and U23144 (N_23144,N_22495,N_20798);
nor U23145 (N_23145,N_21192,N_21238);
nand U23146 (N_23146,N_22133,N_20506);
and U23147 (N_23147,N_20301,N_20008);
xnor U23148 (N_23148,N_21639,N_21067);
nand U23149 (N_23149,N_22297,N_20873);
nand U23150 (N_23150,N_20051,N_22045);
and U23151 (N_23151,N_21148,N_21613);
and U23152 (N_23152,N_20904,N_20032);
xnor U23153 (N_23153,N_20278,N_22441);
nor U23154 (N_23154,N_20743,N_20779);
or U23155 (N_23155,N_21865,N_21559);
xnor U23156 (N_23156,N_20672,N_21590);
xor U23157 (N_23157,N_20698,N_21307);
xnor U23158 (N_23158,N_20241,N_21065);
nand U23159 (N_23159,N_22485,N_20341);
or U23160 (N_23160,N_21477,N_20858);
nand U23161 (N_23161,N_22000,N_21936);
xnor U23162 (N_23162,N_20056,N_22241);
or U23163 (N_23163,N_22061,N_21912);
nand U23164 (N_23164,N_21470,N_20023);
or U23165 (N_23165,N_20129,N_21359);
or U23166 (N_23166,N_20028,N_20728);
and U23167 (N_23167,N_21868,N_22341);
xnor U23168 (N_23168,N_21566,N_22281);
nor U23169 (N_23169,N_21157,N_20295);
nand U23170 (N_23170,N_21361,N_21684);
xor U23171 (N_23171,N_21185,N_22080);
nand U23172 (N_23172,N_22079,N_21314);
xnor U23173 (N_23173,N_21418,N_21556);
nor U23174 (N_23174,N_21855,N_21319);
nand U23175 (N_23175,N_20498,N_20135);
nor U23176 (N_23176,N_22320,N_22330);
and U23177 (N_23177,N_22125,N_20493);
xor U23178 (N_23178,N_21300,N_20956);
or U23179 (N_23179,N_21624,N_21013);
nand U23180 (N_23180,N_21074,N_20622);
nand U23181 (N_23181,N_20782,N_20933);
xor U23182 (N_23182,N_21860,N_22234);
xnor U23183 (N_23183,N_21290,N_21486);
and U23184 (N_23184,N_21187,N_21136);
or U23185 (N_23185,N_21402,N_20106);
or U23186 (N_23186,N_21258,N_20065);
xor U23187 (N_23187,N_20127,N_20163);
or U23188 (N_23188,N_20851,N_20489);
or U23189 (N_23189,N_20463,N_20415);
nor U23190 (N_23190,N_21888,N_21173);
xnor U23191 (N_23191,N_22104,N_21701);
nand U23192 (N_23192,N_20404,N_20780);
or U23193 (N_23193,N_21444,N_21669);
xnor U23194 (N_23194,N_21500,N_21546);
xnor U23195 (N_23195,N_21909,N_21379);
or U23196 (N_23196,N_20043,N_20600);
nor U23197 (N_23197,N_22411,N_20515);
nor U23198 (N_23198,N_22231,N_20533);
nor U23199 (N_23199,N_21336,N_21738);
nor U23200 (N_23200,N_21110,N_21048);
and U23201 (N_23201,N_21831,N_20174);
or U23202 (N_23202,N_21138,N_22469);
nand U23203 (N_23203,N_21823,N_20475);
and U23204 (N_23204,N_20633,N_20544);
nor U23205 (N_23205,N_21410,N_20763);
nor U23206 (N_23206,N_22384,N_21105);
nand U23207 (N_23207,N_20476,N_21676);
or U23208 (N_23208,N_21799,N_21531);
nor U23209 (N_23209,N_20192,N_22385);
nor U23210 (N_23210,N_22130,N_20799);
xnor U23211 (N_23211,N_20685,N_22288);
nand U23212 (N_23212,N_20602,N_22017);
and U23213 (N_23213,N_21235,N_22348);
or U23214 (N_23214,N_22060,N_22108);
and U23215 (N_23215,N_21602,N_21350);
nor U23216 (N_23216,N_22033,N_21230);
xor U23217 (N_23217,N_21133,N_21217);
or U23218 (N_23218,N_20288,N_20219);
nand U23219 (N_23219,N_21124,N_21671);
or U23220 (N_23220,N_21583,N_22322);
nor U23221 (N_23221,N_20381,N_22059);
nor U23222 (N_23222,N_21055,N_21809);
nand U23223 (N_23223,N_20979,N_21589);
xor U23224 (N_23224,N_22449,N_21141);
nor U23225 (N_23225,N_21567,N_21794);
or U23226 (N_23226,N_22025,N_20639);
xnor U23227 (N_23227,N_20286,N_22181);
and U23228 (N_23228,N_21722,N_20038);
xor U23229 (N_23229,N_21405,N_21184);
nor U23230 (N_23230,N_21175,N_20751);
nor U23231 (N_23231,N_20760,N_21553);
or U23232 (N_23232,N_21248,N_22169);
xor U23233 (N_23233,N_22195,N_21693);
and U23234 (N_23234,N_22064,N_22201);
and U23235 (N_23235,N_21351,N_20700);
nand U23236 (N_23236,N_20191,N_20903);
xnor U23237 (N_23237,N_22349,N_22310);
nand U23238 (N_23238,N_20970,N_20399);
or U23239 (N_23239,N_21675,N_20490);
xnor U23240 (N_23240,N_20124,N_22272);
nor U23241 (N_23241,N_21552,N_22156);
and U23242 (N_23242,N_20794,N_21979);
or U23243 (N_23243,N_22374,N_21808);
or U23244 (N_23244,N_22397,N_21827);
xor U23245 (N_23245,N_22158,N_22400);
nand U23246 (N_23246,N_20524,N_22433);
nand U23247 (N_23247,N_20526,N_21885);
or U23248 (N_23248,N_20982,N_22184);
nand U23249 (N_23249,N_22034,N_20091);
nor U23250 (N_23250,N_22293,N_20874);
or U23251 (N_23251,N_22208,N_21193);
xnor U23252 (N_23252,N_22239,N_20525);
xnor U23253 (N_23253,N_21403,N_22413);
nand U23254 (N_23254,N_22233,N_20396);
xor U23255 (N_23255,N_21340,N_21064);
or U23256 (N_23256,N_21463,N_20455);
nand U23257 (N_23257,N_21655,N_21071);
xnor U23258 (N_23258,N_21489,N_21338);
nor U23259 (N_23259,N_20386,N_21279);
or U23260 (N_23260,N_20004,N_20945);
nand U23261 (N_23261,N_22096,N_20424);
xor U23262 (N_23262,N_22403,N_22211);
xor U23263 (N_23263,N_22191,N_20813);
and U23264 (N_23264,N_21862,N_21269);
xnor U23265 (N_23265,N_20371,N_20036);
or U23266 (N_23266,N_20464,N_21617);
xor U23267 (N_23267,N_21660,N_20212);
nor U23268 (N_23268,N_22067,N_22375);
and U23269 (N_23269,N_21719,N_22286);
or U23270 (N_23270,N_21427,N_20930);
or U23271 (N_23271,N_21203,N_21765);
nand U23272 (N_23272,N_20389,N_20235);
xnor U23273 (N_23273,N_21743,N_20059);
nand U23274 (N_23274,N_20485,N_21702);
or U23275 (N_23275,N_20891,N_22040);
or U23276 (N_23276,N_22377,N_22146);
and U23277 (N_23277,N_20442,N_21781);
nand U23278 (N_23278,N_20978,N_21897);
xnor U23279 (N_23279,N_20092,N_21833);
or U23280 (N_23280,N_20854,N_22302);
and U23281 (N_23281,N_20236,N_22451);
and U23282 (N_23282,N_21850,N_20181);
nand U23283 (N_23283,N_22085,N_20765);
and U23284 (N_23284,N_20764,N_21121);
or U23285 (N_23285,N_21986,N_22434);
and U23286 (N_23286,N_22136,N_20603);
nand U23287 (N_23287,N_21570,N_20726);
xor U23288 (N_23288,N_21872,N_21587);
or U23289 (N_23289,N_20567,N_20754);
or U23290 (N_23290,N_20233,N_22139);
and U23291 (N_23291,N_22013,N_22399);
and U23292 (N_23292,N_21004,N_21859);
or U23293 (N_23293,N_22138,N_20585);
or U23294 (N_23294,N_21326,N_21189);
nor U23295 (N_23295,N_21303,N_21715);
xnor U23296 (N_23296,N_20821,N_21261);
and U23297 (N_23297,N_21329,N_20325);
nand U23298 (N_23298,N_20253,N_20132);
and U23299 (N_23299,N_22194,N_21942);
and U23300 (N_23300,N_22481,N_20031);
xnor U23301 (N_23301,N_20398,N_20427);
and U23302 (N_23302,N_20784,N_21680);
xor U23303 (N_23303,N_20513,N_22012);
nor U23304 (N_23304,N_21870,N_22367);
or U23305 (N_23305,N_22246,N_21401);
and U23306 (N_23306,N_21574,N_21645);
and U23307 (N_23307,N_22419,N_21281);
nand U23308 (N_23308,N_22249,N_20642);
or U23309 (N_23309,N_22165,N_22248);
or U23310 (N_23310,N_21045,N_22117);
and U23311 (N_23311,N_21255,N_20082);
or U23312 (N_23312,N_21155,N_20440);
nand U23313 (N_23313,N_22280,N_20257);
or U23314 (N_23314,N_21384,N_21229);
or U23315 (N_23315,N_21991,N_22192);
or U23316 (N_23316,N_20362,N_21412);
or U23317 (N_23317,N_22188,N_20293);
and U23318 (N_23318,N_21152,N_20829);
and U23319 (N_23319,N_20222,N_21241);
nand U23320 (N_23320,N_21415,N_21547);
xor U23321 (N_23321,N_21347,N_21510);
and U23322 (N_23322,N_22238,N_21997);
nand U23323 (N_23323,N_22115,N_21205);
or U23324 (N_23324,N_21520,N_21129);
xor U23325 (N_23325,N_21496,N_21233);
nor U23326 (N_23326,N_20539,N_22380);
or U23327 (N_23327,N_21010,N_21455);
nand U23328 (N_23328,N_20578,N_22076);
nand U23329 (N_23329,N_20859,N_22304);
nor U23330 (N_23330,N_22315,N_21634);
and U23331 (N_23331,N_20793,N_21050);
nand U23332 (N_23332,N_20196,N_21778);
nor U23333 (N_23333,N_20650,N_22387);
xnor U23334 (N_23334,N_21122,N_22335);
xor U23335 (N_23335,N_22049,N_22127);
nand U23336 (N_23336,N_22230,N_22347);
or U23337 (N_23337,N_20708,N_22391);
nor U23338 (N_23338,N_20465,N_22487);
nor U23339 (N_23339,N_21180,N_21854);
nor U23340 (N_23340,N_21242,N_20066);
nor U23341 (N_23341,N_20342,N_21043);
and U23342 (N_23342,N_21822,N_21130);
xnor U23343 (N_23343,N_21572,N_21028);
or U23344 (N_23344,N_20141,N_22202);
and U23345 (N_23345,N_22176,N_21445);
or U23346 (N_23346,N_21421,N_20261);
and U23347 (N_23347,N_22343,N_20548);
and U23348 (N_23348,N_20467,N_22316);
nor U23349 (N_23349,N_20566,N_21678);
or U23350 (N_23350,N_21100,N_20185);
xor U23351 (N_23351,N_22088,N_20422);
and U23352 (N_23352,N_21873,N_20274);
and U23353 (N_23353,N_22216,N_21313);
nand U23354 (N_23354,N_20479,N_21690);
and U23355 (N_23355,N_21803,N_20339);
xor U23356 (N_23356,N_22430,N_22170);
and U23357 (N_23357,N_20139,N_21448);
xor U23358 (N_23358,N_21712,N_20611);
or U23359 (N_23359,N_22493,N_21742);
nor U23360 (N_23360,N_21480,N_21637);
xnor U23361 (N_23361,N_21864,N_21907);
nand U23362 (N_23362,N_20013,N_21773);
or U23363 (N_23363,N_22257,N_20316);
nor U23364 (N_23364,N_20380,N_20923);
or U23365 (N_23365,N_22052,N_21011);
nand U23366 (N_23366,N_22498,N_21297);
nor U23367 (N_23367,N_22376,N_20245);
and U23368 (N_23368,N_21633,N_22346);
and U23369 (N_23369,N_22382,N_22028);
and U23370 (N_23370,N_20641,N_22243);
nor U23371 (N_23371,N_20614,N_20168);
or U23372 (N_23372,N_21364,N_20290);
or U23373 (N_23373,N_21170,N_20173);
and U23374 (N_23374,N_21787,N_21630);
xor U23375 (N_23375,N_20519,N_22144);
or U23376 (N_23376,N_21686,N_21756);
xnor U23377 (N_23377,N_20083,N_22414);
or U23378 (N_23378,N_20796,N_21250);
and U23379 (N_23379,N_20894,N_20206);
nand U23380 (N_23380,N_21285,N_20878);
or U23381 (N_23381,N_20242,N_20770);
or U23382 (N_23382,N_21538,N_20574);
nand U23383 (N_23383,N_20974,N_20299);
or U23384 (N_23384,N_22161,N_20834);
xnor U23385 (N_23385,N_21063,N_21754);
nand U23386 (N_23386,N_20230,N_20756);
or U23387 (N_23387,N_20240,N_21099);
or U23388 (N_23388,N_22471,N_20861);
or U23389 (N_23389,N_21147,N_20802);
nand U23390 (N_23390,N_21335,N_20131);
nor U23391 (N_23391,N_20100,N_22190);
nor U23392 (N_23392,N_20072,N_20101);
and U23393 (N_23393,N_20502,N_22283);
nand U23394 (N_23394,N_20686,N_21254);
or U23395 (N_23395,N_22431,N_21930);
nor U23396 (N_23396,N_22245,N_22101);
or U23397 (N_23397,N_20826,N_20007);
nand U23398 (N_23398,N_20452,N_21755);
nor U23399 (N_23399,N_21334,N_21636);
xor U23400 (N_23400,N_22109,N_21804);
and U23401 (N_23401,N_21513,N_21745);
xor U23402 (N_23402,N_22372,N_22163);
nand U23403 (N_23403,N_22135,N_22226);
or U23404 (N_23404,N_21530,N_21824);
or U23405 (N_23405,N_21181,N_20534);
or U23406 (N_23406,N_21191,N_20070);
or U23407 (N_23407,N_20323,N_21061);
nor U23408 (N_23408,N_20400,N_20656);
xor U23409 (N_23409,N_21108,N_20492);
or U23410 (N_23410,N_21774,N_20959);
nor U23411 (N_23411,N_20197,N_22426);
nand U23412 (N_23412,N_21246,N_20663);
and U23413 (N_23413,N_20523,N_22068);
nand U23414 (N_23414,N_20669,N_20204);
nor U23415 (N_23415,N_20058,N_21423);
nor U23416 (N_23416,N_21150,N_21101);
and U23417 (N_23417,N_21867,N_20916);
or U23418 (N_23418,N_21658,N_20225);
nand U23419 (N_23419,N_20077,N_20251);
nor U23420 (N_23420,N_20645,N_22223);
nand U23421 (N_23421,N_22178,N_21144);
xor U23422 (N_23422,N_21565,N_21757);
nand U23423 (N_23423,N_21509,N_21720);
xnor U23424 (N_23424,N_21009,N_21284);
or U23425 (N_23425,N_22457,N_21343);
nand U23426 (N_23426,N_21694,N_22378);
and U23427 (N_23427,N_22326,N_20046);
nor U23428 (N_23428,N_21091,N_21965);
or U23429 (N_23429,N_20153,N_22056);
and U23430 (N_23430,N_20644,N_21308);
nand U23431 (N_23431,N_20972,N_21644);
xor U23432 (N_23432,N_21288,N_22314);
nand U23433 (N_23433,N_20285,N_21703);
nor U23434 (N_23434,N_21128,N_20366);
nor U23435 (N_23435,N_22252,N_21732);
nor U23436 (N_23436,N_20732,N_20025);
nor U23437 (N_23437,N_21606,N_22100);
nor U23438 (N_23438,N_20969,N_20840);
and U23439 (N_23439,N_20067,N_21725);
nor U23440 (N_23440,N_20333,N_22148);
nand U23441 (N_23441,N_21132,N_20791);
xnor U23442 (N_23442,N_21437,N_20416);
xor U23443 (N_23443,N_22114,N_20434);
nand U23444 (N_23444,N_21324,N_20221);
xnor U23445 (N_23445,N_20734,N_21212);
and U23446 (N_23446,N_21964,N_21943);
and U23447 (N_23447,N_20473,N_20617);
nor U23448 (N_23448,N_20591,N_20609);
or U23449 (N_23449,N_21987,N_22488);
nor U23450 (N_23450,N_20702,N_21368);
xnor U23451 (N_23451,N_20049,N_21161);
and U23452 (N_23452,N_20249,N_20423);
or U23453 (N_23453,N_20774,N_20687);
xnor U23454 (N_23454,N_22083,N_20178);
and U23455 (N_23455,N_21729,N_21815);
and U23456 (N_23456,N_20961,N_21066);
nand U23457 (N_23457,N_20287,N_22011);
nand U23458 (N_23458,N_20211,N_21539);
nand U23459 (N_23459,N_20314,N_20932);
nand U23460 (N_23460,N_21761,N_22065);
and U23461 (N_23461,N_21768,N_20971);
and U23462 (N_23462,N_21452,N_21813);
xor U23463 (N_23463,N_22364,N_20306);
xor U23464 (N_23464,N_21944,N_21228);
nand U23465 (N_23465,N_22290,N_20154);
and U23466 (N_23466,N_22404,N_21078);
or U23467 (N_23467,N_22232,N_20317);
nor U23468 (N_23468,N_20697,N_20118);
nand U23469 (N_23469,N_20330,N_22004);
nand U23470 (N_23470,N_20171,N_21999);
nand U23471 (N_23471,N_21788,N_20847);
nor U23472 (N_23472,N_21790,N_22110);
or U23473 (N_23473,N_20421,N_20263);
nand U23474 (N_23474,N_20392,N_20571);
xor U23475 (N_23475,N_20499,N_21784);
nand U23476 (N_23476,N_20816,N_21234);
and U23477 (N_23477,N_21375,N_20869);
and U23478 (N_23478,N_22209,N_20247);
and U23479 (N_23479,N_21876,N_22373);
nor U23480 (N_23480,N_21954,N_21673);
nor U23481 (N_23481,N_22094,N_22054);
nor U23482 (N_23482,N_20359,N_22058);
xor U23483 (N_23483,N_22070,N_22309);
xor U23484 (N_23484,N_21735,N_21231);
nor U23485 (N_23485,N_21059,N_21726);
nor U23486 (N_23486,N_21302,N_21661);
and U23487 (N_23487,N_21536,N_21404);
or U23488 (N_23488,N_20717,N_21874);
xnor U23489 (N_23489,N_21352,N_22089);
nor U23490 (N_23490,N_20640,N_21266);
nor U23491 (N_23491,N_22292,N_21576);
nor U23492 (N_23492,N_20890,N_22464);
nor U23493 (N_23493,N_22344,N_22455);
and U23494 (N_23494,N_21836,N_22142);
nand U23495 (N_23495,N_22003,N_20284);
nor U23496 (N_23496,N_20612,N_20449);
or U23497 (N_23497,N_20327,N_20999);
xnor U23498 (N_23498,N_21321,N_20758);
and U23499 (N_23499,N_20862,N_21171);
and U23500 (N_23500,N_20073,N_20383);
and U23501 (N_23501,N_20638,N_21259);
nor U23502 (N_23502,N_20673,N_21643);
or U23503 (N_23503,N_21670,N_20014);
and U23504 (N_23504,N_21406,N_21077);
and U23505 (N_23505,N_21177,N_20115);
nand U23506 (N_23506,N_20712,N_21443);
xor U23507 (N_23507,N_21557,N_21310);
and U23508 (N_23508,N_21734,N_20927);
or U23509 (N_23509,N_22149,N_20369);
or U23510 (N_23510,N_21160,N_20158);
nand U23511 (N_23511,N_20030,N_20632);
nand U23512 (N_23512,N_20866,N_21924);
or U23513 (N_23513,N_21515,N_21534);
or U23514 (N_23514,N_22051,N_20931);
or U23515 (N_23515,N_21764,N_20050);
xor U23516 (N_23516,N_20785,N_22466);
nand U23517 (N_23517,N_20134,N_21179);
and U23518 (N_23518,N_21744,N_22247);
or U23519 (N_23519,N_21817,N_21275);
and U23520 (N_23520,N_20557,N_21106);
nand U23521 (N_23521,N_20267,N_20616);
or U23522 (N_23522,N_22463,N_22368);
and U23523 (N_23523,N_21975,N_21656);
nor U23524 (N_23524,N_21163,N_22334);
or U23525 (N_23525,N_21857,N_21893);
nand U23526 (N_23526,N_22221,N_20448);
nand U23527 (N_23527,N_20064,N_21533);
xor U23528 (N_23528,N_21353,N_20409);
and U23529 (N_23529,N_22206,N_22183);
and U23530 (N_23530,N_21332,N_21871);
or U23531 (N_23531,N_22276,N_20011);
and U23532 (N_23532,N_20512,N_20035);
xor U23533 (N_23533,N_22225,N_20395);
nand U23534 (N_23534,N_20658,N_21904);
or U23535 (N_23535,N_21485,N_21526);
nor U23536 (N_23536,N_20119,N_20619);
nor U23537 (N_23537,N_21901,N_20309);
and U23538 (N_23538,N_22103,N_22265);
or U23539 (N_23539,N_21278,N_20117);
nand U23540 (N_23540,N_21283,N_21333);
nor U23541 (N_23541,N_21730,N_21667);
nand U23542 (N_23542,N_21073,N_22187);
xnor U23543 (N_23543,N_20668,N_21723);
or U23544 (N_23544,N_20626,N_21878);
nand U23545 (N_23545,N_20202,N_21550);
or U23546 (N_23546,N_21491,N_20114);
nand U23547 (N_23547,N_20827,N_21505);
or U23548 (N_23548,N_20357,N_21165);
xnor U23549 (N_23549,N_21507,N_22035);
and U23550 (N_23550,N_20905,N_20426);
or U23551 (N_23551,N_22193,N_21442);
nor U23552 (N_23552,N_22145,N_21654);
xor U23553 (N_23553,N_21920,N_21395);
or U23554 (N_23554,N_21075,N_20108);
nand U23555 (N_23555,N_20229,N_21551);
xor U23556 (N_23556,N_20021,N_22361);
nand U23557 (N_23557,N_20358,N_21921);
xor U23558 (N_23558,N_20857,N_21115);
nor U23559 (N_23559,N_21072,N_20104);
nand U23560 (N_23560,N_21511,N_20814);
or U23561 (N_23561,N_21450,N_22333);
xor U23562 (N_23562,N_20938,N_22393);
nand U23563 (N_23563,N_21972,N_20125);
xor U23564 (N_23564,N_22353,N_20291);
nand U23565 (N_23565,N_21989,N_20667);
or U23566 (N_23566,N_21906,N_21441);
or U23567 (N_23567,N_20281,N_20608);
and U23568 (N_23568,N_21149,N_21832);
and U23569 (N_23569,N_20563,N_21433);
and U23570 (N_23570,N_22132,N_20391);
and U23571 (N_23571,N_22462,N_20918);
or U23572 (N_23572,N_20568,N_21400);
and U23573 (N_23573,N_20786,N_20481);
nor U23574 (N_23574,N_20470,N_22102);
or U23575 (N_23575,N_20213,N_20811);
nand U23576 (N_23576,N_20920,N_21058);
nand U23577 (N_23577,N_20146,N_20695);
nand U23578 (N_23578,N_21040,N_21600);
nor U23579 (N_23579,N_22312,N_20201);
or U23580 (N_23580,N_21315,N_20520);
nor U23581 (N_23581,N_21549,N_21062);
xor U23582 (N_23582,N_21555,N_21958);
and U23583 (N_23583,N_21981,N_20177);
and U23584 (N_23584,N_21268,N_20269);
nand U23585 (N_23585,N_22443,N_22454);
nor U23586 (N_23586,N_20488,N_20136);
xor U23587 (N_23587,N_21819,N_21886);
and U23588 (N_23588,N_20889,N_20054);
and U23589 (N_23589,N_20710,N_20745);
xnor U23590 (N_23590,N_21677,N_20344);
nor U23591 (N_23591,N_21312,N_21467);
nand U23592 (N_23592,N_22470,N_20258);
nor U23593 (N_23593,N_21495,N_22010);
nand U23594 (N_23594,N_22105,N_22407);
and U23595 (N_23595,N_20042,N_22055);
and U23596 (N_23596,N_20150,N_21935);
nor U23597 (N_23597,N_21476,N_21591);
and U23598 (N_23598,N_22424,N_20825);
and U23599 (N_23599,N_21098,N_22200);
or U23600 (N_23600,N_21264,N_20112);
nor U23601 (N_23601,N_20592,N_20183);
xor U23602 (N_23602,N_21653,N_22306);
xnor U23603 (N_23603,N_20586,N_20875);
nor U23604 (N_23604,N_20496,N_20818);
and U23605 (N_23605,N_20208,N_22091);
or U23606 (N_23606,N_22383,N_20482);
nor U23607 (N_23607,N_20388,N_20553);
nand U23608 (N_23608,N_21260,N_20162);
nor U23609 (N_23609,N_20405,N_21385);
nand U23610 (N_23610,N_21458,N_21828);
and U23611 (N_23611,N_22027,N_20275);
or U23612 (N_23612,N_22042,N_20705);
xor U23613 (N_23613,N_22299,N_20888);
xnor U23614 (N_23614,N_21425,N_21747);
nor U23615 (N_23615,N_21642,N_22351);
or U23616 (N_23616,N_22236,N_22483);
or U23617 (N_23617,N_21018,N_22439);
nor U23618 (N_23618,N_20659,N_21142);
xor U23619 (N_23619,N_22167,N_21752);
nand U23620 (N_23620,N_20210,N_21367);
xor U23621 (N_23621,N_21017,N_20543);
nand U23622 (N_23622,N_20832,N_20868);
and U23623 (N_23623,N_20549,N_20655);
nor U23624 (N_23624,N_20694,N_20126);
nor U23625 (N_23625,N_20872,N_20155);
nand U23626 (N_23626,N_20315,N_20095);
or U23627 (N_23627,N_22086,N_22030);
nand U23628 (N_23628,N_21188,N_20778);
or U23629 (N_23629,N_20349,N_21687);
nand U23630 (N_23630,N_21304,N_21257);
xnor U23631 (N_23631,N_21593,N_21978);
and U23632 (N_23632,N_20733,N_20677);
nand U23633 (N_23633,N_20804,N_20598);
and U23634 (N_23634,N_22282,N_21164);
nor U23635 (N_23635,N_21488,N_21668);
xnor U23636 (N_23636,N_21006,N_20402);
nor U23637 (N_23637,N_20509,N_22001);
xnor U23638 (N_23638,N_20128,N_21097);
xnor U23639 (N_23639,N_21247,N_22022);
xnor U23640 (N_23640,N_22162,N_22409);
xor U23641 (N_23641,N_20234,N_20572);
xnor U23642 (N_23642,N_20145,N_22204);
nand U23643 (N_23643,N_22066,N_20886);
or U23644 (N_23644,N_21635,N_21236);
xor U23645 (N_23645,N_22175,N_22350);
and U23646 (N_23646,N_20980,N_21416);
nand U23647 (N_23647,N_20629,N_21119);
nor U23648 (N_23648,N_21582,N_20123);
and U23649 (N_23649,N_22396,N_21951);
nand U23650 (N_23650,N_20329,N_22461);
nand U23651 (N_23651,N_20382,N_21451);
nand U23652 (N_23652,N_21767,N_20994);
and U23653 (N_23653,N_20773,N_20018);
and U23654 (N_23654,N_21449,N_21711);
nand U23655 (N_23655,N_20989,N_21362);
xor U23656 (N_23656,N_21377,N_20098);
nor U23657 (N_23657,N_20122,N_21502);
or U23658 (N_23658,N_21139,N_20079);
nor U23659 (N_23659,N_20817,N_20292);
or U23660 (N_23660,N_20823,N_21825);
and U23661 (N_23661,N_21022,N_21093);
xnor U23662 (N_23662,N_22134,N_20346);
or U23663 (N_23663,N_21487,N_21198);
nand U23664 (N_23664,N_20431,N_20934);
and U23665 (N_23665,N_21811,N_20936);
or U23666 (N_23666,N_22355,N_20436);
and U23667 (N_23667,N_20039,N_20942);
xor U23668 (N_23668,N_22262,N_20142);
nand U23669 (N_23669,N_20664,N_20628);
nor U23670 (N_23670,N_21753,N_21934);
or U23671 (N_23671,N_22484,N_20343);
xor U23672 (N_23672,N_20962,N_20849);
or U23673 (N_23673,N_21691,N_21143);
and U23674 (N_23674,N_21512,N_22465);
nand U23675 (N_23675,N_20336,N_21869);
nand U23676 (N_23676,N_21025,N_22038);
xnor U23677 (N_23677,N_21625,N_20613);
xnor U23678 (N_23678,N_20615,N_20882);
xnor U23679 (N_23679,N_21931,N_22496);
or U23680 (N_23680,N_22410,N_22301);
nor U23681 (N_23681,N_20086,N_20977);
nor U23682 (N_23682,N_22428,N_20456);
xor U23683 (N_23683,N_21903,N_22389);
or U23684 (N_23684,N_20718,N_22266);
nor U23685 (N_23685,N_21946,N_20648);
and U23686 (N_23686,N_21962,N_20260);
xnor U23687 (N_23687,N_21629,N_20560);
or U23688 (N_23688,N_21518,N_20684);
nand U23689 (N_23689,N_20109,N_21523);
and U23690 (N_23690,N_20198,N_21770);
nand U23691 (N_23691,N_20721,N_22458);
and U23692 (N_23692,N_20354,N_22256);
and U23693 (N_23693,N_21030,N_20087);
and U23694 (N_23694,N_21342,N_21049);
nor U23695 (N_23695,N_20538,N_21577);
xor U23696 (N_23696,N_21741,N_20044);
nor U23697 (N_23697,N_21956,N_21498);
nand U23698 (N_23698,N_21933,N_21080);
or U23699 (N_23699,N_21910,N_20516);
and U23700 (N_23700,N_21751,N_20588);
and U23701 (N_23701,N_22417,N_22160);
xnor U23702 (N_23702,N_20957,N_20922);
nor U23703 (N_23703,N_20855,N_20300);
xnor U23704 (N_23704,N_21806,N_21672);
nor U23705 (N_23705,N_21221,N_20908);
or U23706 (N_23706,N_22199,N_20217);
or U23707 (N_23707,N_20735,N_20228);
nor U23708 (N_23708,N_21786,N_22444);
xnor U23709 (N_23709,N_21373,N_20093);
nand U23710 (N_23710,N_21501,N_21607);
xor U23711 (N_23711,N_21843,N_21076);
and U23712 (N_23712,N_22448,N_21420);
nor U23713 (N_23713,N_20742,N_20761);
or U23714 (N_23714,N_21689,N_20808);
nand U23715 (N_23715,N_21294,N_21251);
or U23716 (N_23716,N_21024,N_21348);
xnor U23717 (N_23717,N_21118,N_22168);
and U23718 (N_23718,N_22271,N_21916);
and U23719 (N_23719,N_20175,N_20665);
or U23720 (N_23720,N_21084,N_20850);
xnor U23721 (N_23721,N_20692,N_20443);
nor U23722 (N_23722,N_21623,N_22412);
nor U23723 (N_23723,N_21845,N_22014);
or U23724 (N_23724,N_20583,N_20883);
nand U23725 (N_23725,N_20441,N_21810);
or U23726 (N_23726,N_21206,N_20372);
and U23727 (N_23727,N_20411,N_22453);
nor U23728 (N_23728,N_21695,N_21029);
nand U23729 (N_23729,N_20062,N_20822);
or U23730 (N_23730,N_20556,N_20262);
nor U23731 (N_23731,N_20900,N_21456);
xor U23732 (N_23732,N_21609,N_21289);
nor U23733 (N_23733,N_20334,N_20831);
nor U23734 (N_23734,N_20279,N_22390);
nand U23735 (N_23735,N_21573,N_21537);
or U23736 (N_23736,N_20654,N_21866);
nor U23737 (N_23737,N_20200,N_20406);
nor U23738 (N_23738,N_20076,N_22111);
xnor U23739 (N_23739,N_20483,N_20297);
xnor U23740 (N_23740,N_21721,N_21614);
xor U23741 (N_23741,N_21151,N_20003);
nor U23742 (N_23742,N_22098,N_22339);
nor U23743 (N_23743,N_21758,N_20010);
or U23744 (N_23744,N_21622,N_20949);
nor U23745 (N_23745,N_20250,N_21345);
nor U23746 (N_23746,N_21422,N_20194);
nor U23747 (N_23747,N_21923,N_20019);
or U23748 (N_23748,N_22046,N_21183);
or U23749 (N_23749,N_21699,N_20801);
xor U23750 (N_23750,N_21127,N_21944);
or U23751 (N_23751,N_21724,N_22418);
and U23752 (N_23752,N_21133,N_21917);
or U23753 (N_23753,N_21756,N_20891);
or U23754 (N_23754,N_20246,N_20711);
and U23755 (N_23755,N_20968,N_20320);
and U23756 (N_23756,N_20823,N_20126);
nor U23757 (N_23757,N_20583,N_20295);
or U23758 (N_23758,N_21225,N_20415);
or U23759 (N_23759,N_22030,N_20556);
and U23760 (N_23760,N_20580,N_20994);
xnor U23761 (N_23761,N_22323,N_20469);
nor U23762 (N_23762,N_21826,N_20201);
and U23763 (N_23763,N_20444,N_21027);
nand U23764 (N_23764,N_21867,N_20967);
xor U23765 (N_23765,N_22419,N_21261);
and U23766 (N_23766,N_21490,N_21239);
and U23767 (N_23767,N_20415,N_21520);
or U23768 (N_23768,N_20251,N_22389);
nand U23769 (N_23769,N_21608,N_21613);
and U23770 (N_23770,N_20174,N_21103);
xor U23771 (N_23771,N_21102,N_20818);
and U23772 (N_23772,N_22084,N_21222);
and U23773 (N_23773,N_20740,N_21729);
or U23774 (N_23774,N_22010,N_20664);
or U23775 (N_23775,N_22172,N_20080);
nand U23776 (N_23776,N_20580,N_21051);
nand U23777 (N_23777,N_20066,N_20533);
nand U23778 (N_23778,N_21019,N_22318);
or U23779 (N_23779,N_21919,N_21553);
and U23780 (N_23780,N_21312,N_22456);
nor U23781 (N_23781,N_20572,N_22283);
nor U23782 (N_23782,N_20339,N_21716);
nor U23783 (N_23783,N_22484,N_20275);
xor U23784 (N_23784,N_21652,N_20533);
or U23785 (N_23785,N_22492,N_22110);
nand U23786 (N_23786,N_20461,N_21407);
nand U23787 (N_23787,N_22446,N_21531);
or U23788 (N_23788,N_20940,N_21365);
nand U23789 (N_23789,N_21332,N_22269);
or U23790 (N_23790,N_22313,N_20372);
or U23791 (N_23791,N_21385,N_22040);
and U23792 (N_23792,N_20717,N_20040);
xnor U23793 (N_23793,N_20142,N_20490);
and U23794 (N_23794,N_22016,N_21300);
xnor U23795 (N_23795,N_21291,N_20062);
nand U23796 (N_23796,N_21779,N_22462);
nor U23797 (N_23797,N_20601,N_20757);
nand U23798 (N_23798,N_21291,N_21166);
or U23799 (N_23799,N_22116,N_20106);
nor U23800 (N_23800,N_20318,N_20123);
xnor U23801 (N_23801,N_20957,N_20879);
nand U23802 (N_23802,N_20486,N_22034);
nor U23803 (N_23803,N_22349,N_20137);
and U23804 (N_23804,N_21957,N_22134);
and U23805 (N_23805,N_21261,N_20933);
xor U23806 (N_23806,N_21799,N_20380);
or U23807 (N_23807,N_21638,N_21155);
nand U23808 (N_23808,N_20669,N_21882);
nand U23809 (N_23809,N_20628,N_21797);
nand U23810 (N_23810,N_21037,N_20813);
and U23811 (N_23811,N_22163,N_20553);
or U23812 (N_23812,N_21276,N_20326);
xnor U23813 (N_23813,N_21218,N_22494);
and U23814 (N_23814,N_20612,N_20481);
and U23815 (N_23815,N_21655,N_20069);
and U23816 (N_23816,N_22098,N_21318);
nor U23817 (N_23817,N_20685,N_20696);
nand U23818 (N_23818,N_20134,N_22424);
nand U23819 (N_23819,N_22037,N_20702);
xnor U23820 (N_23820,N_20338,N_22242);
or U23821 (N_23821,N_21833,N_20295);
or U23822 (N_23822,N_22270,N_22006);
nand U23823 (N_23823,N_21019,N_21862);
nand U23824 (N_23824,N_21143,N_20733);
nor U23825 (N_23825,N_20107,N_21971);
or U23826 (N_23826,N_20846,N_21191);
nand U23827 (N_23827,N_21703,N_21545);
or U23828 (N_23828,N_21813,N_20939);
and U23829 (N_23829,N_22468,N_20754);
nor U23830 (N_23830,N_21500,N_22174);
xnor U23831 (N_23831,N_20981,N_22240);
and U23832 (N_23832,N_20793,N_21235);
and U23833 (N_23833,N_20462,N_20626);
nor U23834 (N_23834,N_21943,N_21012);
nand U23835 (N_23835,N_21887,N_21502);
nor U23836 (N_23836,N_20040,N_21183);
xor U23837 (N_23837,N_20116,N_21081);
nor U23838 (N_23838,N_20153,N_20877);
xor U23839 (N_23839,N_21166,N_22353);
nor U23840 (N_23840,N_20226,N_21260);
xor U23841 (N_23841,N_20115,N_20116);
nand U23842 (N_23842,N_22456,N_22144);
xor U23843 (N_23843,N_20672,N_22289);
or U23844 (N_23844,N_20198,N_22345);
or U23845 (N_23845,N_22298,N_22049);
xor U23846 (N_23846,N_21098,N_22422);
xor U23847 (N_23847,N_22208,N_20777);
nand U23848 (N_23848,N_21472,N_22438);
nor U23849 (N_23849,N_22011,N_21428);
and U23850 (N_23850,N_22457,N_21328);
xnor U23851 (N_23851,N_20796,N_20184);
and U23852 (N_23852,N_20412,N_22497);
nand U23853 (N_23853,N_21972,N_20013);
nor U23854 (N_23854,N_21423,N_21151);
nand U23855 (N_23855,N_21253,N_21925);
nand U23856 (N_23856,N_20750,N_20761);
nand U23857 (N_23857,N_22096,N_21062);
xnor U23858 (N_23858,N_20389,N_21204);
nor U23859 (N_23859,N_20753,N_22140);
or U23860 (N_23860,N_21204,N_20045);
nor U23861 (N_23861,N_21370,N_21218);
xnor U23862 (N_23862,N_20314,N_21174);
nand U23863 (N_23863,N_21664,N_20572);
and U23864 (N_23864,N_20177,N_21809);
or U23865 (N_23865,N_20885,N_21133);
xor U23866 (N_23866,N_22124,N_22172);
nand U23867 (N_23867,N_20785,N_22153);
nand U23868 (N_23868,N_20143,N_21636);
nor U23869 (N_23869,N_20221,N_22198);
nor U23870 (N_23870,N_20163,N_22365);
and U23871 (N_23871,N_21830,N_20946);
and U23872 (N_23872,N_22339,N_20491);
or U23873 (N_23873,N_21356,N_20867);
xnor U23874 (N_23874,N_22251,N_22391);
and U23875 (N_23875,N_22147,N_20744);
xor U23876 (N_23876,N_20705,N_20416);
nor U23877 (N_23877,N_21872,N_22481);
xnor U23878 (N_23878,N_20543,N_22038);
xnor U23879 (N_23879,N_22131,N_20437);
or U23880 (N_23880,N_20741,N_20979);
xnor U23881 (N_23881,N_21419,N_22259);
xor U23882 (N_23882,N_20961,N_21399);
and U23883 (N_23883,N_20840,N_22118);
and U23884 (N_23884,N_22091,N_20784);
xor U23885 (N_23885,N_21044,N_21331);
or U23886 (N_23886,N_21530,N_20694);
xnor U23887 (N_23887,N_20357,N_21401);
or U23888 (N_23888,N_21311,N_20300);
and U23889 (N_23889,N_22084,N_21524);
nor U23890 (N_23890,N_22461,N_20281);
nand U23891 (N_23891,N_21412,N_22103);
nor U23892 (N_23892,N_21829,N_22167);
nand U23893 (N_23893,N_21787,N_22144);
nor U23894 (N_23894,N_22427,N_21336);
and U23895 (N_23895,N_22146,N_22173);
nor U23896 (N_23896,N_20621,N_20239);
and U23897 (N_23897,N_21344,N_22179);
nand U23898 (N_23898,N_20015,N_21436);
nand U23899 (N_23899,N_20827,N_22156);
xor U23900 (N_23900,N_21343,N_21574);
or U23901 (N_23901,N_20270,N_22039);
nand U23902 (N_23902,N_22410,N_21696);
nor U23903 (N_23903,N_21908,N_22000);
or U23904 (N_23904,N_21256,N_22383);
or U23905 (N_23905,N_21294,N_22024);
and U23906 (N_23906,N_20713,N_22076);
nand U23907 (N_23907,N_21231,N_21004);
or U23908 (N_23908,N_22238,N_20336);
nor U23909 (N_23909,N_21115,N_20024);
or U23910 (N_23910,N_20600,N_22472);
nor U23911 (N_23911,N_20198,N_20764);
and U23912 (N_23912,N_22089,N_21811);
or U23913 (N_23913,N_20321,N_22276);
nor U23914 (N_23914,N_21869,N_22184);
and U23915 (N_23915,N_21331,N_21335);
xor U23916 (N_23916,N_22366,N_20440);
nor U23917 (N_23917,N_20906,N_22280);
xnor U23918 (N_23918,N_20960,N_21581);
nand U23919 (N_23919,N_21471,N_20559);
nand U23920 (N_23920,N_21131,N_21249);
nor U23921 (N_23921,N_20152,N_20900);
or U23922 (N_23922,N_20177,N_20183);
or U23923 (N_23923,N_22391,N_21095);
nor U23924 (N_23924,N_20007,N_21816);
xnor U23925 (N_23925,N_21818,N_20287);
and U23926 (N_23926,N_21577,N_20854);
nor U23927 (N_23927,N_20875,N_20623);
nand U23928 (N_23928,N_21135,N_20847);
xor U23929 (N_23929,N_20166,N_21837);
or U23930 (N_23930,N_20299,N_21484);
and U23931 (N_23931,N_21621,N_21060);
nor U23932 (N_23932,N_21103,N_22368);
nor U23933 (N_23933,N_21107,N_21325);
and U23934 (N_23934,N_21035,N_22348);
or U23935 (N_23935,N_21400,N_21931);
or U23936 (N_23936,N_22434,N_21375);
or U23937 (N_23937,N_20815,N_22002);
and U23938 (N_23938,N_20707,N_21043);
and U23939 (N_23939,N_21360,N_20434);
nand U23940 (N_23940,N_22466,N_22279);
nand U23941 (N_23941,N_21520,N_22255);
and U23942 (N_23942,N_21416,N_22368);
xor U23943 (N_23943,N_20295,N_20020);
or U23944 (N_23944,N_20360,N_21091);
nand U23945 (N_23945,N_21942,N_21240);
and U23946 (N_23946,N_20900,N_22144);
nand U23947 (N_23947,N_20884,N_21378);
nand U23948 (N_23948,N_20178,N_21375);
nand U23949 (N_23949,N_20688,N_21060);
or U23950 (N_23950,N_22023,N_22099);
xor U23951 (N_23951,N_21099,N_21448);
or U23952 (N_23952,N_21781,N_21517);
and U23953 (N_23953,N_22099,N_21156);
nand U23954 (N_23954,N_21231,N_21386);
nor U23955 (N_23955,N_21299,N_21373);
xor U23956 (N_23956,N_22265,N_20270);
and U23957 (N_23957,N_20017,N_21407);
or U23958 (N_23958,N_20750,N_20337);
xnor U23959 (N_23959,N_21196,N_22259);
and U23960 (N_23960,N_20092,N_21180);
nand U23961 (N_23961,N_22227,N_21323);
or U23962 (N_23962,N_20551,N_21167);
and U23963 (N_23963,N_21975,N_22373);
or U23964 (N_23964,N_20321,N_20027);
nand U23965 (N_23965,N_22490,N_22409);
and U23966 (N_23966,N_22284,N_20614);
and U23967 (N_23967,N_20248,N_21642);
xnor U23968 (N_23968,N_20273,N_22480);
and U23969 (N_23969,N_21150,N_21422);
xor U23970 (N_23970,N_21020,N_20208);
xor U23971 (N_23971,N_22454,N_22323);
nand U23972 (N_23972,N_20666,N_21710);
nand U23973 (N_23973,N_21427,N_20904);
and U23974 (N_23974,N_21744,N_21189);
nor U23975 (N_23975,N_20790,N_20304);
and U23976 (N_23976,N_20643,N_22117);
nand U23977 (N_23977,N_21772,N_22140);
nor U23978 (N_23978,N_21051,N_21612);
or U23979 (N_23979,N_21031,N_21981);
xor U23980 (N_23980,N_20448,N_20224);
nand U23981 (N_23981,N_20150,N_21819);
or U23982 (N_23982,N_22049,N_21589);
or U23983 (N_23983,N_22031,N_21029);
nor U23984 (N_23984,N_21579,N_20425);
xor U23985 (N_23985,N_21929,N_20351);
nor U23986 (N_23986,N_21447,N_21569);
and U23987 (N_23987,N_21268,N_21042);
xor U23988 (N_23988,N_22410,N_20057);
nor U23989 (N_23989,N_21467,N_21446);
nand U23990 (N_23990,N_20541,N_21234);
nand U23991 (N_23991,N_21424,N_21869);
and U23992 (N_23992,N_22494,N_20329);
or U23993 (N_23993,N_20844,N_21059);
and U23994 (N_23994,N_20242,N_21976);
xor U23995 (N_23995,N_21966,N_20642);
xnor U23996 (N_23996,N_22399,N_21697);
xnor U23997 (N_23997,N_21222,N_21752);
nor U23998 (N_23998,N_21879,N_22175);
or U23999 (N_23999,N_21564,N_20543);
xor U24000 (N_24000,N_20826,N_20547);
nor U24001 (N_24001,N_21508,N_21638);
xor U24002 (N_24002,N_22454,N_21727);
nor U24003 (N_24003,N_20224,N_22041);
xnor U24004 (N_24004,N_20170,N_21266);
xor U24005 (N_24005,N_20415,N_21542);
or U24006 (N_24006,N_22180,N_21686);
nand U24007 (N_24007,N_21497,N_20642);
and U24008 (N_24008,N_22375,N_20441);
nor U24009 (N_24009,N_20382,N_21540);
and U24010 (N_24010,N_22394,N_21091);
and U24011 (N_24011,N_21624,N_21766);
nor U24012 (N_24012,N_21914,N_21203);
nand U24013 (N_24013,N_22110,N_22244);
nand U24014 (N_24014,N_20756,N_21419);
or U24015 (N_24015,N_21895,N_22148);
or U24016 (N_24016,N_20757,N_20807);
nand U24017 (N_24017,N_21728,N_20984);
and U24018 (N_24018,N_21703,N_21878);
nor U24019 (N_24019,N_21129,N_20529);
nor U24020 (N_24020,N_20197,N_21799);
nand U24021 (N_24021,N_22427,N_20246);
xnor U24022 (N_24022,N_20335,N_21089);
nand U24023 (N_24023,N_20153,N_20559);
xor U24024 (N_24024,N_20191,N_20436);
or U24025 (N_24025,N_20362,N_22267);
and U24026 (N_24026,N_20148,N_21356);
or U24027 (N_24027,N_20617,N_21575);
xnor U24028 (N_24028,N_21976,N_22085);
or U24029 (N_24029,N_20512,N_22161);
xnor U24030 (N_24030,N_22118,N_22473);
nor U24031 (N_24031,N_20650,N_20110);
nand U24032 (N_24032,N_21108,N_20531);
nand U24033 (N_24033,N_22139,N_22234);
nand U24034 (N_24034,N_20700,N_20825);
nor U24035 (N_24035,N_20397,N_21611);
xor U24036 (N_24036,N_20784,N_20786);
xor U24037 (N_24037,N_21281,N_22184);
nand U24038 (N_24038,N_20058,N_20157);
nand U24039 (N_24039,N_21459,N_20542);
xor U24040 (N_24040,N_22109,N_20613);
or U24041 (N_24041,N_20353,N_21235);
nor U24042 (N_24042,N_20795,N_22257);
nor U24043 (N_24043,N_20708,N_22359);
nor U24044 (N_24044,N_20337,N_21638);
nor U24045 (N_24045,N_20008,N_21320);
or U24046 (N_24046,N_22042,N_22340);
or U24047 (N_24047,N_21624,N_21587);
xnor U24048 (N_24048,N_21408,N_20576);
nand U24049 (N_24049,N_20962,N_21064);
nand U24050 (N_24050,N_20332,N_20263);
or U24051 (N_24051,N_21821,N_22043);
nor U24052 (N_24052,N_20030,N_22442);
or U24053 (N_24053,N_21906,N_20574);
and U24054 (N_24054,N_20016,N_20755);
or U24055 (N_24055,N_20364,N_21699);
nand U24056 (N_24056,N_20812,N_20341);
nor U24057 (N_24057,N_21732,N_20611);
and U24058 (N_24058,N_22167,N_22185);
or U24059 (N_24059,N_20250,N_21132);
and U24060 (N_24060,N_21238,N_20088);
or U24061 (N_24061,N_21066,N_20508);
or U24062 (N_24062,N_20885,N_21059);
nand U24063 (N_24063,N_20776,N_21511);
xnor U24064 (N_24064,N_21755,N_21463);
or U24065 (N_24065,N_20828,N_21911);
or U24066 (N_24066,N_20484,N_20899);
nor U24067 (N_24067,N_20184,N_20855);
and U24068 (N_24068,N_20755,N_22333);
or U24069 (N_24069,N_22101,N_20072);
or U24070 (N_24070,N_21859,N_20293);
nor U24071 (N_24071,N_21019,N_22236);
xnor U24072 (N_24072,N_20166,N_21437);
and U24073 (N_24073,N_20390,N_20982);
and U24074 (N_24074,N_21124,N_20956);
xnor U24075 (N_24075,N_22045,N_21877);
and U24076 (N_24076,N_20393,N_21529);
xnor U24077 (N_24077,N_21222,N_21158);
xor U24078 (N_24078,N_20056,N_21757);
xor U24079 (N_24079,N_21171,N_22313);
and U24080 (N_24080,N_21192,N_21338);
or U24081 (N_24081,N_20982,N_22030);
xor U24082 (N_24082,N_20114,N_21463);
xor U24083 (N_24083,N_21260,N_20320);
and U24084 (N_24084,N_20694,N_20045);
and U24085 (N_24085,N_20225,N_21798);
xnor U24086 (N_24086,N_21547,N_21249);
xor U24087 (N_24087,N_20766,N_20885);
nor U24088 (N_24088,N_21425,N_21156);
xnor U24089 (N_24089,N_20836,N_20978);
xnor U24090 (N_24090,N_21742,N_20638);
nor U24091 (N_24091,N_22388,N_22106);
and U24092 (N_24092,N_22072,N_22477);
xnor U24093 (N_24093,N_20489,N_22054);
or U24094 (N_24094,N_20237,N_21234);
nand U24095 (N_24095,N_21170,N_20557);
nor U24096 (N_24096,N_20152,N_22167);
xor U24097 (N_24097,N_21285,N_21761);
nand U24098 (N_24098,N_22364,N_21242);
and U24099 (N_24099,N_20658,N_22075);
nand U24100 (N_24100,N_22084,N_20001);
and U24101 (N_24101,N_22437,N_20607);
nand U24102 (N_24102,N_22106,N_21434);
or U24103 (N_24103,N_20725,N_20236);
nand U24104 (N_24104,N_21620,N_20404);
xor U24105 (N_24105,N_21153,N_22443);
nand U24106 (N_24106,N_21799,N_20483);
xor U24107 (N_24107,N_22162,N_20658);
and U24108 (N_24108,N_20874,N_21115);
or U24109 (N_24109,N_20455,N_20387);
and U24110 (N_24110,N_21915,N_20471);
xor U24111 (N_24111,N_22071,N_20087);
or U24112 (N_24112,N_20798,N_21130);
or U24113 (N_24113,N_20631,N_20817);
nand U24114 (N_24114,N_22464,N_22403);
and U24115 (N_24115,N_21658,N_22203);
nand U24116 (N_24116,N_20090,N_21508);
and U24117 (N_24117,N_21907,N_20189);
nand U24118 (N_24118,N_22105,N_22166);
nand U24119 (N_24119,N_20747,N_21667);
and U24120 (N_24120,N_20265,N_21300);
nand U24121 (N_24121,N_21239,N_21974);
and U24122 (N_24122,N_21292,N_22116);
or U24123 (N_24123,N_20214,N_20217);
nand U24124 (N_24124,N_21921,N_21780);
xnor U24125 (N_24125,N_22304,N_21217);
nand U24126 (N_24126,N_21042,N_21152);
or U24127 (N_24127,N_20860,N_20000);
or U24128 (N_24128,N_20769,N_22023);
xor U24129 (N_24129,N_21143,N_22292);
nor U24130 (N_24130,N_22394,N_20258);
nand U24131 (N_24131,N_22443,N_21458);
xor U24132 (N_24132,N_20830,N_22117);
nand U24133 (N_24133,N_21387,N_21852);
nand U24134 (N_24134,N_22145,N_21704);
and U24135 (N_24135,N_20928,N_21140);
or U24136 (N_24136,N_20530,N_22417);
nor U24137 (N_24137,N_21205,N_21773);
xnor U24138 (N_24138,N_21371,N_20329);
nor U24139 (N_24139,N_21311,N_21227);
nand U24140 (N_24140,N_20372,N_22272);
or U24141 (N_24141,N_21499,N_21971);
nand U24142 (N_24142,N_20480,N_20536);
or U24143 (N_24143,N_20416,N_20208);
xor U24144 (N_24144,N_21287,N_21703);
and U24145 (N_24145,N_20133,N_20789);
and U24146 (N_24146,N_20728,N_21260);
xnor U24147 (N_24147,N_20168,N_20454);
xnor U24148 (N_24148,N_20963,N_21291);
and U24149 (N_24149,N_21753,N_20325);
nor U24150 (N_24150,N_20795,N_21315);
xor U24151 (N_24151,N_22079,N_20255);
nor U24152 (N_24152,N_22059,N_22050);
xor U24153 (N_24153,N_21342,N_21238);
xor U24154 (N_24154,N_21782,N_20980);
xnor U24155 (N_24155,N_20749,N_20998);
nor U24156 (N_24156,N_22033,N_22085);
and U24157 (N_24157,N_20491,N_22341);
nor U24158 (N_24158,N_21517,N_21554);
nor U24159 (N_24159,N_21996,N_20349);
xnor U24160 (N_24160,N_20570,N_21383);
or U24161 (N_24161,N_21748,N_20017);
nand U24162 (N_24162,N_21838,N_21678);
and U24163 (N_24163,N_20654,N_20634);
and U24164 (N_24164,N_21843,N_20297);
nor U24165 (N_24165,N_22213,N_22319);
and U24166 (N_24166,N_20887,N_21633);
nor U24167 (N_24167,N_22480,N_20207);
and U24168 (N_24168,N_22281,N_21341);
and U24169 (N_24169,N_22372,N_21579);
xnor U24170 (N_24170,N_20194,N_21666);
nor U24171 (N_24171,N_22168,N_20802);
nand U24172 (N_24172,N_22038,N_21506);
nand U24173 (N_24173,N_20206,N_21799);
or U24174 (N_24174,N_21763,N_21551);
nor U24175 (N_24175,N_22435,N_20674);
nor U24176 (N_24176,N_20659,N_20164);
nor U24177 (N_24177,N_20088,N_20988);
nand U24178 (N_24178,N_20389,N_21769);
and U24179 (N_24179,N_21300,N_21241);
xnor U24180 (N_24180,N_20397,N_21188);
or U24181 (N_24181,N_20129,N_21892);
nand U24182 (N_24182,N_22328,N_21450);
and U24183 (N_24183,N_20142,N_20781);
and U24184 (N_24184,N_22389,N_22326);
nand U24185 (N_24185,N_22230,N_22081);
nor U24186 (N_24186,N_20654,N_21085);
xor U24187 (N_24187,N_22322,N_21514);
and U24188 (N_24188,N_20908,N_21169);
nand U24189 (N_24189,N_20935,N_22487);
xor U24190 (N_24190,N_21444,N_20874);
nor U24191 (N_24191,N_20768,N_21775);
xor U24192 (N_24192,N_20434,N_21596);
nand U24193 (N_24193,N_21140,N_20690);
nor U24194 (N_24194,N_21714,N_20538);
and U24195 (N_24195,N_22387,N_21301);
nand U24196 (N_24196,N_20490,N_20477);
or U24197 (N_24197,N_21039,N_20874);
or U24198 (N_24198,N_20114,N_20790);
and U24199 (N_24199,N_20662,N_21375);
xor U24200 (N_24200,N_20695,N_20282);
nor U24201 (N_24201,N_21882,N_21176);
and U24202 (N_24202,N_22473,N_21944);
or U24203 (N_24203,N_20740,N_22069);
or U24204 (N_24204,N_21713,N_20987);
xor U24205 (N_24205,N_22173,N_21674);
nand U24206 (N_24206,N_21598,N_21730);
or U24207 (N_24207,N_21013,N_21152);
xor U24208 (N_24208,N_21260,N_22309);
nor U24209 (N_24209,N_22042,N_21912);
nor U24210 (N_24210,N_22243,N_20290);
or U24211 (N_24211,N_20736,N_20967);
xor U24212 (N_24212,N_21311,N_21254);
and U24213 (N_24213,N_21718,N_20357);
or U24214 (N_24214,N_20331,N_21039);
xnor U24215 (N_24215,N_20507,N_21292);
and U24216 (N_24216,N_21041,N_20145);
nor U24217 (N_24217,N_21790,N_22170);
nand U24218 (N_24218,N_20810,N_22000);
or U24219 (N_24219,N_21963,N_20585);
and U24220 (N_24220,N_21131,N_20648);
xor U24221 (N_24221,N_20266,N_21022);
and U24222 (N_24222,N_21552,N_21976);
nand U24223 (N_24223,N_20305,N_20637);
nor U24224 (N_24224,N_22054,N_22150);
nor U24225 (N_24225,N_20331,N_20874);
and U24226 (N_24226,N_21005,N_20287);
nand U24227 (N_24227,N_21930,N_21323);
xnor U24228 (N_24228,N_20364,N_20310);
or U24229 (N_24229,N_22240,N_20481);
xor U24230 (N_24230,N_21065,N_20947);
xnor U24231 (N_24231,N_21678,N_20896);
nor U24232 (N_24232,N_21916,N_21249);
and U24233 (N_24233,N_20564,N_22447);
nor U24234 (N_24234,N_21270,N_22260);
and U24235 (N_24235,N_22474,N_21677);
nor U24236 (N_24236,N_21928,N_20752);
and U24237 (N_24237,N_21778,N_20695);
and U24238 (N_24238,N_21617,N_20103);
xor U24239 (N_24239,N_21358,N_22495);
nor U24240 (N_24240,N_20115,N_21765);
nor U24241 (N_24241,N_21366,N_21955);
nand U24242 (N_24242,N_20419,N_21289);
and U24243 (N_24243,N_20071,N_22415);
nor U24244 (N_24244,N_21899,N_22029);
xnor U24245 (N_24245,N_20978,N_22179);
nand U24246 (N_24246,N_21796,N_21272);
xnor U24247 (N_24247,N_20042,N_21570);
or U24248 (N_24248,N_21298,N_21175);
nor U24249 (N_24249,N_21938,N_20261);
nand U24250 (N_24250,N_22084,N_20952);
nand U24251 (N_24251,N_21316,N_20177);
nand U24252 (N_24252,N_21988,N_20286);
or U24253 (N_24253,N_21387,N_20919);
nand U24254 (N_24254,N_20168,N_21268);
nor U24255 (N_24255,N_20942,N_20777);
nand U24256 (N_24256,N_20721,N_22033);
and U24257 (N_24257,N_20813,N_20892);
or U24258 (N_24258,N_21113,N_20635);
or U24259 (N_24259,N_21730,N_21895);
nor U24260 (N_24260,N_22426,N_20519);
xor U24261 (N_24261,N_21657,N_20829);
xnor U24262 (N_24262,N_20915,N_21872);
nand U24263 (N_24263,N_22050,N_20259);
and U24264 (N_24264,N_21105,N_21317);
nor U24265 (N_24265,N_20673,N_22389);
and U24266 (N_24266,N_20358,N_21428);
nor U24267 (N_24267,N_20994,N_21752);
and U24268 (N_24268,N_21355,N_21210);
or U24269 (N_24269,N_20490,N_20942);
or U24270 (N_24270,N_22443,N_20630);
or U24271 (N_24271,N_20077,N_20320);
nor U24272 (N_24272,N_21979,N_20708);
or U24273 (N_24273,N_20366,N_20903);
or U24274 (N_24274,N_20422,N_21382);
nand U24275 (N_24275,N_22178,N_21349);
or U24276 (N_24276,N_22216,N_20270);
nor U24277 (N_24277,N_20805,N_22084);
nor U24278 (N_24278,N_21517,N_22186);
nand U24279 (N_24279,N_21367,N_21698);
xnor U24280 (N_24280,N_22125,N_20307);
nor U24281 (N_24281,N_20717,N_20803);
or U24282 (N_24282,N_20246,N_20471);
nor U24283 (N_24283,N_20017,N_21714);
nor U24284 (N_24284,N_20029,N_22141);
or U24285 (N_24285,N_21179,N_21754);
xnor U24286 (N_24286,N_20514,N_22136);
or U24287 (N_24287,N_21884,N_21556);
xnor U24288 (N_24288,N_21045,N_21984);
xnor U24289 (N_24289,N_21406,N_21823);
and U24290 (N_24290,N_20441,N_22251);
or U24291 (N_24291,N_21206,N_21652);
or U24292 (N_24292,N_20140,N_20131);
xnor U24293 (N_24293,N_20079,N_20250);
and U24294 (N_24294,N_20379,N_21460);
or U24295 (N_24295,N_21233,N_22465);
nor U24296 (N_24296,N_20865,N_20690);
and U24297 (N_24297,N_20233,N_21040);
nor U24298 (N_24298,N_20180,N_20409);
nor U24299 (N_24299,N_20613,N_20136);
and U24300 (N_24300,N_20979,N_20673);
nand U24301 (N_24301,N_20870,N_20016);
nor U24302 (N_24302,N_21792,N_21118);
and U24303 (N_24303,N_20261,N_20789);
and U24304 (N_24304,N_20584,N_20853);
nor U24305 (N_24305,N_21541,N_21188);
nand U24306 (N_24306,N_21100,N_22219);
xor U24307 (N_24307,N_22486,N_20462);
xor U24308 (N_24308,N_21912,N_22076);
or U24309 (N_24309,N_22394,N_22081);
and U24310 (N_24310,N_22495,N_20617);
and U24311 (N_24311,N_22329,N_21833);
or U24312 (N_24312,N_22180,N_21511);
or U24313 (N_24313,N_21271,N_20626);
nor U24314 (N_24314,N_21317,N_20834);
nand U24315 (N_24315,N_21999,N_20470);
or U24316 (N_24316,N_20019,N_21992);
or U24317 (N_24317,N_22152,N_21334);
nor U24318 (N_24318,N_22386,N_20693);
nand U24319 (N_24319,N_21400,N_21052);
xnor U24320 (N_24320,N_20310,N_22335);
nor U24321 (N_24321,N_20328,N_21734);
nor U24322 (N_24322,N_20592,N_22299);
and U24323 (N_24323,N_20478,N_21353);
nand U24324 (N_24324,N_21235,N_20996);
or U24325 (N_24325,N_21354,N_20026);
nand U24326 (N_24326,N_21736,N_22492);
xnor U24327 (N_24327,N_21440,N_20139);
xnor U24328 (N_24328,N_22480,N_21987);
or U24329 (N_24329,N_20639,N_22149);
nor U24330 (N_24330,N_21014,N_21354);
and U24331 (N_24331,N_20890,N_20653);
or U24332 (N_24332,N_20125,N_21216);
xor U24333 (N_24333,N_22377,N_20268);
or U24334 (N_24334,N_21120,N_21584);
nor U24335 (N_24335,N_20027,N_20193);
and U24336 (N_24336,N_21721,N_21350);
nand U24337 (N_24337,N_21960,N_21789);
xor U24338 (N_24338,N_20248,N_22137);
xor U24339 (N_24339,N_20219,N_21528);
nor U24340 (N_24340,N_20857,N_20383);
or U24341 (N_24341,N_20725,N_20832);
and U24342 (N_24342,N_21373,N_20986);
nand U24343 (N_24343,N_21319,N_22220);
nor U24344 (N_24344,N_21852,N_22323);
and U24345 (N_24345,N_20684,N_21191);
and U24346 (N_24346,N_21504,N_22187);
or U24347 (N_24347,N_21355,N_20334);
and U24348 (N_24348,N_20903,N_20362);
xor U24349 (N_24349,N_20034,N_21773);
or U24350 (N_24350,N_21424,N_22263);
xnor U24351 (N_24351,N_21029,N_21375);
xnor U24352 (N_24352,N_20864,N_21197);
nor U24353 (N_24353,N_21743,N_22326);
or U24354 (N_24354,N_21746,N_22352);
and U24355 (N_24355,N_21571,N_21309);
xor U24356 (N_24356,N_20231,N_21750);
and U24357 (N_24357,N_20283,N_20559);
and U24358 (N_24358,N_21240,N_21366);
nor U24359 (N_24359,N_21507,N_22177);
xnor U24360 (N_24360,N_21194,N_20652);
nor U24361 (N_24361,N_20546,N_21192);
or U24362 (N_24362,N_22205,N_21250);
xor U24363 (N_24363,N_22124,N_20548);
and U24364 (N_24364,N_21440,N_21140);
nor U24365 (N_24365,N_22446,N_21685);
and U24366 (N_24366,N_20250,N_22027);
nand U24367 (N_24367,N_22088,N_22273);
xnor U24368 (N_24368,N_22057,N_21511);
nand U24369 (N_24369,N_21015,N_20196);
xor U24370 (N_24370,N_20928,N_22486);
nor U24371 (N_24371,N_21231,N_20707);
and U24372 (N_24372,N_20943,N_21977);
or U24373 (N_24373,N_21965,N_21050);
or U24374 (N_24374,N_20451,N_20800);
and U24375 (N_24375,N_20336,N_21150);
or U24376 (N_24376,N_22388,N_21206);
xor U24377 (N_24377,N_21508,N_21469);
nor U24378 (N_24378,N_21138,N_21283);
nor U24379 (N_24379,N_22423,N_20763);
nor U24380 (N_24380,N_21425,N_21909);
or U24381 (N_24381,N_20432,N_20035);
xor U24382 (N_24382,N_20020,N_22281);
or U24383 (N_24383,N_21731,N_22118);
nor U24384 (N_24384,N_20007,N_20473);
nand U24385 (N_24385,N_21108,N_21773);
nand U24386 (N_24386,N_20698,N_21604);
nand U24387 (N_24387,N_20986,N_20787);
xnor U24388 (N_24388,N_20178,N_22243);
nand U24389 (N_24389,N_21865,N_22385);
or U24390 (N_24390,N_21138,N_22193);
xor U24391 (N_24391,N_20363,N_21867);
xor U24392 (N_24392,N_21122,N_22096);
nand U24393 (N_24393,N_21365,N_20712);
nand U24394 (N_24394,N_20450,N_20518);
and U24395 (N_24395,N_21385,N_21181);
nand U24396 (N_24396,N_22422,N_20913);
or U24397 (N_24397,N_21630,N_21485);
or U24398 (N_24398,N_20100,N_21905);
nand U24399 (N_24399,N_21322,N_22259);
nand U24400 (N_24400,N_20386,N_20364);
and U24401 (N_24401,N_21433,N_22020);
or U24402 (N_24402,N_20402,N_20514);
xor U24403 (N_24403,N_22020,N_20594);
xor U24404 (N_24404,N_20042,N_20388);
nor U24405 (N_24405,N_21842,N_20047);
xnor U24406 (N_24406,N_21618,N_22161);
xor U24407 (N_24407,N_21727,N_21014);
xor U24408 (N_24408,N_20633,N_20761);
nor U24409 (N_24409,N_22382,N_21499);
and U24410 (N_24410,N_21661,N_22416);
xor U24411 (N_24411,N_21390,N_21748);
xor U24412 (N_24412,N_21608,N_20094);
and U24413 (N_24413,N_22048,N_21732);
nand U24414 (N_24414,N_22291,N_20034);
nand U24415 (N_24415,N_20106,N_20120);
nand U24416 (N_24416,N_21497,N_20463);
nand U24417 (N_24417,N_21480,N_21985);
nand U24418 (N_24418,N_20665,N_21171);
and U24419 (N_24419,N_20715,N_20012);
xnor U24420 (N_24420,N_21584,N_21951);
or U24421 (N_24421,N_22078,N_20016);
xnor U24422 (N_24422,N_21848,N_20467);
nor U24423 (N_24423,N_22077,N_20221);
or U24424 (N_24424,N_21414,N_22159);
nand U24425 (N_24425,N_22386,N_20711);
nand U24426 (N_24426,N_20650,N_20898);
nor U24427 (N_24427,N_21335,N_20165);
or U24428 (N_24428,N_21225,N_22454);
xnor U24429 (N_24429,N_20391,N_21836);
nand U24430 (N_24430,N_20959,N_21684);
nor U24431 (N_24431,N_20672,N_21808);
or U24432 (N_24432,N_21354,N_20904);
xor U24433 (N_24433,N_20771,N_20396);
or U24434 (N_24434,N_22255,N_21693);
xor U24435 (N_24435,N_20250,N_21682);
xor U24436 (N_24436,N_20521,N_20073);
nand U24437 (N_24437,N_22030,N_21791);
nor U24438 (N_24438,N_20908,N_21500);
xnor U24439 (N_24439,N_20760,N_22293);
or U24440 (N_24440,N_20749,N_21513);
nand U24441 (N_24441,N_22139,N_20367);
or U24442 (N_24442,N_22466,N_21155);
xor U24443 (N_24443,N_20016,N_22459);
or U24444 (N_24444,N_20718,N_21875);
or U24445 (N_24445,N_20112,N_22485);
nor U24446 (N_24446,N_20680,N_21029);
nand U24447 (N_24447,N_20027,N_21752);
nand U24448 (N_24448,N_21803,N_21406);
nor U24449 (N_24449,N_22062,N_22098);
nor U24450 (N_24450,N_21880,N_20804);
xor U24451 (N_24451,N_22020,N_21894);
xor U24452 (N_24452,N_20865,N_20234);
nor U24453 (N_24453,N_20362,N_21617);
nor U24454 (N_24454,N_21740,N_20400);
nand U24455 (N_24455,N_22458,N_21491);
nor U24456 (N_24456,N_21742,N_21843);
nor U24457 (N_24457,N_22384,N_20681);
or U24458 (N_24458,N_21190,N_22031);
nor U24459 (N_24459,N_21386,N_21270);
nor U24460 (N_24460,N_21451,N_21935);
nand U24461 (N_24461,N_21087,N_20132);
and U24462 (N_24462,N_21314,N_21310);
nand U24463 (N_24463,N_20602,N_22311);
xor U24464 (N_24464,N_21931,N_20967);
nor U24465 (N_24465,N_22092,N_20239);
xor U24466 (N_24466,N_22421,N_20765);
nor U24467 (N_24467,N_22211,N_20262);
and U24468 (N_24468,N_21722,N_20297);
nand U24469 (N_24469,N_20100,N_21251);
nand U24470 (N_24470,N_21391,N_20218);
nand U24471 (N_24471,N_22160,N_20457);
and U24472 (N_24472,N_20040,N_20832);
nand U24473 (N_24473,N_21240,N_20671);
nor U24474 (N_24474,N_20873,N_20133);
and U24475 (N_24475,N_20582,N_21874);
or U24476 (N_24476,N_20173,N_22127);
xor U24477 (N_24477,N_22016,N_20856);
nor U24478 (N_24478,N_21388,N_20345);
nand U24479 (N_24479,N_22228,N_21630);
and U24480 (N_24480,N_20535,N_20695);
nand U24481 (N_24481,N_22477,N_20543);
and U24482 (N_24482,N_20605,N_21311);
nor U24483 (N_24483,N_20559,N_20476);
nand U24484 (N_24484,N_20245,N_20195);
or U24485 (N_24485,N_21438,N_21252);
and U24486 (N_24486,N_21892,N_21343);
nand U24487 (N_24487,N_21665,N_20005);
nand U24488 (N_24488,N_20805,N_22013);
nand U24489 (N_24489,N_22232,N_21627);
xnor U24490 (N_24490,N_21279,N_20316);
xor U24491 (N_24491,N_21568,N_20793);
or U24492 (N_24492,N_22383,N_20514);
nor U24493 (N_24493,N_20706,N_21585);
nand U24494 (N_24494,N_20384,N_21016);
or U24495 (N_24495,N_20026,N_21086);
nor U24496 (N_24496,N_22292,N_22040);
and U24497 (N_24497,N_21146,N_21529);
nor U24498 (N_24498,N_21979,N_21430);
xor U24499 (N_24499,N_21551,N_21480);
nor U24500 (N_24500,N_20598,N_21358);
xor U24501 (N_24501,N_20162,N_22079);
xnor U24502 (N_24502,N_22455,N_20886);
or U24503 (N_24503,N_20221,N_21008);
or U24504 (N_24504,N_21326,N_20201);
and U24505 (N_24505,N_21272,N_22415);
and U24506 (N_24506,N_21174,N_22256);
nand U24507 (N_24507,N_21595,N_22375);
nor U24508 (N_24508,N_21241,N_21467);
xor U24509 (N_24509,N_20712,N_20926);
and U24510 (N_24510,N_22117,N_21523);
or U24511 (N_24511,N_21530,N_20168);
xor U24512 (N_24512,N_20505,N_20260);
nand U24513 (N_24513,N_21978,N_21422);
and U24514 (N_24514,N_20977,N_21682);
nor U24515 (N_24515,N_21332,N_20651);
nor U24516 (N_24516,N_22280,N_20283);
nand U24517 (N_24517,N_21835,N_21962);
or U24518 (N_24518,N_22356,N_21870);
or U24519 (N_24519,N_21968,N_22285);
xnor U24520 (N_24520,N_21650,N_20505);
or U24521 (N_24521,N_20658,N_20854);
xnor U24522 (N_24522,N_21059,N_21349);
or U24523 (N_24523,N_22462,N_21837);
or U24524 (N_24524,N_21881,N_20806);
xnor U24525 (N_24525,N_20169,N_22413);
or U24526 (N_24526,N_20033,N_20472);
nand U24527 (N_24527,N_20032,N_20622);
or U24528 (N_24528,N_21880,N_20253);
xnor U24529 (N_24529,N_22053,N_20848);
nand U24530 (N_24530,N_20616,N_22498);
xnor U24531 (N_24531,N_21893,N_20286);
xnor U24532 (N_24532,N_20737,N_22304);
and U24533 (N_24533,N_21727,N_22170);
nor U24534 (N_24534,N_20176,N_20011);
xor U24535 (N_24535,N_22287,N_21399);
and U24536 (N_24536,N_20383,N_20370);
xor U24537 (N_24537,N_21271,N_22404);
nand U24538 (N_24538,N_20539,N_21712);
or U24539 (N_24539,N_21267,N_20432);
nor U24540 (N_24540,N_21623,N_20836);
xnor U24541 (N_24541,N_22316,N_21296);
xor U24542 (N_24542,N_20419,N_21810);
nor U24543 (N_24543,N_21123,N_20857);
nand U24544 (N_24544,N_20858,N_22216);
or U24545 (N_24545,N_20228,N_20749);
nand U24546 (N_24546,N_20549,N_20189);
nor U24547 (N_24547,N_21611,N_21935);
or U24548 (N_24548,N_22222,N_20479);
xnor U24549 (N_24549,N_20866,N_22338);
or U24550 (N_24550,N_21158,N_20637);
xor U24551 (N_24551,N_21851,N_21291);
or U24552 (N_24552,N_21202,N_21374);
nand U24553 (N_24553,N_20020,N_21062);
nand U24554 (N_24554,N_21731,N_20680);
nand U24555 (N_24555,N_20474,N_21263);
and U24556 (N_24556,N_22171,N_22260);
or U24557 (N_24557,N_20087,N_20062);
nand U24558 (N_24558,N_21614,N_20889);
xor U24559 (N_24559,N_22138,N_21927);
xor U24560 (N_24560,N_21441,N_22410);
xnor U24561 (N_24561,N_22073,N_20793);
nand U24562 (N_24562,N_21890,N_22263);
and U24563 (N_24563,N_22333,N_22157);
and U24564 (N_24564,N_21252,N_21273);
xnor U24565 (N_24565,N_20076,N_20380);
nor U24566 (N_24566,N_21465,N_20623);
xnor U24567 (N_24567,N_20055,N_20932);
xnor U24568 (N_24568,N_21403,N_21745);
xnor U24569 (N_24569,N_20861,N_20769);
nor U24570 (N_24570,N_20551,N_21949);
xor U24571 (N_24571,N_21022,N_20539);
xnor U24572 (N_24572,N_21897,N_20185);
nor U24573 (N_24573,N_20878,N_21775);
xnor U24574 (N_24574,N_21959,N_22420);
or U24575 (N_24575,N_22385,N_20509);
xnor U24576 (N_24576,N_22224,N_20017);
nand U24577 (N_24577,N_22080,N_21715);
xnor U24578 (N_24578,N_21553,N_22009);
and U24579 (N_24579,N_22476,N_22044);
xor U24580 (N_24580,N_21409,N_20637);
or U24581 (N_24581,N_20003,N_21704);
nand U24582 (N_24582,N_20648,N_21623);
xnor U24583 (N_24583,N_21351,N_21083);
and U24584 (N_24584,N_22443,N_21678);
nand U24585 (N_24585,N_22099,N_21590);
xnor U24586 (N_24586,N_21046,N_22074);
xor U24587 (N_24587,N_20044,N_20170);
xnor U24588 (N_24588,N_21253,N_20283);
nor U24589 (N_24589,N_21035,N_20473);
xnor U24590 (N_24590,N_21133,N_21382);
nand U24591 (N_24591,N_20469,N_22081);
nand U24592 (N_24592,N_21050,N_20043);
or U24593 (N_24593,N_20780,N_21435);
nand U24594 (N_24594,N_20584,N_21315);
and U24595 (N_24595,N_20426,N_21669);
xor U24596 (N_24596,N_20802,N_21070);
nor U24597 (N_24597,N_20018,N_21061);
xor U24598 (N_24598,N_22398,N_22456);
nor U24599 (N_24599,N_21508,N_21804);
nor U24600 (N_24600,N_21100,N_22062);
xnor U24601 (N_24601,N_22089,N_20003);
xnor U24602 (N_24602,N_20718,N_20449);
nand U24603 (N_24603,N_21908,N_20828);
and U24604 (N_24604,N_21730,N_20189);
nor U24605 (N_24605,N_21624,N_21876);
nand U24606 (N_24606,N_21645,N_20821);
nand U24607 (N_24607,N_21160,N_22450);
and U24608 (N_24608,N_20181,N_20248);
nand U24609 (N_24609,N_21062,N_21604);
or U24610 (N_24610,N_21535,N_20595);
and U24611 (N_24611,N_21475,N_21200);
nor U24612 (N_24612,N_21049,N_22215);
xor U24613 (N_24613,N_20354,N_22492);
nand U24614 (N_24614,N_22333,N_22061);
or U24615 (N_24615,N_21612,N_21621);
nor U24616 (N_24616,N_22282,N_20767);
xor U24617 (N_24617,N_20736,N_21666);
nor U24618 (N_24618,N_20873,N_20725);
or U24619 (N_24619,N_21298,N_21075);
nor U24620 (N_24620,N_21317,N_20297);
xor U24621 (N_24621,N_21877,N_21677);
nor U24622 (N_24622,N_21405,N_21499);
nand U24623 (N_24623,N_21324,N_22405);
and U24624 (N_24624,N_21851,N_22234);
and U24625 (N_24625,N_20740,N_20716);
nor U24626 (N_24626,N_21826,N_21013);
and U24627 (N_24627,N_20907,N_20486);
xnor U24628 (N_24628,N_20255,N_22288);
nor U24629 (N_24629,N_20965,N_21621);
nand U24630 (N_24630,N_22337,N_20843);
nand U24631 (N_24631,N_21727,N_22325);
and U24632 (N_24632,N_21569,N_21075);
nand U24633 (N_24633,N_21284,N_20523);
nor U24634 (N_24634,N_21456,N_21972);
and U24635 (N_24635,N_20227,N_22076);
nor U24636 (N_24636,N_22014,N_20184);
nand U24637 (N_24637,N_20347,N_20490);
and U24638 (N_24638,N_20548,N_22239);
and U24639 (N_24639,N_20744,N_20494);
xnor U24640 (N_24640,N_21971,N_21724);
nor U24641 (N_24641,N_21046,N_20688);
and U24642 (N_24642,N_20618,N_20603);
and U24643 (N_24643,N_21600,N_20179);
and U24644 (N_24644,N_21964,N_22216);
and U24645 (N_24645,N_20070,N_20660);
xnor U24646 (N_24646,N_20229,N_20168);
nand U24647 (N_24647,N_21100,N_20910);
and U24648 (N_24648,N_21188,N_21364);
xnor U24649 (N_24649,N_20375,N_20533);
nor U24650 (N_24650,N_22261,N_20184);
nand U24651 (N_24651,N_20985,N_21309);
nor U24652 (N_24652,N_21153,N_21252);
nand U24653 (N_24653,N_21197,N_21182);
and U24654 (N_24654,N_20531,N_22276);
and U24655 (N_24655,N_20782,N_20024);
nor U24656 (N_24656,N_21209,N_21044);
xor U24657 (N_24657,N_20524,N_21881);
and U24658 (N_24658,N_22221,N_21965);
and U24659 (N_24659,N_21752,N_22228);
or U24660 (N_24660,N_20949,N_20832);
nor U24661 (N_24661,N_22212,N_22482);
or U24662 (N_24662,N_21261,N_21801);
and U24663 (N_24663,N_20780,N_20697);
nand U24664 (N_24664,N_20004,N_21564);
xor U24665 (N_24665,N_21486,N_21070);
and U24666 (N_24666,N_20121,N_21287);
and U24667 (N_24667,N_20668,N_22451);
xnor U24668 (N_24668,N_21825,N_20580);
xor U24669 (N_24669,N_21932,N_21976);
or U24670 (N_24670,N_20745,N_21631);
nand U24671 (N_24671,N_20848,N_20446);
and U24672 (N_24672,N_22071,N_21833);
and U24673 (N_24673,N_21844,N_21973);
xor U24674 (N_24674,N_21773,N_20287);
nand U24675 (N_24675,N_22403,N_20017);
xor U24676 (N_24676,N_21193,N_21993);
or U24677 (N_24677,N_20658,N_21849);
or U24678 (N_24678,N_20918,N_21350);
and U24679 (N_24679,N_21334,N_22090);
or U24680 (N_24680,N_21807,N_22485);
xnor U24681 (N_24681,N_22333,N_21772);
or U24682 (N_24682,N_20688,N_20697);
or U24683 (N_24683,N_21099,N_21353);
or U24684 (N_24684,N_21761,N_22309);
or U24685 (N_24685,N_21993,N_21022);
nor U24686 (N_24686,N_21029,N_22267);
xnor U24687 (N_24687,N_22339,N_21732);
xnor U24688 (N_24688,N_21842,N_21971);
or U24689 (N_24689,N_20700,N_21970);
nand U24690 (N_24690,N_22172,N_20832);
nor U24691 (N_24691,N_20558,N_20984);
or U24692 (N_24692,N_20184,N_21904);
nor U24693 (N_24693,N_21891,N_21710);
or U24694 (N_24694,N_20324,N_20929);
xnor U24695 (N_24695,N_22185,N_22171);
nor U24696 (N_24696,N_21889,N_21866);
xnor U24697 (N_24697,N_20539,N_20023);
or U24698 (N_24698,N_21244,N_22135);
or U24699 (N_24699,N_20547,N_20513);
or U24700 (N_24700,N_20452,N_21985);
nor U24701 (N_24701,N_21854,N_21755);
xor U24702 (N_24702,N_20491,N_21873);
xor U24703 (N_24703,N_21436,N_21491);
or U24704 (N_24704,N_21360,N_20821);
nand U24705 (N_24705,N_21333,N_22277);
nor U24706 (N_24706,N_20905,N_20497);
nor U24707 (N_24707,N_20199,N_20056);
and U24708 (N_24708,N_20854,N_21447);
nand U24709 (N_24709,N_22249,N_20422);
or U24710 (N_24710,N_20873,N_20403);
xnor U24711 (N_24711,N_21825,N_20015);
xnor U24712 (N_24712,N_22435,N_20172);
and U24713 (N_24713,N_21668,N_21180);
nand U24714 (N_24714,N_21197,N_21151);
nand U24715 (N_24715,N_20290,N_21866);
nor U24716 (N_24716,N_20582,N_22083);
xnor U24717 (N_24717,N_21937,N_20698);
or U24718 (N_24718,N_21763,N_20633);
xor U24719 (N_24719,N_21752,N_21536);
and U24720 (N_24720,N_22305,N_20913);
or U24721 (N_24721,N_21862,N_20201);
and U24722 (N_24722,N_20500,N_21254);
nand U24723 (N_24723,N_21163,N_20519);
and U24724 (N_24724,N_21670,N_20992);
xnor U24725 (N_24725,N_21157,N_21504);
xnor U24726 (N_24726,N_20110,N_22051);
xor U24727 (N_24727,N_20579,N_20858);
nand U24728 (N_24728,N_22211,N_22345);
xnor U24729 (N_24729,N_20935,N_20095);
or U24730 (N_24730,N_21176,N_21008);
or U24731 (N_24731,N_20974,N_21113);
xnor U24732 (N_24732,N_21859,N_20188);
and U24733 (N_24733,N_20937,N_22452);
or U24734 (N_24734,N_20068,N_20829);
or U24735 (N_24735,N_20741,N_20731);
and U24736 (N_24736,N_20164,N_21970);
nand U24737 (N_24737,N_22317,N_22027);
xnor U24738 (N_24738,N_20485,N_20456);
nand U24739 (N_24739,N_21322,N_21838);
xnor U24740 (N_24740,N_21762,N_20150);
nand U24741 (N_24741,N_21037,N_21985);
or U24742 (N_24742,N_21023,N_22325);
or U24743 (N_24743,N_21543,N_20862);
xnor U24744 (N_24744,N_20143,N_20223);
nor U24745 (N_24745,N_21991,N_20527);
nand U24746 (N_24746,N_22150,N_22225);
or U24747 (N_24747,N_20343,N_21102);
nor U24748 (N_24748,N_22155,N_20257);
nor U24749 (N_24749,N_22125,N_21477);
and U24750 (N_24750,N_20746,N_20802);
nor U24751 (N_24751,N_20036,N_21641);
nand U24752 (N_24752,N_21057,N_21937);
nor U24753 (N_24753,N_21054,N_21712);
and U24754 (N_24754,N_20207,N_20464);
or U24755 (N_24755,N_21183,N_21793);
or U24756 (N_24756,N_22236,N_20421);
nand U24757 (N_24757,N_22444,N_21007);
nand U24758 (N_24758,N_22486,N_22286);
or U24759 (N_24759,N_21819,N_21102);
or U24760 (N_24760,N_21039,N_21953);
nor U24761 (N_24761,N_21917,N_22486);
or U24762 (N_24762,N_22100,N_20358);
and U24763 (N_24763,N_22391,N_21393);
and U24764 (N_24764,N_20732,N_20816);
nand U24765 (N_24765,N_20893,N_22289);
xnor U24766 (N_24766,N_22149,N_20196);
nand U24767 (N_24767,N_21697,N_22070);
xnor U24768 (N_24768,N_21459,N_20255);
and U24769 (N_24769,N_20637,N_22010);
or U24770 (N_24770,N_20064,N_21453);
nor U24771 (N_24771,N_21536,N_20498);
and U24772 (N_24772,N_20262,N_20889);
nand U24773 (N_24773,N_21138,N_21113);
nand U24774 (N_24774,N_21604,N_20260);
and U24775 (N_24775,N_21192,N_21951);
nand U24776 (N_24776,N_20438,N_21533);
nand U24777 (N_24777,N_22309,N_20369);
and U24778 (N_24778,N_20098,N_21906);
nand U24779 (N_24779,N_20154,N_22174);
nor U24780 (N_24780,N_21470,N_21999);
nand U24781 (N_24781,N_20190,N_22422);
xor U24782 (N_24782,N_21661,N_21908);
and U24783 (N_24783,N_21026,N_22108);
or U24784 (N_24784,N_20819,N_20798);
or U24785 (N_24785,N_21453,N_21457);
nor U24786 (N_24786,N_20119,N_22024);
and U24787 (N_24787,N_20465,N_22243);
nor U24788 (N_24788,N_20132,N_22389);
nor U24789 (N_24789,N_20430,N_20766);
xnor U24790 (N_24790,N_20964,N_21165);
xor U24791 (N_24791,N_21124,N_20216);
and U24792 (N_24792,N_21443,N_21664);
or U24793 (N_24793,N_20855,N_20046);
and U24794 (N_24794,N_20271,N_22149);
and U24795 (N_24795,N_22421,N_21353);
or U24796 (N_24796,N_21917,N_20220);
or U24797 (N_24797,N_21181,N_22465);
xor U24798 (N_24798,N_22365,N_22190);
nor U24799 (N_24799,N_22043,N_20811);
and U24800 (N_24800,N_21657,N_21412);
nor U24801 (N_24801,N_21408,N_20100);
nor U24802 (N_24802,N_21531,N_22299);
nor U24803 (N_24803,N_20255,N_21006);
nand U24804 (N_24804,N_21358,N_22451);
nand U24805 (N_24805,N_20398,N_21832);
or U24806 (N_24806,N_22347,N_20377);
nand U24807 (N_24807,N_21635,N_20147);
and U24808 (N_24808,N_21133,N_20732);
nand U24809 (N_24809,N_21541,N_20436);
and U24810 (N_24810,N_20830,N_22154);
xnor U24811 (N_24811,N_20743,N_21784);
xnor U24812 (N_24812,N_20740,N_20268);
nor U24813 (N_24813,N_22473,N_20606);
or U24814 (N_24814,N_20110,N_21978);
or U24815 (N_24815,N_22317,N_20244);
nor U24816 (N_24816,N_20519,N_20802);
nand U24817 (N_24817,N_21630,N_21478);
or U24818 (N_24818,N_20230,N_22146);
and U24819 (N_24819,N_20073,N_20033);
nand U24820 (N_24820,N_21255,N_22107);
xor U24821 (N_24821,N_20651,N_21429);
or U24822 (N_24822,N_21839,N_20416);
or U24823 (N_24823,N_21808,N_21896);
xnor U24824 (N_24824,N_20436,N_20859);
and U24825 (N_24825,N_22036,N_20552);
nor U24826 (N_24826,N_20871,N_20411);
nor U24827 (N_24827,N_20447,N_21193);
or U24828 (N_24828,N_21276,N_20910);
or U24829 (N_24829,N_22272,N_20525);
xnor U24830 (N_24830,N_21197,N_22291);
or U24831 (N_24831,N_21688,N_21699);
xor U24832 (N_24832,N_22420,N_21428);
nand U24833 (N_24833,N_20314,N_22254);
or U24834 (N_24834,N_22232,N_20160);
or U24835 (N_24835,N_22261,N_22273);
or U24836 (N_24836,N_21486,N_20731);
nand U24837 (N_24837,N_20015,N_20142);
or U24838 (N_24838,N_22349,N_21439);
nor U24839 (N_24839,N_22001,N_20189);
and U24840 (N_24840,N_21678,N_21477);
nor U24841 (N_24841,N_21931,N_21641);
or U24842 (N_24842,N_21735,N_22075);
or U24843 (N_24843,N_21423,N_21882);
or U24844 (N_24844,N_20677,N_20512);
and U24845 (N_24845,N_21204,N_21165);
nand U24846 (N_24846,N_20127,N_20410);
nor U24847 (N_24847,N_21204,N_21011);
nor U24848 (N_24848,N_21960,N_21404);
nor U24849 (N_24849,N_22497,N_21112);
and U24850 (N_24850,N_22277,N_22445);
and U24851 (N_24851,N_22040,N_20407);
nor U24852 (N_24852,N_20388,N_20808);
xnor U24853 (N_24853,N_21808,N_20809);
or U24854 (N_24854,N_20698,N_21678);
nand U24855 (N_24855,N_21302,N_20160);
nor U24856 (N_24856,N_21905,N_20213);
xor U24857 (N_24857,N_20601,N_20092);
nor U24858 (N_24858,N_22227,N_20630);
and U24859 (N_24859,N_21847,N_20838);
nor U24860 (N_24860,N_20096,N_22376);
or U24861 (N_24861,N_21173,N_21587);
nand U24862 (N_24862,N_21044,N_22454);
and U24863 (N_24863,N_22491,N_22020);
nor U24864 (N_24864,N_22266,N_22352);
nand U24865 (N_24865,N_20645,N_21669);
xor U24866 (N_24866,N_20559,N_21708);
nand U24867 (N_24867,N_22181,N_22253);
nand U24868 (N_24868,N_20621,N_21348);
nor U24869 (N_24869,N_20225,N_20417);
nor U24870 (N_24870,N_21225,N_22498);
or U24871 (N_24871,N_21194,N_20745);
xor U24872 (N_24872,N_20611,N_21350);
or U24873 (N_24873,N_21651,N_22123);
and U24874 (N_24874,N_22373,N_21243);
nand U24875 (N_24875,N_20364,N_20564);
nand U24876 (N_24876,N_21092,N_20546);
nor U24877 (N_24877,N_22456,N_20984);
and U24878 (N_24878,N_22466,N_21526);
and U24879 (N_24879,N_21010,N_20816);
nand U24880 (N_24880,N_21976,N_21858);
nor U24881 (N_24881,N_20236,N_21315);
xnor U24882 (N_24882,N_20133,N_20354);
nor U24883 (N_24883,N_21190,N_20676);
nor U24884 (N_24884,N_21996,N_21708);
xnor U24885 (N_24885,N_21180,N_22124);
nand U24886 (N_24886,N_21810,N_22203);
xnor U24887 (N_24887,N_20977,N_20850);
nand U24888 (N_24888,N_20461,N_22446);
or U24889 (N_24889,N_21685,N_21686);
nor U24890 (N_24890,N_21390,N_22094);
or U24891 (N_24891,N_21138,N_20058);
or U24892 (N_24892,N_21392,N_20551);
nand U24893 (N_24893,N_21847,N_21260);
nand U24894 (N_24894,N_21167,N_21728);
xor U24895 (N_24895,N_20872,N_20120);
or U24896 (N_24896,N_22446,N_21493);
and U24897 (N_24897,N_21963,N_21118);
xnor U24898 (N_24898,N_22330,N_21863);
nand U24899 (N_24899,N_21184,N_20475);
or U24900 (N_24900,N_21286,N_21513);
xnor U24901 (N_24901,N_20717,N_20898);
or U24902 (N_24902,N_21979,N_22214);
and U24903 (N_24903,N_21932,N_21467);
nand U24904 (N_24904,N_20036,N_22310);
xnor U24905 (N_24905,N_20602,N_21908);
and U24906 (N_24906,N_20646,N_21528);
and U24907 (N_24907,N_21750,N_20422);
or U24908 (N_24908,N_21677,N_22026);
and U24909 (N_24909,N_22325,N_22473);
xnor U24910 (N_24910,N_21825,N_20062);
xor U24911 (N_24911,N_21187,N_20020);
or U24912 (N_24912,N_21775,N_20681);
nand U24913 (N_24913,N_20599,N_20431);
nand U24914 (N_24914,N_21246,N_20674);
or U24915 (N_24915,N_21792,N_21957);
and U24916 (N_24916,N_21794,N_20115);
or U24917 (N_24917,N_20255,N_22021);
nor U24918 (N_24918,N_22029,N_20154);
xnor U24919 (N_24919,N_21726,N_20809);
xor U24920 (N_24920,N_22093,N_21572);
nand U24921 (N_24921,N_21951,N_21509);
nor U24922 (N_24922,N_21839,N_20294);
and U24923 (N_24923,N_22448,N_20824);
or U24924 (N_24924,N_21139,N_20467);
nor U24925 (N_24925,N_21651,N_21298);
nor U24926 (N_24926,N_21400,N_20028);
nor U24927 (N_24927,N_21623,N_22302);
nand U24928 (N_24928,N_20939,N_22328);
or U24929 (N_24929,N_20402,N_21104);
nor U24930 (N_24930,N_22466,N_21745);
xnor U24931 (N_24931,N_21059,N_22421);
nand U24932 (N_24932,N_22211,N_22187);
nor U24933 (N_24933,N_22228,N_20127);
and U24934 (N_24934,N_20741,N_21949);
or U24935 (N_24935,N_21944,N_21357);
or U24936 (N_24936,N_20820,N_21699);
nand U24937 (N_24937,N_20318,N_21100);
nor U24938 (N_24938,N_21727,N_21122);
nor U24939 (N_24939,N_21307,N_21698);
xor U24940 (N_24940,N_21502,N_20820);
or U24941 (N_24941,N_21187,N_22249);
nor U24942 (N_24942,N_21205,N_21788);
and U24943 (N_24943,N_22411,N_21261);
nor U24944 (N_24944,N_22371,N_20497);
or U24945 (N_24945,N_22134,N_21902);
nand U24946 (N_24946,N_20455,N_20737);
or U24947 (N_24947,N_22168,N_20373);
and U24948 (N_24948,N_22237,N_22176);
or U24949 (N_24949,N_22110,N_20700);
nor U24950 (N_24950,N_20915,N_20458);
xnor U24951 (N_24951,N_21122,N_22220);
and U24952 (N_24952,N_21201,N_20159);
or U24953 (N_24953,N_22117,N_22476);
and U24954 (N_24954,N_20645,N_21382);
xnor U24955 (N_24955,N_20078,N_20656);
nand U24956 (N_24956,N_20742,N_21764);
nand U24957 (N_24957,N_20142,N_22158);
nand U24958 (N_24958,N_20454,N_21560);
nand U24959 (N_24959,N_21846,N_22388);
or U24960 (N_24960,N_20402,N_21853);
nor U24961 (N_24961,N_21482,N_21545);
nor U24962 (N_24962,N_20372,N_22299);
and U24963 (N_24963,N_20072,N_20949);
nand U24964 (N_24964,N_20803,N_21125);
or U24965 (N_24965,N_21450,N_20359);
and U24966 (N_24966,N_21817,N_22046);
and U24967 (N_24967,N_21112,N_21991);
nand U24968 (N_24968,N_21708,N_20188);
and U24969 (N_24969,N_21484,N_21472);
or U24970 (N_24970,N_20986,N_22266);
or U24971 (N_24971,N_22216,N_20561);
xor U24972 (N_24972,N_20679,N_22409);
or U24973 (N_24973,N_20488,N_21861);
xnor U24974 (N_24974,N_21533,N_20154);
or U24975 (N_24975,N_20838,N_22239);
nand U24976 (N_24976,N_20752,N_22032);
or U24977 (N_24977,N_22451,N_21984);
and U24978 (N_24978,N_20636,N_21613);
nand U24979 (N_24979,N_21895,N_20436);
and U24980 (N_24980,N_21694,N_21601);
nor U24981 (N_24981,N_20339,N_20744);
nand U24982 (N_24982,N_21271,N_20116);
nor U24983 (N_24983,N_21296,N_21521);
and U24984 (N_24984,N_20437,N_22483);
xor U24985 (N_24985,N_20754,N_22430);
xnor U24986 (N_24986,N_21703,N_21922);
xor U24987 (N_24987,N_20304,N_21248);
nor U24988 (N_24988,N_22432,N_21871);
xnor U24989 (N_24989,N_22030,N_21066);
and U24990 (N_24990,N_20077,N_21367);
xnor U24991 (N_24991,N_20779,N_21211);
and U24992 (N_24992,N_21509,N_22244);
and U24993 (N_24993,N_20921,N_20704);
nand U24994 (N_24994,N_20977,N_21184);
and U24995 (N_24995,N_21291,N_21600);
xor U24996 (N_24996,N_21450,N_21617);
or U24997 (N_24997,N_22128,N_20527);
nand U24998 (N_24998,N_20234,N_21938);
and U24999 (N_24999,N_20532,N_21652);
and UO_0 (O_0,N_24932,N_24668);
and UO_1 (O_1,N_22806,N_24086);
and UO_2 (O_2,N_24113,N_23879);
nor UO_3 (O_3,N_22565,N_24685);
nand UO_4 (O_4,N_23380,N_22980);
xnor UO_5 (O_5,N_24515,N_22679);
and UO_6 (O_6,N_23820,N_24168);
xnor UO_7 (O_7,N_24952,N_23697);
nand UO_8 (O_8,N_23114,N_24410);
and UO_9 (O_9,N_24691,N_24536);
xor UO_10 (O_10,N_24804,N_22705);
nor UO_11 (O_11,N_23957,N_24839);
and UO_12 (O_12,N_23551,N_23797);
and UO_13 (O_13,N_23994,N_22684);
and UO_14 (O_14,N_24366,N_24078);
nor UO_15 (O_15,N_23967,N_24651);
xor UO_16 (O_16,N_22732,N_24429);
nor UO_17 (O_17,N_23586,N_22551);
nand UO_18 (O_18,N_23325,N_22895);
or UO_19 (O_19,N_23106,N_22814);
xnor UO_20 (O_20,N_23687,N_24219);
nor UO_21 (O_21,N_24434,N_24692);
nor UO_22 (O_22,N_23061,N_22623);
nor UO_23 (O_23,N_24484,N_24196);
and UO_24 (O_24,N_24686,N_23269);
xnor UO_25 (O_25,N_24714,N_23230);
nand UO_26 (O_26,N_22636,N_23851);
nor UO_27 (O_27,N_23195,N_23585);
and UO_28 (O_28,N_22571,N_22644);
nor UO_29 (O_29,N_24943,N_23632);
or UO_30 (O_30,N_22745,N_23920);
nor UO_31 (O_31,N_24235,N_24173);
or UO_32 (O_32,N_24549,N_22560);
and UO_33 (O_33,N_23620,N_24676);
nor UO_34 (O_34,N_23467,N_24067);
xnor UO_35 (O_35,N_24285,N_24176);
nand UO_36 (O_36,N_24497,N_23088);
xor UO_37 (O_37,N_22642,N_22601);
nor UO_38 (O_38,N_22610,N_23464);
and UO_39 (O_39,N_24944,N_23649);
or UO_40 (O_40,N_23404,N_24191);
nor UO_41 (O_41,N_22934,N_24684);
or UO_42 (O_42,N_24994,N_22885);
nand UO_43 (O_43,N_22824,N_23117);
or UO_44 (O_44,N_22634,N_23939);
nor UO_45 (O_45,N_23877,N_23615);
nor UO_46 (O_46,N_24328,N_24619);
nand UO_47 (O_47,N_24316,N_23321);
and UO_48 (O_48,N_24566,N_23386);
and UO_49 (O_49,N_24836,N_23223);
and UO_50 (O_50,N_22606,N_23107);
nor UO_51 (O_51,N_22658,N_24520);
and UO_52 (O_52,N_23160,N_24160);
and UO_53 (O_53,N_22817,N_24343);
xnor UO_54 (O_54,N_23574,N_24025);
nand UO_55 (O_55,N_24826,N_22665);
or UO_56 (O_56,N_23528,N_23854);
nor UO_57 (O_57,N_23701,N_23005);
xor UO_58 (O_58,N_23457,N_23392);
or UO_59 (O_59,N_23906,N_24539);
nor UO_60 (O_60,N_24808,N_23788);
nand UO_61 (O_61,N_23739,N_23864);
nor UO_62 (O_62,N_24421,N_24682);
xnor UO_63 (O_63,N_22905,N_24659);
and UO_64 (O_64,N_24217,N_23628);
nand UO_65 (O_65,N_24650,N_23372);
nor UO_66 (O_66,N_23110,N_23575);
and UO_67 (O_67,N_23816,N_24491);
xnor UO_68 (O_68,N_24529,N_24912);
nor UO_69 (O_69,N_24838,N_23388);
and UO_70 (O_70,N_22608,N_23874);
nand UO_71 (O_71,N_24295,N_23358);
nor UO_72 (O_72,N_22585,N_24817);
nor UO_73 (O_73,N_23109,N_23261);
xnor UO_74 (O_74,N_24288,N_24026);
and UO_75 (O_75,N_23071,N_24396);
xnor UO_76 (O_76,N_24260,N_24440);
or UO_77 (O_77,N_22852,N_23095);
nand UO_78 (O_78,N_23985,N_23112);
and UO_79 (O_79,N_22555,N_24679);
nand UO_80 (O_80,N_22762,N_22688);
or UO_81 (O_81,N_24517,N_24381);
nor UO_82 (O_82,N_23813,N_24130);
or UO_83 (O_83,N_22641,N_23278);
nor UO_84 (O_84,N_22740,N_23014);
or UO_85 (O_85,N_23188,N_24828);
or UO_86 (O_86,N_24044,N_22954);
or UO_87 (O_87,N_23393,N_24278);
xor UO_88 (O_88,N_24178,N_24068);
nor UO_89 (O_89,N_23237,N_23431);
or UO_90 (O_90,N_22648,N_24835);
and UO_91 (O_91,N_22906,N_23684);
or UO_92 (O_92,N_23728,N_22540);
nor UO_93 (O_93,N_24174,N_24114);
xnor UO_94 (O_94,N_22556,N_22953);
or UO_95 (O_95,N_22637,N_22982);
nand UO_96 (O_96,N_22780,N_22914);
or UO_97 (O_97,N_24273,N_24494);
nand UO_98 (O_98,N_23795,N_24495);
and UO_99 (O_99,N_23598,N_22963);
nand UO_100 (O_100,N_24030,N_24941);
or UO_101 (O_101,N_24541,N_24865);
or UO_102 (O_102,N_23972,N_24577);
nand UO_103 (O_103,N_24034,N_23113);
and UO_104 (O_104,N_23449,N_23447);
and UO_105 (O_105,N_22561,N_22598);
xor UO_106 (O_106,N_24470,N_23639);
or UO_107 (O_107,N_23724,N_24939);
or UO_108 (O_108,N_23720,N_23206);
nor UO_109 (O_109,N_24351,N_23955);
nor UO_110 (O_110,N_22671,N_23891);
nor UO_111 (O_111,N_23248,N_22809);
nand UO_112 (O_112,N_24562,N_24032);
xnor UO_113 (O_113,N_24527,N_22810);
nor UO_114 (O_114,N_24731,N_24048);
xor UO_115 (O_115,N_23072,N_23881);
nor UO_116 (O_116,N_24853,N_24959);
nor UO_117 (O_117,N_24979,N_24404);
or UO_118 (O_118,N_24813,N_23410);
nand UO_119 (O_119,N_23463,N_23870);
and UO_120 (O_120,N_23159,N_23921);
nor UO_121 (O_121,N_23666,N_24613);
nand UO_122 (O_122,N_23396,N_23763);
xor UO_123 (O_123,N_23013,N_24200);
nand UO_124 (O_124,N_22876,N_23988);
nor UO_125 (O_125,N_24098,N_23260);
or UO_126 (O_126,N_23274,N_23518);
or UO_127 (O_127,N_23568,N_22510);
xor UO_128 (O_128,N_22948,N_23015);
and UO_129 (O_129,N_23187,N_23400);
nand UO_130 (O_130,N_24754,N_23166);
or UO_131 (O_131,N_24490,N_24573);
nor UO_132 (O_132,N_24337,N_24179);
xor UO_133 (O_133,N_22795,N_24166);
or UO_134 (O_134,N_22723,N_24774);
and UO_135 (O_135,N_24043,N_24960);
and UO_136 (O_136,N_23408,N_23613);
and UO_137 (O_137,N_24866,N_23593);
or UO_138 (O_138,N_23902,N_23658);
nand UO_139 (O_139,N_24474,N_23818);
nor UO_140 (O_140,N_23963,N_23180);
nor UO_141 (O_141,N_23706,N_23612);
and UO_142 (O_142,N_24291,N_24307);
or UO_143 (O_143,N_24654,N_22942);
nor UO_144 (O_144,N_24533,N_23983);
and UO_145 (O_145,N_24304,N_24807);
or UO_146 (O_146,N_24252,N_24847);
or UO_147 (O_147,N_24131,N_22908);
nor UO_148 (O_148,N_22656,N_22528);
nor UO_149 (O_149,N_23846,N_24531);
xnor UO_150 (O_150,N_23366,N_23653);
xnor UO_151 (O_151,N_23169,N_24793);
and UO_152 (O_152,N_24906,N_23233);
nor UO_153 (O_153,N_24742,N_24128);
or UO_154 (O_154,N_22760,N_23490);
nor UO_155 (O_155,N_24358,N_23442);
nor UO_156 (O_156,N_23996,N_24698);
nor UO_157 (O_157,N_23297,N_24987);
and UO_158 (O_158,N_22946,N_23554);
nand UO_159 (O_159,N_22964,N_22850);
or UO_160 (O_160,N_24765,N_22902);
xor UO_161 (O_161,N_24053,N_23430);
nor UO_162 (O_162,N_23726,N_24707);
xnor UO_163 (O_163,N_22835,N_24661);
nand UO_164 (O_164,N_24864,N_24171);
or UO_165 (O_165,N_24123,N_23049);
or UO_166 (O_166,N_24559,N_24518);
and UO_167 (O_167,N_23415,N_24112);
nor UO_168 (O_168,N_24587,N_22831);
or UO_169 (O_169,N_24482,N_24596);
or UO_170 (O_170,N_22886,N_22582);
or UO_171 (O_171,N_24700,N_23221);
nor UO_172 (O_172,N_23456,N_23163);
xnor UO_173 (O_173,N_23709,N_22757);
xnor UO_174 (O_174,N_23207,N_23084);
nor UO_175 (O_175,N_23191,N_24747);
or UO_176 (O_176,N_24936,N_23312);
xnor UO_177 (O_177,N_24846,N_23893);
nor UO_178 (O_178,N_22568,N_23525);
or UO_179 (O_179,N_24127,N_24733);
xor UO_180 (O_180,N_23572,N_24869);
nor UO_181 (O_181,N_24095,N_24124);
nor UO_182 (O_182,N_24323,N_23643);
or UO_183 (O_183,N_22931,N_23362);
or UO_184 (O_184,N_24792,N_24418);
or UO_185 (O_185,N_23287,N_22566);
nor UO_186 (O_186,N_22773,N_24362);
and UO_187 (O_187,N_24262,N_24796);
and UO_188 (O_188,N_23129,N_23236);
or UO_189 (O_189,N_24963,N_24672);
or UO_190 (O_190,N_24066,N_23942);
nand UO_191 (O_191,N_24312,N_24221);
xnor UO_192 (O_192,N_24955,N_23521);
and UO_193 (O_193,N_23617,N_24580);
and UO_194 (O_194,N_24354,N_24634);
or UO_195 (O_195,N_24732,N_24333);
or UO_196 (O_196,N_22853,N_23944);
xor UO_197 (O_197,N_24321,N_22748);
and UO_198 (O_198,N_23645,N_22881);
and UO_199 (O_199,N_24775,N_24727);
nor UO_200 (O_200,N_23059,N_24790);
and UO_201 (O_201,N_23412,N_24473);
nand UO_202 (O_202,N_24724,N_24783);
xor UO_203 (O_203,N_24188,N_23611);
or UO_204 (O_204,N_23308,N_24883);
nand UO_205 (O_205,N_23968,N_24085);
and UO_206 (O_206,N_24287,N_23466);
and UO_207 (O_207,N_24371,N_23473);
and UO_208 (O_208,N_22532,N_23975);
nand UO_209 (O_209,N_23503,N_24882);
nand UO_210 (O_210,N_23493,N_23644);
xnor UO_211 (O_211,N_23200,N_22657);
or UO_212 (O_212,N_24310,N_24526);
xor UO_213 (O_213,N_23419,N_23197);
nand UO_214 (O_214,N_22631,N_23642);
and UO_215 (O_215,N_23772,N_23422);
xnor UO_216 (O_216,N_22559,N_23334);
xnor UO_217 (O_217,N_23984,N_23945);
and UO_218 (O_218,N_24194,N_24223);
and UO_219 (O_219,N_22645,N_24528);
and UO_220 (O_220,N_24286,N_23588);
and UO_221 (O_221,N_24855,N_24426);
or UO_222 (O_222,N_23861,N_23142);
nand UO_223 (O_223,N_23783,N_23465);
nand UO_224 (O_224,N_24635,N_23801);
or UO_225 (O_225,N_24555,N_23745);
xnor UO_226 (O_226,N_24175,N_24675);
and UO_227 (O_227,N_24997,N_23776);
nand UO_228 (O_228,N_22678,N_23426);
xor UO_229 (O_229,N_22917,N_23262);
nor UO_230 (O_230,N_24597,N_23686);
and UO_231 (O_231,N_23252,N_23986);
nand UO_232 (O_232,N_23428,N_24225);
xor UO_233 (O_233,N_23699,N_24544);
and UO_234 (O_234,N_22900,N_23799);
nand UO_235 (O_235,N_22668,N_23053);
or UO_236 (O_236,N_23842,N_23479);
nand UO_237 (O_237,N_23173,N_23841);
xnor UO_238 (O_238,N_22974,N_22919);
xnor UO_239 (O_239,N_24207,N_24438);
nand UO_240 (O_240,N_23273,N_22916);
or UO_241 (O_241,N_22769,N_23373);
xor UO_242 (O_242,N_22758,N_22883);
or UO_243 (O_243,N_23011,N_22765);
nand UO_244 (O_244,N_22703,N_24639);
nor UO_245 (O_245,N_24324,N_23682);
nor UO_246 (O_246,N_23276,N_23116);
xor UO_247 (O_247,N_22533,N_23830);
and UO_248 (O_248,N_24852,N_23494);
xor UO_249 (O_249,N_24636,N_22949);
nand UO_250 (O_250,N_24632,N_22801);
nand UO_251 (O_251,N_24002,N_22846);
nand UO_252 (O_252,N_24694,N_22844);
and UO_253 (O_253,N_23217,N_24588);
nor UO_254 (O_254,N_24728,N_22522);
and UO_255 (O_255,N_24688,N_24914);
nand UO_256 (O_256,N_24956,N_22878);
nor UO_257 (O_257,N_24364,N_23520);
xor UO_258 (O_258,N_24970,N_23785);
or UO_259 (O_259,N_24301,N_24598);
and UO_260 (O_260,N_23758,N_24851);
nand UO_261 (O_261,N_24195,N_23685);
or UO_262 (O_262,N_24172,N_24340);
nand UO_263 (O_263,N_22720,N_22874);
nor UO_264 (O_264,N_23285,N_23461);
nand UO_265 (O_265,N_24778,N_23707);
and UO_266 (O_266,N_24144,N_24054);
or UO_267 (O_267,N_23486,N_23244);
nor UO_268 (O_268,N_23452,N_24452);
and UO_269 (O_269,N_23829,N_24663);
nand UO_270 (O_270,N_23213,N_23634);
and UO_271 (O_271,N_23601,N_24844);
xor UO_272 (O_272,N_24388,N_23212);
nand UO_273 (O_273,N_23176,N_24918);
and UO_274 (O_274,N_24090,N_23363);
nand UO_275 (O_275,N_24547,N_23789);
nand UO_276 (O_276,N_22803,N_23310);
or UO_277 (O_277,N_24748,N_22880);
or UO_278 (O_278,N_23669,N_24079);
nand UO_279 (O_279,N_24523,N_24087);
xnor UO_280 (O_280,N_23048,N_24831);
nor UO_281 (O_281,N_23827,N_23171);
nor UO_282 (O_282,N_22713,N_23122);
xnor UO_283 (O_283,N_24193,N_22664);
or UO_284 (O_284,N_22866,N_23040);
nand UO_285 (O_285,N_24135,N_22500);
nor UO_286 (O_286,N_22915,N_24655);
nor UO_287 (O_287,N_24355,N_23606);
nor UO_288 (O_288,N_22797,N_24103);
or UO_289 (O_289,N_22674,N_22896);
or UO_290 (O_290,N_22719,N_23488);
nand UO_291 (O_291,N_23712,N_24208);
and UO_292 (O_292,N_24806,N_23343);
and UO_293 (O_293,N_22513,N_24317);
nand UO_294 (O_294,N_24899,N_23865);
xnor UO_295 (O_295,N_24779,N_24623);
xnor UO_296 (O_296,N_22708,N_24819);
or UO_297 (O_297,N_23327,N_22763);
nand UO_298 (O_298,N_24513,N_23735);
nor UO_299 (O_299,N_24931,N_24590);
nor UO_300 (O_300,N_24848,N_23347);
xor UO_301 (O_301,N_22787,N_22984);
nand UO_302 (O_302,N_23914,N_22518);
or UO_303 (O_303,N_24673,N_24722);
or UO_304 (O_304,N_24109,N_22952);
nand UO_305 (O_305,N_24662,N_23659);
and UO_306 (O_306,N_23876,N_23924);
and UO_307 (O_307,N_24226,N_22932);
xor UO_308 (O_308,N_24416,N_23951);
nand UO_309 (O_309,N_24561,N_24137);
nor UO_310 (O_310,N_24010,N_24772);
nand UO_311 (O_311,N_23516,N_23042);
nand UO_312 (O_312,N_22956,N_22847);
nand UO_313 (O_313,N_24534,N_22816);
nand UO_314 (O_314,N_22981,N_24677);
and UO_315 (O_315,N_23245,N_23766);
xor UO_316 (O_316,N_22659,N_23271);
nor UO_317 (O_317,N_24446,N_24530);
xor UO_318 (O_318,N_24187,N_24795);
nor UO_319 (O_319,N_23616,N_23913);
or UO_320 (O_320,N_24346,N_23900);
xor UO_321 (O_321,N_24063,N_22596);
nand UO_322 (O_322,N_22667,N_24149);
or UO_323 (O_323,N_23296,N_24510);
nor UO_324 (O_324,N_23065,N_22979);
xnor UO_325 (O_325,N_24630,N_23539);
nand UO_326 (O_326,N_23154,N_24671);
or UO_327 (O_327,N_24406,N_24080);
nor UO_328 (O_328,N_22989,N_23101);
and UO_329 (O_329,N_24981,N_23307);
and UO_330 (O_330,N_23134,N_23757);
and UO_331 (O_331,N_23306,N_24600);
nand UO_332 (O_332,N_24105,N_22647);
nand UO_333 (O_333,N_22699,N_24266);
xnor UO_334 (O_334,N_24980,N_23774);
nor UO_335 (O_335,N_23637,N_22807);
xnor UO_336 (O_336,N_23094,N_23663);
xnor UO_337 (O_337,N_22589,N_24075);
and UO_338 (O_338,N_24309,N_23542);
or UO_339 (O_339,N_23204,N_23599);
or UO_340 (O_340,N_23569,N_23375);
or UO_341 (O_341,N_23872,N_23203);
and UO_342 (O_342,N_24665,N_23304);
nand UO_343 (O_343,N_24107,N_23641);
and UO_344 (O_344,N_23246,N_24331);
xnor UO_345 (O_345,N_23499,N_23690);
nand UO_346 (O_346,N_23125,N_23556);
xnor UO_347 (O_347,N_23381,N_23582);
or UO_348 (O_348,N_23771,N_22509);
or UO_349 (O_349,N_22891,N_23469);
nand UO_350 (O_350,N_23597,N_24907);
nor UO_351 (O_351,N_24065,N_24269);
and UO_352 (O_352,N_23406,N_23218);
nor UO_353 (O_353,N_23021,N_24167);
and UO_354 (O_354,N_22965,N_24190);
nor UO_355 (O_355,N_24858,N_22976);
and UO_356 (O_356,N_22843,N_24644);
xor UO_357 (O_357,N_23216,N_24320);
or UO_358 (O_358,N_23522,N_24803);
xor UO_359 (O_359,N_23715,N_23567);
nand UO_360 (O_360,N_24611,N_24435);
nor UO_361 (O_361,N_23622,N_23385);
and UO_362 (O_362,N_24957,N_23662);
xor UO_363 (O_363,N_24432,N_24076);
nand UO_364 (O_364,N_24349,N_23889);
and UO_365 (O_365,N_22635,N_24021);
xor UO_366 (O_366,N_23108,N_22633);
and UO_367 (O_367,N_22800,N_23135);
xnor UO_368 (O_368,N_24061,N_23787);
xor UO_369 (O_369,N_22789,N_22620);
or UO_370 (O_370,N_23577,N_24723);
xnor UO_371 (O_371,N_24378,N_23483);
xnor UO_372 (O_372,N_23198,N_23843);
or UO_373 (O_373,N_24894,N_23661);
xor UO_374 (O_374,N_23727,N_22604);
xor UO_375 (O_375,N_23350,N_23258);
and UO_376 (O_376,N_24220,N_23179);
nand UO_377 (O_377,N_23417,N_24911);
or UO_378 (O_378,N_24845,N_22652);
nand UO_379 (O_379,N_24905,N_23930);
nand UO_380 (O_380,N_24568,N_24360);
xor UO_381 (O_381,N_22783,N_23377);
or UO_382 (O_382,N_24315,N_24624);
xor UO_383 (O_383,N_23062,N_23079);
or UO_384 (O_384,N_22672,N_24903);
or UO_385 (O_385,N_22542,N_23235);
nor UO_386 (O_386,N_23349,N_24570);
or UO_387 (O_387,N_24447,N_23121);
xor UO_388 (O_388,N_22832,N_23768);
nor UO_389 (O_389,N_24966,N_22756);
or UO_390 (O_390,N_24110,N_23150);
or UO_391 (O_391,N_24591,N_23282);
and UO_392 (O_392,N_22863,N_24605);
nor UO_393 (O_393,N_22693,N_22887);
and UO_394 (O_394,N_23806,N_24256);
nand UO_395 (O_395,N_22779,N_23755);
nand UO_396 (O_396,N_23566,N_24007);
and UO_397 (O_397,N_22577,N_24581);
nor UO_398 (O_398,N_23484,N_23770);
and UO_399 (O_399,N_23186,N_22815);
nand UO_400 (O_400,N_23627,N_23681);
nand UO_401 (O_401,N_24117,N_23729);
xor UO_402 (O_402,N_22840,N_23182);
nor UO_403 (O_403,N_23438,N_22534);
and UO_404 (O_404,N_23916,N_24326);
and UO_405 (O_405,N_24824,N_23950);
nand UO_406 (O_406,N_24478,N_22990);
and UO_407 (O_407,N_23012,N_22957);
and UO_408 (O_408,N_24586,N_24119);
and UO_409 (O_409,N_24827,N_23324);
nor UO_410 (O_410,N_22727,N_22753);
nor UO_411 (O_411,N_23589,N_22701);
or UO_412 (O_412,N_24525,N_23032);
xor UO_413 (O_413,N_24186,N_23966);
or UO_414 (O_414,N_23565,N_22625);
and UO_415 (O_415,N_24038,N_24427);
nand UO_416 (O_416,N_22928,N_23127);
xnor UO_417 (O_417,N_23692,N_23812);
xnor UO_418 (O_418,N_23835,N_24919);
xor UO_419 (O_419,N_24916,N_23328);
and UO_420 (O_420,N_23030,N_24560);
xnor UO_421 (O_421,N_24993,N_22677);
xor UO_422 (O_422,N_24431,N_23455);
nor UO_423 (O_423,N_22514,N_23676);
and UO_424 (O_424,N_24535,N_24212);
or UO_425 (O_425,N_22697,N_24185);
xnor UO_426 (O_426,N_22512,N_23839);
xor UO_427 (O_427,N_23552,N_23695);
nand UO_428 (O_428,N_23919,N_23249);
or UO_429 (O_429,N_24270,N_23608);
and UO_430 (O_430,N_24948,N_23524);
and UO_431 (O_431,N_22933,N_23550);
nor UO_432 (O_432,N_24242,N_23086);
nor UO_433 (O_433,N_24202,N_23664);
or UO_434 (O_434,N_23299,N_24678);
and UO_435 (O_435,N_24443,N_24437);
and UO_436 (O_436,N_24382,N_23056);
xnor UO_437 (O_437,N_24083,N_23506);
xnor UO_438 (O_438,N_23626,N_24492);
nand UO_439 (O_439,N_24753,N_22823);
xnor UO_440 (O_440,N_22997,N_23091);
or UO_441 (O_441,N_24592,N_23859);
or UO_442 (O_442,N_23918,N_23177);
or UO_443 (O_443,N_23723,N_22517);
and UO_444 (O_444,N_24729,N_24383);
xor UO_445 (O_445,N_24777,N_22550);
xnor UO_446 (O_446,N_24551,N_24949);
and UO_447 (O_447,N_24282,N_23069);
and UO_448 (O_448,N_24203,N_23540);
nor UO_449 (O_449,N_24913,N_24457);
or UO_450 (O_450,N_23275,N_23409);
xor UO_451 (O_451,N_23781,N_24626);
and UO_452 (O_452,N_23650,N_23534);
xnor UO_453 (O_453,N_23096,N_23845);
or UO_454 (O_454,N_23873,N_23234);
nand UO_455 (O_455,N_24479,N_23962);
and UO_456 (O_456,N_22735,N_24056);
nor UO_457 (O_457,N_24641,N_22836);
nor UO_458 (O_458,N_23884,N_22581);
or UO_459 (O_459,N_24629,N_23536);
xnor UO_460 (O_460,N_23940,N_24511);
nor UO_461 (O_461,N_24472,N_24254);
and UO_462 (O_462,N_23316,N_24990);
nor UO_463 (O_463,N_24829,N_24213);
nand UO_464 (O_464,N_24380,N_23713);
xor UO_465 (O_465,N_24275,N_23747);
nand UO_466 (O_466,N_23847,N_23253);
xnor UO_467 (O_467,N_24646,N_24766);
nor UO_468 (O_468,N_24893,N_24812);
xnor UO_469 (O_469,N_23387,N_24681);
xor UO_470 (O_470,N_23557,N_22873);
nor UO_471 (O_471,N_23161,N_22638);
nor UO_472 (O_472,N_22818,N_24708);
nor UO_473 (O_473,N_23752,N_24322);
and UO_474 (O_474,N_23737,N_22718);
nor UO_475 (O_475,N_23946,N_24101);
xnor UO_476 (O_476,N_23336,N_22618);
or UO_477 (O_477,N_23667,N_24509);
nand UO_478 (O_478,N_24029,N_24537);
or UO_479 (O_479,N_23132,N_23630);
nor UO_480 (O_480,N_23317,N_22670);
nand UO_481 (O_481,N_23383,N_24519);
or UO_482 (O_482,N_24627,N_23093);
xnor UO_483 (O_483,N_24445,N_23264);
nor UO_484 (O_484,N_24003,N_23819);
or UO_485 (O_485,N_23738,N_23498);
xnor UO_486 (O_486,N_24718,N_22988);
or UO_487 (O_487,N_22628,N_22736);
xnor UO_488 (O_488,N_22739,N_24585);
nand UO_489 (O_489,N_23024,N_23318);
xnor UO_490 (O_490,N_24788,N_24341);
and UO_491 (O_491,N_23844,N_24199);
nand UO_492 (O_492,N_24461,N_24142);
nand UO_493 (O_493,N_23595,N_23779);
nand UO_494 (O_494,N_23031,N_24386);
nand UO_495 (O_495,N_22629,N_22940);
nand UO_496 (O_496,N_24617,N_22543);
xor UO_497 (O_497,N_24751,N_22655);
nor UO_498 (O_498,N_22707,N_22698);
and UO_499 (O_499,N_23502,N_23761);
or UO_500 (O_500,N_23917,N_23020);
nand UO_501 (O_501,N_24232,N_22893);
xor UO_502 (O_502,N_23482,N_24391);
and UO_503 (O_503,N_24436,N_24228);
and UO_504 (O_504,N_23688,N_24814);
and UO_505 (O_505,N_24376,N_24502);
or UO_506 (O_506,N_23256,N_23636);
nor UO_507 (O_507,N_23340,N_24524);
or UO_508 (O_508,N_23584,N_22775);
or UO_509 (O_509,N_23485,N_22894);
and UO_510 (O_510,N_22729,N_24569);
nand UO_511 (O_511,N_24878,N_24201);
nor UO_512 (O_512,N_22702,N_24247);
or UO_513 (O_513,N_23866,N_24567);
and UO_514 (O_514,N_24872,N_24738);
and UO_515 (O_515,N_22704,N_23046);
xor UO_516 (O_516,N_24475,N_23671);
nand UO_517 (O_517,N_23345,N_23333);
or UO_518 (O_518,N_24721,N_24216);
nor UO_519 (O_519,N_22955,N_23607);
nor UO_520 (O_520,N_24749,N_24258);
xnor UO_521 (O_521,N_23063,N_23401);
xor UO_522 (O_522,N_24099,N_24928);
or UO_523 (O_523,N_22858,N_23886);
nand UO_524 (O_524,N_23051,N_23290);
nand UO_525 (O_525,N_24757,N_24985);
nor UO_526 (O_526,N_24776,N_23579);
nor UO_527 (O_527,N_23468,N_23267);
and UO_528 (O_528,N_23832,N_24915);
xor UO_529 (O_529,N_23155,N_24859);
nand UO_530 (O_530,N_24231,N_24134);
nand UO_531 (O_531,N_24133,N_22788);
or UO_532 (O_532,N_24177,N_22666);
nor UO_533 (O_533,N_23083,N_24444);
and UO_534 (O_534,N_23784,N_22907);
nand UO_535 (O_535,N_24281,N_24233);
or UO_536 (O_536,N_24045,N_22776);
xnor UO_537 (O_537,N_24209,N_24840);
nand UO_538 (O_538,N_23547,N_24701);
nor UO_539 (O_539,N_22680,N_23689);
xnor UO_540 (O_540,N_23369,N_23105);
nand UO_541 (O_541,N_23382,N_22547);
and UO_542 (O_542,N_24031,N_23300);
xnor UO_543 (O_543,N_24822,N_24132);
nand UO_544 (O_544,N_22587,N_24204);
xor UO_545 (O_545,N_24578,N_24480);
xnor UO_546 (O_546,N_24656,N_23016);
nand UO_547 (O_547,N_23298,N_23270);
nand UO_548 (O_548,N_23635,N_24830);
nand UO_549 (O_549,N_24156,N_23691);
nand UO_550 (O_550,N_24715,N_22972);
or UO_551 (O_551,N_24293,N_23501);
xnor UO_552 (O_552,N_23078,N_24720);
nand UO_553 (O_553,N_23224,N_24385);
or UO_554 (O_554,N_24239,N_24582);
or UO_555 (O_555,N_23698,N_24667);
and UO_556 (O_556,N_24246,N_24162);
and UO_557 (O_557,N_22950,N_22774);
nor UO_558 (O_558,N_24377,N_22985);
nand UO_559 (O_559,N_24532,N_24917);
xnor UO_560 (O_560,N_24849,N_23817);
xor UO_561 (O_561,N_24689,N_22826);
xor UO_562 (O_562,N_23090,N_24885);
nand UO_563 (O_563,N_23175,N_23471);
xor UO_564 (O_564,N_24248,N_22761);
nand UO_565 (O_565,N_23826,N_24923);
nand UO_566 (O_566,N_24521,N_24771);
nor UO_567 (O_567,N_22842,N_24325);
xor UO_568 (O_568,N_24442,N_23814);
nor UO_569 (O_569,N_24347,N_24215);
nor UO_570 (O_570,N_23039,N_24249);
and UO_571 (O_571,N_22875,N_22991);
nor UO_572 (O_572,N_22546,N_23979);
and UO_573 (O_573,N_24967,N_24251);
nor UO_574 (O_574,N_23969,N_22889);
xor UO_575 (O_575,N_22920,N_22939);
nand UO_576 (O_576,N_24895,N_23199);
nor UO_577 (O_577,N_24658,N_24294);
or UO_578 (O_578,N_23131,N_23936);
and UO_579 (O_579,N_24261,N_23210);
and UO_580 (O_580,N_23295,N_23541);
or UO_581 (O_581,N_23778,N_24327);
xor UO_582 (O_582,N_24516,N_23609);
nor UO_583 (O_583,N_24740,N_23741);
and UO_584 (O_584,N_23862,N_22890);
or UO_585 (O_585,N_24481,N_22793);
xor UO_586 (O_586,N_22662,N_23808);
xnor UO_587 (O_587,N_24834,N_24236);
nor UO_588 (O_588,N_22975,N_22683);
xnor UO_589 (O_589,N_24290,N_23280);
xor UO_590 (O_590,N_23378,N_23749);
nand UO_591 (O_591,N_22675,N_22929);
or UO_592 (O_592,N_23510,N_24428);
and UO_593 (O_593,N_23998,N_24071);
nand UO_594 (O_594,N_23100,N_24485);
and UO_595 (O_595,N_23007,N_23359);
nand UO_596 (O_596,N_23151,N_24197);
nand UO_597 (O_597,N_24983,N_22868);
xnor UO_598 (O_598,N_23857,N_23674);
and UO_599 (O_599,N_24574,N_24897);
xnor UO_600 (O_600,N_23578,N_22685);
nor UO_601 (O_601,N_24255,N_24794);
nand UO_602 (O_602,N_24140,N_22626);
and UO_603 (O_603,N_24042,N_24401);
xor UO_604 (O_604,N_23453,N_24820);
and UO_605 (O_605,N_24146,N_24934);
or UO_606 (O_606,N_22695,N_22813);
nor UO_607 (O_607,N_23047,N_23474);
nor UO_608 (O_608,N_23477,N_22754);
and UO_609 (O_609,N_24091,N_22994);
nor UO_610 (O_610,N_23790,N_24308);
xor UO_611 (O_611,N_23008,N_24121);
and UO_612 (O_612,N_24781,N_22686);
or UO_613 (O_613,N_24975,N_23120);
and UO_614 (O_614,N_24904,N_23351);
or UO_615 (O_615,N_24842,N_22621);
nor UO_616 (O_616,N_23162,N_22839);
or UO_617 (O_617,N_23899,N_23544);
and UO_618 (O_618,N_22867,N_23558);
xor UO_619 (O_619,N_23947,N_24504);
or UO_620 (O_620,N_23311,N_24250);
nor UO_621 (O_621,N_22600,N_24628);
xor UO_622 (O_622,N_23811,N_24968);
or UO_623 (O_623,N_23754,N_23102);
nand UO_624 (O_624,N_23929,N_24652);
nand UO_625 (O_625,N_22927,N_23205);
and UO_626 (O_626,N_23943,N_23793);
or UO_627 (O_627,N_22599,N_23515);
or UO_628 (O_628,N_24465,N_24764);
and UO_629 (O_629,N_23834,N_22595);
xor UO_630 (O_630,N_23922,N_24815);
and UO_631 (O_631,N_23066,N_24489);
nand UO_632 (O_632,N_23354,N_24976);
or UO_633 (O_633,N_22710,N_24606);
and UO_634 (O_634,N_24860,N_23077);
and UO_635 (O_635,N_24467,N_22766);
nor UO_636 (O_636,N_24594,N_24150);
or UO_637 (O_637,N_24237,N_23730);
nor UO_638 (O_638,N_23330,N_23026);
xor UO_639 (O_639,N_24958,N_24977);
and UO_640 (O_640,N_22694,N_24725);
and UO_641 (O_641,N_24503,N_23931);
and UO_642 (O_642,N_24240,N_23871);
xor UO_643 (O_643,N_24089,N_23614);
nor UO_644 (O_644,N_24498,N_23446);
or UO_645 (O_645,N_22827,N_24744);
xor UO_646 (O_646,N_24369,N_23027);
xor UO_647 (O_647,N_23580,N_24583);
xnor UO_648 (O_648,N_23938,N_24458);
nand UO_649 (O_649,N_22930,N_24441);
xor UO_650 (O_650,N_24802,N_24088);
nor UO_651 (O_651,N_24760,N_22687);
nand UO_652 (O_652,N_24889,N_23355);
or UO_653 (O_653,N_22535,N_22837);
xnor UO_654 (O_654,N_23292,N_23500);
nor UO_655 (O_655,N_23424,N_24041);
nor UO_656 (O_656,N_22590,N_23365);
or UO_657 (O_657,N_23286,N_24716);
nand UO_658 (O_658,N_24014,N_22924);
and UO_659 (O_659,N_23201,N_23035);
nand UO_660 (O_660,N_22926,N_22584);
and UO_661 (O_661,N_23341,N_24477);
or UO_662 (O_662,N_23831,N_24810);
nand UO_663 (O_663,N_24313,N_24051);
nand UO_664 (O_664,N_24283,N_24218);
or UO_665 (O_665,N_23288,N_22515);
and UO_666 (O_666,N_22822,N_24942);
xor UO_667 (O_667,N_23583,N_23156);
xor UO_668 (O_668,N_24222,N_23992);
xnor UO_669 (O_669,N_23596,N_22849);
nor UO_670 (O_670,N_22944,N_22897);
nor UO_671 (O_671,N_23718,N_24991);
xor UO_672 (O_672,N_24005,N_24375);
or UO_673 (O_673,N_23183,N_23773);
nand UO_674 (O_674,N_22999,N_23974);
xnor UO_675 (O_675,N_24973,N_24548);
and UO_676 (O_676,N_22734,N_23167);
nand UO_677 (O_677,N_23148,N_24785);
nand UO_678 (O_678,N_23999,N_22918);
nor UO_679 (O_679,N_22572,N_23982);
nand UO_680 (O_680,N_24756,N_23880);
or UO_681 (O_681,N_22521,N_24758);
nand UO_682 (O_682,N_23678,N_23941);
and UO_683 (O_683,N_23099,N_24460);
nand UO_684 (O_684,N_24153,N_22573);
and UO_685 (O_685,N_23257,N_23704);
and UO_686 (O_686,N_23398,N_24229);
nand UO_687 (O_687,N_22971,N_23553);
xnor UO_688 (O_688,N_23517,N_23711);
or UO_689 (O_689,N_23923,N_24998);
xnor UO_690 (O_690,N_23309,N_23934);
nand UO_691 (O_691,N_24141,N_24799);
xor UO_692 (O_692,N_23139,N_24035);
nor UO_693 (O_693,N_24506,N_24486);
xnor UO_694 (O_694,N_24338,N_22747);
nand UO_695 (O_695,N_23700,N_24669);
xor UO_696 (O_696,N_22996,N_22531);
and UO_697 (O_697,N_23189,N_22519);
or UO_698 (O_698,N_24336,N_24741);
nand UO_699 (O_699,N_23719,N_24610);
or UO_700 (O_700,N_23708,N_22660);
xnor UO_701 (O_701,N_23696,N_24120);
nand UO_702 (O_702,N_24604,N_22935);
nand UO_703 (O_703,N_23855,N_24049);
nor UO_704 (O_704,N_24158,N_23146);
nand UO_705 (O_705,N_23194,N_23303);
nor UO_706 (O_706,N_24945,N_23868);
nand UO_707 (O_707,N_24908,N_24868);
nand UO_708 (O_708,N_23912,N_22937);
nand UO_709 (O_709,N_24768,N_24092);
nor UO_710 (O_710,N_24988,N_22548);
xnor UO_711 (O_711,N_24695,N_23600);
or UO_712 (O_712,N_24155,N_22841);
xnor UO_713 (O_713,N_23981,N_24040);
nand UO_714 (O_714,N_24306,N_24888);
or UO_715 (O_715,N_24947,N_23673);
xnor UO_716 (O_716,N_24015,N_23371);
or UO_717 (O_717,N_23332,N_24933);
nor UO_718 (O_718,N_23802,N_23184);
and UO_719 (O_719,N_23043,N_23389);
nand UO_720 (O_720,N_23815,N_24962);
and UO_721 (O_721,N_23576,N_24621);
and UO_722 (O_722,N_23909,N_24013);
nand UO_723 (O_723,N_23625,N_22570);
nand UO_724 (O_724,N_22778,N_24660);
or UO_725 (O_725,N_24372,N_24522);
nor UO_726 (O_726,N_23057,N_22588);
xnor UO_727 (O_727,N_23519,N_24234);
xnor UO_728 (O_728,N_23140,N_22709);
and UO_729 (O_729,N_22649,N_23390);
xnor UO_730 (O_730,N_24938,N_23937);
nor UO_731 (O_731,N_23315,N_23523);
xnor UO_732 (O_732,N_23978,N_24786);
nand UO_733 (O_733,N_23933,N_24468);
and UO_734 (O_734,N_24552,N_23472);
and UO_735 (O_735,N_23435,N_23460);
nand UO_736 (O_736,N_22947,N_23775);
xor UO_737 (O_737,N_23897,N_22619);
nand UO_738 (O_738,N_24558,N_24069);
or UO_739 (O_739,N_24986,N_24471);
xnor UO_740 (O_740,N_24037,N_24143);
xnor UO_741 (O_741,N_23581,N_24930);
or UO_742 (O_742,N_24033,N_24816);
and UO_743 (O_743,N_23421,N_24397);
nand UO_744 (O_744,N_24488,N_23680);
nand UO_745 (O_745,N_22613,N_24602);
xor UO_746 (O_746,N_22755,N_23734);
and UO_747 (O_747,N_24395,N_24455);
xnor UO_748 (O_748,N_24837,N_22901);
xor UO_749 (O_749,N_23587,N_24181);
and UO_750 (O_750,N_23782,N_24081);
and UO_751 (O_751,N_23251,N_23651);
nand UO_752 (O_752,N_23748,N_23629);
and UO_753 (O_753,N_23890,N_23672);
nand UO_754 (O_754,N_24399,N_22749);
nand UO_755 (O_755,N_23147,N_22970);
or UO_756 (O_756,N_24345,N_23044);
and UO_757 (O_757,N_22503,N_23128);
nand UO_758 (O_758,N_23480,N_24877);
xor UO_759 (O_759,N_24126,N_24996);
xnor UO_760 (O_760,N_23247,N_22508);
or UO_761 (O_761,N_22770,N_24891);
xnor UO_762 (O_762,N_22583,N_23152);
and UO_763 (O_763,N_23995,N_24575);
and UO_764 (O_764,N_24224,N_22856);
and UO_765 (O_765,N_23807,N_24400);
nand UO_766 (O_766,N_23602,N_23824);
xor UO_767 (O_767,N_23003,N_24439);
or UO_768 (O_768,N_22796,N_24192);
xnor UO_769 (O_769,N_24016,N_22862);
or UO_770 (O_770,N_24615,N_24020);
xor UO_771 (O_771,N_24940,N_24999);
and UO_772 (O_772,N_23856,N_23507);
nor UO_773 (O_773,N_22654,N_24407);
nor UO_774 (O_774,N_23853,N_22505);
nor UO_775 (O_775,N_22855,N_22784);
or UO_776 (O_776,N_23397,N_23904);
and UO_777 (O_777,N_23702,N_23443);
and UO_778 (O_778,N_22772,N_23379);
and UO_779 (O_779,N_24750,N_24387);
xor UO_780 (O_780,N_23432,N_23254);
or UO_781 (O_781,N_24995,N_23211);
or UO_782 (O_782,N_23283,N_24147);
xnor UO_783 (O_783,N_23123,N_22830);
and UO_784 (O_784,N_23118,N_23497);
and UO_785 (O_785,N_24730,N_23395);
and UO_786 (O_786,N_23240,N_23036);
and UO_787 (O_787,N_24926,N_24833);
or UO_788 (O_788,N_22854,N_22828);
or UO_789 (O_789,N_23794,N_24241);
nor UO_790 (O_790,N_23693,N_23002);
nor UO_791 (O_791,N_24106,N_24230);
nand UO_792 (O_792,N_24456,N_22650);
and UO_793 (O_793,N_23075,N_22591);
nor UO_794 (O_794,N_23721,N_23869);
xor UO_795 (O_795,N_24084,N_23756);
nor UO_796 (O_796,N_23265,N_24361);
nor UO_797 (O_797,N_23760,N_24394);
and UO_798 (O_798,N_24640,N_23759);
nand UO_799 (O_799,N_23532,N_23034);
nor UO_800 (O_800,N_24879,N_23322);
and UO_801 (O_801,N_24854,N_24011);
and UO_802 (O_802,N_23823,N_22549);
nor UO_803 (O_803,N_24352,N_23137);
xor UO_804 (O_804,N_24297,N_24450);
nand UO_805 (O_805,N_24104,N_23694);
xor UO_806 (O_806,N_23840,N_23594);
or UO_807 (O_807,N_23925,N_24712);
or UO_808 (O_808,N_22643,N_23905);
nor UO_809 (O_809,N_22923,N_24571);
and UO_810 (O_810,N_24330,N_24703);
and UO_811 (O_811,N_24755,N_24350);
and UO_812 (O_812,N_24739,N_24413);
or UO_813 (O_813,N_23915,N_22812);
nand UO_814 (O_814,N_24136,N_23073);
and UO_815 (O_815,N_24901,N_22799);
nor UO_816 (O_816,N_23242,N_22738);
xnor UO_817 (O_817,N_24373,N_22888);
nor UO_818 (O_818,N_22961,N_23948);
nand UO_819 (O_819,N_23025,N_22663);
and UO_820 (O_820,N_24857,N_23633);
nand UO_821 (O_821,N_24616,N_23418);
nand UO_822 (O_822,N_22646,N_24653);
xnor UO_823 (O_823,N_23989,N_22959);
nor UO_824 (O_824,N_22992,N_23677);
or UO_825 (O_825,N_24402,N_23863);
nor UO_826 (O_826,N_23360,N_24409);
or UO_827 (O_827,N_22611,N_22892);
nor UO_828 (O_828,N_22744,N_23145);
or UO_829 (O_829,N_24198,N_24159);
and UO_830 (O_830,N_23563,N_24565);
or UO_831 (O_831,N_23736,N_24890);
nor UO_832 (O_832,N_23860,N_22616);
nor UO_833 (O_833,N_22791,N_22552);
nor UO_834 (O_834,N_22538,N_24398);
or UO_835 (O_835,N_23022,N_23652);
or UO_836 (O_836,N_24463,N_23746);
nor UO_837 (O_837,N_23987,N_23439);
nor UO_838 (O_838,N_24546,N_23076);
or UO_839 (O_839,N_22750,N_23289);
nor UO_840 (O_840,N_23764,N_22523);
nand UO_841 (O_841,N_24454,N_23956);
nand UO_842 (O_842,N_23804,N_22829);
and UO_843 (O_843,N_22861,N_23828);
or UO_844 (O_844,N_23511,N_24961);
nand UO_845 (O_845,N_24359,N_23888);
xnor UO_846 (O_846,N_24125,N_24664);
xor UO_847 (O_847,N_24334,N_23537);
xnor UO_848 (O_848,N_22593,N_23605);
nor UO_849 (O_849,N_24449,N_22938);
xnor UO_850 (O_850,N_24302,N_22967);
nor UO_851 (O_851,N_23495,N_23476);
or UO_852 (O_852,N_23302,N_22792);
nand UO_853 (O_853,N_22576,N_24782);
nand UO_854 (O_854,N_24514,N_23319);
or UO_855 (O_855,N_23266,N_23977);
nor UO_856 (O_856,N_24116,N_24405);
and UO_857 (O_857,N_22884,N_22877);
and UO_858 (O_858,N_24100,N_23896);
nand UO_859 (O_859,N_23822,N_24726);
nor UO_860 (O_860,N_24206,N_22834);
and UO_861 (O_861,N_24984,N_23170);
and UO_862 (O_862,N_24299,N_23405);
nor UO_863 (O_863,N_22987,N_24704);
nand UO_864 (O_864,N_24875,N_24415);
or UO_865 (O_865,N_23277,N_22977);
and UO_866 (O_866,N_23193,N_23935);
and UO_867 (O_867,N_22904,N_24612);
and UO_868 (O_868,N_23527,N_24697);
xor UO_869 (O_869,N_22502,N_23313);
or UO_870 (O_870,N_24572,N_22882);
or UO_871 (O_871,N_24154,N_24710);
and UO_872 (O_872,N_23543,N_24745);
or UO_873 (O_873,N_23647,N_23136);
xnor UO_874 (O_874,N_23231,N_23153);
nor UO_875 (O_875,N_23448,N_23209);
nor UO_876 (O_876,N_24892,N_23320);
and UO_877 (O_877,N_23604,N_23961);
nand UO_878 (O_878,N_24102,N_22741);
xnor UO_879 (O_879,N_23074,N_23742);
xnor UO_880 (O_880,N_23670,N_23990);
or UO_881 (O_881,N_23202,N_23019);
and UO_882 (O_882,N_24319,N_24595);
nand UO_883 (O_883,N_24850,N_22730);
and UO_884 (O_884,N_22700,N_24856);
xor UO_885 (O_885,N_22768,N_23958);
or UO_886 (O_886,N_23104,N_23219);
xnor UO_887 (O_887,N_24265,N_24389);
nor UO_888 (O_888,N_23849,N_24666);
nor UO_889 (O_889,N_24542,N_23222);
nor UO_890 (O_890,N_22865,N_23703);
xnor UO_891 (O_891,N_22712,N_24072);
nor UO_892 (O_892,N_23364,N_23225);
xnor UO_893 (O_893,N_24759,N_23133);
nor UO_894 (O_894,N_24687,N_23010);
and UO_895 (O_895,N_23050,N_24734);
and UO_896 (O_896,N_23368,N_24680);
xnor UO_897 (O_897,N_23454,N_22804);
or UO_898 (O_898,N_22530,N_24064);
nand UO_899 (O_899,N_22632,N_24353);
nand UO_900 (O_900,N_23965,N_22968);
xnor UO_901 (O_901,N_23852,N_24683);
xnor UO_902 (O_902,N_24148,N_23440);
nand UO_903 (O_903,N_24867,N_24393);
and UO_904 (O_904,N_24073,N_24464);
xnor UO_905 (O_905,N_22986,N_24164);
nor UO_906 (O_906,N_23337,N_24784);
nor UO_907 (O_907,N_22639,N_23903);
nand UO_908 (O_908,N_24693,N_23561);
or UO_909 (O_909,N_23238,N_23144);
nand UO_910 (O_910,N_24335,N_22912);
nor UO_911 (O_911,N_22617,N_24763);
nand UO_912 (O_912,N_23959,N_22794);
nor UO_913 (O_913,N_23926,N_24811);
xor UO_914 (O_914,N_22605,N_24028);
nor UO_915 (O_915,N_23192,N_22767);
nand UO_916 (O_916,N_24564,N_23314);
nor UO_917 (O_917,N_22615,N_23535);
nor UO_918 (O_918,N_23054,N_24910);
nand UO_919 (O_919,N_24298,N_24483);
nand UO_920 (O_920,N_23028,N_23722);
nand UO_921 (O_921,N_23391,N_23429);
and UO_922 (O_922,N_23850,N_23714);
nand UO_923 (O_923,N_24871,N_22669);
and UO_924 (O_924,N_23394,N_24876);
nor UO_925 (O_925,N_22943,N_24743);
xnor UO_926 (O_926,N_24423,N_22603);
and UO_927 (O_927,N_23927,N_23055);
xor UO_928 (O_928,N_24379,N_22821);
nor UO_929 (O_929,N_23215,N_24165);
nor UO_930 (O_930,N_23087,N_23478);
or UO_931 (O_931,N_22790,N_24789);
nand UO_932 (O_932,N_24245,N_24462);
or UO_933 (O_933,N_23882,N_23346);
xor UO_934 (O_934,N_22594,N_24329);
nor UO_935 (O_935,N_23196,N_24339);
xor UO_936 (O_936,N_23124,N_22731);
or UO_937 (O_937,N_24954,N_23158);
or UO_938 (O_938,N_23023,N_22682);
nor UO_939 (O_939,N_23991,N_24356);
nand UO_940 (O_940,N_24296,N_23743);
or UO_941 (O_941,N_23791,N_22969);
and UO_942 (O_942,N_23875,N_24699);
and UO_943 (O_943,N_22870,N_24880);
or UO_944 (O_944,N_22910,N_24705);
and UO_945 (O_945,N_24798,N_23029);
nand UO_946 (O_946,N_23098,N_22516);
and UO_947 (O_947,N_24057,N_24767);
or UO_948 (O_948,N_23413,N_23624);
nand UO_949 (O_949,N_22564,N_24305);
xnor UO_950 (O_950,N_23910,N_24145);
nand UO_951 (O_951,N_22653,N_24805);
and UO_952 (O_952,N_22825,N_24706);
xnor UO_953 (O_953,N_24422,N_23033);
or UO_954 (O_954,N_24268,N_24392);
or UO_955 (O_955,N_24243,N_23848);
or UO_956 (O_956,N_23513,N_23533);
and UO_957 (O_957,N_23399,N_23165);
nor UO_958 (O_958,N_24696,N_22805);
nand UO_959 (O_959,N_24929,N_23339);
or UO_960 (O_960,N_23423,N_22960);
or UO_961 (O_961,N_24965,N_24139);
nor UO_962 (O_962,N_24922,N_22983);
or UO_963 (O_963,N_23509,N_23190);
or UO_964 (O_964,N_24023,N_23725);
nor UO_965 (O_965,N_24920,N_24736);
xor UO_966 (O_966,N_22614,N_22609);
or UO_967 (O_967,N_24161,N_24937);
nand UO_968 (O_968,N_22716,N_24060);
nor UO_969 (O_969,N_22966,N_24303);
and UO_970 (O_970,N_24332,N_23232);
or UO_971 (O_971,N_22945,N_23009);
nor UO_972 (O_972,N_22580,N_24601);
or UO_973 (O_973,N_22998,N_24183);
or UO_974 (O_974,N_23911,N_24556);
or UO_975 (O_975,N_23786,N_23717);
and UO_976 (O_976,N_23250,N_23342);
nor UO_977 (O_977,N_24964,N_22506);
or UO_978 (O_978,N_23623,N_23949);
nand UO_979 (O_979,N_24277,N_23487);
or UO_980 (O_980,N_23335,N_24012);
or UO_981 (O_981,N_24111,N_23052);
and UO_982 (O_982,N_23504,N_24342);
nand UO_983 (O_983,N_22995,N_24896);
or UO_984 (O_984,N_22537,N_23980);
nor UO_985 (O_985,N_23420,N_23993);
and UO_986 (O_986,N_23067,N_24096);
nor UO_987 (O_987,N_24969,N_23226);
and UO_988 (O_988,N_23017,N_23272);
or UO_989 (O_989,N_23895,N_22557);
nor UO_990 (O_990,N_23255,N_23559);
or UO_991 (O_991,N_23130,N_24769);
nor UO_992 (O_992,N_24027,N_24276);
or UO_993 (O_993,N_23018,N_24052);
nor UO_994 (O_994,N_23470,N_22733);
and UO_995 (O_995,N_24702,N_23655);
xnor UO_996 (O_996,N_23411,N_23126);
xnor UO_997 (O_997,N_22501,N_24709);
and UO_998 (O_998,N_22798,N_24770);
xnor UO_999 (O_999,N_23531,N_22622);
or UO_1000 (O_1000,N_23092,N_23894);
nand UO_1001 (O_1001,N_23825,N_24584);
nand UO_1002 (O_1002,N_22802,N_22691);
nor UO_1003 (O_1003,N_23546,N_24873);
and UO_1004 (O_1004,N_22714,N_24900);
nand UO_1005 (O_1005,N_24292,N_24022);
nor UO_1006 (O_1006,N_24384,N_24047);
nand UO_1007 (O_1007,N_24259,N_24951);
xor UO_1008 (O_1008,N_24348,N_23475);
nor UO_1009 (O_1009,N_24752,N_22706);
or UO_1010 (O_1010,N_24898,N_24946);
nor UO_1011 (O_1011,N_22574,N_23733);
and UO_1012 (O_1012,N_23610,N_23344);
nand UO_1013 (O_1013,N_22925,N_23444);
xnor UO_1014 (O_1014,N_24982,N_23796);
xor UO_1015 (O_1015,N_22676,N_22607);
nand UO_1016 (O_1016,N_23590,N_24157);
or UO_1017 (O_1017,N_22743,N_24182);
or UO_1018 (O_1018,N_22726,N_24992);
nand UO_1019 (O_1019,N_24466,N_22563);
nor UO_1020 (O_1020,N_23357,N_23259);
nand UO_1021 (O_1021,N_24670,N_22857);
nor UO_1022 (O_1022,N_23668,N_22539);
nor UO_1023 (O_1023,N_24238,N_24000);
or UO_1024 (O_1024,N_23370,N_23928);
nand UO_1025 (O_1025,N_22673,N_24545);
and UO_1026 (O_1026,N_23353,N_23441);
and UO_1027 (O_1027,N_23710,N_24637);
nand UO_1028 (O_1028,N_23434,N_24314);
and UO_1029 (O_1029,N_24713,N_22562);
xnor UO_1030 (O_1030,N_24184,N_24608);
or UO_1031 (O_1031,N_24717,N_23646);
or UO_1032 (O_1032,N_24674,N_23740);
or UO_1033 (O_1033,N_23115,N_24412);
and UO_1034 (O_1034,N_24004,N_23858);
or UO_1035 (O_1035,N_24550,N_23564);
or UO_1036 (O_1036,N_23809,N_22602);
or UO_1037 (O_1037,N_22869,N_24129);
xnor UO_1038 (O_1038,N_22958,N_23214);
xor UO_1039 (O_1039,N_23323,N_24972);
and UO_1040 (O_1040,N_24039,N_24862);
or UO_1041 (O_1041,N_24214,N_23769);
or UO_1042 (O_1042,N_24284,N_22640);
or UO_1043 (O_1043,N_23997,N_22651);
and UO_1044 (O_1044,N_22851,N_24874);
or UO_1045 (O_1045,N_22612,N_22717);
and UO_1046 (O_1046,N_24499,N_23279);
nor UO_1047 (O_1047,N_23908,N_24210);
nand UO_1048 (O_1048,N_23338,N_24453);
nor UO_1049 (O_1049,N_22724,N_22941);
xor UO_1050 (O_1050,N_24657,N_23433);
or UO_1051 (O_1051,N_24902,N_24609);
nand UO_1052 (O_1052,N_24642,N_24496);
xnor UO_1053 (O_1053,N_24009,N_22903);
and UO_1054 (O_1054,N_23281,N_24046);
nand UO_1055 (O_1055,N_23178,N_24267);
nand UO_1056 (O_1056,N_23038,N_24881);
nand UO_1057 (O_1057,N_24476,N_24050);
nor UO_1058 (O_1058,N_24180,N_24253);
xor UO_1059 (O_1059,N_23081,N_22746);
and UO_1060 (O_1060,N_23555,N_23103);
nor UO_1061 (O_1061,N_22715,N_23451);
xnor UO_1062 (O_1062,N_22529,N_24062);
and UO_1063 (O_1063,N_24927,N_24787);
and UO_1064 (O_1064,N_23491,N_22838);
nand UO_1065 (O_1065,N_23901,N_24279);
nor UO_1066 (O_1066,N_23174,N_23164);
or UO_1067 (O_1067,N_24169,N_23570);
nor UO_1068 (O_1068,N_22520,N_24370);
nand UO_1069 (O_1069,N_24115,N_24797);
xnor UO_1070 (O_1070,N_23425,N_24272);
nor UO_1071 (O_1071,N_22592,N_24690);
nand UO_1072 (O_1072,N_23705,N_23082);
xor UO_1073 (O_1073,N_22973,N_24093);
and UO_1074 (O_1074,N_24649,N_22681);
or UO_1075 (O_1075,N_22771,N_22554);
xnor UO_1076 (O_1076,N_22811,N_24780);
and UO_1077 (O_1077,N_24791,N_23168);
or UO_1078 (O_1078,N_23374,N_23953);
xnor UO_1079 (O_1079,N_24603,N_24607);
or UO_1080 (O_1080,N_24925,N_22845);
xnor UO_1081 (O_1081,N_24761,N_23111);
xor UO_1082 (O_1082,N_23660,N_24257);
or UO_1083 (O_1083,N_23263,N_22569);
and UO_1084 (O_1084,N_23800,N_24576);
xor UO_1085 (O_1085,N_24097,N_23268);
nand UO_1086 (O_1086,N_23037,N_24417);
or UO_1087 (O_1087,N_22978,N_23777);
or UO_1088 (O_1088,N_24414,N_24643);
or UO_1089 (O_1089,N_24036,N_23089);
xnor UO_1090 (O_1090,N_24861,N_22544);
and UO_1091 (O_1091,N_22524,N_22525);
xor UO_1092 (O_1092,N_24024,N_24863);
nand UO_1093 (O_1093,N_22819,N_22860);
and UO_1094 (O_1094,N_23141,N_23331);
nand UO_1095 (O_1095,N_23367,N_24459);
xor UO_1096 (O_1096,N_24094,N_22627);
or UO_1097 (O_1097,N_22879,N_22898);
and UO_1098 (O_1098,N_23462,N_23780);
and UO_1099 (O_1099,N_22808,N_23762);
nor UO_1100 (O_1100,N_23060,N_24493);
or UO_1101 (O_1101,N_24368,N_24118);
nand UO_1102 (O_1102,N_24300,N_22871);
nor UO_1103 (O_1103,N_24374,N_24244);
or UO_1104 (O_1104,N_24357,N_24512);
nor UO_1105 (O_1105,N_23143,N_22782);
and UO_1106 (O_1106,N_23000,N_23508);
nor UO_1107 (O_1107,N_24762,N_24924);
xor UO_1108 (O_1108,N_23045,N_24363);
nand UO_1109 (O_1109,N_22728,N_24579);
nor UO_1110 (O_1110,N_22913,N_24540);
nor UO_1111 (O_1111,N_22864,N_24773);
nor UO_1112 (O_1112,N_23883,N_23427);
and UO_1113 (O_1113,N_24553,N_22526);
and UO_1114 (O_1114,N_23805,N_24719);
xor UO_1115 (O_1115,N_24971,N_22661);
nand UO_1116 (O_1116,N_23603,N_24622);
nand UO_1117 (O_1117,N_23436,N_24711);
or UO_1118 (O_1118,N_23833,N_23591);
or UO_1119 (O_1119,N_23459,N_23291);
nand UO_1120 (O_1120,N_23208,N_23185);
xor UO_1121 (O_1121,N_24800,N_24821);
nand UO_1122 (O_1122,N_24017,N_23971);
nand UO_1123 (O_1123,N_23932,N_24501);
and UO_1124 (O_1124,N_23744,N_22630);
nand UO_1125 (O_1125,N_24884,N_24841);
nand UO_1126 (O_1126,N_23619,N_23631);
xnor UO_1127 (O_1127,N_22722,N_24019);
nand UO_1128 (O_1128,N_24823,N_23181);
nor UO_1129 (O_1129,N_23657,N_24408);
nor UO_1130 (O_1130,N_23538,N_24508);
or UO_1131 (O_1131,N_23458,N_23416);
or UO_1132 (O_1132,N_24843,N_23068);
or UO_1133 (O_1133,N_24505,N_24953);
or UO_1134 (O_1134,N_23767,N_24818);
nand UO_1135 (O_1135,N_24737,N_23887);
and UO_1136 (O_1136,N_23352,N_24543);
or UO_1137 (O_1137,N_23414,N_23753);
xor UO_1138 (O_1138,N_24563,N_23665);
and UO_1139 (O_1139,N_23058,N_22725);
xor UO_1140 (O_1140,N_23648,N_24365);
nand UO_1141 (O_1141,N_24735,N_24008);
or UO_1142 (O_1142,N_24264,N_24274);
or UO_1143 (O_1143,N_23798,N_23654);
and UO_1144 (O_1144,N_24344,N_23765);
nor UO_1145 (O_1145,N_22579,N_22597);
nor UO_1146 (O_1146,N_23560,N_23284);
nand UO_1147 (O_1147,N_22833,N_24420);
or UO_1148 (O_1148,N_24058,N_23489);
nor UO_1149 (O_1149,N_24059,N_24170);
nand UO_1150 (O_1150,N_23437,N_24163);
and UO_1151 (O_1151,N_22689,N_24625);
nand UO_1152 (O_1152,N_23227,N_24921);
or UO_1153 (O_1153,N_24500,N_23229);
and UO_1154 (O_1154,N_23973,N_23683);
or UO_1155 (O_1155,N_23293,N_23329);
or UO_1156 (O_1156,N_24886,N_24978);
xnor UO_1157 (O_1157,N_22777,N_24507);
nand UO_1158 (O_1158,N_24487,N_24280);
nor UO_1159 (O_1159,N_22553,N_23445);
or UO_1160 (O_1160,N_23836,N_23356);
or UO_1161 (O_1161,N_24746,N_22993);
nand UO_1162 (O_1162,N_22899,N_23301);
nand UO_1163 (O_1163,N_24138,N_22820);
or UO_1164 (O_1164,N_22507,N_23821);
or UO_1165 (O_1165,N_24638,N_24205);
nand UO_1166 (O_1166,N_23571,N_23492);
xor UO_1167 (O_1167,N_24403,N_22786);
nor UO_1168 (O_1168,N_23220,N_23070);
xnor UO_1169 (O_1169,N_24887,N_23548);
nor UO_1170 (O_1170,N_24614,N_23640);
nor UO_1171 (O_1171,N_22848,N_22737);
and UO_1172 (O_1172,N_22781,N_23803);
or UO_1173 (O_1173,N_23348,N_23716);
nand UO_1174 (O_1174,N_23679,N_24425);
xor UO_1175 (O_1175,N_24018,N_24648);
or UO_1176 (O_1176,N_23384,N_24070);
and UO_1177 (O_1177,N_24430,N_23562);
or UO_1178 (O_1178,N_23006,N_24271);
nand UO_1179 (O_1179,N_24832,N_23294);
nand UO_1180 (O_1180,N_23085,N_24263);
and UO_1181 (O_1181,N_24077,N_24870);
and UO_1182 (O_1182,N_22578,N_24390);
and UO_1183 (O_1183,N_23907,N_22759);
and UO_1184 (O_1184,N_24618,N_22567);
and UO_1185 (O_1185,N_23001,N_22951);
xnor UO_1186 (O_1186,N_24909,N_23157);
nand UO_1187 (O_1187,N_24599,N_22764);
or UO_1188 (O_1188,N_23618,N_23750);
and UO_1189 (O_1189,N_24989,N_22962);
and UO_1190 (O_1190,N_22696,N_23529);
xor UO_1191 (O_1191,N_24950,N_24589);
or UO_1192 (O_1192,N_23376,N_23326);
or UO_1193 (O_1193,N_23751,N_23885);
nor UO_1194 (O_1194,N_24152,N_23305);
or UO_1195 (O_1195,N_22541,N_24538);
or UO_1196 (O_1196,N_24082,N_23403);
or UO_1197 (O_1197,N_23838,N_23792);
nor UO_1198 (O_1198,N_22624,N_24469);
and UO_1199 (O_1199,N_23402,N_23954);
and UO_1200 (O_1200,N_23481,N_24557);
nand UO_1201 (O_1201,N_23976,N_23041);
nor UO_1202 (O_1202,N_23496,N_22711);
nand UO_1203 (O_1203,N_24645,N_22586);
nor UO_1204 (O_1204,N_23138,N_23810);
and UO_1205 (O_1205,N_22911,N_23952);
nand UO_1206 (O_1206,N_22690,N_24074);
or UO_1207 (O_1207,N_24211,N_23505);
and UO_1208 (O_1208,N_23732,N_23867);
or UO_1209 (O_1209,N_24633,N_24825);
and UO_1210 (O_1210,N_24647,N_24289);
nor UO_1211 (O_1211,N_22922,N_22909);
and UO_1212 (O_1212,N_24433,N_23241);
nand UO_1213 (O_1213,N_24108,N_23228);
or UO_1214 (O_1214,N_24189,N_24935);
nand UO_1215 (O_1215,N_24411,N_23172);
and UO_1216 (O_1216,N_23892,N_24424);
xor UO_1217 (O_1217,N_23080,N_22785);
or UO_1218 (O_1218,N_23837,N_23545);
and UO_1219 (O_1219,N_23064,N_23878);
or UO_1220 (O_1220,N_22527,N_23243);
xnor UO_1221 (O_1221,N_22545,N_22511);
xor UO_1222 (O_1222,N_24151,N_24554);
and UO_1223 (O_1223,N_22558,N_23898);
nor UO_1224 (O_1224,N_23675,N_24001);
xnor UO_1225 (O_1225,N_22504,N_24122);
or UO_1226 (O_1226,N_23621,N_24451);
xor UO_1227 (O_1227,N_22692,N_23530);
or UO_1228 (O_1228,N_24593,N_23960);
nor UO_1229 (O_1229,N_23964,N_22752);
and UO_1230 (O_1230,N_23512,N_22751);
nand UO_1231 (O_1231,N_23549,N_24367);
xor UO_1232 (O_1232,N_24055,N_24227);
or UO_1233 (O_1233,N_23149,N_23731);
and UO_1234 (O_1234,N_23097,N_24631);
nand UO_1235 (O_1235,N_22921,N_24006);
or UO_1236 (O_1236,N_23361,N_24419);
or UO_1237 (O_1237,N_24801,N_24311);
or UO_1238 (O_1238,N_24974,N_24318);
nor UO_1239 (O_1239,N_23638,N_23004);
or UO_1240 (O_1240,N_24620,N_24809);
nand UO_1241 (O_1241,N_23514,N_22872);
nand UO_1242 (O_1242,N_23407,N_22859);
and UO_1243 (O_1243,N_23592,N_24448);
xor UO_1244 (O_1244,N_23970,N_23573);
nor UO_1245 (O_1245,N_23526,N_22742);
or UO_1246 (O_1246,N_22721,N_22936);
nand UO_1247 (O_1247,N_23119,N_23450);
or UO_1248 (O_1248,N_22536,N_22575);
and UO_1249 (O_1249,N_23656,N_23239);
nand UO_1250 (O_1250,N_22698,N_23658);
nand UO_1251 (O_1251,N_23647,N_24727);
xnor UO_1252 (O_1252,N_22964,N_23931);
nor UO_1253 (O_1253,N_23334,N_24040);
nand UO_1254 (O_1254,N_22671,N_22629);
nor UO_1255 (O_1255,N_24601,N_24537);
nor UO_1256 (O_1256,N_23691,N_24657);
and UO_1257 (O_1257,N_24890,N_24742);
nor UO_1258 (O_1258,N_23482,N_22985);
xnor UO_1259 (O_1259,N_22524,N_23945);
and UO_1260 (O_1260,N_22776,N_23480);
nor UO_1261 (O_1261,N_23061,N_24279);
nor UO_1262 (O_1262,N_23436,N_24575);
nor UO_1263 (O_1263,N_23019,N_24854);
and UO_1264 (O_1264,N_23628,N_22726);
or UO_1265 (O_1265,N_23098,N_23845);
nand UO_1266 (O_1266,N_23410,N_23586);
and UO_1267 (O_1267,N_24371,N_24259);
nand UO_1268 (O_1268,N_24786,N_24174);
nand UO_1269 (O_1269,N_22986,N_22921);
nand UO_1270 (O_1270,N_24624,N_22717);
nor UO_1271 (O_1271,N_24998,N_23087);
nand UO_1272 (O_1272,N_22862,N_23737);
and UO_1273 (O_1273,N_24041,N_23805);
nor UO_1274 (O_1274,N_24199,N_23289);
nand UO_1275 (O_1275,N_22985,N_24704);
nand UO_1276 (O_1276,N_22796,N_22620);
nand UO_1277 (O_1277,N_22551,N_23509);
and UO_1278 (O_1278,N_24945,N_23132);
nand UO_1279 (O_1279,N_23341,N_23334);
and UO_1280 (O_1280,N_23534,N_23101);
nor UO_1281 (O_1281,N_22668,N_24208);
nand UO_1282 (O_1282,N_23062,N_24963);
and UO_1283 (O_1283,N_23961,N_23382);
and UO_1284 (O_1284,N_23253,N_22859);
nor UO_1285 (O_1285,N_23886,N_24947);
xnor UO_1286 (O_1286,N_24707,N_22714);
xnor UO_1287 (O_1287,N_24591,N_24643);
xnor UO_1288 (O_1288,N_22715,N_23367);
nand UO_1289 (O_1289,N_22922,N_24478);
or UO_1290 (O_1290,N_23771,N_23464);
or UO_1291 (O_1291,N_24286,N_23509);
or UO_1292 (O_1292,N_23359,N_24996);
nor UO_1293 (O_1293,N_23604,N_23342);
or UO_1294 (O_1294,N_24434,N_24551);
and UO_1295 (O_1295,N_22557,N_24233);
nand UO_1296 (O_1296,N_23501,N_22724);
xnor UO_1297 (O_1297,N_22674,N_23114);
xor UO_1298 (O_1298,N_23492,N_23580);
nor UO_1299 (O_1299,N_24825,N_22912);
xor UO_1300 (O_1300,N_24939,N_22639);
and UO_1301 (O_1301,N_23467,N_22784);
nor UO_1302 (O_1302,N_23235,N_24310);
nand UO_1303 (O_1303,N_24691,N_23464);
or UO_1304 (O_1304,N_23309,N_24083);
and UO_1305 (O_1305,N_23374,N_23041);
or UO_1306 (O_1306,N_24988,N_22558);
nand UO_1307 (O_1307,N_22827,N_24216);
nor UO_1308 (O_1308,N_24208,N_22956);
or UO_1309 (O_1309,N_24554,N_22769);
nor UO_1310 (O_1310,N_22754,N_23962);
xor UO_1311 (O_1311,N_23648,N_22628);
nand UO_1312 (O_1312,N_23988,N_23838);
nand UO_1313 (O_1313,N_23769,N_24001);
or UO_1314 (O_1314,N_23948,N_23327);
xor UO_1315 (O_1315,N_24781,N_24857);
nand UO_1316 (O_1316,N_23974,N_24131);
or UO_1317 (O_1317,N_23222,N_24974);
nor UO_1318 (O_1318,N_24479,N_24935);
and UO_1319 (O_1319,N_23529,N_24995);
nand UO_1320 (O_1320,N_22670,N_23797);
nand UO_1321 (O_1321,N_22912,N_24539);
xnor UO_1322 (O_1322,N_22794,N_24473);
nor UO_1323 (O_1323,N_24020,N_24974);
nor UO_1324 (O_1324,N_23736,N_22529);
and UO_1325 (O_1325,N_24347,N_22760);
xor UO_1326 (O_1326,N_24112,N_24272);
nor UO_1327 (O_1327,N_23534,N_23255);
nand UO_1328 (O_1328,N_23194,N_23794);
or UO_1329 (O_1329,N_23892,N_22663);
xnor UO_1330 (O_1330,N_23240,N_24792);
nand UO_1331 (O_1331,N_24654,N_23064);
or UO_1332 (O_1332,N_24128,N_24733);
nor UO_1333 (O_1333,N_24506,N_24009);
xnor UO_1334 (O_1334,N_23003,N_24017);
nor UO_1335 (O_1335,N_23472,N_22983);
nand UO_1336 (O_1336,N_24967,N_24371);
xor UO_1337 (O_1337,N_23837,N_24305);
nor UO_1338 (O_1338,N_23834,N_23082);
nor UO_1339 (O_1339,N_23208,N_24943);
and UO_1340 (O_1340,N_23948,N_24419);
or UO_1341 (O_1341,N_22946,N_24776);
or UO_1342 (O_1342,N_24834,N_23172);
nor UO_1343 (O_1343,N_24233,N_23539);
xor UO_1344 (O_1344,N_23400,N_24012);
xor UO_1345 (O_1345,N_23793,N_23262);
or UO_1346 (O_1346,N_23647,N_24160);
or UO_1347 (O_1347,N_23524,N_24984);
xor UO_1348 (O_1348,N_23281,N_23872);
or UO_1349 (O_1349,N_23002,N_24788);
xor UO_1350 (O_1350,N_24053,N_24758);
xor UO_1351 (O_1351,N_22721,N_23556);
nand UO_1352 (O_1352,N_23310,N_23576);
nand UO_1353 (O_1353,N_24783,N_24575);
and UO_1354 (O_1354,N_22719,N_23072);
xor UO_1355 (O_1355,N_23278,N_24383);
nand UO_1356 (O_1356,N_23564,N_24918);
and UO_1357 (O_1357,N_24084,N_23214);
or UO_1358 (O_1358,N_23734,N_24316);
nor UO_1359 (O_1359,N_23191,N_23884);
xor UO_1360 (O_1360,N_24685,N_23402);
or UO_1361 (O_1361,N_23390,N_23830);
and UO_1362 (O_1362,N_24327,N_24282);
xnor UO_1363 (O_1363,N_23657,N_23783);
nor UO_1364 (O_1364,N_22796,N_24435);
and UO_1365 (O_1365,N_23651,N_24169);
xnor UO_1366 (O_1366,N_24084,N_23786);
or UO_1367 (O_1367,N_24803,N_23399);
xnor UO_1368 (O_1368,N_24931,N_24058);
nor UO_1369 (O_1369,N_24011,N_22534);
xor UO_1370 (O_1370,N_22816,N_23558);
xnor UO_1371 (O_1371,N_24099,N_23158);
nor UO_1372 (O_1372,N_23590,N_23143);
xnor UO_1373 (O_1373,N_23276,N_22991);
xnor UO_1374 (O_1374,N_23781,N_23239);
and UO_1375 (O_1375,N_23792,N_24223);
nand UO_1376 (O_1376,N_22763,N_23107);
xnor UO_1377 (O_1377,N_22502,N_24493);
xnor UO_1378 (O_1378,N_24387,N_23339);
xnor UO_1379 (O_1379,N_23312,N_24774);
xor UO_1380 (O_1380,N_23408,N_22917);
nor UO_1381 (O_1381,N_23623,N_24420);
xnor UO_1382 (O_1382,N_22641,N_23596);
nand UO_1383 (O_1383,N_22990,N_24199);
nand UO_1384 (O_1384,N_22933,N_23756);
nor UO_1385 (O_1385,N_23628,N_24553);
xor UO_1386 (O_1386,N_23324,N_23377);
xor UO_1387 (O_1387,N_24419,N_22503);
and UO_1388 (O_1388,N_23174,N_23959);
and UO_1389 (O_1389,N_24279,N_23467);
and UO_1390 (O_1390,N_24351,N_24447);
xnor UO_1391 (O_1391,N_23290,N_23772);
or UO_1392 (O_1392,N_23887,N_23757);
or UO_1393 (O_1393,N_23393,N_24263);
xor UO_1394 (O_1394,N_24498,N_24611);
xnor UO_1395 (O_1395,N_23230,N_24457);
and UO_1396 (O_1396,N_22515,N_22636);
and UO_1397 (O_1397,N_24483,N_24806);
xnor UO_1398 (O_1398,N_23087,N_24226);
xnor UO_1399 (O_1399,N_23056,N_22724);
xor UO_1400 (O_1400,N_24662,N_22526);
and UO_1401 (O_1401,N_24595,N_24756);
xnor UO_1402 (O_1402,N_24812,N_24775);
and UO_1403 (O_1403,N_23848,N_23725);
or UO_1404 (O_1404,N_24115,N_23848);
nand UO_1405 (O_1405,N_23180,N_23329);
nor UO_1406 (O_1406,N_24371,N_24296);
or UO_1407 (O_1407,N_24439,N_23640);
xor UO_1408 (O_1408,N_22616,N_24797);
nor UO_1409 (O_1409,N_24940,N_23773);
or UO_1410 (O_1410,N_23358,N_24630);
or UO_1411 (O_1411,N_24698,N_24213);
xnor UO_1412 (O_1412,N_23269,N_23885);
and UO_1413 (O_1413,N_22641,N_22999);
and UO_1414 (O_1414,N_24518,N_24543);
nor UO_1415 (O_1415,N_24015,N_23998);
and UO_1416 (O_1416,N_22796,N_24023);
or UO_1417 (O_1417,N_23003,N_24041);
xnor UO_1418 (O_1418,N_24085,N_22598);
nand UO_1419 (O_1419,N_24292,N_24925);
nand UO_1420 (O_1420,N_24054,N_24164);
nor UO_1421 (O_1421,N_24896,N_23740);
nand UO_1422 (O_1422,N_22757,N_23486);
nor UO_1423 (O_1423,N_24109,N_24478);
nor UO_1424 (O_1424,N_23767,N_22766);
xor UO_1425 (O_1425,N_24359,N_23726);
or UO_1426 (O_1426,N_23942,N_23357);
and UO_1427 (O_1427,N_23972,N_22868);
nand UO_1428 (O_1428,N_22844,N_24839);
nand UO_1429 (O_1429,N_23563,N_22678);
xor UO_1430 (O_1430,N_23430,N_24961);
or UO_1431 (O_1431,N_24267,N_23995);
nand UO_1432 (O_1432,N_22572,N_24158);
xor UO_1433 (O_1433,N_22593,N_24675);
and UO_1434 (O_1434,N_24850,N_22645);
and UO_1435 (O_1435,N_24316,N_24229);
nand UO_1436 (O_1436,N_23253,N_24582);
nand UO_1437 (O_1437,N_23712,N_24710);
xor UO_1438 (O_1438,N_22593,N_22518);
or UO_1439 (O_1439,N_23535,N_24782);
nor UO_1440 (O_1440,N_22811,N_24908);
nand UO_1441 (O_1441,N_24603,N_23960);
xor UO_1442 (O_1442,N_23589,N_23265);
xor UO_1443 (O_1443,N_22862,N_22770);
or UO_1444 (O_1444,N_24898,N_24784);
and UO_1445 (O_1445,N_24700,N_22536);
nand UO_1446 (O_1446,N_24911,N_22723);
nand UO_1447 (O_1447,N_23762,N_24861);
nand UO_1448 (O_1448,N_23394,N_22761);
and UO_1449 (O_1449,N_24951,N_24061);
and UO_1450 (O_1450,N_24586,N_24935);
nand UO_1451 (O_1451,N_24025,N_23589);
xnor UO_1452 (O_1452,N_23798,N_23462);
and UO_1453 (O_1453,N_24537,N_23330);
xnor UO_1454 (O_1454,N_24810,N_24306);
and UO_1455 (O_1455,N_24233,N_23070);
xor UO_1456 (O_1456,N_23340,N_24192);
and UO_1457 (O_1457,N_24404,N_23752);
nand UO_1458 (O_1458,N_23678,N_22720);
nand UO_1459 (O_1459,N_23596,N_23318);
nor UO_1460 (O_1460,N_24861,N_23242);
and UO_1461 (O_1461,N_24183,N_23854);
and UO_1462 (O_1462,N_23598,N_24007);
and UO_1463 (O_1463,N_23612,N_22620);
nand UO_1464 (O_1464,N_24982,N_23392);
or UO_1465 (O_1465,N_24525,N_24724);
or UO_1466 (O_1466,N_24842,N_22660);
or UO_1467 (O_1467,N_23091,N_24737);
or UO_1468 (O_1468,N_24767,N_23533);
and UO_1469 (O_1469,N_24376,N_23064);
and UO_1470 (O_1470,N_22846,N_24261);
nand UO_1471 (O_1471,N_23378,N_23360);
nor UO_1472 (O_1472,N_24658,N_22532);
xor UO_1473 (O_1473,N_23971,N_24891);
xnor UO_1474 (O_1474,N_22528,N_23645);
nand UO_1475 (O_1475,N_22712,N_23844);
nor UO_1476 (O_1476,N_23193,N_24893);
and UO_1477 (O_1477,N_24247,N_24582);
and UO_1478 (O_1478,N_22656,N_22813);
nor UO_1479 (O_1479,N_23312,N_24138);
and UO_1480 (O_1480,N_24029,N_23378);
and UO_1481 (O_1481,N_22769,N_24983);
nor UO_1482 (O_1482,N_24021,N_24200);
xnor UO_1483 (O_1483,N_24263,N_23799);
xnor UO_1484 (O_1484,N_22693,N_23018);
nand UO_1485 (O_1485,N_24292,N_23284);
xnor UO_1486 (O_1486,N_22682,N_22943);
xnor UO_1487 (O_1487,N_23922,N_23900);
or UO_1488 (O_1488,N_23411,N_22883);
or UO_1489 (O_1489,N_24910,N_23335);
xor UO_1490 (O_1490,N_23141,N_23632);
and UO_1491 (O_1491,N_24700,N_24235);
nor UO_1492 (O_1492,N_23241,N_22920);
nor UO_1493 (O_1493,N_24136,N_22547);
nor UO_1494 (O_1494,N_24573,N_22905);
nand UO_1495 (O_1495,N_24239,N_23902);
xor UO_1496 (O_1496,N_23052,N_23856);
xnor UO_1497 (O_1497,N_23861,N_22973);
nand UO_1498 (O_1498,N_24253,N_23802);
nand UO_1499 (O_1499,N_22563,N_23293);
nand UO_1500 (O_1500,N_23198,N_22536);
nor UO_1501 (O_1501,N_23546,N_22848);
and UO_1502 (O_1502,N_23788,N_24562);
and UO_1503 (O_1503,N_22824,N_24986);
xor UO_1504 (O_1504,N_22753,N_24984);
nand UO_1505 (O_1505,N_23107,N_22591);
nor UO_1506 (O_1506,N_24521,N_24791);
nor UO_1507 (O_1507,N_22660,N_24308);
nand UO_1508 (O_1508,N_23242,N_23562);
nor UO_1509 (O_1509,N_22528,N_24584);
and UO_1510 (O_1510,N_23230,N_23885);
or UO_1511 (O_1511,N_24597,N_24109);
nand UO_1512 (O_1512,N_23420,N_24877);
nor UO_1513 (O_1513,N_23310,N_24387);
xnor UO_1514 (O_1514,N_23852,N_23723);
and UO_1515 (O_1515,N_23294,N_22786);
nor UO_1516 (O_1516,N_23521,N_22961);
nor UO_1517 (O_1517,N_24655,N_22796);
xor UO_1518 (O_1518,N_24897,N_22631);
or UO_1519 (O_1519,N_23295,N_23967);
xnor UO_1520 (O_1520,N_22828,N_24313);
xor UO_1521 (O_1521,N_23367,N_23701);
xor UO_1522 (O_1522,N_23730,N_24976);
or UO_1523 (O_1523,N_22616,N_24399);
and UO_1524 (O_1524,N_23744,N_23834);
nor UO_1525 (O_1525,N_24358,N_23485);
xor UO_1526 (O_1526,N_24202,N_24683);
nor UO_1527 (O_1527,N_23459,N_23182);
nand UO_1528 (O_1528,N_24138,N_23089);
xnor UO_1529 (O_1529,N_24068,N_23091);
nand UO_1530 (O_1530,N_23210,N_23163);
or UO_1531 (O_1531,N_22510,N_23903);
or UO_1532 (O_1532,N_23916,N_23171);
xor UO_1533 (O_1533,N_23088,N_22862);
nor UO_1534 (O_1534,N_23697,N_23637);
and UO_1535 (O_1535,N_24235,N_23028);
xor UO_1536 (O_1536,N_24449,N_23522);
xnor UO_1537 (O_1537,N_22911,N_23875);
nand UO_1538 (O_1538,N_24927,N_23230);
nand UO_1539 (O_1539,N_24826,N_23079);
and UO_1540 (O_1540,N_23613,N_22676);
xor UO_1541 (O_1541,N_24586,N_24245);
nand UO_1542 (O_1542,N_22856,N_23639);
and UO_1543 (O_1543,N_22667,N_22540);
nand UO_1544 (O_1544,N_24953,N_22755);
nand UO_1545 (O_1545,N_24201,N_23430);
nor UO_1546 (O_1546,N_23879,N_24351);
xnor UO_1547 (O_1547,N_22844,N_24858);
nor UO_1548 (O_1548,N_23385,N_24201);
nand UO_1549 (O_1549,N_24593,N_23868);
nand UO_1550 (O_1550,N_23590,N_22946);
nor UO_1551 (O_1551,N_23186,N_24552);
nand UO_1552 (O_1552,N_24650,N_23607);
or UO_1553 (O_1553,N_23150,N_23533);
and UO_1554 (O_1554,N_24659,N_22975);
xnor UO_1555 (O_1555,N_23467,N_24599);
nand UO_1556 (O_1556,N_23671,N_23816);
nand UO_1557 (O_1557,N_24798,N_23697);
and UO_1558 (O_1558,N_23466,N_24947);
nand UO_1559 (O_1559,N_23186,N_23442);
nand UO_1560 (O_1560,N_24348,N_24102);
xor UO_1561 (O_1561,N_23455,N_23661);
nand UO_1562 (O_1562,N_22870,N_22506);
xnor UO_1563 (O_1563,N_23953,N_23838);
xnor UO_1564 (O_1564,N_22757,N_24822);
nand UO_1565 (O_1565,N_22680,N_22962);
xnor UO_1566 (O_1566,N_23259,N_24523);
xor UO_1567 (O_1567,N_24854,N_24736);
nand UO_1568 (O_1568,N_24506,N_23094);
or UO_1569 (O_1569,N_24116,N_23787);
nand UO_1570 (O_1570,N_23404,N_24032);
or UO_1571 (O_1571,N_22919,N_24793);
nor UO_1572 (O_1572,N_22917,N_22800);
and UO_1573 (O_1573,N_23202,N_23109);
nor UO_1574 (O_1574,N_23770,N_24140);
and UO_1575 (O_1575,N_22799,N_22574);
and UO_1576 (O_1576,N_23692,N_24427);
or UO_1577 (O_1577,N_23276,N_24191);
nand UO_1578 (O_1578,N_22898,N_24850);
or UO_1579 (O_1579,N_23868,N_24741);
nor UO_1580 (O_1580,N_23631,N_24257);
or UO_1581 (O_1581,N_23439,N_24614);
nor UO_1582 (O_1582,N_22613,N_22939);
nand UO_1583 (O_1583,N_23568,N_24487);
or UO_1584 (O_1584,N_24086,N_22554);
or UO_1585 (O_1585,N_24654,N_23544);
and UO_1586 (O_1586,N_23648,N_24013);
or UO_1587 (O_1587,N_22960,N_23316);
xor UO_1588 (O_1588,N_23033,N_23614);
xor UO_1589 (O_1589,N_22626,N_23126);
and UO_1590 (O_1590,N_24666,N_23222);
and UO_1591 (O_1591,N_23289,N_22937);
or UO_1592 (O_1592,N_24518,N_24612);
or UO_1593 (O_1593,N_24375,N_24158);
nor UO_1594 (O_1594,N_24633,N_23149);
and UO_1595 (O_1595,N_24530,N_23473);
nor UO_1596 (O_1596,N_23790,N_23451);
nand UO_1597 (O_1597,N_24825,N_23927);
and UO_1598 (O_1598,N_24182,N_23731);
nor UO_1599 (O_1599,N_24262,N_22964);
xor UO_1600 (O_1600,N_22911,N_24446);
and UO_1601 (O_1601,N_23368,N_23999);
and UO_1602 (O_1602,N_24960,N_22737);
and UO_1603 (O_1603,N_23105,N_24501);
or UO_1604 (O_1604,N_22793,N_23623);
nand UO_1605 (O_1605,N_24281,N_23259);
nand UO_1606 (O_1606,N_23156,N_24027);
nor UO_1607 (O_1607,N_24003,N_23329);
or UO_1608 (O_1608,N_23398,N_23313);
and UO_1609 (O_1609,N_24106,N_24824);
and UO_1610 (O_1610,N_22996,N_23167);
and UO_1611 (O_1611,N_23515,N_23367);
or UO_1612 (O_1612,N_24733,N_23742);
nor UO_1613 (O_1613,N_24790,N_24597);
nand UO_1614 (O_1614,N_23048,N_24873);
nor UO_1615 (O_1615,N_22943,N_23187);
xnor UO_1616 (O_1616,N_23090,N_24808);
nor UO_1617 (O_1617,N_23779,N_24794);
nor UO_1618 (O_1618,N_22555,N_24921);
nor UO_1619 (O_1619,N_23661,N_24298);
nand UO_1620 (O_1620,N_24625,N_24985);
or UO_1621 (O_1621,N_23214,N_24325);
or UO_1622 (O_1622,N_23765,N_23266);
xor UO_1623 (O_1623,N_22755,N_23902);
or UO_1624 (O_1624,N_24562,N_24776);
nand UO_1625 (O_1625,N_23638,N_22862);
and UO_1626 (O_1626,N_24993,N_22942);
xnor UO_1627 (O_1627,N_22832,N_23555);
nor UO_1628 (O_1628,N_23648,N_24692);
or UO_1629 (O_1629,N_23930,N_24567);
and UO_1630 (O_1630,N_22686,N_24324);
nor UO_1631 (O_1631,N_23920,N_24291);
and UO_1632 (O_1632,N_24907,N_24065);
or UO_1633 (O_1633,N_22794,N_24272);
xnor UO_1634 (O_1634,N_24831,N_23037);
nor UO_1635 (O_1635,N_24298,N_22745);
or UO_1636 (O_1636,N_23115,N_23357);
and UO_1637 (O_1637,N_24538,N_24194);
nand UO_1638 (O_1638,N_23152,N_23390);
or UO_1639 (O_1639,N_24914,N_22599);
nand UO_1640 (O_1640,N_24139,N_22895);
xor UO_1641 (O_1641,N_23411,N_22974);
or UO_1642 (O_1642,N_24773,N_23407);
or UO_1643 (O_1643,N_24415,N_24996);
xor UO_1644 (O_1644,N_23459,N_24489);
nor UO_1645 (O_1645,N_23891,N_24225);
or UO_1646 (O_1646,N_24493,N_24600);
xnor UO_1647 (O_1647,N_24300,N_22867);
xor UO_1648 (O_1648,N_24227,N_23889);
nor UO_1649 (O_1649,N_23265,N_23422);
or UO_1650 (O_1650,N_23310,N_23400);
and UO_1651 (O_1651,N_24366,N_22503);
xor UO_1652 (O_1652,N_24730,N_24675);
and UO_1653 (O_1653,N_24754,N_24556);
nor UO_1654 (O_1654,N_24952,N_24120);
or UO_1655 (O_1655,N_24088,N_23195);
or UO_1656 (O_1656,N_24155,N_23430);
or UO_1657 (O_1657,N_23334,N_23725);
and UO_1658 (O_1658,N_23436,N_22844);
xnor UO_1659 (O_1659,N_24959,N_22690);
nand UO_1660 (O_1660,N_24731,N_23423);
xnor UO_1661 (O_1661,N_23679,N_22726);
nand UO_1662 (O_1662,N_23363,N_24811);
nor UO_1663 (O_1663,N_23952,N_24070);
xnor UO_1664 (O_1664,N_24759,N_22643);
and UO_1665 (O_1665,N_24657,N_24710);
nand UO_1666 (O_1666,N_24898,N_24303);
nand UO_1667 (O_1667,N_23190,N_24847);
nor UO_1668 (O_1668,N_23768,N_24102);
nor UO_1669 (O_1669,N_22538,N_24198);
xnor UO_1670 (O_1670,N_24029,N_23082);
or UO_1671 (O_1671,N_24512,N_24619);
or UO_1672 (O_1672,N_24105,N_22873);
xnor UO_1673 (O_1673,N_23533,N_23038);
xor UO_1674 (O_1674,N_23792,N_22999);
nor UO_1675 (O_1675,N_23188,N_24295);
xor UO_1676 (O_1676,N_22508,N_23785);
nand UO_1677 (O_1677,N_23152,N_24200);
xnor UO_1678 (O_1678,N_24162,N_24842);
nand UO_1679 (O_1679,N_22785,N_24370);
and UO_1680 (O_1680,N_24355,N_24169);
and UO_1681 (O_1681,N_23676,N_23243);
or UO_1682 (O_1682,N_23927,N_23300);
or UO_1683 (O_1683,N_24376,N_22505);
and UO_1684 (O_1684,N_22713,N_24078);
nand UO_1685 (O_1685,N_23747,N_23832);
nand UO_1686 (O_1686,N_24517,N_24200);
or UO_1687 (O_1687,N_22917,N_24670);
and UO_1688 (O_1688,N_23644,N_23185);
and UO_1689 (O_1689,N_23605,N_23924);
xnor UO_1690 (O_1690,N_23659,N_24254);
and UO_1691 (O_1691,N_23054,N_22836);
nor UO_1692 (O_1692,N_24836,N_24767);
nand UO_1693 (O_1693,N_23690,N_24820);
nand UO_1694 (O_1694,N_24891,N_23403);
nand UO_1695 (O_1695,N_23940,N_22625);
or UO_1696 (O_1696,N_23145,N_22674);
and UO_1697 (O_1697,N_24132,N_23056);
nor UO_1698 (O_1698,N_23141,N_24225);
or UO_1699 (O_1699,N_24087,N_22747);
or UO_1700 (O_1700,N_24249,N_23050);
and UO_1701 (O_1701,N_22732,N_24528);
and UO_1702 (O_1702,N_23640,N_24179);
xor UO_1703 (O_1703,N_23583,N_24345);
nor UO_1704 (O_1704,N_23765,N_22678);
and UO_1705 (O_1705,N_24398,N_23042);
xor UO_1706 (O_1706,N_22997,N_23607);
or UO_1707 (O_1707,N_23497,N_23049);
nand UO_1708 (O_1708,N_23099,N_24841);
and UO_1709 (O_1709,N_23094,N_23560);
and UO_1710 (O_1710,N_22501,N_23163);
nand UO_1711 (O_1711,N_22900,N_24644);
nand UO_1712 (O_1712,N_23488,N_24845);
nand UO_1713 (O_1713,N_24352,N_24084);
nand UO_1714 (O_1714,N_22526,N_24109);
or UO_1715 (O_1715,N_23160,N_24817);
and UO_1716 (O_1716,N_23559,N_24022);
nand UO_1717 (O_1717,N_24821,N_24080);
and UO_1718 (O_1718,N_22769,N_24406);
and UO_1719 (O_1719,N_22540,N_23173);
xnor UO_1720 (O_1720,N_24315,N_23324);
and UO_1721 (O_1721,N_24929,N_23154);
nor UO_1722 (O_1722,N_23067,N_24273);
or UO_1723 (O_1723,N_24707,N_22838);
or UO_1724 (O_1724,N_24447,N_23083);
or UO_1725 (O_1725,N_23174,N_24516);
nand UO_1726 (O_1726,N_23746,N_23192);
nand UO_1727 (O_1727,N_23381,N_22638);
xor UO_1728 (O_1728,N_24072,N_24417);
or UO_1729 (O_1729,N_24928,N_23706);
or UO_1730 (O_1730,N_23396,N_23753);
nand UO_1731 (O_1731,N_24233,N_22690);
or UO_1732 (O_1732,N_23486,N_22751);
and UO_1733 (O_1733,N_24482,N_24566);
xnor UO_1734 (O_1734,N_23289,N_22526);
or UO_1735 (O_1735,N_24252,N_24361);
or UO_1736 (O_1736,N_23231,N_23295);
nor UO_1737 (O_1737,N_22745,N_24901);
xnor UO_1738 (O_1738,N_23099,N_23365);
and UO_1739 (O_1739,N_23112,N_22629);
nor UO_1740 (O_1740,N_23308,N_24722);
and UO_1741 (O_1741,N_24966,N_24273);
and UO_1742 (O_1742,N_23180,N_23513);
nand UO_1743 (O_1743,N_24082,N_22875);
or UO_1744 (O_1744,N_24991,N_24071);
or UO_1745 (O_1745,N_23813,N_23842);
nand UO_1746 (O_1746,N_23457,N_23287);
nor UO_1747 (O_1747,N_24172,N_23445);
nor UO_1748 (O_1748,N_24239,N_22578);
nor UO_1749 (O_1749,N_23244,N_24292);
and UO_1750 (O_1750,N_23767,N_23277);
nor UO_1751 (O_1751,N_22560,N_24306);
nand UO_1752 (O_1752,N_24081,N_24812);
and UO_1753 (O_1753,N_22869,N_23190);
and UO_1754 (O_1754,N_22764,N_22635);
and UO_1755 (O_1755,N_24594,N_22763);
nor UO_1756 (O_1756,N_23409,N_23296);
or UO_1757 (O_1757,N_22847,N_24552);
nand UO_1758 (O_1758,N_23051,N_23554);
xor UO_1759 (O_1759,N_22732,N_24045);
or UO_1760 (O_1760,N_23542,N_23028);
and UO_1761 (O_1761,N_23832,N_23924);
and UO_1762 (O_1762,N_22761,N_22810);
xnor UO_1763 (O_1763,N_24161,N_24909);
or UO_1764 (O_1764,N_24413,N_24448);
nor UO_1765 (O_1765,N_23657,N_24012);
or UO_1766 (O_1766,N_24547,N_24426);
nand UO_1767 (O_1767,N_22795,N_23855);
and UO_1768 (O_1768,N_24300,N_23779);
or UO_1769 (O_1769,N_22738,N_24216);
or UO_1770 (O_1770,N_23166,N_23356);
and UO_1771 (O_1771,N_24660,N_24542);
nor UO_1772 (O_1772,N_24816,N_24114);
or UO_1773 (O_1773,N_24865,N_22716);
nor UO_1774 (O_1774,N_22767,N_23457);
nand UO_1775 (O_1775,N_23068,N_22635);
and UO_1776 (O_1776,N_24682,N_24667);
and UO_1777 (O_1777,N_24879,N_23688);
xnor UO_1778 (O_1778,N_23784,N_24432);
nand UO_1779 (O_1779,N_24236,N_22552);
nand UO_1780 (O_1780,N_22777,N_24527);
xor UO_1781 (O_1781,N_23745,N_23316);
xor UO_1782 (O_1782,N_23557,N_24407);
and UO_1783 (O_1783,N_22544,N_24706);
nor UO_1784 (O_1784,N_23433,N_22898);
or UO_1785 (O_1785,N_23298,N_24438);
or UO_1786 (O_1786,N_24264,N_22863);
or UO_1787 (O_1787,N_23017,N_22872);
and UO_1788 (O_1788,N_24222,N_22716);
nand UO_1789 (O_1789,N_24057,N_23874);
nor UO_1790 (O_1790,N_22743,N_23001);
xnor UO_1791 (O_1791,N_22563,N_24499);
nor UO_1792 (O_1792,N_24386,N_24455);
or UO_1793 (O_1793,N_24545,N_23633);
and UO_1794 (O_1794,N_23626,N_22533);
and UO_1795 (O_1795,N_24119,N_22876);
or UO_1796 (O_1796,N_24931,N_23202);
or UO_1797 (O_1797,N_23534,N_23140);
nor UO_1798 (O_1798,N_24157,N_22662);
nand UO_1799 (O_1799,N_22992,N_24720);
or UO_1800 (O_1800,N_23048,N_23152);
xnor UO_1801 (O_1801,N_24079,N_24402);
xor UO_1802 (O_1802,N_24161,N_22986);
xnor UO_1803 (O_1803,N_24955,N_22560);
nor UO_1804 (O_1804,N_24030,N_23966);
and UO_1805 (O_1805,N_24154,N_24675);
nor UO_1806 (O_1806,N_23929,N_22821);
nand UO_1807 (O_1807,N_22735,N_24411);
nand UO_1808 (O_1808,N_24611,N_23877);
nor UO_1809 (O_1809,N_22568,N_22677);
xor UO_1810 (O_1810,N_23366,N_24092);
xor UO_1811 (O_1811,N_24806,N_24911);
xnor UO_1812 (O_1812,N_23853,N_24625);
or UO_1813 (O_1813,N_24074,N_24465);
and UO_1814 (O_1814,N_24014,N_24321);
xnor UO_1815 (O_1815,N_23689,N_24336);
or UO_1816 (O_1816,N_23592,N_22812);
nand UO_1817 (O_1817,N_24336,N_23562);
xor UO_1818 (O_1818,N_24150,N_24857);
nor UO_1819 (O_1819,N_22655,N_22563);
or UO_1820 (O_1820,N_24983,N_24539);
nor UO_1821 (O_1821,N_23026,N_23340);
and UO_1822 (O_1822,N_23306,N_23878);
or UO_1823 (O_1823,N_23306,N_23616);
and UO_1824 (O_1824,N_23161,N_23701);
nor UO_1825 (O_1825,N_23613,N_24003);
or UO_1826 (O_1826,N_24871,N_22618);
nor UO_1827 (O_1827,N_22862,N_24579);
or UO_1828 (O_1828,N_23224,N_24503);
xnor UO_1829 (O_1829,N_22757,N_24012);
and UO_1830 (O_1830,N_24426,N_24856);
or UO_1831 (O_1831,N_22758,N_24922);
and UO_1832 (O_1832,N_23354,N_23517);
and UO_1833 (O_1833,N_23876,N_22690);
nor UO_1834 (O_1834,N_23921,N_24325);
or UO_1835 (O_1835,N_23218,N_22904);
nand UO_1836 (O_1836,N_22833,N_24094);
or UO_1837 (O_1837,N_24967,N_23296);
xnor UO_1838 (O_1838,N_23720,N_24289);
nor UO_1839 (O_1839,N_23730,N_24277);
xor UO_1840 (O_1840,N_23922,N_24707);
or UO_1841 (O_1841,N_23417,N_23508);
or UO_1842 (O_1842,N_23807,N_22790);
or UO_1843 (O_1843,N_23371,N_22506);
nand UO_1844 (O_1844,N_23231,N_24722);
and UO_1845 (O_1845,N_24634,N_24149);
nand UO_1846 (O_1846,N_23363,N_23740);
and UO_1847 (O_1847,N_22858,N_24759);
nor UO_1848 (O_1848,N_24836,N_24107);
xor UO_1849 (O_1849,N_22938,N_24709);
nor UO_1850 (O_1850,N_23405,N_22517);
xor UO_1851 (O_1851,N_23991,N_24649);
or UO_1852 (O_1852,N_22825,N_24504);
or UO_1853 (O_1853,N_23461,N_22811);
and UO_1854 (O_1854,N_23884,N_24295);
nor UO_1855 (O_1855,N_24803,N_24837);
xnor UO_1856 (O_1856,N_23600,N_24925);
and UO_1857 (O_1857,N_22823,N_24776);
and UO_1858 (O_1858,N_22700,N_23659);
nor UO_1859 (O_1859,N_23302,N_24188);
nand UO_1860 (O_1860,N_24143,N_24205);
nor UO_1861 (O_1861,N_23858,N_23486);
and UO_1862 (O_1862,N_24085,N_24612);
and UO_1863 (O_1863,N_24472,N_24224);
xnor UO_1864 (O_1864,N_24704,N_22755);
nand UO_1865 (O_1865,N_22847,N_24581);
nor UO_1866 (O_1866,N_23449,N_24566);
nor UO_1867 (O_1867,N_24659,N_24916);
nand UO_1868 (O_1868,N_24848,N_24261);
nor UO_1869 (O_1869,N_22907,N_24876);
xnor UO_1870 (O_1870,N_22564,N_23358);
xor UO_1871 (O_1871,N_23764,N_22968);
xnor UO_1872 (O_1872,N_22983,N_22930);
nor UO_1873 (O_1873,N_23523,N_23918);
or UO_1874 (O_1874,N_24372,N_24506);
and UO_1875 (O_1875,N_24545,N_23550);
xor UO_1876 (O_1876,N_24675,N_22732);
nor UO_1877 (O_1877,N_23004,N_23596);
or UO_1878 (O_1878,N_24230,N_22985);
nor UO_1879 (O_1879,N_22815,N_23169);
nand UO_1880 (O_1880,N_22542,N_22990);
nand UO_1881 (O_1881,N_24451,N_24533);
or UO_1882 (O_1882,N_23015,N_22942);
xor UO_1883 (O_1883,N_24099,N_23805);
nand UO_1884 (O_1884,N_22614,N_22987);
xnor UO_1885 (O_1885,N_24370,N_24323);
or UO_1886 (O_1886,N_24925,N_24717);
nand UO_1887 (O_1887,N_23233,N_24079);
or UO_1888 (O_1888,N_24889,N_24490);
nand UO_1889 (O_1889,N_23549,N_23109);
or UO_1890 (O_1890,N_23919,N_23089);
nand UO_1891 (O_1891,N_22767,N_24817);
xor UO_1892 (O_1892,N_23405,N_24497);
nand UO_1893 (O_1893,N_23556,N_23534);
or UO_1894 (O_1894,N_23858,N_23113);
xor UO_1895 (O_1895,N_22873,N_22646);
nor UO_1896 (O_1896,N_24367,N_23452);
xor UO_1897 (O_1897,N_22980,N_23260);
and UO_1898 (O_1898,N_23397,N_24681);
nand UO_1899 (O_1899,N_24593,N_23880);
nor UO_1900 (O_1900,N_24176,N_23593);
xor UO_1901 (O_1901,N_24197,N_22688);
xor UO_1902 (O_1902,N_24458,N_24672);
xnor UO_1903 (O_1903,N_24668,N_23187);
xnor UO_1904 (O_1904,N_24642,N_23305);
nand UO_1905 (O_1905,N_23005,N_22856);
nor UO_1906 (O_1906,N_23612,N_23289);
nor UO_1907 (O_1907,N_22611,N_24748);
nor UO_1908 (O_1908,N_24167,N_24666);
nand UO_1909 (O_1909,N_22939,N_23649);
nor UO_1910 (O_1910,N_24221,N_23880);
xnor UO_1911 (O_1911,N_23006,N_23629);
or UO_1912 (O_1912,N_22580,N_24020);
xnor UO_1913 (O_1913,N_24435,N_22673);
or UO_1914 (O_1914,N_22583,N_23018);
xor UO_1915 (O_1915,N_23033,N_23057);
nand UO_1916 (O_1916,N_24182,N_23596);
nand UO_1917 (O_1917,N_23375,N_24742);
nand UO_1918 (O_1918,N_22563,N_23659);
xor UO_1919 (O_1919,N_24336,N_24342);
xnor UO_1920 (O_1920,N_23081,N_24704);
xor UO_1921 (O_1921,N_24267,N_24399);
and UO_1922 (O_1922,N_22608,N_24902);
nor UO_1923 (O_1923,N_24136,N_24539);
nand UO_1924 (O_1924,N_24995,N_23488);
or UO_1925 (O_1925,N_24069,N_23684);
nor UO_1926 (O_1926,N_22659,N_24949);
xor UO_1927 (O_1927,N_23951,N_23771);
and UO_1928 (O_1928,N_23964,N_23919);
nand UO_1929 (O_1929,N_23144,N_23274);
and UO_1930 (O_1930,N_23680,N_24244);
nand UO_1931 (O_1931,N_23323,N_24422);
nand UO_1932 (O_1932,N_22715,N_22738);
nand UO_1933 (O_1933,N_24255,N_24495);
nand UO_1934 (O_1934,N_23141,N_23534);
nor UO_1935 (O_1935,N_23842,N_24750);
xor UO_1936 (O_1936,N_24516,N_22804);
nor UO_1937 (O_1937,N_23215,N_23183);
or UO_1938 (O_1938,N_23332,N_23480);
nor UO_1939 (O_1939,N_22692,N_23954);
nor UO_1940 (O_1940,N_23841,N_24536);
xnor UO_1941 (O_1941,N_22972,N_23731);
nand UO_1942 (O_1942,N_24911,N_24119);
xnor UO_1943 (O_1943,N_24320,N_24639);
or UO_1944 (O_1944,N_24561,N_23817);
and UO_1945 (O_1945,N_23687,N_22717);
nor UO_1946 (O_1946,N_23321,N_23047);
nor UO_1947 (O_1947,N_23740,N_22890);
nor UO_1948 (O_1948,N_23415,N_24784);
xor UO_1949 (O_1949,N_22630,N_24555);
nor UO_1950 (O_1950,N_23376,N_24935);
or UO_1951 (O_1951,N_24743,N_23025);
and UO_1952 (O_1952,N_24494,N_23062);
xnor UO_1953 (O_1953,N_24503,N_23237);
and UO_1954 (O_1954,N_24086,N_24022);
or UO_1955 (O_1955,N_22961,N_23908);
or UO_1956 (O_1956,N_23655,N_24974);
and UO_1957 (O_1957,N_24729,N_23500);
xnor UO_1958 (O_1958,N_24503,N_23426);
and UO_1959 (O_1959,N_23254,N_24989);
xnor UO_1960 (O_1960,N_22515,N_24657);
xnor UO_1961 (O_1961,N_24127,N_24766);
or UO_1962 (O_1962,N_24263,N_22738);
nand UO_1963 (O_1963,N_23307,N_23244);
nor UO_1964 (O_1964,N_23473,N_24291);
xnor UO_1965 (O_1965,N_22640,N_24545);
nand UO_1966 (O_1966,N_22576,N_24245);
xnor UO_1967 (O_1967,N_24068,N_24105);
nand UO_1968 (O_1968,N_23459,N_23185);
or UO_1969 (O_1969,N_23391,N_23479);
nand UO_1970 (O_1970,N_24243,N_22888);
or UO_1971 (O_1971,N_23409,N_23954);
nand UO_1972 (O_1972,N_22583,N_24227);
or UO_1973 (O_1973,N_22800,N_23363);
nor UO_1974 (O_1974,N_23071,N_24726);
or UO_1975 (O_1975,N_23646,N_23633);
xnor UO_1976 (O_1976,N_22589,N_22991);
xnor UO_1977 (O_1977,N_24932,N_22790);
and UO_1978 (O_1978,N_24906,N_24963);
and UO_1979 (O_1979,N_23086,N_23493);
xor UO_1980 (O_1980,N_23763,N_24495);
nand UO_1981 (O_1981,N_23610,N_24784);
xnor UO_1982 (O_1982,N_23129,N_23314);
nor UO_1983 (O_1983,N_24936,N_24459);
nand UO_1984 (O_1984,N_22628,N_24068);
xnor UO_1985 (O_1985,N_22903,N_24768);
or UO_1986 (O_1986,N_24995,N_24949);
and UO_1987 (O_1987,N_23358,N_23855);
nor UO_1988 (O_1988,N_22761,N_23611);
or UO_1989 (O_1989,N_23707,N_24004);
nand UO_1990 (O_1990,N_24373,N_23812);
and UO_1991 (O_1991,N_24919,N_22692);
nand UO_1992 (O_1992,N_24369,N_24763);
and UO_1993 (O_1993,N_24757,N_24957);
nor UO_1994 (O_1994,N_24837,N_24240);
nand UO_1995 (O_1995,N_24485,N_24730);
nand UO_1996 (O_1996,N_23707,N_22560);
nor UO_1997 (O_1997,N_24906,N_24128);
nand UO_1998 (O_1998,N_22524,N_24485);
or UO_1999 (O_1999,N_23712,N_22853);
or UO_2000 (O_2000,N_22761,N_22725);
nor UO_2001 (O_2001,N_23069,N_22501);
and UO_2002 (O_2002,N_24430,N_23701);
nand UO_2003 (O_2003,N_24803,N_23957);
or UO_2004 (O_2004,N_22517,N_23788);
and UO_2005 (O_2005,N_23063,N_23897);
or UO_2006 (O_2006,N_23555,N_24286);
nor UO_2007 (O_2007,N_23155,N_24513);
nand UO_2008 (O_2008,N_24473,N_24144);
nor UO_2009 (O_2009,N_23058,N_24936);
or UO_2010 (O_2010,N_22920,N_23262);
and UO_2011 (O_2011,N_23259,N_23474);
nand UO_2012 (O_2012,N_23434,N_24724);
xnor UO_2013 (O_2013,N_23585,N_23032);
nor UO_2014 (O_2014,N_24050,N_22996);
and UO_2015 (O_2015,N_24268,N_23268);
nor UO_2016 (O_2016,N_23301,N_24648);
nand UO_2017 (O_2017,N_22973,N_24459);
nor UO_2018 (O_2018,N_23225,N_24860);
nor UO_2019 (O_2019,N_22916,N_23386);
nand UO_2020 (O_2020,N_23875,N_23052);
and UO_2021 (O_2021,N_23495,N_23964);
nor UO_2022 (O_2022,N_24555,N_24161);
or UO_2023 (O_2023,N_24456,N_24263);
nand UO_2024 (O_2024,N_22667,N_23393);
nand UO_2025 (O_2025,N_23059,N_22789);
nand UO_2026 (O_2026,N_23890,N_22735);
and UO_2027 (O_2027,N_24401,N_22915);
or UO_2028 (O_2028,N_24390,N_24283);
nor UO_2029 (O_2029,N_23002,N_24965);
or UO_2030 (O_2030,N_23045,N_23254);
xnor UO_2031 (O_2031,N_23848,N_24001);
nand UO_2032 (O_2032,N_24668,N_24557);
xor UO_2033 (O_2033,N_24124,N_24603);
and UO_2034 (O_2034,N_24660,N_23890);
or UO_2035 (O_2035,N_23645,N_24059);
nor UO_2036 (O_2036,N_23416,N_23301);
xnor UO_2037 (O_2037,N_22969,N_24884);
nand UO_2038 (O_2038,N_23827,N_22810);
nand UO_2039 (O_2039,N_22756,N_24834);
xor UO_2040 (O_2040,N_24706,N_23185);
and UO_2041 (O_2041,N_24091,N_22500);
xor UO_2042 (O_2042,N_24191,N_23966);
nor UO_2043 (O_2043,N_23500,N_24206);
and UO_2044 (O_2044,N_23337,N_24426);
nand UO_2045 (O_2045,N_24876,N_22549);
or UO_2046 (O_2046,N_22794,N_23666);
nand UO_2047 (O_2047,N_23376,N_22872);
and UO_2048 (O_2048,N_24640,N_23285);
nand UO_2049 (O_2049,N_23880,N_24344);
nand UO_2050 (O_2050,N_24654,N_24352);
nand UO_2051 (O_2051,N_23583,N_23181);
xor UO_2052 (O_2052,N_23770,N_24165);
nor UO_2053 (O_2053,N_22881,N_23649);
nor UO_2054 (O_2054,N_24169,N_24806);
and UO_2055 (O_2055,N_24574,N_23131);
or UO_2056 (O_2056,N_23244,N_23409);
or UO_2057 (O_2057,N_24650,N_24645);
xnor UO_2058 (O_2058,N_23179,N_22502);
and UO_2059 (O_2059,N_23773,N_23678);
nand UO_2060 (O_2060,N_23173,N_22514);
nor UO_2061 (O_2061,N_22828,N_23321);
nor UO_2062 (O_2062,N_24234,N_22622);
nor UO_2063 (O_2063,N_24619,N_24811);
nand UO_2064 (O_2064,N_22586,N_22695);
and UO_2065 (O_2065,N_22986,N_23097);
xor UO_2066 (O_2066,N_23339,N_23425);
xnor UO_2067 (O_2067,N_22616,N_22916);
xnor UO_2068 (O_2068,N_22678,N_23059);
nand UO_2069 (O_2069,N_22776,N_23560);
or UO_2070 (O_2070,N_23813,N_24718);
nand UO_2071 (O_2071,N_24006,N_23929);
or UO_2072 (O_2072,N_24210,N_24603);
nand UO_2073 (O_2073,N_24428,N_24312);
nand UO_2074 (O_2074,N_23853,N_24650);
and UO_2075 (O_2075,N_24021,N_23029);
or UO_2076 (O_2076,N_23621,N_23984);
nand UO_2077 (O_2077,N_24172,N_23212);
nand UO_2078 (O_2078,N_24786,N_22694);
nor UO_2079 (O_2079,N_22602,N_24910);
nor UO_2080 (O_2080,N_22716,N_23791);
xor UO_2081 (O_2081,N_23466,N_23036);
or UO_2082 (O_2082,N_23191,N_22905);
or UO_2083 (O_2083,N_23646,N_24232);
nor UO_2084 (O_2084,N_23975,N_24630);
and UO_2085 (O_2085,N_23759,N_24218);
xnor UO_2086 (O_2086,N_22807,N_23269);
xor UO_2087 (O_2087,N_24441,N_22780);
or UO_2088 (O_2088,N_22955,N_24497);
and UO_2089 (O_2089,N_24395,N_24009);
nand UO_2090 (O_2090,N_23685,N_22764);
or UO_2091 (O_2091,N_23253,N_24417);
nor UO_2092 (O_2092,N_22631,N_24437);
nor UO_2093 (O_2093,N_24807,N_23181);
and UO_2094 (O_2094,N_24876,N_22861);
or UO_2095 (O_2095,N_24148,N_24961);
nand UO_2096 (O_2096,N_23335,N_24735);
nand UO_2097 (O_2097,N_24532,N_24528);
nand UO_2098 (O_2098,N_24712,N_24180);
xor UO_2099 (O_2099,N_23992,N_23202);
or UO_2100 (O_2100,N_22512,N_23529);
nand UO_2101 (O_2101,N_22759,N_23115);
and UO_2102 (O_2102,N_23983,N_23962);
nor UO_2103 (O_2103,N_22640,N_23455);
nor UO_2104 (O_2104,N_24876,N_23663);
nand UO_2105 (O_2105,N_24081,N_22680);
nand UO_2106 (O_2106,N_24551,N_23754);
nor UO_2107 (O_2107,N_24982,N_24432);
xnor UO_2108 (O_2108,N_24414,N_23915);
nand UO_2109 (O_2109,N_24626,N_23549);
nor UO_2110 (O_2110,N_23566,N_24380);
nor UO_2111 (O_2111,N_23407,N_23277);
nor UO_2112 (O_2112,N_23856,N_24020);
nand UO_2113 (O_2113,N_23456,N_24165);
nand UO_2114 (O_2114,N_24577,N_24329);
or UO_2115 (O_2115,N_24174,N_23505);
nand UO_2116 (O_2116,N_23492,N_23380);
or UO_2117 (O_2117,N_24316,N_24794);
and UO_2118 (O_2118,N_24812,N_23569);
nor UO_2119 (O_2119,N_23423,N_24678);
nand UO_2120 (O_2120,N_23372,N_22533);
and UO_2121 (O_2121,N_23278,N_23123);
or UO_2122 (O_2122,N_24240,N_23647);
nor UO_2123 (O_2123,N_22977,N_23044);
nand UO_2124 (O_2124,N_23916,N_24249);
nor UO_2125 (O_2125,N_23182,N_22982);
or UO_2126 (O_2126,N_23690,N_23591);
nor UO_2127 (O_2127,N_22836,N_23373);
nor UO_2128 (O_2128,N_22968,N_24554);
nand UO_2129 (O_2129,N_22636,N_24733);
and UO_2130 (O_2130,N_23423,N_24663);
nand UO_2131 (O_2131,N_23294,N_24198);
or UO_2132 (O_2132,N_23396,N_23164);
xor UO_2133 (O_2133,N_22829,N_24805);
xor UO_2134 (O_2134,N_23409,N_24779);
or UO_2135 (O_2135,N_24295,N_24806);
and UO_2136 (O_2136,N_24770,N_24665);
nand UO_2137 (O_2137,N_23483,N_23167);
nor UO_2138 (O_2138,N_22897,N_24500);
and UO_2139 (O_2139,N_24360,N_22603);
nand UO_2140 (O_2140,N_24387,N_24580);
nand UO_2141 (O_2141,N_23250,N_24359);
or UO_2142 (O_2142,N_24725,N_23590);
nand UO_2143 (O_2143,N_23939,N_24108);
xnor UO_2144 (O_2144,N_23105,N_24904);
and UO_2145 (O_2145,N_23992,N_22818);
or UO_2146 (O_2146,N_24957,N_23542);
nand UO_2147 (O_2147,N_22890,N_23122);
xor UO_2148 (O_2148,N_23964,N_22552);
and UO_2149 (O_2149,N_23746,N_23512);
nand UO_2150 (O_2150,N_24256,N_23586);
xor UO_2151 (O_2151,N_24188,N_23519);
xnor UO_2152 (O_2152,N_24803,N_24844);
nor UO_2153 (O_2153,N_22654,N_23050);
nor UO_2154 (O_2154,N_23520,N_23992);
and UO_2155 (O_2155,N_24974,N_23290);
or UO_2156 (O_2156,N_23321,N_22932);
and UO_2157 (O_2157,N_22703,N_24029);
nand UO_2158 (O_2158,N_24957,N_24771);
nor UO_2159 (O_2159,N_24252,N_23473);
xor UO_2160 (O_2160,N_24361,N_23041);
and UO_2161 (O_2161,N_22997,N_24364);
or UO_2162 (O_2162,N_23823,N_23837);
xor UO_2163 (O_2163,N_24384,N_23323);
xnor UO_2164 (O_2164,N_23131,N_24087);
or UO_2165 (O_2165,N_23595,N_23404);
xor UO_2166 (O_2166,N_24622,N_24965);
nand UO_2167 (O_2167,N_22948,N_23924);
nor UO_2168 (O_2168,N_24947,N_22711);
nor UO_2169 (O_2169,N_23990,N_24172);
or UO_2170 (O_2170,N_24568,N_24450);
xnor UO_2171 (O_2171,N_23380,N_23809);
nor UO_2172 (O_2172,N_23390,N_22591);
nor UO_2173 (O_2173,N_22562,N_23406);
or UO_2174 (O_2174,N_24181,N_23726);
or UO_2175 (O_2175,N_23048,N_24062);
nor UO_2176 (O_2176,N_22975,N_22942);
or UO_2177 (O_2177,N_22901,N_23280);
xor UO_2178 (O_2178,N_24190,N_22922);
xnor UO_2179 (O_2179,N_24521,N_24708);
xnor UO_2180 (O_2180,N_22750,N_24997);
or UO_2181 (O_2181,N_22851,N_23330);
nand UO_2182 (O_2182,N_24952,N_23095);
nand UO_2183 (O_2183,N_23458,N_24705);
xor UO_2184 (O_2184,N_23346,N_23401);
and UO_2185 (O_2185,N_23341,N_24307);
and UO_2186 (O_2186,N_23322,N_23152);
nor UO_2187 (O_2187,N_22901,N_23292);
and UO_2188 (O_2188,N_23798,N_23120);
nand UO_2189 (O_2189,N_23784,N_22753);
xor UO_2190 (O_2190,N_24377,N_23614);
and UO_2191 (O_2191,N_24083,N_23798);
xnor UO_2192 (O_2192,N_23581,N_23584);
nor UO_2193 (O_2193,N_22639,N_24299);
or UO_2194 (O_2194,N_23306,N_23922);
nor UO_2195 (O_2195,N_24620,N_23597);
nor UO_2196 (O_2196,N_23035,N_24457);
xnor UO_2197 (O_2197,N_24131,N_22817);
nor UO_2198 (O_2198,N_24124,N_24418);
xnor UO_2199 (O_2199,N_24565,N_24940);
and UO_2200 (O_2200,N_24695,N_23900);
and UO_2201 (O_2201,N_23788,N_24564);
nor UO_2202 (O_2202,N_24157,N_24700);
nand UO_2203 (O_2203,N_22805,N_23529);
xor UO_2204 (O_2204,N_23493,N_23398);
or UO_2205 (O_2205,N_23378,N_24439);
nor UO_2206 (O_2206,N_22950,N_23947);
nand UO_2207 (O_2207,N_22510,N_22994);
or UO_2208 (O_2208,N_23333,N_23972);
and UO_2209 (O_2209,N_23241,N_24301);
xnor UO_2210 (O_2210,N_23061,N_24518);
or UO_2211 (O_2211,N_24187,N_23236);
nor UO_2212 (O_2212,N_24719,N_22905);
nor UO_2213 (O_2213,N_23840,N_23158);
and UO_2214 (O_2214,N_22990,N_24881);
and UO_2215 (O_2215,N_23108,N_23464);
nor UO_2216 (O_2216,N_23189,N_24603);
and UO_2217 (O_2217,N_23147,N_24814);
and UO_2218 (O_2218,N_24058,N_23548);
nand UO_2219 (O_2219,N_23506,N_24637);
nor UO_2220 (O_2220,N_23841,N_24776);
or UO_2221 (O_2221,N_24589,N_23779);
and UO_2222 (O_2222,N_24086,N_22585);
xnor UO_2223 (O_2223,N_22599,N_22860);
nand UO_2224 (O_2224,N_24378,N_23938);
nand UO_2225 (O_2225,N_24933,N_23386);
nand UO_2226 (O_2226,N_23822,N_23319);
nor UO_2227 (O_2227,N_24551,N_24478);
nor UO_2228 (O_2228,N_24190,N_23451);
xnor UO_2229 (O_2229,N_24092,N_23774);
or UO_2230 (O_2230,N_24180,N_23820);
or UO_2231 (O_2231,N_23495,N_23405);
nand UO_2232 (O_2232,N_24543,N_24205);
or UO_2233 (O_2233,N_22723,N_23849);
xor UO_2234 (O_2234,N_24800,N_23194);
nor UO_2235 (O_2235,N_22608,N_23047);
nor UO_2236 (O_2236,N_24231,N_22831);
nand UO_2237 (O_2237,N_23882,N_23630);
nand UO_2238 (O_2238,N_23402,N_23897);
or UO_2239 (O_2239,N_24652,N_23697);
nand UO_2240 (O_2240,N_23644,N_24488);
or UO_2241 (O_2241,N_23613,N_24986);
or UO_2242 (O_2242,N_23347,N_24833);
and UO_2243 (O_2243,N_22815,N_23297);
nor UO_2244 (O_2244,N_24377,N_23476);
or UO_2245 (O_2245,N_23878,N_23809);
and UO_2246 (O_2246,N_23264,N_23978);
and UO_2247 (O_2247,N_24046,N_22717);
nor UO_2248 (O_2248,N_24724,N_22798);
or UO_2249 (O_2249,N_23992,N_23760);
nor UO_2250 (O_2250,N_23106,N_24680);
or UO_2251 (O_2251,N_22580,N_22952);
nand UO_2252 (O_2252,N_22648,N_24071);
and UO_2253 (O_2253,N_24335,N_23892);
or UO_2254 (O_2254,N_24507,N_24609);
nand UO_2255 (O_2255,N_24615,N_24751);
nor UO_2256 (O_2256,N_23919,N_23786);
and UO_2257 (O_2257,N_22752,N_22906);
or UO_2258 (O_2258,N_24759,N_23145);
and UO_2259 (O_2259,N_24926,N_23777);
nand UO_2260 (O_2260,N_22826,N_24257);
xnor UO_2261 (O_2261,N_24703,N_22853);
or UO_2262 (O_2262,N_23111,N_22557);
and UO_2263 (O_2263,N_23908,N_22520);
and UO_2264 (O_2264,N_23653,N_23144);
nand UO_2265 (O_2265,N_23969,N_22525);
nor UO_2266 (O_2266,N_22985,N_23053);
nand UO_2267 (O_2267,N_24082,N_23590);
and UO_2268 (O_2268,N_24990,N_24240);
or UO_2269 (O_2269,N_24748,N_23644);
and UO_2270 (O_2270,N_24127,N_23216);
and UO_2271 (O_2271,N_22663,N_24137);
nand UO_2272 (O_2272,N_23676,N_24039);
nand UO_2273 (O_2273,N_23623,N_23052);
xor UO_2274 (O_2274,N_23322,N_24170);
nor UO_2275 (O_2275,N_23685,N_24530);
and UO_2276 (O_2276,N_23919,N_22557);
or UO_2277 (O_2277,N_24710,N_24927);
xnor UO_2278 (O_2278,N_23107,N_23325);
nor UO_2279 (O_2279,N_24423,N_22524);
or UO_2280 (O_2280,N_23412,N_23210);
nor UO_2281 (O_2281,N_23412,N_23215);
and UO_2282 (O_2282,N_23345,N_24372);
nor UO_2283 (O_2283,N_24314,N_23156);
nor UO_2284 (O_2284,N_24436,N_23197);
nor UO_2285 (O_2285,N_24659,N_23739);
nand UO_2286 (O_2286,N_23246,N_23177);
nor UO_2287 (O_2287,N_22893,N_23410);
xnor UO_2288 (O_2288,N_24273,N_23509);
nor UO_2289 (O_2289,N_23698,N_22650);
or UO_2290 (O_2290,N_24836,N_24704);
xor UO_2291 (O_2291,N_23123,N_24661);
or UO_2292 (O_2292,N_23255,N_22605);
nor UO_2293 (O_2293,N_23745,N_22923);
nand UO_2294 (O_2294,N_22574,N_24367);
nand UO_2295 (O_2295,N_23023,N_23076);
nor UO_2296 (O_2296,N_24173,N_24670);
xor UO_2297 (O_2297,N_23033,N_23143);
nand UO_2298 (O_2298,N_22788,N_23585);
nor UO_2299 (O_2299,N_22973,N_22937);
xnor UO_2300 (O_2300,N_23727,N_22777);
nor UO_2301 (O_2301,N_23576,N_23476);
nor UO_2302 (O_2302,N_24435,N_24759);
nor UO_2303 (O_2303,N_23765,N_24855);
or UO_2304 (O_2304,N_24897,N_23590);
nor UO_2305 (O_2305,N_22803,N_23273);
and UO_2306 (O_2306,N_23820,N_23348);
nand UO_2307 (O_2307,N_22566,N_23926);
nand UO_2308 (O_2308,N_24903,N_23057);
xnor UO_2309 (O_2309,N_23031,N_23293);
nor UO_2310 (O_2310,N_24448,N_23238);
nor UO_2311 (O_2311,N_24469,N_24560);
and UO_2312 (O_2312,N_24620,N_23156);
and UO_2313 (O_2313,N_22519,N_22628);
nand UO_2314 (O_2314,N_24392,N_22840);
and UO_2315 (O_2315,N_24031,N_23929);
xnor UO_2316 (O_2316,N_24611,N_22763);
and UO_2317 (O_2317,N_23687,N_22688);
or UO_2318 (O_2318,N_24291,N_23625);
and UO_2319 (O_2319,N_24508,N_23915);
or UO_2320 (O_2320,N_24342,N_24499);
and UO_2321 (O_2321,N_24954,N_24490);
or UO_2322 (O_2322,N_22973,N_23721);
xor UO_2323 (O_2323,N_23458,N_24704);
xnor UO_2324 (O_2324,N_24220,N_23044);
or UO_2325 (O_2325,N_23036,N_22948);
and UO_2326 (O_2326,N_23491,N_23505);
xnor UO_2327 (O_2327,N_23229,N_22969);
or UO_2328 (O_2328,N_23082,N_24611);
nor UO_2329 (O_2329,N_24553,N_24497);
and UO_2330 (O_2330,N_24840,N_24130);
or UO_2331 (O_2331,N_24847,N_23827);
nand UO_2332 (O_2332,N_22621,N_23122);
nor UO_2333 (O_2333,N_22821,N_23813);
xnor UO_2334 (O_2334,N_23453,N_22607);
nor UO_2335 (O_2335,N_22627,N_22733);
nand UO_2336 (O_2336,N_24299,N_22976);
or UO_2337 (O_2337,N_24439,N_22875);
and UO_2338 (O_2338,N_24066,N_22900);
nand UO_2339 (O_2339,N_23192,N_23824);
nor UO_2340 (O_2340,N_24651,N_24746);
nor UO_2341 (O_2341,N_24026,N_24773);
or UO_2342 (O_2342,N_24814,N_23895);
xnor UO_2343 (O_2343,N_24507,N_24843);
or UO_2344 (O_2344,N_24044,N_23131);
xnor UO_2345 (O_2345,N_23467,N_24882);
nor UO_2346 (O_2346,N_24052,N_24748);
or UO_2347 (O_2347,N_24848,N_23702);
and UO_2348 (O_2348,N_23740,N_22893);
xor UO_2349 (O_2349,N_24422,N_23224);
nor UO_2350 (O_2350,N_24312,N_23797);
nor UO_2351 (O_2351,N_24129,N_23694);
xor UO_2352 (O_2352,N_23651,N_23905);
and UO_2353 (O_2353,N_23303,N_23739);
nand UO_2354 (O_2354,N_24509,N_23112);
nor UO_2355 (O_2355,N_23447,N_22896);
nand UO_2356 (O_2356,N_23544,N_23299);
or UO_2357 (O_2357,N_22673,N_24108);
and UO_2358 (O_2358,N_24951,N_23747);
and UO_2359 (O_2359,N_23125,N_22886);
xor UO_2360 (O_2360,N_23223,N_23751);
nand UO_2361 (O_2361,N_23047,N_24639);
nor UO_2362 (O_2362,N_23101,N_23645);
and UO_2363 (O_2363,N_22696,N_23331);
or UO_2364 (O_2364,N_24683,N_23324);
or UO_2365 (O_2365,N_23869,N_24579);
nand UO_2366 (O_2366,N_23351,N_24890);
or UO_2367 (O_2367,N_24866,N_22622);
nor UO_2368 (O_2368,N_24806,N_22603);
xor UO_2369 (O_2369,N_23566,N_24976);
nor UO_2370 (O_2370,N_24509,N_22576);
and UO_2371 (O_2371,N_24567,N_24659);
or UO_2372 (O_2372,N_24120,N_23516);
nor UO_2373 (O_2373,N_22507,N_23193);
xnor UO_2374 (O_2374,N_24360,N_24238);
and UO_2375 (O_2375,N_23609,N_24116);
nor UO_2376 (O_2376,N_23545,N_22990);
nand UO_2377 (O_2377,N_23232,N_22951);
xor UO_2378 (O_2378,N_23045,N_24097);
and UO_2379 (O_2379,N_23641,N_22810);
nand UO_2380 (O_2380,N_24138,N_24316);
or UO_2381 (O_2381,N_24929,N_23327);
nor UO_2382 (O_2382,N_22564,N_23058);
and UO_2383 (O_2383,N_24543,N_24789);
or UO_2384 (O_2384,N_24041,N_24443);
xnor UO_2385 (O_2385,N_22874,N_23685);
and UO_2386 (O_2386,N_23679,N_24919);
xnor UO_2387 (O_2387,N_24408,N_23805);
nor UO_2388 (O_2388,N_24558,N_23955);
nand UO_2389 (O_2389,N_24513,N_23070);
nor UO_2390 (O_2390,N_22877,N_23917);
nor UO_2391 (O_2391,N_23299,N_23103);
xnor UO_2392 (O_2392,N_22934,N_24695);
nor UO_2393 (O_2393,N_23520,N_24716);
nor UO_2394 (O_2394,N_24375,N_23912);
and UO_2395 (O_2395,N_22687,N_24014);
xor UO_2396 (O_2396,N_23813,N_24065);
and UO_2397 (O_2397,N_23127,N_23936);
nand UO_2398 (O_2398,N_24592,N_22515);
nor UO_2399 (O_2399,N_23319,N_22550);
and UO_2400 (O_2400,N_23587,N_23105);
nor UO_2401 (O_2401,N_23641,N_24689);
xnor UO_2402 (O_2402,N_23632,N_22772);
or UO_2403 (O_2403,N_24232,N_22863);
nand UO_2404 (O_2404,N_22639,N_23481);
and UO_2405 (O_2405,N_23545,N_22672);
or UO_2406 (O_2406,N_23160,N_24620);
xnor UO_2407 (O_2407,N_23547,N_23576);
xor UO_2408 (O_2408,N_24268,N_22949);
xor UO_2409 (O_2409,N_24519,N_24847);
or UO_2410 (O_2410,N_22836,N_23267);
nand UO_2411 (O_2411,N_23103,N_24786);
xor UO_2412 (O_2412,N_22538,N_24140);
nand UO_2413 (O_2413,N_22787,N_22829);
or UO_2414 (O_2414,N_24569,N_22924);
or UO_2415 (O_2415,N_24675,N_22573);
nor UO_2416 (O_2416,N_24481,N_23317);
and UO_2417 (O_2417,N_23544,N_24485);
nor UO_2418 (O_2418,N_23451,N_23753);
xor UO_2419 (O_2419,N_24220,N_23173);
nor UO_2420 (O_2420,N_23689,N_24531);
nand UO_2421 (O_2421,N_23185,N_23880);
nand UO_2422 (O_2422,N_24627,N_23575);
or UO_2423 (O_2423,N_23830,N_23138);
nor UO_2424 (O_2424,N_24529,N_22684);
and UO_2425 (O_2425,N_24718,N_23723);
nand UO_2426 (O_2426,N_24769,N_22507);
or UO_2427 (O_2427,N_23049,N_24719);
and UO_2428 (O_2428,N_24718,N_22676);
and UO_2429 (O_2429,N_22776,N_22658);
and UO_2430 (O_2430,N_24516,N_24133);
or UO_2431 (O_2431,N_24164,N_23980);
and UO_2432 (O_2432,N_24880,N_24623);
nor UO_2433 (O_2433,N_24783,N_24243);
and UO_2434 (O_2434,N_22523,N_23132);
and UO_2435 (O_2435,N_22527,N_24731);
and UO_2436 (O_2436,N_22842,N_24936);
or UO_2437 (O_2437,N_22901,N_23939);
nor UO_2438 (O_2438,N_22752,N_22760);
xor UO_2439 (O_2439,N_23547,N_23832);
or UO_2440 (O_2440,N_24235,N_24668);
nor UO_2441 (O_2441,N_22788,N_22925);
or UO_2442 (O_2442,N_24034,N_24620);
nand UO_2443 (O_2443,N_23928,N_23840);
or UO_2444 (O_2444,N_22885,N_23079);
and UO_2445 (O_2445,N_24260,N_24599);
and UO_2446 (O_2446,N_23875,N_23652);
nand UO_2447 (O_2447,N_22520,N_22990);
nor UO_2448 (O_2448,N_23492,N_24865);
and UO_2449 (O_2449,N_24416,N_24789);
nor UO_2450 (O_2450,N_22909,N_23033);
xor UO_2451 (O_2451,N_24344,N_24430);
and UO_2452 (O_2452,N_22533,N_22907);
or UO_2453 (O_2453,N_24270,N_24931);
or UO_2454 (O_2454,N_22827,N_24462);
nor UO_2455 (O_2455,N_24280,N_22787);
or UO_2456 (O_2456,N_22669,N_23287);
xor UO_2457 (O_2457,N_22899,N_24399);
or UO_2458 (O_2458,N_24933,N_24125);
nand UO_2459 (O_2459,N_24839,N_22917);
nand UO_2460 (O_2460,N_24631,N_23389);
and UO_2461 (O_2461,N_22800,N_23550);
xor UO_2462 (O_2462,N_24132,N_23676);
nor UO_2463 (O_2463,N_24196,N_24265);
xor UO_2464 (O_2464,N_24923,N_23175);
xnor UO_2465 (O_2465,N_23557,N_22712);
nand UO_2466 (O_2466,N_22970,N_23780);
nor UO_2467 (O_2467,N_24277,N_23942);
or UO_2468 (O_2468,N_22502,N_24658);
nand UO_2469 (O_2469,N_23185,N_23178);
xnor UO_2470 (O_2470,N_22811,N_23551);
or UO_2471 (O_2471,N_24452,N_23554);
or UO_2472 (O_2472,N_23562,N_23056);
and UO_2473 (O_2473,N_24660,N_24124);
nor UO_2474 (O_2474,N_24420,N_23405);
nand UO_2475 (O_2475,N_23295,N_23543);
nand UO_2476 (O_2476,N_24356,N_22715);
and UO_2477 (O_2477,N_23304,N_22716);
nor UO_2478 (O_2478,N_23713,N_23849);
xnor UO_2479 (O_2479,N_24891,N_23056);
and UO_2480 (O_2480,N_23477,N_22939);
xor UO_2481 (O_2481,N_24463,N_23754);
xor UO_2482 (O_2482,N_23050,N_24900);
nor UO_2483 (O_2483,N_23073,N_24093);
or UO_2484 (O_2484,N_22962,N_23625);
nor UO_2485 (O_2485,N_22733,N_23590);
xnor UO_2486 (O_2486,N_24133,N_23838);
nor UO_2487 (O_2487,N_24937,N_22531);
and UO_2488 (O_2488,N_24155,N_23637);
nand UO_2489 (O_2489,N_24738,N_22945);
and UO_2490 (O_2490,N_23093,N_24534);
and UO_2491 (O_2491,N_24773,N_24465);
and UO_2492 (O_2492,N_22501,N_23841);
xnor UO_2493 (O_2493,N_24905,N_23129);
nand UO_2494 (O_2494,N_22718,N_23292);
and UO_2495 (O_2495,N_22887,N_23720);
xor UO_2496 (O_2496,N_24241,N_23071);
nand UO_2497 (O_2497,N_22976,N_22740);
and UO_2498 (O_2498,N_22582,N_23863);
and UO_2499 (O_2499,N_24373,N_24638);
xor UO_2500 (O_2500,N_24261,N_22609);
or UO_2501 (O_2501,N_22691,N_22791);
xnor UO_2502 (O_2502,N_23770,N_24251);
nand UO_2503 (O_2503,N_23249,N_24559);
nand UO_2504 (O_2504,N_24241,N_24312);
and UO_2505 (O_2505,N_23685,N_23380);
nand UO_2506 (O_2506,N_24788,N_22621);
xor UO_2507 (O_2507,N_24225,N_22980);
nor UO_2508 (O_2508,N_22687,N_22931);
and UO_2509 (O_2509,N_23612,N_24278);
nand UO_2510 (O_2510,N_22741,N_23053);
and UO_2511 (O_2511,N_23828,N_24609);
nor UO_2512 (O_2512,N_24180,N_24981);
or UO_2513 (O_2513,N_23750,N_23720);
xor UO_2514 (O_2514,N_23106,N_23835);
or UO_2515 (O_2515,N_23927,N_24539);
nand UO_2516 (O_2516,N_22779,N_23887);
nor UO_2517 (O_2517,N_24745,N_23309);
nand UO_2518 (O_2518,N_23273,N_24849);
or UO_2519 (O_2519,N_23371,N_22608);
xnor UO_2520 (O_2520,N_22977,N_22502);
nand UO_2521 (O_2521,N_23876,N_24149);
xnor UO_2522 (O_2522,N_24053,N_24114);
and UO_2523 (O_2523,N_24162,N_24467);
nor UO_2524 (O_2524,N_24263,N_24415);
nor UO_2525 (O_2525,N_24351,N_24163);
nor UO_2526 (O_2526,N_23757,N_22735);
nand UO_2527 (O_2527,N_23986,N_23663);
or UO_2528 (O_2528,N_24345,N_23646);
and UO_2529 (O_2529,N_24144,N_23268);
nand UO_2530 (O_2530,N_24818,N_23214);
or UO_2531 (O_2531,N_22908,N_24219);
or UO_2532 (O_2532,N_22538,N_23218);
nand UO_2533 (O_2533,N_23114,N_23229);
and UO_2534 (O_2534,N_22560,N_22537);
or UO_2535 (O_2535,N_23677,N_23001);
and UO_2536 (O_2536,N_24541,N_22732);
nor UO_2537 (O_2537,N_22774,N_23417);
xnor UO_2538 (O_2538,N_24233,N_22646);
xnor UO_2539 (O_2539,N_24861,N_24978);
nand UO_2540 (O_2540,N_23667,N_22560);
xnor UO_2541 (O_2541,N_24794,N_22728);
and UO_2542 (O_2542,N_24716,N_24269);
nor UO_2543 (O_2543,N_22956,N_24551);
or UO_2544 (O_2544,N_23940,N_22699);
or UO_2545 (O_2545,N_24432,N_23441);
or UO_2546 (O_2546,N_23794,N_22842);
and UO_2547 (O_2547,N_24735,N_24629);
nand UO_2548 (O_2548,N_24794,N_24324);
or UO_2549 (O_2549,N_23975,N_24528);
and UO_2550 (O_2550,N_23745,N_24293);
and UO_2551 (O_2551,N_23798,N_24293);
nor UO_2552 (O_2552,N_23189,N_22901);
or UO_2553 (O_2553,N_23865,N_24258);
nor UO_2554 (O_2554,N_23833,N_23567);
or UO_2555 (O_2555,N_23021,N_24017);
nor UO_2556 (O_2556,N_23153,N_24782);
xor UO_2557 (O_2557,N_24874,N_24092);
or UO_2558 (O_2558,N_24474,N_23065);
and UO_2559 (O_2559,N_23101,N_22896);
nor UO_2560 (O_2560,N_23877,N_22697);
or UO_2561 (O_2561,N_23511,N_22800);
nor UO_2562 (O_2562,N_23287,N_23222);
nand UO_2563 (O_2563,N_23250,N_23491);
nor UO_2564 (O_2564,N_24505,N_23061);
and UO_2565 (O_2565,N_23741,N_24284);
nor UO_2566 (O_2566,N_24622,N_24401);
or UO_2567 (O_2567,N_23496,N_24276);
nor UO_2568 (O_2568,N_23470,N_23656);
nor UO_2569 (O_2569,N_24080,N_22559);
nor UO_2570 (O_2570,N_22882,N_24766);
or UO_2571 (O_2571,N_23463,N_24308);
and UO_2572 (O_2572,N_22948,N_23869);
nand UO_2573 (O_2573,N_23899,N_24557);
nor UO_2574 (O_2574,N_23260,N_23309);
nor UO_2575 (O_2575,N_23766,N_23020);
and UO_2576 (O_2576,N_24515,N_24639);
nand UO_2577 (O_2577,N_22727,N_22708);
nor UO_2578 (O_2578,N_23002,N_23283);
nor UO_2579 (O_2579,N_23553,N_22692);
and UO_2580 (O_2580,N_23268,N_23458);
or UO_2581 (O_2581,N_24583,N_24488);
nor UO_2582 (O_2582,N_23394,N_23560);
and UO_2583 (O_2583,N_24189,N_23453);
or UO_2584 (O_2584,N_24876,N_22628);
and UO_2585 (O_2585,N_23575,N_22644);
xnor UO_2586 (O_2586,N_24565,N_24402);
nor UO_2587 (O_2587,N_24164,N_22867);
and UO_2588 (O_2588,N_22691,N_24450);
or UO_2589 (O_2589,N_23363,N_23407);
and UO_2590 (O_2590,N_23656,N_24935);
nor UO_2591 (O_2591,N_23176,N_23499);
and UO_2592 (O_2592,N_22528,N_23175);
and UO_2593 (O_2593,N_24422,N_22716);
nand UO_2594 (O_2594,N_24739,N_24310);
nand UO_2595 (O_2595,N_24680,N_24034);
xor UO_2596 (O_2596,N_22865,N_24566);
nand UO_2597 (O_2597,N_23010,N_24091);
nor UO_2598 (O_2598,N_24123,N_22575);
and UO_2599 (O_2599,N_24619,N_22946);
nor UO_2600 (O_2600,N_23519,N_24522);
or UO_2601 (O_2601,N_23831,N_22847);
nor UO_2602 (O_2602,N_22624,N_24375);
nor UO_2603 (O_2603,N_23998,N_23269);
nor UO_2604 (O_2604,N_23380,N_24615);
or UO_2605 (O_2605,N_22855,N_22681);
nand UO_2606 (O_2606,N_23608,N_23153);
or UO_2607 (O_2607,N_24144,N_23359);
xor UO_2608 (O_2608,N_24806,N_23474);
or UO_2609 (O_2609,N_24456,N_22614);
and UO_2610 (O_2610,N_22756,N_24677);
and UO_2611 (O_2611,N_23909,N_24392);
nor UO_2612 (O_2612,N_23323,N_24354);
or UO_2613 (O_2613,N_24996,N_23468);
or UO_2614 (O_2614,N_22862,N_22872);
nand UO_2615 (O_2615,N_22658,N_22727);
nor UO_2616 (O_2616,N_22548,N_22927);
xnor UO_2617 (O_2617,N_22578,N_22609);
or UO_2618 (O_2618,N_23968,N_23079);
nand UO_2619 (O_2619,N_24464,N_23714);
and UO_2620 (O_2620,N_23939,N_23198);
and UO_2621 (O_2621,N_24503,N_24808);
xor UO_2622 (O_2622,N_24283,N_23411);
nor UO_2623 (O_2623,N_24341,N_24537);
nor UO_2624 (O_2624,N_24393,N_22814);
xnor UO_2625 (O_2625,N_23482,N_23517);
nor UO_2626 (O_2626,N_23385,N_23983);
nand UO_2627 (O_2627,N_23773,N_23875);
xor UO_2628 (O_2628,N_23753,N_24727);
xnor UO_2629 (O_2629,N_23097,N_24258);
xnor UO_2630 (O_2630,N_24389,N_24403);
nand UO_2631 (O_2631,N_23896,N_23369);
and UO_2632 (O_2632,N_22682,N_23307);
xor UO_2633 (O_2633,N_24794,N_24887);
or UO_2634 (O_2634,N_24306,N_22709);
nand UO_2635 (O_2635,N_23853,N_23172);
nor UO_2636 (O_2636,N_23847,N_24769);
xor UO_2637 (O_2637,N_24717,N_24313);
and UO_2638 (O_2638,N_23376,N_24568);
nand UO_2639 (O_2639,N_23608,N_22965);
and UO_2640 (O_2640,N_24540,N_23898);
xor UO_2641 (O_2641,N_24116,N_23195);
nand UO_2642 (O_2642,N_23934,N_22761);
xor UO_2643 (O_2643,N_23617,N_24900);
xor UO_2644 (O_2644,N_23128,N_24941);
xnor UO_2645 (O_2645,N_23155,N_22972);
or UO_2646 (O_2646,N_23720,N_24333);
xor UO_2647 (O_2647,N_23634,N_23881);
or UO_2648 (O_2648,N_23392,N_22543);
xnor UO_2649 (O_2649,N_24994,N_24423);
or UO_2650 (O_2650,N_23787,N_23318);
or UO_2651 (O_2651,N_24693,N_22847);
nor UO_2652 (O_2652,N_22706,N_24731);
nand UO_2653 (O_2653,N_22515,N_24744);
and UO_2654 (O_2654,N_24642,N_22584);
and UO_2655 (O_2655,N_24696,N_23805);
xor UO_2656 (O_2656,N_22512,N_24676);
or UO_2657 (O_2657,N_24885,N_24715);
nor UO_2658 (O_2658,N_22597,N_24202);
nand UO_2659 (O_2659,N_23056,N_23319);
xnor UO_2660 (O_2660,N_23533,N_22511);
nand UO_2661 (O_2661,N_24544,N_24222);
xor UO_2662 (O_2662,N_23966,N_23683);
xor UO_2663 (O_2663,N_23789,N_22828);
nand UO_2664 (O_2664,N_23042,N_23082);
nor UO_2665 (O_2665,N_22942,N_22921);
xnor UO_2666 (O_2666,N_24481,N_24169);
and UO_2667 (O_2667,N_23625,N_23806);
or UO_2668 (O_2668,N_22529,N_24577);
and UO_2669 (O_2669,N_23524,N_23988);
xnor UO_2670 (O_2670,N_24638,N_23582);
xnor UO_2671 (O_2671,N_23166,N_24710);
xnor UO_2672 (O_2672,N_24568,N_23674);
or UO_2673 (O_2673,N_24320,N_23294);
or UO_2674 (O_2674,N_22828,N_23967);
xnor UO_2675 (O_2675,N_22830,N_24438);
and UO_2676 (O_2676,N_24490,N_23665);
xor UO_2677 (O_2677,N_24949,N_24449);
nand UO_2678 (O_2678,N_22660,N_23494);
or UO_2679 (O_2679,N_24193,N_24667);
xnor UO_2680 (O_2680,N_23374,N_23608);
xnor UO_2681 (O_2681,N_24181,N_24372);
nand UO_2682 (O_2682,N_24965,N_23305);
or UO_2683 (O_2683,N_24786,N_22714);
and UO_2684 (O_2684,N_22634,N_22872);
or UO_2685 (O_2685,N_22760,N_23538);
or UO_2686 (O_2686,N_24845,N_24043);
nor UO_2687 (O_2687,N_24787,N_23214);
nand UO_2688 (O_2688,N_24595,N_23443);
nand UO_2689 (O_2689,N_23992,N_23198);
nor UO_2690 (O_2690,N_23747,N_24361);
or UO_2691 (O_2691,N_22904,N_23761);
or UO_2692 (O_2692,N_24064,N_23582);
nor UO_2693 (O_2693,N_24788,N_23939);
and UO_2694 (O_2694,N_24941,N_24836);
xnor UO_2695 (O_2695,N_22809,N_23408);
nand UO_2696 (O_2696,N_23817,N_22922);
xor UO_2697 (O_2697,N_22706,N_23679);
nand UO_2698 (O_2698,N_23482,N_23519);
nor UO_2699 (O_2699,N_24685,N_24390);
or UO_2700 (O_2700,N_23688,N_22640);
or UO_2701 (O_2701,N_24540,N_24437);
nor UO_2702 (O_2702,N_23751,N_23796);
xnor UO_2703 (O_2703,N_22704,N_22921);
nand UO_2704 (O_2704,N_23410,N_22758);
or UO_2705 (O_2705,N_22775,N_22623);
nor UO_2706 (O_2706,N_23532,N_24899);
nand UO_2707 (O_2707,N_22721,N_24989);
and UO_2708 (O_2708,N_23841,N_23809);
and UO_2709 (O_2709,N_22906,N_23286);
and UO_2710 (O_2710,N_23994,N_22557);
or UO_2711 (O_2711,N_24085,N_24950);
xnor UO_2712 (O_2712,N_22805,N_24983);
or UO_2713 (O_2713,N_23119,N_24312);
xnor UO_2714 (O_2714,N_23246,N_22580);
xnor UO_2715 (O_2715,N_22948,N_24919);
nand UO_2716 (O_2716,N_23881,N_23432);
nor UO_2717 (O_2717,N_24086,N_22663);
or UO_2718 (O_2718,N_22924,N_24120);
or UO_2719 (O_2719,N_23211,N_23142);
and UO_2720 (O_2720,N_24005,N_22868);
xnor UO_2721 (O_2721,N_24298,N_23845);
nor UO_2722 (O_2722,N_22686,N_22968);
xor UO_2723 (O_2723,N_22715,N_23392);
or UO_2724 (O_2724,N_23300,N_24484);
and UO_2725 (O_2725,N_24719,N_22967);
xor UO_2726 (O_2726,N_24238,N_23094);
xnor UO_2727 (O_2727,N_23098,N_23299);
or UO_2728 (O_2728,N_23532,N_24593);
or UO_2729 (O_2729,N_24432,N_24189);
nor UO_2730 (O_2730,N_23355,N_23170);
nor UO_2731 (O_2731,N_22742,N_24304);
and UO_2732 (O_2732,N_24592,N_23066);
and UO_2733 (O_2733,N_23292,N_23870);
nor UO_2734 (O_2734,N_24968,N_24687);
nand UO_2735 (O_2735,N_24185,N_24147);
nand UO_2736 (O_2736,N_23874,N_24398);
or UO_2737 (O_2737,N_22958,N_22670);
nor UO_2738 (O_2738,N_23675,N_24881);
nand UO_2739 (O_2739,N_22848,N_24881);
or UO_2740 (O_2740,N_24330,N_24042);
or UO_2741 (O_2741,N_22557,N_23183);
nor UO_2742 (O_2742,N_23522,N_23041);
or UO_2743 (O_2743,N_24064,N_23977);
xnor UO_2744 (O_2744,N_24870,N_24442);
or UO_2745 (O_2745,N_22734,N_23455);
nor UO_2746 (O_2746,N_23628,N_24573);
nand UO_2747 (O_2747,N_24543,N_23361);
nor UO_2748 (O_2748,N_23162,N_23896);
nand UO_2749 (O_2749,N_22956,N_23770);
nor UO_2750 (O_2750,N_22870,N_22659);
or UO_2751 (O_2751,N_24193,N_23641);
xnor UO_2752 (O_2752,N_23967,N_23423);
nand UO_2753 (O_2753,N_23285,N_23346);
xor UO_2754 (O_2754,N_24497,N_22708);
xor UO_2755 (O_2755,N_23615,N_23051);
or UO_2756 (O_2756,N_24928,N_24364);
and UO_2757 (O_2757,N_24325,N_23338);
and UO_2758 (O_2758,N_24250,N_23997);
or UO_2759 (O_2759,N_24700,N_24329);
nand UO_2760 (O_2760,N_24617,N_23221);
and UO_2761 (O_2761,N_23517,N_22500);
nor UO_2762 (O_2762,N_22819,N_23965);
or UO_2763 (O_2763,N_23509,N_24604);
nand UO_2764 (O_2764,N_24113,N_22764);
and UO_2765 (O_2765,N_22974,N_24239);
xnor UO_2766 (O_2766,N_23506,N_24296);
or UO_2767 (O_2767,N_24134,N_23519);
nand UO_2768 (O_2768,N_24711,N_24693);
and UO_2769 (O_2769,N_22839,N_24916);
xnor UO_2770 (O_2770,N_23858,N_24335);
nor UO_2771 (O_2771,N_23041,N_23665);
and UO_2772 (O_2772,N_23255,N_23378);
xnor UO_2773 (O_2773,N_23978,N_24673);
or UO_2774 (O_2774,N_23926,N_23703);
nand UO_2775 (O_2775,N_23590,N_24539);
xnor UO_2776 (O_2776,N_24535,N_23823);
or UO_2777 (O_2777,N_23644,N_24679);
or UO_2778 (O_2778,N_23345,N_24070);
xnor UO_2779 (O_2779,N_24876,N_24553);
or UO_2780 (O_2780,N_24827,N_24573);
or UO_2781 (O_2781,N_24364,N_23296);
nand UO_2782 (O_2782,N_23982,N_24066);
and UO_2783 (O_2783,N_24661,N_24507);
or UO_2784 (O_2784,N_22911,N_22958);
nor UO_2785 (O_2785,N_23278,N_23637);
xnor UO_2786 (O_2786,N_24736,N_24584);
and UO_2787 (O_2787,N_24748,N_23871);
xnor UO_2788 (O_2788,N_22555,N_23606);
or UO_2789 (O_2789,N_22800,N_24963);
or UO_2790 (O_2790,N_23982,N_24230);
xnor UO_2791 (O_2791,N_22763,N_23965);
nor UO_2792 (O_2792,N_22815,N_24075);
nor UO_2793 (O_2793,N_23080,N_24642);
or UO_2794 (O_2794,N_24176,N_24815);
and UO_2795 (O_2795,N_23649,N_23892);
or UO_2796 (O_2796,N_22967,N_24328);
or UO_2797 (O_2797,N_23035,N_24828);
and UO_2798 (O_2798,N_24589,N_24573);
nand UO_2799 (O_2799,N_24266,N_24529);
or UO_2800 (O_2800,N_22671,N_23310);
nor UO_2801 (O_2801,N_24641,N_23808);
xor UO_2802 (O_2802,N_24716,N_23753);
nor UO_2803 (O_2803,N_23751,N_23541);
xor UO_2804 (O_2804,N_23645,N_23591);
or UO_2805 (O_2805,N_24746,N_24726);
or UO_2806 (O_2806,N_23284,N_23481);
nor UO_2807 (O_2807,N_23098,N_22975);
or UO_2808 (O_2808,N_24101,N_24501);
or UO_2809 (O_2809,N_23390,N_24761);
and UO_2810 (O_2810,N_24944,N_23438);
or UO_2811 (O_2811,N_23358,N_23389);
nand UO_2812 (O_2812,N_22853,N_23888);
xor UO_2813 (O_2813,N_24160,N_24124);
xor UO_2814 (O_2814,N_24699,N_23730);
xor UO_2815 (O_2815,N_22830,N_23410);
and UO_2816 (O_2816,N_22777,N_22938);
nand UO_2817 (O_2817,N_24216,N_24789);
xnor UO_2818 (O_2818,N_23783,N_23606);
or UO_2819 (O_2819,N_22796,N_24778);
nand UO_2820 (O_2820,N_24819,N_24386);
nor UO_2821 (O_2821,N_24269,N_22708);
nor UO_2822 (O_2822,N_23235,N_24562);
nand UO_2823 (O_2823,N_23660,N_23530);
xor UO_2824 (O_2824,N_23529,N_23025);
nand UO_2825 (O_2825,N_24712,N_24162);
or UO_2826 (O_2826,N_23918,N_24560);
nand UO_2827 (O_2827,N_24966,N_23562);
and UO_2828 (O_2828,N_22553,N_22562);
xnor UO_2829 (O_2829,N_23706,N_23844);
or UO_2830 (O_2830,N_23374,N_23682);
nand UO_2831 (O_2831,N_23557,N_24114);
nand UO_2832 (O_2832,N_23528,N_24117);
or UO_2833 (O_2833,N_22554,N_24150);
and UO_2834 (O_2834,N_24958,N_24270);
xnor UO_2835 (O_2835,N_24532,N_24912);
nor UO_2836 (O_2836,N_23560,N_22913);
or UO_2837 (O_2837,N_22714,N_22565);
nand UO_2838 (O_2838,N_23463,N_24819);
nand UO_2839 (O_2839,N_23705,N_24777);
or UO_2840 (O_2840,N_23240,N_23050);
and UO_2841 (O_2841,N_22701,N_24404);
nand UO_2842 (O_2842,N_22812,N_24427);
and UO_2843 (O_2843,N_24186,N_24785);
xnor UO_2844 (O_2844,N_23411,N_23129);
xor UO_2845 (O_2845,N_23593,N_23257);
or UO_2846 (O_2846,N_24549,N_23196);
or UO_2847 (O_2847,N_23271,N_24527);
nor UO_2848 (O_2848,N_24663,N_24181);
nor UO_2849 (O_2849,N_23290,N_22951);
nor UO_2850 (O_2850,N_23407,N_22559);
and UO_2851 (O_2851,N_23476,N_23134);
xnor UO_2852 (O_2852,N_22973,N_23165);
nand UO_2853 (O_2853,N_22782,N_24034);
xnor UO_2854 (O_2854,N_23255,N_23423);
and UO_2855 (O_2855,N_24785,N_24758);
nor UO_2856 (O_2856,N_23150,N_23108);
and UO_2857 (O_2857,N_24942,N_24914);
and UO_2858 (O_2858,N_24110,N_24641);
nor UO_2859 (O_2859,N_23989,N_23451);
xnor UO_2860 (O_2860,N_24236,N_22601);
and UO_2861 (O_2861,N_23662,N_22876);
nand UO_2862 (O_2862,N_23983,N_24410);
and UO_2863 (O_2863,N_24105,N_22848);
and UO_2864 (O_2864,N_22993,N_24098);
nor UO_2865 (O_2865,N_24127,N_23371);
nand UO_2866 (O_2866,N_22615,N_23217);
nor UO_2867 (O_2867,N_24347,N_24118);
nor UO_2868 (O_2868,N_24048,N_24413);
and UO_2869 (O_2869,N_24074,N_23327);
xnor UO_2870 (O_2870,N_24526,N_22714);
and UO_2871 (O_2871,N_23001,N_24563);
nor UO_2872 (O_2872,N_24989,N_22895);
nand UO_2873 (O_2873,N_24975,N_22508);
and UO_2874 (O_2874,N_23506,N_23156);
or UO_2875 (O_2875,N_24636,N_24619);
nand UO_2876 (O_2876,N_24366,N_23220);
nand UO_2877 (O_2877,N_24372,N_24061);
and UO_2878 (O_2878,N_23470,N_24974);
or UO_2879 (O_2879,N_23420,N_24346);
and UO_2880 (O_2880,N_22912,N_24454);
and UO_2881 (O_2881,N_23014,N_23215);
or UO_2882 (O_2882,N_24852,N_22587);
nand UO_2883 (O_2883,N_24215,N_24024);
nor UO_2884 (O_2884,N_22753,N_23729);
nand UO_2885 (O_2885,N_24777,N_24458);
or UO_2886 (O_2886,N_24499,N_24871);
nand UO_2887 (O_2887,N_23234,N_24599);
nor UO_2888 (O_2888,N_23022,N_23612);
nand UO_2889 (O_2889,N_24949,N_22513);
or UO_2890 (O_2890,N_23265,N_23429);
or UO_2891 (O_2891,N_24609,N_24583);
xor UO_2892 (O_2892,N_24294,N_24888);
and UO_2893 (O_2893,N_23817,N_23880);
nor UO_2894 (O_2894,N_22613,N_23738);
xnor UO_2895 (O_2895,N_23445,N_22999);
nand UO_2896 (O_2896,N_24551,N_24533);
and UO_2897 (O_2897,N_24734,N_23189);
nor UO_2898 (O_2898,N_24176,N_23865);
nand UO_2899 (O_2899,N_23394,N_23557);
nor UO_2900 (O_2900,N_22716,N_24348);
xor UO_2901 (O_2901,N_24558,N_23635);
nand UO_2902 (O_2902,N_23282,N_24051);
nor UO_2903 (O_2903,N_24594,N_22944);
nand UO_2904 (O_2904,N_24810,N_23051);
nor UO_2905 (O_2905,N_22730,N_22952);
and UO_2906 (O_2906,N_22793,N_24963);
xnor UO_2907 (O_2907,N_22668,N_24960);
or UO_2908 (O_2908,N_22509,N_24312);
nor UO_2909 (O_2909,N_23881,N_24442);
or UO_2910 (O_2910,N_24163,N_24562);
nand UO_2911 (O_2911,N_23492,N_23421);
and UO_2912 (O_2912,N_23999,N_22695);
xnor UO_2913 (O_2913,N_23126,N_24006);
xor UO_2914 (O_2914,N_23271,N_24455);
and UO_2915 (O_2915,N_24892,N_23798);
or UO_2916 (O_2916,N_23519,N_24734);
and UO_2917 (O_2917,N_22688,N_22786);
nor UO_2918 (O_2918,N_24115,N_23150);
nand UO_2919 (O_2919,N_23595,N_24336);
xor UO_2920 (O_2920,N_22637,N_23729);
nand UO_2921 (O_2921,N_24374,N_22985);
or UO_2922 (O_2922,N_22530,N_22543);
nor UO_2923 (O_2923,N_22693,N_23392);
nor UO_2924 (O_2924,N_24226,N_23211);
and UO_2925 (O_2925,N_23879,N_24635);
xnor UO_2926 (O_2926,N_24738,N_24113);
nor UO_2927 (O_2927,N_24125,N_24181);
or UO_2928 (O_2928,N_23365,N_23039);
xnor UO_2929 (O_2929,N_23794,N_23270);
xnor UO_2930 (O_2930,N_24510,N_23477);
xor UO_2931 (O_2931,N_23342,N_23976);
and UO_2932 (O_2932,N_24729,N_24180);
xnor UO_2933 (O_2933,N_24636,N_24361);
or UO_2934 (O_2934,N_22634,N_23645);
xnor UO_2935 (O_2935,N_24024,N_24266);
nor UO_2936 (O_2936,N_23205,N_23156);
xnor UO_2937 (O_2937,N_23409,N_23362);
xnor UO_2938 (O_2938,N_22537,N_24001);
and UO_2939 (O_2939,N_23731,N_23325);
or UO_2940 (O_2940,N_23161,N_23357);
nor UO_2941 (O_2941,N_22610,N_23655);
nand UO_2942 (O_2942,N_22613,N_22769);
nand UO_2943 (O_2943,N_23026,N_24080);
nand UO_2944 (O_2944,N_24326,N_24381);
and UO_2945 (O_2945,N_24447,N_23224);
or UO_2946 (O_2946,N_23591,N_24651);
nor UO_2947 (O_2947,N_23450,N_23688);
nand UO_2948 (O_2948,N_23257,N_24731);
xnor UO_2949 (O_2949,N_23076,N_23026);
nand UO_2950 (O_2950,N_23670,N_22756);
nand UO_2951 (O_2951,N_23613,N_23492);
nor UO_2952 (O_2952,N_24554,N_23500);
nand UO_2953 (O_2953,N_22997,N_22891);
or UO_2954 (O_2954,N_23676,N_23895);
xnor UO_2955 (O_2955,N_23400,N_24648);
and UO_2956 (O_2956,N_24377,N_24903);
nor UO_2957 (O_2957,N_24319,N_24108);
and UO_2958 (O_2958,N_24196,N_22709);
nand UO_2959 (O_2959,N_24286,N_24235);
and UO_2960 (O_2960,N_23983,N_24591);
xor UO_2961 (O_2961,N_22853,N_22558);
and UO_2962 (O_2962,N_24225,N_23550);
and UO_2963 (O_2963,N_22822,N_24030);
and UO_2964 (O_2964,N_23098,N_24773);
nand UO_2965 (O_2965,N_24688,N_24222);
nand UO_2966 (O_2966,N_23560,N_23826);
nand UO_2967 (O_2967,N_22709,N_24230);
or UO_2968 (O_2968,N_23675,N_23838);
and UO_2969 (O_2969,N_23667,N_24812);
xnor UO_2970 (O_2970,N_24936,N_24793);
xor UO_2971 (O_2971,N_24520,N_24982);
and UO_2972 (O_2972,N_23969,N_23478);
nand UO_2973 (O_2973,N_22614,N_24497);
nand UO_2974 (O_2974,N_22561,N_23672);
xnor UO_2975 (O_2975,N_24878,N_23671);
xnor UO_2976 (O_2976,N_22951,N_23033);
and UO_2977 (O_2977,N_24715,N_24724);
or UO_2978 (O_2978,N_23903,N_23367);
nand UO_2979 (O_2979,N_23953,N_23786);
xnor UO_2980 (O_2980,N_23411,N_24755);
xor UO_2981 (O_2981,N_24397,N_24627);
or UO_2982 (O_2982,N_22710,N_24125);
or UO_2983 (O_2983,N_24077,N_24263);
or UO_2984 (O_2984,N_23355,N_23536);
nor UO_2985 (O_2985,N_22660,N_23974);
nor UO_2986 (O_2986,N_22879,N_23484);
nand UO_2987 (O_2987,N_23541,N_23226);
nand UO_2988 (O_2988,N_23657,N_22788);
nand UO_2989 (O_2989,N_24232,N_23909);
nand UO_2990 (O_2990,N_22926,N_23273);
xnor UO_2991 (O_2991,N_24824,N_23094);
or UO_2992 (O_2992,N_23925,N_23493);
nor UO_2993 (O_2993,N_23758,N_23453);
and UO_2994 (O_2994,N_23911,N_23692);
and UO_2995 (O_2995,N_22845,N_22989);
nor UO_2996 (O_2996,N_23802,N_23648);
xnor UO_2997 (O_2997,N_24171,N_23935);
nand UO_2998 (O_2998,N_22535,N_24056);
or UO_2999 (O_2999,N_24310,N_24406);
endmodule