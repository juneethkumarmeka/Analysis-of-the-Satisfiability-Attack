module basic_500_3000_500_15_levels_2xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_493,In_363);
or U1 (N_1,In_467,In_77);
nand U2 (N_2,In_419,In_41);
nor U3 (N_3,In_9,In_123);
nor U4 (N_4,In_390,In_12);
xnor U5 (N_5,In_164,In_298);
or U6 (N_6,In_206,In_483);
nand U7 (N_7,In_362,In_299);
and U8 (N_8,In_212,In_340);
and U9 (N_9,In_310,In_496);
nand U10 (N_10,In_51,In_480);
nor U11 (N_11,In_109,In_413);
and U12 (N_12,In_21,In_414);
or U13 (N_13,In_293,In_424);
nand U14 (N_14,In_331,In_246);
nor U15 (N_15,In_470,In_17);
and U16 (N_16,In_469,In_321);
or U17 (N_17,In_175,In_198);
nor U18 (N_18,In_440,In_396);
and U19 (N_19,In_292,In_410);
or U20 (N_20,In_497,In_124);
and U21 (N_21,In_63,In_380);
nand U22 (N_22,In_209,In_107);
nor U23 (N_23,In_393,In_316);
nand U24 (N_24,In_400,In_32);
and U25 (N_25,In_157,In_121);
nor U26 (N_26,In_456,In_317);
nand U27 (N_27,In_241,In_301);
nand U28 (N_28,In_348,In_314);
nand U29 (N_29,In_471,In_457);
nor U30 (N_30,In_454,In_217);
nor U31 (N_31,In_382,In_499);
or U32 (N_32,In_487,In_196);
or U33 (N_33,In_200,In_481);
or U34 (N_34,In_59,In_190);
and U35 (N_35,In_171,In_14);
nand U36 (N_36,In_168,In_227);
nand U37 (N_37,In_489,In_139);
nor U38 (N_38,In_287,In_34);
nand U39 (N_39,In_412,In_486);
nor U40 (N_40,In_237,In_182);
or U41 (N_41,In_229,In_436);
nand U42 (N_42,In_374,In_27);
nand U43 (N_43,In_401,In_408);
and U44 (N_44,In_52,In_16);
xnor U45 (N_45,In_148,In_88);
or U46 (N_46,In_322,In_304);
and U47 (N_47,In_71,In_265);
or U48 (N_48,In_22,In_389);
and U49 (N_49,In_365,In_201);
and U50 (N_50,In_294,In_67);
or U51 (N_51,In_319,In_238);
and U52 (N_52,In_330,In_267);
nand U53 (N_53,In_335,In_387);
and U54 (N_54,In_129,In_90);
xor U55 (N_55,In_285,In_482);
or U56 (N_56,In_133,In_431);
and U57 (N_57,In_465,In_233);
nor U58 (N_58,In_367,In_208);
and U59 (N_59,In_307,In_189);
or U60 (N_60,In_268,In_485);
or U61 (N_61,In_74,In_156);
and U62 (N_62,In_395,In_179);
xor U63 (N_63,In_366,In_118);
or U64 (N_64,In_49,In_38);
nand U65 (N_65,In_136,In_42);
or U66 (N_66,In_347,In_441);
or U67 (N_67,In_86,In_281);
nand U68 (N_68,In_353,In_255);
or U69 (N_69,In_50,In_327);
nor U70 (N_70,In_384,In_339);
or U71 (N_71,In_165,In_250);
nand U72 (N_72,In_418,In_388);
nand U73 (N_73,In_249,In_120);
nand U74 (N_74,In_93,In_214);
nand U75 (N_75,In_188,In_141);
nand U76 (N_76,In_448,In_111);
and U77 (N_77,In_442,In_404);
nor U78 (N_78,In_76,In_296);
xor U79 (N_79,In_272,In_96);
and U80 (N_80,In_279,In_55);
nor U81 (N_81,In_194,In_75);
and U82 (N_82,In_333,In_94);
nor U83 (N_83,In_460,In_358);
and U84 (N_84,In_213,In_427);
or U85 (N_85,In_283,In_385);
nand U86 (N_86,In_459,In_100);
and U87 (N_87,In_463,In_172);
nand U88 (N_88,In_159,In_302);
and U89 (N_89,In_167,In_24);
or U90 (N_90,In_352,In_324);
nand U91 (N_91,In_342,In_259);
or U92 (N_92,In_429,In_166);
and U93 (N_93,In_420,In_140);
and U94 (N_94,In_376,In_473);
nand U95 (N_95,In_318,In_343);
and U96 (N_96,In_33,In_476);
and U97 (N_97,In_170,In_355);
nor U98 (N_98,In_223,In_328);
or U99 (N_99,In_58,In_54);
nand U100 (N_100,In_433,In_432);
nand U101 (N_101,In_492,In_313);
and U102 (N_102,In_210,In_325);
and U103 (N_103,In_407,In_153);
nor U104 (N_104,In_297,In_247);
nor U105 (N_105,In_402,In_137);
nand U106 (N_106,In_243,In_360);
nor U107 (N_107,In_435,In_125);
nand U108 (N_108,In_72,In_490);
nor U109 (N_109,In_288,In_79);
or U110 (N_110,In_180,In_472);
xor U111 (N_111,In_146,In_261);
or U112 (N_112,In_452,In_278);
or U113 (N_113,In_202,In_303);
or U114 (N_114,In_178,In_494);
or U115 (N_115,In_434,In_235);
and U116 (N_116,In_462,In_228);
nor U117 (N_117,In_3,In_323);
and U118 (N_118,In_305,In_428);
nand U119 (N_119,In_132,In_369);
or U120 (N_120,In_386,In_193);
and U121 (N_121,In_204,In_44);
nand U122 (N_122,In_336,In_357);
or U123 (N_123,In_47,In_69);
nand U124 (N_124,In_350,In_498);
and U125 (N_125,In_104,In_144);
xnor U126 (N_126,In_425,In_370);
nand U127 (N_127,In_216,In_359);
nor U128 (N_128,In_82,In_91);
and U129 (N_129,In_252,In_280);
nand U130 (N_130,In_332,In_113);
nor U131 (N_131,In_119,In_275);
nor U132 (N_132,In_383,In_143);
nor U133 (N_133,In_92,In_491);
nand U134 (N_134,In_344,In_320);
and U135 (N_135,In_234,In_8);
and U136 (N_136,In_258,In_240);
and U137 (N_137,In_394,In_195);
nand U138 (N_138,In_273,In_7);
nand U139 (N_139,In_361,In_416);
nor U140 (N_140,In_68,In_83);
nor U141 (N_141,In_446,In_80);
and U142 (N_142,In_36,In_161);
nand U143 (N_143,In_105,In_53);
nand U144 (N_144,In_371,In_15);
nand U145 (N_145,In_373,In_149);
or U146 (N_146,In_423,In_99);
nand U147 (N_147,In_290,In_315);
or U148 (N_148,In_114,In_438);
nand U149 (N_149,In_199,In_20);
and U150 (N_150,In_274,In_37);
nor U151 (N_151,In_306,In_57);
nand U152 (N_152,In_269,In_421);
nand U153 (N_153,In_176,In_447);
nor U154 (N_154,In_102,In_455);
xnor U155 (N_155,In_232,In_312);
nand U156 (N_156,In_134,In_254);
or U157 (N_157,In_349,In_181);
or U158 (N_158,In_449,In_122);
nor U159 (N_159,In_488,In_253);
nand U160 (N_160,In_25,In_375);
nor U161 (N_161,In_231,In_207);
and U162 (N_162,In_158,In_126);
nand U163 (N_163,In_224,In_392);
nand U164 (N_164,In_177,In_130);
or U165 (N_165,In_115,In_399);
or U166 (N_166,In_162,In_284);
or U167 (N_167,In_276,In_108);
and U168 (N_168,In_117,In_346);
nor U169 (N_169,In_403,In_257);
or U170 (N_170,In_106,In_31);
nand U171 (N_171,In_337,In_354);
nand U172 (N_172,In_291,In_341);
nand U173 (N_173,In_110,In_295);
or U174 (N_174,In_39,In_411);
or U175 (N_175,In_222,In_184);
or U176 (N_176,In_101,In_225);
or U177 (N_177,In_1,In_4);
or U178 (N_178,In_98,In_85);
nand U179 (N_179,In_73,In_81);
or U180 (N_180,In_169,In_150);
nand U181 (N_181,In_187,In_474);
or U182 (N_182,In_48,In_154);
nand U183 (N_183,In_405,In_309);
and U184 (N_184,In_484,In_308);
xor U185 (N_185,In_131,In_218);
nor U186 (N_186,In_192,In_135);
nor U187 (N_187,In_334,In_453);
nor U188 (N_188,In_245,In_244);
and U189 (N_189,In_368,In_64);
nand U190 (N_190,In_466,In_66);
nor U191 (N_191,In_185,In_263);
and U192 (N_192,In_338,In_391);
or U193 (N_193,In_89,In_356);
nand U194 (N_194,In_282,In_163);
nor U195 (N_195,In_26,In_220);
nor U196 (N_196,In_468,In_183);
nor U197 (N_197,In_372,In_242);
or U198 (N_198,In_256,In_377);
or U199 (N_199,In_5,In_46);
and U200 (N_200,N_19,In_236);
nor U201 (N_201,In_97,N_102);
nand U202 (N_202,N_157,N_42);
nor U203 (N_203,N_55,N_9);
nand U204 (N_204,In_445,In_112);
nand U205 (N_205,N_186,N_85);
nand U206 (N_206,N_58,N_40);
nand U207 (N_207,N_45,In_364);
and U208 (N_208,N_114,In_95);
nand U209 (N_209,N_133,In_197);
nand U210 (N_210,N_194,N_127);
nor U211 (N_211,N_23,N_173);
or U212 (N_212,In_61,In_10);
and U213 (N_213,N_162,N_138);
and U214 (N_214,N_92,N_132);
nor U215 (N_215,N_71,In_128);
nand U216 (N_216,N_165,In_142);
or U217 (N_217,In_326,N_119);
and U218 (N_218,In_6,N_100);
nor U219 (N_219,In_264,N_116);
or U220 (N_220,In_221,N_123);
nand U221 (N_221,N_60,In_87);
nand U222 (N_222,N_151,N_128);
nor U223 (N_223,N_150,In_286);
and U224 (N_224,In_437,In_351);
or U225 (N_225,In_345,N_110);
nor U226 (N_226,In_479,In_11);
or U227 (N_227,N_17,N_158);
nand U228 (N_228,N_73,N_15);
and U229 (N_229,N_129,N_122);
and U230 (N_230,N_37,In_40);
nand U231 (N_231,N_166,N_164);
nand U232 (N_232,In_226,N_44);
and U233 (N_233,N_36,In_443);
or U234 (N_234,In_289,In_78);
nor U235 (N_235,In_478,N_117);
and U236 (N_236,In_277,In_417);
or U237 (N_237,N_6,In_450);
and U238 (N_238,N_181,N_198);
and U239 (N_239,In_60,N_65);
or U240 (N_240,N_147,N_105);
nor U241 (N_241,N_88,N_139);
and U242 (N_242,In_329,N_191);
nor U243 (N_243,In_160,N_176);
and U244 (N_244,N_79,N_97);
and U245 (N_245,In_230,N_14);
nand U246 (N_246,In_495,N_112);
or U247 (N_247,N_90,In_444);
nand U248 (N_248,N_149,In_2);
nand U249 (N_249,N_51,N_48);
nand U250 (N_250,In_475,N_56);
and U251 (N_251,In_65,In_379);
nor U252 (N_252,N_167,In_155);
nand U253 (N_253,In_422,N_10);
or U254 (N_254,In_300,N_61);
nor U255 (N_255,N_29,N_134);
or U256 (N_256,In_203,In_186);
and U257 (N_257,In_461,N_103);
nor U258 (N_258,N_32,N_141);
nand U259 (N_259,In_409,N_188);
and U260 (N_260,N_190,N_84);
or U261 (N_261,N_1,In_116);
and U262 (N_262,N_136,N_13);
nand U263 (N_263,In_29,N_67);
nand U264 (N_264,N_124,In_30);
and U265 (N_265,N_24,N_75);
nand U266 (N_266,N_22,N_159);
or U267 (N_267,N_155,N_185);
or U268 (N_268,N_46,N_35);
nor U269 (N_269,N_77,N_50);
nor U270 (N_270,N_74,N_131);
and U271 (N_271,N_57,N_98);
nor U272 (N_272,N_156,N_3);
or U273 (N_273,N_80,N_152);
or U274 (N_274,N_93,N_39);
xnor U275 (N_275,In_145,N_120);
nand U276 (N_276,N_0,N_2);
nand U277 (N_277,N_163,N_30);
and U278 (N_278,In_147,N_38);
nor U279 (N_279,N_96,N_183);
or U280 (N_280,N_168,In_311);
nand U281 (N_281,N_21,In_43);
or U282 (N_282,N_82,N_101);
or U283 (N_283,N_81,In_56);
nand U284 (N_284,N_199,N_66);
nand U285 (N_285,N_28,In_270);
and U286 (N_286,N_27,N_178);
and U287 (N_287,N_113,In_103);
nor U288 (N_288,N_26,In_127);
nand U289 (N_289,In_219,In_458);
nor U290 (N_290,In_398,In_271);
and U291 (N_291,In_477,N_94);
and U292 (N_292,N_111,N_78);
nand U293 (N_293,N_125,N_41);
nand U294 (N_294,N_121,N_86);
nor U295 (N_295,N_4,N_144);
nor U296 (N_296,In_70,N_146);
xor U297 (N_297,N_148,N_64);
nor U298 (N_298,In_464,N_16);
nand U299 (N_299,N_143,N_72);
and U300 (N_300,N_177,N_172);
nor U301 (N_301,N_175,N_12);
or U302 (N_302,In_239,N_197);
and U303 (N_303,N_68,In_0);
nand U304 (N_304,N_135,In_381);
nor U305 (N_305,N_109,In_13);
nand U306 (N_306,N_99,In_426);
nor U307 (N_307,N_49,N_187);
and U308 (N_308,N_179,In_19);
and U309 (N_309,N_43,In_151);
nor U310 (N_310,N_115,In_18);
nor U311 (N_311,N_7,In_191);
nor U312 (N_312,N_192,N_154);
nand U313 (N_313,N_130,N_70);
and U314 (N_314,N_137,N_196);
nand U315 (N_315,N_31,N_47);
or U316 (N_316,N_59,N_180);
and U317 (N_317,N_11,N_20);
or U318 (N_318,N_171,In_174);
nand U319 (N_319,N_161,In_260);
and U320 (N_320,In_415,N_108);
and U321 (N_321,N_25,N_182);
or U322 (N_322,N_62,In_138);
and U323 (N_323,N_53,N_95);
or U324 (N_324,In_266,N_63);
and U325 (N_325,N_33,In_215);
nor U326 (N_326,N_189,N_107);
nor U327 (N_327,In_378,In_173);
or U328 (N_328,In_406,N_160);
xor U329 (N_329,N_54,N_184);
nor U330 (N_330,N_145,N_118);
nor U331 (N_331,N_52,N_87);
and U332 (N_332,N_140,In_45);
nor U333 (N_333,N_89,N_76);
or U334 (N_334,In_62,In_35);
and U335 (N_335,In_397,In_251);
or U336 (N_336,In_23,In_430);
nor U337 (N_337,N_153,In_262);
or U338 (N_338,N_126,In_439);
nand U339 (N_339,In_28,N_18);
nor U340 (N_340,In_451,N_8);
and U341 (N_341,N_83,N_195);
nand U342 (N_342,N_169,N_170);
or U343 (N_343,N_142,In_152);
or U344 (N_344,N_104,N_5);
or U345 (N_345,N_174,In_205);
and U346 (N_346,In_248,In_211);
nand U347 (N_347,N_69,N_91);
and U348 (N_348,In_84,N_106);
nor U349 (N_349,N_34,N_193);
nor U350 (N_350,N_37,N_154);
and U351 (N_351,N_78,N_110);
and U352 (N_352,N_81,N_60);
nor U353 (N_353,N_93,N_117);
and U354 (N_354,In_35,In_138);
nand U355 (N_355,N_149,N_140);
and U356 (N_356,N_54,N_189);
and U357 (N_357,N_67,In_0);
nor U358 (N_358,N_52,In_23);
nand U359 (N_359,N_88,In_226);
nand U360 (N_360,N_151,N_26);
nand U361 (N_361,N_141,In_300);
or U362 (N_362,N_133,N_137);
nand U363 (N_363,N_95,N_194);
nor U364 (N_364,N_137,In_381);
nand U365 (N_365,In_84,N_186);
nor U366 (N_366,N_155,In_329);
xnor U367 (N_367,N_95,N_2);
or U368 (N_368,N_107,In_479);
nand U369 (N_369,N_88,In_458);
or U370 (N_370,In_142,N_153);
or U371 (N_371,In_329,N_111);
and U372 (N_372,N_136,In_230);
nand U373 (N_373,N_173,N_95);
and U374 (N_374,N_89,In_406);
nand U375 (N_375,N_41,N_2);
and U376 (N_376,N_133,N_111);
or U377 (N_377,N_31,N_176);
and U378 (N_378,N_90,N_30);
or U379 (N_379,N_13,N_88);
nor U380 (N_380,N_41,N_189);
xor U381 (N_381,N_185,In_495);
or U382 (N_382,N_177,N_196);
nand U383 (N_383,N_177,N_155);
and U384 (N_384,N_142,In_445);
or U385 (N_385,N_134,N_55);
nand U386 (N_386,N_113,N_38);
nand U387 (N_387,N_179,N_31);
nor U388 (N_388,N_49,N_60);
nand U389 (N_389,N_171,In_142);
nand U390 (N_390,In_62,N_47);
nor U391 (N_391,N_53,N_3);
and U392 (N_392,N_156,N_50);
and U393 (N_393,N_171,N_122);
nand U394 (N_394,N_169,In_479);
nor U395 (N_395,In_11,In_197);
or U396 (N_396,In_28,In_60);
or U397 (N_397,N_158,N_3);
or U398 (N_398,N_192,N_118);
or U399 (N_399,In_6,N_81);
and U400 (N_400,N_311,N_365);
and U401 (N_401,N_339,N_298);
nor U402 (N_402,N_256,N_215);
or U403 (N_403,N_314,N_398);
nor U404 (N_404,N_348,N_377);
and U405 (N_405,N_237,N_336);
nor U406 (N_406,N_393,N_276);
nor U407 (N_407,N_244,N_259);
and U408 (N_408,N_257,N_304);
nand U409 (N_409,N_219,N_380);
or U410 (N_410,N_204,N_223);
nor U411 (N_411,N_356,N_310);
nand U412 (N_412,N_296,N_373);
and U413 (N_413,N_246,N_224);
or U414 (N_414,N_233,N_382);
and U415 (N_415,N_289,N_331);
xor U416 (N_416,N_273,N_333);
nand U417 (N_417,N_258,N_355);
and U418 (N_418,N_260,N_302);
nor U419 (N_419,N_201,N_369);
or U420 (N_420,N_230,N_313);
nand U421 (N_421,N_252,N_375);
nor U422 (N_422,N_278,N_294);
nand U423 (N_423,N_324,N_293);
or U424 (N_424,N_280,N_290);
nor U425 (N_425,N_255,N_345);
nor U426 (N_426,N_216,N_297);
nor U427 (N_427,N_226,N_202);
nand U428 (N_428,N_270,N_374);
nand U429 (N_429,N_272,N_330);
or U430 (N_430,N_378,N_238);
and U431 (N_431,N_225,N_325);
or U432 (N_432,N_389,N_207);
nand U433 (N_433,N_309,N_337);
or U434 (N_434,N_267,N_291);
nor U435 (N_435,N_399,N_274);
nand U436 (N_436,N_253,N_396);
nand U437 (N_437,N_240,N_248);
nand U438 (N_438,N_303,N_235);
and U439 (N_439,N_221,N_352);
nand U440 (N_440,N_367,N_364);
nor U441 (N_441,N_227,N_203);
nor U442 (N_442,N_301,N_214);
nor U443 (N_443,N_218,N_368);
or U444 (N_444,N_229,N_329);
xor U445 (N_445,N_359,N_236);
and U446 (N_446,N_379,N_288);
nor U447 (N_447,N_323,N_232);
nor U448 (N_448,N_354,N_350);
and U449 (N_449,N_322,N_360);
nand U450 (N_450,N_390,N_231);
or U451 (N_451,N_282,N_334);
nor U452 (N_452,N_284,N_318);
nand U453 (N_453,N_279,N_383);
or U454 (N_454,N_264,N_209);
nor U455 (N_455,N_239,N_315);
nor U456 (N_456,N_287,N_376);
and U457 (N_457,N_372,N_254);
and U458 (N_458,N_245,N_327);
and U459 (N_459,N_312,N_205);
and U460 (N_460,N_361,N_387);
nand U461 (N_461,N_261,N_321);
nand U462 (N_462,N_332,N_307);
or U463 (N_463,N_292,N_249);
and U464 (N_464,N_341,N_206);
nor U465 (N_465,N_308,N_281);
nand U466 (N_466,N_299,N_271);
or U467 (N_467,N_262,N_358);
nand U468 (N_468,N_228,N_338);
nand U469 (N_469,N_397,N_266);
or U470 (N_470,N_384,N_320);
nor U471 (N_471,N_328,N_213);
and U472 (N_472,N_222,N_316);
nand U473 (N_473,N_392,N_212);
or U474 (N_474,N_295,N_286);
nor U475 (N_475,N_394,N_351);
nand U476 (N_476,N_251,N_388);
nand U477 (N_477,N_317,N_347);
or U478 (N_478,N_217,N_241);
and U479 (N_479,N_268,N_305);
or U480 (N_480,N_391,N_371);
nor U481 (N_481,N_386,N_342);
nor U482 (N_482,N_269,N_340);
or U483 (N_483,N_250,N_319);
or U484 (N_484,N_335,N_275);
nand U485 (N_485,N_349,N_208);
nor U486 (N_486,N_243,N_381);
nor U487 (N_487,N_283,N_343);
nor U488 (N_488,N_395,N_242);
and U489 (N_489,N_211,N_200);
xor U490 (N_490,N_344,N_363);
nor U491 (N_491,N_326,N_385);
nor U492 (N_492,N_234,N_220);
xor U493 (N_493,N_306,N_366);
nor U494 (N_494,N_210,N_247);
nor U495 (N_495,N_277,N_357);
and U496 (N_496,N_370,N_346);
nand U497 (N_497,N_263,N_362);
xnor U498 (N_498,N_265,N_300);
or U499 (N_499,N_353,N_285);
nand U500 (N_500,N_379,N_256);
nand U501 (N_501,N_217,N_338);
and U502 (N_502,N_210,N_348);
and U503 (N_503,N_332,N_337);
and U504 (N_504,N_300,N_251);
nand U505 (N_505,N_384,N_281);
or U506 (N_506,N_205,N_267);
nand U507 (N_507,N_339,N_340);
and U508 (N_508,N_351,N_345);
nand U509 (N_509,N_205,N_327);
and U510 (N_510,N_251,N_223);
nor U511 (N_511,N_222,N_243);
or U512 (N_512,N_299,N_346);
and U513 (N_513,N_279,N_351);
and U514 (N_514,N_214,N_236);
or U515 (N_515,N_333,N_334);
nor U516 (N_516,N_219,N_394);
or U517 (N_517,N_346,N_209);
and U518 (N_518,N_301,N_360);
nand U519 (N_519,N_371,N_239);
nand U520 (N_520,N_322,N_201);
xnor U521 (N_521,N_226,N_270);
or U522 (N_522,N_334,N_386);
and U523 (N_523,N_278,N_349);
and U524 (N_524,N_253,N_382);
and U525 (N_525,N_337,N_286);
or U526 (N_526,N_204,N_393);
and U527 (N_527,N_202,N_372);
and U528 (N_528,N_328,N_226);
or U529 (N_529,N_344,N_302);
and U530 (N_530,N_238,N_231);
or U531 (N_531,N_371,N_235);
or U532 (N_532,N_377,N_311);
or U533 (N_533,N_212,N_281);
or U534 (N_534,N_297,N_392);
and U535 (N_535,N_204,N_363);
nand U536 (N_536,N_231,N_355);
nor U537 (N_537,N_386,N_210);
and U538 (N_538,N_214,N_225);
and U539 (N_539,N_300,N_327);
nand U540 (N_540,N_263,N_378);
nor U541 (N_541,N_269,N_226);
or U542 (N_542,N_393,N_271);
or U543 (N_543,N_366,N_284);
and U544 (N_544,N_358,N_391);
nor U545 (N_545,N_285,N_271);
and U546 (N_546,N_218,N_328);
or U547 (N_547,N_362,N_314);
nand U548 (N_548,N_379,N_382);
or U549 (N_549,N_399,N_324);
and U550 (N_550,N_281,N_341);
and U551 (N_551,N_286,N_206);
nor U552 (N_552,N_230,N_271);
nor U553 (N_553,N_205,N_277);
nor U554 (N_554,N_332,N_308);
nand U555 (N_555,N_214,N_229);
nand U556 (N_556,N_256,N_309);
or U557 (N_557,N_271,N_344);
or U558 (N_558,N_377,N_252);
and U559 (N_559,N_381,N_291);
or U560 (N_560,N_385,N_261);
or U561 (N_561,N_378,N_374);
or U562 (N_562,N_364,N_336);
nor U563 (N_563,N_308,N_220);
or U564 (N_564,N_313,N_287);
and U565 (N_565,N_323,N_388);
or U566 (N_566,N_255,N_268);
or U567 (N_567,N_321,N_305);
or U568 (N_568,N_346,N_285);
nand U569 (N_569,N_260,N_272);
and U570 (N_570,N_370,N_252);
nand U571 (N_571,N_360,N_200);
nor U572 (N_572,N_348,N_239);
or U573 (N_573,N_341,N_222);
nand U574 (N_574,N_229,N_358);
or U575 (N_575,N_351,N_300);
or U576 (N_576,N_263,N_357);
and U577 (N_577,N_326,N_265);
nand U578 (N_578,N_392,N_314);
nor U579 (N_579,N_262,N_283);
nand U580 (N_580,N_373,N_378);
nand U581 (N_581,N_367,N_368);
or U582 (N_582,N_234,N_284);
nor U583 (N_583,N_399,N_360);
or U584 (N_584,N_373,N_251);
nor U585 (N_585,N_233,N_300);
nand U586 (N_586,N_307,N_326);
or U587 (N_587,N_278,N_338);
and U588 (N_588,N_221,N_241);
and U589 (N_589,N_306,N_245);
nand U590 (N_590,N_373,N_238);
and U591 (N_591,N_377,N_230);
or U592 (N_592,N_245,N_314);
nand U593 (N_593,N_304,N_242);
nand U594 (N_594,N_200,N_295);
and U595 (N_595,N_248,N_251);
and U596 (N_596,N_322,N_304);
nor U597 (N_597,N_384,N_361);
or U598 (N_598,N_317,N_253);
and U599 (N_599,N_293,N_253);
xnor U600 (N_600,N_404,N_474);
and U601 (N_601,N_458,N_594);
nor U602 (N_602,N_540,N_445);
or U603 (N_603,N_542,N_441);
nor U604 (N_604,N_553,N_522);
and U605 (N_605,N_541,N_578);
or U606 (N_606,N_572,N_454);
nand U607 (N_607,N_567,N_519);
nor U608 (N_608,N_480,N_587);
nor U609 (N_609,N_536,N_426);
nand U610 (N_610,N_537,N_510);
nor U611 (N_611,N_416,N_509);
nor U612 (N_612,N_478,N_508);
nor U613 (N_613,N_492,N_422);
nor U614 (N_614,N_483,N_588);
nor U615 (N_615,N_462,N_581);
nor U616 (N_616,N_544,N_576);
nand U617 (N_617,N_534,N_439);
and U618 (N_618,N_423,N_412);
nor U619 (N_619,N_453,N_438);
and U620 (N_620,N_477,N_402);
or U621 (N_621,N_475,N_467);
and U622 (N_622,N_575,N_433);
nand U623 (N_623,N_507,N_463);
and U624 (N_624,N_574,N_531);
nand U625 (N_625,N_599,N_443);
and U626 (N_626,N_484,N_500);
or U627 (N_627,N_409,N_499);
nand U628 (N_628,N_518,N_473);
nand U629 (N_629,N_569,N_494);
nand U630 (N_630,N_429,N_592);
nand U631 (N_631,N_414,N_558);
and U632 (N_632,N_425,N_591);
nor U633 (N_633,N_543,N_551);
nand U634 (N_634,N_504,N_403);
xor U635 (N_635,N_456,N_582);
nor U636 (N_636,N_580,N_472);
nand U637 (N_637,N_464,N_546);
or U638 (N_638,N_550,N_589);
nor U639 (N_639,N_503,N_552);
nand U640 (N_640,N_530,N_523);
nand U641 (N_641,N_533,N_513);
or U642 (N_642,N_532,N_469);
or U643 (N_643,N_459,N_535);
or U644 (N_644,N_421,N_548);
nand U645 (N_645,N_547,N_496);
and U646 (N_646,N_442,N_579);
or U647 (N_647,N_559,N_471);
nand U648 (N_648,N_596,N_420);
and U649 (N_649,N_562,N_432);
or U650 (N_650,N_526,N_449);
nor U651 (N_651,N_498,N_495);
nor U652 (N_652,N_525,N_529);
or U653 (N_653,N_448,N_466);
nor U654 (N_654,N_512,N_515);
nor U655 (N_655,N_517,N_407);
xnor U656 (N_656,N_460,N_430);
and U657 (N_657,N_410,N_444);
nor U658 (N_658,N_408,N_447);
nor U659 (N_659,N_598,N_501);
nand U660 (N_660,N_584,N_493);
and U661 (N_661,N_557,N_417);
nand U662 (N_662,N_406,N_590);
or U663 (N_663,N_468,N_450);
nand U664 (N_664,N_524,N_505);
and U665 (N_665,N_565,N_497);
or U666 (N_666,N_405,N_597);
nor U667 (N_667,N_465,N_489);
nand U668 (N_668,N_427,N_586);
nand U669 (N_669,N_506,N_573);
nor U670 (N_670,N_555,N_440);
xor U671 (N_671,N_561,N_485);
or U672 (N_672,N_539,N_560);
nor U673 (N_673,N_491,N_437);
or U674 (N_674,N_446,N_455);
and U675 (N_675,N_556,N_424);
and U676 (N_676,N_470,N_434);
xnor U677 (N_677,N_564,N_511);
or U678 (N_678,N_593,N_585);
or U679 (N_679,N_419,N_538);
nand U680 (N_680,N_583,N_413);
nand U681 (N_681,N_514,N_487);
nor U682 (N_682,N_479,N_566);
and U683 (N_683,N_482,N_481);
and U684 (N_684,N_570,N_502);
nand U685 (N_685,N_435,N_418);
nand U686 (N_686,N_521,N_461);
nand U687 (N_687,N_545,N_488);
or U688 (N_688,N_490,N_415);
and U689 (N_689,N_520,N_411);
or U690 (N_690,N_595,N_428);
and U691 (N_691,N_568,N_476);
nor U692 (N_692,N_436,N_571);
nand U693 (N_693,N_528,N_516);
nand U694 (N_694,N_549,N_486);
or U695 (N_695,N_431,N_401);
and U696 (N_696,N_457,N_577);
nor U697 (N_697,N_452,N_400);
and U698 (N_698,N_554,N_527);
or U699 (N_699,N_563,N_451);
nor U700 (N_700,N_514,N_442);
and U701 (N_701,N_570,N_584);
and U702 (N_702,N_481,N_415);
or U703 (N_703,N_512,N_493);
nand U704 (N_704,N_441,N_448);
or U705 (N_705,N_510,N_482);
nor U706 (N_706,N_538,N_497);
or U707 (N_707,N_493,N_454);
and U708 (N_708,N_583,N_521);
or U709 (N_709,N_562,N_445);
or U710 (N_710,N_557,N_564);
or U711 (N_711,N_431,N_406);
nand U712 (N_712,N_485,N_407);
nand U713 (N_713,N_533,N_450);
nand U714 (N_714,N_526,N_508);
or U715 (N_715,N_433,N_410);
nor U716 (N_716,N_579,N_411);
nand U717 (N_717,N_538,N_568);
or U718 (N_718,N_436,N_425);
nor U719 (N_719,N_477,N_464);
and U720 (N_720,N_444,N_438);
nor U721 (N_721,N_560,N_417);
and U722 (N_722,N_497,N_559);
nor U723 (N_723,N_555,N_419);
or U724 (N_724,N_596,N_482);
and U725 (N_725,N_437,N_447);
nand U726 (N_726,N_430,N_594);
or U727 (N_727,N_463,N_530);
or U728 (N_728,N_481,N_456);
nor U729 (N_729,N_456,N_453);
nand U730 (N_730,N_405,N_455);
nand U731 (N_731,N_416,N_537);
or U732 (N_732,N_547,N_475);
nand U733 (N_733,N_453,N_579);
and U734 (N_734,N_469,N_596);
nand U735 (N_735,N_494,N_499);
and U736 (N_736,N_492,N_476);
nand U737 (N_737,N_595,N_567);
nand U738 (N_738,N_453,N_546);
and U739 (N_739,N_530,N_527);
or U740 (N_740,N_540,N_447);
or U741 (N_741,N_446,N_462);
and U742 (N_742,N_561,N_589);
or U743 (N_743,N_585,N_594);
nand U744 (N_744,N_467,N_483);
and U745 (N_745,N_498,N_435);
nor U746 (N_746,N_412,N_508);
and U747 (N_747,N_543,N_482);
nand U748 (N_748,N_563,N_497);
and U749 (N_749,N_411,N_499);
or U750 (N_750,N_444,N_477);
and U751 (N_751,N_579,N_440);
or U752 (N_752,N_598,N_507);
nor U753 (N_753,N_464,N_589);
or U754 (N_754,N_578,N_588);
or U755 (N_755,N_474,N_511);
nor U756 (N_756,N_580,N_443);
nor U757 (N_757,N_571,N_520);
nand U758 (N_758,N_583,N_520);
xnor U759 (N_759,N_592,N_556);
nand U760 (N_760,N_458,N_583);
nor U761 (N_761,N_509,N_505);
xnor U762 (N_762,N_579,N_506);
nor U763 (N_763,N_500,N_466);
xnor U764 (N_764,N_438,N_577);
nor U765 (N_765,N_576,N_407);
nor U766 (N_766,N_518,N_464);
nand U767 (N_767,N_472,N_410);
nand U768 (N_768,N_567,N_438);
and U769 (N_769,N_529,N_492);
nand U770 (N_770,N_452,N_530);
nand U771 (N_771,N_473,N_558);
or U772 (N_772,N_554,N_448);
nand U773 (N_773,N_458,N_402);
nor U774 (N_774,N_494,N_529);
nor U775 (N_775,N_510,N_591);
nand U776 (N_776,N_521,N_589);
nand U777 (N_777,N_530,N_587);
nor U778 (N_778,N_456,N_512);
and U779 (N_779,N_431,N_468);
nor U780 (N_780,N_457,N_471);
nand U781 (N_781,N_436,N_536);
nand U782 (N_782,N_583,N_472);
or U783 (N_783,N_541,N_560);
or U784 (N_784,N_440,N_490);
nor U785 (N_785,N_594,N_451);
or U786 (N_786,N_478,N_496);
or U787 (N_787,N_406,N_591);
and U788 (N_788,N_445,N_590);
nand U789 (N_789,N_582,N_564);
nand U790 (N_790,N_408,N_464);
and U791 (N_791,N_572,N_555);
xnor U792 (N_792,N_538,N_547);
nor U793 (N_793,N_521,N_439);
nor U794 (N_794,N_524,N_534);
xor U795 (N_795,N_439,N_557);
or U796 (N_796,N_576,N_496);
nor U797 (N_797,N_583,N_484);
nor U798 (N_798,N_555,N_431);
nand U799 (N_799,N_570,N_524);
nor U800 (N_800,N_636,N_744);
nand U801 (N_801,N_656,N_667);
nand U802 (N_802,N_726,N_645);
or U803 (N_803,N_790,N_612);
nand U804 (N_804,N_725,N_673);
and U805 (N_805,N_628,N_663);
and U806 (N_806,N_601,N_642);
and U807 (N_807,N_788,N_686);
nor U808 (N_808,N_734,N_662);
nand U809 (N_809,N_660,N_730);
or U810 (N_810,N_649,N_614);
and U811 (N_811,N_625,N_650);
nand U812 (N_812,N_707,N_626);
nand U813 (N_813,N_631,N_613);
nor U814 (N_814,N_709,N_648);
nor U815 (N_815,N_701,N_798);
nor U816 (N_816,N_705,N_685);
nor U817 (N_817,N_780,N_756);
nor U818 (N_818,N_671,N_658);
and U819 (N_819,N_773,N_794);
xnor U820 (N_820,N_721,N_779);
and U821 (N_821,N_682,N_711);
or U822 (N_822,N_633,N_742);
nor U823 (N_823,N_710,N_670);
and U824 (N_824,N_740,N_616);
or U825 (N_825,N_694,N_702);
nor U826 (N_826,N_713,N_715);
and U827 (N_827,N_760,N_785);
nor U828 (N_828,N_706,N_752);
xnor U829 (N_829,N_789,N_718);
and U830 (N_830,N_659,N_772);
nand U831 (N_831,N_623,N_606);
nand U832 (N_832,N_716,N_723);
nor U833 (N_833,N_704,N_635);
or U834 (N_834,N_683,N_765);
or U835 (N_835,N_728,N_666);
nor U836 (N_836,N_607,N_754);
nor U837 (N_837,N_678,N_796);
nand U838 (N_838,N_675,N_768);
and U839 (N_839,N_687,N_783);
nand U840 (N_840,N_620,N_795);
nand U841 (N_841,N_605,N_776);
or U842 (N_842,N_655,N_712);
nor U843 (N_843,N_639,N_689);
nor U844 (N_844,N_755,N_695);
xnor U845 (N_845,N_745,N_753);
nand U846 (N_846,N_698,N_781);
nand U847 (N_847,N_684,N_646);
nor U848 (N_848,N_652,N_799);
xnor U849 (N_849,N_750,N_629);
and U850 (N_850,N_737,N_632);
nand U851 (N_851,N_643,N_657);
or U852 (N_852,N_699,N_722);
or U853 (N_853,N_778,N_630);
nor U854 (N_854,N_791,N_664);
and U855 (N_855,N_770,N_775);
nand U856 (N_856,N_681,N_729);
or U857 (N_857,N_766,N_787);
and U858 (N_858,N_792,N_677);
and U859 (N_859,N_661,N_761);
and U860 (N_860,N_604,N_622);
nor U861 (N_861,N_621,N_708);
and U862 (N_862,N_724,N_700);
nand U863 (N_863,N_774,N_647);
or U864 (N_864,N_600,N_674);
or U865 (N_865,N_786,N_609);
nand U866 (N_866,N_692,N_727);
or U867 (N_867,N_797,N_651);
nand U868 (N_868,N_793,N_668);
nor U869 (N_869,N_624,N_676);
and U870 (N_870,N_617,N_777);
and U871 (N_871,N_736,N_611);
and U872 (N_872,N_743,N_746);
nand U873 (N_873,N_720,N_738);
nand U874 (N_874,N_619,N_690);
nor U875 (N_875,N_758,N_782);
or U876 (N_876,N_618,N_747);
nand U877 (N_877,N_771,N_693);
and U878 (N_878,N_769,N_669);
nand U879 (N_879,N_731,N_732);
or U880 (N_880,N_688,N_757);
nor U881 (N_881,N_653,N_665);
nor U882 (N_882,N_759,N_640);
nand U883 (N_883,N_679,N_641);
nand U884 (N_884,N_719,N_638);
and U885 (N_885,N_784,N_691);
nor U886 (N_886,N_697,N_696);
and U887 (N_887,N_735,N_703);
and U888 (N_888,N_748,N_672);
or U889 (N_889,N_739,N_634);
nand U890 (N_890,N_717,N_615);
nor U891 (N_891,N_603,N_749);
nand U892 (N_892,N_762,N_637);
or U893 (N_893,N_680,N_654);
xor U894 (N_894,N_763,N_602);
nand U895 (N_895,N_714,N_764);
nand U896 (N_896,N_644,N_767);
nand U897 (N_897,N_751,N_627);
nor U898 (N_898,N_608,N_741);
nor U899 (N_899,N_610,N_733);
or U900 (N_900,N_785,N_629);
or U901 (N_901,N_714,N_648);
nor U902 (N_902,N_793,N_792);
nand U903 (N_903,N_768,N_747);
and U904 (N_904,N_619,N_623);
nor U905 (N_905,N_685,N_683);
nor U906 (N_906,N_742,N_741);
and U907 (N_907,N_606,N_696);
nand U908 (N_908,N_661,N_627);
xnor U909 (N_909,N_774,N_799);
and U910 (N_910,N_639,N_732);
nor U911 (N_911,N_741,N_663);
nor U912 (N_912,N_686,N_663);
nor U913 (N_913,N_782,N_718);
nor U914 (N_914,N_766,N_651);
nor U915 (N_915,N_683,N_630);
and U916 (N_916,N_665,N_715);
and U917 (N_917,N_773,N_734);
nand U918 (N_918,N_654,N_746);
nor U919 (N_919,N_630,N_691);
nor U920 (N_920,N_790,N_765);
nor U921 (N_921,N_772,N_790);
nand U922 (N_922,N_798,N_717);
nor U923 (N_923,N_702,N_721);
or U924 (N_924,N_664,N_781);
and U925 (N_925,N_656,N_735);
and U926 (N_926,N_629,N_704);
nand U927 (N_927,N_633,N_660);
or U928 (N_928,N_790,N_731);
nor U929 (N_929,N_616,N_796);
and U930 (N_930,N_698,N_719);
and U931 (N_931,N_730,N_711);
and U932 (N_932,N_783,N_713);
and U933 (N_933,N_665,N_756);
or U934 (N_934,N_651,N_625);
nand U935 (N_935,N_763,N_791);
nand U936 (N_936,N_703,N_627);
nand U937 (N_937,N_786,N_717);
and U938 (N_938,N_708,N_616);
and U939 (N_939,N_673,N_690);
or U940 (N_940,N_700,N_626);
nor U941 (N_941,N_771,N_732);
nor U942 (N_942,N_711,N_742);
and U943 (N_943,N_680,N_763);
nand U944 (N_944,N_776,N_672);
and U945 (N_945,N_741,N_616);
nand U946 (N_946,N_624,N_798);
nand U947 (N_947,N_744,N_781);
and U948 (N_948,N_607,N_619);
or U949 (N_949,N_781,N_674);
nand U950 (N_950,N_779,N_653);
or U951 (N_951,N_795,N_670);
nor U952 (N_952,N_659,N_603);
xnor U953 (N_953,N_762,N_746);
nor U954 (N_954,N_787,N_611);
nor U955 (N_955,N_767,N_635);
nor U956 (N_956,N_760,N_744);
nor U957 (N_957,N_669,N_698);
and U958 (N_958,N_633,N_786);
and U959 (N_959,N_792,N_687);
or U960 (N_960,N_632,N_616);
and U961 (N_961,N_638,N_683);
or U962 (N_962,N_782,N_779);
and U963 (N_963,N_651,N_693);
nand U964 (N_964,N_736,N_708);
nand U965 (N_965,N_620,N_694);
nand U966 (N_966,N_601,N_759);
or U967 (N_967,N_719,N_633);
or U968 (N_968,N_701,N_720);
xnor U969 (N_969,N_615,N_771);
nor U970 (N_970,N_771,N_686);
nor U971 (N_971,N_712,N_746);
or U972 (N_972,N_611,N_752);
xor U973 (N_973,N_606,N_669);
nand U974 (N_974,N_695,N_639);
and U975 (N_975,N_702,N_637);
nor U976 (N_976,N_656,N_694);
nand U977 (N_977,N_628,N_635);
or U978 (N_978,N_706,N_739);
nor U979 (N_979,N_611,N_648);
nor U980 (N_980,N_637,N_686);
and U981 (N_981,N_685,N_726);
and U982 (N_982,N_621,N_640);
and U983 (N_983,N_789,N_731);
or U984 (N_984,N_734,N_690);
nor U985 (N_985,N_604,N_712);
and U986 (N_986,N_762,N_640);
or U987 (N_987,N_745,N_731);
and U988 (N_988,N_697,N_760);
or U989 (N_989,N_765,N_662);
nand U990 (N_990,N_654,N_767);
nand U991 (N_991,N_614,N_688);
and U992 (N_992,N_716,N_638);
nor U993 (N_993,N_652,N_606);
nand U994 (N_994,N_730,N_742);
and U995 (N_995,N_747,N_674);
nor U996 (N_996,N_745,N_797);
nor U997 (N_997,N_789,N_741);
or U998 (N_998,N_699,N_615);
nand U999 (N_999,N_755,N_715);
and U1000 (N_1000,N_896,N_839);
or U1001 (N_1001,N_851,N_833);
nor U1002 (N_1002,N_980,N_892);
and U1003 (N_1003,N_921,N_803);
nor U1004 (N_1004,N_885,N_850);
or U1005 (N_1005,N_966,N_869);
nand U1006 (N_1006,N_877,N_832);
nand U1007 (N_1007,N_829,N_905);
nand U1008 (N_1008,N_801,N_842);
and U1009 (N_1009,N_820,N_827);
and U1010 (N_1010,N_819,N_918);
nor U1011 (N_1011,N_947,N_909);
nor U1012 (N_1012,N_985,N_828);
or U1013 (N_1013,N_906,N_917);
and U1014 (N_1014,N_907,N_922);
and U1015 (N_1015,N_945,N_899);
nor U1016 (N_1016,N_826,N_807);
nor U1017 (N_1017,N_900,N_957);
nor U1018 (N_1018,N_843,N_935);
or U1019 (N_1019,N_903,N_952);
or U1020 (N_1020,N_870,N_949);
and U1021 (N_1021,N_914,N_848);
or U1022 (N_1022,N_808,N_859);
nand U1023 (N_1023,N_997,N_974);
nor U1024 (N_1024,N_920,N_973);
xor U1025 (N_1025,N_816,N_874);
and U1026 (N_1026,N_844,N_897);
nand U1027 (N_1027,N_982,N_963);
and U1028 (N_1028,N_994,N_845);
or U1029 (N_1029,N_979,N_858);
or U1030 (N_1030,N_872,N_888);
or U1031 (N_1031,N_999,N_913);
and U1032 (N_1032,N_958,N_898);
nand U1033 (N_1033,N_887,N_800);
nand U1034 (N_1034,N_881,N_821);
nand U1035 (N_1035,N_970,N_884);
nor U1036 (N_1036,N_878,N_838);
and U1037 (N_1037,N_811,N_910);
or U1038 (N_1038,N_946,N_965);
and U1039 (N_1039,N_993,N_865);
or U1040 (N_1040,N_901,N_849);
nor U1041 (N_1041,N_831,N_818);
nand U1042 (N_1042,N_893,N_825);
or U1043 (N_1043,N_936,N_853);
or U1044 (N_1044,N_996,N_912);
nor U1045 (N_1045,N_840,N_925);
and U1046 (N_1046,N_988,N_856);
and U1047 (N_1047,N_986,N_991);
nor U1048 (N_1048,N_951,N_989);
or U1049 (N_1049,N_880,N_961);
nor U1050 (N_1050,N_817,N_889);
and U1051 (N_1051,N_871,N_868);
and U1052 (N_1052,N_972,N_924);
nor U1053 (N_1053,N_954,N_864);
nor U1054 (N_1054,N_928,N_948);
nor U1055 (N_1055,N_908,N_911);
and U1056 (N_1056,N_943,N_861);
nor U1057 (N_1057,N_919,N_866);
or U1058 (N_1058,N_975,N_983);
nor U1059 (N_1059,N_882,N_971);
or U1060 (N_1060,N_823,N_802);
xnor U1061 (N_1061,N_830,N_834);
and U1062 (N_1062,N_886,N_860);
nand U1063 (N_1063,N_959,N_812);
and U1064 (N_1064,N_883,N_969);
and U1065 (N_1065,N_894,N_956);
nand U1066 (N_1066,N_814,N_944);
nand U1067 (N_1067,N_976,N_934);
or U1068 (N_1068,N_810,N_852);
and U1069 (N_1069,N_806,N_932);
nand U1070 (N_1070,N_929,N_837);
and U1071 (N_1071,N_841,N_937);
and U1072 (N_1072,N_895,N_930);
or U1073 (N_1073,N_953,N_835);
nor U1074 (N_1074,N_977,N_863);
nand U1075 (N_1075,N_809,N_968);
nor U1076 (N_1076,N_987,N_824);
or U1077 (N_1077,N_992,N_822);
nand U1078 (N_1078,N_978,N_984);
and U1079 (N_1079,N_967,N_990);
nand U1080 (N_1080,N_891,N_938);
nand U1081 (N_1081,N_855,N_942);
nand U1082 (N_1082,N_950,N_939);
nor U1083 (N_1083,N_867,N_836);
nor U1084 (N_1084,N_854,N_879);
or U1085 (N_1085,N_904,N_805);
nor U1086 (N_1086,N_923,N_960);
nor U1087 (N_1087,N_875,N_995);
nand U1088 (N_1088,N_862,N_813);
nand U1089 (N_1089,N_915,N_998);
nor U1090 (N_1090,N_927,N_916);
or U1091 (N_1091,N_964,N_890);
or U1092 (N_1092,N_902,N_962);
or U1093 (N_1093,N_876,N_857);
or U1094 (N_1094,N_931,N_815);
or U1095 (N_1095,N_981,N_846);
nor U1096 (N_1096,N_926,N_933);
and U1097 (N_1097,N_955,N_847);
or U1098 (N_1098,N_873,N_941);
xor U1099 (N_1099,N_804,N_940);
and U1100 (N_1100,N_875,N_902);
and U1101 (N_1101,N_985,N_846);
nor U1102 (N_1102,N_955,N_815);
and U1103 (N_1103,N_953,N_942);
and U1104 (N_1104,N_982,N_858);
and U1105 (N_1105,N_824,N_940);
or U1106 (N_1106,N_826,N_980);
and U1107 (N_1107,N_824,N_875);
and U1108 (N_1108,N_855,N_915);
nand U1109 (N_1109,N_899,N_838);
and U1110 (N_1110,N_862,N_887);
and U1111 (N_1111,N_820,N_873);
or U1112 (N_1112,N_812,N_924);
nand U1113 (N_1113,N_883,N_805);
and U1114 (N_1114,N_989,N_971);
nor U1115 (N_1115,N_926,N_994);
and U1116 (N_1116,N_826,N_854);
or U1117 (N_1117,N_828,N_940);
and U1118 (N_1118,N_892,N_887);
or U1119 (N_1119,N_899,N_982);
nand U1120 (N_1120,N_998,N_958);
and U1121 (N_1121,N_827,N_973);
nor U1122 (N_1122,N_845,N_870);
nor U1123 (N_1123,N_996,N_980);
nor U1124 (N_1124,N_925,N_806);
and U1125 (N_1125,N_898,N_999);
or U1126 (N_1126,N_996,N_849);
and U1127 (N_1127,N_976,N_808);
nand U1128 (N_1128,N_944,N_803);
or U1129 (N_1129,N_913,N_992);
nand U1130 (N_1130,N_895,N_945);
or U1131 (N_1131,N_887,N_951);
nor U1132 (N_1132,N_822,N_964);
nand U1133 (N_1133,N_886,N_864);
or U1134 (N_1134,N_956,N_927);
and U1135 (N_1135,N_813,N_887);
or U1136 (N_1136,N_875,N_913);
nor U1137 (N_1137,N_816,N_864);
or U1138 (N_1138,N_996,N_979);
nor U1139 (N_1139,N_887,N_838);
and U1140 (N_1140,N_980,N_952);
nand U1141 (N_1141,N_888,N_984);
nor U1142 (N_1142,N_881,N_917);
and U1143 (N_1143,N_826,N_949);
or U1144 (N_1144,N_801,N_993);
nor U1145 (N_1145,N_882,N_884);
and U1146 (N_1146,N_844,N_987);
and U1147 (N_1147,N_928,N_855);
nor U1148 (N_1148,N_985,N_817);
nor U1149 (N_1149,N_940,N_838);
and U1150 (N_1150,N_865,N_935);
nor U1151 (N_1151,N_834,N_945);
or U1152 (N_1152,N_836,N_905);
nand U1153 (N_1153,N_834,N_884);
and U1154 (N_1154,N_931,N_823);
or U1155 (N_1155,N_930,N_877);
xor U1156 (N_1156,N_877,N_956);
nor U1157 (N_1157,N_807,N_887);
or U1158 (N_1158,N_986,N_861);
nor U1159 (N_1159,N_845,N_803);
and U1160 (N_1160,N_959,N_993);
nor U1161 (N_1161,N_808,N_843);
nor U1162 (N_1162,N_803,N_922);
and U1163 (N_1163,N_958,N_810);
or U1164 (N_1164,N_919,N_931);
or U1165 (N_1165,N_975,N_856);
or U1166 (N_1166,N_943,N_823);
or U1167 (N_1167,N_829,N_938);
nor U1168 (N_1168,N_982,N_971);
nor U1169 (N_1169,N_836,N_889);
nor U1170 (N_1170,N_819,N_812);
nand U1171 (N_1171,N_875,N_864);
nor U1172 (N_1172,N_883,N_877);
nand U1173 (N_1173,N_955,N_836);
and U1174 (N_1174,N_875,N_801);
nand U1175 (N_1175,N_823,N_970);
and U1176 (N_1176,N_932,N_813);
nand U1177 (N_1177,N_966,N_890);
nand U1178 (N_1178,N_804,N_958);
nand U1179 (N_1179,N_885,N_803);
nor U1180 (N_1180,N_912,N_941);
and U1181 (N_1181,N_801,N_981);
or U1182 (N_1182,N_851,N_870);
nand U1183 (N_1183,N_844,N_817);
nor U1184 (N_1184,N_947,N_899);
nand U1185 (N_1185,N_992,N_989);
nor U1186 (N_1186,N_804,N_963);
or U1187 (N_1187,N_938,N_973);
and U1188 (N_1188,N_856,N_924);
or U1189 (N_1189,N_947,N_935);
xor U1190 (N_1190,N_911,N_997);
nand U1191 (N_1191,N_886,N_960);
xor U1192 (N_1192,N_822,N_803);
nand U1193 (N_1193,N_883,N_867);
or U1194 (N_1194,N_928,N_856);
nor U1195 (N_1195,N_982,N_890);
or U1196 (N_1196,N_980,N_989);
or U1197 (N_1197,N_947,N_998);
or U1198 (N_1198,N_944,N_890);
nand U1199 (N_1199,N_922,N_860);
nand U1200 (N_1200,N_1024,N_1059);
nor U1201 (N_1201,N_1145,N_1178);
nand U1202 (N_1202,N_1193,N_1101);
nand U1203 (N_1203,N_1163,N_1017);
nor U1204 (N_1204,N_1199,N_1097);
nor U1205 (N_1205,N_1098,N_1061);
nand U1206 (N_1206,N_1026,N_1170);
or U1207 (N_1207,N_1140,N_1057);
nand U1208 (N_1208,N_1111,N_1006);
nor U1209 (N_1209,N_1056,N_1181);
nand U1210 (N_1210,N_1001,N_1087);
nor U1211 (N_1211,N_1106,N_1169);
nor U1212 (N_1212,N_1162,N_1195);
or U1213 (N_1213,N_1037,N_1109);
nor U1214 (N_1214,N_1002,N_1019);
nand U1215 (N_1215,N_1187,N_1089);
and U1216 (N_1216,N_1058,N_1069);
nand U1217 (N_1217,N_1023,N_1034);
nor U1218 (N_1218,N_1031,N_1009);
nand U1219 (N_1219,N_1192,N_1117);
or U1220 (N_1220,N_1115,N_1104);
nor U1221 (N_1221,N_1194,N_1110);
xnor U1222 (N_1222,N_1112,N_1004);
xor U1223 (N_1223,N_1011,N_1039);
nor U1224 (N_1224,N_1100,N_1042);
or U1225 (N_1225,N_1167,N_1148);
or U1226 (N_1226,N_1022,N_1118);
nand U1227 (N_1227,N_1040,N_1007);
and U1228 (N_1228,N_1177,N_1091);
and U1229 (N_1229,N_1119,N_1171);
nand U1230 (N_1230,N_1094,N_1173);
or U1231 (N_1231,N_1139,N_1124);
and U1232 (N_1232,N_1071,N_1136);
nor U1233 (N_1233,N_1076,N_1044);
nor U1234 (N_1234,N_1068,N_1079);
and U1235 (N_1235,N_1014,N_1120);
or U1236 (N_1236,N_1186,N_1072);
nor U1237 (N_1237,N_1131,N_1154);
or U1238 (N_1238,N_1147,N_1066);
or U1239 (N_1239,N_1015,N_1176);
and U1240 (N_1240,N_1159,N_1165);
nand U1241 (N_1241,N_1065,N_1129);
or U1242 (N_1242,N_1102,N_1095);
nor U1243 (N_1243,N_1133,N_1125);
and U1244 (N_1244,N_1126,N_1161);
or U1245 (N_1245,N_1123,N_1051);
nand U1246 (N_1246,N_1018,N_1128);
and U1247 (N_1247,N_1141,N_1143);
or U1248 (N_1248,N_1137,N_1127);
or U1249 (N_1249,N_1081,N_1180);
nor U1250 (N_1250,N_1030,N_1174);
or U1251 (N_1251,N_1188,N_1064);
xor U1252 (N_1252,N_1077,N_1084);
and U1253 (N_1253,N_1116,N_1121);
and U1254 (N_1254,N_1114,N_1080);
and U1255 (N_1255,N_1074,N_1168);
and U1256 (N_1256,N_1045,N_1062);
nand U1257 (N_1257,N_1043,N_1103);
nand U1258 (N_1258,N_1164,N_1038);
or U1259 (N_1259,N_1189,N_1153);
and U1260 (N_1260,N_1055,N_1085);
nand U1261 (N_1261,N_1012,N_1016);
or U1262 (N_1262,N_1025,N_1198);
and U1263 (N_1263,N_1050,N_1185);
nand U1264 (N_1264,N_1096,N_1158);
or U1265 (N_1265,N_1035,N_1105);
and U1266 (N_1266,N_1191,N_1020);
or U1267 (N_1267,N_1130,N_1052);
or U1268 (N_1268,N_1108,N_1082);
or U1269 (N_1269,N_1144,N_1155);
nor U1270 (N_1270,N_1197,N_1060);
and U1271 (N_1271,N_1086,N_1010);
nand U1272 (N_1272,N_1138,N_1183);
nor U1273 (N_1273,N_1142,N_1041);
nand U1274 (N_1274,N_1113,N_1036);
nor U1275 (N_1275,N_1150,N_1054);
xnor U1276 (N_1276,N_1107,N_1156);
xnor U1277 (N_1277,N_1160,N_1053);
or U1278 (N_1278,N_1047,N_1048);
and U1279 (N_1279,N_1078,N_1157);
nand U1280 (N_1280,N_1008,N_1088);
nor U1281 (N_1281,N_1092,N_1146);
or U1282 (N_1282,N_1152,N_1073);
nor U1283 (N_1283,N_1028,N_1099);
nand U1284 (N_1284,N_1070,N_1003);
or U1285 (N_1285,N_1172,N_1166);
nand U1286 (N_1286,N_1067,N_1135);
nand U1287 (N_1287,N_1063,N_1083);
and U1288 (N_1288,N_1151,N_1190);
and U1289 (N_1289,N_1175,N_1184);
nand U1290 (N_1290,N_1029,N_1134);
and U1291 (N_1291,N_1049,N_1075);
nor U1292 (N_1292,N_1033,N_1149);
nand U1293 (N_1293,N_1005,N_1132);
or U1294 (N_1294,N_1090,N_1013);
nand U1295 (N_1295,N_1179,N_1032);
and U1296 (N_1296,N_1027,N_1021);
or U1297 (N_1297,N_1046,N_1000);
nand U1298 (N_1298,N_1122,N_1093);
and U1299 (N_1299,N_1196,N_1182);
or U1300 (N_1300,N_1089,N_1002);
and U1301 (N_1301,N_1049,N_1069);
or U1302 (N_1302,N_1055,N_1100);
nor U1303 (N_1303,N_1155,N_1066);
nor U1304 (N_1304,N_1192,N_1077);
or U1305 (N_1305,N_1199,N_1111);
nand U1306 (N_1306,N_1010,N_1113);
nand U1307 (N_1307,N_1115,N_1161);
xor U1308 (N_1308,N_1192,N_1042);
and U1309 (N_1309,N_1049,N_1151);
or U1310 (N_1310,N_1099,N_1073);
or U1311 (N_1311,N_1054,N_1100);
nand U1312 (N_1312,N_1182,N_1184);
nand U1313 (N_1313,N_1006,N_1009);
nand U1314 (N_1314,N_1183,N_1040);
nand U1315 (N_1315,N_1004,N_1136);
xnor U1316 (N_1316,N_1158,N_1116);
or U1317 (N_1317,N_1053,N_1073);
and U1318 (N_1318,N_1099,N_1132);
nand U1319 (N_1319,N_1057,N_1115);
and U1320 (N_1320,N_1129,N_1067);
nand U1321 (N_1321,N_1174,N_1199);
or U1322 (N_1322,N_1052,N_1034);
nor U1323 (N_1323,N_1151,N_1034);
or U1324 (N_1324,N_1145,N_1095);
nand U1325 (N_1325,N_1147,N_1133);
or U1326 (N_1326,N_1043,N_1059);
or U1327 (N_1327,N_1088,N_1011);
nand U1328 (N_1328,N_1083,N_1134);
nor U1329 (N_1329,N_1113,N_1157);
nand U1330 (N_1330,N_1141,N_1036);
and U1331 (N_1331,N_1012,N_1183);
or U1332 (N_1332,N_1098,N_1185);
or U1333 (N_1333,N_1144,N_1040);
nor U1334 (N_1334,N_1152,N_1009);
nor U1335 (N_1335,N_1097,N_1060);
and U1336 (N_1336,N_1174,N_1183);
nor U1337 (N_1337,N_1105,N_1109);
or U1338 (N_1338,N_1186,N_1031);
and U1339 (N_1339,N_1150,N_1106);
nand U1340 (N_1340,N_1037,N_1132);
or U1341 (N_1341,N_1186,N_1181);
and U1342 (N_1342,N_1027,N_1046);
or U1343 (N_1343,N_1057,N_1013);
nor U1344 (N_1344,N_1064,N_1098);
and U1345 (N_1345,N_1176,N_1084);
or U1346 (N_1346,N_1199,N_1017);
or U1347 (N_1347,N_1185,N_1116);
xor U1348 (N_1348,N_1062,N_1122);
and U1349 (N_1349,N_1009,N_1150);
nor U1350 (N_1350,N_1175,N_1079);
nor U1351 (N_1351,N_1149,N_1054);
or U1352 (N_1352,N_1031,N_1064);
nand U1353 (N_1353,N_1079,N_1041);
or U1354 (N_1354,N_1109,N_1187);
or U1355 (N_1355,N_1191,N_1050);
or U1356 (N_1356,N_1000,N_1163);
and U1357 (N_1357,N_1190,N_1074);
nand U1358 (N_1358,N_1049,N_1121);
and U1359 (N_1359,N_1138,N_1002);
or U1360 (N_1360,N_1112,N_1187);
nand U1361 (N_1361,N_1010,N_1180);
or U1362 (N_1362,N_1108,N_1035);
and U1363 (N_1363,N_1138,N_1157);
nor U1364 (N_1364,N_1126,N_1157);
or U1365 (N_1365,N_1122,N_1115);
and U1366 (N_1366,N_1192,N_1030);
or U1367 (N_1367,N_1184,N_1179);
nand U1368 (N_1368,N_1184,N_1017);
nor U1369 (N_1369,N_1051,N_1049);
and U1370 (N_1370,N_1126,N_1140);
and U1371 (N_1371,N_1046,N_1155);
nor U1372 (N_1372,N_1065,N_1022);
nand U1373 (N_1373,N_1127,N_1059);
nor U1374 (N_1374,N_1138,N_1150);
nor U1375 (N_1375,N_1050,N_1170);
nand U1376 (N_1376,N_1029,N_1159);
nor U1377 (N_1377,N_1147,N_1113);
and U1378 (N_1378,N_1057,N_1176);
or U1379 (N_1379,N_1151,N_1057);
nand U1380 (N_1380,N_1090,N_1117);
nand U1381 (N_1381,N_1095,N_1044);
nand U1382 (N_1382,N_1097,N_1162);
or U1383 (N_1383,N_1140,N_1186);
or U1384 (N_1384,N_1124,N_1050);
or U1385 (N_1385,N_1138,N_1132);
and U1386 (N_1386,N_1023,N_1170);
or U1387 (N_1387,N_1139,N_1083);
nor U1388 (N_1388,N_1021,N_1142);
nor U1389 (N_1389,N_1013,N_1167);
and U1390 (N_1390,N_1192,N_1084);
nor U1391 (N_1391,N_1146,N_1109);
nand U1392 (N_1392,N_1094,N_1128);
nand U1393 (N_1393,N_1188,N_1069);
and U1394 (N_1394,N_1007,N_1109);
and U1395 (N_1395,N_1171,N_1141);
nand U1396 (N_1396,N_1035,N_1057);
or U1397 (N_1397,N_1178,N_1073);
nand U1398 (N_1398,N_1003,N_1047);
nor U1399 (N_1399,N_1076,N_1176);
nor U1400 (N_1400,N_1209,N_1391);
or U1401 (N_1401,N_1332,N_1250);
xor U1402 (N_1402,N_1259,N_1257);
nor U1403 (N_1403,N_1269,N_1333);
and U1404 (N_1404,N_1238,N_1321);
nor U1405 (N_1405,N_1346,N_1339);
nand U1406 (N_1406,N_1360,N_1350);
nor U1407 (N_1407,N_1288,N_1312);
nor U1408 (N_1408,N_1331,N_1394);
and U1409 (N_1409,N_1347,N_1241);
or U1410 (N_1410,N_1377,N_1320);
nand U1411 (N_1411,N_1336,N_1334);
nor U1412 (N_1412,N_1319,N_1385);
and U1413 (N_1413,N_1303,N_1289);
nor U1414 (N_1414,N_1351,N_1236);
xor U1415 (N_1415,N_1311,N_1270);
or U1416 (N_1416,N_1239,N_1248);
or U1417 (N_1417,N_1228,N_1285);
and U1418 (N_1418,N_1326,N_1307);
nand U1419 (N_1419,N_1398,N_1314);
nand U1420 (N_1420,N_1220,N_1363);
or U1421 (N_1421,N_1308,N_1274);
nor U1422 (N_1422,N_1355,N_1358);
nor U1423 (N_1423,N_1234,N_1330);
and U1424 (N_1424,N_1343,N_1263);
nand U1425 (N_1425,N_1252,N_1337);
or U1426 (N_1426,N_1295,N_1335);
or U1427 (N_1427,N_1362,N_1258);
nor U1428 (N_1428,N_1246,N_1310);
and U1429 (N_1429,N_1202,N_1229);
and U1430 (N_1430,N_1207,N_1386);
and U1431 (N_1431,N_1268,N_1367);
or U1432 (N_1432,N_1203,N_1325);
and U1433 (N_1433,N_1397,N_1287);
nand U1434 (N_1434,N_1206,N_1226);
nor U1435 (N_1435,N_1211,N_1341);
and U1436 (N_1436,N_1297,N_1204);
and U1437 (N_1437,N_1224,N_1352);
or U1438 (N_1438,N_1291,N_1221);
or U1439 (N_1439,N_1237,N_1345);
xnor U1440 (N_1440,N_1282,N_1348);
nand U1441 (N_1441,N_1253,N_1217);
or U1442 (N_1442,N_1324,N_1271);
nand U1443 (N_1443,N_1309,N_1370);
nand U1444 (N_1444,N_1261,N_1260);
nand U1445 (N_1445,N_1390,N_1281);
nor U1446 (N_1446,N_1200,N_1293);
or U1447 (N_1447,N_1212,N_1275);
nor U1448 (N_1448,N_1276,N_1243);
and U1449 (N_1449,N_1374,N_1232);
nor U1450 (N_1450,N_1249,N_1368);
and U1451 (N_1451,N_1233,N_1284);
or U1452 (N_1452,N_1219,N_1280);
and U1453 (N_1453,N_1364,N_1356);
and U1454 (N_1454,N_1389,N_1283);
and U1455 (N_1455,N_1264,N_1372);
or U1456 (N_1456,N_1382,N_1205);
and U1457 (N_1457,N_1361,N_1301);
nor U1458 (N_1458,N_1277,N_1244);
nand U1459 (N_1459,N_1384,N_1208);
and U1460 (N_1460,N_1279,N_1323);
or U1461 (N_1461,N_1298,N_1255);
or U1462 (N_1462,N_1292,N_1380);
nor U1463 (N_1463,N_1265,N_1227);
and U1464 (N_1464,N_1216,N_1305);
nor U1465 (N_1465,N_1344,N_1396);
nor U1466 (N_1466,N_1267,N_1290);
or U1467 (N_1467,N_1381,N_1375);
nor U1468 (N_1468,N_1315,N_1225);
nor U1469 (N_1469,N_1373,N_1299);
nand U1470 (N_1470,N_1222,N_1218);
and U1471 (N_1471,N_1296,N_1354);
and U1472 (N_1472,N_1349,N_1230);
and U1473 (N_1473,N_1338,N_1240);
nand U1474 (N_1474,N_1340,N_1266);
and U1475 (N_1475,N_1213,N_1328);
nand U1476 (N_1476,N_1378,N_1342);
and U1477 (N_1477,N_1322,N_1392);
and U1478 (N_1478,N_1300,N_1304);
and U1479 (N_1479,N_1387,N_1327);
or U1480 (N_1480,N_1379,N_1254);
and U1481 (N_1481,N_1294,N_1278);
nand U1482 (N_1482,N_1245,N_1214);
nand U1483 (N_1483,N_1247,N_1273);
or U1484 (N_1484,N_1357,N_1383);
nand U1485 (N_1485,N_1366,N_1262);
or U1486 (N_1486,N_1388,N_1306);
and U1487 (N_1487,N_1365,N_1376);
nor U1488 (N_1488,N_1272,N_1223);
xor U1489 (N_1489,N_1359,N_1329);
nor U1490 (N_1490,N_1369,N_1316);
and U1491 (N_1491,N_1231,N_1242);
xnor U1492 (N_1492,N_1313,N_1215);
or U1493 (N_1493,N_1210,N_1256);
nand U1494 (N_1494,N_1395,N_1393);
and U1495 (N_1495,N_1235,N_1201);
nor U1496 (N_1496,N_1317,N_1399);
nand U1497 (N_1497,N_1318,N_1251);
nor U1498 (N_1498,N_1371,N_1302);
and U1499 (N_1499,N_1286,N_1353);
and U1500 (N_1500,N_1213,N_1342);
nor U1501 (N_1501,N_1270,N_1264);
nor U1502 (N_1502,N_1382,N_1211);
nand U1503 (N_1503,N_1359,N_1341);
and U1504 (N_1504,N_1319,N_1219);
nor U1505 (N_1505,N_1393,N_1309);
and U1506 (N_1506,N_1246,N_1279);
or U1507 (N_1507,N_1200,N_1211);
and U1508 (N_1508,N_1310,N_1242);
or U1509 (N_1509,N_1256,N_1374);
and U1510 (N_1510,N_1390,N_1312);
nand U1511 (N_1511,N_1351,N_1332);
and U1512 (N_1512,N_1252,N_1219);
and U1513 (N_1513,N_1358,N_1303);
nand U1514 (N_1514,N_1275,N_1325);
nand U1515 (N_1515,N_1205,N_1221);
and U1516 (N_1516,N_1271,N_1255);
nand U1517 (N_1517,N_1215,N_1226);
nand U1518 (N_1518,N_1285,N_1234);
and U1519 (N_1519,N_1243,N_1257);
nor U1520 (N_1520,N_1347,N_1271);
nand U1521 (N_1521,N_1369,N_1229);
nand U1522 (N_1522,N_1330,N_1399);
nor U1523 (N_1523,N_1383,N_1367);
and U1524 (N_1524,N_1306,N_1206);
nor U1525 (N_1525,N_1276,N_1360);
nor U1526 (N_1526,N_1335,N_1226);
and U1527 (N_1527,N_1331,N_1263);
or U1528 (N_1528,N_1307,N_1239);
nor U1529 (N_1529,N_1399,N_1207);
xor U1530 (N_1530,N_1372,N_1364);
xnor U1531 (N_1531,N_1368,N_1392);
and U1532 (N_1532,N_1388,N_1399);
nand U1533 (N_1533,N_1254,N_1266);
and U1534 (N_1534,N_1290,N_1398);
or U1535 (N_1535,N_1221,N_1200);
or U1536 (N_1536,N_1241,N_1249);
nor U1537 (N_1537,N_1286,N_1391);
and U1538 (N_1538,N_1294,N_1212);
nor U1539 (N_1539,N_1308,N_1369);
and U1540 (N_1540,N_1224,N_1334);
nand U1541 (N_1541,N_1236,N_1273);
and U1542 (N_1542,N_1377,N_1329);
nor U1543 (N_1543,N_1315,N_1309);
or U1544 (N_1544,N_1333,N_1314);
nor U1545 (N_1545,N_1392,N_1366);
and U1546 (N_1546,N_1225,N_1386);
and U1547 (N_1547,N_1397,N_1304);
and U1548 (N_1548,N_1214,N_1359);
nor U1549 (N_1549,N_1266,N_1231);
nor U1550 (N_1550,N_1262,N_1267);
nor U1551 (N_1551,N_1295,N_1357);
nor U1552 (N_1552,N_1214,N_1288);
nor U1553 (N_1553,N_1214,N_1263);
nand U1554 (N_1554,N_1316,N_1211);
and U1555 (N_1555,N_1373,N_1235);
nand U1556 (N_1556,N_1353,N_1214);
nor U1557 (N_1557,N_1310,N_1306);
and U1558 (N_1558,N_1228,N_1321);
and U1559 (N_1559,N_1339,N_1371);
nand U1560 (N_1560,N_1343,N_1373);
or U1561 (N_1561,N_1389,N_1219);
and U1562 (N_1562,N_1295,N_1287);
and U1563 (N_1563,N_1251,N_1374);
and U1564 (N_1564,N_1230,N_1267);
nor U1565 (N_1565,N_1393,N_1293);
or U1566 (N_1566,N_1352,N_1246);
and U1567 (N_1567,N_1262,N_1347);
and U1568 (N_1568,N_1209,N_1214);
and U1569 (N_1569,N_1270,N_1256);
nor U1570 (N_1570,N_1241,N_1233);
or U1571 (N_1571,N_1204,N_1230);
nor U1572 (N_1572,N_1204,N_1398);
and U1573 (N_1573,N_1235,N_1236);
nor U1574 (N_1574,N_1201,N_1215);
or U1575 (N_1575,N_1220,N_1335);
nand U1576 (N_1576,N_1391,N_1359);
nand U1577 (N_1577,N_1235,N_1338);
nand U1578 (N_1578,N_1368,N_1241);
and U1579 (N_1579,N_1213,N_1200);
nor U1580 (N_1580,N_1352,N_1315);
nand U1581 (N_1581,N_1331,N_1287);
nand U1582 (N_1582,N_1228,N_1227);
and U1583 (N_1583,N_1202,N_1225);
nand U1584 (N_1584,N_1388,N_1390);
nor U1585 (N_1585,N_1211,N_1278);
or U1586 (N_1586,N_1244,N_1232);
nand U1587 (N_1587,N_1265,N_1382);
or U1588 (N_1588,N_1383,N_1229);
or U1589 (N_1589,N_1265,N_1320);
and U1590 (N_1590,N_1273,N_1336);
and U1591 (N_1591,N_1289,N_1376);
or U1592 (N_1592,N_1365,N_1328);
or U1593 (N_1593,N_1317,N_1284);
nand U1594 (N_1594,N_1285,N_1316);
nor U1595 (N_1595,N_1210,N_1399);
nor U1596 (N_1596,N_1222,N_1211);
nor U1597 (N_1597,N_1246,N_1230);
nand U1598 (N_1598,N_1386,N_1371);
or U1599 (N_1599,N_1261,N_1355);
nor U1600 (N_1600,N_1412,N_1557);
nor U1601 (N_1601,N_1443,N_1471);
and U1602 (N_1602,N_1463,N_1411);
and U1603 (N_1603,N_1490,N_1590);
and U1604 (N_1604,N_1470,N_1568);
or U1605 (N_1605,N_1572,N_1461);
or U1606 (N_1606,N_1524,N_1452);
and U1607 (N_1607,N_1466,N_1556);
nor U1608 (N_1608,N_1507,N_1529);
and U1609 (N_1609,N_1563,N_1585);
and U1610 (N_1610,N_1464,N_1543);
or U1611 (N_1611,N_1539,N_1431);
nand U1612 (N_1612,N_1521,N_1582);
or U1613 (N_1613,N_1561,N_1552);
xnor U1614 (N_1614,N_1406,N_1574);
or U1615 (N_1615,N_1535,N_1555);
and U1616 (N_1616,N_1503,N_1525);
xnor U1617 (N_1617,N_1597,N_1550);
or U1618 (N_1618,N_1577,N_1413);
or U1619 (N_1619,N_1509,N_1460);
nor U1620 (N_1620,N_1586,N_1445);
nor U1621 (N_1621,N_1514,N_1484);
and U1622 (N_1622,N_1435,N_1593);
and U1623 (N_1623,N_1537,N_1419);
nor U1624 (N_1624,N_1576,N_1579);
nand U1625 (N_1625,N_1491,N_1438);
and U1626 (N_1626,N_1459,N_1486);
nor U1627 (N_1627,N_1564,N_1544);
or U1628 (N_1628,N_1533,N_1434);
nand U1629 (N_1629,N_1497,N_1496);
and U1630 (N_1630,N_1441,N_1513);
nor U1631 (N_1631,N_1522,N_1498);
and U1632 (N_1632,N_1462,N_1575);
nand U1633 (N_1633,N_1587,N_1440);
nor U1634 (N_1634,N_1457,N_1591);
and U1635 (N_1635,N_1429,N_1505);
nor U1636 (N_1636,N_1430,N_1517);
nor U1637 (N_1637,N_1558,N_1494);
nor U1638 (N_1638,N_1421,N_1488);
nand U1639 (N_1639,N_1404,N_1588);
and U1640 (N_1640,N_1454,N_1504);
nor U1641 (N_1641,N_1405,N_1477);
or U1642 (N_1642,N_1481,N_1547);
or U1643 (N_1643,N_1500,N_1594);
nor U1644 (N_1644,N_1569,N_1415);
or U1645 (N_1645,N_1472,N_1570);
and U1646 (N_1646,N_1483,N_1553);
nand U1647 (N_1647,N_1403,N_1518);
and U1648 (N_1648,N_1548,N_1566);
and U1649 (N_1649,N_1455,N_1424);
nand U1650 (N_1650,N_1581,N_1428);
nand U1651 (N_1651,N_1541,N_1512);
nand U1652 (N_1652,N_1478,N_1465);
nand U1653 (N_1653,N_1499,N_1467);
nand U1654 (N_1654,N_1515,N_1567);
and U1655 (N_1655,N_1565,N_1407);
nand U1656 (N_1656,N_1436,N_1542);
and U1657 (N_1657,N_1458,N_1451);
or U1658 (N_1658,N_1469,N_1401);
nand U1659 (N_1659,N_1416,N_1502);
and U1660 (N_1660,N_1501,N_1426);
nand U1661 (N_1661,N_1508,N_1446);
or U1662 (N_1662,N_1584,N_1456);
or U1663 (N_1663,N_1479,N_1487);
nand U1664 (N_1664,N_1523,N_1449);
nand U1665 (N_1665,N_1526,N_1519);
and U1666 (N_1666,N_1489,N_1474);
and U1667 (N_1667,N_1527,N_1473);
and U1668 (N_1668,N_1598,N_1480);
nand U1669 (N_1669,N_1423,N_1589);
nor U1670 (N_1670,N_1540,N_1439);
nand U1671 (N_1671,N_1432,N_1444);
nand U1672 (N_1672,N_1595,N_1583);
nand U1673 (N_1673,N_1596,N_1536);
and U1674 (N_1674,N_1418,N_1549);
and U1675 (N_1675,N_1551,N_1571);
or U1676 (N_1676,N_1573,N_1468);
nor U1677 (N_1677,N_1442,N_1546);
and U1678 (N_1678,N_1433,N_1580);
nor U1679 (N_1679,N_1417,N_1495);
nor U1680 (N_1680,N_1414,N_1528);
or U1681 (N_1681,N_1400,N_1562);
nor U1682 (N_1682,N_1520,N_1599);
and U1683 (N_1683,N_1402,N_1560);
and U1684 (N_1684,N_1476,N_1485);
xnor U1685 (N_1685,N_1409,N_1506);
nor U1686 (N_1686,N_1592,N_1475);
and U1687 (N_1687,N_1554,N_1420);
or U1688 (N_1688,N_1532,N_1531);
and U1689 (N_1689,N_1530,N_1492);
nor U1690 (N_1690,N_1447,N_1511);
nor U1691 (N_1691,N_1410,N_1538);
nor U1692 (N_1692,N_1516,N_1534);
or U1693 (N_1693,N_1427,N_1448);
nor U1694 (N_1694,N_1437,N_1559);
nand U1695 (N_1695,N_1545,N_1422);
nand U1696 (N_1696,N_1453,N_1450);
and U1697 (N_1697,N_1493,N_1510);
or U1698 (N_1698,N_1425,N_1578);
nor U1699 (N_1699,N_1482,N_1408);
or U1700 (N_1700,N_1413,N_1464);
nor U1701 (N_1701,N_1432,N_1413);
nor U1702 (N_1702,N_1516,N_1425);
and U1703 (N_1703,N_1564,N_1451);
nand U1704 (N_1704,N_1405,N_1581);
and U1705 (N_1705,N_1465,N_1430);
and U1706 (N_1706,N_1487,N_1486);
and U1707 (N_1707,N_1480,N_1526);
and U1708 (N_1708,N_1496,N_1555);
nand U1709 (N_1709,N_1509,N_1523);
nor U1710 (N_1710,N_1500,N_1475);
and U1711 (N_1711,N_1437,N_1511);
nor U1712 (N_1712,N_1585,N_1570);
nor U1713 (N_1713,N_1527,N_1453);
nand U1714 (N_1714,N_1505,N_1592);
or U1715 (N_1715,N_1597,N_1450);
nand U1716 (N_1716,N_1503,N_1450);
or U1717 (N_1717,N_1501,N_1519);
xor U1718 (N_1718,N_1422,N_1582);
nand U1719 (N_1719,N_1586,N_1495);
nand U1720 (N_1720,N_1416,N_1514);
and U1721 (N_1721,N_1442,N_1521);
and U1722 (N_1722,N_1543,N_1454);
nand U1723 (N_1723,N_1532,N_1494);
nand U1724 (N_1724,N_1463,N_1571);
or U1725 (N_1725,N_1430,N_1521);
or U1726 (N_1726,N_1544,N_1469);
or U1727 (N_1727,N_1594,N_1468);
nand U1728 (N_1728,N_1494,N_1540);
nor U1729 (N_1729,N_1487,N_1499);
and U1730 (N_1730,N_1568,N_1491);
nand U1731 (N_1731,N_1526,N_1427);
and U1732 (N_1732,N_1551,N_1546);
nor U1733 (N_1733,N_1524,N_1434);
nand U1734 (N_1734,N_1464,N_1443);
nor U1735 (N_1735,N_1561,N_1546);
and U1736 (N_1736,N_1459,N_1564);
or U1737 (N_1737,N_1543,N_1559);
and U1738 (N_1738,N_1509,N_1543);
and U1739 (N_1739,N_1452,N_1434);
and U1740 (N_1740,N_1492,N_1436);
and U1741 (N_1741,N_1402,N_1420);
nand U1742 (N_1742,N_1448,N_1410);
or U1743 (N_1743,N_1510,N_1462);
or U1744 (N_1744,N_1547,N_1474);
and U1745 (N_1745,N_1527,N_1449);
or U1746 (N_1746,N_1498,N_1442);
and U1747 (N_1747,N_1440,N_1548);
or U1748 (N_1748,N_1574,N_1434);
xnor U1749 (N_1749,N_1539,N_1587);
nand U1750 (N_1750,N_1465,N_1467);
nand U1751 (N_1751,N_1505,N_1502);
and U1752 (N_1752,N_1425,N_1495);
or U1753 (N_1753,N_1419,N_1510);
or U1754 (N_1754,N_1535,N_1418);
nor U1755 (N_1755,N_1521,N_1555);
or U1756 (N_1756,N_1409,N_1578);
nand U1757 (N_1757,N_1446,N_1443);
nor U1758 (N_1758,N_1596,N_1567);
nor U1759 (N_1759,N_1474,N_1448);
and U1760 (N_1760,N_1549,N_1450);
or U1761 (N_1761,N_1471,N_1462);
and U1762 (N_1762,N_1544,N_1575);
and U1763 (N_1763,N_1403,N_1449);
nor U1764 (N_1764,N_1456,N_1596);
nor U1765 (N_1765,N_1457,N_1579);
or U1766 (N_1766,N_1438,N_1572);
or U1767 (N_1767,N_1540,N_1467);
nor U1768 (N_1768,N_1423,N_1552);
and U1769 (N_1769,N_1409,N_1463);
nor U1770 (N_1770,N_1416,N_1441);
nor U1771 (N_1771,N_1464,N_1454);
nand U1772 (N_1772,N_1542,N_1494);
nand U1773 (N_1773,N_1510,N_1475);
nand U1774 (N_1774,N_1562,N_1489);
nor U1775 (N_1775,N_1530,N_1575);
nor U1776 (N_1776,N_1443,N_1589);
nand U1777 (N_1777,N_1449,N_1567);
and U1778 (N_1778,N_1414,N_1423);
and U1779 (N_1779,N_1420,N_1581);
nand U1780 (N_1780,N_1455,N_1516);
nor U1781 (N_1781,N_1467,N_1579);
or U1782 (N_1782,N_1572,N_1403);
and U1783 (N_1783,N_1598,N_1470);
nand U1784 (N_1784,N_1547,N_1404);
or U1785 (N_1785,N_1454,N_1412);
nor U1786 (N_1786,N_1537,N_1563);
and U1787 (N_1787,N_1507,N_1408);
nor U1788 (N_1788,N_1488,N_1557);
nor U1789 (N_1789,N_1495,N_1553);
nor U1790 (N_1790,N_1504,N_1469);
or U1791 (N_1791,N_1494,N_1413);
or U1792 (N_1792,N_1497,N_1471);
or U1793 (N_1793,N_1476,N_1471);
or U1794 (N_1794,N_1486,N_1550);
and U1795 (N_1795,N_1444,N_1547);
nand U1796 (N_1796,N_1501,N_1464);
or U1797 (N_1797,N_1472,N_1592);
nor U1798 (N_1798,N_1452,N_1404);
xnor U1799 (N_1799,N_1469,N_1524);
and U1800 (N_1800,N_1718,N_1693);
or U1801 (N_1801,N_1666,N_1685);
nand U1802 (N_1802,N_1783,N_1774);
xor U1803 (N_1803,N_1660,N_1686);
nand U1804 (N_1804,N_1767,N_1733);
nand U1805 (N_1805,N_1664,N_1768);
nand U1806 (N_1806,N_1631,N_1638);
and U1807 (N_1807,N_1713,N_1659);
or U1808 (N_1808,N_1653,N_1798);
xor U1809 (N_1809,N_1748,N_1618);
nand U1810 (N_1810,N_1626,N_1765);
nand U1811 (N_1811,N_1648,N_1647);
nor U1812 (N_1812,N_1633,N_1764);
nand U1813 (N_1813,N_1641,N_1730);
and U1814 (N_1814,N_1739,N_1636);
nand U1815 (N_1815,N_1625,N_1716);
or U1816 (N_1816,N_1699,N_1753);
xor U1817 (N_1817,N_1789,N_1634);
or U1818 (N_1818,N_1793,N_1670);
nand U1819 (N_1819,N_1607,N_1704);
or U1820 (N_1820,N_1672,N_1757);
nand U1821 (N_1821,N_1743,N_1771);
nand U1822 (N_1822,N_1796,N_1649);
and U1823 (N_1823,N_1637,N_1787);
nand U1824 (N_1824,N_1781,N_1687);
nand U1825 (N_1825,N_1601,N_1688);
and U1826 (N_1826,N_1749,N_1705);
nand U1827 (N_1827,N_1663,N_1605);
or U1828 (N_1828,N_1620,N_1734);
or U1829 (N_1829,N_1691,N_1747);
nor U1830 (N_1830,N_1727,N_1770);
or U1831 (N_1831,N_1777,N_1766);
and U1832 (N_1832,N_1642,N_1639);
and U1833 (N_1833,N_1681,N_1797);
nor U1834 (N_1834,N_1720,N_1617);
and U1835 (N_1835,N_1711,N_1600);
and U1836 (N_1836,N_1623,N_1611);
and U1837 (N_1837,N_1752,N_1763);
nor U1838 (N_1838,N_1657,N_1608);
and U1839 (N_1839,N_1782,N_1635);
or U1840 (N_1840,N_1724,N_1609);
or U1841 (N_1841,N_1744,N_1755);
nand U1842 (N_1842,N_1694,N_1695);
nand U1843 (N_1843,N_1671,N_1684);
or U1844 (N_1844,N_1732,N_1702);
nand U1845 (N_1845,N_1624,N_1708);
nand U1846 (N_1846,N_1750,N_1761);
and U1847 (N_1847,N_1779,N_1622);
or U1848 (N_1848,N_1717,N_1745);
and U1849 (N_1849,N_1788,N_1772);
and U1850 (N_1850,N_1604,N_1795);
and U1851 (N_1851,N_1714,N_1709);
nor U1852 (N_1852,N_1728,N_1627);
and U1853 (N_1853,N_1615,N_1619);
nand U1854 (N_1854,N_1701,N_1721);
or U1855 (N_1855,N_1629,N_1773);
nand U1856 (N_1856,N_1786,N_1697);
nand U1857 (N_1857,N_1736,N_1703);
nor U1858 (N_1858,N_1654,N_1651);
and U1859 (N_1859,N_1644,N_1692);
nor U1860 (N_1860,N_1689,N_1630);
nor U1861 (N_1861,N_1759,N_1612);
nand U1862 (N_1862,N_1726,N_1769);
or U1863 (N_1863,N_1658,N_1632);
nor U1864 (N_1864,N_1791,N_1621);
nand U1865 (N_1865,N_1758,N_1616);
nand U1866 (N_1866,N_1628,N_1712);
nand U1867 (N_1867,N_1794,N_1683);
or U1868 (N_1868,N_1784,N_1700);
or U1869 (N_1869,N_1762,N_1662);
or U1870 (N_1870,N_1719,N_1735);
nor U1871 (N_1871,N_1690,N_1667);
nor U1872 (N_1872,N_1722,N_1706);
or U1873 (N_1873,N_1661,N_1751);
nand U1874 (N_1874,N_1656,N_1738);
nand U1875 (N_1875,N_1646,N_1679);
nand U1876 (N_1876,N_1746,N_1799);
nand U1877 (N_1877,N_1776,N_1678);
nand U1878 (N_1878,N_1673,N_1731);
nor U1879 (N_1879,N_1778,N_1645);
nand U1880 (N_1880,N_1602,N_1775);
and U1881 (N_1881,N_1674,N_1643);
and U1882 (N_1882,N_1741,N_1603);
or U1883 (N_1883,N_1655,N_1675);
nand U1884 (N_1884,N_1725,N_1614);
and U1885 (N_1885,N_1606,N_1780);
and U1886 (N_1886,N_1740,N_1715);
xor U1887 (N_1887,N_1785,N_1760);
nand U1888 (N_1888,N_1652,N_1676);
nand U1889 (N_1889,N_1613,N_1665);
nor U1890 (N_1890,N_1792,N_1742);
and U1891 (N_1891,N_1610,N_1707);
or U1892 (N_1892,N_1698,N_1737);
nand U1893 (N_1893,N_1677,N_1668);
and U1894 (N_1894,N_1650,N_1723);
or U1895 (N_1895,N_1682,N_1754);
nand U1896 (N_1896,N_1640,N_1729);
and U1897 (N_1897,N_1680,N_1756);
or U1898 (N_1898,N_1790,N_1669);
or U1899 (N_1899,N_1710,N_1696);
nor U1900 (N_1900,N_1753,N_1762);
xnor U1901 (N_1901,N_1705,N_1713);
nor U1902 (N_1902,N_1742,N_1788);
and U1903 (N_1903,N_1662,N_1672);
or U1904 (N_1904,N_1750,N_1714);
and U1905 (N_1905,N_1668,N_1705);
nor U1906 (N_1906,N_1791,N_1789);
and U1907 (N_1907,N_1762,N_1719);
and U1908 (N_1908,N_1716,N_1670);
or U1909 (N_1909,N_1772,N_1766);
nor U1910 (N_1910,N_1655,N_1688);
or U1911 (N_1911,N_1767,N_1788);
nor U1912 (N_1912,N_1788,N_1635);
or U1913 (N_1913,N_1788,N_1608);
or U1914 (N_1914,N_1689,N_1741);
nor U1915 (N_1915,N_1634,N_1691);
nor U1916 (N_1916,N_1670,N_1660);
nand U1917 (N_1917,N_1692,N_1662);
and U1918 (N_1918,N_1790,N_1622);
nand U1919 (N_1919,N_1765,N_1601);
or U1920 (N_1920,N_1686,N_1781);
and U1921 (N_1921,N_1761,N_1798);
and U1922 (N_1922,N_1722,N_1614);
and U1923 (N_1923,N_1737,N_1675);
and U1924 (N_1924,N_1646,N_1694);
nand U1925 (N_1925,N_1682,N_1779);
and U1926 (N_1926,N_1639,N_1723);
and U1927 (N_1927,N_1693,N_1630);
nor U1928 (N_1928,N_1629,N_1722);
or U1929 (N_1929,N_1717,N_1785);
and U1930 (N_1930,N_1618,N_1636);
nand U1931 (N_1931,N_1697,N_1704);
and U1932 (N_1932,N_1702,N_1774);
nand U1933 (N_1933,N_1798,N_1782);
and U1934 (N_1934,N_1709,N_1680);
and U1935 (N_1935,N_1697,N_1626);
nand U1936 (N_1936,N_1738,N_1799);
nand U1937 (N_1937,N_1662,N_1744);
or U1938 (N_1938,N_1679,N_1650);
or U1939 (N_1939,N_1788,N_1669);
and U1940 (N_1940,N_1685,N_1683);
and U1941 (N_1941,N_1792,N_1754);
or U1942 (N_1942,N_1656,N_1669);
nor U1943 (N_1943,N_1711,N_1705);
or U1944 (N_1944,N_1612,N_1600);
nor U1945 (N_1945,N_1724,N_1758);
and U1946 (N_1946,N_1670,N_1718);
xnor U1947 (N_1947,N_1769,N_1709);
nand U1948 (N_1948,N_1749,N_1679);
nor U1949 (N_1949,N_1694,N_1721);
and U1950 (N_1950,N_1693,N_1657);
nand U1951 (N_1951,N_1781,N_1779);
or U1952 (N_1952,N_1637,N_1705);
and U1953 (N_1953,N_1785,N_1648);
and U1954 (N_1954,N_1683,N_1708);
nor U1955 (N_1955,N_1603,N_1681);
nor U1956 (N_1956,N_1762,N_1649);
nor U1957 (N_1957,N_1664,N_1765);
nor U1958 (N_1958,N_1782,N_1619);
nor U1959 (N_1959,N_1603,N_1632);
nor U1960 (N_1960,N_1651,N_1733);
nand U1961 (N_1961,N_1767,N_1713);
and U1962 (N_1962,N_1737,N_1655);
and U1963 (N_1963,N_1649,N_1755);
or U1964 (N_1964,N_1682,N_1668);
nand U1965 (N_1965,N_1761,N_1629);
nand U1966 (N_1966,N_1689,N_1639);
or U1967 (N_1967,N_1634,N_1607);
or U1968 (N_1968,N_1698,N_1651);
and U1969 (N_1969,N_1778,N_1795);
nand U1970 (N_1970,N_1707,N_1720);
nor U1971 (N_1971,N_1679,N_1643);
and U1972 (N_1972,N_1664,N_1789);
nand U1973 (N_1973,N_1693,N_1699);
or U1974 (N_1974,N_1719,N_1699);
or U1975 (N_1975,N_1676,N_1757);
nand U1976 (N_1976,N_1613,N_1673);
or U1977 (N_1977,N_1739,N_1651);
nor U1978 (N_1978,N_1682,N_1750);
xnor U1979 (N_1979,N_1716,N_1701);
or U1980 (N_1980,N_1782,N_1754);
nor U1981 (N_1981,N_1796,N_1616);
and U1982 (N_1982,N_1615,N_1623);
nor U1983 (N_1983,N_1756,N_1778);
or U1984 (N_1984,N_1778,N_1730);
nor U1985 (N_1985,N_1708,N_1766);
and U1986 (N_1986,N_1759,N_1630);
nand U1987 (N_1987,N_1638,N_1676);
nand U1988 (N_1988,N_1654,N_1693);
nand U1989 (N_1989,N_1798,N_1755);
and U1990 (N_1990,N_1638,N_1772);
nand U1991 (N_1991,N_1730,N_1603);
nor U1992 (N_1992,N_1792,N_1679);
nor U1993 (N_1993,N_1647,N_1787);
nor U1994 (N_1994,N_1631,N_1772);
and U1995 (N_1995,N_1613,N_1694);
and U1996 (N_1996,N_1674,N_1798);
nand U1997 (N_1997,N_1686,N_1698);
or U1998 (N_1998,N_1780,N_1639);
nand U1999 (N_1999,N_1798,N_1608);
and U2000 (N_2000,N_1847,N_1830);
or U2001 (N_2001,N_1863,N_1822);
nor U2002 (N_2002,N_1894,N_1910);
or U2003 (N_2003,N_1990,N_1834);
or U2004 (N_2004,N_1920,N_1867);
nor U2005 (N_2005,N_1877,N_1911);
nand U2006 (N_2006,N_1996,N_1876);
nand U2007 (N_2007,N_1905,N_1917);
nand U2008 (N_2008,N_1970,N_1831);
or U2009 (N_2009,N_1921,N_1811);
and U2010 (N_2010,N_1854,N_1852);
xnor U2011 (N_2011,N_1860,N_1967);
or U2012 (N_2012,N_1875,N_1940);
nor U2013 (N_2013,N_1907,N_1869);
nand U2014 (N_2014,N_1801,N_1950);
or U2015 (N_2015,N_1953,N_1906);
or U2016 (N_2016,N_1955,N_1957);
and U2017 (N_2017,N_1952,N_1971);
or U2018 (N_2018,N_1930,N_1839);
nand U2019 (N_2019,N_1820,N_1880);
nand U2020 (N_2020,N_1954,N_1825);
nor U2021 (N_2021,N_1848,N_1844);
nand U2022 (N_2022,N_1896,N_1926);
nor U2023 (N_2023,N_1937,N_1829);
and U2024 (N_2024,N_1814,N_1807);
and U2025 (N_2025,N_1895,N_1851);
nand U2026 (N_2026,N_1984,N_1832);
nor U2027 (N_2027,N_1964,N_1802);
nand U2028 (N_2028,N_1972,N_1841);
nand U2029 (N_2029,N_1865,N_1938);
or U2030 (N_2030,N_1886,N_1891);
or U2031 (N_2031,N_1871,N_1857);
and U2032 (N_2032,N_1838,N_1900);
or U2033 (N_2033,N_1809,N_1925);
or U2034 (N_2034,N_1846,N_1824);
and U2035 (N_2035,N_1947,N_1804);
nor U2036 (N_2036,N_1960,N_1962);
nand U2037 (N_2037,N_1874,N_1982);
and U2038 (N_2038,N_1870,N_1916);
nand U2039 (N_2039,N_1988,N_1919);
nand U2040 (N_2040,N_1859,N_1823);
and U2041 (N_2041,N_1902,N_1861);
nor U2042 (N_2042,N_1800,N_1993);
nor U2043 (N_2043,N_1965,N_1977);
or U2044 (N_2044,N_1966,N_1944);
and U2045 (N_2045,N_1855,N_1806);
nor U2046 (N_2046,N_1866,N_1909);
or U2047 (N_2047,N_1961,N_1819);
nor U2048 (N_2048,N_1968,N_1979);
and U2049 (N_2049,N_1978,N_1849);
and U2050 (N_2050,N_1897,N_1959);
nor U2051 (N_2051,N_1812,N_1827);
nor U2052 (N_2052,N_1883,N_1890);
xor U2053 (N_2053,N_1980,N_1974);
and U2054 (N_2054,N_1934,N_1922);
nand U2055 (N_2055,N_1836,N_1803);
nor U2056 (N_2056,N_1892,N_1884);
nand U2057 (N_2057,N_1864,N_1915);
nor U2058 (N_2058,N_1945,N_1912);
and U2059 (N_2059,N_1948,N_1932);
nand U2060 (N_2060,N_1929,N_1885);
nor U2061 (N_2061,N_1997,N_1949);
nand U2062 (N_2062,N_1837,N_1987);
and U2063 (N_2063,N_1914,N_1951);
and U2064 (N_2064,N_1958,N_1941);
and U2065 (N_2065,N_1936,N_1878);
nor U2066 (N_2066,N_1933,N_1998);
or U2067 (N_2067,N_1815,N_1821);
nand U2068 (N_2068,N_1942,N_1858);
or U2069 (N_2069,N_1918,N_1816);
or U2070 (N_2070,N_1999,N_1969);
or U2071 (N_2071,N_1924,N_1981);
xnor U2072 (N_2072,N_1882,N_1985);
nand U2073 (N_2073,N_1850,N_1872);
and U2074 (N_2074,N_1973,N_1893);
xnor U2075 (N_2075,N_1956,N_1992);
nor U2076 (N_2076,N_1901,N_1975);
nand U2077 (N_2077,N_1928,N_1889);
nor U2078 (N_2078,N_1931,N_1826);
nand U2079 (N_2079,N_1983,N_1908);
nand U2080 (N_2080,N_1833,N_1943);
nor U2081 (N_2081,N_1810,N_1904);
xor U2082 (N_2082,N_1853,N_1887);
and U2083 (N_2083,N_1828,N_1888);
nor U2084 (N_2084,N_1903,N_1913);
nand U2085 (N_2085,N_1840,N_1995);
nor U2086 (N_2086,N_1817,N_1873);
or U2087 (N_2087,N_1923,N_1989);
xnor U2088 (N_2088,N_1856,N_1963);
nand U2089 (N_2089,N_1939,N_1986);
nor U2090 (N_2090,N_1991,N_1881);
or U2091 (N_2091,N_1927,N_1845);
and U2092 (N_2092,N_1813,N_1862);
or U2093 (N_2093,N_1935,N_1879);
or U2094 (N_2094,N_1946,N_1898);
nand U2095 (N_2095,N_1835,N_1976);
and U2096 (N_2096,N_1818,N_1842);
and U2097 (N_2097,N_1808,N_1868);
and U2098 (N_2098,N_1805,N_1899);
and U2099 (N_2099,N_1994,N_1843);
nand U2100 (N_2100,N_1895,N_1967);
or U2101 (N_2101,N_1978,N_1831);
nand U2102 (N_2102,N_1816,N_1909);
nor U2103 (N_2103,N_1917,N_1970);
nor U2104 (N_2104,N_1944,N_1895);
nand U2105 (N_2105,N_1905,N_1999);
nand U2106 (N_2106,N_1955,N_1968);
or U2107 (N_2107,N_1830,N_1837);
nand U2108 (N_2108,N_1838,N_1853);
nor U2109 (N_2109,N_1921,N_1978);
nor U2110 (N_2110,N_1922,N_1850);
or U2111 (N_2111,N_1838,N_1982);
nor U2112 (N_2112,N_1856,N_1803);
xnor U2113 (N_2113,N_1886,N_1982);
nor U2114 (N_2114,N_1879,N_1909);
and U2115 (N_2115,N_1802,N_1991);
or U2116 (N_2116,N_1997,N_1810);
nor U2117 (N_2117,N_1881,N_1836);
and U2118 (N_2118,N_1800,N_1912);
and U2119 (N_2119,N_1825,N_1966);
nand U2120 (N_2120,N_1852,N_1809);
and U2121 (N_2121,N_1873,N_1962);
or U2122 (N_2122,N_1928,N_1869);
nor U2123 (N_2123,N_1818,N_1827);
nand U2124 (N_2124,N_1820,N_1803);
nor U2125 (N_2125,N_1839,N_1985);
xor U2126 (N_2126,N_1991,N_1959);
or U2127 (N_2127,N_1804,N_1929);
or U2128 (N_2128,N_1968,N_1990);
or U2129 (N_2129,N_1907,N_1917);
and U2130 (N_2130,N_1982,N_1988);
or U2131 (N_2131,N_1969,N_1895);
nand U2132 (N_2132,N_1956,N_1837);
and U2133 (N_2133,N_1958,N_1880);
or U2134 (N_2134,N_1888,N_1995);
nand U2135 (N_2135,N_1852,N_1923);
or U2136 (N_2136,N_1962,N_1853);
nand U2137 (N_2137,N_1874,N_1836);
nand U2138 (N_2138,N_1937,N_1877);
nor U2139 (N_2139,N_1979,N_1997);
nand U2140 (N_2140,N_1885,N_1915);
nand U2141 (N_2141,N_1894,N_1840);
or U2142 (N_2142,N_1868,N_1984);
nand U2143 (N_2143,N_1827,N_1865);
and U2144 (N_2144,N_1937,N_1982);
and U2145 (N_2145,N_1802,N_1946);
and U2146 (N_2146,N_1952,N_1813);
and U2147 (N_2147,N_1958,N_1909);
and U2148 (N_2148,N_1940,N_1883);
or U2149 (N_2149,N_1889,N_1831);
and U2150 (N_2150,N_1876,N_1906);
or U2151 (N_2151,N_1992,N_1841);
or U2152 (N_2152,N_1933,N_1815);
and U2153 (N_2153,N_1944,N_1945);
and U2154 (N_2154,N_1869,N_1966);
and U2155 (N_2155,N_1943,N_1834);
or U2156 (N_2156,N_1887,N_1992);
nand U2157 (N_2157,N_1970,N_1914);
and U2158 (N_2158,N_1947,N_1989);
and U2159 (N_2159,N_1848,N_1857);
nand U2160 (N_2160,N_1809,N_1998);
nand U2161 (N_2161,N_1957,N_1823);
nand U2162 (N_2162,N_1932,N_1986);
and U2163 (N_2163,N_1927,N_1838);
nand U2164 (N_2164,N_1872,N_1982);
nor U2165 (N_2165,N_1969,N_1982);
and U2166 (N_2166,N_1844,N_1817);
or U2167 (N_2167,N_1944,N_1886);
or U2168 (N_2168,N_1947,N_1842);
or U2169 (N_2169,N_1918,N_1896);
and U2170 (N_2170,N_1971,N_1950);
nor U2171 (N_2171,N_1882,N_1873);
nand U2172 (N_2172,N_1916,N_1958);
nand U2173 (N_2173,N_1858,N_1873);
nand U2174 (N_2174,N_1923,N_1819);
nand U2175 (N_2175,N_1961,N_1937);
or U2176 (N_2176,N_1950,N_1826);
and U2177 (N_2177,N_1919,N_1860);
nor U2178 (N_2178,N_1963,N_1838);
and U2179 (N_2179,N_1995,N_1959);
nor U2180 (N_2180,N_1951,N_1943);
or U2181 (N_2181,N_1938,N_1994);
and U2182 (N_2182,N_1943,N_1923);
or U2183 (N_2183,N_1885,N_1900);
or U2184 (N_2184,N_1875,N_1870);
nand U2185 (N_2185,N_1960,N_1913);
and U2186 (N_2186,N_1868,N_1837);
nand U2187 (N_2187,N_1812,N_1950);
and U2188 (N_2188,N_1809,N_1805);
nand U2189 (N_2189,N_1915,N_1841);
nand U2190 (N_2190,N_1895,N_1919);
and U2191 (N_2191,N_1929,N_1883);
or U2192 (N_2192,N_1870,N_1944);
nor U2193 (N_2193,N_1846,N_1931);
nand U2194 (N_2194,N_1981,N_1828);
and U2195 (N_2195,N_1891,N_1939);
nor U2196 (N_2196,N_1903,N_1921);
and U2197 (N_2197,N_1853,N_1951);
nand U2198 (N_2198,N_1983,N_1826);
nor U2199 (N_2199,N_1815,N_1924);
or U2200 (N_2200,N_2014,N_2145);
and U2201 (N_2201,N_2165,N_2179);
nor U2202 (N_2202,N_2151,N_2170);
and U2203 (N_2203,N_2088,N_2186);
or U2204 (N_2204,N_2099,N_2160);
nand U2205 (N_2205,N_2002,N_2068);
or U2206 (N_2206,N_2150,N_2178);
nand U2207 (N_2207,N_2032,N_2140);
nand U2208 (N_2208,N_2197,N_2015);
nor U2209 (N_2209,N_2110,N_2091);
and U2210 (N_2210,N_2082,N_2117);
nor U2211 (N_2211,N_2005,N_2004);
nor U2212 (N_2212,N_2113,N_2102);
nand U2213 (N_2213,N_2001,N_2153);
nor U2214 (N_2214,N_2027,N_2062);
and U2215 (N_2215,N_2146,N_2035);
nand U2216 (N_2216,N_2006,N_2003);
nand U2217 (N_2217,N_2087,N_2038);
nor U2218 (N_2218,N_2126,N_2132);
nand U2219 (N_2219,N_2022,N_2046);
nand U2220 (N_2220,N_2135,N_2115);
nor U2221 (N_2221,N_2129,N_2039);
and U2222 (N_2222,N_2095,N_2007);
or U2223 (N_2223,N_2085,N_2118);
or U2224 (N_2224,N_2109,N_2112);
and U2225 (N_2225,N_2180,N_2111);
nand U2226 (N_2226,N_2021,N_2159);
or U2227 (N_2227,N_2028,N_2065);
or U2228 (N_2228,N_2054,N_2144);
or U2229 (N_2229,N_2121,N_2119);
or U2230 (N_2230,N_2056,N_2097);
and U2231 (N_2231,N_2012,N_2025);
nand U2232 (N_2232,N_2076,N_2107);
xor U2233 (N_2233,N_2174,N_2182);
or U2234 (N_2234,N_2125,N_2059);
nand U2235 (N_2235,N_2023,N_2133);
and U2236 (N_2236,N_2008,N_2199);
nand U2237 (N_2237,N_2123,N_2024);
nor U2238 (N_2238,N_2010,N_2169);
nand U2239 (N_2239,N_2173,N_2164);
or U2240 (N_2240,N_2189,N_2079);
nand U2241 (N_2241,N_2000,N_2116);
nor U2242 (N_2242,N_2185,N_2093);
nand U2243 (N_2243,N_2090,N_2053);
and U2244 (N_2244,N_2018,N_2019);
or U2245 (N_2245,N_2016,N_2149);
nand U2246 (N_2246,N_2073,N_2063);
and U2247 (N_2247,N_2049,N_2100);
or U2248 (N_2248,N_2136,N_2128);
or U2249 (N_2249,N_2086,N_2171);
nand U2250 (N_2250,N_2080,N_2193);
and U2251 (N_2251,N_2196,N_2184);
or U2252 (N_2252,N_2114,N_2131);
nand U2253 (N_2253,N_2198,N_2029);
nand U2254 (N_2254,N_2120,N_2094);
or U2255 (N_2255,N_2147,N_2168);
and U2256 (N_2256,N_2083,N_2181);
nand U2257 (N_2257,N_2195,N_2074);
and U2258 (N_2258,N_2044,N_2089);
nor U2259 (N_2259,N_2122,N_2011);
and U2260 (N_2260,N_2130,N_2167);
nand U2261 (N_2261,N_2177,N_2139);
nand U2262 (N_2262,N_2047,N_2098);
or U2263 (N_2263,N_2137,N_2043);
or U2264 (N_2264,N_2141,N_2105);
and U2265 (N_2265,N_2134,N_2162);
and U2266 (N_2266,N_2101,N_2072);
nor U2267 (N_2267,N_2048,N_2172);
nor U2268 (N_2268,N_2052,N_2108);
nor U2269 (N_2269,N_2096,N_2064);
nor U2270 (N_2270,N_2084,N_2051);
or U2271 (N_2271,N_2050,N_2166);
nand U2272 (N_2272,N_2157,N_2081);
or U2273 (N_2273,N_2138,N_2030);
and U2274 (N_2274,N_2034,N_2127);
or U2275 (N_2275,N_2192,N_2156);
and U2276 (N_2276,N_2066,N_2055);
nand U2277 (N_2277,N_2026,N_2040);
nand U2278 (N_2278,N_2042,N_2183);
or U2279 (N_2279,N_2077,N_2124);
nand U2280 (N_2280,N_2033,N_2154);
and U2281 (N_2281,N_2092,N_2152);
nor U2282 (N_2282,N_2037,N_2075);
and U2283 (N_2283,N_2041,N_2106);
nor U2284 (N_2284,N_2057,N_2163);
nand U2285 (N_2285,N_2142,N_2103);
or U2286 (N_2286,N_2017,N_2143);
or U2287 (N_2287,N_2031,N_2104);
nand U2288 (N_2288,N_2187,N_2070);
and U2289 (N_2289,N_2148,N_2190);
and U2290 (N_2290,N_2013,N_2158);
or U2291 (N_2291,N_2009,N_2061);
and U2292 (N_2292,N_2069,N_2194);
or U2293 (N_2293,N_2036,N_2155);
or U2294 (N_2294,N_2078,N_2045);
and U2295 (N_2295,N_2175,N_2161);
nand U2296 (N_2296,N_2058,N_2020);
nand U2297 (N_2297,N_2191,N_2060);
nor U2298 (N_2298,N_2071,N_2176);
and U2299 (N_2299,N_2067,N_2188);
nand U2300 (N_2300,N_2072,N_2018);
nand U2301 (N_2301,N_2131,N_2083);
and U2302 (N_2302,N_2052,N_2049);
nor U2303 (N_2303,N_2091,N_2039);
or U2304 (N_2304,N_2043,N_2116);
and U2305 (N_2305,N_2126,N_2008);
and U2306 (N_2306,N_2053,N_2043);
nor U2307 (N_2307,N_2171,N_2054);
and U2308 (N_2308,N_2077,N_2111);
and U2309 (N_2309,N_2157,N_2165);
nand U2310 (N_2310,N_2026,N_2054);
nor U2311 (N_2311,N_2085,N_2128);
nand U2312 (N_2312,N_2195,N_2056);
nor U2313 (N_2313,N_2133,N_2098);
nand U2314 (N_2314,N_2105,N_2172);
nor U2315 (N_2315,N_2111,N_2091);
nor U2316 (N_2316,N_2079,N_2057);
and U2317 (N_2317,N_2106,N_2095);
nand U2318 (N_2318,N_2046,N_2031);
nand U2319 (N_2319,N_2004,N_2041);
nand U2320 (N_2320,N_2112,N_2188);
and U2321 (N_2321,N_2116,N_2186);
nor U2322 (N_2322,N_2170,N_2154);
nor U2323 (N_2323,N_2089,N_2155);
or U2324 (N_2324,N_2138,N_2037);
and U2325 (N_2325,N_2017,N_2112);
or U2326 (N_2326,N_2049,N_2067);
nor U2327 (N_2327,N_2152,N_2166);
nor U2328 (N_2328,N_2102,N_2039);
and U2329 (N_2329,N_2062,N_2078);
and U2330 (N_2330,N_2027,N_2170);
or U2331 (N_2331,N_2062,N_2151);
nor U2332 (N_2332,N_2144,N_2197);
nor U2333 (N_2333,N_2054,N_2037);
nand U2334 (N_2334,N_2010,N_2152);
xnor U2335 (N_2335,N_2144,N_2081);
nor U2336 (N_2336,N_2190,N_2071);
or U2337 (N_2337,N_2010,N_2071);
or U2338 (N_2338,N_2182,N_2000);
and U2339 (N_2339,N_2001,N_2083);
or U2340 (N_2340,N_2161,N_2109);
nand U2341 (N_2341,N_2173,N_2070);
or U2342 (N_2342,N_2163,N_2061);
nand U2343 (N_2343,N_2041,N_2105);
or U2344 (N_2344,N_2032,N_2025);
nor U2345 (N_2345,N_2065,N_2024);
nand U2346 (N_2346,N_2126,N_2097);
or U2347 (N_2347,N_2060,N_2021);
nor U2348 (N_2348,N_2120,N_2167);
nand U2349 (N_2349,N_2042,N_2047);
or U2350 (N_2350,N_2008,N_2010);
and U2351 (N_2351,N_2108,N_2039);
nand U2352 (N_2352,N_2079,N_2154);
or U2353 (N_2353,N_2084,N_2069);
or U2354 (N_2354,N_2128,N_2071);
nand U2355 (N_2355,N_2026,N_2177);
nor U2356 (N_2356,N_2057,N_2175);
and U2357 (N_2357,N_2172,N_2126);
xor U2358 (N_2358,N_2172,N_2085);
or U2359 (N_2359,N_2049,N_2169);
nor U2360 (N_2360,N_2169,N_2066);
nand U2361 (N_2361,N_2155,N_2105);
or U2362 (N_2362,N_2068,N_2088);
or U2363 (N_2363,N_2137,N_2133);
and U2364 (N_2364,N_2185,N_2131);
nand U2365 (N_2365,N_2082,N_2187);
and U2366 (N_2366,N_2187,N_2045);
nor U2367 (N_2367,N_2099,N_2107);
or U2368 (N_2368,N_2165,N_2110);
and U2369 (N_2369,N_2006,N_2014);
xor U2370 (N_2370,N_2064,N_2152);
nand U2371 (N_2371,N_2020,N_2047);
nand U2372 (N_2372,N_2067,N_2172);
nand U2373 (N_2373,N_2118,N_2102);
nor U2374 (N_2374,N_2070,N_2192);
nor U2375 (N_2375,N_2174,N_2058);
nand U2376 (N_2376,N_2001,N_2167);
or U2377 (N_2377,N_2045,N_2091);
nand U2378 (N_2378,N_2090,N_2181);
and U2379 (N_2379,N_2132,N_2056);
nand U2380 (N_2380,N_2035,N_2150);
nand U2381 (N_2381,N_2091,N_2116);
nor U2382 (N_2382,N_2197,N_2057);
nand U2383 (N_2383,N_2178,N_2185);
nand U2384 (N_2384,N_2009,N_2141);
and U2385 (N_2385,N_2198,N_2189);
nor U2386 (N_2386,N_2157,N_2163);
and U2387 (N_2387,N_2035,N_2106);
nor U2388 (N_2388,N_2025,N_2107);
nand U2389 (N_2389,N_2104,N_2109);
nand U2390 (N_2390,N_2156,N_2167);
nand U2391 (N_2391,N_2029,N_2046);
nor U2392 (N_2392,N_2134,N_2015);
nor U2393 (N_2393,N_2067,N_2141);
nand U2394 (N_2394,N_2049,N_2095);
nand U2395 (N_2395,N_2046,N_2149);
or U2396 (N_2396,N_2188,N_2024);
nand U2397 (N_2397,N_2061,N_2162);
and U2398 (N_2398,N_2066,N_2076);
or U2399 (N_2399,N_2117,N_2106);
and U2400 (N_2400,N_2290,N_2297);
or U2401 (N_2401,N_2247,N_2209);
nand U2402 (N_2402,N_2382,N_2293);
nand U2403 (N_2403,N_2278,N_2397);
and U2404 (N_2404,N_2248,N_2213);
nand U2405 (N_2405,N_2203,N_2358);
nor U2406 (N_2406,N_2372,N_2264);
and U2407 (N_2407,N_2243,N_2379);
or U2408 (N_2408,N_2391,N_2318);
nand U2409 (N_2409,N_2289,N_2217);
nand U2410 (N_2410,N_2356,N_2255);
nand U2411 (N_2411,N_2368,N_2244);
or U2412 (N_2412,N_2266,N_2326);
nor U2413 (N_2413,N_2251,N_2359);
xor U2414 (N_2414,N_2336,N_2281);
or U2415 (N_2415,N_2328,N_2259);
and U2416 (N_2416,N_2257,N_2219);
or U2417 (N_2417,N_2341,N_2369);
and U2418 (N_2418,N_2307,N_2348);
or U2419 (N_2419,N_2256,N_2253);
nor U2420 (N_2420,N_2238,N_2353);
nor U2421 (N_2421,N_2323,N_2267);
or U2422 (N_2422,N_2395,N_2374);
and U2423 (N_2423,N_2245,N_2313);
nand U2424 (N_2424,N_2349,N_2310);
nor U2425 (N_2425,N_2311,N_2325);
nand U2426 (N_2426,N_2304,N_2284);
nand U2427 (N_2427,N_2333,N_2319);
xnor U2428 (N_2428,N_2301,N_2321);
nand U2429 (N_2429,N_2373,N_2399);
and U2430 (N_2430,N_2363,N_2335);
nand U2431 (N_2431,N_2233,N_2366);
nand U2432 (N_2432,N_2392,N_2210);
nand U2433 (N_2433,N_2312,N_2381);
or U2434 (N_2434,N_2222,N_2367);
nor U2435 (N_2435,N_2226,N_2246);
nor U2436 (N_2436,N_2296,N_2240);
or U2437 (N_2437,N_2320,N_2273);
and U2438 (N_2438,N_2388,N_2308);
nand U2439 (N_2439,N_2270,N_2315);
or U2440 (N_2440,N_2235,N_2282);
or U2441 (N_2441,N_2221,N_2331);
xor U2442 (N_2442,N_2287,N_2355);
nand U2443 (N_2443,N_2241,N_2305);
or U2444 (N_2444,N_2364,N_2227);
or U2445 (N_2445,N_2211,N_2370);
or U2446 (N_2446,N_2228,N_2215);
nor U2447 (N_2447,N_2218,N_2280);
or U2448 (N_2448,N_2276,N_2376);
nand U2449 (N_2449,N_2380,N_2236);
nand U2450 (N_2450,N_2277,N_2342);
nand U2451 (N_2451,N_2384,N_2263);
nand U2452 (N_2452,N_2377,N_2229);
nor U2453 (N_2453,N_2258,N_2204);
nand U2454 (N_2454,N_2343,N_2324);
or U2455 (N_2455,N_2250,N_2272);
and U2456 (N_2456,N_2274,N_2352);
and U2457 (N_2457,N_2294,N_2214);
xnor U2458 (N_2458,N_2354,N_2316);
and U2459 (N_2459,N_2286,N_2309);
or U2460 (N_2460,N_2393,N_2351);
and U2461 (N_2461,N_2216,N_2299);
nand U2462 (N_2462,N_2298,N_2302);
or U2463 (N_2463,N_2242,N_2231);
nand U2464 (N_2464,N_2317,N_2327);
nand U2465 (N_2465,N_2260,N_2350);
or U2466 (N_2466,N_2371,N_2337);
or U2467 (N_2467,N_2279,N_2254);
nor U2468 (N_2468,N_2334,N_2205);
and U2469 (N_2469,N_2360,N_2265);
and U2470 (N_2470,N_2292,N_2398);
and U2471 (N_2471,N_2232,N_2361);
and U2472 (N_2472,N_2295,N_2249);
or U2473 (N_2473,N_2224,N_2306);
nor U2474 (N_2474,N_2230,N_2362);
or U2475 (N_2475,N_2346,N_2212);
or U2476 (N_2476,N_2252,N_2357);
xnor U2477 (N_2477,N_2303,N_2261);
nor U2478 (N_2478,N_2207,N_2288);
and U2479 (N_2479,N_2268,N_2208);
or U2480 (N_2480,N_2386,N_2378);
nand U2481 (N_2481,N_2220,N_2345);
and U2482 (N_2482,N_2330,N_2375);
or U2483 (N_2483,N_2262,N_2340);
nand U2484 (N_2484,N_2383,N_2385);
nor U2485 (N_2485,N_2300,N_2223);
xnor U2486 (N_2486,N_2237,N_2314);
nor U2487 (N_2487,N_2239,N_2347);
nor U2488 (N_2488,N_2202,N_2234);
nor U2489 (N_2489,N_2344,N_2339);
or U2490 (N_2490,N_2200,N_2285);
nand U2491 (N_2491,N_2338,N_2283);
xnor U2492 (N_2492,N_2365,N_2389);
nor U2493 (N_2493,N_2396,N_2322);
or U2494 (N_2494,N_2225,N_2394);
or U2495 (N_2495,N_2269,N_2390);
nor U2496 (N_2496,N_2201,N_2332);
and U2497 (N_2497,N_2271,N_2291);
nand U2498 (N_2498,N_2329,N_2275);
or U2499 (N_2499,N_2387,N_2206);
or U2500 (N_2500,N_2376,N_2321);
and U2501 (N_2501,N_2375,N_2312);
or U2502 (N_2502,N_2204,N_2365);
nand U2503 (N_2503,N_2366,N_2235);
nand U2504 (N_2504,N_2392,N_2360);
or U2505 (N_2505,N_2350,N_2381);
nor U2506 (N_2506,N_2339,N_2276);
nor U2507 (N_2507,N_2394,N_2338);
nor U2508 (N_2508,N_2254,N_2325);
and U2509 (N_2509,N_2318,N_2324);
and U2510 (N_2510,N_2223,N_2376);
nand U2511 (N_2511,N_2280,N_2251);
nand U2512 (N_2512,N_2346,N_2325);
and U2513 (N_2513,N_2332,N_2282);
or U2514 (N_2514,N_2212,N_2206);
nand U2515 (N_2515,N_2252,N_2354);
nor U2516 (N_2516,N_2230,N_2225);
nand U2517 (N_2517,N_2360,N_2208);
nor U2518 (N_2518,N_2323,N_2326);
nor U2519 (N_2519,N_2325,N_2359);
or U2520 (N_2520,N_2219,N_2290);
nand U2521 (N_2521,N_2390,N_2321);
nor U2522 (N_2522,N_2352,N_2285);
and U2523 (N_2523,N_2254,N_2241);
and U2524 (N_2524,N_2247,N_2235);
nand U2525 (N_2525,N_2295,N_2316);
nand U2526 (N_2526,N_2374,N_2361);
or U2527 (N_2527,N_2209,N_2225);
nor U2528 (N_2528,N_2350,N_2324);
and U2529 (N_2529,N_2218,N_2226);
nand U2530 (N_2530,N_2307,N_2304);
and U2531 (N_2531,N_2304,N_2234);
nor U2532 (N_2532,N_2362,N_2251);
or U2533 (N_2533,N_2398,N_2399);
nor U2534 (N_2534,N_2392,N_2246);
and U2535 (N_2535,N_2393,N_2291);
or U2536 (N_2536,N_2375,N_2365);
nand U2537 (N_2537,N_2241,N_2222);
nor U2538 (N_2538,N_2214,N_2218);
and U2539 (N_2539,N_2385,N_2371);
or U2540 (N_2540,N_2206,N_2307);
nor U2541 (N_2541,N_2242,N_2337);
nor U2542 (N_2542,N_2211,N_2350);
nand U2543 (N_2543,N_2248,N_2246);
and U2544 (N_2544,N_2370,N_2326);
nand U2545 (N_2545,N_2249,N_2332);
nand U2546 (N_2546,N_2394,N_2325);
and U2547 (N_2547,N_2384,N_2302);
nand U2548 (N_2548,N_2278,N_2213);
and U2549 (N_2549,N_2353,N_2285);
nand U2550 (N_2550,N_2342,N_2226);
nand U2551 (N_2551,N_2383,N_2258);
nor U2552 (N_2552,N_2269,N_2330);
and U2553 (N_2553,N_2212,N_2256);
nor U2554 (N_2554,N_2257,N_2341);
nor U2555 (N_2555,N_2261,N_2391);
or U2556 (N_2556,N_2294,N_2289);
and U2557 (N_2557,N_2246,N_2326);
nand U2558 (N_2558,N_2240,N_2396);
nor U2559 (N_2559,N_2214,N_2339);
nand U2560 (N_2560,N_2304,N_2326);
nor U2561 (N_2561,N_2302,N_2231);
nor U2562 (N_2562,N_2382,N_2379);
nand U2563 (N_2563,N_2264,N_2320);
nor U2564 (N_2564,N_2343,N_2305);
nand U2565 (N_2565,N_2361,N_2228);
nand U2566 (N_2566,N_2267,N_2350);
and U2567 (N_2567,N_2387,N_2362);
nor U2568 (N_2568,N_2234,N_2355);
nand U2569 (N_2569,N_2379,N_2340);
nand U2570 (N_2570,N_2263,N_2378);
nor U2571 (N_2571,N_2264,N_2390);
nand U2572 (N_2572,N_2234,N_2210);
and U2573 (N_2573,N_2213,N_2377);
nor U2574 (N_2574,N_2269,N_2234);
and U2575 (N_2575,N_2219,N_2284);
and U2576 (N_2576,N_2268,N_2343);
and U2577 (N_2577,N_2242,N_2219);
nor U2578 (N_2578,N_2209,N_2275);
nand U2579 (N_2579,N_2345,N_2225);
or U2580 (N_2580,N_2234,N_2236);
and U2581 (N_2581,N_2232,N_2358);
and U2582 (N_2582,N_2252,N_2334);
or U2583 (N_2583,N_2286,N_2317);
or U2584 (N_2584,N_2264,N_2237);
nor U2585 (N_2585,N_2205,N_2361);
or U2586 (N_2586,N_2309,N_2306);
nor U2587 (N_2587,N_2289,N_2357);
nand U2588 (N_2588,N_2377,N_2225);
nor U2589 (N_2589,N_2258,N_2271);
and U2590 (N_2590,N_2273,N_2322);
or U2591 (N_2591,N_2378,N_2363);
or U2592 (N_2592,N_2302,N_2300);
nand U2593 (N_2593,N_2312,N_2243);
and U2594 (N_2594,N_2236,N_2247);
nand U2595 (N_2595,N_2236,N_2338);
and U2596 (N_2596,N_2305,N_2315);
or U2597 (N_2597,N_2266,N_2244);
nand U2598 (N_2598,N_2294,N_2350);
and U2599 (N_2599,N_2254,N_2220);
and U2600 (N_2600,N_2504,N_2483);
and U2601 (N_2601,N_2484,N_2417);
nor U2602 (N_2602,N_2427,N_2497);
or U2603 (N_2603,N_2446,N_2403);
xor U2604 (N_2604,N_2480,N_2586);
nand U2605 (N_2605,N_2521,N_2459);
nor U2606 (N_2606,N_2486,N_2493);
or U2607 (N_2607,N_2428,N_2490);
or U2608 (N_2608,N_2592,N_2482);
xor U2609 (N_2609,N_2538,N_2550);
nand U2610 (N_2610,N_2407,N_2501);
nand U2611 (N_2611,N_2476,N_2429);
nand U2612 (N_2612,N_2460,N_2442);
xor U2613 (N_2613,N_2587,N_2522);
or U2614 (N_2614,N_2597,N_2581);
or U2615 (N_2615,N_2579,N_2444);
or U2616 (N_2616,N_2599,N_2445);
and U2617 (N_2617,N_2533,N_2544);
or U2618 (N_2618,N_2479,N_2435);
nand U2619 (N_2619,N_2489,N_2472);
nor U2620 (N_2620,N_2448,N_2548);
or U2621 (N_2621,N_2546,N_2594);
nand U2622 (N_2622,N_2547,N_2418);
and U2623 (N_2623,N_2573,N_2541);
nor U2624 (N_2624,N_2539,N_2419);
nand U2625 (N_2625,N_2416,N_2457);
or U2626 (N_2626,N_2583,N_2474);
or U2627 (N_2627,N_2465,N_2540);
or U2628 (N_2628,N_2409,N_2576);
and U2629 (N_2629,N_2405,N_2414);
nand U2630 (N_2630,N_2590,N_2462);
nor U2631 (N_2631,N_2450,N_2568);
nand U2632 (N_2632,N_2567,N_2505);
or U2633 (N_2633,N_2578,N_2437);
or U2634 (N_2634,N_2454,N_2469);
or U2635 (N_2635,N_2595,N_2570);
nand U2636 (N_2636,N_2481,N_2434);
nor U2637 (N_2637,N_2464,N_2534);
or U2638 (N_2638,N_2408,N_2485);
nor U2639 (N_2639,N_2488,N_2562);
or U2640 (N_2640,N_2496,N_2468);
nand U2641 (N_2641,N_2526,N_2451);
nor U2642 (N_2642,N_2543,N_2421);
and U2643 (N_2643,N_2512,N_2478);
and U2644 (N_2644,N_2574,N_2467);
or U2645 (N_2645,N_2580,N_2412);
or U2646 (N_2646,N_2514,N_2425);
and U2647 (N_2647,N_2402,N_2528);
nor U2648 (N_2648,N_2436,N_2525);
and U2649 (N_2649,N_2532,N_2545);
and U2650 (N_2650,N_2572,N_2558);
or U2651 (N_2651,N_2423,N_2598);
and U2652 (N_2652,N_2589,N_2537);
and U2653 (N_2653,N_2564,N_2531);
and U2654 (N_2654,N_2500,N_2438);
and U2655 (N_2655,N_2499,N_2404);
or U2656 (N_2656,N_2461,N_2523);
nor U2657 (N_2657,N_2432,N_2455);
or U2658 (N_2658,N_2536,N_2506);
and U2659 (N_2659,N_2413,N_2494);
nor U2660 (N_2660,N_2571,N_2440);
nor U2661 (N_2661,N_2400,N_2466);
and U2662 (N_2662,N_2430,N_2519);
nor U2663 (N_2663,N_2591,N_2529);
and U2664 (N_2664,N_2577,N_2458);
or U2665 (N_2665,N_2553,N_2441);
nand U2666 (N_2666,N_2552,N_2565);
nand U2667 (N_2667,N_2551,N_2516);
nand U2668 (N_2668,N_2566,N_2503);
or U2669 (N_2669,N_2433,N_2563);
and U2670 (N_2670,N_2406,N_2509);
nor U2671 (N_2671,N_2511,N_2517);
and U2672 (N_2672,N_2453,N_2561);
nor U2673 (N_2673,N_2492,N_2471);
or U2674 (N_2674,N_2507,N_2575);
nand U2675 (N_2675,N_2498,N_2508);
nor U2676 (N_2676,N_2530,N_2447);
or U2677 (N_2677,N_2582,N_2456);
or U2678 (N_2678,N_2473,N_2470);
nor U2679 (N_2679,N_2554,N_2452);
or U2680 (N_2680,N_2510,N_2410);
or U2681 (N_2681,N_2559,N_2556);
and U2682 (N_2682,N_2513,N_2518);
nor U2683 (N_2683,N_2585,N_2415);
nand U2684 (N_2684,N_2477,N_2596);
or U2685 (N_2685,N_2593,N_2535);
or U2686 (N_2686,N_2401,N_2569);
nor U2687 (N_2687,N_2555,N_2588);
nor U2688 (N_2688,N_2439,N_2475);
nand U2689 (N_2689,N_2515,N_2557);
and U2690 (N_2690,N_2502,N_2431);
and U2691 (N_2691,N_2424,N_2491);
and U2692 (N_2692,N_2520,N_2584);
nor U2693 (N_2693,N_2527,N_2487);
and U2694 (N_2694,N_2560,N_2463);
nand U2695 (N_2695,N_2411,N_2426);
and U2696 (N_2696,N_2549,N_2449);
or U2697 (N_2697,N_2443,N_2495);
nand U2698 (N_2698,N_2524,N_2420);
nor U2699 (N_2699,N_2542,N_2422);
and U2700 (N_2700,N_2579,N_2432);
nor U2701 (N_2701,N_2412,N_2459);
nand U2702 (N_2702,N_2481,N_2528);
nor U2703 (N_2703,N_2483,N_2549);
xnor U2704 (N_2704,N_2500,N_2538);
nor U2705 (N_2705,N_2473,N_2406);
nand U2706 (N_2706,N_2458,N_2533);
and U2707 (N_2707,N_2586,N_2594);
or U2708 (N_2708,N_2401,N_2445);
and U2709 (N_2709,N_2525,N_2440);
and U2710 (N_2710,N_2529,N_2451);
nor U2711 (N_2711,N_2417,N_2539);
nor U2712 (N_2712,N_2591,N_2423);
nand U2713 (N_2713,N_2570,N_2464);
nand U2714 (N_2714,N_2562,N_2586);
or U2715 (N_2715,N_2445,N_2458);
or U2716 (N_2716,N_2494,N_2439);
nor U2717 (N_2717,N_2500,N_2564);
nand U2718 (N_2718,N_2473,N_2519);
or U2719 (N_2719,N_2476,N_2499);
nor U2720 (N_2720,N_2508,N_2555);
or U2721 (N_2721,N_2532,N_2427);
and U2722 (N_2722,N_2533,N_2589);
and U2723 (N_2723,N_2569,N_2487);
nand U2724 (N_2724,N_2445,N_2487);
nand U2725 (N_2725,N_2417,N_2469);
nand U2726 (N_2726,N_2539,N_2529);
nor U2727 (N_2727,N_2508,N_2533);
nor U2728 (N_2728,N_2416,N_2473);
nand U2729 (N_2729,N_2593,N_2460);
or U2730 (N_2730,N_2564,N_2417);
nand U2731 (N_2731,N_2510,N_2472);
nand U2732 (N_2732,N_2461,N_2430);
or U2733 (N_2733,N_2573,N_2403);
xor U2734 (N_2734,N_2454,N_2579);
and U2735 (N_2735,N_2428,N_2565);
nor U2736 (N_2736,N_2448,N_2525);
and U2737 (N_2737,N_2517,N_2484);
nand U2738 (N_2738,N_2528,N_2455);
and U2739 (N_2739,N_2423,N_2546);
and U2740 (N_2740,N_2481,N_2554);
nor U2741 (N_2741,N_2472,N_2430);
or U2742 (N_2742,N_2468,N_2440);
nand U2743 (N_2743,N_2406,N_2479);
and U2744 (N_2744,N_2460,N_2539);
or U2745 (N_2745,N_2530,N_2475);
xnor U2746 (N_2746,N_2415,N_2590);
nor U2747 (N_2747,N_2537,N_2474);
xnor U2748 (N_2748,N_2456,N_2415);
nor U2749 (N_2749,N_2422,N_2583);
xor U2750 (N_2750,N_2581,N_2556);
or U2751 (N_2751,N_2424,N_2593);
nor U2752 (N_2752,N_2421,N_2431);
or U2753 (N_2753,N_2505,N_2515);
nor U2754 (N_2754,N_2536,N_2527);
or U2755 (N_2755,N_2509,N_2569);
or U2756 (N_2756,N_2567,N_2447);
and U2757 (N_2757,N_2585,N_2430);
or U2758 (N_2758,N_2444,N_2577);
nor U2759 (N_2759,N_2504,N_2448);
nor U2760 (N_2760,N_2409,N_2447);
or U2761 (N_2761,N_2548,N_2405);
and U2762 (N_2762,N_2526,N_2504);
xnor U2763 (N_2763,N_2477,N_2409);
and U2764 (N_2764,N_2588,N_2491);
or U2765 (N_2765,N_2506,N_2504);
or U2766 (N_2766,N_2544,N_2516);
or U2767 (N_2767,N_2512,N_2497);
nand U2768 (N_2768,N_2599,N_2524);
or U2769 (N_2769,N_2543,N_2558);
nor U2770 (N_2770,N_2504,N_2515);
nand U2771 (N_2771,N_2517,N_2443);
and U2772 (N_2772,N_2554,N_2550);
nand U2773 (N_2773,N_2577,N_2485);
nor U2774 (N_2774,N_2463,N_2578);
or U2775 (N_2775,N_2593,N_2597);
and U2776 (N_2776,N_2552,N_2475);
or U2777 (N_2777,N_2542,N_2431);
and U2778 (N_2778,N_2548,N_2493);
or U2779 (N_2779,N_2462,N_2564);
nor U2780 (N_2780,N_2567,N_2546);
xnor U2781 (N_2781,N_2485,N_2513);
or U2782 (N_2782,N_2539,N_2494);
nor U2783 (N_2783,N_2401,N_2523);
or U2784 (N_2784,N_2444,N_2591);
nand U2785 (N_2785,N_2429,N_2430);
and U2786 (N_2786,N_2525,N_2549);
or U2787 (N_2787,N_2565,N_2595);
nor U2788 (N_2788,N_2486,N_2512);
nor U2789 (N_2789,N_2573,N_2413);
or U2790 (N_2790,N_2459,N_2577);
nor U2791 (N_2791,N_2598,N_2547);
or U2792 (N_2792,N_2538,N_2591);
nand U2793 (N_2793,N_2411,N_2536);
nor U2794 (N_2794,N_2497,N_2528);
nand U2795 (N_2795,N_2509,N_2414);
and U2796 (N_2796,N_2577,N_2512);
nand U2797 (N_2797,N_2494,N_2448);
and U2798 (N_2798,N_2547,N_2533);
and U2799 (N_2799,N_2505,N_2550);
and U2800 (N_2800,N_2779,N_2662);
nor U2801 (N_2801,N_2735,N_2665);
or U2802 (N_2802,N_2768,N_2691);
nand U2803 (N_2803,N_2618,N_2601);
nor U2804 (N_2804,N_2666,N_2743);
nand U2805 (N_2805,N_2647,N_2639);
or U2806 (N_2806,N_2713,N_2635);
nor U2807 (N_2807,N_2751,N_2786);
nor U2808 (N_2808,N_2798,N_2692);
or U2809 (N_2809,N_2678,N_2625);
nand U2810 (N_2810,N_2795,N_2773);
and U2811 (N_2811,N_2796,N_2634);
and U2812 (N_2812,N_2734,N_2696);
nor U2813 (N_2813,N_2753,N_2704);
nor U2814 (N_2814,N_2623,N_2684);
nand U2815 (N_2815,N_2643,N_2648);
and U2816 (N_2816,N_2785,N_2714);
or U2817 (N_2817,N_2663,N_2730);
or U2818 (N_2818,N_2664,N_2650);
and U2819 (N_2819,N_2789,N_2737);
nand U2820 (N_2820,N_2661,N_2780);
or U2821 (N_2821,N_2695,N_2660);
or U2822 (N_2822,N_2712,N_2640);
nor U2823 (N_2823,N_2788,N_2631);
and U2824 (N_2824,N_2705,N_2668);
and U2825 (N_2825,N_2703,N_2769);
and U2826 (N_2826,N_2702,N_2670);
or U2827 (N_2827,N_2701,N_2711);
nand U2828 (N_2828,N_2629,N_2641);
or U2829 (N_2829,N_2699,N_2633);
nand U2830 (N_2830,N_2676,N_2693);
or U2831 (N_2831,N_2775,N_2729);
nand U2832 (N_2832,N_2642,N_2607);
and U2833 (N_2833,N_2709,N_2638);
and U2834 (N_2834,N_2742,N_2716);
and U2835 (N_2835,N_2739,N_2762);
or U2836 (N_2836,N_2710,N_2609);
and U2837 (N_2837,N_2763,N_2784);
and U2838 (N_2838,N_2671,N_2694);
nor U2839 (N_2839,N_2604,N_2690);
or U2840 (N_2840,N_2681,N_2777);
or U2841 (N_2841,N_2677,N_2752);
nand U2842 (N_2842,N_2636,N_2760);
and U2843 (N_2843,N_2700,N_2720);
nand U2844 (N_2844,N_2630,N_2611);
and U2845 (N_2845,N_2799,N_2746);
or U2846 (N_2846,N_2721,N_2610);
or U2847 (N_2847,N_2603,N_2717);
and U2848 (N_2848,N_2637,N_2715);
and U2849 (N_2849,N_2680,N_2787);
nand U2850 (N_2850,N_2645,N_2756);
nor U2851 (N_2851,N_2605,N_2616);
nand U2852 (N_2852,N_2600,N_2657);
nor U2853 (N_2853,N_2646,N_2778);
and U2854 (N_2854,N_2765,N_2672);
or U2855 (N_2855,N_2740,N_2653);
nor U2856 (N_2856,N_2685,N_2621);
nand U2857 (N_2857,N_2741,N_2736);
nor U2858 (N_2858,N_2669,N_2602);
or U2859 (N_2859,N_2770,N_2683);
and U2860 (N_2860,N_2651,N_2745);
nand U2861 (N_2861,N_2771,N_2744);
and U2862 (N_2862,N_2731,N_2649);
nand U2863 (N_2863,N_2759,N_2679);
and U2864 (N_2864,N_2761,N_2726);
or U2865 (N_2865,N_2733,N_2624);
and U2866 (N_2866,N_2619,N_2675);
and U2867 (N_2867,N_2686,N_2772);
or U2868 (N_2868,N_2755,N_2622);
and U2869 (N_2869,N_2767,N_2764);
xor U2870 (N_2870,N_2688,N_2632);
nor U2871 (N_2871,N_2738,N_2724);
nor U2872 (N_2872,N_2781,N_2750);
nand U2873 (N_2873,N_2725,N_2783);
or U2874 (N_2874,N_2774,N_2689);
and U2875 (N_2875,N_2732,N_2612);
or U2876 (N_2876,N_2727,N_2707);
or U2877 (N_2877,N_2687,N_2708);
nor U2878 (N_2878,N_2748,N_2656);
or U2879 (N_2879,N_2794,N_2791);
nor U2880 (N_2880,N_2614,N_2682);
nand U2881 (N_2881,N_2644,N_2793);
nor U2882 (N_2882,N_2613,N_2674);
and U2883 (N_2883,N_2790,N_2728);
or U2884 (N_2884,N_2749,N_2615);
and U2885 (N_2885,N_2627,N_2617);
or U2886 (N_2886,N_2620,N_2658);
and U2887 (N_2887,N_2608,N_2766);
or U2888 (N_2888,N_2655,N_2757);
or U2889 (N_2889,N_2776,N_2654);
nand U2890 (N_2890,N_2667,N_2673);
and U2891 (N_2891,N_2719,N_2628);
or U2892 (N_2892,N_2797,N_2754);
or U2893 (N_2893,N_2606,N_2718);
and U2894 (N_2894,N_2747,N_2723);
nand U2895 (N_2895,N_2659,N_2697);
and U2896 (N_2896,N_2782,N_2706);
and U2897 (N_2897,N_2792,N_2758);
nand U2898 (N_2898,N_2626,N_2698);
or U2899 (N_2899,N_2652,N_2722);
or U2900 (N_2900,N_2622,N_2672);
nand U2901 (N_2901,N_2674,N_2629);
nor U2902 (N_2902,N_2759,N_2641);
nand U2903 (N_2903,N_2731,N_2674);
and U2904 (N_2904,N_2757,N_2695);
or U2905 (N_2905,N_2782,N_2724);
or U2906 (N_2906,N_2676,N_2777);
nor U2907 (N_2907,N_2674,N_2634);
nand U2908 (N_2908,N_2654,N_2799);
or U2909 (N_2909,N_2653,N_2615);
or U2910 (N_2910,N_2603,N_2606);
nor U2911 (N_2911,N_2721,N_2709);
or U2912 (N_2912,N_2601,N_2689);
or U2913 (N_2913,N_2733,N_2727);
nand U2914 (N_2914,N_2696,N_2685);
and U2915 (N_2915,N_2772,N_2736);
nand U2916 (N_2916,N_2700,N_2607);
and U2917 (N_2917,N_2616,N_2622);
nor U2918 (N_2918,N_2658,N_2714);
or U2919 (N_2919,N_2719,N_2662);
nor U2920 (N_2920,N_2767,N_2630);
and U2921 (N_2921,N_2772,N_2703);
nor U2922 (N_2922,N_2637,N_2677);
or U2923 (N_2923,N_2601,N_2657);
nand U2924 (N_2924,N_2733,N_2741);
and U2925 (N_2925,N_2643,N_2781);
nand U2926 (N_2926,N_2727,N_2637);
or U2927 (N_2927,N_2759,N_2790);
nand U2928 (N_2928,N_2653,N_2799);
nand U2929 (N_2929,N_2669,N_2611);
or U2930 (N_2930,N_2646,N_2631);
or U2931 (N_2931,N_2616,N_2779);
and U2932 (N_2932,N_2655,N_2770);
or U2933 (N_2933,N_2765,N_2799);
nand U2934 (N_2934,N_2733,N_2791);
or U2935 (N_2935,N_2626,N_2664);
xor U2936 (N_2936,N_2775,N_2657);
or U2937 (N_2937,N_2664,N_2622);
nor U2938 (N_2938,N_2706,N_2662);
nand U2939 (N_2939,N_2652,N_2641);
and U2940 (N_2940,N_2744,N_2706);
nand U2941 (N_2941,N_2680,N_2770);
nor U2942 (N_2942,N_2693,N_2633);
nand U2943 (N_2943,N_2677,N_2672);
and U2944 (N_2944,N_2617,N_2741);
nor U2945 (N_2945,N_2637,N_2601);
or U2946 (N_2946,N_2647,N_2605);
nand U2947 (N_2947,N_2767,N_2780);
nand U2948 (N_2948,N_2747,N_2610);
nor U2949 (N_2949,N_2630,N_2605);
nand U2950 (N_2950,N_2707,N_2795);
nand U2951 (N_2951,N_2665,N_2778);
or U2952 (N_2952,N_2668,N_2650);
nand U2953 (N_2953,N_2694,N_2685);
nand U2954 (N_2954,N_2636,N_2721);
nor U2955 (N_2955,N_2774,N_2728);
nand U2956 (N_2956,N_2716,N_2684);
or U2957 (N_2957,N_2784,N_2641);
or U2958 (N_2958,N_2731,N_2719);
and U2959 (N_2959,N_2644,N_2721);
or U2960 (N_2960,N_2631,N_2658);
or U2961 (N_2961,N_2782,N_2722);
nor U2962 (N_2962,N_2760,N_2656);
and U2963 (N_2963,N_2603,N_2657);
and U2964 (N_2964,N_2694,N_2691);
and U2965 (N_2965,N_2786,N_2642);
or U2966 (N_2966,N_2636,N_2674);
xor U2967 (N_2967,N_2759,N_2765);
and U2968 (N_2968,N_2694,N_2798);
and U2969 (N_2969,N_2721,N_2626);
and U2970 (N_2970,N_2644,N_2629);
or U2971 (N_2971,N_2667,N_2637);
nor U2972 (N_2972,N_2772,N_2603);
nand U2973 (N_2973,N_2623,N_2604);
and U2974 (N_2974,N_2747,N_2641);
xnor U2975 (N_2975,N_2721,N_2701);
and U2976 (N_2976,N_2742,N_2634);
nor U2977 (N_2977,N_2655,N_2765);
or U2978 (N_2978,N_2754,N_2612);
nor U2979 (N_2979,N_2667,N_2741);
or U2980 (N_2980,N_2795,N_2618);
nand U2981 (N_2981,N_2729,N_2602);
and U2982 (N_2982,N_2735,N_2773);
nor U2983 (N_2983,N_2619,N_2760);
and U2984 (N_2984,N_2665,N_2601);
nand U2985 (N_2985,N_2684,N_2698);
or U2986 (N_2986,N_2774,N_2760);
nand U2987 (N_2987,N_2631,N_2707);
or U2988 (N_2988,N_2604,N_2687);
or U2989 (N_2989,N_2791,N_2631);
nor U2990 (N_2990,N_2664,N_2764);
nand U2991 (N_2991,N_2736,N_2629);
and U2992 (N_2992,N_2672,N_2682);
nor U2993 (N_2993,N_2722,N_2727);
or U2994 (N_2994,N_2765,N_2735);
or U2995 (N_2995,N_2693,N_2665);
nand U2996 (N_2996,N_2793,N_2755);
and U2997 (N_2997,N_2783,N_2722);
or U2998 (N_2998,N_2641,N_2632);
xor U2999 (N_2999,N_2767,N_2615);
or UO_0 (O_0,N_2962,N_2836);
and UO_1 (O_1,N_2942,N_2975);
or UO_2 (O_2,N_2988,N_2832);
or UO_3 (O_3,N_2810,N_2896);
nor UO_4 (O_4,N_2841,N_2901);
or UO_5 (O_5,N_2869,N_2818);
nand UO_6 (O_6,N_2976,N_2813);
or UO_7 (O_7,N_2827,N_2912);
nand UO_8 (O_8,N_2982,N_2862);
nor UO_9 (O_9,N_2989,N_2898);
and UO_10 (O_10,N_2908,N_2829);
nand UO_11 (O_11,N_2801,N_2890);
nor UO_12 (O_12,N_2899,N_2949);
or UO_13 (O_13,N_2874,N_2876);
nor UO_14 (O_14,N_2958,N_2947);
nor UO_15 (O_15,N_2815,N_2806);
and UO_16 (O_16,N_2822,N_2918);
nor UO_17 (O_17,N_2994,N_2968);
and UO_18 (O_18,N_2933,N_2940);
nor UO_19 (O_19,N_2845,N_2819);
nand UO_20 (O_20,N_2807,N_2866);
nand UO_21 (O_21,N_2846,N_2973);
and UO_22 (O_22,N_2914,N_2858);
nor UO_23 (O_23,N_2946,N_2930);
or UO_24 (O_24,N_2906,N_2931);
nor UO_25 (O_25,N_2916,N_2999);
nand UO_26 (O_26,N_2978,N_2913);
nand UO_27 (O_27,N_2991,N_2888);
nor UO_28 (O_28,N_2844,N_2969);
and UO_29 (O_29,N_2996,N_2941);
nor UO_30 (O_30,N_2920,N_2902);
and UO_31 (O_31,N_2824,N_2970);
and UO_32 (O_32,N_2826,N_2909);
or UO_33 (O_33,N_2803,N_2850);
or UO_34 (O_34,N_2963,N_2839);
or UO_35 (O_35,N_2873,N_2922);
nand UO_36 (O_36,N_2915,N_2879);
nand UO_37 (O_37,N_2883,N_2848);
nor UO_38 (O_38,N_2871,N_2838);
and UO_39 (O_39,N_2800,N_2894);
nand UO_40 (O_40,N_2997,N_2837);
nand UO_41 (O_41,N_2972,N_2878);
nand UO_42 (O_42,N_2959,N_2863);
and UO_43 (O_43,N_2855,N_2884);
or UO_44 (O_44,N_2980,N_2971);
or UO_45 (O_45,N_2814,N_2811);
nor UO_46 (O_46,N_2937,N_2965);
and UO_47 (O_47,N_2833,N_2842);
nor UO_48 (O_48,N_2923,N_2917);
and UO_49 (O_49,N_2910,N_2950);
or UO_50 (O_50,N_2864,N_2919);
or UO_51 (O_51,N_2956,N_2992);
or UO_52 (O_52,N_2926,N_2820);
or UO_53 (O_53,N_2979,N_2854);
nor UO_54 (O_54,N_2867,N_2875);
or UO_55 (O_55,N_2828,N_2944);
and UO_56 (O_56,N_2857,N_2924);
nand UO_57 (O_57,N_2843,N_2840);
nor UO_58 (O_58,N_2851,N_2952);
or UO_59 (O_59,N_2966,N_2987);
xnor UO_60 (O_60,N_2895,N_2823);
or UO_61 (O_61,N_2974,N_2877);
or UO_62 (O_62,N_2961,N_2904);
nand UO_63 (O_63,N_2900,N_2954);
nor UO_64 (O_64,N_2897,N_2903);
nor UO_65 (O_65,N_2891,N_2804);
or UO_66 (O_66,N_2886,N_2849);
and UO_67 (O_67,N_2967,N_2868);
or UO_68 (O_68,N_2925,N_2808);
nor UO_69 (O_69,N_2831,N_2834);
nor UO_70 (O_70,N_2860,N_2935);
or UO_71 (O_71,N_2932,N_2943);
nor UO_72 (O_72,N_2847,N_2889);
nand UO_73 (O_73,N_2921,N_2859);
nor UO_74 (O_74,N_2939,N_2852);
and UO_75 (O_75,N_2957,N_2835);
nand UO_76 (O_76,N_2955,N_2882);
and UO_77 (O_77,N_2983,N_2853);
or UO_78 (O_78,N_2936,N_2984);
or UO_79 (O_79,N_2893,N_2981);
or UO_80 (O_80,N_2830,N_2887);
nand UO_81 (O_81,N_2977,N_2964);
and UO_82 (O_82,N_2990,N_2805);
or UO_83 (O_83,N_2960,N_2928);
nand UO_84 (O_84,N_2872,N_2985);
nand UO_85 (O_85,N_2934,N_2995);
and UO_86 (O_86,N_2948,N_2802);
or UO_87 (O_87,N_2911,N_2938);
nor UO_88 (O_88,N_2880,N_2945);
xnor UO_89 (O_89,N_2951,N_2812);
and UO_90 (O_90,N_2998,N_2929);
nor UO_91 (O_91,N_2809,N_2816);
nor UO_92 (O_92,N_2907,N_2927);
nor UO_93 (O_93,N_2892,N_2861);
or UO_94 (O_94,N_2993,N_2821);
nor UO_95 (O_95,N_2856,N_2986);
and UO_96 (O_96,N_2870,N_2885);
nand UO_97 (O_97,N_2825,N_2817);
or UO_98 (O_98,N_2953,N_2905);
and UO_99 (O_99,N_2881,N_2865);
nand UO_100 (O_100,N_2884,N_2979);
nor UO_101 (O_101,N_2917,N_2989);
or UO_102 (O_102,N_2941,N_2828);
nand UO_103 (O_103,N_2817,N_2940);
nand UO_104 (O_104,N_2832,N_2938);
or UO_105 (O_105,N_2911,N_2939);
nand UO_106 (O_106,N_2832,N_2866);
nor UO_107 (O_107,N_2807,N_2883);
or UO_108 (O_108,N_2897,N_2917);
and UO_109 (O_109,N_2842,N_2814);
nand UO_110 (O_110,N_2846,N_2986);
nor UO_111 (O_111,N_2849,N_2864);
or UO_112 (O_112,N_2865,N_2809);
nor UO_113 (O_113,N_2827,N_2989);
nor UO_114 (O_114,N_2814,N_2896);
nand UO_115 (O_115,N_2887,N_2954);
nand UO_116 (O_116,N_2836,N_2812);
and UO_117 (O_117,N_2957,N_2942);
or UO_118 (O_118,N_2859,N_2880);
nor UO_119 (O_119,N_2969,N_2938);
and UO_120 (O_120,N_2998,N_2875);
and UO_121 (O_121,N_2869,N_2979);
xnor UO_122 (O_122,N_2967,N_2817);
or UO_123 (O_123,N_2981,N_2826);
nor UO_124 (O_124,N_2876,N_2808);
nor UO_125 (O_125,N_2897,N_2922);
or UO_126 (O_126,N_2957,N_2992);
nor UO_127 (O_127,N_2879,N_2817);
or UO_128 (O_128,N_2903,N_2893);
nor UO_129 (O_129,N_2811,N_2935);
nand UO_130 (O_130,N_2964,N_2892);
nand UO_131 (O_131,N_2816,N_2975);
nand UO_132 (O_132,N_2841,N_2978);
nor UO_133 (O_133,N_2802,N_2876);
xor UO_134 (O_134,N_2803,N_2916);
nor UO_135 (O_135,N_2918,N_2924);
nand UO_136 (O_136,N_2848,N_2935);
xor UO_137 (O_137,N_2914,N_2885);
or UO_138 (O_138,N_2875,N_2921);
and UO_139 (O_139,N_2933,N_2979);
nor UO_140 (O_140,N_2808,N_2956);
nor UO_141 (O_141,N_2981,N_2938);
or UO_142 (O_142,N_2884,N_2853);
nor UO_143 (O_143,N_2819,N_2862);
nor UO_144 (O_144,N_2902,N_2948);
nand UO_145 (O_145,N_2925,N_2965);
and UO_146 (O_146,N_2872,N_2870);
nand UO_147 (O_147,N_2820,N_2846);
xor UO_148 (O_148,N_2966,N_2814);
xnor UO_149 (O_149,N_2802,N_2945);
nor UO_150 (O_150,N_2960,N_2959);
xnor UO_151 (O_151,N_2832,N_2950);
and UO_152 (O_152,N_2955,N_2952);
nand UO_153 (O_153,N_2810,N_2856);
and UO_154 (O_154,N_2801,N_2989);
or UO_155 (O_155,N_2894,N_2873);
or UO_156 (O_156,N_2863,N_2877);
nand UO_157 (O_157,N_2954,N_2862);
or UO_158 (O_158,N_2970,N_2898);
nor UO_159 (O_159,N_2945,N_2957);
and UO_160 (O_160,N_2882,N_2897);
nand UO_161 (O_161,N_2989,N_2836);
nor UO_162 (O_162,N_2874,N_2964);
nor UO_163 (O_163,N_2987,N_2989);
or UO_164 (O_164,N_2878,N_2850);
nand UO_165 (O_165,N_2831,N_2966);
and UO_166 (O_166,N_2950,N_2874);
or UO_167 (O_167,N_2894,N_2839);
nor UO_168 (O_168,N_2871,N_2805);
nor UO_169 (O_169,N_2954,N_2905);
nand UO_170 (O_170,N_2800,N_2896);
nand UO_171 (O_171,N_2971,N_2966);
and UO_172 (O_172,N_2915,N_2855);
nand UO_173 (O_173,N_2854,N_2874);
or UO_174 (O_174,N_2890,N_2812);
or UO_175 (O_175,N_2851,N_2902);
xnor UO_176 (O_176,N_2887,N_2815);
nand UO_177 (O_177,N_2965,N_2894);
and UO_178 (O_178,N_2999,N_2955);
nor UO_179 (O_179,N_2984,N_2807);
nand UO_180 (O_180,N_2964,N_2827);
or UO_181 (O_181,N_2872,N_2806);
nor UO_182 (O_182,N_2869,N_2996);
and UO_183 (O_183,N_2805,N_2969);
and UO_184 (O_184,N_2864,N_2983);
xnor UO_185 (O_185,N_2856,N_2929);
nand UO_186 (O_186,N_2975,N_2885);
nand UO_187 (O_187,N_2876,N_2932);
and UO_188 (O_188,N_2900,N_2873);
and UO_189 (O_189,N_2911,N_2928);
or UO_190 (O_190,N_2882,N_2947);
and UO_191 (O_191,N_2806,N_2972);
or UO_192 (O_192,N_2870,N_2810);
and UO_193 (O_193,N_2989,N_2922);
and UO_194 (O_194,N_2850,N_2860);
nor UO_195 (O_195,N_2889,N_2824);
and UO_196 (O_196,N_2800,N_2950);
and UO_197 (O_197,N_2814,N_2853);
nor UO_198 (O_198,N_2959,N_2950);
xnor UO_199 (O_199,N_2852,N_2807);
and UO_200 (O_200,N_2960,N_2996);
or UO_201 (O_201,N_2886,N_2882);
nor UO_202 (O_202,N_2951,N_2911);
or UO_203 (O_203,N_2967,N_2823);
or UO_204 (O_204,N_2899,N_2897);
nor UO_205 (O_205,N_2982,N_2949);
or UO_206 (O_206,N_2987,N_2916);
nor UO_207 (O_207,N_2877,N_2819);
nand UO_208 (O_208,N_2891,N_2868);
nand UO_209 (O_209,N_2925,N_2836);
nor UO_210 (O_210,N_2929,N_2951);
nand UO_211 (O_211,N_2822,N_2897);
nor UO_212 (O_212,N_2928,N_2912);
nor UO_213 (O_213,N_2887,N_2971);
nand UO_214 (O_214,N_2840,N_2810);
nor UO_215 (O_215,N_2981,N_2869);
nor UO_216 (O_216,N_2978,N_2980);
nand UO_217 (O_217,N_2946,N_2970);
nor UO_218 (O_218,N_2932,N_2848);
nand UO_219 (O_219,N_2806,N_2855);
nand UO_220 (O_220,N_2910,N_2807);
nand UO_221 (O_221,N_2947,N_2995);
or UO_222 (O_222,N_2813,N_2860);
nor UO_223 (O_223,N_2925,N_2888);
or UO_224 (O_224,N_2861,N_2986);
and UO_225 (O_225,N_2802,N_2854);
or UO_226 (O_226,N_2974,N_2930);
nand UO_227 (O_227,N_2825,N_2904);
or UO_228 (O_228,N_2852,N_2918);
nor UO_229 (O_229,N_2829,N_2904);
or UO_230 (O_230,N_2850,N_2909);
and UO_231 (O_231,N_2956,N_2863);
and UO_232 (O_232,N_2800,N_2843);
and UO_233 (O_233,N_2972,N_2856);
nor UO_234 (O_234,N_2997,N_2864);
and UO_235 (O_235,N_2910,N_2922);
and UO_236 (O_236,N_2922,N_2866);
nor UO_237 (O_237,N_2920,N_2844);
nand UO_238 (O_238,N_2866,N_2959);
nor UO_239 (O_239,N_2897,N_2905);
or UO_240 (O_240,N_2929,N_2876);
xnor UO_241 (O_241,N_2838,N_2947);
nor UO_242 (O_242,N_2968,N_2920);
nor UO_243 (O_243,N_2837,N_2993);
nand UO_244 (O_244,N_2905,N_2932);
nand UO_245 (O_245,N_2948,N_2950);
and UO_246 (O_246,N_2826,N_2952);
or UO_247 (O_247,N_2927,N_2817);
nand UO_248 (O_248,N_2894,N_2908);
and UO_249 (O_249,N_2817,N_2995);
nor UO_250 (O_250,N_2882,N_2939);
nand UO_251 (O_251,N_2891,N_2887);
nor UO_252 (O_252,N_2857,N_2804);
and UO_253 (O_253,N_2914,N_2886);
and UO_254 (O_254,N_2817,N_2996);
and UO_255 (O_255,N_2898,N_2872);
or UO_256 (O_256,N_2972,N_2990);
nor UO_257 (O_257,N_2872,N_2849);
nor UO_258 (O_258,N_2877,N_2800);
and UO_259 (O_259,N_2894,N_2802);
and UO_260 (O_260,N_2840,N_2927);
and UO_261 (O_261,N_2915,N_2951);
nor UO_262 (O_262,N_2937,N_2930);
or UO_263 (O_263,N_2802,N_2885);
nand UO_264 (O_264,N_2807,N_2834);
nor UO_265 (O_265,N_2873,N_2996);
nor UO_266 (O_266,N_2823,N_2828);
and UO_267 (O_267,N_2863,N_2908);
and UO_268 (O_268,N_2978,N_2917);
nand UO_269 (O_269,N_2852,N_2878);
and UO_270 (O_270,N_2938,N_2828);
or UO_271 (O_271,N_2938,N_2887);
nand UO_272 (O_272,N_2948,N_2899);
and UO_273 (O_273,N_2870,N_2890);
xor UO_274 (O_274,N_2924,N_2862);
or UO_275 (O_275,N_2959,N_2900);
xor UO_276 (O_276,N_2992,N_2844);
nor UO_277 (O_277,N_2860,N_2909);
or UO_278 (O_278,N_2925,N_2866);
and UO_279 (O_279,N_2966,N_2809);
or UO_280 (O_280,N_2961,N_2850);
nor UO_281 (O_281,N_2942,N_2952);
nand UO_282 (O_282,N_2983,N_2928);
nand UO_283 (O_283,N_2850,N_2920);
and UO_284 (O_284,N_2954,N_2801);
nor UO_285 (O_285,N_2956,N_2944);
or UO_286 (O_286,N_2951,N_2823);
nand UO_287 (O_287,N_2959,N_2986);
nor UO_288 (O_288,N_2862,N_2883);
or UO_289 (O_289,N_2827,N_2889);
or UO_290 (O_290,N_2813,N_2935);
and UO_291 (O_291,N_2908,N_2978);
nand UO_292 (O_292,N_2953,N_2981);
nand UO_293 (O_293,N_2946,N_2904);
nor UO_294 (O_294,N_2987,N_2985);
or UO_295 (O_295,N_2988,N_2915);
nand UO_296 (O_296,N_2905,N_2836);
nand UO_297 (O_297,N_2965,N_2960);
nor UO_298 (O_298,N_2841,N_2804);
and UO_299 (O_299,N_2958,N_2979);
or UO_300 (O_300,N_2950,N_2845);
or UO_301 (O_301,N_2808,N_2944);
nand UO_302 (O_302,N_2911,N_2829);
nand UO_303 (O_303,N_2952,N_2973);
and UO_304 (O_304,N_2823,N_2881);
nor UO_305 (O_305,N_2834,N_2808);
and UO_306 (O_306,N_2981,N_2824);
and UO_307 (O_307,N_2930,N_2892);
nor UO_308 (O_308,N_2993,N_2896);
and UO_309 (O_309,N_2982,N_2888);
xnor UO_310 (O_310,N_2949,N_2881);
nor UO_311 (O_311,N_2879,N_2897);
or UO_312 (O_312,N_2991,N_2885);
nand UO_313 (O_313,N_2850,N_2852);
nand UO_314 (O_314,N_2864,N_2975);
nand UO_315 (O_315,N_2909,N_2815);
nand UO_316 (O_316,N_2898,N_2862);
nand UO_317 (O_317,N_2867,N_2948);
nand UO_318 (O_318,N_2924,N_2901);
nor UO_319 (O_319,N_2958,N_2806);
and UO_320 (O_320,N_2940,N_2991);
nand UO_321 (O_321,N_2915,N_2956);
and UO_322 (O_322,N_2961,N_2838);
xnor UO_323 (O_323,N_2812,N_2942);
nor UO_324 (O_324,N_2917,N_2882);
nand UO_325 (O_325,N_2826,N_2925);
nand UO_326 (O_326,N_2822,N_2998);
nor UO_327 (O_327,N_2966,N_2954);
or UO_328 (O_328,N_2961,N_2945);
nor UO_329 (O_329,N_2841,N_2871);
nand UO_330 (O_330,N_2847,N_2803);
and UO_331 (O_331,N_2918,N_2940);
and UO_332 (O_332,N_2986,N_2923);
or UO_333 (O_333,N_2895,N_2809);
nand UO_334 (O_334,N_2907,N_2966);
xor UO_335 (O_335,N_2810,N_2885);
nor UO_336 (O_336,N_2982,N_2844);
nand UO_337 (O_337,N_2906,N_2832);
nand UO_338 (O_338,N_2976,N_2905);
and UO_339 (O_339,N_2986,N_2918);
nor UO_340 (O_340,N_2807,N_2879);
nor UO_341 (O_341,N_2908,N_2890);
nor UO_342 (O_342,N_2952,N_2874);
nor UO_343 (O_343,N_2833,N_2820);
and UO_344 (O_344,N_2844,N_2874);
nand UO_345 (O_345,N_2984,N_2819);
and UO_346 (O_346,N_2818,N_2846);
and UO_347 (O_347,N_2928,N_2986);
and UO_348 (O_348,N_2831,N_2841);
or UO_349 (O_349,N_2838,N_2932);
xnor UO_350 (O_350,N_2902,N_2954);
and UO_351 (O_351,N_2842,N_2930);
nor UO_352 (O_352,N_2893,N_2806);
or UO_353 (O_353,N_2967,N_2856);
and UO_354 (O_354,N_2991,N_2870);
or UO_355 (O_355,N_2973,N_2950);
nor UO_356 (O_356,N_2866,N_2926);
and UO_357 (O_357,N_2970,N_2906);
nand UO_358 (O_358,N_2923,N_2948);
or UO_359 (O_359,N_2896,N_2965);
nand UO_360 (O_360,N_2979,N_2987);
nand UO_361 (O_361,N_2827,N_2839);
xnor UO_362 (O_362,N_2895,N_2892);
xor UO_363 (O_363,N_2814,N_2802);
nor UO_364 (O_364,N_2902,N_2930);
or UO_365 (O_365,N_2997,N_2854);
and UO_366 (O_366,N_2842,N_2977);
nand UO_367 (O_367,N_2910,N_2842);
nor UO_368 (O_368,N_2947,N_2875);
nand UO_369 (O_369,N_2946,N_2861);
nor UO_370 (O_370,N_2932,N_2927);
or UO_371 (O_371,N_2818,N_2939);
nor UO_372 (O_372,N_2872,N_2877);
nor UO_373 (O_373,N_2966,N_2949);
nor UO_374 (O_374,N_2906,N_2838);
nand UO_375 (O_375,N_2869,N_2937);
and UO_376 (O_376,N_2926,N_2922);
or UO_377 (O_377,N_2896,N_2923);
or UO_378 (O_378,N_2969,N_2953);
nand UO_379 (O_379,N_2891,N_2924);
and UO_380 (O_380,N_2994,N_2989);
nor UO_381 (O_381,N_2818,N_2882);
or UO_382 (O_382,N_2954,N_2880);
nand UO_383 (O_383,N_2891,N_2935);
xor UO_384 (O_384,N_2922,N_2902);
and UO_385 (O_385,N_2978,N_2867);
or UO_386 (O_386,N_2821,N_2970);
or UO_387 (O_387,N_2958,N_2959);
nand UO_388 (O_388,N_2882,N_2830);
or UO_389 (O_389,N_2803,N_2950);
or UO_390 (O_390,N_2970,N_2825);
nor UO_391 (O_391,N_2999,N_2806);
or UO_392 (O_392,N_2975,N_2919);
and UO_393 (O_393,N_2944,N_2805);
and UO_394 (O_394,N_2928,N_2985);
nand UO_395 (O_395,N_2963,N_2940);
nor UO_396 (O_396,N_2865,N_2998);
nand UO_397 (O_397,N_2806,N_2987);
or UO_398 (O_398,N_2995,N_2843);
nand UO_399 (O_399,N_2944,N_2985);
nor UO_400 (O_400,N_2957,N_2805);
nand UO_401 (O_401,N_2852,N_2933);
and UO_402 (O_402,N_2988,N_2943);
and UO_403 (O_403,N_2937,N_2964);
or UO_404 (O_404,N_2907,N_2822);
nand UO_405 (O_405,N_2965,N_2978);
or UO_406 (O_406,N_2994,N_2824);
and UO_407 (O_407,N_2901,N_2886);
nor UO_408 (O_408,N_2851,N_2934);
or UO_409 (O_409,N_2885,N_2869);
or UO_410 (O_410,N_2826,N_2972);
nand UO_411 (O_411,N_2842,N_2871);
or UO_412 (O_412,N_2903,N_2961);
nand UO_413 (O_413,N_2922,N_2823);
nor UO_414 (O_414,N_2979,N_2816);
nor UO_415 (O_415,N_2847,N_2947);
nand UO_416 (O_416,N_2808,N_2889);
nor UO_417 (O_417,N_2881,N_2845);
or UO_418 (O_418,N_2996,N_2994);
nor UO_419 (O_419,N_2923,N_2807);
or UO_420 (O_420,N_2813,N_2918);
or UO_421 (O_421,N_2901,N_2875);
nand UO_422 (O_422,N_2805,N_2891);
xor UO_423 (O_423,N_2922,N_2986);
nand UO_424 (O_424,N_2823,N_2864);
nand UO_425 (O_425,N_2978,N_2910);
nand UO_426 (O_426,N_2984,N_2842);
or UO_427 (O_427,N_2824,N_2925);
nor UO_428 (O_428,N_2948,N_2897);
and UO_429 (O_429,N_2895,N_2822);
nand UO_430 (O_430,N_2980,N_2955);
or UO_431 (O_431,N_2942,N_2876);
and UO_432 (O_432,N_2969,N_2941);
nand UO_433 (O_433,N_2907,N_2805);
or UO_434 (O_434,N_2996,N_2804);
nor UO_435 (O_435,N_2891,N_2952);
nor UO_436 (O_436,N_2885,N_2867);
nor UO_437 (O_437,N_2920,N_2936);
and UO_438 (O_438,N_2928,N_2800);
and UO_439 (O_439,N_2915,N_2830);
nor UO_440 (O_440,N_2857,N_2983);
and UO_441 (O_441,N_2862,N_2994);
or UO_442 (O_442,N_2909,N_2824);
nand UO_443 (O_443,N_2977,N_2887);
or UO_444 (O_444,N_2839,N_2876);
and UO_445 (O_445,N_2948,N_2837);
nand UO_446 (O_446,N_2803,N_2894);
nand UO_447 (O_447,N_2823,N_2811);
nand UO_448 (O_448,N_2921,N_2950);
and UO_449 (O_449,N_2904,N_2802);
or UO_450 (O_450,N_2897,N_2901);
and UO_451 (O_451,N_2867,N_2931);
nor UO_452 (O_452,N_2852,N_2818);
and UO_453 (O_453,N_2985,N_2951);
xor UO_454 (O_454,N_2804,N_2893);
and UO_455 (O_455,N_2966,N_2882);
or UO_456 (O_456,N_2964,N_2844);
nor UO_457 (O_457,N_2998,N_2921);
and UO_458 (O_458,N_2829,N_2919);
and UO_459 (O_459,N_2930,N_2987);
and UO_460 (O_460,N_2869,N_2820);
and UO_461 (O_461,N_2924,N_2904);
xnor UO_462 (O_462,N_2805,N_2926);
nor UO_463 (O_463,N_2808,N_2949);
nor UO_464 (O_464,N_2820,N_2847);
nand UO_465 (O_465,N_2829,N_2999);
nand UO_466 (O_466,N_2802,N_2831);
or UO_467 (O_467,N_2951,N_2845);
and UO_468 (O_468,N_2856,N_2832);
nand UO_469 (O_469,N_2934,N_2886);
nor UO_470 (O_470,N_2819,N_2970);
xnor UO_471 (O_471,N_2902,N_2955);
or UO_472 (O_472,N_2973,N_2847);
nor UO_473 (O_473,N_2905,N_2827);
nand UO_474 (O_474,N_2826,N_2970);
or UO_475 (O_475,N_2909,N_2827);
and UO_476 (O_476,N_2950,N_2876);
or UO_477 (O_477,N_2869,N_2806);
and UO_478 (O_478,N_2850,N_2889);
nor UO_479 (O_479,N_2955,N_2946);
and UO_480 (O_480,N_2920,N_2852);
nand UO_481 (O_481,N_2962,N_2933);
and UO_482 (O_482,N_2869,N_2946);
and UO_483 (O_483,N_2861,N_2965);
nand UO_484 (O_484,N_2835,N_2818);
and UO_485 (O_485,N_2912,N_2932);
nor UO_486 (O_486,N_2812,N_2956);
and UO_487 (O_487,N_2855,N_2995);
and UO_488 (O_488,N_2916,N_2885);
or UO_489 (O_489,N_2913,N_2811);
or UO_490 (O_490,N_2880,N_2830);
or UO_491 (O_491,N_2965,N_2813);
nor UO_492 (O_492,N_2860,N_2806);
nand UO_493 (O_493,N_2835,N_2946);
and UO_494 (O_494,N_2949,N_2973);
nand UO_495 (O_495,N_2951,N_2905);
and UO_496 (O_496,N_2967,N_2833);
or UO_497 (O_497,N_2838,N_2956);
nor UO_498 (O_498,N_2918,N_2978);
or UO_499 (O_499,N_2994,N_2963);
endmodule