module basic_750_5000_1000_50_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
or U0 (N_0,In_418,In_430);
or U1 (N_1,In_159,In_282);
xnor U2 (N_2,In_300,In_467);
or U3 (N_3,In_709,In_315);
nor U4 (N_4,In_223,In_453);
xor U5 (N_5,In_407,In_131);
nor U6 (N_6,In_263,In_555);
xnor U7 (N_7,In_334,In_594);
nor U8 (N_8,In_231,In_224);
xor U9 (N_9,In_563,In_400);
or U10 (N_10,In_83,In_689);
xnor U11 (N_11,In_139,In_180);
and U12 (N_12,In_616,In_416);
nand U13 (N_13,In_218,In_659);
or U14 (N_14,In_299,In_185);
nor U15 (N_15,In_373,In_646);
nor U16 (N_16,In_370,In_245);
nor U17 (N_17,In_423,In_623);
xor U18 (N_18,In_253,In_130);
nand U19 (N_19,In_177,In_437);
xor U20 (N_20,In_698,In_55);
or U21 (N_21,In_236,In_265);
nor U22 (N_22,In_431,In_643);
and U23 (N_23,In_404,In_70);
nor U24 (N_24,In_192,In_444);
nor U25 (N_25,In_511,In_560);
or U26 (N_26,In_483,In_655);
and U27 (N_27,In_741,In_417);
and U28 (N_28,In_533,In_266);
and U29 (N_29,In_637,In_516);
or U30 (N_30,In_743,In_474);
nor U31 (N_31,In_550,In_612);
and U32 (N_32,In_35,In_119);
and U33 (N_33,In_175,In_4);
nand U34 (N_34,In_96,In_471);
or U35 (N_35,In_145,In_584);
or U36 (N_36,In_552,In_269);
nand U37 (N_37,In_522,In_675);
and U38 (N_38,In_41,In_439);
nand U39 (N_39,In_667,In_480);
nand U40 (N_40,In_498,In_127);
or U41 (N_41,In_290,In_335);
or U42 (N_42,In_491,In_461);
or U43 (N_43,In_733,In_559);
nand U44 (N_44,In_607,In_206);
nor U45 (N_45,In_604,In_90);
or U46 (N_46,In_247,In_71);
or U47 (N_47,In_7,In_688);
or U48 (N_48,In_62,In_634);
nor U49 (N_49,In_5,In_78);
nor U50 (N_50,In_387,In_57);
or U51 (N_51,In_451,In_295);
and U52 (N_52,In_297,In_326);
or U53 (N_53,In_46,In_557);
nand U54 (N_54,In_617,In_500);
xnor U55 (N_55,In_434,In_54);
xor U56 (N_56,In_399,In_221);
nand U57 (N_57,In_599,In_720);
xor U58 (N_58,In_731,In_31);
nand U59 (N_59,In_531,In_580);
nand U60 (N_60,In_254,In_1);
and U61 (N_61,In_314,In_454);
and U62 (N_62,In_678,In_135);
or U63 (N_63,In_296,In_190);
or U64 (N_64,In_261,In_229);
nand U65 (N_65,In_548,In_134);
nor U66 (N_66,In_279,In_18);
and U67 (N_67,In_450,In_647);
or U68 (N_68,In_302,In_16);
and U69 (N_69,In_132,In_22);
and U70 (N_70,In_694,In_242);
xor U71 (N_71,In_74,In_39);
or U72 (N_72,In_631,In_150);
nand U73 (N_73,In_736,In_167);
or U74 (N_74,In_87,In_285);
and U75 (N_75,In_625,In_528);
nor U76 (N_76,In_686,In_85);
nand U77 (N_77,In_475,In_657);
xnor U78 (N_78,In_244,In_158);
or U79 (N_79,In_88,In_69);
nor U80 (N_80,In_38,In_252);
and U81 (N_81,In_372,In_495);
nand U82 (N_82,In_421,In_432);
and U83 (N_83,In_577,In_457);
nand U84 (N_84,In_298,In_628);
nor U85 (N_85,In_730,In_144);
nand U86 (N_86,In_609,In_316);
nor U87 (N_87,In_642,In_734);
nor U88 (N_88,In_259,In_355);
or U89 (N_89,In_749,In_714);
and U90 (N_90,In_228,In_148);
nor U91 (N_91,In_358,In_389);
and U92 (N_92,In_72,In_492);
and U93 (N_93,In_402,In_436);
nand U94 (N_94,In_11,In_391);
xor U95 (N_95,In_225,In_708);
nand U96 (N_96,In_582,In_411);
nor U97 (N_97,In_43,In_571);
nor U98 (N_98,In_705,In_465);
xnor U99 (N_99,In_307,In_497);
nor U100 (N_100,In_204,In_652);
nand U101 (N_101,In_321,In_469);
and U102 (N_102,In_517,In_745);
and U103 (N_103,In_293,N_20);
nand U104 (N_104,In_63,In_210);
nor U105 (N_105,In_674,In_502);
nand U106 (N_106,In_360,In_510);
xor U107 (N_107,In_546,In_726);
nor U108 (N_108,In_352,In_662);
xor U109 (N_109,N_53,N_46);
or U110 (N_110,In_565,In_157);
nand U111 (N_111,In_92,In_633);
or U112 (N_112,In_128,In_410);
nor U113 (N_113,N_36,In_15);
nand U114 (N_114,In_408,In_716);
and U115 (N_115,In_320,N_24);
nand U116 (N_116,In_84,N_45);
and U117 (N_117,In_424,N_86);
nand U118 (N_118,In_137,In_112);
or U119 (N_119,In_45,In_549);
nor U120 (N_120,In_386,In_147);
or U121 (N_121,In_178,In_611);
nor U122 (N_122,In_380,In_508);
or U123 (N_123,N_54,N_14);
nor U124 (N_124,In_171,N_30);
xor U125 (N_125,N_70,In_684);
or U126 (N_126,In_537,In_356);
and U127 (N_127,In_354,In_196);
xor U128 (N_128,In_328,In_523);
and U129 (N_129,In_205,N_49);
or U130 (N_130,In_473,In_717);
nor U131 (N_131,In_213,In_547);
nor U132 (N_132,In_448,In_362);
xor U133 (N_133,In_273,In_108);
or U134 (N_134,In_327,N_58);
and U135 (N_135,In_110,In_215);
nor U136 (N_136,In_479,In_258);
nor U137 (N_137,In_692,In_207);
or U138 (N_138,In_375,In_673);
nor U139 (N_139,In_233,In_696);
or U140 (N_140,N_5,In_458);
nand U141 (N_141,In_301,In_388);
or U142 (N_142,In_313,In_366);
nand U143 (N_143,In_650,In_154);
nor U144 (N_144,In_590,In_406);
and U145 (N_145,N_66,In_239);
and U146 (N_146,In_163,N_15);
xnor U147 (N_147,In_525,In_262);
and U148 (N_148,In_341,In_371);
or U149 (N_149,In_182,In_166);
nor U150 (N_150,In_146,N_90);
and U151 (N_151,In_200,In_34);
or U152 (N_152,In_735,In_660);
or U153 (N_153,In_82,In_707);
or U154 (N_154,In_597,In_447);
and U155 (N_155,In_61,In_287);
nand U156 (N_156,In_427,In_428);
nand U157 (N_157,In_484,In_713);
and U158 (N_158,In_250,In_544);
xor U159 (N_159,In_2,N_43);
nor U160 (N_160,In_197,In_32);
nand U161 (N_161,In_703,In_203);
xnor U162 (N_162,In_746,In_656);
xor U163 (N_163,In_649,In_398);
or U164 (N_164,In_103,In_700);
and U165 (N_165,In_379,In_68);
or U166 (N_166,In_569,In_573);
and U167 (N_167,N_93,In_710);
and U168 (N_168,N_37,In_575);
and U169 (N_169,In_173,In_91);
and U170 (N_170,In_246,In_73);
nand U171 (N_171,In_440,In_121);
nor U172 (N_172,In_363,In_169);
xnor U173 (N_173,N_3,In_392);
and U174 (N_174,In_13,N_60);
nor U175 (N_175,In_396,In_638);
nor U176 (N_176,In_564,In_319);
or U177 (N_177,In_568,In_585);
and U178 (N_178,In_101,In_455);
nand U179 (N_179,In_342,In_501);
nor U180 (N_180,In_219,In_118);
and U181 (N_181,In_477,In_76);
nand U182 (N_182,In_142,In_325);
nor U183 (N_183,In_340,In_3);
nand U184 (N_184,N_99,In_438);
or U185 (N_185,In_309,In_286);
or U186 (N_186,In_586,In_227);
and U187 (N_187,In_504,In_385);
nor U188 (N_188,In_317,N_75);
or U189 (N_189,In_8,N_6);
or U190 (N_190,N_27,N_55);
nand U191 (N_191,In_681,In_718);
nor U192 (N_192,N_4,In_330);
or U193 (N_193,In_291,In_125);
or U194 (N_194,N_21,N_2);
nand U195 (N_195,In_645,In_728);
xnor U196 (N_196,In_737,In_111);
or U197 (N_197,In_742,In_562);
or U198 (N_198,In_126,N_79);
and U199 (N_199,In_499,In_530);
nor U200 (N_200,In_419,N_31);
nor U201 (N_201,In_202,In_496);
or U202 (N_202,In_30,N_134);
xnor U203 (N_203,In_676,In_622);
and U204 (N_204,N_128,In_217);
or U205 (N_205,In_351,N_82);
nor U206 (N_206,N_153,In_214);
and U207 (N_207,In_632,In_220);
and U208 (N_208,N_144,In_48);
or U209 (N_209,N_171,In_506);
xor U210 (N_210,N_0,In_394);
nand U211 (N_211,In_64,N_72);
or U212 (N_212,N_42,In_268);
nand U213 (N_213,In_605,In_165);
and U214 (N_214,In_603,In_472);
and U215 (N_215,In_486,In_89);
or U216 (N_216,In_318,In_117);
and U217 (N_217,In_711,In_106);
nor U218 (N_218,In_280,In_168);
nand U219 (N_219,N_56,In_635);
nand U220 (N_220,In_536,In_312);
nand U221 (N_221,In_255,In_264);
nand U222 (N_222,In_271,In_114);
nor U223 (N_223,N_71,In_294);
and U224 (N_224,N_109,In_687);
or U225 (N_225,In_376,N_156);
and U226 (N_226,N_125,N_91);
or U227 (N_227,In_435,In_143);
or U228 (N_228,N_40,In_727);
and U229 (N_229,In_683,N_8);
and U230 (N_230,In_24,In_725);
nand U231 (N_231,In_129,In_413);
xor U232 (N_232,In_50,In_589);
nand U233 (N_233,In_658,In_212);
nand U234 (N_234,In_397,In_606);
and U235 (N_235,In_378,In_403);
nor U236 (N_236,In_67,In_724);
or U237 (N_237,In_100,In_27);
nand U238 (N_238,In_598,In_627);
xnor U239 (N_239,In_482,N_136);
and U240 (N_240,In_693,N_157);
nor U241 (N_241,N_183,In_574);
or U242 (N_242,In_140,N_39);
nand U243 (N_243,In_97,In_256);
or U244 (N_244,In_554,N_123);
or U245 (N_245,N_154,In_579);
and U246 (N_246,In_591,In_561);
xor U247 (N_247,In_476,N_139);
xnor U248 (N_248,In_60,In_353);
nand U249 (N_249,N_11,In_518);
and U250 (N_250,N_104,In_304);
or U251 (N_251,In_104,In_14);
or U252 (N_252,In_270,In_524);
nor U253 (N_253,In_519,N_41);
xor U254 (N_254,N_197,In_748);
and U255 (N_255,In_234,N_165);
and U256 (N_256,In_512,In_534);
nor U257 (N_257,In_503,In_695);
or U258 (N_258,In_374,In_174);
and U259 (N_259,In_93,In_654);
and U260 (N_260,In_542,N_68);
and U261 (N_261,In_505,In_42);
and U262 (N_262,N_63,In_209);
xnor U263 (N_263,In_723,In_420);
nor U264 (N_264,In_226,In_0);
xor U265 (N_265,In_583,N_110);
and U266 (N_266,In_629,In_529);
or U267 (N_267,N_89,N_181);
nand U268 (N_268,In_669,In_729);
nand U269 (N_269,In_237,In_288);
or U270 (N_270,In_36,N_147);
xor U271 (N_271,In_333,In_551);
or U272 (N_272,N_13,N_169);
or U273 (N_273,In_156,In_464);
xnor U274 (N_274,In_80,In_164);
or U275 (N_275,N_25,N_103);
or U276 (N_276,N_199,In_614);
and U277 (N_277,In_59,N_150);
nand U278 (N_278,In_682,In_665);
or U279 (N_279,In_47,In_115);
xor U280 (N_280,In_558,In_161);
nand U281 (N_281,In_367,N_191);
xnor U282 (N_282,N_112,In_459);
or U283 (N_283,N_194,In_640);
and U284 (N_284,In_429,N_61);
and U285 (N_285,In_541,In_198);
and U286 (N_286,N_67,In_556);
or U287 (N_287,In_332,In_740);
nand U288 (N_288,In_278,N_163);
xnor U289 (N_289,In_240,In_193);
xor U290 (N_290,In_608,N_155);
and U291 (N_291,In_699,N_159);
and U292 (N_292,In_677,In_306);
or U293 (N_293,In_343,N_160);
and U294 (N_294,In_535,In_425);
and U295 (N_295,N_77,In_243);
nor U296 (N_296,In_572,In_216);
xor U297 (N_297,In_109,In_593);
and U298 (N_298,In_17,In_347);
or U299 (N_299,N_118,In_383);
and U300 (N_300,In_415,N_166);
and U301 (N_301,In_576,In_641);
and U302 (N_302,In_162,N_140);
nor U303 (N_303,In_702,In_160);
nor U304 (N_304,In_81,N_272);
and U305 (N_305,N_88,N_265);
nor U306 (N_306,In_25,In_172);
or U307 (N_307,N_278,N_216);
or U308 (N_308,In_666,N_202);
nand U309 (N_309,In_412,N_106);
and U310 (N_310,N_117,N_64);
xnor U311 (N_311,In_445,In_113);
nand U312 (N_312,In_222,N_222);
or U313 (N_313,In_201,N_207);
nor U314 (N_314,In_191,In_630);
nand U315 (N_315,N_241,N_224);
and U316 (N_316,N_257,N_95);
nor U317 (N_317,In_53,N_213);
nor U318 (N_318,In_520,N_279);
nor U319 (N_319,In_618,In_456);
xor U320 (N_320,N_271,In_697);
nand U321 (N_321,In_323,In_284);
nand U322 (N_322,N_275,N_115);
nand U323 (N_323,In_671,N_261);
and U324 (N_324,N_253,N_227);
and U325 (N_325,N_196,In_600);
and U326 (N_326,N_290,In_116);
and U327 (N_327,In_248,N_195);
nand U328 (N_328,In_712,N_244);
nand U329 (N_329,In_377,N_149);
nor U330 (N_330,N_220,In_208);
nor U331 (N_331,In_149,N_208);
and U332 (N_332,N_284,In_189);
nand U333 (N_333,In_20,N_18);
xnor U334 (N_334,In_545,In_283);
or U335 (N_335,In_251,In_365);
xnor U336 (N_336,N_262,In_310);
nand U337 (N_337,N_83,In_526);
nor U338 (N_338,In_732,N_175);
nor U339 (N_339,N_269,N_137);
or U340 (N_340,In_357,In_706);
nor U341 (N_341,In_513,In_442);
nand U342 (N_342,N_289,N_38);
nor U343 (N_343,In_449,In_680);
and U344 (N_344,In_107,In_170);
nor U345 (N_345,In_744,In_303);
nor U346 (N_346,N_172,N_287);
and U347 (N_347,In_540,N_236);
xnor U348 (N_348,In_663,In_94);
nor U349 (N_349,N_142,N_246);
and U350 (N_350,In_99,In_685);
and U351 (N_351,N_254,N_80);
xnor U352 (N_352,N_17,N_260);
and U353 (N_353,N_215,In_183);
xnor U354 (N_354,In_601,In_514);
nor U355 (N_355,N_288,N_48);
nand U356 (N_356,In_120,In_691);
xnor U357 (N_357,N_273,N_107);
nand U358 (N_358,N_111,In_260);
and U359 (N_359,N_209,In_179);
and U360 (N_360,In_701,N_131);
or U361 (N_361,N_205,N_250);
or U362 (N_362,N_62,N_186);
nand U363 (N_363,N_285,In_308);
nand U364 (N_364,In_747,N_276);
nand U365 (N_365,In_468,In_493);
nand U366 (N_366,In_141,N_81);
nand U367 (N_367,In_739,N_247);
nand U368 (N_368,In_23,In_274);
xnor U369 (N_369,In_602,N_235);
nor U370 (N_370,N_180,N_74);
nor U371 (N_371,In_267,In_305);
xor U372 (N_372,In_384,In_452);
nor U373 (N_373,In_336,N_239);
nand U374 (N_374,In_653,N_19);
xor U375 (N_375,N_167,In_136);
or U376 (N_376,N_228,N_78);
nand U377 (N_377,N_277,In_329);
nand U378 (N_378,N_263,In_348);
nor U379 (N_379,N_264,In_10);
or U380 (N_380,N_85,In_19);
and U381 (N_381,In_199,In_77);
nand U382 (N_382,N_162,N_210);
nand U383 (N_383,N_286,In_485);
xor U384 (N_384,In_52,N_174);
nor U385 (N_385,N_124,N_76);
and U386 (N_386,In_238,In_588);
or U387 (N_387,In_395,N_258);
or U388 (N_388,In_66,N_179);
and U389 (N_389,In_344,N_242);
and U390 (N_390,N_29,In_393);
nor U391 (N_391,N_192,In_369);
or U392 (N_392,In_44,In_578);
and U393 (N_393,N_32,In_49);
nor U394 (N_394,N_141,In_672);
nor U395 (N_395,N_151,In_257);
xor U396 (N_396,N_59,In_401);
nand U397 (N_397,In_521,In_409);
nor U398 (N_398,In_721,In_211);
and U399 (N_399,In_382,N_267);
nor U400 (N_400,N_308,In_338);
xnor U401 (N_401,N_152,In_194);
or U402 (N_402,In_639,N_292);
nand U403 (N_403,N_399,N_35);
nor U404 (N_404,In_592,N_204);
nand U405 (N_405,N_301,In_232);
and U406 (N_406,In_184,N_302);
nor U407 (N_407,N_190,In_668);
xnor U408 (N_408,N_395,In_28);
and U409 (N_409,N_105,In_487);
or U410 (N_410,N_296,N_353);
or U411 (N_411,N_316,In_426);
and U412 (N_412,In_79,In_626);
or U413 (N_413,In_292,N_252);
nand U414 (N_414,N_33,N_359);
and U415 (N_415,N_374,N_217);
or U416 (N_416,N_300,In_651);
and U417 (N_417,N_304,N_309);
or U418 (N_418,N_297,N_321);
and U419 (N_419,N_211,In_241);
nand U420 (N_420,In_345,In_181);
nor U421 (N_421,N_231,In_478);
nand U422 (N_422,In_176,N_384);
or U423 (N_423,N_237,N_346);
and U424 (N_424,In_613,In_414);
nor U425 (N_425,N_341,N_7);
and U426 (N_426,In_98,In_422);
nand U427 (N_427,N_87,N_355);
xor U428 (N_428,N_393,In_75);
nor U429 (N_429,N_331,N_92);
and U430 (N_430,N_363,N_303);
nand U431 (N_431,In_507,N_396);
and U432 (N_432,N_361,N_102);
or U433 (N_433,In_102,In_187);
or U434 (N_434,N_184,N_193);
nand U435 (N_435,N_378,In_364);
nand U436 (N_436,In_704,In_494);
and U437 (N_437,N_338,N_73);
xor U438 (N_438,N_130,N_12);
or U439 (N_439,N_357,N_214);
nand U440 (N_440,N_376,N_323);
nand U441 (N_441,N_266,In_311);
nand U442 (N_442,N_94,In_124);
nand U443 (N_443,In_230,N_203);
nand U444 (N_444,In_65,N_101);
nand U445 (N_445,N_291,In_610);
and U446 (N_446,N_343,N_379);
nor U447 (N_447,N_337,N_294);
and U448 (N_448,In_532,N_344);
nand U449 (N_449,In_539,N_315);
or U450 (N_450,N_348,N_234);
or U451 (N_451,N_188,In_123);
nor U452 (N_452,N_219,N_114);
or U453 (N_453,N_282,In_339);
nand U454 (N_454,N_375,In_470);
or U455 (N_455,In_719,N_397);
and U456 (N_456,In_26,N_340);
or U457 (N_457,N_122,In_481);
or U458 (N_458,N_248,N_176);
xnor U459 (N_459,In_490,N_119);
nor U460 (N_460,N_365,N_394);
and U461 (N_461,In_289,N_386);
and U462 (N_462,N_358,In_488);
nor U463 (N_463,N_9,N_281);
or U464 (N_464,In_276,In_58);
nand U465 (N_465,N_377,N_34);
and U466 (N_466,N_10,N_121);
and U467 (N_467,N_69,In_138);
nand U468 (N_468,N_178,N_373);
nor U469 (N_469,In_433,N_135);
nand U470 (N_470,N_310,In_443);
and U471 (N_471,In_466,In_21);
nand U472 (N_472,N_47,N_326);
nand U473 (N_473,N_317,In_619);
and U474 (N_474,N_382,In_272);
xnor U475 (N_475,N_116,In_570);
nand U476 (N_476,In_56,N_295);
nor U477 (N_477,N_245,N_177);
and U478 (N_478,N_387,N_356);
or U479 (N_479,N_372,N_280);
nor U480 (N_480,N_330,N_311);
nand U481 (N_481,N_133,In_441);
nand U482 (N_482,N_232,In_661);
nand U483 (N_483,N_170,N_84);
nor U484 (N_484,In_133,N_367);
xnor U485 (N_485,In_621,N_333);
and U486 (N_486,N_100,In_463);
nor U487 (N_487,In_33,N_336);
and U488 (N_488,N_371,N_50);
nand U489 (N_489,N_240,N_398);
and U490 (N_490,N_380,In_664);
nand U491 (N_491,In_6,N_327);
nand U492 (N_492,N_226,In_346);
or U493 (N_493,N_249,N_345);
nor U494 (N_494,In_644,N_364);
nand U495 (N_495,In_543,In_636);
or U496 (N_496,N_324,N_366);
and U497 (N_497,N_65,N_352);
and U498 (N_498,N_225,N_293);
nor U499 (N_499,In_151,N_158);
nor U500 (N_500,N_230,N_16);
xnor U501 (N_501,N_26,N_489);
and U502 (N_502,N_385,N_475);
nand U503 (N_503,N_256,N_1);
or U504 (N_504,N_187,N_435);
or U505 (N_505,N_497,In_281);
xnor U506 (N_506,In_349,N_498);
nand U507 (N_507,N_437,N_132);
or U508 (N_508,In_515,N_462);
or U509 (N_509,N_441,N_415);
and U510 (N_510,N_113,N_270);
or U511 (N_511,In_509,N_318);
and U512 (N_512,N_108,N_447);
nand U513 (N_513,In_405,In_648);
and U514 (N_514,N_454,N_419);
and U515 (N_515,N_305,N_476);
nand U516 (N_516,N_468,N_459);
nand U517 (N_517,N_450,N_362);
or U518 (N_518,N_238,N_201);
and U519 (N_519,N_51,In_624);
or U520 (N_520,N_413,N_168);
nor U521 (N_521,In_152,In_105);
and U522 (N_522,N_464,N_423);
xnor U523 (N_523,N_456,In_381);
or U524 (N_524,N_416,N_442);
nand U525 (N_525,N_421,N_138);
or U526 (N_526,N_471,In_581);
nor U527 (N_527,N_313,N_97);
nand U528 (N_528,N_306,N_329);
and U529 (N_529,N_255,N_392);
or U530 (N_530,N_492,In_337);
and U531 (N_531,N_482,In_324);
xor U532 (N_532,In_188,N_325);
xor U533 (N_533,N_438,N_161);
xor U534 (N_534,N_467,N_409);
nand U535 (N_535,N_443,N_173);
and U536 (N_536,In_446,N_446);
or U537 (N_537,In_331,N_406);
and U538 (N_538,N_453,In_715);
nor U539 (N_539,N_390,N_473);
nand U540 (N_540,In_153,N_460);
or U541 (N_541,In_738,N_414);
xor U542 (N_542,N_455,N_274);
nand U543 (N_543,N_314,N_320);
and U544 (N_544,N_432,N_477);
xnor U545 (N_545,In_690,N_200);
nand U546 (N_546,In_277,N_470);
or U547 (N_547,In_566,N_469);
and U548 (N_548,In_37,N_120);
xor U549 (N_549,N_212,N_407);
or U550 (N_550,N_347,N_299);
or U551 (N_551,N_143,N_480);
nor U552 (N_552,In_368,N_436);
nand U553 (N_553,N_420,N_445);
nand U554 (N_554,N_488,N_332);
nand U555 (N_555,N_218,In_275);
nor U556 (N_556,In_489,N_28);
nor U557 (N_557,N_221,In_553);
nor U558 (N_558,N_448,N_449);
and U559 (N_559,N_391,N_185);
nand U560 (N_560,N_368,N_418);
nand U561 (N_561,N_412,N_342);
and U562 (N_562,N_461,N_52);
or U563 (N_563,N_444,N_478);
or U564 (N_564,N_351,N_319);
nand U565 (N_565,In_9,N_322);
nor U566 (N_566,N_381,N_431);
and U567 (N_567,In_86,In_95);
xnor U568 (N_568,N_494,In_596);
and U569 (N_569,N_268,In_51);
or U570 (N_570,N_23,N_410);
or U571 (N_571,N_388,N_433);
or U572 (N_572,N_457,N_44);
or U573 (N_573,N_428,N_298);
nor U574 (N_574,In_29,N_490);
and U575 (N_575,In_460,N_312);
or U576 (N_576,N_426,N_430);
nand U577 (N_577,N_96,In_390);
and U578 (N_578,N_339,N_145);
or U579 (N_579,N_486,N_370);
or U580 (N_580,N_440,In_40);
nor U581 (N_581,In_195,N_483);
nor U582 (N_582,N_463,N_148);
and U583 (N_583,In_567,N_400);
and U584 (N_584,N_127,N_402);
and U585 (N_585,N_350,N_243);
and U586 (N_586,N_429,N_389);
and U587 (N_587,N_427,In_122);
or U588 (N_588,In_361,N_401);
or U589 (N_589,In_722,N_485);
and U590 (N_590,N_354,In_679);
nor U591 (N_591,In_670,In_538);
or U592 (N_592,N_451,In_249);
xor U593 (N_593,N_335,In_12);
and U594 (N_594,In_615,N_182);
and U595 (N_595,N_499,N_479);
nor U596 (N_596,N_452,In_359);
nand U597 (N_597,N_233,N_474);
xnor U598 (N_598,N_434,N_493);
nor U599 (N_599,N_408,N_458);
xnor U600 (N_600,N_558,N_328);
or U601 (N_601,N_405,N_129);
and U602 (N_602,N_583,N_576);
or U603 (N_603,N_548,N_544);
nand U604 (N_604,N_568,N_307);
nor U605 (N_605,N_525,N_570);
nand U606 (N_606,In_186,N_502);
and U607 (N_607,N_553,N_503);
and U608 (N_608,N_487,N_543);
nand U609 (N_609,In_322,N_526);
and U610 (N_610,N_550,N_519);
or U611 (N_611,N_417,N_561);
and U612 (N_612,N_562,In_462);
xnor U613 (N_613,N_508,N_565);
or U614 (N_614,N_595,N_589);
nand U615 (N_615,N_511,N_514);
or U616 (N_616,N_555,N_572);
nor U617 (N_617,N_575,N_557);
nand U618 (N_618,N_422,N_198);
nand U619 (N_619,In_155,N_439);
or U620 (N_620,N_596,N_594);
and U621 (N_621,N_404,N_528);
nor U622 (N_622,N_527,N_425);
or U623 (N_623,N_569,N_598);
xor U624 (N_624,N_573,N_529);
and U625 (N_625,N_229,In_350);
nand U626 (N_626,N_530,N_556);
or U627 (N_627,N_403,N_559);
nor U628 (N_628,N_538,N_540);
or U629 (N_629,N_466,N_523);
nand U630 (N_630,N_554,N_251);
nand U631 (N_631,N_532,N_484);
or U632 (N_632,N_520,N_424);
nor U633 (N_633,N_500,N_551);
nor U634 (N_634,N_146,N_360);
nor U635 (N_635,In_527,N_584);
or U636 (N_636,N_537,N_512);
nand U637 (N_637,N_521,N_411);
or U638 (N_638,N_465,N_593);
or U639 (N_639,N_547,N_599);
or U640 (N_640,N_126,N_588);
or U641 (N_641,N_507,N_515);
or U642 (N_642,N_334,N_546);
and U643 (N_643,N_189,N_542);
and U644 (N_644,N_524,N_513);
or U645 (N_645,N_586,N_491);
nand U646 (N_646,N_579,N_574);
or U647 (N_647,N_369,N_531);
and U648 (N_648,N_481,N_517);
or U649 (N_649,N_535,N_501);
nand U650 (N_650,N_496,N_98);
or U651 (N_651,N_563,N_534);
xnor U652 (N_652,N_581,N_564);
nand U653 (N_653,In_620,N_545);
nor U654 (N_654,N_597,N_472);
and U655 (N_655,In_587,N_164);
xnor U656 (N_656,N_578,N_567);
nand U657 (N_657,N_591,N_560);
nor U658 (N_658,N_552,N_283);
nor U659 (N_659,N_592,N_577);
or U660 (N_660,N_349,N_504);
xor U661 (N_661,N_590,N_571);
nor U662 (N_662,N_495,N_383);
and U663 (N_663,N_536,N_259);
or U664 (N_664,N_223,N_509);
xnor U665 (N_665,N_57,N_587);
or U666 (N_666,In_235,N_522);
nand U667 (N_667,N_549,N_585);
nand U668 (N_668,N_506,N_580);
nor U669 (N_669,N_516,N_505);
nor U670 (N_670,N_539,N_206);
nor U671 (N_671,N_541,N_582);
nand U672 (N_672,N_566,In_595);
nor U673 (N_673,N_533,N_518);
and U674 (N_674,N_510,N_22);
and U675 (N_675,N_546,N_592);
nand U676 (N_676,N_535,N_547);
or U677 (N_677,N_565,N_404);
and U678 (N_678,N_403,N_587);
xnor U679 (N_679,N_496,In_595);
nor U680 (N_680,N_534,N_129);
xor U681 (N_681,N_513,N_546);
and U682 (N_682,N_495,N_505);
nand U683 (N_683,N_500,N_504);
xnor U684 (N_684,N_424,N_541);
nand U685 (N_685,N_411,N_558);
or U686 (N_686,N_543,N_552);
and U687 (N_687,N_540,N_537);
and U688 (N_688,N_562,N_98);
nor U689 (N_689,N_542,N_544);
xor U690 (N_690,N_592,N_349);
xor U691 (N_691,N_512,N_405);
or U692 (N_692,N_504,N_559);
nand U693 (N_693,N_404,N_509);
nand U694 (N_694,N_514,N_500);
or U695 (N_695,N_189,N_508);
nand U696 (N_696,N_564,N_551);
nor U697 (N_697,N_529,N_425);
or U698 (N_698,N_547,N_516);
nand U699 (N_699,N_206,N_531);
nand U700 (N_700,N_638,N_655);
or U701 (N_701,N_663,N_699);
or U702 (N_702,N_680,N_695);
and U703 (N_703,N_600,N_615);
nand U704 (N_704,N_619,N_634);
xnor U705 (N_705,N_647,N_618);
nand U706 (N_706,N_681,N_696);
nand U707 (N_707,N_612,N_661);
nand U708 (N_708,N_668,N_630);
or U709 (N_709,N_694,N_679);
and U710 (N_710,N_617,N_691);
or U711 (N_711,N_689,N_658);
and U712 (N_712,N_651,N_627);
nor U713 (N_713,N_625,N_610);
nor U714 (N_714,N_666,N_664);
nand U715 (N_715,N_646,N_649);
xnor U716 (N_716,N_674,N_698);
or U717 (N_717,N_611,N_603);
or U718 (N_718,N_673,N_653);
and U719 (N_719,N_688,N_693);
nor U720 (N_720,N_670,N_648);
or U721 (N_721,N_684,N_676);
or U722 (N_722,N_609,N_665);
and U723 (N_723,N_687,N_635);
nand U724 (N_724,N_644,N_607);
nand U725 (N_725,N_604,N_685);
and U726 (N_726,N_690,N_629);
or U727 (N_727,N_623,N_643);
and U728 (N_728,N_620,N_652);
and U729 (N_729,N_654,N_669);
or U730 (N_730,N_605,N_650);
and U731 (N_731,N_677,N_683);
and U732 (N_732,N_675,N_660);
or U733 (N_733,N_616,N_667);
or U734 (N_734,N_672,N_640);
nand U735 (N_735,N_613,N_601);
or U736 (N_736,N_657,N_639);
and U737 (N_737,N_622,N_608);
xnor U738 (N_738,N_628,N_606);
nor U739 (N_739,N_642,N_637);
or U740 (N_740,N_686,N_678);
xnor U741 (N_741,N_626,N_682);
and U742 (N_742,N_645,N_662);
xnor U743 (N_743,N_624,N_641);
xor U744 (N_744,N_633,N_631);
or U745 (N_745,N_602,N_632);
nor U746 (N_746,N_692,N_671);
and U747 (N_747,N_697,N_656);
xor U748 (N_748,N_621,N_636);
nor U749 (N_749,N_659,N_614);
or U750 (N_750,N_673,N_686);
nand U751 (N_751,N_649,N_650);
xor U752 (N_752,N_634,N_657);
and U753 (N_753,N_661,N_689);
nor U754 (N_754,N_626,N_629);
nor U755 (N_755,N_618,N_631);
nor U756 (N_756,N_631,N_684);
nor U757 (N_757,N_604,N_637);
or U758 (N_758,N_659,N_692);
xnor U759 (N_759,N_659,N_655);
and U760 (N_760,N_641,N_692);
nor U761 (N_761,N_627,N_656);
or U762 (N_762,N_678,N_689);
xor U763 (N_763,N_659,N_691);
and U764 (N_764,N_687,N_657);
xor U765 (N_765,N_622,N_660);
nor U766 (N_766,N_633,N_636);
or U767 (N_767,N_692,N_685);
nor U768 (N_768,N_606,N_676);
or U769 (N_769,N_634,N_641);
and U770 (N_770,N_612,N_652);
nand U771 (N_771,N_640,N_639);
or U772 (N_772,N_626,N_642);
xor U773 (N_773,N_616,N_626);
or U774 (N_774,N_681,N_691);
and U775 (N_775,N_683,N_644);
or U776 (N_776,N_619,N_653);
or U777 (N_777,N_684,N_697);
xnor U778 (N_778,N_676,N_627);
nand U779 (N_779,N_657,N_673);
or U780 (N_780,N_604,N_672);
or U781 (N_781,N_661,N_672);
or U782 (N_782,N_601,N_607);
and U783 (N_783,N_667,N_658);
xnor U784 (N_784,N_651,N_641);
nor U785 (N_785,N_606,N_699);
or U786 (N_786,N_665,N_638);
nand U787 (N_787,N_612,N_648);
nand U788 (N_788,N_641,N_644);
xor U789 (N_789,N_644,N_671);
or U790 (N_790,N_685,N_676);
and U791 (N_791,N_668,N_611);
nand U792 (N_792,N_672,N_649);
xor U793 (N_793,N_629,N_639);
nor U794 (N_794,N_612,N_620);
nor U795 (N_795,N_686,N_639);
or U796 (N_796,N_663,N_624);
nand U797 (N_797,N_670,N_694);
xor U798 (N_798,N_682,N_618);
or U799 (N_799,N_656,N_692);
nor U800 (N_800,N_725,N_783);
and U801 (N_801,N_723,N_737);
and U802 (N_802,N_796,N_754);
nand U803 (N_803,N_735,N_760);
and U804 (N_804,N_788,N_731);
nor U805 (N_805,N_739,N_752);
nand U806 (N_806,N_706,N_755);
xnor U807 (N_807,N_756,N_718);
nand U808 (N_808,N_779,N_708);
or U809 (N_809,N_734,N_789);
nand U810 (N_810,N_702,N_763);
nand U811 (N_811,N_780,N_709);
nand U812 (N_812,N_743,N_749);
or U813 (N_813,N_728,N_717);
nor U814 (N_814,N_701,N_773);
nor U815 (N_815,N_753,N_765);
nand U816 (N_816,N_757,N_707);
xnor U817 (N_817,N_738,N_766);
and U818 (N_818,N_792,N_774);
or U819 (N_819,N_713,N_730);
and U820 (N_820,N_772,N_726);
or U821 (N_821,N_750,N_724);
and U822 (N_822,N_790,N_732);
nor U823 (N_823,N_744,N_714);
nor U824 (N_824,N_747,N_751);
xor U825 (N_825,N_733,N_741);
nor U826 (N_826,N_715,N_722);
and U827 (N_827,N_721,N_704);
nand U828 (N_828,N_712,N_795);
nand U829 (N_829,N_791,N_775);
nand U830 (N_830,N_711,N_786);
nand U831 (N_831,N_798,N_748);
or U832 (N_832,N_799,N_727);
nor U833 (N_833,N_787,N_793);
nand U834 (N_834,N_742,N_736);
or U835 (N_835,N_758,N_716);
or U836 (N_836,N_777,N_784);
nor U837 (N_837,N_781,N_785);
and U838 (N_838,N_705,N_769);
nand U839 (N_839,N_764,N_778);
nand U840 (N_840,N_782,N_746);
and U841 (N_841,N_771,N_719);
nor U842 (N_842,N_794,N_745);
nand U843 (N_843,N_759,N_729);
xnor U844 (N_844,N_776,N_700);
and U845 (N_845,N_761,N_710);
and U846 (N_846,N_770,N_720);
xnor U847 (N_847,N_768,N_703);
nor U848 (N_848,N_767,N_797);
and U849 (N_849,N_740,N_762);
xnor U850 (N_850,N_707,N_793);
or U851 (N_851,N_782,N_703);
or U852 (N_852,N_769,N_789);
xnor U853 (N_853,N_764,N_707);
nor U854 (N_854,N_728,N_734);
and U855 (N_855,N_711,N_753);
nand U856 (N_856,N_731,N_774);
and U857 (N_857,N_729,N_730);
nor U858 (N_858,N_786,N_700);
nor U859 (N_859,N_724,N_776);
xor U860 (N_860,N_704,N_765);
or U861 (N_861,N_793,N_743);
nor U862 (N_862,N_735,N_764);
and U863 (N_863,N_736,N_715);
nor U864 (N_864,N_704,N_768);
nand U865 (N_865,N_727,N_791);
nand U866 (N_866,N_726,N_794);
nand U867 (N_867,N_774,N_709);
nor U868 (N_868,N_777,N_773);
or U869 (N_869,N_767,N_710);
or U870 (N_870,N_736,N_754);
nor U871 (N_871,N_757,N_763);
or U872 (N_872,N_721,N_720);
and U873 (N_873,N_766,N_755);
or U874 (N_874,N_700,N_701);
nor U875 (N_875,N_731,N_790);
nor U876 (N_876,N_700,N_737);
nor U877 (N_877,N_795,N_722);
and U878 (N_878,N_752,N_771);
or U879 (N_879,N_783,N_743);
nor U880 (N_880,N_708,N_762);
nand U881 (N_881,N_791,N_747);
or U882 (N_882,N_740,N_703);
and U883 (N_883,N_790,N_725);
nor U884 (N_884,N_704,N_726);
or U885 (N_885,N_763,N_747);
nand U886 (N_886,N_782,N_744);
and U887 (N_887,N_758,N_774);
or U888 (N_888,N_700,N_703);
nand U889 (N_889,N_703,N_714);
nand U890 (N_890,N_728,N_762);
or U891 (N_891,N_781,N_730);
or U892 (N_892,N_741,N_731);
or U893 (N_893,N_751,N_711);
and U894 (N_894,N_739,N_744);
nand U895 (N_895,N_721,N_711);
and U896 (N_896,N_731,N_799);
and U897 (N_897,N_787,N_701);
or U898 (N_898,N_772,N_780);
or U899 (N_899,N_798,N_753);
and U900 (N_900,N_849,N_888);
nor U901 (N_901,N_880,N_829);
and U902 (N_902,N_845,N_832);
and U903 (N_903,N_864,N_808);
and U904 (N_904,N_852,N_815);
and U905 (N_905,N_813,N_873);
nor U906 (N_906,N_836,N_817);
or U907 (N_907,N_853,N_844);
nor U908 (N_908,N_827,N_893);
or U909 (N_909,N_865,N_820);
and U910 (N_910,N_833,N_851);
and U911 (N_911,N_822,N_874);
nand U912 (N_912,N_859,N_802);
or U913 (N_913,N_841,N_805);
or U914 (N_914,N_892,N_819);
nor U915 (N_915,N_838,N_830);
and U916 (N_916,N_810,N_826);
nand U917 (N_917,N_870,N_898);
and U918 (N_918,N_882,N_894);
nand U919 (N_919,N_890,N_828);
nand U920 (N_920,N_866,N_884);
and U921 (N_921,N_855,N_809);
nor U922 (N_922,N_839,N_856);
and U923 (N_923,N_848,N_877);
and U924 (N_924,N_834,N_886);
and U925 (N_925,N_842,N_812);
and U926 (N_926,N_897,N_850);
and U927 (N_927,N_895,N_879);
or U928 (N_928,N_825,N_862);
or U929 (N_929,N_814,N_869);
or U930 (N_930,N_867,N_860);
nand U931 (N_931,N_891,N_875);
and U932 (N_932,N_824,N_847);
or U933 (N_933,N_887,N_821);
or U934 (N_934,N_885,N_868);
nand U935 (N_935,N_846,N_818);
or U936 (N_936,N_889,N_816);
xor U937 (N_937,N_823,N_863);
and U938 (N_938,N_800,N_871);
or U939 (N_939,N_831,N_872);
nand U940 (N_940,N_843,N_835);
or U941 (N_941,N_801,N_857);
xnor U942 (N_942,N_881,N_807);
xor U943 (N_943,N_861,N_811);
or U944 (N_944,N_858,N_876);
and U945 (N_945,N_806,N_837);
xnor U946 (N_946,N_854,N_883);
nand U947 (N_947,N_878,N_804);
and U948 (N_948,N_803,N_899);
xnor U949 (N_949,N_840,N_896);
nand U950 (N_950,N_849,N_868);
or U951 (N_951,N_876,N_859);
nor U952 (N_952,N_847,N_898);
nand U953 (N_953,N_843,N_850);
or U954 (N_954,N_819,N_809);
nor U955 (N_955,N_860,N_861);
or U956 (N_956,N_826,N_845);
or U957 (N_957,N_891,N_898);
and U958 (N_958,N_814,N_834);
or U959 (N_959,N_898,N_864);
nand U960 (N_960,N_878,N_821);
nand U961 (N_961,N_897,N_843);
nand U962 (N_962,N_882,N_897);
and U963 (N_963,N_875,N_826);
nor U964 (N_964,N_845,N_893);
or U965 (N_965,N_877,N_891);
nor U966 (N_966,N_826,N_809);
nor U967 (N_967,N_847,N_897);
and U968 (N_968,N_868,N_850);
and U969 (N_969,N_819,N_894);
nand U970 (N_970,N_865,N_896);
or U971 (N_971,N_836,N_888);
nor U972 (N_972,N_875,N_856);
nor U973 (N_973,N_839,N_855);
xor U974 (N_974,N_822,N_834);
or U975 (N_975,N_846,N_826);
or U976 (N_976,N_895,N_817);
nand U977 (N_977,N_843,N_896);
xor U978 (N_978,N_838,N_865);
xor U979 (N_979,N_889,N_895);
nand U980 (N_980,N_821,N_851);
nor U981 (N_981,N_880,N_823);
and U982 (N_982,N_831,N_840);
nand U983 (N_983,N_805,N_822);
or U984 (N_984,N_877,N_859);
or U985 (N_985,N_861,N_804);
or U986 (N_986,N_814,N_896);
xor U987 (N_987,N_814,N_839);
or U988 (N_988,N_828,N_878);
or U989 (N_989,N_803,N_842);
nand U990 (N_990,N_855,N_823);
and U991 (N_991,N_829,N_855);
nand U992 (N_992,N_872,N_850);
nor U993 (N_993,N_865,N_834);
and U994 (N_994,N_838,N_867);
or U995 (N_995,N_870,N_820);
or U996 (N_996,N_853,N_835);
nand U997 (N_997,N_868,N_896);
and U998 (N_998,N_854,N_846);
xor U999 (N_999,N_870,N_810);
xnor U1000 (N_1000,N_994,N_936);
nand U1001 (N_1001,N_929,N_922);
nor U1002 (N_1002,N_972,N_966);
or U1003 (N_1003,N_900,N_934);
nor U1004 (N_1004,N_909,N_937);
nand U1005 (N_1005,N_950,N_968);
and U1006 (N_1006,N_982,N_945);
nor U1007 (N_1007,N_985,N_960);
xor U1008 (N_1008,N_998,N_919);
nand U1009 (N_1009,N_925,N_959);
and U1010 (N_1010,N_992,N_974);
nand U1011 (N_1011,N_970,N_944);
nand U1012 (N_1012,N_902,N_978);
xor U1013 (N_1013,N_951,N_952);
nor U1014 (N_1014,N_935,N_933);
or U1015 (N_1015,N_958,N_903);
and U1016 (N_1016,N_942,N_918);
nand U1017 (N_1017,N_956,N_997);
nand U1018 (N_1018,N_957,N_986);
nand U1019 (N_1019,N_916,N_914);
xor U1020 (N_1020,N_908,N_989);
nand U1021 (N_1021,N_948,N_995);
or U1022 (N_1022,N_977,N_955);
or U1023 (N_1023,N_975,N_904);
or U1024 (N_1024,N_973,N_947);
or U1025 (N_1025,N_910,N_984);
nor U1026 (N_1026,N_917,N_930);
or U1027 (N_1027,N_939,N_928);
nand U1028 (N_1028,N_940,N_932);
xor U1029 (N_1029,N_980,N_954);
and U1030 (N_1030,N_938,N_953);
and U1031 (N_1031,N_924,N_907);
nand U1032 (N_1032,N_964,N_971);
and U1033 (N_1033,N_979,N_927);
nand U1034 (N_1034,N_961,N_926);
nor U1035 (N_1035,N_949,N_931);
or U1036 (N_1036,N_983,N_991);
and U1037 (N_1037,N_906,N_988);
nand U1038 (N_1038,N_921,N_923);
or U1039 (N_1039,N_962,N_901);
and U1040 (N_1040,N_987,N_993);
and U1041 (N_1041,N_911,N_999);
and U1042 (N_1042,N_963,N_981);
nor U1043 (N_1043,N_912,N_905);
or U1044 (N_1044,N_920,N_913);
or U1045 (N_1045,N_969,N_976);
nor U1046 (N_1046,N_915,N_965);
and U1047 (N_1047,N_996,N_967);
nor U1048 (N_1048,N_946,N_990);
nor U1049 (N_1049,N_941,N_943);
nor U1050 (N_1050,N_984,N_953);
nor U1051 (N_1051,N_936,N_907);
or U1052 (N_1052,N_971,N_952);
and U1053 (N_1053,N_973,N_946);
nor U1054 (N_1054,N_936,N_960);
nor U1055 (N_1055,N_982,N_991);
xor U1056 (N_1056,N_917,N_985);
and U1057 (N_1057,N_993,N_901);
nor U1058 (N_1058,N_937,N_932);
or U1059 (N_1059,N_950,N_946);
or U1060 (N_1060,N_965,N_964);
nor U1061 (N_1061,N_974,N_906);
xor U1062 (N_1062,N_978,N_910);
nand U1063 (N_1063,N_927,N_998);
nor U1064 (N_1064,N_960,N_973);
and U1065 (N_1065,N_929,N_912);
nand U1066 (N_1066,N_906,N_992);
nor U1067 (N_1067,N_908,N_955);
xor U1068 (N_1068,N_958,N_915);
nor U1069 (N_1069,N_991,N_935);
nor U1070 (N_1070,N_954,N_979);
nor U1071 (N_1071,N_969,N_925);
or U1072 (N_1072,N_919,N_936);
or U1073 (N_1073,N_958,N_939);
nand U1074 (N_1074,N_977,N_989);
nor U1075 (N_1075,N_990,N_906);
nand U1076 (N_1076,N_991,N_959);
nor U1077 (N_1077,N_981,N_984);
or U1078 (N_1078,N_988,N_939);
xnor U1079 (N_1079,N_977,N_947);
and U1080 (N_1080,N_999,N_950);
nand U1081 (N_1081,N_933,N_902);
nand U1082 (N_1082,N_909,N_991);
and U1083 (N_1083,N_906,N_920);
nand U1084 (N_1084,N_964,N_984);
nand U1085 (N_1085,N_907,N_990);
or U1086 (N_1086,N_929,N_948);
nand U1087 (N_1087,N_901,N_946);
and U1088 (N_1088,N_918,N_935);
nand U1089 (N_1089,N_935,N_968);
xor U1090 (N_1090,N_947,N_961);
nor U1091 (N_1091,N_958,N_931);
and U1092 (N_1092,N_931,N_928);
or U1093 (N_1093,N_962,N_961);
nand U1094 (N_1094,N_957,N_941);
or U1095 (N_1095,N_917,N_997);
nor U1096 (N_1096,N_966,N_959);
and U1097 (N_1097,N_990,N_926);
nand U1098 (N_1098,N_993,N_964);
and U1099 (N_1099,N_938,N_920);
nor U1100 (N_1100,N_1039,N_1061);
nand U1101 (N_1101,N_1037,N_1058);
nor U1102 (N_1102,N_1009,N_1019);
nor U1103 (N_1103,N_1057,N_1026);
nor U1104 (N_1104,N_1092,N_1064);
nand U1105 (N_1105,N_1051,N_1006);
nand U1106 (N_1106,N_1073,N_1022);
and U1107 (N_1107,N_1046,N_1029);
or U1108 (N_1108,N_1089,N_1030);
nor U1109 (N_1109,N_1094,N_1042);
xnor U1110 (N_1110,N_1093,N_1040);
and U1111 (N_1111,N_1084,N_1070);
nand U1112 (N_1112,N_1025,N_1027);
and U1113 (N_1113,N_1033,N_1008);
and U1114 (N_1114,N_1097,N_1004);
nand U1115 (N_1115,N_1000,N_1048);
nand U1116 (N_1116,N_1060,N_1062);
nor U1117 (N_1117,N_1032,N_1053);
and U1118 (N_1118,N_1077,N_1079);
and U1119 (N_1119,N_1071,N_1083);
and U1120 (N_1120,N_1028,N_1082);
nor U1121 (N_1121,N_1091,N_1013);
and U1122 (N_1122,N_1031,N_1095);
and U1123 (N_1123,N_1075,N_1016);
xor U1124 (N_1124,N_1047,N_1081);
and U1125 (N_1125,N_1076,N_1018);
or U1126 (N_1126,N_1087,N_1056);
or U1127 (N_1127,N_1038,N_1036);
and U1128 (N_1128,N_1069,N_1014);
and U1129 (N_1129,N_1043,N_1067);
nand U1130 (N_1130,N_1020,N_1050);
or U1131 (N_1131,N_1049,N_1068);
nand U1132 (N_1132,N_1011,N_1072);
nand U1133 (N_1133,N_1044,N_1096);
or U1134 (N_1134,N_1005,N_1088);
or U1135 (N_1135,N_1085,N_1024);
xor U1136 (N_1136,N_1041,N_1066);
nand U1137 (N_1137,N_1099,N_1059);
or U1138 (N_1138,N_1098,N_1002);
nand U1139 (N_1139,N_1054,N_1021);
or U1140 (N_1140,N_1074,N_1063);
and U1141 (N_1141,N_1035,N_1015);
and U1142 (N_1142,N_1090,N_1023);
or U1143 (N_1143,N_1017,N_1010);
nand U1144 (N_1144,N_1080,N_1001);
nor U1145 (N_1145,N_1012,N_1086);
xor U1146 (N_1146,N_1003,N_1078);
nor U1147 (N_1147,N_1045,N_1052);
nor U1148 (N_1148,N_1065,N_1055);
xnor U1149 (N_1149,N_1034,N_1007);
and U1150 (N_1150,N_1023,N_1070);
nand U1151 (N_1151,N_1043,N_1044);
or U1152 (N_1152,N_1043,N_1078);
and U1153 (N_1153,N_1074,N_1043);
nand U1154 (N_1154,N_1022,N_1001);
and U1155 (N_1155,N_1054,N_1031);
or U1156 (N_1156,N_1084,N_1019);
and U1157 (N_1157,N_1059,N_1079);
nor U1158 (N_1158,N_1035,N_1048);
nor U1159 (N_1159,N_1041,N_1035);
and U1160 (N_1160,N_1010,N_1005);
and U1161 (N_1161,N_1055,N_1081);
nor U1162 (N_1162,N_1000,N_1042);
and U1163 (N_1163,N_1072,N_1001);
nor U1164 (N_1164,N_1025,N_1020);
and U1165 (N_1165,N_1072,N_1084);
or U1166 (N_1166,N_1077,N_1087);
xnor U1167 (N_1167,N_1085,N_1017);
and U1168 (N_1168,N_1032,N_1025);
nand U1169 (N_1169,N_1078,N_1041);
nor U1170 (N_1170,N_1060,N_1055);
nor U1171 (N_1171,N_1022,N_1093);
or U1172 (N_1172,N_1005,N_1047);
xor U1173 (N_1173,N_1060,N_1097);
nand U1174 (N_1174,N_1082,N_1017);
or U1175 (N_1175,N_1080,N_1002);
nand U1176 (N_1176,N_1021,N_1096);
nor U1177 (N_1177,N_1048,N_1084);
and U1178 (N_1178,N_1047,N_1035);
nor U1179 (N_1179,N_1003,N_1055);
nor U1180 (N_1180,N_1026,N_1023);
or U1181 (N_1181,N_1021,N_1039);
nor U1182 (N_1182,N_1075,N_1064);
nand U1183 (N_1183,N_1070,N_1054);
nand U1184 (N_1184,N_1006,N_1071);
nor U1185 (N_1185,N_1058,N_1066);
and U1186 (N_1186,N_1002,N_1069);
nand U1187 (N_1187,N_1089,N_1083);
nand U1188 (N_1188,N_1006,N_1057);
nor U1189 (N_1189,N_1038,N_1076);
nand U1190 (N_1190,N_1062,N_1086);
or U1191 (N_1191,N_1027,N_1017);
nor U1192 (N_1192,N_1036,N_1030);
or U1193 (N_1193,N_1078,N_1069);
nor U1194 (N_1194,N_1096,N_1045);
or U1195 (N_1195,N_1003,N_1084);
or U1196 (N_1196,N_1008,N_1039);
or U1197 (N_1197,N_1046,N_1052);
nand U1198 (N_1198,N_1044,N_1006);
nand U1199 (N_1199,N_1090,N_1020);
nand U1200 (N_1200,N_1126,N_1146);
nand U1201 (N_1201,N_1156,N_1187);
or U1202 (N_1202,N_1193,N_1135);
nor U1203 (N_1203,N_1133,N_1117);
and U1204 (N_1204,N_1119,N_1141);
or U1205 (N_1205,N_1194,N_1132);
nand U1206 (N_1206,N_1198,N_1170);
nand U1207 (N_1207,N_1197,N_1104);
and U1208 (N_1208,N_1174,N_1151);
and U1209 (N_1209,N_1157,N_1144);
nand U1210 (N_1210,N_1114,N_1162);
xor U1211 (N_1211,N_1159,N_1166);
or U1212 (N_1212,N_1100,N_1158);
nand U1213 (N_1213,N_1161,N_1122);
or U1214 (N_1214,N_1188,N_1185);
nor U1215 (N_1215,N_1189,N_1148);
xnor U1216 (N_1216,N_1129,N_1186);
and U1217 (N_1217,N_1150,N_1113);
nor U1218 (N_1218,N_1123,N_1149);
or U1219 (N_1219,N_1178,N_1105);
nand U1220 (N_1220,N_1139,N_1102);
or U1221 (N_1221,N_1152,N_1168);
and U1222 (N_1222,N_1121,N_1101);
or U1223 (N_1223,N_1167,N_1134);
nor U1224 (N_1224,N_1191,N_1180);
nor U1225 (N_1225,N_1183,N_1112);
and U1226 (N_1226,N_1145,N_1160);
nor U1227 (N_1227,N_1165,N_1111);
or U1228 (N_1228,N_1118,N_1199);
and U1229 (N_1229,N_1173,N_1130);
nand U1230 (N_1230,N_1154,N_1155);
or U1231 (N_1231,N_1136,N_1147);
or U1232 (N_1232,N_1142,N_1140);
and U1233 (N_1233,N_1106,N_1110);
nand U1234 (N_1234,N_1163,N_1196);
nor U1235 (N_1235,N_1175,N_1120);
or U1236 (N_1236,N_1177,N_1128);
nand U1237 (N_1237,N_1107,N_1109);
and U1238 (N_1238,N_1131,N_1137);
or U1239 (N_1239,N_1116,N_1182);
and U1240 (N_1240,N_1195,N_1184);
nand U1241 (N_1241,N_1190,N_1127);
or U1242 (N_1242,N_1138,N_1176);
nor U1243 (N_1243,N_1125,N_1192);
and U1244 (N_1244,N_1172,N_1164);
and U1245 (N_1245,N_1179,N_1169);
xor U1246 (N_1246,N_1153,N_1124);
or U1247 (N_1247,N_1103,N_1143);
or U1248 (N_1248,N_1181,N_1171);
and U1249 (N_1249,N_1115,N_1108);
and U1250 (N_1250,N_1127,N_1146);
nand U1251 (N_1251,N_1189,N_1110);
or U1252 (N_1252,N_1148,N_1136);
and U1253 (N_1253,N_1152,N_1120);
xnor U1254 (N_1254,N_1127,N_1131);
or U1255 (N_1255,N_1188,N_1107);
xor U1256 (N_1256,N_1179,N_1124);
or U1257 (N_1257,N_1141,N_1131);
nor U1258 (N_1258,N_1109,N_1120);
xor U1259 (N_1259,N_1182,N_1198);
nand U1260 (N_1260,N_1110,N_1129);
and U1261 (N_1261,N_1119,N_1123);
nand U1262 (N_1262,N_1135,N_1183);
and U1263 (N_1263,N_1130,N_1125);
or U1264 (N_1264,N_1128,N_1198);
or U1265 (N_1265,N_1153,N_1196);
nor U1266 (N_1266,N_1126,N_1156);
or U1267 (N_1267,N_1157,N_1197);
xor U1268 (N_1268,N_1187,N_1102);
and U1269 (N_1269,N_1193,N_1198);
or U1270 (N_1270,N_1103,N_1186);
nor U1271 (N_1271,N_1172,N_1121);
nor U1272 (N_1272,N_1150,N_1198);
nor U1273 (N_1273,N_1133,N_1160);
nand U1274 (N_1274,N_1170,N_1167);
xor U1275 (N_1275,N_1101,N_1175);
nand U1276 (N_1276,N_1106,N_1142);
nor U1277 (N_1277,N_1126,N_1108);
nand U1278 (N_1278,N_1197,N_1119);
nor U1279 (N_1279,N_1144,N_1141);
nand U1280 (N_1280,N_1177,N_1111);
or U1281 (N_1281,N_1140,N_1183);
or U1282 (N_1282,N_1129,N_1104);
xnor U1283 (N_1283,N_1144,N_1182);
and U1284 (N_1284,N_1168,N_1103);
xor U1285 (N_1285,N_1142,N_1181);
or U1286 (N_1286,N_1194,N_1141);
nor U1287 (N_1287,N_1159,N_1176);
or U1288 (N_1288,N_1167,N_1166);
and U1289 (N_1289,N_1176,N_1157);
or U1290 (N_1290,N_1152,N_1124);
xnor U1291 (N_1291,N_1100,N_1162);
xnor U1292 (N_1292,N_1145,N_1140);
or U1293 (N_1293,N_1144,N_1129);
nand U1294 (N_1294,N_1150,N_1151);
nand U1295 (N_1295,N_1199,N_1154);
nand U1296 (N_1296,N_1184,N_1177);
nor U1297 (N_1297,N_1188,N_1118);
and U1298 (N_1298,N_1158,N_1173);
nor U1299 (N_1299,N_1120,N_1198);
and U1300 (N_1300,N_1214,N_1286);
nand U1301 (N_1301,N_1236,N_1243);
or U1302 (N_1302,N_1226,N_1235);
or U1303 (N_1303,N_1247,N_1292);
or U1304 (N_1304,N_1248,N_1253);
and U1305 (N_1305,N_1218,N_1205);
nand U1306 (N_1306,N_1216,N_1203);
nand U1307 (N_1307,N_1211,N_1277);
and U1308 (N_1308,N_1266,N_1239);
nand U1309 (N_1309,N_1240,N_1227);
or U1310 (N_1310,N_1228,N_1260);
nand U1311 (N_1311,N_1244,N_1206);
nand U1312 (N_1312,N_1219,N_1231);
and U1313 (N_1313,N_1246,N_1252);
nor U1314 (N_1314,N_1281,N_1200);
or U1315 (N_1315,N_1285,N_1215);
or U1316 (N_1316,N_1262,N_1233);
nand U1317 (N_1317,N_1249,N_1224);
and U1318 (N_1318,N_1234,N_1256);
nand U1319 (N_1319,N_1272,N_1270);
or U1320 (N_1320,N_1297,N_1221);
or U1321 (N_1321,N_1288,N_1222);
nand U1322 (N_1322,N_1251,N_1230);
and U1323 (N_1323,N_1202,N_1282);
or U1324 (N_1324,N_1237,N_1264);
nor U1325 (N_1325,N_1254,N_1293);
or U1326 (N_1326,N_1268,N_1269);
and U1327 (N_1327,N_1294,N_1275);
and U1328 (N_1328,N_1279,N_1242);
nand U1329 (N_1329,N_1287,N_1263);
xnor U1330 (N_1330,N_1290,N_1241);
or U1331 (N_1331,N_1232,N_1208);
and U1332 (N_1332,N_1283,N_1229);
nor U1333 (N_1333,N_1207,N_1265);
or U1334 (N_1334,N_1299,N_1276);
xnor U1335 (N_1335,N_1250,N_1238);
nor U1336 (N_1336,N_1217,N_1271);
nand U1337 (N_1337,N_1295,N_1298);
nor U1338 (N_1338,N_1212,N_1225);
nand U1339 (N_1339,N_1296,N_1261);
nor U1340 (N_1340,N_1273,N_1201);
nand U1341 (N_1341,N_1291,N_1223);
or U1342 (N_1342,N_1267,N_1257);
nand U1343 (N_1343,N_1280,N_1289);
nand U1344 (N_1344,N_1210,N_1204);
nor U1345 (N_1345,N_1209,N_1284);
and U1346 (N_1346,N_1259,N_1274);
and U1347 (N_1347,N_1220,N_1245);
nand U1348 (N_1348,N_1258,N_1255);
nand U1349 (N_1349,N_1213,N_1278);
nand U1350 (N_1350,N_1230,N_1247);
nand U1351 (N_1351,N_1256,N_1238);
nand U1352 (N_1352,N_1226,N_1295);
nor U1353 (N_1353,N_1287,N_1220);
and U1354 (N_1354,N_1292,N_1269);
nor U1355 (N_1355,N_1265,N_1205);
nor U1356 (N_1356,N_1261,N_1267);
and U1357 (N_1357,N_1249,N_1257);
nor U1358 (N_1358,N_1270,N_1200);
nand U1359 (N_1359,N_1207,N_1242);
nand U1360 (N_1360,N_1288,N_1207);
nand U1361 (N_1361,N_1210,N_1223);
and U1362 (N_1362,N_1279,N_1218);
nand U1363 (N_1363,N_1238,N_1295);
or U1364 (N_1364,N_1264,N_1279);
and U1365 (N_1365,N_1243,N_1245);
nand U1366 (N_1366,N_1215,N_1271);
or U1367 (N_1367,N_1213,N_1226);
or U1368 (N_1368,N_1201,N_1229);
or U1369 (N_1369,N_1204,N_1271);
nand U1370 (N_1370,N_1236,N_1269);
or U1371 (N_1371,N_1297,N_1220);
nand U1372 (N_1372,N_1224,N_1290);
nand U1373 (N_1373,N_1263,N_1222);
nand U1374 (N_1374,N_1288,N_1227);
nand U1375 (N_1375,N_1259,N_1246);
and U1376 (N_1376,N_1260,N_1204);
or U1377 (N_1377,N_1281,N_1293);
or U1378 (N_1378,N_1242,N_1209);
and U1379 (N_1379,N_1250,N_1242);
nand U1380 (N_1380,N_1274,N_1247);
and U1381 (N_1381,N_1293,N_1268);
nor U1382 (N_1382,N_1293,N_1275);
or U1383 (N_1383,N_1285,N_1290);
nand U1384 (N_1384,N_1281,N_1267);
nor U1385 (N_1385,N_1291,N_1219);
or U1386 (N_1386,N_1208,N_1263);
and U1387 (N_1387,N_1298,N_1259);
nor U1388 (N_1388,N_1230,N_1200);
nor U1389 (N_1389,N_1239,N_1208);
or U1390 (N_1390,N_1266,N_1254);
nand U1391 (N_1391,N_1239,N_1298);
or U1392 (N_1392,N_1236,N_1298);
nand U1393 (N_1393,N_1276,N_1216);
nor U1394 (N_1394,N_1282,N_1247);
and U1395 (N_1395,N_1259,N_1221);
nand U1396 (N_1396,N_1286,N_1245);
nand U1397 (N_1397,N_1290,N_1255);
nor U1398 (N_1398,N_1207,N_1211);
and U1399 (N_1399,N_1280,N_1259);
and U1400 (N_1400,N_1317,N_1320);
and U1401 (N_1401,N_1329,N_1341);
xnor U1402 (N_1402,N_1308,N_1309);
nand U1403 (N_1403,N_1374,N_1399);
xor U1404 (N_1404,N_1378,N_1377);
nand U1405 (N_1405,N_1385,N_1393);
nand U1406 (N_1406,N_1390,N_1383);
and U1407 (N_1407,N_1396,N_1340);
nor U1408 (N_1408,N_1369,N_1382);
nor U1409 (N_1409,N_1314,N_1310);
or U1410 (N_1410,N_1349,N_1306);
and U1411 (N_1411,N_1386,N_1331);
nor U1412 (N_1412,N_1334,N_1350);
nor U1413 (N_1413,N_1361,N_1343);
and U1414 (N_1414,N_1321,N_1397);
xnor U1415 (N_1415,N_1328,N_1357);
or U1416 (N_1416,N_1381,N_1379);
and U1417 (N_1417,N_1359,N_1388);
and U1418 (N_1418,N_1365,N_1366);
nand U1419 (N_1419,N_1363,N_1394);
and U1420 (N_1420,N_1364,N_1344);
nand U1421 (N_1421,N_1324,N_1318);
nor U1422 (N_1422,N_1387,N_1323);
nor U1423 (N_1423,N_1351,N_1304);
and U1424 (N_1424,N_1362,N_1395);
xor U1425 (N_1425,N_1305,N_1337);
nor U1426 (N_1426,N_1335,N_1356);
or U1427 (N_1427,N_1333,N_1392);
nand U1428 (N_1428,N_1313,N_1342);
nand U1429 (N_1429,N_1371,N_1376);
xnor U1430 (N_1430,N_1345,N_1322);
or U1431 (N_1431,N_1384,N_1301);
and U1432 (N_1432,N_1311,N_1360);
and U1433 (N_1433,N_1368,N_1302);
nand U1434 (N_1434,N_1315,N_1316);
and U1435 (N_1435,N_1319,N_1332);
nand U1436 (N_1436,N_1338,N_1336);
nor U1437 (N_1437,N_1339,N_1372);
and U1438 (N_1438,N_1312,N_1367);
nor U1439 (N_1439,N_1352,N_1355);
or U1440 (N_1440,N_1303,N_1300);
xor U1441 (N_1441,N_1326,N_1370);
or U1442 (N_1442,N_1330,N_1373);
xnor U1443 (N_1443,N_1346,N_1398);
and U1444 (N_1444,N_1375,N_1353);
and U1445 (N_1445,N_1391,N_1389);
and U1446 (N_1446,N_1307,N_1380);
xnor U1447 (N_1447,N_1327,N_1325);
and U1448 (N_1448,N_1348,N_1354);
nand U1449 (N_1449,N_1347,N_1358);
and U1450 (N_1450,N_1311,N_1335);
nor U1451 (N_1451,N_1383,N_1311);
nand U1452 (N_1452,N_1381,N_1370);
and U1453 (N_1453,N_1305,N_1367);
nor U1454 (N_1454,N_1331,N_1318);
and U1455 (N_1455,N_1367,N_1369);
or U1456 (N_1456,N_1362,N_1373);
xnor U1457 (N_1457,N_1378,N_1346);
nand U1458 (N_1458,N_1331,N_1302);
and U1459 (N_1459,N_1323,N_1351);
nand U1460 (N_1460,N_1398,N_1337);
nand U1461 (N_1461,N_1302,N_1379);
and U1462 (N_1462,N_1389,N_1353);
nor U1463 (N_1463,N_1314,N_1327);
or U1464 (N_1464,N_1342,N_1366);
nand U1465 (N_1465,N_1305,N_1393);
nor U1466 (N_1466,N_1373,N_1389);
xnor U1467 (N_1467,N_1332,N_1352);
or U1468 (N_1468,N_1316,N_1374);
or U1469 (N_1469,N_1305,N_1399);
nor U1470 (N_1470,N_1328,N_1337);
and U1471 (N_1471,N_1392,N_1311);
and U1472 (N_1472,N_1338,N_1362);
nor U1473 (N_1473,N_1351,N_1380);
or U1474 (N_1474,N_1310,N_1393);
nand U1475 (N_1475,N_1375,N_1360);
nor U1476 (N_1476,N_1307,N_1346);
nor U1477 (N_1477,N_1370,N_1399);
or U1478 (N_1478,N_1316,N_1331);
or U1479 (N_1479,N_1369,N_1326);
and U1480 (N_1480,N_1301,N_1307);
and U1481 (N_1481,N_1352,N_1342);
nand U1482 (N_1482,N_1308,N_1387);
nand U1483 (N_1483,N_1375,N_1351);
nor U1484 (N_1484,N_1373,N_1325);
or U1485 (N_1485,N_1356,N_1348);
or U1486 (N_1486,N_1382,N_1388);
nand U1487 (N_1487,N_1316,N_1371);
nor U1488 (N_1488,N_1347,N_1376);
nand U1489 (N_1489,N_1335,N_1312);
or U1490 (N_1490,N_1315,N_1320);
nor U1491 (N_1491,N_1376,N_1342);
nand U1492 (N_1492,N_1347,N_1324);
and U1493 (N_1493,N_1326,N_1392);
or U1494 (N_1494,N_1390,N_1377);
or U1495 (N_1495,N_1303,N_1320);
and U1496 (N_1496,N_1372,N_1378);
nor U1497 (N_1497,N_1373,N_1326);
xnor U1498 (N_1498,N_1389,N_1345);
or U1499 (N_1499,N_1313,N_1380);
nor U1500 (N_1500,N_1473,N_1470);
nor U1501 (N_1501,N_1431,N_1486);
nand U1502 (N_1502,N_1409,N_1451);
and U1503 (N_1503,N_1414,N_1460);
or U1504 (N_1504,N_1436,N_1475);
and U1505 (N_1505,N_1477,N_1405);
xor U1506 (N_1506,N_1491,N_1472);
or U1507 (N_1507,N_1498,N_1487);
or U1508 (N_1508,N_1441,N_1427);
or U1509 (N_1509,N_1439,N_1484);
or U1510 (N_1510,N_1417,N_1406);
and U1511 (N_1511,N_1463,N_1465);
nor U1512 (N_1512,N_1488,N_1404);
or U1513 (N_1513,N_1403,N_1420);
nor U1514 (N_1514,N_1426,N_1411);
or U1515 (N_1515,N_1480,N_1462);
and U1516 (N_1516,N_1494,N_1458);
or U1517 (N_1517,N_1430,N_1453);
nand U1518 (N_1518,N_1464,N_1402);
or U1519 (N_1519,N_1459,N_1482);
or U1520 (N_1520,N_1432,N_1449);
nand U1521 (N_1521,N_1401,N_1428);
and U1522 (N_1522,N_1440,N_1483);
and U1523 (N_1523,N_1442,N_1450);
and U1524 (N_1524,N_1433,N_1461);
nor U1525 (N_1525,N_1478,N_1457);
nor U1526 (N_1526,N_1421,N_1400);
or U1527 (N_1527,N_1466,N_1467);
or U1528 (N_1528,N_1444,N_1425);
nand U1529 (N_1529,N_1413,N_1471);
or U1530 (N_1530,N_1438,N_1410);
and U1531 (N_1531,N_1423,N_1485);
and U1532 (N_1532,N_1474,N_1481);
nand U1533 (N_1533,N_1424,N_1407);
nand U1534 (N_1534,N_1452,N_1476);
nand U1535 (N_1535,N_1499,N_1448);
and U1536 (N_1536,N_1479,N_1497);
nor U1537 (N_1537,N_1446,N_1415);
nor U1538 (N_1538,N_1493,N_1422);
or U1539 (N_1539,N_1437,N_1416);
and U1540 (N_1540,N_1469,N_1408);
xor U1541 (N_1541,N_1456,N_1447);
nand U1542 (N_1542,N_1412,N_1454);
nand U1543 (N_1543,N_1468,N_1434);
nand U1544 (N_1544,N_1435,N_1489);
xor U1545 (N_1545,N_1496,N_1492);
nor U1546 (N_1546,N_1445,N_1490);
nand U1547 (N_1547,N_1418,N_1419);
nand U1548 (N_1548,N_1443,N_1495);
nand U1549 (N_1549,N_1455,N_1429);
and U1550 (N_1550,N_1489,N_1417);
or U1551 (N_1551,N_1430,N_1438);
nor U1552 (N_1552,N_1489,N_1411);
nor U1553 (N_1553,N_1450,N_1402);
nand U1554 (N_1554,N_1416,N_1448);
nand U1555 (N_1555,N_1417,N_1415);
or U1556 (N_1556,N_1479,N_1445);
or U1557 (N_1557,N_1403,N_1484);
nand U1558 (N_1558,N_1422,N_1419);
or U1559 (N_1559,N_1479,N_1410);
nor U1560 (N_1560,N_1487,N_1467);
and U1561 (N_1561,N_1461,N_1474);
and U1562 (N_1562,N_1402,N_1485);
and U1563 (N_1563,N_1450,N_1435);
nand U1564 (N_1564,N_1428,N_1495);
or U1565 (N_1565,N_1401,N_1495);
and U1566 (N_1566,N_1469,N_1487);
and U1567 (N_1567,N_1440,N_1408);
or U1568 (N_1568,N_1491,N_1428);
xnor U1569 (N_1569,N_1468,N_1410);
nand U1570 (N_1570,N_1498,N_1421);
nor U1571 (N_1571,N_1479,N_1469);
or U1572 (N_1572,N_1496,N_1422);
xor U1573 (N_1573,N_1410,N_1459);
nand U1574 (N_1574,N_1492,N_1498);
or U1575 (N_1575,N_1431,N_1492);
nor U1576 (N_1576,N_1414,N_1469);
nor U1577 (N_1577,N_1413,N_1463);
nand U1578 (N_1578,N_1471,N_1483);
xor U1579 (N_1579,N_1427,N_1401);
nand U1580 (N_1580,N_1445,N_1485);
nor U1581 (N_1581,N_1409,N_1491);
or U1582 (N_1582,N_1468,N_1401);
or U1583 (N_1583,N_1428,N_1422);
and U1584 (N_1584,N_1469,N_1430);
or U1585 (N_1585,N_1450,N_1496);
nor U1586 (N_1586,N_1457,N_1451);
or U1587 (N_1587,N_1451,N_1495);
or U1588 (N_1588,N_1467,N_1435);
nand U1589 (N_1589,N_1421,N_1484);
and U1590 (N_1590,N_1409,N_1429);
nor U1591 (N_1591,N_1424,N_1456);
nor U1592 (N_1592,N_1471,N_1491);
nor U1593 (N_1593,N_1436,N_1429);
nand U1594 (N_1594,N_1404,N_1462);
xor U1595 (N_1595,N_1418,N_1404);
nor U1596 (N_1596,N_1400,N_1486);
xor U1597 (N_1597,N_1447,N_1450);
nor U1598 (N_1598,N_1447,N_1419);
nand U1599 (N_1599,N_1416,N_1427);
or U1600 (N_1600,N_1534,N_1502);
nand U1601 (N_1601,N_1552,N_1511);
or U1602 (N_1602,N_1500,N_1572);
or U1603 (N_1603,N_1547,N_1551);
and U1604 (N_1604,N_1578,N_1556);
nand U1605 (N_1605,N_1562,N_1579);
and U1606 (N_1606,N_1519,N_1543);
nand U1607 (N_1607,N_1513,N_1506);
or U1608 (N_1608,N_1553,N_1559);
xnor U1609 (N_1609,N_1581,N_1573);
xor U1610 (N_1610,N_1523,N_1544);
nor U1611 (N_1611,N_1555,N_1536);
or U1612 (N_1612,N_1515,N_1517);
and U1613 (N_1613,N_1529,N_1541);
nor U1614 (N_1614,N_1505,N_1509);
or U1615 (N_1615,N_1525,N_1597);
nor U1616 (N_1616,N_1560,N_1586);
nand U1617 (N_1617,N_1528,N_1599);
nor U1618 (N_1618,N_1571,N_1512);
nor U1619 (N_1619,N_1577,N_1566);
nand U1620 (N_1620,N_1522,N_1520);
nand U1621 (N_1621,N_1595,N_1526);
nor U1622 (N_1622,N_1530,N_1587);
and U1623 (N_1623,N_1576,N_1564);
and U1624 (N_1624,N_1507,N_1568);
nand U1625 (N_1625,N_1549,N_1545);
nor U1626 (N_1626,N_1533,N_1591);
nor U1627 (N_1627,N_1594,N_1514);
and U1628 (N_1628,N_1557,N_1501);
and U1629 (N_1629,N_1588,N_1535);
and U1630 (N_1630,N_1538,N_1584);
or U1631 (N_1631,N_1503,N_1596);
nor U1632 (N_1632,N_1590,N_1585);
or U1633 (N_1633,N_1521,N_1580);
xor U1634 (N_1634,N_1546,N_1563);
xnor U1635 (N_1635,N_1569,N_1508);
and U1636 (N_1636,N_1524,N_1575);
or U1637 (N_1637,N_1583,N_1510);
nand U1638 (N_1638,N_1574,N_1527);
nor U1639 (N_1639,N_1532,N_1592);
and U1640 (N_1640,N_1540,N_1582);
nand U1641 (N_1641,N_1531,N_1550);
and U1642 (N_1642,N_1554,N_1542);
nor U1643 (N_1643,N_1598,N_1589);
nor U1644 (N_1644,N_1516,N_1593);
and U1645 (N_1645,N_1518,N_1570);
or U1646 (N_1646,N_1539,N_1565);
nand U1647 (N_1647,N_1537,N_1558);
nor U1648 (N_1648,N_1504,N_1567);
and U1649 (N_1649,N_1561,N_1548);
nor U1650 (N_1650,N_1506,N_1575);
nor U1651 (N_1651,N_1553,N_1520);
nand U1652 (N_1652,N_1503,N_1560);
and U1653 (N_1653,N_1533,N_1550);
and U1654 (N_1654,N_1566,N_1508);
or U1655 (N_1655,N_1543,N_1592);
nand U1656 (N_1656,N_1504,N_1585);
nor U1657 (N_1657,N_1504,N_1516);
or U1658 (N_1658,N_1519,N_1534);
and U1659 (N_1659,N_1540,N_1579);
and U1660 (N_1660,N_1507,N_1534);
or U1661 (N_1661,N_1523,N_1592);
nor U1662 (N_1662,N_1569,N_1528);
or U1663 (N_1663,N_1587,N_1531);
nand U1664 (N_1664,N_1521,N_1567);
and U1665 (N_1665,N_1529,N_1518);
nand U1666 (N_1666,N_1563,N_1552);
nor U1667 (N_1667,N_1542,N_1593);
xor U1668 (N_1668,N_1534,N_1503);
nand U1669 (N_1669,N_1595,N_1576);
nand U1670 (N_1670,N_1551,N_1545);
nand U1671 (N_1671,N_1582,N_1594);
nand U1672 (N_1672,N_1593,N_1525);
nand U1673 (N_1673,N_1544,N_1539);
and U1674 (N_1674,N_1547,N_1508);
xnor U1675 (N_1675,N_1519,N_1500);
or U1676 (N_1676,N_1562,N_1535);
and U1677 (N_1677,N_1573,N_1504);
and U1678 (N_1678,N_1513,N_1559);
or U1679 (N_1679,N_1520,N_1562);
nand U1680 (N_1680,N_1538,N_1501);
or U1681 (N_1681,N_1532,N_1547);
xor U1682 (N_1682,N_1545,N_1537);
nand U1683 (N_1683,N_1532,N_1530);
xnor U1684 (N_1684,N_1502,N_1580);
and U1685 (N_1685,N_1531,N_1512);
nand U1686 (N_1686,N_1579,N_1557);
nand U1687 (N_1687,N_1510,N_1597);
or U1688 (N_1688,N_1530,N_1555);
or U1689 (N_1689,N_1533,N_1559);
or U1690 (N_1690,N_1526,N_1541);
xor U1691 (N_1691,N_1543,N_1520);
xnor U1692 (N_1692,N_1584,N_1595);
or U1693 (N_1693,N_1513,N_1591);
and U1694 (N_1694,N_1570,N_1564);
or U1695 (N_1695,N_1599,N_1506);
or U1696 (N_1696,N_1520,N_1507);
nand U1697 (N_1697,N_1591,N_1540);
and U1698 (N_1698,N_1570,N_1571);
nor U1699 (N_1699,N_1544,N_1509);
nor U1700 (N_1700,N_1639,N_1602);
nand U1701 (N_1701,N_1645,N_1695);
or U1702 (N_1702,N_1667,N_1640);
nor U1703 (N_1703,N_1641,N_1662);
nand U1704 (N_1704,N_1673,N_1643);
and U1705 (N_1705,N_1649,N_1670);
and U1706 (N_1706,N_1614,N_1694);
nor U1707 (N_1707,N_1692,N_1619);
nor U1708 (N_1708,N_1669,N_1635);
nor U1709 (N_1709,N_1690,N_1656);
and U1710 (N_1710,N_1621,N_1609);
and U1711 (N_1711,N_1618,N_1674);
xnor U1712 (N_1712,N_1653,N_1638);
nor U1713 (N_1713,N_1617,N_1628);
and U1714 (N_1714,N_1661,N_1696);
nor U1715 (N_1715,N_1697,N_1648);
and U1716 (N_1716,N_1647,N_1637);
or U1717 (N_1717,N_1675,N_1632);
or U1718 (N_1718,N_1616,N_1698);
xor U1719 (N_1719,N_1629,N_1608);
nor U1720 (N_1720,N_1620,N_1606);
nor U1721 (N_1721,N_1607,N_1681);
and U1722 (N_1722,N_1677,N_1678);
and U1723 (N_1723,N_1600,N_1646);
or U1724 (N_1724,N_1687,N_1611);
nand U1725 (N_1725,N_1686,N_1689);
nor U1726 (N_1726,N_1642,N_1626);
and U1727 (N_1727,N_1685,N_1624);
nor U1728 (N_1728,N_1683,N_1630);
and U1729 (N_1729,N_1633,N_1657);
nand U1730 (N_1730,N_1680,N_1651);
and U1731 (N_1731,N_1631,N_1654);
or U1732 (N_1732,N_1655,N_1663);
nor U1733 (N_1733,N_1622,N_1664);
and U1734 (N_1734,N_1665,N_1691);
nor U1735 (N_1735,N_1671,N_1676);
and U1736 (N_1736,N_1652,N_1636);
and U1737 (N_1737,N_1682,N_1634);
and U1738 (N_1738,N_1612,N_1693);
nor U1739 (N_1739,N_1679,N_1650);
and U1740 (N_1740,N_1699,N_1688);
nand U1741 (N_1741,N_1604,N_1644);
or U1742 (N_1742,N_1660,N_1684);
and U1743 (N_1743,N_1625,N_1672);
nand U1744 (N_1744,N_1610,N_1613);
nand U1745 (N_1745,N_1615,N_1601);
xnor U1746 (N_1746,N_1623,N_1603);
xnor U1747 (N_1747,N_1666,N_1668);
or U1748 (N_1748,N_1605,N_1658);
xor U1749 (N_1749,N_1627,N_1659);
nor U1750 (N_1750,N_1679,N_1647);
nor U1751 (N_1751,N_1635,N_1638);
nand U1752 (N_1752,N_1668,N_1632);
and U1753 (N_1753,N_1614,N_1619);
and U1754 (N_1754,N_1680,N_1659);
nand U1755 (N_1755,N_1645,N_1604);
or U1756 (N_1756,N_1637,N_1670);
and U1757 (N_1757,N_1634,N_1669);
nand U1758 (N_1758,N_1697,N_1668);
nand U1759 (N_1759,N_1631,N_1677);
nor U1760 (N_1760,N_1674,N_1623);
and U1761 (N_1761,N_1681,N_1638);
nor U1762 (N_1762,N_1646,N_1608);
nor U1763 (N_1763,N_1648,N_1606);
nand U1764 (N_1764,N_1616,N_1694);
and U1765 (N_1765,N_1625,N_1697);
nand U1766 (N_1766,N_1602,N_1668);
nor U1767 (N_1767,N_1603,N_1610);
nor U1768 (N_1768,N_1666,N_1620);
nand U1769 (N_1769,N_1602,N_1669);
nor U1770 (N_1770,N_1618,N_1663);
and U1771 (N_1771,N_1675,N_1612);
nand U1772 (N_1772,N_1663,N_1684);
nand U1773 (N_1773,N_1623,N_1602);
nand U1774 (N_1774,N_1691,N_1677);
or U1775 (N_1775,N_1621,N_1655);
nand U1776 (N_1776,N_1696,N_1612);
nand U1777 (N_1777,N_1646,N_1664);
and U1778 (N_1778,N_1699,N_1682);
or U1779 (N_1779,N_1645,N_1623);
nor U1780 (N_1780,N_1698,N_1674);
nor U1781 (N_1781,N_1697,N_1690);
nand U1782 (N_1782,N_1643,N_1615);
nand U1783 (N_1783,N_1670,N_1658);
nand U1784 (N_1784,N_1624,N_1664);
nor U1785 (N_1785,N_1616,N_1614);
and U1786 (N_1786,N_1667,N_1673);
or U1787 (N_1787,N_1671,N_1699);
or U1788 (N_1788,N_1646,N_1638);
nor U1789 (N_1789,N_1673,N_1659);
nor U1790 (N_1790,N_1611,N_1623);
xor U1791 (N_1791,N_1673,N_1625);
or U1792 (N_1792,N_1674,N_1696);
nor U1793 (N_1793,N_1693,N_1662);
xor U1794 (N_1794,N_1634,N_1625);
nor U1795 (N_1795,N_1608,N_1664);
nand U1796 (N_1796,N_1642,N_1689);
nand U1797 (N_1797,N_1637,N_1632);
xor U1798 (N_1798,N_1661,N_1663);
nand U1799 (N_1799,N_1633,N_1606);
and U1800 (N_1800,N_1720,N_1701);
nand U1801 (N_1801,N_1775,N_1780);
nand U1802 (N_1802,N_1777,N_1782);
or U1803 (N_1803,N_1774,N_1766);
and U1804 (N_1804,N_1781,N_1753);
or U1805 (N_1805,N_1754,N_1725);
or U1806 (N_1806,N_1711,N_1772);
xor U1807 (N_1807,N_1783,N_1712);
nor U1808 (N_1808,N_1719,N_1793);
and U1809 (N_1809,N_1724,N_1773);
nand U1810 (N_1810,N_1759,N_1798);
or U1811 (N_1811,N_1742,N_1749);
nor U1812 (N_1812,N_1713,N_1731);
nand U1813 (N_1813,N_1760,N_1735);
xor U1814 (N_1814,N_1791,N_1708);
or U1815 (N_1815,N_1750,N_1737);
and U1816 (N_1816,N_1716,N_1704);
nand U1817 (N_1817,N_1768,N_1733);
or U1818 (N_1818,N_1746,N_1743);
nor U1819 (N_1819,N_1769,N_1751);
and U1820 (N_1820,N_1789,N_1717);
xor U1821 (N_1821,N_1752,N_1715);
or U1822 (N_1822,N_1799,N_1718);
nor U1823 (N_1823,N_1744,N_1796);
or U1824 (N_1824,N_1787,N_1765);
nor U1825 (N_1825,N_1723,N_1757);
nand U1826 (N_1826,N_1790,N_1706);
nor U1827 (N_1827,N_1707,N_1763);
or U1828 (N_1828,N_1700,N_1729);
nor U1829 (N_1829,N_1732,N_1758);
or U1830 (N_1830,N_1755,N_1770);
nand U1831 (N_1831,N_1710,N_1794);
or U1832 (N_1832,N_1764,N_1741);
or U1833 (N_1833,N_1727,N_1702);
nand U1834 (N_1834,N_1739,N_1721);
xnor U1835 (N_1835,N_1785,N_1738);
xor U1836 (N_1836,N_1748,N_1709);
nand U1837 (N_1837,N_1730,N_1705);
and U1838 (N_1838,N_1771,N_1761);
nor U1839 (N_1839,N_1784,N_1788);
nand U1840 (N_1840,N_1779,N_1795);
and U1841 (N_1841,N_1762,N_1734);
nand U1842 (N_1842,N_1747,N_1703);
or U1843 (N_1843,N_1726,N_1792);
and U1844 (N_1844,N_1722,N_1740);
xnor U1845 (N_1845,N_1778,N_1736);
and U1846 (N_1846,N_1714,N_1786);
nor U1847 (N_1847,N_1797,N_1767);
xor U1848 (N_1848,N_1756,N_1745);
or U1849 (N_1849,N_1728,N_1776);
nand U1850 (N_1850,N_1767,N_1736);
nor U1851 (N_1851,N_1723,N_1791);
nand U1852 (N_1852,N_1751,N_1757);
and U1853 (N_1853,N_1729,N_1796);
and U1854 (N_1854,N_1707,N_1747);
nand U1855 (N_1855,N_1764,N_1717);
and U1856 (N_1856,N_1734,N_1700);
nor U1857 (N_1857,N_1715,N_1760);
nand U1858 (N_1858,N_1740,N_1742);
nand U1859 (N_1859,N_1716,N_1703);
nor U1860 (N_1860,N_1790,N_1794);
or U1861 (N_1861,N_1700,N_1780);
nor U1862 (N_1862,N_1791,N_1751);
or U1863 (N_1863,N_1777,N_1759);
or U1864 (N_1864,N_1767,N_1720);
and U1865 (N_1865,N_1751,N_1762);
nor U1866 (N_1866,N_1745,N_1737);
or U1867 (N_1867,N_1709,N_1728);
nand U1868 (N_1868,N_1739,N_1753);
xor U1869 (N_1869,N_1716,N_1713);
or U1870 (N_1870,N_1778,N_1709);
or U1871 (N_1871,N_1782,N_1789);
nand U1872 (N_1872,N_1733,N_1736);
xor U1873 (N_1873,N_1719,N_1715);
nor U1874 (N_1874,N_1708,N_1790);
nor U1875 (N_1875,N_1733,N_1732);
or U1876 (N_1876,N_1769,N_1756);
or U1877 (N_1877,N_1701,N_1716);
nor U1878 (N_1878,N_1742,N_1754);
and U1879 (N_1879,N_1760,N_1764);
and U1880 (N_1880,N_1733,N_1724);
or U1881 (N_1881,N_1715,N_1782);
and U1882 (N_1882,N_1763,N_1756);
xor U1883 (N_1883,N_1732,N_1740);
and U1884 (N_1884,N_1789,N_1788);
or U1885 (N_1885,N_1749,N_1751);
nand U1886 (N_1886,N_1791,N_1730);
nand U1887 (N_1887,N_1723,N_1750);
and U1888 (N_1888,N_1711,N_1726);
and U1889 (N_1889,N_1782,N_1737);
and U1890 (N_1890,N_1700,N_1777);
and U1891 (N_1891,N_1753,N_1715);
or U1892 (N_1892,N_1788,N_1777);
and U1893 (N_1893,N_1775,N_1713);
or U1894 (N_1894,N_1732,N_1727);
xnor U1895 (N_1895,N_1790,N_1726);
xor U1896 (N_1896,N_1712,N_1723);
nor U1897 (N_1897,N_1734,N_1787);
or U1898 (N_1898,N_1785,N_1752);
nor U1899 (N_1899,N_1773,N_1770);
or U1900 (N_1900,N_1887,N_1843);
nor U1901 (N_1901,N_1855,N_1858);
xnor U1902 (N_1902,N_1882,N_1808);
xnor U1903 (N_1903,N_1883,N_1800);
and U1904 (N_1904,N_1863,N_1867);
or U1905 (N_1905,N_1815,N_1810);
or U1906 (N_1906,N_1868,N_1878);
xor U1907 (N_1907,N_1884,N_1847);
nor U1908 (N_1908,N_1820,N_1854);
or U1909 (N_1909,N_1865,N_1864);
nor U1910 (N_1910,N_1888,N_1895);
or U1911 (N_1911,N_1848,N_1830);
nor U1912 (N_1912,N_1874,N_1892);
nor U1913 (N_1913,N_1871,N_1838);
nand U1914 (N_1914,N_1852,N_1856);
nand U1915 (N_1915,N_1826,N_1876);
or U1916 (N_1916,N_1801,N_1827);
and U1917 (N_1917,N_1879,N_1845);
nor U1918 (N_1918,N_1893,N_1859);
and U1919 (N_1919,N_1802,N_1872);
nand U1920 (N_1920,N_1829,N_1840);
and U1921 (N_1921,N_1818,N_1823);
and U1922 (N_1922,N_1891,N_1898);
xor U1923 (N_1923,N_1803,N_1833);
or U1924 (N_1924,N_1875,N_1899);
nor U1925 (N_1925,N_1870,N_1821);
nor U1926 (N_1926,N_1862,N_1846);
nor U1927 (N_1927,N_1842,N_1873);
nand U1928 (N_1928,N_1836,N_1894);
and U1929 (N_1929,N_1881,N_1851);
or U1930 (N_1930,N_1849,N_1839);
nor U1931 (N_1931,N_1817,N_1809);
or U1932 (N_1932,N_1832,N_1831);
or U1933 (N_1933,N_1857,N_1860);
xor U1934 (N_1934,N_1813,N_1869);
xor U1935 (N_1935,N_1896,N_1841);
nand U1936 (N_1936,N_1861,N_1822);
xor U1937 (N_1937,N_1866,N_1816);
nand U1938 (N_1938,N_1850,N_1889);
nor U1939 (N_1939,N_1844,N_1819);
and U1940 (N_1940,N_1804,N_1824);
or U1941 (N_1941,N_1806,N_1885);
nand U1942 (N_1942,N_1834,N_1825);
nand U1943 (N_1943,N_1837,N_1807);
nor U1944 (N_1944,N_1897,N_1828);
nand U1945 (N_1945,N_1890,N_1814);
nor U1946 (N_1946,N_1886,N_1835);
and U1947 (N_1947,N_1811,N_1805);
and U1948 (N_1948,N_1880,N_1877);
xor U1949 (N_1949,N_1812,N_1853);
and U1950 (N_1950,N_1809,N_1874);
nand U1951 (N_1951,N_1803,N_1840);
nand U1952 (N_1952,N_1884,N_1860);
and U1953 (N_1953,N_1885,N_1860);
nand U1954 (N_1954,N_1843,N_1882);
nor U1955 (N_1955,N_1804,N_1888);
nor U1956 (N_1956,N_1884,N_1820);
and U1957 (N_1957,N_1834,N_1851);
xor U1958 (N_1958,N_1881,N_1820);
and U1959 (N_1959,N_1849,N_1870);
xor U1960 (N_1960,N_1840,N_1895);
and U1961 (N_1961,N_1834,N_1891);
and U1962 (N_1962,N_1816,N_1814);
and U1963 (N_1963,N_1878,N_1836);
or U1964 (N_1964,N_1822,N_1802);
and U1965 (N_1965,N_1866,N_1896);
nor U1966 (N_1966,N_1897,N_1898);
nand U1967 (N_1967,N_1817,N_1869);
or U1968 (N_1968,N_1876,N_1865);
and U1969 (N_1969,N_1822,N_1880);
xnor U1970 (N_1970,N_1887,N_1815);
nor U1971 (N_1971,N_1886,N_1807);
xor U1972 (N_1972,N_1875,N_1815);
nand U1973 (N_1973,N_1833,N_1865);
nor U1974 (N_1974,N_1839,N_1878);
or U1975 (N_1975,N_1800,N_1828);
and U1976 (N_1976,N_1851,N_1849);
and U1977 (N_1977,N_1842,N_1824);
nor U1978 (N_1978,N_1850,N_1849);
nor U1979 (N_1979,N_1874,N_1885);
xnor U1980 (N_1980,N_1807,N_1885);
and U1981 (N_1981,N_1821,N_1862);
nand U1982 (N_1982,N_1852,N_1848);
nand U1983 (N_1983,N_1836,N_1871);
nor U1984 (N_1984,N_1834,N_1893);
xnor U1985 (N_1985,N_1846,N_1830);
or U1986 (N_1986,N_1830,N_1820);
nand U1987 (N_1987,N_1836,N_1891);
and U1988 (N_1988,N_1860,N_1810);
or U1989 (N_1989,N_1861,N_1835);
or U1990 (N_1990,N_1807,N_1870);
or U1991 (N_1991,N_1896,N_1831);
and U1992 (N_1992,N_1801,N_1820);
or U1993 (N_1993,N_1802,N_1842);
nand U1994 (N_1994,N_1833,N_1802);
and U1995 (N_1995,N_1857,N_1880);
and U1996 (N_1996,N_1810,N_1850);
nand U1997 (N_1997,N_1801,N_1860);
or U1998 (N_1998,N_1809,N_1816);
nand U1999 (N_1999,N_1847,N_1851);
xnor U2000 (N_2000,N_1981,N_1906);
or U2001 (N_2001,N_1902,N_1999);
nor U2002 (N_2002,N_1936,N_1911);
nor U2003 (N_2003,N_1961,N_1942);
nand U2004 (N_2004,N_1928,N_1924);
or U2005 (N_2005,N_1949,N_1955);
or U2006 (N_2006,N_1984,N_1945);
nand U2007 (N_2007,N_1957,N_1917);
and U2008 (N_2008,N_1920,N_1925);
nor U2009 (N_2009,N_1974,N_1964);
nand U2010 (N_2010,N_1913,N_1940);
nand U2011 (N_2011,N_1980,N_1990);
and U2012 (N_2012,N_1988,N_1927);
and U2013 (N_2013,N_1909,N_1907);
xor U2014 (N_2014,N_1975,N_1979);
and U2015 (N_2015,N_1959,N_1992);
or U2016 (N_2016,N_1954,N_1908);
or U2017 (N_2017,N_1951,N_1941);
or U2018 (N_2018,N_1921,N_1983);
nor U2019 (N_2019,N_1929,N_1969);
xnor U2020 (N_2020,N_1944,N_1965);
or U2021 (N_2021,N_1976,N_1994);
or U2022 (N_2022,N_1987,N_1916);
or U2023 (N_2023,N_1958,N_1931);
nand U2024 (N_2024,N_1900,N_1934);
or U2025 (N_2025,N_1950,N_1991);
nor U2026 (N_2026,N_1963,N_1986);
or U2027 (N_2027,N_1962,N_1995);
nor U2028 (N_2028,N_1989,N_1996);
nand U2029 (N_2029,N_1977,N_1923);
and U2030 (N_2030,N_1912,N_1946);
nand U2031 (N_2031,N_1982,N_1953);
nor U2032 (N_2032,N_1938,N_1915);
and U2033 (N_2033,N_1904,N_1937);
xnor U2034 (N_2034,N_1973,N_1935);
nor U2035 (N_2035,N_1905,N_1930);
and U2036 (N_2036,N_1910,N_1993);
nand U2037 (N_2037,N_1967,N_1948);
or U2038 (N_2038,N_1901,N_1918);
xor U2039 (N_2039,N_1997,N_1985);
or U2040 (N_2040,N_1956,N_1971);
nor U2041 (N_2041,N_1943,N_1922);
and U2042 (N_2042,N_1952,N_1978);
and U2043 (N_2043,N_1972,N_1926);
and U2044 (N_2044,N_1960,N_1998);
nor U2045 (N_2045,N_1947,N_1903);
nand U2046 (N_2046,N_1919,N_1970);
and U2047 (N_2047,N_1939,N_1966);
or U2048 (N_2048,N_1914,N_1933);
and U2049 (N_2049,N_1968,N_1932);
or U2050 (N_2050,N_1971,N_1946);
xnor U2051 (N_2051,N_1924,N_1953);
or U2052 (N_2052,N_1967,N_1936);
nor U2053 (N_2053,N_1962,N_1941);
nor U2054 (N_2054,N_1966,N_1992);
or U2055 (N_2055,N_1995,N_1977);
nor U2056 (N_2056,N_1966,N_1961);
nor U2057 (N_2057,N_1933,N_1987);
nor U2058 (N_2058,N_1998,N_1949);
and U2059 (N_2059,N_1979,N_1918);
nand U2060 (N_2060,N_1937,N_1901);
nand U2061 (N_2061,N_1920,N_1995);
and U2062 (N_2062,N_1997,N_1977);
nor U2063 (N_2063,N_1973,N_1902);
or U2064 (N_2064,N_1907,N_1986);
nor U2065 (N_2065,N_1946,N_1952);
nor U2066 (N_2066,N_1989,N_1915);
and U2067 (N_2067,N_1954,N_1910);
nor U2068 (N_2068,N_1908,N_1941);
nor U2069 (N_2069,N_1970,N_1927);
nand U2070 (N_2070,N_1901,N_1935);
xnor U2071 (N_2071,N_1923,N_1942);
nor U2072 (N_2072,N_1958,N_1921);
nor U2073 (N_2073,N_1920,N_1938);
nor U2074 (N_2074,N_1939,N_1990);
or U2075 (N_2075,N_1911,N_1951);
nand U2076 (N_2076,N_1907,N_1966);
nand U2077 (N_2077,N_1971,N_1911);
and U2078 (N_2078,N_1911,N_1981);
and U2079 (N_2079,N_1994,N_1931);
and U2080 (N_2080,N_1998,N_1962);
nand U2081 (N_2081,N_1943,N_1996);
or U2082 (N_2082,N_1936,N_1907);
nand U2083 (N_2083,N_1912,N_1929);
and U2084 (N_2084,N_1990,N_1994);
nor U2085 (N_2085,N_1965,N_1999);
and U2086 (N_2086,N_1978,N_1992);
nor U2087 (N_2087,N_1917,N_1935);
and U2088 (N_2088,N_1987,N_1902);
or U2089 (N_2089,N_1942,N_1925);
or U2090 (N_2090,N_1948,N_1915);
or U2091 (N_2091,N_1973,N_1913);
xnor U2092 (N_2092,N_1926,N_1933);
nor U2093 (N_2093,N_1925,N_1955);
and U2094 (N_2094,N_1977,N_1921);
nor U2095 (N_2095,N_1947,N_1978);
and U2096 (N_2096,N_1982,N_1902);
nor U2097 (N_2097,N_1900,N_1904);
nor U2098 (N_2098,N_1913,N_1979);
or U2099 (N_2099,N_1932,N_1908);
or U2100 (N_2100,N_2044,N_2059);
nand U2101 (N_2101,N_2003,N_2007);
and U2102 (N_2102,N_2032,N_2041);
nor U2103 (N_2103,N_2034,N_2078);
and U2104 (N_2104,N_2023,N_2083);
or U2105 (N_2105,N_2058,N_2021);
or U2106 (N_2106,N_2049,N_2091);
nand U2107 (N_2107,N_2082,N_2063);
nor U2108 (N_2108,N_2000,N_2079);
nand U2109 (N_2109,N_2026,N_2071);
xnor U2110 (N_2110,N_2085,N_2068);
or U2111 (N_2111,N_2054,N_2090);
or U2112 (N_2112,N_2099,N_2040);
xor U2113 (N_2113,N_2043,N_2069);
nor U2114 (N_2114,N_2012,N_2053);
or U2115 (N_2115,N_2039,N_2006);
or U2116 (N_2116,N_2076,N_2013);
or U2117 (N_2117,N_2051,N_2092);
or U2118 (N_2118,N_2020,N_2008);
or U2119 (N_2119,N_2019,N_2022);
nand U2120 (N_2120,N_2017,N_2065);
nand U2121 (N_2121,N_2070,N_2005);
nor U2122 (N_2122,N_2025,N_2095);
nor U2123 (N_2123,N_2050,N_2073);
and U2124 (N_2124,N_2087,N_2094);
and U2125 (N_2125,N_2061,N_2030);
xor U2126 (N_2126,N_2014,N_2088);
nand U2127 (N_2127,N_2060,N_2015);
nor U2128 (N_2128,N_2081,N_2033);
and U2129 (N_2129,N_2057,N_2042);
and U2130 (N_2130,N_2052,N_2046);
or U2131 (N_2131,N_2077,N_2056);
nor U2132 (N_2132,N_2035,N_2072);
nand U2133 (N_2133,N_2004,N_2002);
or U2134 (N_2134,N_2064,N_2097);
nand U2135 (N_2135,N_2075,N_2001);
and U2136 (N_2136,N_2011,N_2031);
and U2137 (N_2137,N_2067,N_2027);
and U2138 (N_2138,N_2045,N_2024);
and U2139 (N_2139,N_2048,N_2096);
or U2140 (N_2140,N_2028,N_2036);
or U2141 (N_2141,N_2055,N_2009);
and U2142 (N_2142,N_2047,N_2086);
and U2143 (N_2143,N_2089,N_2074);
or U2144 (N_2144,N_2016,N_2062);
nor U2145 (N_2145,N_2093,N_2098);
xor U2146 (N_2146,N_2084,N_2038);
xnor U2147 (N_2147,N_2029,N_2037);
or U2148 (N_2148,N_2080,N_2018);
nand U2149 (N_2149,N_2010,N_2066);
xor U2150 (N_2150,N_2063,N_2024);
or U2151 (N_2151,N_2026,N_2055);
or U2152 (N_2152,N_2076,N_2091);
or U2153 (N_2153,N_2002,N_2022);
or U2154 (N_2154,N_2090,N_2018);
nor U2155 (N_2155,N_2008,N_2087);
nand U2156 (N_2156,N_2087,N_2053);
nor U2157 (N_2157,N_2085,N_2050);
or U2158 (N_2158,N_2073,N_2035);
nor U2159 (N_2159,N_2045,N_2020);
xnor U2160 (N_2160,N_2062,N_2026);
and U2161 (N_2161,N_2018,N_2061);
nor U2162 (N_2162,N_2001,N_2015);
or U2163 (N_2163,N_2039,N_2003);
and U2164 (N_2164,N_2058,N_2090);
xor U2165 (N_2165,N_2018,N_2082);
and U2166 (N_2166,N_2013,N_2088);
nand U2167 (N_2167,N_2033,N_2054);
nand U2168 (N_2168,N_2098,N_2085);
and U2169 (N_2169,N_2007,N_2081);
nand U2170 (N_2170,N_2086,N_2012);
nand U2171 (N_2171,N_2060,N_2083);
or U2172 (N_2172,N_2017,N_2045);
or U2173 (N_2173,N_2032,N_2064);
nor U2174 (N_2174,N_2038,N_2080);
nand U2175 (N_2175,N_2075,N_2090);
nor U2176 (N_2176,N_2082,N_2086);
nor U2177 (N_2177,N_2029,N_2012);
nor U2178 (N_2178,N_2092,N_2081);
or U2179 (N_2179,N_2071,N_2036);
and U2180 (N_2180,N_2043,N_2080);
or U2181 (N_2181,N_2067,N_2008);
nor U2182 (N_2182,N_2088,N_2038);
or U2183 (N_2183,N_2042,N_2058);
nor U2184 (N_2184,N_2020,N_2013);
nor U2185 (N_2185,N_2058,N_2018);
and U2186 (N_2186,N_2082,N_2088);
and U2187 (N_2187,N_2024,N_2097);
nor U2188 (N_2188,N_2025,N_2086);
nand U2189 (N_2189,N_2021,N_2090);
nor U2190 (N_2190,N_2029,N_2034);
or U2191 (N_2191,N_2027,N_2014);
or U2192 (N_2192,N_2030,N_2046);
or U2193 (N_2193,N_2050,N_2042);
nor U2194 (N_2194,N_2093,N_2031);
nor U2195 (N_2195,N_2080,N_2053);
nor U2196 (N_2196,N_2084,N_2044);
nand U2197 (N_2197,N_2022,N_2039);
nor U2198 (N_2198,N_2098,N_2043);
nand U2199 (N_2199,N_2091,N_2097);
nand U2200 (N_2200,N_2165,N_2171);
nand U2201 (N_2201,N_2143,N_2175);
or U2202 (N_2202,N_2166,N_2112);
nand U2203 (N_2203,N_2109,N_2162);
xor U2204 (N_2204,N_2153,N_2135);
nor U2205 (N_2205,N_2137,N_2134);
and U2206 (N_2206,N_2148,N_2114);
nor U2207 (N_2207,N_2110,N_2123);
and U2208 (N_2208,N_2176,N_2189);
nor U2209 (N_2209,N_2130,N_2106);
or U2210 (N_2210,N_2121,N_2152);
and U2211 (N_2211,N_2173,N_2149);
or U2212 (N_2212,N_2124,N_2151);
nand U2213 (N_2213,N_2194,N_2182);
or U2214 (N_2214,N_2188,N_2128);
nand U2215 (N_2215,N_2111,N_2199);
nand U2216 (N_2216,N_2172,N_2169);
and U2217 (N_2217,N_2187,N_2132);
or U2218 (N_2218,N_2144,N_2158);
nand U2219 (N_2219,N_2104,N_2160);
or U2220 (N_2220,N_2113,N_2100);
and U2221 (N_2221,N_2125,N_2161);
nand U2222 (N_2222,N_2138,N_2177);
xor U2223 (N_2223,N_2164,N_2180);
and U2224 (N_2224,N_2181,N_2133);
or U2225 (N_2225,N_2139,N_2178);
xnor U2226 (N_2226,N_2150,N_2195);
or U2227 (N_2227,N_2167,N_2131);
and U2228 (N_2228,N_2103,N_2126);
nor U2229 (N_2229,N_2193,N_2156);
and U2230 (N_2230,N_2185,N_2191);
or U2231 (N_2231,N_2129,N_2116);
nand U2232 (N_2232,N_2192,N_2145);
nor U2233 (N_2233,N_2183,N_2105);
and U2234 (N_2234,N_2118,N_2184);
nor U2235 (N_2235,N_2127,N_2154);
xnor U2236 (N_2236,N_2136,N_2117);
nor U2237 (N_2237,N_2179,N_2101);
nand U2238 (N_2238,N_2157,N_2107);
or U2239 (N_2239,N_2120,N_2102);
and U2240 (N_2240,N_2115,N_2140);
nand U2241 (N_2241,N_2190,N_2186);
and U2242 (N_2242,N_2163,N_2119);
or U2243 (N_2243,N_2147,N_2198);
or U2244 (N_2244,N_2146,N_2197);
nand U2245 (N_2245,N_2196,N_2170);
and U2246 (N_2246,N_2122,N_2142);
nor U2247 (N_2247,N_2159,N_2141);
nor U2248 (N_2248,N_2174,N_2155);
and U2249 (N_2249,N_2168,N_2108);
nand U2250 (N_2250,N_2101,N_2131);
or U2251 (N_2251,N_2124,N_2196);
xnor U2252 (N_2252,N_2172,N_2184);
or U2253 (N_2253,N_2198,N_2171);
or U2254 (N_2254,N_2160,N_2171);
and U2255 (N_2255,N_2135,N_2178);
nand U2256 (N_2256,N_2107,N_2142);
and U2257 (N_2257,N_2175,N_2114);
xnor U2258 (N_2258,N_2113,N_2130);
or U2259 (N_2259,N_2160,N_2189);
or U2260 (N_2260,N_2108,N_2190);
nor U2261 (N_2261,N_2108,N_2164);
nand U2262 (N_2262,N_2117,N_2146);
nor U2263 (N_2263,N_2126,N_2190);
and U2264 (N_2264,N_2160,N_2119);
nand U2265 (N_2265,N_2131,N_2148);
and U2266 (N_2266,N_2166,N_2168);
xnor U2267 (N_2267,N_2114,N_2145);
and U2268 (N_2268,N_2188,N_2139);
nor U2269 (N_2269,N_2158,N_2140);
nand U2270 (N_2270,N_2137,N_2193);
or U2271 (N_2271,N_2117,N_2198);
and U2272 (N_2272,N_2131,N_2168);
and U2273 (N_2273,N_2140,N_2198);
nand U2274 (N_2274,N_2191,N_2196);
and U2275 (N_2275,N_2160,N_2143);
or U2276 (N_2276,N_2117,N_2100);
or U2277 (N_2277,N_2138,N_2156);
or U2278 (N_2278,N_2162,N_2188);
xnor U2279 (N_2279,N_2159,N_2169);
nand U2280 (N_2280,N_2159,N_2100);
nand U2281 (N_2281,N_2143,N_2162);
and U2282 (N_2282,N_2119,N_2196);
and U2283 (N_2283,N_2119,N_2172);
nor U2284 (N_2284,N_2105,N_2167);
or U2285 (N_2285,N_2125,N_2148);
xor U2286 (N_2286,N_2155,N_2124);
or U2287 (N_2287,N_2146,N_2185);
or U2288 (N_2288,N_2111,N_2129);
and U2289 (N_2289,N_2188,N_2167);
and U2290 (N_2290,N_2114,N_2146);
or U2291 (N_2291,N_2163,N_2177);
nand U2292 (N_2292,N_2197,N_2160);
nor U2293 (N_2293,N_2119,N_2108);
nand U2294 (N_2294,N_2178,N_2188);
nor U2295 (N_2295,N_2123,N_2147);
nor U2296 (N_2296,N_2132,N_2128);
nand U2297 (N_2297,N_2164,N_2115);
nor U2298 (N_2298,N_2176,N_2165);
nor U2299 (N_2299,N_2122,N_2129);
or U2300 (N_2300,N_2204,N_2255);
nor U2301 (N_2301,N_2235,N_2274);
and U2302 (N_2302,N_2236,N_2224);
or U2303 (N_2303,N_2272,N_2291);
nor U2304 (N_2304,N_2242,N_2282);
xnor U2305 (N_2305,N_2222,N_2220);
xnor U2306 (N_2306,N_2268,N_2207);
or U2307 (N_2307,N_2244,N_2232);
or U2308 (N_2308,N_2248,N_2289);
and U2309 (N_2309,N_2283,N_2249);
or U2310 (N_2310,N_2221,N_2257);
or U2311 (N_2311,N_2214,N_2265);
and U2312 (N_2312,N_2234,N_2203);
nand U2313 (N_2313,N_2208,N_2278);
nor U2314 (N_2314,N_2299,N_2211);
nor U2315 (N_2315,N_2284,N_2266);
nor U2316 (N_2316,N_2205,N_2271);
xor U2317 (N_2317,N_2276,N_2240);
nand U2318 (N_2318,N_2215,N_2286);
nand U2319 (N_2319,N_2201,N_2213);
or U2320 (N_2320,N_2275,N_2262);
nand U2321 (N_2321,N_2228,N_2200);
nor U2322 (N_2322,N_2239,N_2269);
nor U2323 (N_2323,N_2285,N_2258);
nand U2324 (N_2324,N_2238,N_2287);
nor U2325 (N_2325,N_2253,N_2295);
nor U2326 (N_2326,N_2233,N_2259);
nor U2327 (N_2327,N_2277,N_2260);
xor U2328 (N_2328,N_2293,N_2273);
and U2329 (N_2329,N_2227,N_2254);
nor U2330 (N_2330,N_2296,N_2251);
nor U2331 (N_2331,N_2237,N_2297);
nor U2332 (N_2332,N_2210,N_2264);
and U2333 (N_2333,N_2217,N_2209);
nand U2334 (N_2334,N_2247,N_2294);
or U2335 (N_2335,N_2298,N_2212);
nor U2336 (N_2336,N_2219,N_2280);
xor U2337 (N_2337,N_2206,N_2270);
nor U2338 (N_2338,N_2225,N_2261);
nand U2339 (N_2339,N_2288,N_2243);
or U2340 (N_2340,N_2226,N_2246);
nor U2341 (N_2341,N_2290,N_2229);
or U2342 (N_2342,N_2267,N_2241);
and U2343 (N_2343,N_2231,N_2223);
xnor U2344 (N_2344,N_2292,N_2202);
and U2345 (N_2345,N_2230,N_2218);
xor U2346 (N_2346,N_2281,N_2245);
or U2347 (N_2347,N_2250,N_2252);
and U2348 (N_2348,N_2216,N_2256);
nand U2349 (N_2349,N_2279,N_2263);
or U2350 (N_2350,N_2251,N_2218);
and U2351 (N_2351,N_2230,N_2228);
nand U2352 (N_2352,N_2295,N_2233);
nor U2353 (N_2353,N_2284,N_2260);
xor U2354 (N_2354,N_2204,N_2262);
or U2355 (N_2355,N_2202,N_2203);
nor U2356 (N_2356,N_2291,N_2204);
or U2357 (N_2357,N_2295,N_2223);
nand U2358 (N_2358,N_2290,N_2299);
nor U2359 (N_2359,N_2226,N_2231);
and U2360 (N_2360,N_2228,N_2247);
nor U2361 (N_2361,N_2220,N_2250);
and U2362 (N_2362,N_2225,N_2227);
nor U2363 (N_2363,N_2202,N_2281);
and U2364 (N_2364,N_2290,N_2200);
and U2365 (N_2365,N_2294,N_2236);
or U2366 (N_2366,N_2212,N_2232);
nor U2367 (N_2367,N_2263,N_2292);
and U2368 (N_2368,N_2278,N_2266);
nand U2369 (N_2369,N_2283,N_2231);
nand U2370 (N_2370,N_2284,N_2203);
nor U2371 (N_2371,N_2295,N_2200);
nand U2372 (N_2372,N_2219,N_2255);
and U2373 (N_2373,N_2218,N_2264);
xor U2374 (N_2374,N_2277,N_2250);
nand U2375 (N_2375,N_2273,N_2246);
xor U2376 (N_2376,N_2279,N_2231);
or U2377 (N_2377,N_2202,N_2233);
nand U2378 (N_2378,N_2241,N_2212);
nor U2379 (N_2379,N_2283,N_2252);
and U2380 (N_2380,N_2280,N_2227);
nand U2381 (N_2381,N_2233,N_2232);
nand U2382 (N_2382,N_2219,N_2237);
and U2383 (N_2383,N_2217,N_2242);
or U2384 (N_2384,N_2204,N_2210);
and U2385 (N_2385,N_2286,N_2283);
xor U2386 (N_2386,N_2290,N_2237);
nand U2387 (N_2387,N_2270,N_2208);
nor U2388 (N_2388,N_2263,N_2249);
or U2389 (N_2389,N_2298,N_2294);
nor U2390 (N_2390,N_2241,N_2266);
and U2391 (N_2391,N_2288,N_2275);
and U2392 (N_2392,N_2222,N_2228);
and U2393 (N_2393,N_2242,N_2255);
and U2394 (N_2394,N_2211,N_2259);
nand U2395 (N_2395,N_2209,N_2223);
or U2396 (N_2396,N_2221,N_2238);
nor U2397 (N_2397,N_2203,N_2246);
and U2398 (N_2398,N_2200,N_2297);
and U2399 (N_2399,N_2288,N_2289);
xnor U2400 (N_2400,N_2327,N_2388);
nand U2401 (N_2401,N_2348,N_2334);
or U2402 (N_2402,N_2340,N_2305);
nand U2403 (N_2403,N_2338,N_2352);
nand U2404 (N_2404,N_2331,N_2317);
or U2405 (N_2405,N_2350,N_2328);
or U2406 (N_2406,N_2313,N_2367);
or U2407 (N_2407,N_2363,N_2333);
and U2408 (N_2408,N_2337,N_2311);
xor U2409 (N_2409,N_2319,N_2358);
or U2410 (N_2410,N_2391,N_2339);
and U2411 (N_2411,N_2355,N_2375);
or U2412 (N_2412,N_2394,N_2324);
nor U2413 (N_2413,N_2360,N_2378);
and U2414 (N_2414,N_2326,N_2349);
nand U2415 (N_2415,N_2309,N_2345);
and U2416 (N_2416,N_2368,N_2392);
nor U2417 (N_2417,N_2332,N_2310);
nand U2418 (N_2418,N_2336,N_2399);
xor U2419 (N_2419,N_2369,N_2323);
nand U2420 (N_2420,N_2370,N_2380);
and U2421 (N_2421,N_2353,N_2372);
and U2422 (N_2422,N_2390,N_2325);
nor U2423 (N_2423,N_2354,N_2308);
and U2424 (N_2424,N_2362,N_2377);
nand U2425 (N_2425,N_2321,N_2351);
or U2426 (N_2426,N_2383,N_2389);
nand U2427 (N_2427,N_2374,N_2307);
and U2428 (N_2428,N_2396,N_2306);
or U2429 (N_2429,N_2330,N_2304);
and U2430 (N_2430,N_2300,N_2364);
and U2431 (N_2431,N_2373,N_2316);
or U2432 (N_2432,N_2393,N_2329);
or U2433 (N_2433,N_2397,N_2314);
or U2434 (N_2434,N_2385,N_2315);
nand U2435 (N_2435,N_2343,N_2301);
nand U2436 (N_2436,N_2318,N_2342);
nand U2437 (N_2437,N_2366,N_2357);
nand U2438 (N_2438,N_2371,N_2312);
nor U2439 (N_2439,N_2395,N_2347);
or U2440 (N_2440,N_2359,N_2341);
nand U2441 (N_2441,N_2346,N_2303);
nand U2442 (N_2442,N_2384,N_2322);
or U2443 (N_2443,N_2398,N_2379);
or U2444 (N_2444,N_2365,N_2344);
or U2445 (N_2445,N_2381,N_2387);
and U2446 (N_2446,N_2320,N_2376);
or U2447 (N_2447,N_2361,N_2382);
nor U2448 (N_2448,N_2356,N_2335);
nor U2449 (N_2449,N_2386,N_2302);
xor U2450 (N_2450,N_2387,N_2302);
nor U2451 (N_2451,N_2376,N_2373);
and U2452 (N_2452,N_2322,N_2305);
or U2453 (N_2453,N_2309,N_2398);
xnor U2454 (N_2454,N_2300,N_2322);
or U2455 (N_2455,N_2369,N_2300);
nor U2456 (N_2456,N_2303,N_2317);
nor U2457 (N_2457,N_2354,N_2352);
nor U2458 (N_2458,N_2358,N_2303);
nand U2459 (N_2459,N_2351,N_2330);
or U2460 (N_2460,N_2372,N_2334);
nor U2461 (N_2461,N_2386,N_2309);
nand U2462 (N_2462,N_2378,N_2364);
nand U2463 (N_2463,N_2371,N_2313);
nor U2464 (N_2464,N_2323,N_2328);
and U2465 (N_2465,N_2319,N_2374);
nand U2466 (N_2466,N_2347,N_2366);
xnor U2467 (N_2467,N_2361,N_2369);
nand U2468 (N_2468,N_2399,N_2310);
nand U2469 (N_2469,N_2366,N_2334);
nor U2470 (N_2470,N_2359,N_2328);
or U2471 (N_2471,N_2317,N_2397);
or U2472 (N_2472,N_2352,N_2314);
xor U2473 (N_2473,N_2323,N_2307);
xnor U2474 (N_2474,N_2394,N_2311);
or U2475 (N_2475,N_2314,N_2355);
nor U2476 (N_2476,N_2394,N_2316);
xnor U2477 (N_2477,N_2370,N_2324);
or U2478 (N_2478,N_2370,N_2335);
nor U2479 (N_2479,N_2355,N_2358);
nor U2480 (N_2480,N_2355,N_2333);
nor U2481 (N_2481,N_2345,N_2384);
nor U2482 (N_2482,N_2334,N_2374);
and U2483 (N_2483,N_2305,N_2347);
nor U2484 (N_2484,N_2385,N_2317);
or U2485 (N_2485,N_2354,N_2397);
and U2486 (N_2486,N_2325,N_2310);
and U2487 (N_2487,N_2386,N_2344);
nand U2488 (N_2488,N_2305,N_2316);
nor U2489 (N_2489,N_2394,N_2308);
nor U2490 (N_2490,N_2392,N_2369);
and U2491 (N_2491,N_2315,N_2379);
or U2492 (N_2492,N_2377,N_2346);
nand U2493 (N_2493,N_2393,N_2366);
nor U2494 (N_2494,N_2313,N_2398);
nor U2495 (N_2495,N_2316,N_2367);
nand U2496 (N_2496,N_2364,N_2311);
and U2497 (N_2497,N_2380,N_2369);
nor U2498 (N_2498,N_2378,N_2335);
and U2499 (N_2499,N_2347,N_2311);
nor U2500 (N_2500,N_2494,N_2476);
nand U2501 (N_2501,N_2477,N_2499);
nor U2502 (N_2502,N_2446,N_2489);
nor U2503 (N_2503,N_2427,N_2420);
nor U2504 (N_2504,N_2449,N_2480);
and U2505 (N_2505,N_2414,N_2471);
or U2506 (N_2506,N_2437,N_2490);
xor U2507 (N_2507,N_2419,N_2473);
nand U2508 (N_2508,N_2497,N_2434);
and U2509 (N_2509,N_2488,N_2469);
or U2510 (N_2510,N_2412,N_2439);
nand U2511 (N_2511,N_2400,N_2428);
or U2512 (N_2512,N_2461,N_2426);
or U2513 (N_2513,N_2451,N_2424);
nand U2514 (N_2514,N_2498,N_2467);
or U2515 (N_2515,N_2452,N_2465);
and U2516 (N_2516,N_2422,N_2423);
or U2517 (N_2517,N_2453,N_2466);
nand U2518 (N_2518,N_2425,N_2450);
nand U2519 (N_2519,N_2486,N_2492);
or U2520 (N_2520,N_2493,N_2478);
or U2521 (N_2521,N_2416,N_2455);
and U2522 (N_2522,N_2447,N_2484);
nor U2523 (N_2523,N_2458,N_2482);
or U2524 (N_2524,N_2463,N_2454);
or U2525 (N_2525,N_2474,N_2448);
or U2526 (N_2526,N_2436,N_2457);
and U2527 (N_2527,N_2432,N_2460);
nor U2528 (N_2528,N_2418,N_2487);
and U2529 (N_2529,N_2408,N_2456);
or U2530 (N_2530,N_2435,N_2411);
nor U2531 (N_2531,N_2475,N_2470);
and U2532 (N_2532,N_2445,N_2462);
nor U2533 (N_2533,N_2433,N_2495);
or U2534 (N_2534,N_2440,N_2402);
nand U2535 (N_2535,N_2444,N_2443);
nand U2536 (N_2536,N_2401,N_2479);
and U2537 (N_2537,N_2415,N_2442);
nand U2538 (N_2538,N_2485,N_2429);
nand U2539 (N_2539,N_2417,N_2410);
nor U2540 (N_2540,N_2406,N_2468);
and U2541 (N_2541,N_2441,N_2496);
and U2542 (N_2542,N_2481,N_2438);
nor U2543 (N_2543,N_2405,N_2407);
xnor U2544 (N_2544,N_2409,N_2491);
nand U2545 (N_2545,N_2459,N_2483);
nand U2546 (N_2546,N_2421,N_2464);
nor U2547 (N_2547,N_2403,N_2404);
and U2548 (N_2548,N_2413,N_2430);
xnor U2549 (N_2549,N_2431,N_2472);
nor U2550 (N_2550,N_2435,N_2476);
nor U2551 (N_2551,N_2416,N_2478);
and U2552 (N_2552,N_2455,N_2418);
nor U2553 (N_2553,N_2413,N_2451);
and U2554 (N_2554,N_2466,N_2464);
nand U2555 (N_2555,N_2467,N_2436);
and U2556 (N_2556,N_2499,N_2470);
nor U2557 (N_2557,N_2442,N_2404);
xnor U2558 (N_2558,N_2456,N_2401);
nor U2559 (N_2559,N_2441,N_2407);
and U2560 (N_2560,N_2478,N_2434);
nor U2561 (N_2561,N_2437,N_2409);
and U2562 (N_2562,N_2449,N_2496);
and U2563 (N_2563,N_2403,N_2487);
nand U2564 (N_2564,N_2444,N_2465);
xor U2565 (N_2565,N_2460,N_2423);
nor U2566 (N_2566,N_2496,N_2420);
nand U2567 (N_2567,N_2406,N_2479);
or U2568 (N_2568,N_2479,N_2488);
and U2569 (N_2569,N_2420,N_2404);
nor U2570 (N_2570,N_2463,N_2442);
xor U2571 (N_2571,N_2411,N_2463);
nor U2572 (N_2572,N_2407,N_2414);
or U2573 (N_2573,N_2468,N_2444);
nand U2574 (N_2574,N_2400,N_2425);
xor U2575 (N_2575,N_2454,N_2482);
nand U2576 (N_2576,N_2494,N_2491);
nor U2577 (N_2577,N_2489,N_2449);
and U2578 (N_2578,N_2467,N_2477);
xor U2579 (N_2579,N_2441,N_2405);
nor U2580 (N_2580,N_2426,N_2412);
and U2581 (N_2581,N_2406,N_2422);
or U2582 (N_2582,N_2442,N_2423);
nor U2583 (N_2583,N_2407,N_2489);
and U2584 (N_2584,N_2404,N_2418);
nor U2585 (N_2585,N_2449,N_2458);
xnor U2586 (N_2586,N_2489,N_2445);
or U2587 (N_2587,N_2475,N_2400);
or U2588 (N_2588,N_2424,N_2474);
nor U2589 (N_2589,N_2452,N_2438);
nand U2590 (N_2590,N_2477,N_2471);
nor U2591 (N_2591,N_2481,N_2452);
or U2592 (N_2592,N_2498,N_2469);
nor U2593 (N_2593,N_2448,N_2435);
xnor U2594 (N_2594,N_2422,N_2475);
nand U2595 (N_2595,N_2410,N_2463);
xor U2596 (N_2596,N_2441,N_2423);
or U2597 (N_2597,N_2463,N_2465);
nor U2598 (N_2598,N_2408,N_2411);
and U2599 (N_2599,N_2452,N_2416);
or U2600 (N_2600,N_2539,N_2528);
or U2601 (N_2601,N_2553,N_2585);
nand U2602 (N_2602,N_2525,N_2540);
nor U2603 (N_2603,N_2591,N_2517);
nor U2604 (N_2604,N_2554,N_2588);
nand U2605 (N_2605,N_2560,N_2522);
nand U2606 (N_2606,N_2558,N_2504);
or U2607 (N_2607,N_2513,N_2567);
nand U2608 (N_2608,N_2543,N_2520);
nand U2609 (N_2609,N_2523,N_2530);
nand U2610 (N_2610,N_2555,N_2551);
nand U2611 (N_2611,N_2597,N_2536);
nor U2612 (N_2612,N_2573,N_2569);
and U2613 (N_2613,N_2589,N_2531);
or U2614 (N_2614,N_2586,N_2561);
xor U2615 (N_2615,N_2581,N_2521);
or U2616 (N_2616,N_2512,N_2549);
nand U2617 (N_2617,N_2534,N_2529);
and U2618 (N_2618,N_2565,N_2583);
nor U2619 (N_2619,N_2535,N_2584);
or U2620 (N_2620,N_2527,N_2577);
or U2621 (N_2621,N_2587,N_2545);
nand U2622 (N_2622,N_2510,N_2515);
or U2623 (N_2623,N_2500,N_2506);
and U2624 (N_2624,N_2566,N_2578);
nand U2625 (N_2625,N_2537,N_2544);
and U2626 (N_2626,N_2575,N_2593);
nor U2627 (N_2627,N_2595,N_2562);
or U2628 (N_2628,N_2598,N_2596);
xor U2629 (N_2629,N_2546,N_2574);
nand U2630 (N_2630,N_2599,N_2568);
and U2631 (N_2631,N_2563,N_2571);
and U2632 (N_2632,N_2503,N_2580);
nand U2633 (N_2633,N_2572,N_2559);
or U2634 (N_2634,N_2590,N_2548);
and U2635 (N_2635,N_2542,N_2524);
nand U2636 (N_2636,N_2547,N_2564);
nand U2637 (N_2637,N_2594,N_2518);
and U2638 (N_2638,N_2550,N_2556);
and U2639 (N_2639,N_2505,N_2532);
or U2640 (N_2640,N_2508,N_2511);
nor U2641 (N_2641,N_2557,N_2507);
nor U2642 (N_2642,N_2552,N_2509);
and U2643 (N_2643,N_2516,N_2576);
nor U2644 (N_2644,N_2541,N_2579);
or U2645 (N_2645,N_2502,N_2592);
or U2646 (N_2646,N_2526,N_2533);
and U2647 (N_2647,N_2570,N_2582);
and U2648 (N_2648,N_2514,N_2538);
nor U2649 (N_2649,N_2501,N_2519);
xor U2650 (N_2650,N_2533,N_2575);
nor U2651 (N_2651,N_2550,N_2599);
or U2652 (N_2652,N_2559,N_2599);
nor U2653 (N_2653,N_2598,N_2503);
and U2654 (N_2654,N_2565,N_2587);
nor U2655 (N_2655,N_2523,N_2515);
or U2656 (N_2656,N_2501,N_2566);
and U2657 (N_2657,N_2549,N_2520);
and U2658 (N_2658,N_2518,N_2582);
nand U2659 (N_2659,N_2525,N_2595);
nand U2660 (N_2660,N_2531,N_2588);
and U2661 (N_2661,N_2517,N_2508);
and U2662 (N_2662,N_2504,N_2539);
or U2663 (N_2663,N_2527,N_2590);
or U2664 (N_2664,N_2530,N_2519);
nor U2665 (N_2665,N_2521,N_2565);
nand U2666 (N_2666,N_2506,N_2537);
nand U2667 (N_2667,N_2552,N_2589);
nand U2668 (N_2668,N_2511,N_2542);
nor U2669 (N_2669,N_2504,N_2500);
nand U2670 (N_2670,N_2587,N_2541);
nor U2671 (N_2671,N_2566,N_2579);
xor U2672 (N_2672,N_2588,N_2545);
and U2673 (N_2673,N_2501,N_2593);
xor U2674 (N_2674,N_2549,N_2558);
or U2675 (N_2675,N_2515,N_2544);
nor U2676 (N_2676,N_2529,N_2535);
nor U2677 (N_2677,N_2577,N_2574);
and U2678 (N_2678,N_2551,N_2508);
and U2679 (N_2679,N_2591,N_2529);
nand U2680 (N_2680,N_2518,N_2584);
nor U2681 (N_2681,N_2541,N_2551);
and U2682 (N_2682,N_2574,N_2534);
xor U2683 (N_2683,N_2569,N_2536);
nor U2684 (N_2684,N_2543,N_2556);
nand U2685 (N_2685,N_2519,N_2536);
nand U2686 (N_2686,N_2547,N_2592);
nor U2687 (N_2687,N_2573,N_2571);
and U2688 (N_2688,N_2544,N_2584);
nand U2689 (N_2689,N_2587,N_2555);
nand U2690 (N_2690,N_2594,N_2508);
nor U2691 (N_2691,N_2521,N_2556);
nand U2692 (N_2692,N_2594,N_2597);
or U2693 (N_2693,N_2500,N_2531);
or U2694 (N_2694,N_2507,N_2598);
xnor U2695 (N_2695,N_2558,N_2521);
nand U2696 (N_2696,N_2501,N_2571);
and U2697 (N_2697,N_2537,N_2556);
nand U2698 (N_2698,N_2543,N_2570);
nand U2699 (N_2699,N_2575,N_2542);
or U2700 (N_2700,N_2693,N_2611);
nand U2701 (N_2701,N_2675,N_2619);
nand U2702 (N_2702,N_2610,N_2615);
nor U2703 (N_2703,N_2666,N_2600);
nand U2704 (N_2704,N_2644,N_2630);
and U2705 (N_2705,N_2638,N_2680);
or U2706 (N_2706,N_2691,N_2685);
or U2707 (N_2707,N_2616,N_2682);
or U2708 (N_2708,N_2618,N_2690);
nor U2709 (N_2709,N_2697,N_2653);
xnor U2710 (N_2710,N_2604,N_2652);
and U2711 (N_2711,N_2602,N_2614);
nor U2712 (N_2712,N_2687,N_2608);
nor U2713 (N_2713,N_2668,N_2617);
nand U2714 (N_2714,N_2674,N_2677);
nor U2715 (N_2715,N_2643,N_2692);
xor U2716 (N_2716,N_2649,N_2694);
nor U2717 (N_2717,N_2665,N_2655);
or U2718 (N_2718,N_2678,N_2622);
nand U2719 (N_2719,N_2607,N_2636);
nand U2720 (N_2720,N_2679,N_2645);
xor U2721 (N_2721,N_2683,N_2684);
or U2722 (N_2722,N_2635,N_2681);
and U2723 (N_2723,N_2613,N_2664);
and U2724 (N_2724,N_2688,N_2627);
nand U2725 (N_2725,N_2628,N_2672);
nor U2726 (N_2726,N_2612,N_2625);
nand U2727 (N_2727,N_2651,N_2632);
or U2728 (N_2728,N_2601,N_2695);
nor U2729 (N_2729,N_2661,N_2670);
nor U2730 (N_2730,N_2698,N_2641);
nor U2731 (N_2731,N_2667,N_2609);
nor U2732 (N_2732,N_2642,N_2629);
xnor U2733 (N_2733,N_2640,N_2650);
and U2734 (N_2734,N_2631,N_2634);
nand U2735 (N_2735,N_2646,N_2620);
and U2736 (N_2736,N_2657,N_2676);
or U2737 (N_2737,N_2605,N_2671);
nor U2738 (N_2738,N_2663,N_2660);
and U2739 (N_2739,N_2656,N_2686);
or U2740 (N_2740,N_2648,N_2673);
and U2741 (N_2741,N_2624,N_2669);
nand U2742 (N_2742,N_2603,N_2662);
nand U2743 (N_2743,N_2696,N_2639);
and U2744 (N_2744,N_2659,N_2699);
nor U2745 (N_2745,N_2606,N_2621);
nor U2746 (N_2746,N_2633,N_2647);
nor U2747 (N_2747,N_2654,N_2623);
nor U2748 (N_2748,N_2689,N_2658);
and U2749 (N_2749,N_2626,N_2637);
nand U2750 (N_2750,N_2629,N_2646);
or U2751 (N_2751,N_2625,N_2676);
and U2752 (N_2752,N_2621,N_2609);
or U2753 (N_2753,N_2677,N_2647);
nand U2754 (N_2754,N_2650,N_2629);
nand U2755 (N_2755,N_2634,N_2693);
and U2756 (N_2756,N_2664,N_2649);
or U2757 (N_2757,N_2688,N_2634);
or U2758 (N_2758,N_2626,N_2604);
or U2759 (N_2759,N_2628,N_2661);
or U2760 (N_2760,N_2603,N_2682);
nor U2761 (N_2761,N_2603,N_2613);
nor U2762 (N_2762,N_2635,N_2673);
xnor U2763 (N_2763,N_2603,N_2624);
xnor U2764 (N_2764,N_2666,N_2635);
nor U2765 (N_2765,N_2660,N_2603);
and U2766 (N_2766,N_2616,N_2684);
nand U2767 (N_2767,N_2627,N_2683);
nor U2768 (N_2768,N_2697,N_2690);
nand U2769 (N_2769,N_2660,N_2601);
or U2770 (N_2770,N_2651,N_2689);
nand U2771 (N_2771,N_2606,N_2631);
nand U2772 (N_2772,N_2635,N_2661);
and U2773 (N_2773,N_2608,N_2664);
and U2774 (N_2774,N_2603,N_2686);
and U2775 (N_2775,N_2684,N_2679);
and U2776 (N_2776,N_2672,N_2627);
or U2777 (N_2777,N_2689,N_2611);
or U2778 (N_2778,N_2619,N_2660);
or U2779 (N_2779,N_2624,N_2646);
and U2780 (N_2780,N_2669,N_2652);
or U2781 (N_2781,N_2669,N_2675);
nor U2782 (N_2782,N_2622,N_2682);
and U2783 (N_2783,N_2692,N_2617);
and U2784 (N_2784,N_2695,N_2651);
or U2785 (N_2785,N_2648,N_2609);
nand U2786 (N_2786,N_2669,N_2699);
nand U2787 (N_2787,N_2676,N_2604);
nand U2788 (N_2788,N_2633,N_2613);
or U2789 (N_2789,N_2688,N_2603);
nand U2790 (N_2790,N_2673,N_2689);
nor U2791 (N_2791,N_2623,N_2601);
and U2792 (N_2792,N_2605,N_2689);
nor U2793 (N_2793,N_2633,N_2621);
nand U2794 (N_2794,N_2668,N_2643);
nor U2795 (N_2795,N_2651,N_2698);
and U2796 (N_2796,N_2624,N_2692);
and U2797 (N_2797,N_2604,N_2635);
nand U2798 (N_2798,N_2640,N_2689);
xnor U2799 (N_2799,N_2697,N_2601);
nor U2800 (N_2800,N_2778,N_2783);
and U2801 (N_2801,N_2700,N_2787);
nand U2802 (N_2802,N_2791,N_2725);
and U2803 (N_2803,N_2766,N_2769);
nand U2804 (N_2804,N_2799,N_2710);
nor U2805 (N_2805,N_2711,N_2771);
or U2806 (N_2806,N_2759,N_2768);
nand U2807 (N_2807,N_2795,N_2770);
nor U2808 (N_2808,N_2788,N_2749);
nand U2809 (N_2809,N_2767,N_2798);
nand U2810 (N_2810,N_2717,N_2714);
nor U2811 (N_2811,N_2719,N_2730);
nand U2812 (N_2812,N_2774,N_2753);
xnor U2813 (N_2813,N_2723,N_2752);
nand U2814 (N_2814,N_2709,N_2748);
and U2815 (N_2815,N_2706,N_2720);
and U2816 (N_2816,N_2793,N_2764);
and U2817 (N_2817,N_2790,N_2712);
xnor U2818 (N_2818,N_2747,N_2703);
nand U2819 (N_2819,N_2781,N_2796);
nand U2820 (N_2820,N_2794,N_2718);
or U2821 (N_2821,N_2775,N_2777);
and U2822 (N_2822,N_2708,N_2702);
nand U2823 (N_2823,N_2743,N_2705);
or U2824 (N_2824,N_2754,N_2701);
xnor U2825 (N_2825,N_2761,N_2782);
nand U2826 (N_2826,N_2756,N_2744);
and U2827 (N_2827,N_2739,N_2750);
xor U2828 (N_2828,N_2751,N_2738);
nor U2829 (N_2829,N_2740,N_2762);
and U2830 (N_2830,N_2742,N_2776);
nand U2831 (N_2831,N_2780,N_2728);
nand U2832 (N_2832,N_2789,N_2735);
nand U2833 (N_2833,N_2758,N_2746);
or U2834 (N_2834,N_2732,N_2726);
or U2835 (N_2835,N_2707,N_2704);
nor U2836 (N_2836,N_2734,N_2713);
nand U2837 (N_2837,N_2716,N_2715);
xor U2838 (N_2838,N_2736,N_2729);
nand U2839 (N_2839,N_2760,N_2797);
or U2840 (N_2840,N_2733,N_2721);
nor U2841 (N_2841,N_2772,N_2786);
or U2842 (N_2842,N_2779,N_2737);
nor U2843 (N_2843,N_2773,N_2757);
and U2844 (N_2844,N_2763,N_2755);
nor U2845 (N_2845,N_2731,N_2741);
xor U2846 (N_2846,N_2724,N_2792);
nor U2847 (N_2847,N_2745,N_2727);
nand U2848 (N_2848,N_2765,N_2722);
nor U2849 (N_2849,N_2784,N_2785);
nor U2850 (N_2850,N_2769,N_2791);
or U2851 (N_2851,N_2761,N_2754);
nor U2852 (N_2852,N_2792,N_2736);
or U2853 (N_2853,N_2767,N_2768);
and U2854 (N_2854,N_2707,N_2752);
nand U2855 (N_2855,N_2736,N_2716);
nor U2856 (N_2856,N_2784,N_2735);
or U2857 (N_2857,N_2763,N_2742);
nor U2858 (N_2858,N_2768,N_2745);
and U2859 (N_2859,N_2730,N_2767);
xnor U2860 (N_2860,N_2710,N_2763);
xnor U2861 (N_2861,N_2736,N_2791);
and U2862 (N_2862,N_2716,N_2781);
nand U2863 (N_2863,N_2778,N_2714);
xor U2864 (N_2864,N_2788,N_2742);
nand U2865 (N_2865,N_2724,N_2787);
nor U2866 (N_2866,N_2768,N_2763);
nor U2867 (N_2867,N_2799,N_2791);
xnor U2868 (N_2868,N_2723,N_2760);
nor U2869 (N_2869,N_2753,N_2735);
nor U2870 (N_2870,N_2775,N_2737);
nand U2871 (N_2871,N_2735,N_2751);
nor U2872 (N_2872,N_2709,N_2730);
nand U2873 (N_2873,N_2752,N_2716);
and U2874 (N_2874,N_2700,N_2702);
nor U2875 (N_2875,N_2763,N_2756);
nand U2876 (N_2876,N_2719,N_2746);
or U2877 (N_2877,N_2747,N_2773);
nand U2878 (N_2878,N_2780,N_2724);
or U2879 (N_2879,N_2735,N_2723);
and U2880 (N_2880,N_2792,N_2706);
nand U2881 (N_2881,N_2762,N_2735);
xnor U2882 (N_2882,N_2730,N_2744);
xnor U2883 (N_2883,N_2709,N_2768);
or U2884 (N_2884,N_2718,N_2765);
xnor U2885 (N_2885,N_2777,N_2767);
nand U2886 (N_2886,N_2709,N_2741);
nor U2887 (N_2887,N_2716,N_2725);
or U2888 (N_2888,N_2785,N_2709);
or U2889 (N_2889,N_2739,N_2777);
nand U2890 (N_2890,N_2730,N_2711);
or U2891 (N_2891,N_2742,N_2766);
nor U2892 (N_2892,N_2753,N_2747);
nor U2893 (N_2893,N_2713,N_2771);
or U2894 (N_2894,N_2730,N_2759);
nor U2895 (N_2895,N_2714,N_2742);
nand U2896 (N_2896,N_2700,N_2797);
or U2897 (N_2897,N_2719,N_2760);
and U2898 (N_2898,N_2740,N_2717);
nor U2899 (N_2899,N_2792,N_2713);
nand U2900 (N_2900,N_2893,N_2842);
or U2901 (N_2901,N_2853,N_2847);
nor U2902 (N_2902,N_2852,N_2816);
nor U2903 (N_2903,N_2872,N_2851);
or U2904 (N_2904,N_2811,N_2854);
nand U2905 (N_2905,N_2849,N_2826);
and U2906 (N_2906,N_2818,N_2806);
or U2907 (N_2907,N_2877,N_2860);
nor U2908 (N_2908,N_2878,N_2824);
nand U2909 (N_2909,N_2807,N_2899);
nor U2910 (N_2910,N_2813,N_2819);
nand U2911 (N_2911,N_2812,N_2817);
nor U2912 (N_2912,N_2843,N_2839);
nor U2913 (N_2913,N_2876,N_2810);
nor U2914 (N_2914,N_2850,N_2863);
and U2915 (N_2915,N_2861,N_2882);
xnor U2916 (N_2916,N_2829,N_2848);
or U2917 (N_2917,N_2894,N_2805);
nand U2918 (N_2918,N_2822,N_2865);
xnor U2919 (N_2919,N_2840,N_2857);
nor U2920 (N_2920,N_2887,N_2823);
and U2921 (N_2921,N_2875,N_2830);
or U2922 (N_2922,N_2891,N_2800);
and U2923 (N_2923,N_2886,N_2866);
or U2924 (N_2924,N_2833,N_2888);
or U2925 (N_2925,N_2844,N_2895);
and U2926 (N_2926,N_2870,N_2867);
and U2927 (N_2927,N_2858,N_2831);
nor U2928 (N_2928,N_2873,N_2803);
or U2929 (N_2929,N_2846,N_2884);
nor U2930 (N_2930,N_2809,N_2862);
nand U2931 (N_2931,N_2856,N_2855);
nor U2932 (N_2932,N_2837,N_2836);
nor U2933 (N_2933,N_2821,N_2859);
or U2934 (N_2934,N_2880,N_2832);
or U2935 (N_2935,N_2820,N_2896);
and U2936 (N_2936,N_2890,N_2897);
and U2937 (N_2937,N_2835,N_2801);
xnor U2938 (N_2938,N_2883,N_2802);
nor U2939 (N_2939,N_2827,N_2889);
and U2940 (N_2940,N_2874,N_2881);
or U2941 (N_2941,N_2864,N_2845);
nand U2942 (N_2942,N_2898,N_2885);
and U2943 (N_2943,N_2869,N_2871);
and U2944 (N_2944,N_2868,N_2892);
xor U2945 (N_2945,N_2814,N_2808);
or U2946 (N_2946,N_2879,N_2841);
xnor U2947 (N_2947,N_2834,N_2828);
and U2948 (N_2948,N_2825,N_2815);
and U2949 (N_2949,N_2838,N_2804);
xor U2950 (N_2950,N_2833,N_2869);
or U2951 (N_2951,N_2861,N_2887);
xnor U2952 (N_2952,N_2856,N_2829);
nand U2953 (N_2953,N_2826,N_2809);
and U2954 (N_2954,N_2835,N_2883);
nand U2955 (N_2955,N_2829,N_2896);
or U2956 (N_2956,N_2858,N_2803);
or U2957 (N_2957,N_2824,N_2869);
nor U2958 (N_2958,N_2859,N_2894);
or U2959 (N_2959,N_2835,N_2807);
nor U2960 (N_2960,N_2820,N_2823);
or U2961 (N_2961,N_2805,N_2823);
and U2962 (N_2962,N_2863,N_2831);
and U2963 (N_2963,N_2859,N_2836);
nand U2964 (N_2964,N_2816,N_2865);
or U2965 (N_2965,N_2849,N_2862);
or U2966 (N_2966,N_2846,N_2863);
and U2967 (N_2967,N_2858,N_2841);
nor U2968 (N_2968,N_2884,N_2815);
nor U2969 (N_2969,N_2853,N_2897);
nor U2970 (N_2970,N_2875,N_2801);
nor U2971 (N_2971,N_2816,N_2844);
nand U2972 (N_2972,N_2888,N_2815);
nand U2973 (N_2973,N_2892,N_2826);
and U2974 (N_2974,N_2846,N_2841);
or U2975 (N_2975,N_2894,N_2843);
nor U2976 (N_2976,N_2860,N_2870);
or U2977 (N_2977,N_2860,N_2888);
and U2978 (N_2978,N_2882,N_2886);
nor U2979 (N_2979,N_2815,N_2802);
nor U2980 (N_2980,N_2804,N_2815);
or U2981 (N_2981,N_2877,N_2807);
and U2982 (N_2982,N_2814,N_2863);
nor U2983 (N_2983,N_2887,N_2868);
nand U2984 (N_2984,N_2831,N_2855);
or U2985 (N_2985,N_2860,N_2820);
and U2986 (N_2986,N_2865,N_2883);
or U2987 (N_2987,N_2845,N_2806);
nand U2988 (N_2988,N_2882,N_2863);
nor U2989 (N_2989,N_2832,N_2888);
and U2990 (N_2990,N_2850,N_2866);
nand U2991 (N_2991,N_2810,N_2858);
xor U2992 (N_2992,N_2833,N_2854);
nand U2993 (N_2993,N_2821,N_2871);
nand U2994 (N_2994,N_2862,N_2846);
or U2995 (N_2995,N_2846,N_2870);
and U2996 (N_2996,N_2833,N_2821);
and U2997 (N_2997,N_2817,N_2896);
xnor U2998 (N_2998,N_2840,N_2823);
and U2999 (N_2999,N_2862,N_2838);
and U3000 (N_3000,N_2983,N_2989);
and U3001 (N_3001,N_2946,N_2936);
or U3002 (N_3002,N_2954,N_2968);
nor U3003 (N_3003,N_2957,N_2963);
and U3004 (N_3004,N_2907,N_2950);
xor U3005 (N_3005,N_2917,N_2927);
nand U3006 (N_3006,N_2944,N_2999);
nand U3007 (N_3007,N_2928,N_2978);
nand U3008 (N_3008,N_2984,N_2960);
and U3009 (N_3009,N_2947,N_2996);
and U3010 (N_3010,N_2991,N_2921);
xor U3011 (N_3011,N_2967,N_2923);
nand U3012 (N_3012,N_2924,N_2998);
nand U3013 (N_3013,N_2945,N_2915);
xnor U3014 (N_3014,N_2911,N_2920);
xor U3015 (N_3015,N_2993,N_2912);
xor U3016 (N_3016,N_2961,N_2941);
or U3017 (N_3017,N_2901,N_2982);
nand U3018 (N_3018,N_2943,N_2974);
nor U3019 (N_3019,N_2940,N_2972);
and U3020 (N_3020,N_2900,N_2938);
and U3021 (N_3021,N_2977,N_2987);
nor U3022 (N_3022,N_2962,N_2918);
and U3023 (N_3023,N_2966,N_2990);
nand U3024 (N_3024,N_2956,N_2931);
nor U3025 (N_3025,N_2906,N_2910);
xor U3026 (N_3026,N_2970,N_2932);
nand U3027 (N_3027,N_2992,N_2958);
or U3028 (N_3028,N_2934,N_2929);
nor U3029 (N_3029,N_2976,N_2926);
and U3030 (N_3030,N_2930,N_2971);
or U3031 (N_3031,N_2988,N_2986);
nor U3032 (N_3032,N_2975,N_2953);
and U3033 (N_3033,N_2937,N_2952);
nor U3034 (N_3034,N_2965,N_2969);
or U3035 (N_3035,N_2964,N_2908);
nor U3036 (N_3036,N_2949,N_2914);
xor U3037 (N_3037,N_2905,N_2925);
and U3038 (N_3038,N_2942,N_2933);
nor U3039 (N_3039,N_2916,N_2948);
xnor U3040 (N_3040,N_2955,N_2903);
or U3041 (N_3041,N_2981,N_2935);
and U3042 (N_3042,N_2902,N_2913);
or U3043 (N_3043,N_2951,N_2995);
nand U3044 (N_3044,N_2979,N_2904);
xor U3045 (N_3045,N_2922,N_2939);
nor U3046 (N_3046,N_2997,N_2959);
and U3047 (N_3047,N_2973,N_2919);
and U3048 (N_3048,N_2980,N_2994);
or U3049 (N_3049,N_2909,N_2985);
or U3050 (N_3050,N_2949,N_2911);
nor U3051 (N_3051,N_2915,N_2982);
nand U3052 (N_3052,N_2940,N_2902);
or U3053 (N_3053,N_2921,N_2942);
and U3054 (N_3054,N_2962,N_2949);
nand U3055 (N_3055,N_2995,N_2930);
and U3056 (N_3056,N_2950,N_2914);
nor U3057 (N_3057,N_2997,N_2944);
nand U3058 (N_3058,N_2978,N_2920);
nand U3059 (N_3059,N_2926,N_2920);
xnor U3060 (N_3060,N_2929,N_2924);
nand U3061 (N_3061,N_2973,N_2994);
or U3062 (N_3062,N_2947,N_2939);
and U3063 (N_3063,N_2964,N_2961);
nand U3064 (N_3064,N_2902,N_2926);
xnor U3065 (N_3065,N_2913,N_2980);
nor U3066 (N_3066,N_2950,N_2900);
nor U3067 (N_3067,N_2982,N_2971);
nand U3068 (N_3068,N_2908,N_2921);
nand U3069 (N_3069,N_2964,N_2950);
nand U3070 (N_3070,N_2931,N_2914);
or U3071 (N_3071,N_2939,N_2911);
xnor U3072 (N_3072,N_2928,N_2979);
nand U3073 (N_3073,N_2992,N_2903);
and U3074 (N_3074,N_2977,N_2976);
or U3075 (N_3075,N_2996,N_2987);
nor U3076 (N_3076,N_2942,N_2917);
nor U3077 (N_3077,N_2906,N_2977);
nor U3078 (N_3078,N_2968,N_2997);
xor U3079 (N_3079,N_2974,N_2994);
xnor U3080 (N_3080,N_2968,N_2926);
or U3081 (N_3081,N_2903,N_2913);
and U3082 (N_3082,N_2966,N_2984);
nor U3083 (N_3083,N_2914,N_2966);
or U3084 (N_3084,N_2993,N_2943);
or U3085 (N_3085,N_2965,N_2921);
nor U3086 (N_3086,N_2975,N_2901);
xor U3087 (N_3087,N_2961,N_2939);
nand U3088 (N_3088,N_2982,N_2957);
and U3089 (N_3089,N_2982,N_2930);
and U3090 (N_3090,N_2929,N_2994);
nand U3091 (N_3091,N_2939,N_2929);
or U3092 (N_3092,N_2992,N_2980);
nand U3093 (N_3093,N_2910,N_2922);
nor U3094 (N_3094,N_2931,N_2947);
nor U3095 (N_3095,N_2979,N_2915);
xnor U3096 (N_3096,N_2906,N_2914);
xnor U3097 (N_3097,N_2992,N_2951);
or U3098 (N_3098,N_2937,N_2941);
and U3099 (N_3099,N_2928,N_2934);
nor U3100 (N_3100,N_3071,N_3031);
nor U3101 (N_3101,N_3077,N_3050);
and U3102 (N_3102,N_3063,N_3010);
nor U3103 (N_3103,N_3090,N_3009);
and U3104 (N_3104,N_3068,N_3037);
nand U3105 (N_3105,N_3016,N_3030);
and U3106 (N_3106,N_3086,N_3032);
nand U3107 (N_3107,N_3035,N_3099);
nand U3108 (N_3108,N_3093,N_3011);
or U3109 (N_3109,N_3038,N_3049);
nand U3110 (N_3110,N_3087,N_3005);
xnor U3111 (N_3111,N_3069,N_3047);
nand U3112 (N_3112,N_3008,N_3060);
nor U3113 (N_3113,N_3039,N_3024);
xnor U3114 (N_3114,N_3082,N_3085);
or U3115 (N_3115,N_3029,N_3006);
nor U3116 (N_3116,N_3021,N_3002);
nand U3117 (N_3117,N_3078,N_3084);
or U3118 (N_3118,N_3022,N_3043);
or U3119 (N_3119,N_3097,N_3000);
nand U3120 (N_3120,N_3076,N_3003);
and U3121 (N_3121,N_3052,N_3023);
or U3122 (N_3122,N_3051,N_3019);
nor U3123 (N_3123,N_3036,N_3083);
or U3124 (N_3124,N_3026,N_3057);
nor U3125 (N_3125,N_3067,N_3053);
and U3126 (N_3126,N_3095,N_3061);
nor U3127 (N_3127,N_3062,N_3013);
and U3128 (N_3128,N_3020,N_3046);
nand U3129 (N_3129,N_3080,N_3058);
or U3130 (N_3130,N_3042,N_3096);
nand U3131 (N_3131,N_3017,N_3075);
and U3132 (N_3132,N_3066,N_3041);
nand U3133 (N_3133,N_3001,N_3028);
or U3134 (N_3134,N_3088,N_3074);
nor U3135 (N_3135,N_3007,N_3064);
nand U3136 (N_3136,N_3025,N_3089);
and U3137 (N_3137,N_3054,N_3012);
and U3138 (N_3138,N_3081,N_3059);
and U3139 (N_3139,N_3072,N_3034);
nand U3140 (N_3140,N_3073,N_3092);
nor U3141 (N_3141,N_3070,N_3018);
nand U3142 (N_3142,N_3079,N_3091);
nand U3143 (N_3143,N_3044,N_3040);
xor U3144 (N_3144,N_3056,N_3015);
nor U3145 (N_3145,N_3004,N_3045);
nor U3146 (N_3146,N_3065,N_3098);
or U3147 (N_3147,N_3048,N_3055);
nor U3148 (N_3148,N_3094,N_3033);
or U3149 (N_3149,N_3027,N_3014);
or U3150 (N_3150,N_3040,N_3061);
nor U3151 (N_3151,N_3046,N_3074);
or U3152 (N_3152,N_3001,N_3008);
and U3153 (N_3153,N_3068,N_3077);
or U3154 (N_3154,N_3028,N_3083);
or U3155 (N_3155,N_3091,N_3046);
and U3156 (N_3156,N_3016,N_3006);
xor U3157 (N_3157,N_3029,N_3050);
nand U3158 (N_3158,N_3056,N_3038);
and U3159 (N_3159,N_3051,N_3041);
and U3160 (N_3160,N_3010,N_3061);
and U3161 (N_3161,N_3037,N_3088);
and U3162 (N_3162,N_3039,N_3076);
and U3163 (N_3163,N_3068,N_3009);
or U3164 (N_3164,N_3068,N_3019);
or U3165 (N_3165,N_3048,N_3010);
and U3166 (N_3166,N_3092,N_3071);
and U3167 (N_3167,N_3034,N_3022);
or U3168 (N_3168,N_3087,N_3031);
and U3169 (N_3169,N_3061,N_3009);
nand U3170 (N_3170,N_3028,N_3063);
nand U3171 (N_3171,N_3009,N_3008);
nand U3172 (N_3172,N_3077,N_3064);
nor U3173 (N_3173,N_3099,N_3095);
nand U3174 (N_3174,N_3012,N_3066);
xnor U3175 (N_3175,N_3093,N_3041);
nor U3176 (N_3176,N_3016,N_3093);
or U3177 (N_3177,N_3027,N_3029);
and U3178 (N_3178,N_3027,N_3030);
or U3179 (N_3179,N_3046,N_3005);
nor U3180 (N_3180,N_3097,N_3054);
or U3181 (N_3181,N_3018,N_3012);
xor U3182 (N_3182,N_3003,N_3000);
nand U3183 (N_3183,N_3043,N_3044);
nor U3184 (N_3184,N_3073,N_3098);
nand U3185 (N_3185,N_3029,N_3079);
nor U3186 (N_3186,N_3003,N_3096);
nor U3187 (N_3187,N_3074,N_3079);
nand U3188 (N_3188,N_3004,N_3081);
or U3189 (N_3189,N_3084,N_3090);
nand U3190 (N_3190,N_3090,N_3051);
nor U3191 (N_3191,N_3099,N_3000);
nand U3192 (N_3192,N_3030,N_3051);
and U3193 (N_3193,N_3074,N_3010);
or U3194 (N_3194,N_3013,N_3057);
nor U3195 (N_3195,N_3076,N_3048);
or U3196 (N_3196,N_3045,N_3023);
and U3197 (N_3197,N_3084,N_3086);
or U3198 (N_3198,N_3083,N_3043);
nand U3199 (N_3199,N_3095,N_3091);
or U3200 (N_3200,N_3138,N_3189);
nand U3201 (N_3201,N_3184,N_3101);
and U3202 (N_3202,N_3190,N_3130);
nand U3203 (N_3203,N_3162,N_3183);
nand U3204 (N_3204,N_3144,N_3132);
or U3205 (N_3205,N_3139,N_3124);
xor U3206 (N_3206,N_3187,N_3137);
or U3207 (N_3207,N_3142,N_3131);
nand U3208 (N_3208,N_3146,N_3178);
or U3209 (N_3209,N_3149,N_3164);
nor U3210 (N_3210,N_3182,N_3151);
nand U3211 (N_3211,N_3169,N_3143);
nor U3212 (N_3212,N_3157,N_3107);
nand U3213 (N_3213,N_3128,N_3192);
and U3214 (N_3214,N_3100,N_3109);
or U3215 (N_3215,N_3147,N_3119);
nand U3216 (N_3216,N_3129,N_3140);
and U3217 (N_3217,N_3161,N_3148);
and U3218 (N_3218,N_3134,N_3112);
and U3219 (N_3219,N_3122,N_3116);
or U3220 (N_3220,N_3176,N_3170);
and U3221 (N_3221,N_3188,N_3174);
nand U3222 (N_3222,N_3177,N_3199);
and U3223 (N_3223,N_3197,N_3154);
nor U3224 (N_3224,N_3181,N_3196);
or U3225 (N_3225,N_3121,N_3166);
nand U3226 (N_3226,N_3126,N_3167);
nand U3227 (N_3227,N_3179,N_3155);
nand U3228 (N_3228,N_3171,N_3106);
and U3229 (N_3229,N_3168,N_3103);
xor U3230 (N_3230,N_3194,N_3145);
and U3231 (N_3231,N_3123,N_3105);
or U3232 (N_3232,N_3113,N_3125);
and U3233 (N_3233,N_3195,N_3108);
nor U3234 (N_3234,N_3110,N_3120);
or U3235 (N_3235,N_3141,N_3111);
xor U3236 (N_3236,N_3173,N_3156);
nand U3237 (N_3237,N_3150,N_3104);
and U3238 (N_3238,N_3152,N_3193);
and U3239 (N_3239,N_3127,N_3160);
nand U3240 (N_3240,N_3191,N_3115);
and U3241 (N_3241,N_3135,N_3180);
nand U3242 (N_3242,N_3158,N_3172);
and U3243 (N_3243,N_3175,N_3153);
nor U3244 (N_3244,N_3133,N_3136);
and U3245 (N_3245,N_3159,N_3102);
nand U3246 (N_3246,N_3163,N_3165);
xnor U3247 (N_3247,N_3114,N_3118);
nand U3248 (N_3248,N_3186,N_3117);
or U3249 (N_3249,N_3198,N_3185);
nand U3250 (N_3250,N_3114,N_3174);
nor U3251 (N_3251,N_3132,N_3119);
and U3252 (N_3252,N_3116,N_3108);
nand U3253 (N_3253,N_3105,N_3154);
or U3254 (N_3254,N_3162,N_3148);
nor U3255 (N_3255,N_3155,N_3168);
or U3256 (N_3256,N_3100,N_3113);
and U3257 (N_3257,N_3191,N_3123);
and U3258 (N_3258,N_3173,N_3110);
nand U3259 (N_3259,N_3158,N_3170);
or U3260 (N_3260,N_3131,N_3175);
xnor U3261 (N_3261,N_3104,N_3160);
nor U3262 (N_3262,N_3150,N_3148);
nor U3263 (N_3263,N_3181,N_3106);
or U3264 (N_3264,N_3179,N_3132);
nor U3265 (N_3265,N_3154,N_3129);
and U3266 (N_3266,N_3133,N_3170);
or U3267 (N_3267,N_3138,N_3176);
and U3268 (N_3268,N_3162,N_3151);
or U3269 (N_3269,N_3125,N_3107);
or U3270 (N_3270,N_3140,N_3139);
nor U3271 (N_3271,N_3150,N_3149);
nand U3272 (N_3272,N_3184,N_3122);
nand U3273 (N_3273,N_3114,N_3138);
and U3274 (N_3274,N_3108,N_3173);
nor U3275 (N_3275,N_3188,N_3152);
nand U3276 (N_3276,N_3182,N_3173);
nor U3277 (N_3277,N_3108,N_3179);
nand U3278 (N_3278,N_3194,N_3120);
nand U3279 (N_3279,N_3144,N_3163);
or U3280 (N_3280,N_3112,N_3169);
or U3281 (N_3281,N_3156,N_3172);
or U3282 (N_3282,N_3136,N_3150);
nor U3283 (N_3283,N_3128,N_3130);
nand U3284 (N_3284,N_3129,N_3197);
or U3285 (N_3285,N_3167,N_3173);
or U3286 (N_3286,N_3153,N_3181);
and U3287 (N_3287,N_3125,N_3198);
nor U3288 (N_3288,N_3165,N_3181);
or U3289 (N_3289,N_3173,N_3188);
and U3290 (N_3290,N_3113,N_3191);
and U3291 (N_3291,N_3175,N_3151);
nand U3292 (N_3292,N_3171,N_3169);
and U3293 (N_3293,N_3177,N_3153);
and U3294 (N_3294,N_3148,N_3119);
xor U3295 (N_3295,N_3190,N_3126);
nor U3296 (N_3296,N_3143,N_3103);
and U3297 (N_3297,N_3100,N_3191);
or U3298 (N_3298,N_3147,N_3157);
nor U3299 (N_3299,N_3129,N_3150);
nor U3300 (N_3300,N_3287,N_3246);
nor U3301 (N_3301,N_3202,N_3270);
nand U3302 (N_3302,N_3205,N_3239);
or U3303 (N_3303,N_3214,N_3231);
or U3304 (N_3304,N_3242,N_3258);
nand U3305 (N_3305,N_3225,N_3211);
xor U3306 (N_3306,N_3277,N_3292);
or U3307 (N_3307,N_3235,N_3200);
or U3308 (N_3308,N_3217,N_3245);
and U3309 (N_3309,N_3250,N_3255);
nor U3310 (N_3310,N_3296,N_3268);
and U3311 (N_3311,N_3273,N_3238);
xnor U3312 (N_3312,N_3212,N_3234);
nand U3313 (N_3313,N_3271,N_3216);
or U3314 (N_3314,N_3281,N_3213);
nor U3315 (N_3315,N_3262,N_3227);
nand U3316 (N_3316,N_3233,N_3215);
xor U3317 (N_3317,N_3228,N_3229);
or U3318 (N_3318,N_3201,N_3290);
nand U3319 (N_3319,N_3264,N_3256);
or U3320 (N_3320,N_3283,N_3203);
nand U3321 (N_3321,N_3275,N_3223);
or U3322 (N_3322,N_3272,N_3279);
nand U3323 (N_3323,N_3298,N_3237);
or U3324 (N_3324,N_3222,N_3220);
and U3325 (N_3325,N_3208,N_3247);
nor U3326 (N_3326,N_3221,N_3224);
nand U3327 (N_3327,N_3266,N_3280);
or U3328 (N_3328,N_3218,N_3204);
or U3329 (N_3329,N_3226,N_3276);
or U3330 (N_3330,N_3248,N_3269);
or U3331 (N_3331,N_3282,N_3230);
nor U3332 (N_3332,N_3252,N_3254);
or U3333 (N_3333,N_3236,N_3241);
nand U3334 (N_3334,N_3206,N_3243);
or U3335 (N_3335,N_3253,N_3297);
or U3336 (N_3336,N_3285,N_3207);
and U3337 (N_3337,N_3259,N_3274);
or U3338 (N_3338,N_3265,N_3284);
nand U3339 (N_3339,N_3257,N_3291);
and U3340 (N_3340,N_3263,N_3260);
nor U3341 (N_3341,N_3286,N_3210);
nand U3342 (N_3342,N_3240,N_3293);
and U3343 (N_3343,N_3244,N_3209);
nor U3344 (N_3344,N_3288,N_3267);
and U3345 (N_3345,N_3278,N_3249);
or U3346 (N_3346,N_3251,N_3219);
and U3347 (N_3347,N_3261,N_3289);
nor U3348 (N_3348,N_3299,N_3232);
nand U3349 (N_3349,N_3294,N_3295);
nand U3350 (N_3350,N_3249,N_3208);
nand U3351 (N_3351,N_3263,N_3224);
or U3352 (N_3352,N_3206,N_3259);
nand U3353 (N_3353,N_3224,N_3243);
nand U3354 (N_3354,N_3274,N_3295);
nand U3355 (N_3355,N_3271,N_3231);
and U3356 (N_3356,N_3254,N_3291);
or U3357 (N_3357,N_3270,N_3208);
nand U3358 (N_3358,N_3284,N_3255);
nor U3359 (N_3359,N_3204,N_3264);
nor U3360 (N_3360,N_3211,N_3207);
and U3361 (N_3361,N_3250,N_3210);
nor U3362 (N_3362,N_3214,N_3299);
nand U3363 (N_3363,N_3239,N_3275);
or U3364 (N_3364,N_3273,N_3249);
or U3365 (N_3365,N_3230,N_3209);
xnor U3366 (N_3366,N_3219,N_3227);
and U3367 (N_3367,N_3228,N_3263);
nor U3368 (N_3368,N_3268,N_3272);
and U3369 (N_3369,N_3270,N_3253);
nand U3370 (N_3370,N_3253,N_3240);
nor U3371 (N_3371,N_3246,N_3241);
or U3372 (N_3372,N_3239,N_3230);
and U3373 (N_3373,N_3259,N_3219);
nor U3374 (N_3374,N_3275,N_3266);
and U3375 (N_3375,N_3261,N_3287);
nor U3376 (N_3376,N_3298,N_3219);
nand U3377 (N_3377,N_3212,N_3279);
and U3378 (N_3378,N_3282,N_3268);
nor U3379 (N_3379,N_3294,N_3243);
or U3380 (N_3380,N_3265,N_3243);
or U3381 (N_3381,N_3273,N_3274);
and U3382 (N_3382,N_3275,N_3211);
xor U3383 (N_3383,N_3241,N_3218);
nor U3384 (N_3384,N_3282,N_3269);
or U3385 (N_3385,N_3257,N_3262);
and U3386 (N_3386,N_3261,N_3284);
and U3387 (N_3387,N_3226,N_3204);
xnor U3388 (N_3388,N_3220,N_3283);
nor U3389 (N_3389,N_3268,N_3292);
xor U3390 (N_3390,N_3259,N_3291);
and U3391 (N_3391,N_3292,N_3255);
nor U3392 (N_3392,N_3200,N_3257);
nor U3393 (N_3393,N_3282,N_3271);
nor U3394 (N_3394,N_3296,N_3234);
and U3395 (N_3395,N_3269,N_3289);
nor U3396 (N_3396,N_3244,N_3228);
and U3397 (N_3397,N_3262,N_3234);
and U3398 (N_3398,N_3266,N_3258);
and U3399 (N_3399,N_3216,N_3266);
and U3400 (N_3400,N_3301,N_3375);
and U3401 (N_3401,N_3384,N_3343);
or U3402 (N_3402,N_3364,N_3338);
or U3403 (N_3403,N_3321,N_3387);
and U3404 (N_3404,N_3374,N_3334);
or U3405 (N_3405,N_3389,N_3309);
or U3406 (N_3406,N_3367,N_3383);
nor U3407 (N_3407,N_3313,N_3327);
nor U3408 (N_3408,N_3312,N_3377);
nand U3409 (N_3409,N_3380,N_3324);
nand U3410 (N_3410,N_3349,N_3303);
or U3411 (N_3411,N_3333,N_3373);
nor U3412 (N_3412,N_3385,N_3330);
xor U3413 (N_3413,N_3342,N_3351);
nand U3414 (N_3414,N_3356,N_3329);
nor U3415 (N_3415,N_3306,N_3358);
or U3416 (N_3416,N_3308,N_3350);
xor U3417 (N_3417,N_3378,N_3368);
or U3418 (N_3418,N_3369,N_3355);
xnor U3419 (N_3419,N_3386,N_3391);
and U3420 (N_3420,N_3357,N_3315);
and U3421 (N_3421,N_3360,N_3316);
nor U3422 (N_3422,N_3310,N_3344);
or U3423 (N_3423,N_3390,N_3371);
or U3424 (N_3424,N_3336,N_3388);
nand U3425 (N_3425,N_3370,N_3396);
or U3426 (N_3426,N_3323,N_3361);
or U3427 (N_3427,N_3392,N_3362);
nor U3428 (N_3428,N_3337,N_3314);
xnor U3429 (N_3429,N_3335,N_3366);
nor U3430 (N_3430,N_3372,N_3340);
nor U3431 (N_3431,N_3318,N_3331);
nand U3432 (N_3432,N_3382,N_3365);
nand U3433 (N_3433,N_3317,N_3376);
nor U3434 (N_3434,N_3363,N_3332);
and U3435 (N_3435,N_3302,N_3399);
nand U3436 (N_3436,N_3300,N_3393);
nand U3437 (N_3437,N_3320,N_3311);
nand U3438 (N_3438,N_3354,N_3339);
or U3439 (N_3439,N_3347,N_3322);
and U3440 (N_3440,N_3353,N_3304);
nand U3441 (N_3441,N_3352,N_3319);
or U3442 (N_3442,N_3359,N_3394);
and U3443 (N_3443,N_3345,N_3379);
nand U3444 (N_3444,N_3381,N_3325);
and U3445 (N_3445,N_3341,N_3305);
nor U3446 (N_3446,N_3348,N_3328);
or U3447 (N_3447,N_3346,N_3326);
nor U3448 (N_3448,N_3398,N_3397);
and U3449 (N_3449,N_3307,N_3395);
nand U3450 (N_3450,N_3331,N_3373);
and U3451 (N_3451,N_3360,N_3374);
or U3452 (N_3452,N_3304,N_3377);
nand U3453 (N_3453,N_3303,N_3346);
or U3454 (N_3454,N_3379,N_3326);
nand U3455 (N_3455,N_3364,N_3352);
xor U3456 (N_3456,N_3349,N_3394);
or U3457 (N_3457,N_3352,N_3339);
nor U3458 (N_3458,N_3308,N_3370);
or U3459 (N_3459,N_3325,N_3383);
nor U3460 (N_3460,N_3355,N_3385);
or U3461 (N_3461,N_3308,N_3368);
and U3462 (N_3462,N_3370,N_3363);
and U3463 (N_3463,N_3380,N_3335);
nand U3464 (N_3464,N_3338,N_3316);
and U3465 (N_3465,N_3303,N_3389);
nand U3466 (N_3466,N_3348,N_3369);
nand U3467 (N_3467,N_3322,N_3390);
and U3468 (N_3468,N_3361,N_3364);
and U3469 (N_3469,N_3306,N_3315);
or U3470 (N_3470,N_3332,N_3357);
and U3471 (N_3471,N_3343,N_3338);
and U3472 (N_3472,N_3384,N_3327);
nand U3473 (N_3473,N_3322,N_3358);
nor U3474 (N_3474,N_3358,N_3315);
or U3475 (N_3475,N_3371,N_3327);
and U3476 (N_3476,N_3364,N_3357);
or U3477 (N_3477,N_3374,N_3358);
or U3478 (N_3478,N_3327,N_3353);
nand U3479 (N_3479,N_3330,N_3327);
nand U3480 (N_3480,N_3363,N_3356);
xor U3481 (N_3481,N_3339,N_3327);
and U3482 (N_3482,N_3315,N_3364);
nor U3483 (N_3483,N_3316,N_3348);
nand U3484 (N_3484,N_3398,N_3355);
and U3485 (N_3485,N_3350,N_3320);
nand U3486 (N_3486,N_3371,N_3341);
xor U3487 (N_3487,N_3380,N_3341);
or U3488 (N_3488,N_3326,N_3398);
nor U3489 (N_3489,N_3337,N_3376);
and U3490 (N_3490,N_3330,N_3329);
nand U3491 (N_3491,N_3389,N_3323);
nor U3492 (N_3492,N_3321,N_3376);
nor U3493 (N_3493,N_3387,N_3343);
xor U3494 (N_3494,N_3324,N_3351);
nand U3495 (N_3495,N_3327,N_3386);
nand U3496 (N_3496,N_3382,N_3383);
xnor U3497 (N_3497,N_3364,N_3378);
or U3498 (N_3498,N_3318,N_3338);
or U3499 (N_3499,N_3389,N_3307);
or U3500 (N_3500,N_3411,N_3442);
or U3501 (N_3501,N_3487,N_3451);
or U3502 (N_3502,N_3498,N_3422);
and U3503 (N_3503,N_3445,N_3461);
nand U3504 (N_3504,N_3437,N_3429);
nand U3505 (N_3505,N_3458,N_3465);
xor U3506 (N_3506,N_3462,N_3405);
nor U3507 (N_3507,N_3443,N_3435);
or U3508 (N_3508,N_3480,N_3494);
nand U3509 (N_3509,N_3463,N_3468);
or U3510 (N_3510,N_3496,N_3459);
or U3511 (N_3511,N_3402,N_3428);
and U3512 (N_3512,N_3434,N_3491);
nand U3513 (N_3513,N_3441,N_3452);
and U3514 (N_3514,N_3479,N_3436);
nor U3515 (N_3515,N_3489,N_3419);
nand U3516 (N_3516,N_3406,N_3495);
and U3517 (N_3517,N_3433,N_3432);
nor U3518 (N_3518,N_3425,N_3497);
or U3519 (N_3519,N_3440,N_3414);
nand U3520 (N_3520,N_3424,N_3412);
nand U3521 (N_3521,N_3460,N_3403);
or U3522 (N_3522,N_3482,N_3488);
nor U3523 (N_3523,N_3477,N_3475);
or U3524 (N_3524,N_3447,N_3400);
nand U3525 (N_3525,N_3464,N_3448);
nor U3526 (N_3526,N_3455,N_3420);
xnor U3527 (N_3527,N_3430,N_3431);
nand U3528 (N_3528,N_3421,N_3439);
or U3529 (N_3529,N_3444,N_3410);
and U3530 (N_3530,N_3418,N_3457);
nand U3531 (N_3531,N_3416,N_3415);
and U3532 (N_3532,N_3454,N_3483);
or U3533 (N_3533,N_3453,N_3404);
and U3534 (N_3534,N_3490,N_3469);
and U3535 (N_3535,N_3466,N_3481);
nand U3536 (N_3536,N_3478,N_3438);
and U3537 (N_3537,N_3471,N_3409);
and U3538 (N_3538,N_3401,N_3423);
xnor U3539 (N_3539,N_3470,N_3456);
and U3540 (N_3540,N_3417,N_3485);
nand U3541 (N_3541,N_3413,N_3473);
nor U3542 (N_3542,N_3407,N_3499);
nor U3543 (N_3543,N_3408,N_3484);
nand U3544 (N_3544,N_3450,N_3472);
or U3545 (N_3545,N_3467,N_3474);
nand U3546 (N_3546,N_3476,N_3449);
and U3547 (N_3547,N_3486,N_3493);
nor U3548 (N_3548,N_3427,N_3492);
and U3549 (N_3549,N_3426,N_3446);
nand U3550 (N_3550,N_3448,N_3470);
and U3551 (N_3551,N_3439,N_3497);
xor U3552 (N_3552,N_3441,N_3450);
nand U3553 (N_3553,N_3423,N_3479);
nand U3554 (N_3554,N_3407,N_3430);
nand U3555 (N_3555,N_3470,N_3426);
or U3556 (N_3556,N_3498,N_3465);
and U3557 (N_3557,N_3455,N_3422);
or U3558 (N_3558,N_3443,N_3415);
nor U3559 (N_3559,N_3480,N_3418);
nand U3560 (N_3560,N_3408,N_3482);
nor U3561 (N_3561,N_3448,N_3486);
nand U3562 (N_3562,N_3490,N_3430);
nor U3563 (N_3563,N_3472,N_3455);
and U3564 (N_3564,N_3435,N_3492);
or U3565 (N_3565,N_3409,N_3490);
nand U3566 (N_3566,N_3479,N_3453);
and U3567 (N_3567,N_3455,N_3476);
or U3568 (N_3568,N_3463,N_3430);
nor U3569 (N_3569,N_3429,N_3461);
or U3570 (N_3570,N_3418,N_3444);
and U3571 (N_3571,N_3422,N_3402);
nor U3572 (N_3572,N_3402,N_3412);
or U3573 (N_3573,N_3491,N_3468);
nand U3574 (N_3574,N_3410,N_3452);
and U3575 (N_3575,N_3494,N_3435);
nor U3576 (N_3576,N_3464,N_3443);
xor U3577 (N_3577,N_3469,N_3483);
xnor U3578 (N_3578,N_3435,N_3429);
nor U3579 (N_3579,N_3436,N_3462);
xor U3580 (N_3580,N_3430,N_3496);
nand U3581 (N_3581,N_3451,N_3431);
or U3582 (N_3582,N_3470,N_3433);
and U3583 (N_3583,N_3449,N_3430);
and U3584 (N_3584,N_3409,N_3481);
and U3585 (N_3585,N_3434,N_3417);
nor U3586 (N_3586,N_3412,N_3464);
or U3587 (N_3587,N_3407,N_3478);
nand U3588 (N_3588,N_3460,N_3489);
xor U3589 (N_3589,N_3480,N_3433);
nor U3590 (N_3590,N_3494,N_3405);
xnor U3591 (N_3591,N_3473,N_3412);
xnor U3592 (N_3592,N_3460,N_3449);
or U3593 (N_3593,N_3412,N_3475);
nand U3594 (N_3594,N_3409,N_3404);
nor U3595 (N_3595,N_3484,N_3413);
nor U3596 (N_3596,N_3419,N_3496);
nor U3597 (N_3597,N_3454,N_3458);
nor U3598 (N_3598,N_3463,N_3441);
or U3599 (N_3599,N_3477,N_3441);
xor U3600 (N_3600,N_3521,N_3575);
nor U3601 (N_3601,N_3503,N_3540);
xor U3602 (N_3602,N_3566,N_3576);
and U3603 (N_3603,N_3595,N_3517);
nor U3604 (N_3604,N_3586,N_3594);
and U3605 (N_3605,N_3536,N_3581);
nand U3606 (N_3606,N_3550,N_3545);
nor U3607 (N_3607,N_3562,N_3542);
nand U3608 (N_3608,N_3515,N_3578);
and U3609 (N_3609,N_3500,N_3599);
and U3610 (N_3610,N_3524,N_3559);
and U3611 (N_3611,N_3563,N_3585);
or U3612 (N_3612,N_3546,N_3557);
nand U3613 (N_3613,N_3551,N_3547);
nor U3614 (N_3614,N_3590,N_3506);
and U3615 (N_3615,N_3597,N_3577);
or U3616 (N_3616,N_3514,N_3548);
and U3617 (N_3617,N_3570,N_3573);
nor U3618 (N_3618,N_3504,N_3520);
or U3619 (N_3619,N_3582,N_3560);
or U3620 (N_3620,N_3502,N_3593);
or U3621 (N_3621,N_3583,N_3564);
nand U3622 (N_3622,N_3516,N_3537);
nor U3623 (N_3623,N_3589,N_3509);
nor U3624 (N_3624,N_3529,N_3567);
nand U3625 (N_3625,N_3588,N_3584);
or U3626 (N_3626,N_3526,N_3534);
xnor U3627 (N_3627,N_3569,N_3555);
nand U3628 (N_3628,N_3553,N_3531);
nand U3629 (N_3629,N_3571,N_3544);
or U3630 (N_3630,N_3541,N_3512);
or U3631 (N_3631,N_3530,N_3532);
nor U3632 (N_3632,N_3510,N_3525);
or U3633 (N_3633,N_3508,N_3527);
nand U3634 (N_3634,N_3568,N_3572);
nand U3635 (N_3635,N_3556,N_3511);
nor U3636 (N_3636,N_3587,N_3574);
or U3637 (N_3637,N_3507,N_3596);
and U3638 (N_3638,N_3539,N_3501);
nor U3639 (N_3639,N_3535,N_3579);
and U3640 (N_3640,N_3561,N_3519);
nand U3641 (N_3641,N_3522,N_3554);
nor U3642 (N_3642,N_3543,N_3552);
nand U3643 (N_3643,N_3598,N_3558);
and U3644 (N_3644,N_3513,N_3591);
xnor U3645 (N_3645,N_3528,N_3538);
nand U3646 (N_3646,N_3580,N_3518);
and U3647 (N_3647,N_3592,N_3523);
or U3648 (N_3648,N_3549,N_3505);
nor U3649 (N_3649,N_3533,N_3565);
or U3650 (N_3650,N_3527,N_3552);
and U3651 (N_3651,N_3504,N_3595);
or U3652 (N_3652,N_3562,N_3529);
nand U3653 (N_3653,N_3597,N_3513);
and U3654 (N_3654,N_3581,N_3582);
and U3655 (N_3655,N_3579,N_3524);
nor U3656 (N_3656,N_3573,N_3578);
nand U3657 (N_3657,N_3566,N_3572);
or U3658 (N_3658,N_3534,N_3569);
nand U3659 (N_3659,N_3507,N_3542);
and U3660 (N_3660,N_3540,N_3505);
or U3661 (N_3661,N_3528,N_3561);
nor U3662 (N_3662,N_3542,N_3524);
and U3663 (N_3663,N_3595,N_3528);
nor U3664 (N_3664,N_3585,N_3537);
nand U3665 (N_3665,N_3566,N_3584);
nand U3666 (N_3666,N_3539,N_3557);
nand U3667 (N_3667,N_3506,N_3562);
nand U3668 (N_3668,N_3546,N_3578);
nor U3669 (N_3669,N_3587,N_3573);
xnor U3670 (N_3670,N_3527,N_3578);
nand U3671 (N_3671,N_3505,N_3518);
or U3672 (N_3672,N_3563,N_3516);
nor U3673 (N_3673,N_3597,N_3582);
nor U3674 (N_3674,N_3567,N_3573);
and U3675 (N_3675,N_3574,N_3528);
or U3676 (N_3676,N_3569,N_3541);
nor U3677 (N_3677,N_3595,N_3549);
and U3678 (N_3678,N_3587,N_3561);
or U3679 (N_3679,N_3570,N_3546);
and U3680 (N_3680,N_3532,N_3587);
and U3681 (N_3681,N_3550,N_3564);
and U3682 (N_3682,N_3560,N_3544);
nand U3683 (N_3683,N_3571,N_3586);
or U3684 (N_3684,N_3543,N_3513);
nor U3685 (N_3685,N_3559,N_3553);
or U3686 (N_3686,N_3559,N_3503);
or U3687 (N_3687,N_3541,N_3530);
or U3688 (N_3688,N_3566,N_3525);
xnor U3689 (N_3689,N_3571,N_3517);
and U3690 (N_3690,N_3583,N_3588);
xor U3691 (N_3691,N_3540,N_3514);
or U3692 (N_3692,N_3526,N_3584);
xor U3693 (N_3693,N_3541,N_3555);
nand U3694 (N_3694,N_3590,N_3503);
nor U3695 (N_3695,N_3529,N_3592);
or U3696 (N_3696,N_3535,N_3569);
nor U3697 (N_3697,N_3520,N_3546);
and U3698 (N_3698,N_3596,N_3554);
nand U3699 (N_3699,N_3592,N_3589);
nor U3700 (N_3700,N_3603,N_3606);
or U3701 (N_3701,N_3652,N_3614);
or U3702 (N_3702,N_3630,N_3669);
and U3703 (N_3703,N_3696,N_3633);
and U3704 (N_3704,N_3667,N_3659);
xor U3705 (N_3705,N_3656,N_3651);
nand U3706 (N_3706,N_3625,N_3657);
and U3707 (N_3707,N_3671,N_3681);
xor U3708 (N_3708,N_3695,N_3686);
nand U3709 (N_3709,N_3672,N_3626);
and U3710 (N_3710,N_3661,N_3632);
nor U3711 (N_3711,N_3654,N_3668);
and U3712 (N_3712,N_3638,N_3688);
and U3713 (N_3713,N_3660,N_3604);
nand U3714 (N_3714,N_3655,N_3665);
nand U3715 (N_3715,N_3653,N_3637);
or U3716 (N_3716,N_3676,N_3624);
nor U3717 (N_3717,N_3642,N_3639);
nor U3718 (N_3718,N_3635,N_3616);
or U3719 (N_3719,N_3608,N_3699);
or U3720 (N_3720,N_3620,N_3698);
and U3721 (N_3721,N_3673,N_3693);
nand U3722 (N_3722,N_3697,N_3611);
nor U3723 (N_3723,N_3623,N_3648);
nor U3724 (N_3724,N_3627,N_3607);
xnor U3725 (N_3725,N_3684,N_3663);
nor U3726 (N_3726,N_3600,N_3615);
and U3727 (N_3727,N_3618,N_3649);
and U3728 (N_3728,N_3629,N_3644);
and U3729 (N_3729,N_3650,N_3617);
nor U3730 (N_3730,N_3646,N_3675);
or U3731 (N_3731,N_3602,N_3687);
nand U3732 (N_3732,N_3609,N_3643);
and U3733 (N_3733,N_3674,N_3645);
nand U3734 (N_3734,N_3677,N_3610);
or U3735 (N_3735,N_3692,N_3680);
xor U3736 (N_3736,N_3678,N_3694);
nand U3737 (N_3737,N_3690,N_3621);
or U3738 (N_3738,N_3640,N_3601);
and U3739 (N_3739,N_3679,N_3682);
nor U3740 (N_3740,N_3685,N_3613);
and U3741 (N_3741,N_3666,N_3664);
and U3742 (N_3742,N_3612,N_3689);
and U3743 (N_3743,N_3634,N_3658);
nand U3744 (N_3744,N_3605,N_3670);
and U3745 (N_3745,N_3647,N_3691);
nand U3746 (N_3746,N_3636,N_3662);
nor U3747 (N_3747,N_3628,N_3631);
nor U3748 (N_3748,N_3619,N_3641);
nand U3749 (N_3749,N_3622,N_3683);
nor U3750 (N_3750,N_3636,N_3697);
and U3751 (N_3751,N_3685,N_3638);
nand U3752 (N_3752,N_3675,N_3605);
and U3753 (N_3753,N_3651,N_3611);
and U3754 (N_3754,N_3605,N_3613);
or U3755 (N_3755,N_3607,N_3655);
xor U3756 (N_3756,N_3693,N_3624);
or U3757 (N_3757,N_3621,N_3627);
or U3758 (N_3758,N_3681,N_3662);
or U3759 (N_3759,N_3634,N_3645);
xor U3760 (N_3760,N_3623,N_3652);
nand U3761 (N_3761,N_3654,N_3642);
and U3762 (N_3762,N_3677,N_3690);
nor U3763 (N_3763,N_3672,N_3664);
and U3764 (N_3764,N_3649,N_3688);
nor U3765 (N_3765,N_3668,N_3639);
nor U3766 (N_3766,N_3639,N_3631);
nor U3767 (N_3767,N_3664,N_3648);
nand U3768 (N_3768,N_3639,N_3681);
and U3769 (N_3769,N_3670,N_3614);
or U3770 (N_3770,N_3666,N_3662);
or U3771 (N_3771,N_3615,N_3603);
nand U3772 (N_3772,N_3671,N_3678);
or U3773 (N_3773,N_3616,N_3697);
nand U3774 (N_3774,N_3605,N_3657);
nor U3775 (N_3775,N_3691,N_3685);
nand U3776 (N_3776,N_3695,N_3654);
or U3777 (N_3777,N_3601,N_3661);
or U3778 (N_3778,N_3621,N_3629);
and U3779 (N_3779,N_3635,N_3604);
nor U3780 (N_3780,N_3695,N_3679);
nand U3781 (N_3781,N_3696,N_3663);
and U3782 (N_3782,N_3690,N_3673);
nor U3783 (N_3783,N_3641,N_3617);
nor U3784 (N_3784,N_3615,N_3649);
nor U3785 (N_3785,N_3623,N_3678);
nand U3786 (N_3786,N_3695,N_3617);
or U3787 (N_3787,N_3612,N_3633);
nor U3788 (N_3788,N_3679,N_3614);
nand U3789 (N_3789,N_3682,N_3653);
and U3790 (N_3790,N_3668,N_3619);
xnor U3791 (N_3791,N_3691,N_3679);
nor U3792 (N_3792,N_3696,N_3674);
xnor U3793 (N_3793,N_3662,N_3651);
nor U3794 (N_3794,N_3679,N_3603);
and U3795 (N_3795,N_3623,N_3641);
or U3796 (N_3796,N_3653,N_3669);
or U3797 (N_3797,N_3674,N_3671);
or U3798 (N_3798,N_3617,N_3622);
nor U3799 (N_3799,N_3699,N_3647);
xor U3800 (N_3800,N_3789,N_3702);
and U3801 (N_3801,N_3710,N_3734);
or U3802 (N_3802,N_3740,N_3766);
and U3803 (N_3803,N_3790,N_3785);
nand U3804 (N_3804,N_3707,N_3738);
or U3805 (N_3805,N_3746,N_3720);
xnor U3806 (N_3806,N_3721,N_3757);
nand U3807 (N_3807,N_3705,N_3714);
nand U3808 (N_3808,N_3730,N_3795);
or U3809 (N_3809,N_3771,N_3731);
or U3810 (N_3810,N_3756,N_3786);
or U3811 (N_3811,N_3717,N_3778);
nand U3812 (N_3812,N_3779,N_3733);
nand U3813 (N_3813,N_3716,N_3767);
or U3814 (N_3814,N_3743,N_3781);
nand U3815 (N_3815,N_3703,N_3788);
xnor U3816 (N_3816,N_3725,N_3715);
and U3817 (N_3817,N_3706,N_3713);
xor U3818 (N_3818,N_3797,N_3732);
nor U3819 (N_3819,N_3752,N_3708);
nand U3820 (N_3820,N_3736,N_3760);
nand U3821 (N_3821,N_3700,N_3769);
or U3822 (N_3822,N_3722,N_3727);
or U3823 (N_3823,N_3765,N_3780);
nor U3824 (N_3824,N_3739,N_3745);
or U3825 (N_3825,N_3799,N_3755);
and U3826 (N_3826,N_3787,N_3753);
and U3827 (N_3827,N_3784,N_3701);
or U3828 (N_3828,N_3758,N_3773);
nor U3829 (N_3829,N_3711,N_3770);
or U3830 (N_3830,N_3793,N_3776);
or U3831 (N_3831,N_3748,N_3792);
xnor U3832 (N_3832,N_3751,N_3791);
nand U3833 (N_3833,N_3704,N_3750);
and U3834 (N_3834,N_3764,N_3723);
nor U3835 (N_3835,N_3796,N_3728);
nor U3836 (N_3836,N_3744,N_3772);
nand U3837 (N_3837,N_3763,N_3762);
and U3838 (N_3838,N_3794,N_3747);
or U3839 (N_3839,N_3798,N_3774);
and U3840 (N_3840,N_3735,N_3726);
or U3841 (N_3841,N_3777,N_3737);
or U3842 (N_3842,N_3741,N_3742);
and U3843 (N_3843,N_3719,N_3729);
or U3844 (N_3844,N_3754,N_3724);
nand U3845 (N_3845,N_3783,N_3768);
nand U3846 (N_3846,N_3775,N_3749);
nor U3847 (N_3847,N_3782,N_3718);
and U3848 (N_3848,N_3709,N_3761);
or U3849 (N_3849,N_3712,N_3759);
and U3850 (N_3850,N_3787,N_3760);
and U3851 (N_3851,N_3763,N_3752);
or U3852 (N_3852,N_3743,N_3738);
or U3853 (N_3853,N_3763,N_3731);
nand U3854 (N_3854,N_3704,N_3772);
nand U3855 (N_3855,N_3707,N_3786);
and U3856 (N_3856,N_3719,N_3780);
or U3857 (N_3857,N_3712,N_3776);
and U3858 (N_3858,N_3797,N_3729);
nor U3859 (N_3859,N_3748,N_3733);
nand U3860 (N_3860,N_3730,N_3728);
nor U3861 (N_3861,N_3752,N_3798);
or U3862 (N_3862,N_3718,N_3748);
nor U3863 (N_3863,N_3777,N_3728);
or U3864 (N_3864,N_3785,N_3700);
nand U3865 (N_3865,N_3768,N_3751);
or U3866 (N_3866,N_3711,N_3777);
and U3867 (N_3867,N_3760,N_3761);
nand U3868 (N_3868,N_3799,N_3765);
nand U3869 (N_3869,N_3721,N_3771);
nor U3870 (N_3870,N_3775,N_3763);
nand U3871 (N_3871,N_3706,N_3756);
xor U3872 (N_3872,N_3780,N_3737);
or U3873 (N_3873,N_3740,N_3727);
nor U3874 (N_3874,N_3717,N_3752);
xnor U3875 (N_3875,N_3748,N_3701);
or U3876 (N_3876,N_3798,N_3720);
nor U3877 (N_3877,N_3757,N_3728);
nor U3878 (N_3878,N_3744,N_3711);
xor U3879 (N_3879,N_3705,N_3780);
or U3880 (N_3880,N_3782,N_3776);
or U3881 (N_3881,N_3721,N_3712);
nand U3882 (N_3882,N_3795,N_3764);
xor U3883 (N_3883,N_3792,N_3782);
xnor U3884 (N_3884,N_3768,N_3752);
xor U3885 (N_3885,N_3710,N_3773);
nor U3886 (N_3886,N_3733,N_3717);
and U3887 (N_3887,N_3739,N_3740);
or U3888 (N_3888,N_3722,N_3720);
nand U3889 (N_3889,N_3712,N_3729);
and U3890 (N_3890,N_3729,N_3756);
nand U3891 (N_3891,N_3717,N_3774);
nor U3892 (N_3892,N_3776,N_3748);
nand U3893 (N_3893,N_3768,N_3797);
nand U3894 (N_3894,N_3764,N_3751);
xor U3895 (N_3895,N_3749,N_3718);
and U3896 (N_3896,N_3749,N_3770);
nand U3897 (N_3897,N_3760,N_3722);
nand U3898 (N_3898,N_3748,N_3756);
xor U3899 (N_3899,N_3790,N_3715);
nand U3900 (N_3900,N_3878,N_3885);
or U3901 (N_3901,N_3818,N_3870);
nand U3902 (N_3902,N_3865,N_3895);
and U3903 (N_3903,N_3867,N_3894);
or U3904 (N_3904,N_3873,N_3886);
and U3905 (N_3905,N_3863,N_3871);
and U3906 (N_3906,N_3826,N_3821);
or U3907 (N_3907,N_3855,N_3880);
and U3908 (N_3908,N_3875,N_3808);
nand U3909 (N_3909,N_3814,N_3819);
or U3910 (N_3910,N_3872,N_3899);
nor U3911 (N_3911,N_3858,N_3893);
and U3912 (N_3912,N_3854,N_3806);
and U3913 (N_3913,N_3844,N_3849);
nor U3914 (N_3914,N_3887,N_3862);
nor U3915 (N_3915,N_3838,N_3809);
or U3916 (N_3916,N_3846,N_3801);
nor U3917 (N_3917,N_3829,N_3824);
nand U3918 (N_3918,N_3827,N_3805);
or U3919 (N_3919,N_3845,N_3820);
and U3920 (N_3920,N_3816,N_3881);
xor U3921 (N_3921,N_3811,N_3840);
or U3922 (N_3922,N_3832,N_3892);
nor U3923 (N_3923,N_3807,N_3848);
nor U3924 (N_3924,N_3836,N_3837);
nand U3925 (N_3925,N_3891,N_3822);
or U3926 (N_3926,N_3882,N_3802);
and U3927 (N_3927,N_3884,N_3889);
or U3928 (N_3928,N_3843,N_3890);
nor U3929 (N_3929,N_3823,N_3803);
nand U3930 (N_3930,N_3861,N_3842);
xor U3931 (N_3931,N_3864,N_3813);
nand U3932 (N_3932,N_3877,N_3839);
or U3933 (N_3933,N_3874,N_3815);
xnor U3934 (N_3934,N_3850,N_3896);
nor U3935 (N_3935,N_3853,N_3847);
xor U3936 (N_3936,N_3879,N_3804);
xnor U3937 (N_3937,N_3869,N_3841);
nor U3938 (N_3938,N_3856,N_3852);
nand U3939 (N_3939,N_3897,N_3857);
nand U3940 (N_3940,N_3876,N_3851);
or U3941 (N_3941,N_3817,N_3830);
nor U3942 (N_3942,N_3834,N_3883);
or U3943 (N_3943,N_3859,N_3866);
and U3944 (N_3944,N_3825,N_3860);
or U3945 (N_3945,N_3800,N_3833);
nor U3946 (N_3946,N_3868,N_3812);
nor U3947 (N_3947,N_3888,N_3835);
nor U3948 (N_3948,N_3898,N_3831);
xor U3949 (N_3949,N_3810,N_3828);
nor U3950 (N_3950,N_3803,N_3807);
nor U3951 (N_3951,N_3869,N_3836);
nand U3952 (N_3952,N_3825,N_3881);
nor U3953 (N_3953,N_3871,N_3891);
nand U3954 (N_3954,N_3850,N_3802);
or U3955 (N_3955,N_3898,N_3874);
and U3956 (N_3956,N_3831,N_3888);
xor U3957 (N_3957,N_3861,N_3879);
or U3958 (N_3958,N_3828,N_3886);
or U3959 (N_3959,N_3884,N_3862);
nand U3960 (N_3960,N_3850,N_3814);
nand U3961 (N_3961,N_3876,N_3841);
nand U3962 (N_3962,N_3885,N_3847);
nor U3963 (N_3963,N_3854,N_3841);
nand U3964 (N_3964,N_3898,N_3865);
nor U3965 (N_3965,N_3882,N_3817);
xor U3966 (N_3966,N_3814,N_3878);
nand U3967 (N_3967,N_3854,N_3886);
xnor U3968 (N_3968,N_3854,N_3830);
nand U3969 (N_3969,N_3843,N_3834);
nor U3970 (N_3970,N_3898,N_3857);
and U3971 (N_3971,N_3848,N_3895);
nor U3972 (N_3972,N_3875,N_3869);
or U3973 (N_3973,N_3872,N_3879);
nor U3974 (N_3974,N_3885,N_3845);
xor U3975 (N_3975,N_3856,N_3829);
nor U3976 (N_3976,N_3887,N_3809);
nand U3977 (N_3977,N_3892,N_3801);
nand U3978 (N_3978,N_3808,N_3889);
or U3979 (N_3979,N_3808,N_3895);
or U3980 (N_3980,N_3872,N_3817);
nor U3981 (N_3981,N_3889,N_3812);
and U3982 (N_3982,N_3839,N_3861);
and U3983 (N_3983,N_3829,N_3869);
nor U3984 (N_3984,N_3891,N_3842);
nor U3985 (N_3985,N_3899,N_3829);
nor U3986 (N_3986,N_3804,N_3830);
or U3987 (N_3987,N_3845,N_3859);
nor U3988 (N_3988,N_3839,N_3824);
nand U3989 (N_3989,N_3853,N_3818);
nor U3990 (N_3990,N_3805,N_3868);
nand U3991 (N_3991,N_3835,N_3842);
and U3992 (N_3992,N_3886,N_3862);
nand U3993 (N_3993,N_3890,N_3820);
nand U3994 (N_3994,N_3884,N_3821);
nor U3995 (N_3995,N_3843,N_3895);
and U3996 (N_3996,N_3872,N_3833);
nand U3997 (N_3997,N_3865,N_3870);
or U3998 (N_3998,N_3837,N_3845);
and U3999 (N_3999,N_3894,N_3892);
and U4000 (N_4000,N_3919,N_3998);
or U4001 (N_4001,N_3972,N_3949);
and U4002 (N_4002,N_3965,N_3978);
nor U4003 (N_4003,N_3928,N_3964);
nand U4004 (N_4004,N_3979,N_3975);
and U4005 (N_4005,N_3980,N_3901);
nand U4006 (N_4006,N_3962,N_3973);
xor U4007 (N_4007,N_3959,N_3932);
nor U4008 (N_4008,N_3988,N_3970);
or U4009 (N_4009,N_3924,N_3927);
nor U4010 (N_4010,N_3939,N_3940);
or U4011 (N_4011,N_3957,N_3991);
nor U4012 (N_4012,N_3914,N_3907);
nand U4013 (N_4013,N_3944,N_3995);
nor U4014 (N_4014,N_3953,N_3961);
and U4015 (N_4015,N_3926,N_3909);
xnor U4016 (N_4016,N_3925,N_3967);
xnor U4017 (N_4017,N_3992,N_3951);
and U4018 (N_4018,N_3941,N_3955);
nor U4019 (N_4019,N_3915,N_3969);
nor U4020 (N_4020,N_3929,N_3997);
nand U4021 (N_4021,N_3923,N_3946);
xor U4022 (N_4022,N_3954,N_3981);
nand U4023 (N_4023,N_3963,N_3999);
nor U4024 (N_4024,N_3931,N_3920);
and U4025 (N_4025,N_3906,N_3911);
and U4026 (N_4026,N_3910,N_3982);
xor U4027 (N_4027,N_3933,N_3930);
or U4028 (N_4028,N_3987,N_3908);
and U4029 (N_4029,N_3900,N_3922);
or U4030 (N_4030,N_3971,N_3993);
nand U4031 (N_4031,N_3936,N_3983);
or U4032 (N_4032,N_3912,N_3921);
or U4033 (N_4033,N_3916,N_3977);
xnor U4034 (N_4034,N_3958,N_3942);
xnor U4035 (N_4035,N_3974,N_3948);
nor U4036 (N_4036,N_3990,N_3976);
nand U4037 (N_4037,N_3902,N_3984);
xnor U4038 (N_4038,N_3952,N_3956);
or U4039 (N_4039,N_3950,N_3918);
nor U4040 (N_4040,N_3913,N_3934);
nor U4041 (N_4041,N_3986,N_3905);
and U4042 (N_4042,N_3968,N_3938);
or U4043 (N_4043,N_3960,N_3994);
nand U4044 (N_4044,N_3903,N_3904);
and U4045 (N_4045,N_3947,N_3966);
nor U4046 (N_4046,N_3996,N_3989);
nand U4047 (N_4047,N_3945,N_3985);
nor U4048 (N_4048,N_3943,N_3917);
and U4049 (N_4049,N_3935,N_3937);
nand U4050 (N_4050,N_3972,N_3915);
or U4051 (N_4051,N_3902,N_3930);
and U4052 (N_4052,N_3965,N_3999);
xnor U4053 (N_4053,N_3961,N_3981);
nand U4054 (N_4054,N_3955,N_3943);
nor U4055 (N_4055,N_3975,N_3941);
nor U4056 (N_4056,N_3943,N_3967);
xnor U4057 (N_4057,N_3990,N_3956);
and U4058 (N_4058,N_3927,N_3993);
or U4059 (N_4059,N_3900,N_3945);
nand U4060 (N_4060,N_3974,N_3984);
and U4061 (N_4061,N_3983,N_3993);
nand U4062 (N_4062,N_3922,N_3923);
or U4063 (N_4063,N_3910,N_3940);
xnor U4064 (N_4064,N_3956,N_3989);
nand U4065 (N_4065,N_3932,N_3990);
nor U4066 (N_4066,N_3925,N_3952);
or U4067 (N_4067,N_3924,N_3906);
or U4068 (N_4068,N_3971,N_3965);
nor U4069 (N_4069,N_3902,N_3983);
nor U4070 (N_4070,N_3900,N_3948);
nand U4071 (N_4071,N_3945,N_3964);
nand U4072 (N_4072,N_3978,N_3964);
and U4073 (N_4073,N_3991,N_3905);
xnor U4074 (N_4074,N_3904,N_3925);
or U4075 (N_4075,N_3909,N_3911);
or U4076 (N_4076,N_3948,N_3960);
or U4077 (N_4077,N_3905,N_3951);
nand U4078 (N_4078,N_3981,N_3970);
nand U4079 (N_4079,N_3970,N_3998);
and U4080 (N_4080,N_3909,N_3959);
xor U4081 (N_4081,N_3992,N_3938);
or U4082 (N_4082,N_3911,N_3975);
or U4083 (N_4083,N_3989,N_3995);
or U4084 (N_4084,N_3934,N_3922);
nor U4085 (N_4085,N_3995,N_3977);
or U4086 (N_4086,N_3958,N_3926);
nand U4087 (N_4087,N_3959,N_3907);
and U4088 (N_4088,N_3916,N_3903);
nor U4089 (N_4089,N_3937,N_3980);
nand U4090 (N_4090,N_3976,N_3904);
and U4091 (N_4091,N_3971,N_3997);
nor U4092 (N_4092,N_3960,N_3969);
nand U4093 (N_4093,N_3960,N_3959);
nor U4094 (N_4094,N_3911,N_3913);
or U4095 (N_4095,N_3993,N_3979);
and U4096 (N_4096,N_3932,N_3997);
xor U4097 (N_4097,N_3919,N_3996);
xor U4098 (N_4098,N_3941,N_3931);
nand U4099 (N_4099,N_3901,N_3942);
or U4100 (N_4100,N_4051,N_4075);
and U4101 (N_4101,N_4063,N_4016);
nand U4102 (N_4102,N_4093,N_4084);
xor U4103 (N_4103,N_4028,N_4033);
or U4104 (N_4104,N_4095,N_4030);
nand U4105 (N_4105,N_4005,N_4007);
or U4106 (N_4106,N_4099,N_4059);
and U4107 (N_4107,N_4044,N_4076);
and U4108 (N_4108,N_4069,N_4024);
xor U4109 (N_4109,N_4022,N_4068);
xor U4110 (N_4110,N_4073,N_4077);
and U4111 (N_4111,N_4000,N_4055);
and U4112 (N_4112,N_4015,N_4078);
or U4113 (N_4113,N_4066,N_4090);
or U4114 (N_4114,N_4064,N_4011);
and U4115 (N_4115,N_4056,N_4074);
and U4116 (N_4116,N_4094,N_4081);
nor U4117 (N_4117,N_4083,N_4023);
nand U4118 (N_4118,N_4097,N_4003);
nand U4119 (N_4119,N_4092,N_4045);
nand U4120 (N_4120,N_4014,N_4019);
nor U4121 (N_4121,N_4043,N_4047);
nor U4122 (N_4122,N_4082,N_4067);
and U4123 (N_4123,N_4036,N_4054);
and U4124 (N_4124,N_4089,N_4088);
nand U4125 (N_4125,N_4032,N_4001);
nor U4126 (N_4126,N_4087,N_4026);
and U4127 (N_4127,N_4025,N_4070);
and U4128 (N_4128,N_4062,N_4035);
xnor U4129 (N_4129,N_4071,N_4009);
or U4130 (N_4130,N_4031,N_4039);
or U4131 (N_4131,N_4027,N_4006);
or U4132 (N_4132,N_4091,N_4029);
nor U4133 (N_4133,N_4050,N_4021);
nor U4134 (N_4134,N_4034,N_4042);
nand U4135 (N_4135,N_4098,N_4080);
nand U4136 (N_4136,N_4053,N_4013);
and U4137 (N_4137,N_4012,N_4004);
and U4138 (N_4138,N_4046,N_4085);
nand U4139 (N_4139,N_4002,N_4079);
nand U4140 (N_4140,N_4058,N_4086);
or U4141 (N_4141,N_4061,N_4017);
xor U4142 (N_4142,N_4057,N_4018);
or U4143 (N_4143,N_4048,N_4096);
xnor U4144 (N_4144,N_4040,N_4008);
nor U4145 (N_4145,N_4060,N_4065);
nand U4146 (N_4146,N_4041,N_4052);
and U4147 (N_4147,N_4020,N_4010);
or U4148 (N_4148,N_4072,N_4049);
nand U4149 (N_4149,N_4037,N_4038);
and U4150 (N_4150,N_4037,N_4030);
xor U4151 (N_4151,N_4026,N_4093);
or U4152 (N_4152,N_4071,N_4070);
xnor U4153 (N_4153,N_4089,N_4021);
nand U4154 (N_4154,N_4089,N_4006);
nand U4155 (N_4155,N_4002,N_4010);
nand U4156 (N_4156,N_4045,N_4011);
xnor U4157 (N_4157,N_4029,N_4018);
or U4158 (N_4158,N_4094,N_4044);
or U4159 (N_4159,N_4010,N_4034);
or U4160 (N_4160,N_4091,N_4063);
or U4161 (N_4161,N_4059,N_4026);
or U4162 (N_4162,N_4003,N_4099);
nor U4163 (N_4163,N_4056,N_4000);
or U4164 (N_4164,N_4040,N_4095);
or U4165 (N_4165,N_4027,N_4031);
nor U4166 (N_4166,N_4036,N_4064);
and U4167 (N_4167,N_4074,N_4090);
and U4168 (N_4168,N_4074,N_4000);
nor U4169 (N_4169,N_4055,N_4016);
nor U4170 (N_4170,N_4082,N_4099);
nor U4171 (N_4171,N_4076,N_4079);
or U4172 (N_4172,N_4012,N_4040);
nand U4173 (N_4173,N_4066,N_4092);
xnor U4174 (N_4174,N_4094,N_4058);
or U4175 (N_4175,N_4058,N_4095);
nor U4176 (N_4176,N_4079,N_4063);
and U4177 (N_4177,N_4016,N_4036);
and U4178 (N_4178,N_4097,N_4024);
xor U4179 (N_4179,N_4083,N_4004);
nand U4180 (N_4180,N_4028,N_4078);
xnor U4181 (N_4181,N_4055,N_4024);
or U4182 (N_4182,N_4034,N_4091);
and U4183 (N_4183,N_4004,N_4033);
xor U4184 (N_4184,N_4065,N_4010);
nand U4185 (N_4185,N_4072,N_4082);
nand U4186 (N_4186,N_4046,N_4069);
nand U4187 (N_4187,N_4042,N_4044);
nor U4188 (N_4188,N_4086,N_4018);
nor U4189 (N_4189,N_4013,N_4007);
nor U4190 (N_4190,N_4090,N_4022);
nor U4191 (N_4191,N_4013,N_4012);
nor U4192 (N_4192,N_4043,N_4038);
nand U4193 (N_4193,N_4016,N_4053);
xor U4194 (N_4194,N_4049,N_4006);
and U4195 (N_4195,N_4062,N_4041);
or U4196 (N_4196,N_4065,N_4004);
nand U4197 (N_4197,N_4009,N_4025);
nand U4198 (N_4198,N_4056,N_4052);
or U4199 (N_4199,N_4087,N_4036);
nand U4200 (N_4200,N_4145,N_4131);
and U4201 (N_4201,N_4149,N_4158);
and U4202 (N_4202,N_4162,N_4104);
nand U4203 (N_4203,N_4138,N_4112);
nor U4204 (N_4204,N_4178,N_4180);
or U4205 (N_4205,N_4111,N_4160);
nor U4206 (N_4206,N_4172,N_4173);
and U4207 (N_4207,N_4109,N_4197);
nand U4208 (N_4208,N_4190,N_4194);
nor U4209 (N_4209,N_4128,N_4191);
nand U4210 (N_4210,N_4116,N_4189);
and U4211 (N_4211,N_4148,N_4141);
or U4212 (N_4212,N_4139,N_4166);
or U4213 (N_4213,N_4134,N_4101);
nand U4214 (N_4214,N_4118,N_4143);
nor U4215 (N_4215,N_4151,N_4195);
nand U4216 (N_4216,N_4163,N_4103);
nor U4217 (N_4217,N_4165,N_4100);
and U4218 (N_4218,N_4115,N_4198);
and U4219 (N_4219,N_4102,N_4175);
nor U4220 (N_4220,N_4126,N_4132);
nand U4221 (N_4221,N_4129,N_4147);
or U4222 (N_4222,N_4127,N_4186);
nand U4223 (N_4223,N_4196,N_4114);
and U4224 (N_4224,N_4174,N_4154);
or U4225 (N_4225,N_4110,N_4171);
xor U4226 (N_4226,N_4193,N_4133);
and U4227 (N_4227,N_4161,N_4176);
or U4228 (N_4228,N_4188,N_4144);
nand U4229 (N_4229,N_4140,N_4168);
and U4230 (N_4230,N_4187,N_4169);
and U4231 (N_4231,N_4108,N_4177);
and U4232 (N_4232,N_4199,N_4159);
nand U4233 (N_4233,N_4182,N_4120);
xnor U4234 (N_4234,N_4105,N_4123);
or U4235 (N_4235,N_4184,N_4124);
xnor U4236 (N_4236,N_4122,N_4167);
and U4237 (N_4237,N_4150,N_4113);
xor U4238 (N_4238,N_4181,N_4117);
xnor U4239 (N_4239,N_4130,N_4106);
nor U4240 (N_4240,N_4152,N_4121);
and U4241 (N_4241,N_4183,N_4119);
nor U4242 (N_4242,N_4137,N_4153);
or U4243 (N_4243,N_4164,N_4156);
nand U4244 (N_4244,N_4179,N_4146);
or U4245 (N_4245,N_4142,N_4135);
nand U4246 (N_4246,N_4185,N_4155);
and U4247 (N_4247,N_4157,N_4170);
nor U4248 (N_4248,N_4136,N_4125);
xnor U4249 (N_4249,N_4192,N_4107);
nand U4250 (N_4250,N_4102,N_4196);
and U4251 (N_4251,N_4172,N_4197);
and U4252 (N_4252,N_4146,N_4136);
nor U4253 (N_4253,N_4111,N_4158);
nand U4254 (N_4254,N_4103,N_4110);
nand U4255 (N_4255,N_4118,N_4189);
or U4256 (N_4256,N_4131,N_4127);
nand U4257 (N_4257,N_4118,N_4172);
and U4258 (N_4258,N_4107,N_4137);
nor U4259 (N_4259,N_4133,N_4115);
nor U4260 (N_4260,N_4120,N_4115);
xnor U4261 (N_4261,N_4134,N_4164);
nor U4262 (N_4262,N_4130,N_4183);
nor U4263 (N_4263,N_4142,N_4166);
or U4264 (N_4264,N_4175,N_4192);
xnor U4265 (N_4265,N_4166,N_4110);
nand U4266 (N_4266,N_4167,N_4149);
xor U4267 (N_4267,N_4162,N_4126);
and U4268 (N_4268,N_4106,N_4178);
or U4269 (N_4269,N_4141,N_4125);
or U4270 (N_4270,N_4192,N_4157);
and U4271 (N_4271,N_4189,N_4137);
nand U4272 (N_4272,N_4199,N_4161);
and U4273 (N_4273,N_4109,N_4135);
nand U4274 (N_4274,N_4118,N_4154);
xnor U4275 (N_4275,N_4146,N_4126);
nand U4276 (N_4276,N_4168,N_4158);
or U4277 (N_4277,N_4104,N_4152);
or U4278 (N_4278,N_4169,N_4194);
and U4279 (N_4279,N_4162,N_4181);
or U4280 (N_4280,N_4187,N_4178);
nor U4281 (N_4281,N_4196,N_4163);
nand U4282 (N_4282,N_4185,N_4136);
or U4283 (N_4283,N_4174,N_4116);
or U4284 (N_4284,N_4138,N_4143);
and U4285 (N_4285,N_4114,N_4156);
and U4286 (N_4286,N_4155,N_4138);
and U4287 (N_4287,N_4147,N_4149);
or U4288 (N_4288,N_4121,N_4166);
or U4289 (N_4289,N_4131,N_4126);
nor U4290 (N_4290,N_4136,N_4164);
nor U4291 (N_4291,N_4170,N_4192);
nor U4292 (N_4292,N_4128,N_4172);
and U4293 (N_4293,N_4127,N_4155);
xnor U4294 (N_4294,N_4119,N_4117);
and U4295 (N_4295,N_4163,N_4118);
or U4296 (N_4296,N_4198,N_4141);
and U4297 (N_4297,N_4130,N_4168);
xnor U4298 (N_4298,N_4102,N_4178);
xnor U4299 (N_4299,N_4150,N_4156);
nor U4300 (N_4300,N_4204,N_4269);
and U4301 (N_4301,N_4282,N_4252);
or U4302 (N_4302,N_4226,N_4268);
nor U4303 (N_4303,N_4240,N_4202);
nand U4304 (N_4304,N_4218,N_4288);
nand U4305 (N_4305,N_4255,N_4208);
nor U4306 (N_4306,N_4250,N_4227);
nor U4307 (N_4307,N_4206,N_4287);
nand U4308 (N_4308,N_4271,N_4294);
or U4309 (N_4309,N_4216,N_4246);
and U4310 (N_4310,N_4258,N_4281);
and U4311 (N_4311,N_4290,N_4275);
and U4312 (N_4312,N_4222,N_4225);
nand U4313 (N_4313,N_4265,N_4245);
or U4314 (N_4314,N_4215,N_4297);
and U4315 (N_4315,N_4277,N_4241);
and U4316 (N_4316,N_4283,N_4223);
nor U4317 (N_4317,N_4264,N_4217);
xnor U4318 (N_4318,N_4211,N_4232);
nor U4319 (N_4319,N_4273,N_4296);
nor U4320 (N_4320,N_4298,N_4231);
nand U4321 (N_4321,N_4286,N_4209);
nand U4322 (N_4322,N_4249,N_4234);
xnor U4323 (N_4323,N_4285,N_4243);
nor U4324 (N_4324,N_4228,N_4293);
nand U4325 (N_4325,N_4205,N_4230);
nor U4326 (N_4326,N_4261,N_4262);
and U4327 (N_4327,N_4221,N_4248);
or U4328 (N_4328,N_4229,N_4214);
nor U4329 (N_4329,N_4274,N_4219);
nand U4330 (N_4330,N_4295,N_4212);
and U4331 (N_4331,N_4259,N_4236);
nor U4332 (N_4332,N_4233,N_4251);
nand U4333 (N_4333,N_4213,N_4201);
and U4334 (N_4334,N_4256,N_4276);
and U4335 (N_4335,N_4279,N_4224);
xnor U4336 (N_4336,N_4203,N_4237);
nor U4337 (N_4337,N_4270,N_4253);
nor U4338 (N_4338,N_4235,N_4267);
nand U4339 (N_4339,N_4291,N_4289);
and U4340 (N_4340,N_4278,N_4266);
or U4341 (N_4341,N_4238,N_4239);
nor U4342 (N_4342,N_4299,N_4207);
nand U4343 (N_4343,N_4210,N_4284);
nor U4344 (N_4344,N_4263,N_4220);
or U4345 (N_4345,N_4254,N_4292);
nor U4346 (N_4346,N_4272,N_4280);
or U4347 (N_4347,N_4244,N_4247);
nor U4348 (N_4348,N_4260,N_4242);
nand U4349 (N_4349,N_4257,N_4200);
and U4350 (N_4350,N_4248,N_4280);
nand U4351 (N_4351,N_4263,N_4203);
nand U4352 (N_4352,N_4257,N_4239);
nand U4353 (N_4353,N_4253,N_4289);
nor U4354 (N_4354,N_4289,N_4205);
xnor U4355 (N_4355,N_4245,N_4249);
nor U4356 (N_4356,N_4245,N_4268);
xnor U4357 (N_4357,N_4292,N_4209);
nand U4358 (N_4358,N_4250,N_4286);
nor U4359 (N_4359,N_4226,N_4253);
nor U4360 (N_4360,N_4289,N_4235);
or U4361 (N_4361,N_4208,N_4289);
or U4362 (N_4362,N_4252,N_4200);
nor U4363 (N_4363,N_4224,N_4289);
nand U4364 (N_4364,N_4240,N_4250);
or U4365 (N_4365,N_4234,N_4282);
xor U4366 (N_4366,N_4281,N_4227);
nor U4367 (N_4367,N_4215,N_4250);
nor U4368 (N_4368,N_4201,N_4218);
nand U4369 (N_4369,N_4224,N_4268);
nand U4370 (N_4370,N_4203,N_4206);
or U4371 (N_4371,N_4240,N_4234);
nor U4372 (N_4372,N_4212,N_4241);
or U4373 (N_4373,N_4273,N_4254);
nor U4374 (N_4374,N_4250,N_4205);
nor U4375 (N_4375,N_4240,N_4286);
or U4376 (N_4376,N_4233,N_4263);
or U4377 (N_4377,N_4206,N_4298);
nand U4378 (N_4378,N_4226,N_4298);
nand U4379 (N_4379,N_4225,N_4297);
or U4380 (N_4380,N_4201,N_4297);
xor U4381 (N_4381,N_4212,N_4249);
nor U4382 (N_4382,N_4265,N_4230);
nand U4383 (N_4383,N_4227,N_4233);
xnor U4384 (N_4384,N_4294,N_4242);
nor U4385 (N_4385,N_4277,N_4295);
and U4386 (N_4386,N_4283,N_4297);
or U4387 (N_4387,N_4214,N_4239);
and U4388 (N_4388,N_4253,N_4284);
and U4389 (N_4389,N_4267,N_4273);
and U4390 (N_4390,N_4222,N_4215);
and U4391 (N_4391,N_4256,N_4219);
or U4392 (N_4392,N_4255,N_4261);
and U4393 (N_4393,N_4295,N_4278);
or U4394 (N_4394,N_4287,N_4251);
or U4395 (N_4395,N_4247,N_4252);
nor U4396 (N_4396,N_4227,N_4219);
nand U4397 (N_4397,N_4249,N_4226);
nor U4398 (N_4398,N_4254,N_4271);
nor U4399 (N_4399,N_4211,N_4231);
or U4400 (N_4400,N_4331,N_4317);
nor U4401 (N_4401,N_4305,N_4389);
nor U4402 (N_4402,N_4324,N_4341);
nand U4403 (N_4403,N_4307,N_4326);
and U4404 (N_4404,N_4361,N_4381);
or U4405 (N_4405,N_4396,N_4316);
xor U4406 (N_4406,N_4335,N_4328);
and U4407 (N_4407,N_4339,N_4363);
and U4408 (N_4408,N_4332,N_4378);
or U4409 (N_4409,N_4311,N_4346);
and U4410 (N_4410,N_4382,N_4380);
and U4411 (N_4411,N_4373,N_4351);
and U4412 (N_4412,N_4372,N_4347);
and U4413 (N_4413,N_4375,N_4393);
nand U4414 (N_4414,N_4308,N_4354);
nand U4415 (N_4415,N_4333,N_4303);
xnor U4416 (N_4416,N_4336,N_4366);
xor U4417 (N_4417,N_4313,N_4370);
nand U4418 (N_4418,N_4349,N_4338);
nand U4419 (N_4419,N_4352,N_4365);
nand U4420 (N_4420,N_4379,N_4319);
nor U4421 (N_4421,N_4357,N_4399);
nand U4422 (N_4422,N_4350,N_4345);
nand U4423 (N_4423,N_4358,N_4329);
and U4424 (N_4424,N_4360,N_4356);
and U4425 (N_4425,N_4321,N_4377);
nor U4426 (N_4426,N_4355,N_4309);
nor U4427 (N_4427,N_4325,N_4302);
and U4428 (N_4428,N_4314,N_4374);
and U4429 (N_4429,N_4300,N_4304);
and U4430 (N_4430,N_4320,N_4390);
nor U4431 (N_4431,N_4383,N_4397);
or U4432 (N_4432,N_4359,N_4384);
nand U4433 (N_4433,N_4368,N_4312);
and U4434 (N_4434,N_4315,N_4392);
nand U4435 (N_4435,N_4391,N_4395);
or U4436 (N_4436,N_4306,N_4340);
nor U4437 (N_4437,N_4385,N_4369);
nand U4438 (N_4438,N_4353,N_4394);
nor U4439 (N_4439,N_4323,N_4371);
or U4440 (N_4440,N_4310,N_4327);
or U4441 (N_4441,N_4322,N_4348);
and U4442 (N_4442,N_4342,N_4386);
or U4443 (N_4443,N_4398,N_4330);
and U4444 (N_4444,N_4334,N_4344);
and U4445 (N_4445,N_4364,N_4376);
nand U4446 (N_4446,N_4343,N_4388);
nand U4447 (N_4447,N_4337,N_4362);
and U4448 (N_4448,N_4318,N_4301);
or U4449 (N_4449,N_4387,N_4367);
or U4450 (N_4450,N_4323,N_4300);
and U4451 (N_4451,N_4318,N_4339);
and U4452 (N_4452,N_4355,N_4352);
nand U4453 (N_4453,N_4396,N_4325);
nor U4454 (N_4454,N_4304,N_4388);
nand U4455 (N_4455,N_4316,N_4342);
xor U4456 (N_4456,N_4305,N_4352);
xnor U4457 (N_4457,N_4366,N_4384);
nor U4458 (N_4458,N_4331,N_4395);
or U4459 (N_4459,N_4397,N_4350);
and U4460 (N_4460,N_4344,N_4308);
or U4461 (N_4461,N_4341,N_4339);
or U4462 (N_4462,N_4391,N_4396);
and U4463 (N_4463,N_4372,N_4321);
nor U4464 (N_4464,N_4319,N_4318);
nor U4465 (N_4465,N_4363,N_4371);
nand U4466 (N_4466,N_4342,N_4392);
or U4467 (N_4467,N_4319,N_4307);
nand U4468 (N_4468,N_4364,N_4317);
nand U4469 (N_4469,N_4367,N_4383);
xnor U4470 (N_4470,N_4300,N_4341);
nor U4471 (N_4471,N_4381,N_4363);
nor U4472 (N_4472,N_4326,N_4360);
and U4473 (N_4473,N_4372,N_4332);
or U4474 (N_4474,N_4395,N_4333);
and U4475 (N_4475,N_4354,N_4338);
nor U4476 (N_4476,N_4309,N_4302);
nor U4477 (N_4477,N_4363,N_4313);
nand U4478 (N_4478,N_4392,N_4301);
nor U4479 (N_4479,N_4324,N_4359);
or U4480 (N_4480,N_4340,N_4389);
or U4481 (N_4481,N_4354,N_4337);
and U4482 (N_4482,N_4369,N_4343);
and U4483 (N_4483,N_4328,N_4330);
nand U4484 (N_4484,N_4383,N_4336);
nand U4485 (N_4485,N_4376,N_4301);
nand U4486 (N_4486,N_4326,N_4314);
or U4487 (N_4487,N_4305,N_4328);
and U4488 (N_4488,N_4347,N_4308);
xnor U4489 (N_4489,N_4314,N_4334);
xor U4490 (N_4490,N_4374,N_4351);
nand U4491 (N_4491,N_4314,N_4339);
nand U4492 (N_4492,N_4380,N_4357);
nor U4493 (N_4493,N_4326,N_4311);
nor U4494 (N_4494,N_4302,N_4353);
nor U4495 (N_4495,N_4337,N_4332);
and U4496 (N_4496,N_4383,N_4306);
or U4497 (N_4497,N_4338,N_4361);
and U4498 (N_4498,N_4373,N_4307);
and U4499 (N_4499,N_4390,N_4354);
and U4500 (N_4500,N_4498,N_4409);
xnor U4501 (N_4501,N_4454,N_4424);
xor U4502 (N_4502,N_4434,N_4456);
and U4503 (N_4503,N_4426,N_4462);
nand U4504 (N_4504,N_4473,N_4437);
nand U4505 (N_4505,N_4481,N_4489);
or U4506 (N_4506,N_4440,N_4461);
and U4507 (N_4507,N_4430,N_4482);
or U4508 (N_4508,N_4468,N_4414);
and U4509 (N_4509,N_4488,N_4421);
or U4510 (N_4510,N_4444,N_4493);
and U4511 (N_4511,N_4495,N_4439);
and U4512 (N_4512,N_4427,N_4405);
or U4513 (N_4513,N_4445,N_4433);
or U4514 (N_4514,N_4429,N_4487);
and U4515 (N_4515,N_4435,N_4447);
and U4516 (N_4516,N_4455,N_4486);
nor U4517 (N_4517,N_4404,N_4406);
and U4518 (N_4518,N_4413,N_4460);
or U4519 (N_4519,N_4419,N_4496);
or U4520 (N_4520,N_4479,N_4476);
and U4521 (N_4521,N_4446,N_4410);
xor U4522 (N_4522,N_4420,N_4449);
or U4523 (N_4523,N_4459,N_4499);
nand U4524 (N_4524,N_4497,N_4418);
or U4525 (N_4525,N_4480,N_4485);
nand U4526 (N_4526,N_4490,N_4494);
or U4527 (N_4527,N_4428,N_4450);
or U4528 (N_4528,N_4464,N_4463);
nor U4529 (N_4529,N_4458,N_4422);
and U4530 (N_4530,N_4451,N_4477);
xnor U4531 (N_4531,N_4467,N_4400);
or U4532 (N_4532,N_4432,N_4407);
or U4533 (N_4533,N_4483,N_4475);
and U4534 (N_4534,N_4416,N_4452);
nand U4535 (N_4535,N_4457,N_4425);
or U4536 (N_4536,N_4471,N_4465);
or U4537 (N_4537,N_4448,N_4478);
xor U4538 (N_4538,N_4431,N_4491);
nand U4539 (N_4539,N_4408,N_4403);
nor U4540 (N_4540,N_4466,N_4470);
nor U4541 (N_4541,N_4472,N_4442);
or U4542 (N_4542,N_4415,N_4438);
nor U4543 (N_4543,N_4492,N_4401);
nor U4544 (N_4544,N_4469,N_4484);
xor U4545 (N_4545,N_4402,N_4441);
nand U4546 (N_4546,N_4443,N_4436);
or U4547 (N_4547,N_4411,N_4453);
and U4548 (N_4548,N_4474,N_4423);
or U4549 (N_4549,N_4412,N_4417);
nor U4550 (N_4550,N_4450,N_4433);
or U4551 (N_4551,N_4427,N_4478);
nor U4552 (N_4552,N_4468,N_4489);
or U4553 (N_4553,N_4406,N_4495);
nor U4554 (N_4554,N_4412,N_4480);
or U4555 (N_4555,N_4408,N_4465);
nor U4556 (N_4556,N_4497,N_4441);
or U4557 (N_4557,N_4426,N_4408);
and U4558 (N_4558,N_4424,N_4450);
nor U4559 (N_4559,N_4436,N_4469);
nor U4560 (N_4560,N_4426,N_4429);
or U4561 (N_4561,N_4495,N_4458);
nand U4562 (N_4562,N_4405,N_4412);
nand U4563 (N_4563,N_4449,N_4412);
nand U4564 (N_4564,N_4459,N_4479);
and U4565 (N_4565,N_4492,N_4407);
nor U4566 (N_4566,N_4411,N_4410);
or U4567 (N_4567,N_4456,N_4478);
nor U4568 (N_4568,N_4460,N_4405);
nand U4569 (N_4569,N_4464,N_4475);
nor U4570 (N_4570,N_4468,N_4438);
nand U4571 (N_4571,N_4400,N_4491);
or U4572 (N_4572,N_4431,N_4408);
and U4573 (N_4573,N_4409,N_4448);
or U4574 (N_4574,N_4468,N_4430);
and U4575 (N_4575,N_4412,N_4478);
or U4576 (N_4576,N_4430,N_4493);
nand U4577 (N_4577,N_4402,N_4483);
nor U4578 (N_4578,N_4439,N_4447);
or U4579 (N_4579,N_4425,N_4466);
and U4580 (N_4580,N_4428,N_4460);
nor U4581 (N_4581,N_4415,N_4417);
nand U4582 (N_4582,N_4423,N_4455);
and U4583 (N_4583,N_4416,N_4499);
nand U4584 (N_4584,N_4401,N_4434);
nor U4585 (N_4585,N_4447,N_4497);
xnor U4586 (N_4586,N_4454,N_4420);
or U4587 (N_4587,N_4490,N_4440);
nor U4588 (N_4588,N_4457,N_4406);
nor U4589 (N_4589,N_4453,N_4488);
nor U4590 (N_4590,N_4455,N_4438);
and U4591 (N_4591,N_4460,N_4468);
nor U4592 (N_4592,N_4459,N_4462);
xnor U4593 (N_4593,N_4469,N_4449);
or U4594 (N_4594,N_4453,N_4495);
nor U4595 (N_4595,N_4454,N_4497);
nand U4596 (N_4596,N_4425,N_4406);
nand U4597 (N_4597,N_4465,N_4458);
xnor U4598 (N_4598,N_4494,N_4473);
nor U4599 (N_4599,N_4473,N_4487);
nand U4600 (N_4600,N_4531,N_4529);
nand U4601 (N_4601,N_4569,N_4578);
nand U4602 (N_4602,N_4526,N_4535);
nand U4603 (N_4603,N_4547,N_4596);
nand U4604 (N_4604,N_4552,N_4528);
nor U4605 (N_4605,N_4502,N_4509);
nand U4606 (N_4606,N_4520,N_4567);
nand U4607 (N_4607,N_4574,N_4548);
nand U4608 (N_4608,N_4522,N_4572);
and U4609 (N_4609,N_4539,N_4586);
and U4610 (N_4610,N_4500,N_4582);
nand U4611 (N_4611,N_4512,N_4564);
or U4612 (N_4612,N_4516,N_4598);
or U4613 (N_4613,N_4560,N_4518);
or U4614 (N_4614,N_4558,N_4555);
and U4615 (N_4615,N_4565,N_4562);
xnor U4616 (N_4616,N_4561,N_4514);
xnor U4617 (N_4617,N_4549,N_4517);
nand U4618 (N_4618,N_4545,N_4557);
nor U4619 (N_4619,N_4599,N_4544);
and U4620 (N_4620,N_4551,N_4550);
nand U4621 (N_4621,N_4505,N_4541);
xor U4622 (N_4622,N_4563,N_4527);
or U4623 (N_4623,N_4590,N_4534);
nor U4624 (N_4624,N_4585,N_4538);
or U4625 (N_4625,N_4537,N_4583);
or U4626 (N_4626,N_4543,N_4553);
or U4627 (N_4627,N_4595,N_4524);
nor U4628 (N_4628,N_4581,N_4597);
nand U4629 (N_4629,N_4576,N_4515);
xor U4630 (N_4630,N_4559,N_4536);
or U4631 (N_4631,N_4510,N_4521);
and U4632 (N_4632,N_4594,N_4504);
nand U4633 (N_4633,N_4570,N_4508);
or U4634 (N_4634,N_4566,N_4532);
nor U4635 (N_4635,N_4554,N_4511);
xnor U4636 (N_4636,N_4507,N_4519);
nand U4637 (N_4637,N_4556,N_4589);
or U4638 (N_4638,N_4533,N_4587);
and U4639 (N_4639,N_4540,N_4588);
nor U4640 (N_4640,N_4593,N_4568);
and U4641 (N_4641,N_4577,N_4573);
and U4642 (N_4642,N_4530,N_4506);
and U4643 (N_4643,N_4584,N_4580);
nor U4644 (N_4644,N_4542,N_4513);
or U4645 (N_4645,N_4525,N_4575);
nor U4646 (N_4646,N_4579,N_4503);
or U4647 (N_4647,N_4523,N_4591);
or U4648 (N_4648,N_4546,N_4571);
nand U4649 (N_4649,N_4592,N_4501);
or U4650 (N_4650,N_4534,N_4556);
or U4651 (N_4651,N_4558,N_4522);
nor U4652 (N_4652,N_4536,N_4546);
nor U4653 (N_4653,N_4560,N_4515);
or U4654 (N_4654,N_4568,N_4504);
nor U4655 (N_4655,N_4555,N_4525);
nor U4656 (N_4656,N_4502,N_4579);
and U4657 (N_4657,N_4584,N_4563);
and U4658 (N_4658,N_4509,N_4518);
nand U4659 (N_4659,N_4567,N_4582);
nand U4660 (N_4660,N_4559,N_4546);
nand U4661 (N_4661,N_4592,N_4595);
nand U4662 (N_4662,N_4598,N_4599);
nand U4663 (N_4663,N_4550,N_4548);
xor U4664 (N_4664,N_4519,N_4591);
or U4665 (N_4665,N_4522,N_4544);
nand U4666 (N_4666,N_4540,N_4510);
or U4667 (N_4667,N_4521,N_4573);
nand U4668 (N_4668,N_4569,N_4551);
nor U4669 (N_4669,N_4562,N_4544);
nor U4670 (N_4670,N_4510,N_4539);
nand U4671 (N_4671,N_4594,N_4593);
and U4672 (N_4672,N_4574,N_4530);
xor U4673 (N_4673,N_4554,N_4522);
or U4674 (N_4674,N_4543,N_4523);
and U4675 (N_4675,N_4507,N_4527);
nand U4676 (N_4676,N_4514,N_4512);
or U4677 (N_4677,N_4593,N_4532);
nor U4678 (N_4678,N_4534,N_4547);
nor U4679 (N_4679,N_4590,N_4559);
xor U4680 (N_4680,N_4533,N_4595);
nand U4681 (N_4681,N_4581,N_4585);
nand U4682 (N_4682,N_4572,N_4595);
or U4683 (N_4683,N_4506,N_4584);
nand U4684 (N_4684,N_4564,N_4508);
xnor U4685 (N_4685,N_4594,N_4560);
nand U4686 (N_4686,N_4593,N_4553);
or U4687 (N_4687,N_4564,N_4593);
nor U4688 (N_4688,N_4584,N_4514);
xor U4689 (N_4689,N_4546,N_4552);
nor U4690 (N_4690,N_4533,N_4525);
and U4691 (N_4691,N_4549,N_4523);
nor U4692 (N_4692,N_4522,N_4590);
nor U4693 (N_4693,N_4533,N_4537);
or U4694 (N_4694,N_4533,N_4554);
nor U4695 (N_4695,N_4573,N_4527);
nand U4696 (N_4696,N_4545,N_4595);
nor U4697 (N_4697,N_4574,N_4595);
or U4698 (N_4698,N_4597,N_4502);
and U4699 (N_4699,N_4500,N_4594);
xnor U4700 (N_4700,N_4658,N_4636);
and U4701 (N_4701,N_4679,N_4651);
and U4702 (N_4702,N_4690,N_4677);
xor U4703 (N_4703,N_4610,N_4607);
or U4704 (N_4704,N_4647,N_4631);
or U4705 (N_4705,N_4606,N_4638);
or U4706 (N_4706,N_4613,N_4650);
or U4707 (N_4707,N_4687,N_4669);
and U4708 (N_4708,N_4622,N_4642);
and U4709 (N_4709,N_4624,N_4657);
nor U4710 (N_4710,N_4614,N_4693);
nand U4711 (N_4711,N_4686,N_4692);
nor U4712 (N_4712,N_4628,N_4655);
or U4713 (N_4713,N_4629,N_4620);
nor U4714 (N_4714,N_4640,N_4649);
or U4715 (N_4715,N_4632,N_4608);
or U4716 (N_4716,N_4666,N_4619);
or U4717 (N_4717,N_4605,N_4667);
and U4718 (N_4718,N_4644,N_4695);
nand U4719 (N_4719,N_4621,N_4670);
nand U4720 (N_4720,N_4625,N_4656);
nor U4721 (N_4721,N_4671,N_4681);
or U4722 (N_4722,N_4618,N_4682);
nand U4723 (N_4723,N_4661,N_4648);
and U4724 (N_4724,N_4659,N_4639);
or U4725 (N_4725,N_4696,N_4699);
xor U4726 (N_4726,N_4623,N_4630);
xnor U4727 (N_4727,N_4665,N_4676);
xor U4728 (N_4728,N_4611,N_4685);
nand U4729 (N_4729,N_4694,N_4680);
nor U4730 (N_4730,N_4641,N_4616);
xor U4731 (N_4731,N_4654,N_4678);
and U4732 (N_4732,N_4634,N_4637);
nand U4733 (N_4733,N_4689,N_4627);
or U4734 (N_4734,N_4653,N_4664);
nor U4735 (N_4735,N_4674,N_4698);
nor U4736 (N_4736,N_4633,N_4673);
nand U4737 (N_4737,N_4609,N_4675);
or U4738 (N_4738,N_4660,N_4601);
and U4739 (N_4739,N_4645,N_4668);
and U4740 (N_4740,N_4602,N_4603);
or U4741 (N_4741,N_4646,N_4697);
and U4742 (N_4742,N_4663,N_4643);
nand U4743 (N_4743,N_4688,N_4635);
or U4744 (N_4744,N_4604,N_4612);
and U4745 (N_4745,N_4652,N_4600);
xor U4746 (N_4746,N_4691,N_4683);
or U4747 (N_4747,N_4626,N_4617);
nor U4748 (N_4748,N_4615,N_4684);
nand U4749 (N_4749,N_4672,N_4662);
or U4750 (N_4750,N_4644,N_4646);
or U4751 (N_4751,N_4633,N_4656);
nand U4752 (N_4752,N_4673,N_4660);
and U4753 (N_4753,N_4621,N_4680);
or U4754 (N_4754,N_4650,N_4630);
and U4755 (N_4755,N_4692,N_4663);
or U4756 (N_4756,N_4639,N_4638);
and U4757 (N_4757,N_4675,N_4680);
and U4758 (N_4758,N_4649,N_4621);
or U4759 (N_4759,N_4613,N_4618);
nor U4760 (N_4760,N_4635,N_4656);
xor U4761 (N_4761,N_4621,N_4687);
nand U4762 (N_4762,N_4674,N_4697);
or U4763 (N_4763,N_4667,N_4633);
nor U4764 (N_4764,N_4679,N_4671);
xor U4765 (N_4765,N_4600,N_4688);
and U4766 (N_4766,N_4648,N_4687);
xor U4767 (N_4767,N_4677,N_4658);
or U4768 (N_4768,N_4675,N_4626);
nor U4769 (N_4769,N_4637,N_4601);
or U4770 (N_4770,N_4656,N_4612);
and U4771 (N_4771,N_4601,N_4615);
nor U4772 (N_4772,N_4612,N_4632);
or U4773 (N_4773,N_4630,N_4686);
and U4774 (N_4774,N_4601,N_4646);
or U4775 (N_4775,N_4667,N_4623);
nor U4776 (N_4776,N_4613,N_4623);
nor U4777 (N_4777,N_4699,N_4651);
xnor U4778 (N_4778,N_4658,N_4629);
nand U4779 (N_4779,N_4618,N_4649);
nor U4780 (N_4780,N_4643,N_4641);
nor U4781 (N_4781,N_4662,N_4625);
and U4782 (N_4782,N_4670,N_4646);
or U4783 (N_4783,N_4686,N_4663);
nor U4784 (N_4784,N_4675,N_4677);
xor U4785 (N_4785,N_4607,N_4669);
nand U4786 (N_4786,N_4622,N_4606);
xor U4787 (N_4787,N_4677,N_4616);
xor U4788 (N_4788,N_4685,N_4619);
nand U4789 (N_4789,N_4657,N_4699);
or U4790 (N_4790,N_4685,N_4690);
nand U4791 (N_4791,N_4620,N_4692);
or U4792 (N_4792,N_4631,N_4660);
xnor U4793 (N_4793,N_4641,N_4630);
or U4794 (N_4794,N_4697,N_4698);
and U4795 (N_4795,N_4632,N_4624);
nand U4796 (N_4796,N_4696,N_4691);
nor U4797 (N_4797,N_4667,N_4698);
xnor U4798 (N_4798,N_4683,N_4607);
and U4799 (N_4799,N_4648,N_4656);
nor U4800 (N_4800,N_4726,N_4770);
nor U4801 (N_4801,N_4712,N_4753);
xor U4802 (N_4802,N_4749,N_4767);
nand U4803 (N_4803,N_4701,N_4750);
or U4804 (N_4804,N_4705,N_4708);
and U4805 (N_4805,N_4799,N_4747);
and U4806 (N_4806,N_4731,N_4702);
nand U4807 (N_4807,N_4782,N_4763);
or U4808 (N_4808,N_4758,N_4785);
and U4809 (N_4809,N_4789,N_4793);
and U4810 (N_4810,N_4716,N_4778);
or U4811 (N_4811,N_4722,N_4729);
nor U4812 (N_4812,N_4715,N_4768);
nor U4813 (N_4813,N_4703,N_4714);
nand U4814 (N_4814,N_4756,N_4786);
nand U4815 (N_4815,N_4711,N_4700);
nor U4816 (N_4816,N_4732,N_4775);
or U4817 (N_4817,N_4740,N_4704);
and U4818 (N_4818,N_4798,N_4764);
and U4819 (N_4819,N_4733,N_4779);
xnor U4820 (N_4820,N_4772,N_4706);
or U4821 (N_4821,N_4790,N_4736);
nand U4822 (N_4822,N_4718,N_4777);
or U4823 (N_4823,N_4752,N_4781);
nor U4824 (N_4824,N_4757,N_4727);
and U4825 (N_4825,N_4797,N_4773);
and U4826 (N_4826,N_4784,N_4780);
nand U4827 (N_4827,N_4751,N_4759);
nor U4828 (N_4828,N_4734,N_4719);
and U4829 (N_4829,N_4709,N_4755);
and U4830 (N_4830,N_4745,N_4730);
nor U4831 (N_4831,N_4746,N_4707);
nor U4832 (N_4832,N_4761,N_4744);
xnor U4833 (N_4833,N_4725,N_4774);
nand U4834 (N_4834,N_4796,N_4735);
nor U4835 (N_4835,N_4787,N_4760);
and U4836 (N_4836,N_4728,N_4783);
and U4837 (N_4837,N_4776,N_4737);
and U4838 (N_4838,N_4791,N_4762);
nor U4839 (N_4839,N_4792,N_4795);
nand U4840 (N_4840,N_4748,N_4713);
nand U4841 (N_4841,N_4765,N_4741);
and U4842 (N_4842,N_4738,N_4720);
or U4843 (N_4843,N_4742,N_4717);
and U4844 (N_4844,N_4739,N_4769);
or U4845 (N_4845,N_4788,N_4724);
nand U4846 (N_4846,N_4721,N_4754);
xnor U4847 (N_4847,N_4771,N_4710);
and U4848 (N_4848,N_4723,N_4743);
nor U4849 (N_4849,N_4766,N_4794);
or U4850 (N_4850,N_4784,N_4738);
or U4851 (N_4851,N_4756,N_4719);
xor U4852 (N_4852,N_4763,N_4776);
nor U4853 (N_4853,N_4799,N_4765);
nor U4854 (N_4854,N_4729,N_4720);
nand U4855 (N_4855,N_4745,N_4720);
and U4856 (N_4856,N_4702,N_4753);
xor U4857 (N_4857,N_4707,N_4713);
nand U4858 (N_4858,N_4750,N_4746);
and U4859 (N_4859,N_4779,N_4708);
and U4860 (N_4860,N_4764,N_4745);
nor U4861 (N_4861,N_4770,N_4794);
xor U4862 (N_4862,N_4768,N_4769);
nand U4863 (N_4863,N_4732,N_4796);
or U4864 (N_4864,N_4706,N_4742);
nand U4865 (N_4865,N_4797,N_4774);
nor U4866 (N_4866,N_4743,N_4763);
or U4867 (N_4867,N_4714,N_4759);
nor U4868 (N_4868,N_4772,N_4748);
nor U4869 (N_4869,N_4790,N_4796);
nand U4870 (N_4870,N_4768,N_4789);
or U4871 (N_4871,N_4731,N_4700);
nand U4872 (N_4872,N_4733,N_4758);
nand U4873 (N_4873,N_4764,N_4749);
nor U4874 (N_4874,N_4738,N_4771);
nand U4875 (N_4875,N_4711,N_4782);
and U4876 (N_4876,N_4771,N_4799);
nand U4877 (N_4877,N_4765,N_4752);
or U4878 (N_4878,N_4790,N_4792);
nand U4879 (N_4879,N_4768,N_4746);
nand U4880 (N_4880,N_4732,N_4718);
nor U4881 (N_4881,N_4712,N_4742);
nor U4882 (N_4882,N_4724,N_4787);
or U4883 (N_4883,N_4758,N_4784);
or U4884 (N_4884,N_4778,N_4721);
nor U4885 (N_4885,N_4756,N_4793);
and U4886 (N_4886,N_4708,N_4715);
or U4887 (N_4887,N_4721,N_4755);
nor U4888 (N_4888,N_4785,N_4702);
nor U4889 (N_4889,N_4753,N_4797);
xnor U4890 (N_4890,N_4711,N_4794);
and U4891 (N_4891,N_4774,N_4701);
nand U4892 (N_4892,N_4707,N_4728);
or U4893 (N_4893,N_4743,N_4734);
and U4894 (N_4894,N_4711,N_4706);
nor U4895 (N_4895,N_4708,N_4702);
nor U4896 (N_4896,N_4754,N_4764);
nor U4897 (N_4897,N_4780,N_4717);
nand U4898 (N_4898,N_4766,N_4702);
xnor U4899 (N_4899,N_4793,N_4779);
nand U4900 (N_4900,N_4808,N_4825);
or U4901 (N_4901,N_4845,N_4815);
xnor U4902 (N_4902,N_4840,N_4846);
and U4903 (N_4903,N_4874,N_4816);
or U4904 (N_4904,N_4892,N_4896);
nand U4905 (N_4905,N_4828,N_4810);
and U4906 (N_4906,N_4832,N_4823);
nor U4907 (N_4907,N_4879,N_4868);
and U4908 (N_4908,N_4889,N_4863);
and U4909 (N_4909,N_4844,N_4830);
and U4910 (N_4910,N_4897,N_4861);
and U4911 (N_4911,N_4857,N_4820);
and U4912 (N_4912,N_4847,N_4821);
nand U4913 (N_4913,N_4843,N_4859);
or U4914 (N_4914,N_4827,N_4806);
nand U4915 (N_4915,N_4875,N_4864);
or U4916 (N_4916,N_4802,N_4885);
and U4917 (N_4917,N_4814,N_4805);
and U4918 (N_4918,N_4899,N_4807);
nand U4919 (N_4919,N_4848,N_4865);
or U4920 (N_4920,N_4833,N_4831);
or U4921 (N_4921,N_4866,N_4838);
or U4922 (N_4922,N_4882,N_4886);
nand U4923 (N_4923,N_4818,N_4804);
nand U4924 (N_4924,N_4860,N_4849);
nand U4925 (N_4925,N_4851,N_4839);
or U4926 (N_4926,N_4894,N_4856);
or U4927 (N_4927,N_4883,N_4824);
nor U4928 (N_4928,N_4835,N_4855);
and U4929 (N_4929,N_4812,N_4817);
nand U4930 (N_4930,N_4853,N_4803);
nand U4931 (N_4931,N_4880,N_4854);
nor U4932 (N_4932,N_4887,N_4884);
or U4933 (N_4933,N_4822,N_4869);
or U4934 (N_4934,N_4819,N_4858);
or U4935 (N_4935,N_4890,N_4841);
and U4936 (N_4936,N_4826,N_4811);
or U4937 (N_4937,N_4813,N_4801);
nor U4938 (N_4938,N_4872,N_4837);
and U4939 (N_4939,N_4871,N_4829);
and U4940 (N_4940,N_4877,N_4881);
and U4941 (N_4941,N_4873,N_4891);
or U4942 (N_4942,N_4893,N_4834);
and U4943 (N_4943,N_4809,N_4867);
nor U4944 (N_4944,N_4878,N_4895);
nand U4945 (N_4945,N_4862,N_4876);
xor U4946 (N_4946,N_4888,N_4852);
nor U4947 (N_4947,N_4850,N_4842);
and U4948 (N_4948,N_4800,N_4870);
nor U4949 (N_4949,N_4836,N_4898);
nor U4950 (N_4950,N_4847,N_4816);
nor U4951 (N_4951,N_4889,N_4898);
nor U4952 (N_4952,N_4882,N_4853);
or U4953 (N_4953,N_4839,N_4835);
nand U4954 (N_4954,N_4870,N_4844);
and U4955 (N_4955,N_4880,N_4835);
nand U4956 (N_4956,N_4824,N_4897);
and U4957 (N_4957,N_4819,N_4851);
nand U4958 (N_4958,N_4846,N_4802);
and U4959 (N_4959,N_4846,N_4884);
or U4960 (N_4960,N_4894,N_4872);
and U4961 (N_4961,N_4863,N_4846);
nand U4962 (N_4962,N_4873,N_4806);
xor U4963 (N_4963,N_4855,N_4877);
nor U4964 (N_4964,N_4896,N_4801);
xor U4965 (N_4965,N_4810,N_4848);
and U4966 (N_4966,N_4804,N_4857);
xnor U4967 (N_4967,N_4821,N_4850);
or U4968 (N_4968,N_4819,N_4868);
nor U4969 (N_4969,N_4877,N_4836);
or U4970 (N_4970,N_4838,N_4872);
and U4971 (N_4971,N_4839,N_4872);
nor U4972 (N_4972,N_4844,N_4828);
nand U4973 (N_4973,N_4844,N_4889);
nand U4974 (N_4974,N_4854,N_4839);
or U4975 (N_4975,N_4842,N_4868);
or U4976 (N_4976,N_4859,N_4885);
or U4977 (N_4977,N_4879,N_4855);
and U4978 (N_4978,N_4825,N_4854);
or U4979 (N_4979,N_4872,N_4864);
or U4980 (N_4980,N_4816,N_4851);
or U4981 (N_4981,N_4867,N_4836);
and U4982 (N_4982,N_4814,N_4862);
nor U4983 (N_4983,N_4887,N_4811);
nand U4984 (N_4984,N_4887,N_4899);
nor U4985 (N_4985,N_4886,N_4848);
or U4986 (N_4986,N_4853,N_4883);
or U4987 (N_4987,N_4859,N_4891);
nor U4988 (N_4988,N_4891,N_4836);
or U4989 (N_4989,N_4831,N_4872);
or U4990 (N_4990,N_4875,N_4893);
or U4991 (N_4991,N_4879,N_4881);
xor U4992 (N_4992,N_4846,N_4869);
or U4993 (N_4993,N_4886,N_4822);
nor U4994 (N_4994,N_4864,N_4877);
nor U4995 (N_4995,N_4883,N_4803);
nand U4996 (N_4996,N_4813,N_4822);
or U4997 (N_4997,N_4889,N_4871);
nand U4998 (N_4998,N_4884,N_4824);
or U4999 (N_4999,N_4881,N_4851);
nand UO_0 (O_0,N_4908,N_4978);
nand UO_1 (O_1,N_4904,N_4954);
and UO_2 (O_2,N_4907,N_4952);
and UO_3 (O_3,N_4957,N_4937);
nor UO_4 (O_4,N_4985,N_4972);
nor UO_5 (O_5,N_4943,N_4991);
nand UO_6 (O_6,N_4928,N_4930);
and UO_7 (O_7,N_4909,N_4920);
nor UO_8 (O_8,N_4990,N_4905);
nor UO_9 (O_9,N_4971,N_4950);
or UO_10 (O_10,N_4984,N_4996);
xor UO_11 (O_11,N_4955,N_4913);
nor UO_12 (O_12,N_4962,N_4923);
or UO_13 (O_13,N_4924,N_4967);
or UO_14 (O_14,N_4949,N_4959);
xor UO_15 (O_15,N_4938,N_4917);
nand UO_16 (O_16,N_4914,N_4931);
nor UO_17 (O_17,N_4915,N_4941);
nand UO_18 (O_18,N_4911,N_4922);
or UO_19 (O_19,N_4994,N_4921);
xor UO_20 (O_20,N_4977,N_4983);
nor UO_21 (O_21,N_4970,N_4976);
nor UO_22 (O_22,N_4934,N_4942);
or UO_23 (O_23,N_4906,N_4956);
or UO_24 (O_24,N_4965,N_4981);
and UO_25 (O_25,N_4964,N_4963);
and UO_26 (O_26,N_4988,N_4960);
nand UO_27 (O_27,N_4980,N_4951);
nor UO_28 (O_28,N_4966,N_4900);
nand UO_29 (O_29,N_4961,N_4986);
or UO_30 (O_30,N_4929,N_4999);
or UO_31 (O_31,N_4903,N_4974);
nand UO_32 (O_32,N_4945,N_4940);
and UO_33 (O_33,N_4919,N_4947);
and UO_34 (O_34,N_4901,N_4912);
xnor UO_35 (O_35,N_4958,N_4989);
and UO_36 (O_36,N_4935,N_4979);
nand UO_37 (O_37,N_4932,N_4995);
nand UO_38 (O_38,N_4992,N_4946);
and UO_39 (O_39,N_4973,N_4993);
nor UO_40 (O_40,N_4918,N_4982);
xor UO_41 (O_41,N_4936,N_4968);
nor UO_42 (O_42,N_4910,N_4902);
or UO_43 (O_43,N_4969,N_4975);
xor UO_44 (O_44,N_4916,N_4939);
and UO_45 (O_45,N_4987,N_4926);
nor UO_46 (O_46,N_4953,N_4997);
nor UO_47 (O_47,N_4925,N_4998);
xnor UO_48 (O_48,N_4933,N_4944);
and UO_49 (O_49,N_4948,N_4927);
and UO_50 (O_50,N_4982,N_4912);
nand UO_51 (O_51,N_4900,N_4986);
nor UO_52 (O_52,N_4971,N_4962);
or UO_53 (O_53,N_4993,N_4940);
nor UO_54 (O_54,N_4963,N_4947);
nor UO_55 (O_55,N_4945,N_4958);
or UO_56 (O_56,N_4987,N_4970);
and UO_57 (O_57,N_4925,N_4978);
and UO_58 (O_58,N_4955,N_4988);
nor UO_59 (O_59,N_4910,N_4905);
nand UO_60 (O_60,N_4941,N_4937);
and UO_61 (O_61,N_4921,N_4931);
nor UO_62 (O_62,N_4977,N_4937);
and UO_63 (O_63,N_4926,N_4969);
nor UO_64 (O_64,N_4906,N_4933);
or UO_65 (O_65,N_4915,N_4983);
nor UO_66 (O_66,N_4908,N_4949);
nand UO_67 (O_67,N_4900,N_4953);
and UO_68 (O_68,N_4934,N_4901);
xnor UO_69 (O_69,N_4982,N_4919);
nand UO_70 (O_70,N_4973,N_4980);
or UO_71 (O_71,N_4918,N_4995);
nand UO_72 (O_72,N_4928,N_4948);
or UO_73 (O_73,N_4908,N_4917);
nand UO_74 (O_74,N_4993,N_4980);
nor UO_75 (O_75,N_4988,N_4927);
nor UO_76 (O_76,N_4970,N_4983);
nor UO_77 (O_77,N_4913,N_4979);
xnor UO_78 (O_78,N_4989,N_4966);
and UO_79 (O_79,N_4985,N_4951);
xnor UO_80 (O_80,N_4934,N_4960);
or UO_81 (O_81,N_4925,N_4912);
and UO_82 (O_82,N_4944,N_4965);
and UO_83 (O_83,N_4995,N_4978);
and UO_84 (O_84,N_4991,N_4940);
or UO_85 (O_85,N_4909,N_4905);
or UO_86 (O_86,N_4950,N_4955);
and UO_87 (O_87,N_4960,N_4952);
and UO_88 (O_88,N_4928,N_4976);
nand UO_89 (O_89,N_4954,N_4903);
and UO_90 (O_90,N_4963,N_4988);
xor UO_91 (O_91,N_4978,N_4909);
nand UO_92 (O_92,N_4940,N_4972);
nand UO_93 (O_93,N_4920,N_4902);
nor UO_94 (O_94,N_4900,N_4943);
xor UO_95 (O_95,N_4986,N_4913);
nand UO_96 (O_96,N_4980,N_4974);
xor UO_97 (O_97,N_4970,N_4992);
nor UO_98 (O_98,N_4916,N_4975);
or UO_99 (O_99,N_4941,N_4930);
nor UO_100 (O_100,N_4954,N_4968);
or UO_101 (O_101,N_4942,N_4990);
nand UO_102 (O_102,N_4974,N_4948);
or UO_103 (O_103,N_4936,N_4917);
or UO_104 (O_104,N_4984,N_4934);
xnor UO_105 (O_105,N_4912,N_4971);
nand UO_106 (O_106,N_4952,N_4926);
and UO_107 (O_107,N_4916,N_4900);
nand UO_108 (O_108,N_4951,N_4967);
nor UO_109 (O_109,N_4948,N_4952);
nand UO_110 (O_110,N_4957,N_4901);
and UO_111 (O_111,N_4963,N_4907);
nor UO_112 (O_112,N_4916,N_4950);
xor UO_113 (O_113,N_4906,N_4914);
xor UO_114 (O_114,N_4980,N_4928);
or UO_115 (O_115,N_4975,N_4964);
xnor UO_116 (O_116,N_4963,N_4989);
xor UO_117 (O_117,N_4903,N_4902);
and UO_118 (O_118,N_4981,N_4973);
and UO_119 (O_119,N_4945,N_4939);
xnor UO_120 (O_120,N_4978,N_4951);
or UO_121 (O_121,N_4957,N_4979);
nand UO_122 (O_122,N_4917,N_4962);
and UO_123 (O_123,N_4970,N_4916);
and UO_124 (O_124,N_4919,N_4998);
nor UO_125 (O_125,N_4976,N_4902);
or UO_126 (O_126,N_4989,N_4943);
or UO_127 (O_127,N_4935,N_4945);
nand UO_128 (O_128,N_4929,N_4915);
nor UO_129 (O_129,N_4941,N_4904);
nand UO_130 (O_130,N_4912,N_4906);
nand UO_131 (O_131,N_4973,N_4975);
or UO_132 (O_132,N_4955,N_4922);
xnor UO_133 (O_133,N_4954,N_4993);
and UO_134 (O_134,N_4973,N_4919);
or UO_135 (O_135,N_4919,N_4991);
and UO_136 (O_136,N_4936,N_4964);
nor UO_137 (O_137,N_4938,N_4951);
and UO_138 (O_138,N_4992,N_4975);
xnor UO_139 (O_139,N_4901,N_4916);
and UO_140 (O_140,N_4943,N_4912);
or UO_141 (O_141,N_4908,N_4925);
nor UO_142 (O_142,N_4971,N_4947);
xor UO_143 (O_143,N_4970,N_4985);
or UO_144 (O_144,N_4968,N_4937);
and UO_145 (O_145,N_4973,N_4989);
nor UO_146 (O_146,N_4904,N_4985);
and UO_147 (O_147,N_4974,N_4978);
nand UO_148 (O_148,N_4908,N_4956);
nand UO_149 (O_149,N_4959,N_4922);
nand UO_150 (O_150,N_4949,N_4912);
nand UO_151 (O_151,N_4919,N_4988);
and UO_152 (O_152,N_4963,N_4962);
or UO_153 (O_153,N_4936,N_4983);
nor UO_154 (O_154,N_4960,N_4996);
xor UO_155 (O_155,N_4903,N_4923);
and UO_156 (O_156,N_4984,N_4906);
or UO_157 (O_157,N_4986,N_4976);
and UO_158 (O_158,N_4904,N_4926);
xnor UO_159 (O_159,N_4967,N_4954);
and UO_160 (O_160,N_4950,N_4960);
and UO_161 (O_161,N_4903,N_4998);
nor UO_162 (O_162,N_4996,N_4955);
nand UO_163 (O_163,N_4962,N_4976);
and UO_164 (O_164,N_4901,N_4986);
nor UO_165 (O_165,N_4974,N_4920);
or UO_166 (O_166,N_4950,N_4943);
or UO_167 (O_167,N_4913,N_4975);
and UO_168 (O_168,N_4975,N_4939);
and UO_169 (O_169,N_4934,N_4964);
and UO_170 (O_170,N_4936,N_4935);
or UO_171 (O_171,N_4947,N_4929);
nor UO_172 (O_172,N_4942,N_4939);
nor UO_173 (O_173,N_4990,N_4914);
nor UO_174 (O_174,N_4906,N_4965);
xor UO_175 (O_175,N_4923,N_4983);
nor UO_176 (O_176,N_4989,N_4933);
and UO_177 (O_177,N_4950,N_4913);
and UO_178 (O_178,N_4951,N_4958);
and UO_179 (O_179,N_4911,N_4959);
and UO_180 (O_180,N_4923,N_4998);
nand UO_181 (O_181,N_4989,N_4979);
and UO_182 (O_182,N_4941,N_4902);
nand UO_183 (O_183,N_4941,N_4994);
nand UO_184 (O_184,N_4977,N_4969);
or UO_185 (O_185,N_4939,N_4908);
xnor UO_186 (O_186,N_4969,N_4911);
and UO_187 (O_187,N_4921,N_4929);
nor UO_188 (O_188,N_4909,N_4989);
or UO_189 (O_189,N_4938,N_4918);
nor UO_190 (O_190,N_4967,N_4965);
or UO_191 (O_191,N_4985,N_4941);
nand UO_192 (O_192,N_4986,N_4958);
and UO_193 (O_193,N_4998,N_4970);
or UO_194 (O_194,N_4971,N_4917);
and UO_195 (O_195,N_4990,N_4984);
and UO_196 (O_196,N_4932,N_4942);
nor UO_197 (O_197,N_4902,N_4942);
nand UO_198 (O_198,N_4952,N_4966);
nand UO_199 (O_199,N_4922,N_4954);
nor UO_200 (O_200,N_4959,N_4981);
and UO_201 (O_201,N_4989,N_4907);
nor UO_202 (O_202,N_4912,N_4966);
or UO_203 (O_203,N_4966,N_4996);
xor UO_204 (O_204,N_4904,N_4901);
and UO_205 (O_205,N_4928,N_4968);
nand UO_206 (O_206,N_4983,N_4957);
and UO_207 (O_207,N_4918,N_4947);
and UO_208 (O_208,N_4916,N_4994);
and UO_209 (O_209,N_4960,N_4918);
or UO_210 (O_210,N_4977,N_4921);
and UO_211 (O_211,N_4909,N_4987);
or UO_212 (O_212,N_4967,N_4914);
or UO_213 (O_213,N_4990,N_4945);
xnor UO_214 (O_214,N_4978,N_4928);
and UO_215 (O_215,N_4944,N_4958);
or UO_216 (O_216,N_4955,N_4917);
xor UO_217 (O_217,N_4997,N_4991);
nand UO_218 (O_218,N_4999,N_4940);
or UO_219 (O_219,N_4922,N_4918);
nand UO_220 (O_220,N_4928,N_4987);
nand UO_221 (O_221,N_4973,N_4900);
or UO_222 (O_222,N_4957,N_4906);
nand UO_223 (O_223,N_4982,N_4986);
or UO_224 (O_224,N_4983,N_4907);
nor UO_225 (O_225,N_4926,N_4937);
nor UO_226 (O_226,N_4991,N_4923);
nor UO_227 (O_227,N_4936,N_4906);
nand UO_228 (O_228,N_4927,N_4942);
and UO_229 (O_229,N_4966,N_4997);
nand UO_230 (O_230,N_4921,N_4942);
nor UO_231 (O_231,N_4932,N_4905);
or UO_232 (O_232,N_4908,N_4905);
nor UO_233 (O_233,N_4961,N_4919);
or UO_234 (O_234,N_4903,N_4911);
and UO_235 (O_235,N_4992,N_4933);
and UO_236 (O_236,N_4985,N_4947);
nor UO_237 (O_237,N_4904,N_4998);
or UO_238 (O_238,N_4912,N_4947);
or UO_239 (O_239,N_4988,N_4966);
or UO_240 (O_240,N_4995,N_4987);
or UO_241 (O_241,N_4934,N_4927);
or UO_242 (O_242,N_4935,N_4968);
nand UO_243 (O_243,N_4956,N_4951);
and UO_244 (O_244,N_4956,N_4965);
and UO_245 (O_245,N_4930,N_4965);
nor UO_246 (O_246,N_4993,N_4974);
nand UO_247 (O_247,N_4935,N_4912);
or UO_248 (O_248,N_4938,N_4936);
or UO_249 (O_249,N_4951,N_4982);
xor UO_250 (O_250,N_4992,N_4934);
and UO_251 (O_251,N_4974,N_4995);
nor UO_252 (O_252,N_4903,N_4958);
nor UO_253 (O_253,N_4981,N_4952);
or UO_254 (O_254,N_4914,N_4988);
nor UO_255 (O_255,N_4921,N_4987);
nand UO_256 (O_256,N_4908,N_4915);
or UO_257 (O_257,N_4929,N_4954);
nand UO_258 (O_258,N_4984,N_4901);
or UO_259 (O_259,N_4908,N_4957);
and UO_260 (O_260,N_4947,N_4943);
xor UO_261 (O_261,N_4929,N_4973);
nor UO_262 (O_262,N_4950,N_4995);
or UO_263 (O_263,N_4914,N_4994);
and UO_264 (O_264,N_4984,N_4980);
or UO_265 (O_265,N_4986,N_4914);
xor UO_266 (O_266,N_4974,N_4902);
xor UO_267 (O_267,N_4971,N_4909);
nand UO_268 (O_268,N_4930,N_4995);
nand UO_269 (O_269,N_4994,N_4915);
or UO_270 (O_270,N_4942,N_4952);
nand UO_271 (O_271,N_4987,N_4994);
or UO_272 (O_272,N_4918,N_4908);
and UO_273 (O_273,N_4931,N_4994);
nor UO_274 (O_274,N_4986,N_4937);
xor UO_275 (O_275,N_4954,N_4992);
or UO_276 (O_276,N_4976,N_4965);
and UO_277 (O_277,N_4926,N_4923);
or UO_278 (O_278,N_4928,N_4921);
nand UO_279 (O_279,N_4976,N_4939);
nand UO_280 (O_280,N_4918,N_4992);
or UO_281 (O_281,N_4917,N_4937);
xnor UO_282 (O_282,N_4915,N_4909);
and UO_283 (O_283,N_4934,N_4937);
nor UO_284 (O_284,N_4958,N_4959);
nand UO_285 (O_285,N_4921,N_4988);
nor UO_286 (O_286,N_4972,N_4988);
nand UO_287 (O_287,N_4980,N_4934);
nand UO_288 (O_288,N_4928,N_4935);
xnor UO_289 (O_289,N_4904,N_4966);
xnor UO_290 (O_290,N_4928,N_4981);
nand UO_291 (O_291,N_4928,N_4997);
nand UO_292 (O_292,N_4939,N_4993);
nor UO_293 (O_293,N_4907,N_4928);
and UO_294 (O_294,N_4974,N_4966);
nor UO_295 (O_295,N_4997,N_4930);
and UO_296 (O_296,N_4964,N_4989);
or UO_297 (O_297,N_4978,N_4940);
and UO_298 (O_298,N_4911,N_4990);
or UO_299 (O_299,N_4933,N_4958);
nor UO_300 (O_300,N_4967,N_4922);
nand UO_301 (O_301,N_4934,N_4989);
nand UO_302 (O_302,N_4914,N_4971);
nand UO_303 (O_303,N_4950,N_4981);
or UO_304 (O_304,N_4921,N_4930);
nand UO_305 (O_305,N_4990,N_4947);
nand UO_306 (O_306,N_4909,N_4911);
nand UO_307 (O_307,N_4963,N_4936);
or UO_308 (O_308,N_4990,N_4960);
or UO_309 (O_309,N_4989,N_4996);
or UO_310 (O_310,N_4905,N_4959);
nor UO_311 (O_311,N_4904,N_4989);
nor UO_312 (O_312,N_4907,N_4974);
and UO_313 (O_313,N_4974,N_4916);
nor UO_314 (O_314,N_4996,N_4990);
nand UO_315 (O_315,N_4908,N_4990);
nor UO_316 (O_316,N_4911,N_4998);
and UO_317 (O_317,N_4950,N_4979);
nand UO_318 (O_318,N_4906,N_4976);
and UO_319 (O_319,N_4909,N_4976);
and UO_320 (O_320,N_4916,N_4904);
or UO_321 (O_321,N_4982,N_4936);
nand UO_322 (O_322,N_4966,N_4941);
or UO_323 (O_323,N_4945,N_4934);
or UO_324 (O_324,N_4949,N_4929);
nor UO_325 (O_325,N_4963,N_4973);
nand UO_326 (O_326,N_4913,N_4938);
xnor UO_327 (O_327,N_4949,N_4943);
or UO_328 (O_328,N_4960,N_4985);
nand UO_329 (O_329,N_4942,N_4994);
nor UO_330 (O_330,N_4967,N_4923);
and UO_331 (O_331,N_4927,N_4994);
and UO_332 (O_332,N_4969,N_4935);
or UO_333 (O_333,N_4938,N_4967);
nand UO_334 (O_334,N_4960,N_4972);
nand UO_335 (O_335,N_4907,N_4905);
nand UO_336 (O_336,N_4900,N_4915);
nand UO_337 (O_337,N_4992,N_4997);
or UO_338 (O_338,N_4977,N_4915);
and UO_339 (O_339,N_4928,N_4973);
or UO_340 (O_340,N_4943,N_4972);
nor UO_341 (O_341,N_4993,N_4990);
nand UO_342 (O_342,N_4999,N_4977);
or UO_343 (O_343,N_4957,N_4932);
and UO_344 (O_344,N_4985,N_4912);
and UO_345 (O_345,N_4921,N_4941);
nor UO_346 (O_346,N_4916,N_4942);
nor UO_347 (O_347,N_4974,N_4931);
and UO_348 (O_348,N_4915,N_4903);
or UO_349 (O_349,N_4964,N_4900);
nor UO_350 (O_350,N_4977,N_4962);
and UO_351 (O_351,N_4949,N_4919);
and UO_352 (O_352,N_4913,N_4931);
or UO_353 (O_353,N_4936,N_4916);
nor UO_354 (O_354,N_4956,N_4959);
and UO_355 (O_355,N_4941,N_4935);
or UO_356 (O_356,N_4961,N_4945);
or UO_357 (O_357,N_4974,N_4971);
or UO_358 (O_358,N_4945,N_4968);
or UO_359 (O_359,N_4959,N_4945);
nor UO_360 (O_360,N_4936,N_4979);
nand UO_361 (O_361,N_4938,N_4968);
xor UO_362 (O_362,N_4934,N_4972);
or UO_363 (O_363,N_4970,N_4903);
xnor UO_364 (O_364,N_4960,N_4906);
and UO_365 (O_365,N_4911,N_4985);
xor UO_366 (O_366,N_4943,N_4954);
and UO_367 (O_367,N_4945,N_4933);
nor UO_368 (O_368,N_4961,N_4911);
nor UO_369 (O_369,N_4914,N_4998);
and UO_370 (O_370,N_4933,N_4995);
and UO_371 (O_371,N_4931,N_4944);
and UO_372 (O_372,N_4942,N_4972);
nor UO_373 (O_373,N_4993,N_4912);
nand UO_374 (O_374,N_4982,N_4957);
and UO_375 (O_375,N_4932,N_4951);
nor UO_376 (O_376,N_4976,N_4966);
nor UO_377 (O_377,N_4917,N_4990);
and UO_378 (O_378,N_4937,N_4948);
or UO_379 (O_379,N_4922,N_4983);
or UO_380 (O_380,N_4936,N_4973);
or UO_381 (O_381,N_4997,N_4927);
nor UO_382 (O_382,N_4951,N_4900);
and UO_383 (O_383,N_4937,N_4911);
nand UO_384 (O_384,N_4907,N_4916);
and UO_385 (O_385,N_4995,N_4966);
or UO_386 (O_386,N_4985,N_4962);
nor UO_387 (O_387,N_4938,N_4996);
nand UO_388 (O_388,N_4900,N_4940);
and UO_389 (O_389,N_4987,N_4923);
nor UO_390 (O_390,N_4994,N_4982);
and UO_391 (O_391,N_4977,N_4994);
and UO_392 (O_392,N_4984,N_4933);
xnor UO_393 (O_393,N_4934,N_4998);
nor UO_394 (O_394,N_4950,N_4948);
nand UO_395 (O_395,N_4930,N_4961);
xnor UO_396 (O_396,N_4941,N_4999);
nand UO_397 (O_397,N_4948,N_4914);
or UO_398 (O_398,N_4900,N_4911);
and UO_399 (O_399,N_4922,N_4958);
or UO_400 (O_400,N_4953,N_4941);
nand UO_401 (O_401,N_4921,N_4918);
nand UO_402 (O_402,N_4929,N_4924);
nor UO_403 (O_403,N_4930,N_4972);
and UO_404 (O_404,N_4941,N_4940);
and UO_405 (O_405,N_4976,N_4998);
nor UO_406 (O_406,N_4944,N_4903);
nor UO_407 (O_407,N_4982,N_4917);
and UO_408 (O_408,N_4976,N_4987);
xor UO_409 (O_409,N_4957,N_4911);
nor UO_410 (O_410,N_4996,N_4909);
nor UO_411 (O_411,N_4999,N_4922);
or UO_412 (O_412,N_4940,N_4944);
or UO_413 (O_413,N_4958,N_4936);
and UO_414 (O_414,N_4901,N_4994);
or UO_415 (O_415,N_4997,N_4963);
nand UO_416 (O_416,N_4984,N_4902);
or UO_417 (O_417,N_4959,N_4998);
and UO_418 (O_418,N_4993,N_4979);
nand UO_419 (O_419,N_4905,N_4924);
nand UO_420 (O_420,N_4980,N_4915);
and UO_421 (O_421,N_4926,N_4939);
or UO_422 (O_422,N_4928,N_4929);
and UO_423 (O_423,N_4931,N_4962);
and UO_424 (O_424,N_4942,N_4973);
nor UO_425 (O_425,N_4962,N_4987);
or UO_426 (O_426,N_4967,N_4947);
or UO_427 (O_427,N_4975,N_4927);
xor UO_428 (O_428,N_4981,N_4940);
and UO_429 (O_429,N_4981,N_4958);
or UO_430 (O_430,N_4997,N_4908);
and UO_431 (O_431,N_4968,N_4915);
or UO_432 (O_432,N_4962,N_4979);
nand UO_433 (O_433,N_4990,N_4931);
nor UO_434 (O_434,N_4913,N_4939);
nor UO_435 (O_435,N_4964,N_4985);
and UO_436 (O_436,N_4917,N_4993);
nand UO_437 (O_437,N_4976,N_4919);
nor UO_438 (O_438,N_4979,N_4976);
nor UO_439 (O_439,N_4946,N_4954);
nor UO_440 (O_440,N_4922,N_4985);
or UO_441 (O_441,N_4942,N_4903);
and UO_442 (O_442,N_4988,N_4977);
nor UO_443 (O_443,N_4930,N_4977);
nor UO_444 (O_444,N_4995,N_4988);
and UO_445 (O_445,N_4902,N_4986);
nor UO_446 (O_446,N_4932,N_4990);
and UO_447 (O_447,N_4903,N_4945);
and UO_448 (O_448,N_4904,N_4919);
xnor UO_449 (O_449,N_4905,N_4915);
xor UO_450 (O_450,N_4989,N_4936);
and UO_451 (O_451,N_4919,N_4944);
and UO_452 (O_452,N_4971,N_4932);
and UO_453 (O_453,N_4975,N_4970);
and UO_454 (O_454,N_4932,N_4931);
or UO_455 (O_455,N_4939,N_4924);
nand UO_456 (O_456,N_4983,N_4987);
or UO_457 (O_457,N_4964,N_4946);
xnor UO_458 (O_458,N_4952,N_4956);
or UO_459 (O_459,N_4929,N_4943);
or UO_460 (O_460,N_4973,N_4913);
nand UO_461 (O_461,N_4985,N_4984);
nor UO_462 (O_462,N_4906,N_4945);
nand UO_463 (O_463,N_4948,N_4963);
and UO_464 (O_464,N_4986,N_4940);
nor UO_465 (O_465,N_4925,N_4923);
or UO_466 (O_466,N_4905,N_4918);
and UO_467 (O_467,N_4925,N_4946);
or UO_468 (O_468,N_4959,N_4963);
or UO_469 (O_469,N_4972,N_4959);
nand UO_470 (O_470,N_4998,N_4957);
nand UO_471 (O_471,N_4958,N_4948);
nand UO_472 (O_472,N_4903,N_4973);
nor UO_473 (O_473,N_4904,N_4911);
and UO_474 (O_474,N_4959,N_4912);
nor UO_475 (O_475,N_4953,N_4933);
nand UO_476 (O_476,N_4906,N_4953);
or UO_477 (O_477,N_4968,N_4969);
nor UO_478 (O_478,N_4918,N_4920);
or UO_479 (O_479,N_4956,N_4939);
nor UO_480 (O_480,N_4963,N_4901);
nor UO_481 (O_481,N_4957,N_4945);
xnor UO_482 (O_482,N_4937,N_4965);
xor UO_483 (O_483,N_4919,N_4942);
nand UO_484 (O_484,N_4914,N_4927);
nand UO_485 (O_485,N_4931,N_4915);
nor UO_486 (O_486,N_4914,N_4976);
or UO_487 (O_487,N_4923,N_4906);
and UO_488 (O_488,N_4929,N_4944);
or UO_489 (O_489,N_4995,N_4937);
nand UO_490 (O_490,N_4996,N_4978);
or UO_491 (O_491,N_4926,N_4914);
nor UO_492 (O_492,N_4951,N_4994);
nand UO_493 (O_493,N_4931,N_4912);
or UO_494 (O_494,N_4963,N_4968);
or UO_495 (O_495,N_4975,N_4918);
nand UO_496 (O_496,N_4959,N_4914);
xor UO_497 (O_497,N_4960,N_4962);
nand UO_498 (O_498,N_4957,N_4967);
nand UO_499 (O_499,N_4922,N_4900);
or UO_500 (O_500,N_4997,N_4918);
nor UO_501 (O_501,N_4967,N_4997);
or UO_502 (O_502,N_4972,N_4976);
or UO_503 (O_503,N_4935,N_4992);
xor UO_504 (O_504,N_4940,N_4903);
and UO_505 (O_505,N_4930,N_4942);
or UO_506 (O_506,N_4907,N_4996);
and UO_507 (O_507,N_4988,N_4997);
nor UO_508 (O_508,N_4977,N_4957);
or UO_509 (O_509,N_4989,N_4926);
nand UO_510 (O_510,N_4906,N_4961);
nand UO_511 (O_511,N_4917,N_4965);
and UO_512 (O_512,N_4986,N_4993);
nand UO_513 (O_513,N_4953,N_4919);
xor UO_514 (O_514,N_4948,N_4939);
nand UO_515 (O_515,N_4989,N_4995);
nor UO_516 (O_516,N_4940,N_4975);
or UO_517 (O_517,N_4910,N_4987);
and UO_518 (O_518,N_4998,N_4955);
or UO_519 (O_519,N_4916,N_4918);
nor UO_520 (O_520,N_4981,N_4936);
nand UO_521 (O_521,N_4999,N_4974);
nand UO_522 (O_522,N_4943,N_4960);
or UO_523 (O_523,N_4987,N_4949);
and UO_524 (O_524,N_4982,N_4946);
nand UO_525 (O_525,N_4999,N_4991);
xor UO_526 (O_526,N_4950,N_4974);
xor UO_527 (O_527,N_4999,N_4978);
or UO_528 (O_528,N_4958,N_4987);
nor UO_529 (O_529,N_4952,N_4902);
and UO_530 (O_530,N_4967,N_4916);
nor UO_531 (O_531,N_4964,N_4931);
xnor UO_532 (O_532,N_4965,N_4905);
or UO_533 (O_533,N_4906,N_4986);
or UO_534 (O_534,N_4987,N_4999);
and UO_535 (O_535,N_4971,N_4988);
nand UO_536 (O_536,N_4923,N_4956);
and UO_537 (O_537,N_4925,N_4972);
and UO_538 (O_538,N_4923,N_4922);
nand UO_539 (O_539,N_4902,N_4916);
and UO_540 (O_540,N_4911,N_4930);
nor UO_541 (O_541,N_4965,N_4923);
nand UO_542 (O_542,N_4902,N_4964);
or UO_543 (O_543,N_4940,N_4931);
or UO_544 (O_544,N_4925,N_4930);
nand UO_545 (O_545,N_4958,N_4908);
and UO_546 (O_546,N_4998,N_4926);
nand UO_547 (O_547,N_4914,N_4983);
nor UO_548 (O_548,N_4992,N_4906);
and UO_549 (O_549,N_4922,N_4989);
or UO_550 (O_550,N_4956,N_4941);
nand UO_551 (O_551,N_4962,N_4940);
and UO_552 (O_552,N_4943,N_4990);
nand UO_553 (O_553,N_4991,N_4986);
nor UO_554 (O_554,N_4924,N_4933);
and UO_555 (O_555,N_4918,N_4926);
or UO_556 (O_556,N_4983,N_4986);
and UO_557 (O_557,N_4959,N_4971);
nand UO_558 (O_558,N_4993,N_4910);
and UO_559 (O_559,N_4990,N_4937);
and UO_560 (O_560,N_4917,N_4928);
and UO_561 (O_561,N_4967,N_4976);
and UO_562 (O_562,N_4991,N_4980);
or UO_563 (O_563,N_4936,N_4925);
and UO_564 (O_564,N_4955,N_4940);
or UO_565 (O_565,N_4950,N_4954);
and UO_566 (O_566,N_4922,N_4971);
nor UO_567 (O_567,N_4903,N_4938);
nor UO_568 (O_568,N_4948,N_4907);
or UO_569 (O_569,N_4906,N_4938);
nand UO_570 (O_570,N_4939,N_4911);
and UO_571 (O_571,N_4922,N_4907);
and UO_572 (O_572,N_4956,N_4979);
and UO_573 (O_573,N_4954,N_4910);
or UO_574 (O_574,N_4996,N_4952);
nor UO_575 (O_575,N_4989,N_4990);
nand UO_576 (O_576,N_4957,N_4971);
and UO_577 (O_577,N_4997,N_4948);
or UO_578 (O_578,N_4980,N_4914);
nor UO_579 (O_579,N_4904,N_4928);
and UO_580 (O_580,N_4911,N_4908);
and UO_581 (O_581,N_4974,N_4987);
and UO_582 (O_582,N_4903,N_4982);
xor UO_583 (O_583,N_4939,N_4963);
and UO_584 (O_584,N_4924,N_4906);
nand UO_585 (O_585,N_4958,N_4974);
nor UO_586 (O_586,N_4917,N_4942);
nor UO_587 (O_587,N_4969,N_4958);
nor UO_588 (O_588,N_4921,N_4965);
nor UO_589 (O_589,N_4933,N_4964);
nor UO_590 (O_590,N_4943,N_4907);
and UO_591 (O_591,N_4947,N_4922);
or UO_592 (O_592,N_4960,N_4913);
nand UO_593 (O_593,N_4951,N_4981);
or UO_594 (O_594,N_4986,N_4951);
and UO_595 (O_595,N_4923,N_4970);
nor UO_596 (O_596,N_4981,N_4984);
and UO_597 (O_597,N_4967,N_4955);
or UO_598 (O_598,N_4974,N_4928);
and UO_599 (O_599,N_4991,N_4998);
and UO_600 (O_600,N_4922,N_4977);
or UO_601 (O_601,N_4991,N_4954);
xor UO_602 (O_602,N_4901,N_4924);
or UO_603 (O_603,N_4993,N_4934);
xor UO_604 (O_604,N_4977,N_4964);
nor UO_605 (O_605,N_4975,N_4999);
nor UO_606 (O_606,N_4961,N_4931);
nor UO_607 (O_607,N_4913,N_4991);
nand UO_608 (O_608,N_4961,N_4941);
nand UO_609 (O_609,N_4963,N_4994);
nand UO_610 (O_610,N_4955,N_4918);
and UO_611 (O_611,N_4937,N_4914);
nor UO_612 (O_612,N_4926,N_4971);
nand UO_613 (O_613,N_4953,N_4996);
nand UO_614 (O_614,N_4998,N_4938);
nand UO_615 (O_615,N_4910,N_4963);
nor UO_616 (O_616,N_4927,N_4989);
or UO_617 (O_617,N_4909,N_4995);
nor UO_618 (O_618,N_4918,N_4983);
nand UO_619 (O_619,N_4985,N_4979);
and UO_620 (O_620,N_4960,N_4975);
and UO_621 (O_621,N_4952,N_4963);
nand UO_622 (O_622,N_4913,N_4965);
nand UO_623 (O_623,N_4990,N_4915);
nor UO_624 (O_624,N_4994,N_4910);
xor UO_625 (O_625,N_4981,N_4978);
nand UO_626 (O_626,N_4907,N_4933);
or UO_627 (O_627,N_4928,N_4994);
nand UO_628 (O_628,N_4944,N_4977);
nor UO_629 (O_629,N_4957,N_4975);
nand UO_630 (O_630,N_4966,N_4970);
nor UO_631 (O_631,N_4994,N_4902);
or UO_632 (O_632,N_4969,N_4956);
nor UO_633 (O_633,N_4968,N_4993);
nand UO_634 (O_634,N_4977,N_4991);
nand UO_635 (O_635,N_4971,N_4983);
or UO_636 (O_636,N_4924,N_4989);
nand UO_637 (O_637,N_4995,N_4913);
nand UO_638 (O_638,N_4916,N_4998);
or UO_639 (O_639,N_4929,N_4959);
nor UO_640 (O_640,N_4953,N_4938);
and UO_641 (O_641,N_4959,N_4976);
nand UO_642 (O_642,N_4905,N_4964);
and UO_643 (O_643,N_4947,N_4962);
xor UO_644 (O_644,N_4951,N_4995);
and UO_645 (O_645,N_4914,N_4951);
nand UO_646 (O_646,N_4993,N_4955);
nor UO_647 (O_647,N_4970,N_4921);
xor UO_648 (O_648,N_4989,N_4998);
nor UO_649 (O_649,N_4919,N_4986);
or UO_650 (O_650,N_4923,N_4911);
nand UO_651 (O_651,N_4950,N_4908);
nand UO_652 (O_652,N_4906,N_4952);
or UO_653 (O_653,N_4990,N_4974);
nor UO_654 (O_654,N_4946,N_4943);
nor UO_655 (O_655,N_4913,N_4924);
nor UO_656 (O_656,N_4967,N_4906);
and UO_657 (O_657,N_4920,N_4985);
nor UO_658 (O_658,N_4996,N_4943);
or UO_659 (O_659,N_4932,N_4919);
and UO_660 (O_660,N_4925,N_4995);
or UO_661 (O_661,N_4978,N_4905);
nor UO_662 (O_662,N_4953,N_4989);
or UO_663 (O_663,N_4982,N_4914);
nor UO_664 (O_664,N_4994,N_4939);
nor UO_665 (O_665,N_4970,N_4941);
nor UO_666 (O_666,N_4918,N_4977);
or UO_667 (O_667,N_4937,N_4902);
nor UO_668 (O_668,N_4949,N_4906);
nor UO_669 (O_669,N_4978,N_4969);
nor UO_670 (O_670,N_4913,N_4908);
and UO_671 (O_671,N_4917,N_4979);
or UO_672 (O_672,N_4965,N_4934);
nand UO_673 (O_673,N_4971,N_4943);
and UO_674 (O_674,N_4969,N_4947);
and UO_675 (O_675,N_4998,N_4950);
nor UO_676 (O_676,N_4912,N_4905);
or UO_677 (O_677,N_4961,N_4982);
nand UO_678 (O_678,N_4983,N_4900);
nor UO_679 (O_679,N_4973,N_4904);
nor UO_680 (O_680,N_4975,N_4994);
xnor UO_681 (O_681,N_4928,N_4924);
nand UO_682 (O_682,N_4947,N_4921);
nor UO_683 (O_683,N_4962,N_4984);
or UO_684 (O_684,N_4945,N_4904);
or UO_685 (O_685,N_4963,N_4934);
or UO_686 (O_686,N_4903,N_4965);
nor UO_687 (O_687,N_4974,N_4922);
nor UO_688 (O_688,N_4918,N_4936);
nor UO_689 (O_689,N_4920,N_4966);
xnor UO_690 (O_690,N_4987,N_4902);
and UO_691 (O_691,N_4945,N_4981);
nor UO_692 (O_692,N_4994,N_4961);
nand UO_693 (O_693,N_4992,N_4925);
and UO_694 (O_694,N_4906,N_4995);
nor UO_695 (O_695,N_4985,N_4943);
nor UO_696 (O_696,N_4938,N_4900);
nor UO_697 (O_697,N_4919,N_4970);
or UO_698 (O_698,N_4945,N_4993);
xnor UO_699 (O_699,N_4994,N_4948);
or UO_700 (O_700,N_4939,N_4967);
nor UO_701 (O_701,N_4968,N_4977);
nand UO_702 (O_702,N_4930,N_4956);
or UO_703 (O_703,N_4920,N_4927);
nand UO_704 (O_704,N_4923,N_4975);
and UO_705 (O_705,N_4959,N_4939);
or UO_706 (O_706,N_4912,N_4979);
and UO_707 (O_707,N_4995,N_4946);
nand UO_708 (O_708,N_4934,N_4976);
nor UO_709 (O_709,N_4905,N_4921);
and UO_710 (O_710,N_4931,N_4986);
or UO_711 (O_711,N_4978,N_4979);
nand UO_712 (O_712,N_4950,N_4985);
or UO_713 (O_713,N_4937,N_4983);
or UO_714 (O_714,N_4961,N_4976);
or UO_715 (O_715,N_4955,N_4946);
nor UO_716 (O_716,N_4969,N_4999);
or UO_717 (O_717,N_4991,N_4947);
xnor UO_718 (O_718,N_4909,N_4999);
nor UO_719 (O_719,N_4964,N_4909);
nand UO_720 (O_720,N_4946,N_4941);
and UO_721 (O_721,N_4908,N_4953);
nor UO_722 (O_722,N_4947,N_4904);
nand UO_723 (O_723,N_4910,N_4926);
and UO_724 (O_724,N_4961,N_4960);
nand UO_725 (O_725,N_4915,N_4992);
nand UO_726 (O_726,N_4943,N_4940);
and UO_727 (O_727,N_4901,N_4917);
nand UO_728 (O_728,N_4943,N_4993);
xnor UO_729 (O_729,N_4902,N_4981);
or UO_730 (O_730,N_4962,N_4969);
and UO_731 (O_731,N_4968,N_4970);
nor UO_732 (O_732,N_4948,N_4971);
and UO_733 (O_733,N_4998,N_4947);
nand UO_734 (O_734,N_4907,N_4975);
or UO_735 (O_735,N_4986,N_4930);
or UO_736 (O_736,N_4948,N_4925);
and UO_737 (O_737,N_4957,N_4935);
and UO_738 (O_738,N_4900,N_4988);
xnor UO_739 (O_739,N_4958,N_4980);
xnor UO_740 (O_740,N_4936,N_4988);
xnor UO_741 (O_741,N_4914,N_4900);
or UO_742 (O_742,N_4933,N_4926);
or UO_743 (O_743,N_4976,N_4925);
and UO_744 (O_744,N_4920,N_4946);
and UO_745 (O_745,N_4900,N_4936);
and UO_746 (O_746,N_4995,N_4963);
nor UO_747 (O_747,N_4940,N_4911);
nand UO_748 (O_748,N_4919,N_4992);
and UO_749 (O_749,N_4928,N_4941);
nor UO_750 (O_750,N_4984,N_4905);
xor UO_751 (O_751,N_4996,N_4944);
nor UO_752 (O_752,N_4920,N_4948);
or UO_753 (O_753,N_4963,N_4982);
nor UO_754 (O_754,N_4965,N_4914);
xor UO_755 (O_755,N_4968,N_4950);
nand UO_756 (O_756,N_4910,N_4952);
nor UO_757 (O_757,N_4947,N_4942);
nand UO_758 (O_758,N_4998,N_4948);
or UO_759 (O_759,N_4935,N_4963);
nand UO_760 (O_760,N_4905,N_4963);
nor UO_761 (O_761,N_4969,N_4953);
and UO_762 (O_762,N_4938,N_4919);
and UO_763 (O_763,N_4912,N_4978);
and UO_764 (O_764,N_4938,N_4969);
and UO_765 (O_765,N_4960,N_4916);
nand UO_766 (O_766,N_4920,N_4954);
nand UO_767 (O_767,N_4903,N_4941);
nor UO_768 (O_768,N_4985,N_4939);
xnor UO_769 (O_769,N_4932,N_4916);
xnor UO_770 (O_770,N_4948,N_4970);
nor UO_771 (O_771,N_4992,N_4911);
or UO_772 (O_772,N_4922,N_4987);
or UO_773 (O_773,N_4957,N_4909);
xnor UO_774 (O_774,N_4991,N_4989);
nor UO_775 (O_775,N_4926,N_4913);
and UO_776 (O_776,N_4978,N_4958);
or UO_777 (O_777,N_4996,N_4900);
and UO_778 (O_778,N_4952,N_4989);
and UO_779 (O_779,N_4994,N_4944);
or UO_780 (O_780,N_4919,N_4975);
and UO_781 (O_781,N_4918,N_4911);
and UO_782 (O_782,N_4938,N_4924);
or UO_783 (O_783,N_4932,N_4981);
and UO_784 (O_784,N_4990,N_4906);
or UO_785 (O_785,N_4959,N_4970);
or UO_786 (O_786,N_4930,N_4968);
xor UO_787 (O_787,N_4962,N_4968);
and UO_788 (O_788,N_4922,N_4913);
and UO_789 (O_789,N_4977,N_4901);
and UO_790 (O_790,N_4973,N_4977);
nand UO_791 (O_791,N_4903,N_4933);
xnor UO_792 (O_792,N_4974,N_4972);
nor UO_793 (O_793,N_4959,N_4950);
nand UO_794 (O_794,N_4971,N_4944);
xor UO_795 (O_795,N_4911,N_4984);
or UO_796 (O_796,N_4959,N_4982);
or UO_797 (O_797,N_4963,N_4971);
xor UO_798 (O_798,N_4908,N_4980);
nor UO_799 (O_799,N_4990,N_4964);
and UO_800 (O_800,N_4945,N_4992);
and UO_801 (O_801,N_4936,N_4919);
and UO_802 (O_802,N_4953,N_4902);
and UO_803 (O_803,N_4962,N_4900);
nor UO_804 (O_804,N_4910,N_4965);
nand UO_805 (O_805,N_4923,N_4907);
nand UO_806 (O_806,N_4922,N_4906);
and UO_807 (O_807,N_4959,N_4903);
nand UO_808 (O_808,N_4925,N_4970);
or UO_809 (O_809,N_4969,N_4992);
or UO_810 (O_810,N_4963,N_4938);
nand UO_811 (O_811,N_4905,N_4961);
nor UO_812 (O_812,N_4920,N_4964);
or UO_813 (O_813,N_4942,N_4922);
and UO_814 (O_814,N_4983,N_4995);
xor UO_815 (O_815,N_4947,N_4978);
and UO_816 (O_816,N_4908,N_4985);
and UO_817 (O_817,N_4902,N_4963);
xnor UO_818 (O_818,N_4949,N_4930);
xor UO_819 (O_819,N_4973,N_4927);
nand UO_820 (O_820,N_4903,N_4934);
nor UO_821 (O_821,N_4987,N_4956);
and UO_822 (O_822,N_4917,N_4927);
nor UO_823 (O_823,N_4924,N_4920);
xnor UO_824 (O_824,N_4981,N_4937);
or UO_825 (O_825,N_4981,N_4997);
or UO_826 (O_826,N_4951,N_4987);
or UO_827 (O_827,N_4921,N_4971);
nand UO_828 (O_828,N_4916,N_4956);
nand UO_829 (O_829,N_4938,N_4910);
or UO_830 (O_830,N_4977,N_4927);
and UO_831 (O_831,N_4979,N_4991);
nor UO_832 (O_832,N_4953,N_4918);
nor UO_833 (O_833,N_4988,N_4950);
and UO_834 (O_834,N_4912,N_4972);
or UO_835 (O_835,N_4996,N_4980);
and UO_836 (O_836,N_4913,N_4914);
or UO_837 (O_837,N_4987,N_4941);
or UO_838 (O_838,N_4928,N_4927);
or UO_839 (O_839,N_4950,N_4992);
or UO_840 (O_840,N_4923,N_4945);
nand UO_841 (O_841,N_4936,N_4952);
or UO_842 (O_842,N_4936,N_4972);
xor UO_843 (O_843,N_4923,N_4964);
xor UO_844 (O_844,N_4924,N_4978);
and UO_845 (O_845,N_4904,N_4992);
nand UO_846 (O_846,N_4911,N_4982);
nor UO_847 (O_847,N_4910,N_4961);
and UO_848 (O_848,N_4923,N_4996);
nand UO_849 (O_849,N_4944,N_4997);
and UO_850 (O_850,N_4977,N_4993);
nor UO_851 (O_851,N_4908,N_4986);
or UO_852 (O_852,N_4961,N_4958);
nand UO_853 (O_853,N_4931,N_4933);
nor UO_854 (O_854,N_4964,N_4903);
nand UO_855 (O_855,N_4956,N_4976);
nand UO_856 (O_856,N_4954,N_4994);
or UO_857 (O_857,N_4916,N_4903);
nor UO_858 (O_858,N_4941,N_4952);
and UO_859 (O_859,N_4935,N_4918);
xor UO_860 (O_860,N_4982,N_4954);
nand UO_861 (O_861,N_4967,N_4962);
nand UO_862 (O_862,N_4954,N_4979);
nand UO_863 (O_863,N_4977,N_4911);
or UO_864 (O_864,N_4999,N_4959);
nor UO_865 (O_865,N_4950,N_4945);
nor UO_866 (O_866,N_4982,N_4988);
nand UO_867 (O_867,N_4987,N_4982);
nand UO_868 (O_868,N_4945,N_4942);
nand UO_869 (O_869,N_4939,N_4909);
or UO_870 (O_870,N_4946,N_4907);
and UO_871 (O_871,N_4953,N_4921);
or UO_872 (O_872,N_4945,N_4919);
nor UO_873 (O_873,N_4983,N_4910);
and UO_874 (O_874,N_4946,N_4965);
and UO_875 (O_875,N_4930,N_4951);
and UO_876 (O_876,N_4992,N_4913);
and UO_877 (O_877,N_4944,N_4959);
nor UO_878 (O_878,N_4965,N_4989);
and UO_879 (O_879,N_4923,N_4913);
and UO_880 (O_880,N_4975,N_4922);
xor UO_881 (O_881,N_4992,N_4944);
or UO_882 (O_882,N_4910,N_4904);
nand UO_883 (O_883,N_4925,N_4907);
nand UO_884 (O_884,N_4911,N_4974);
or UO_885 (O_885,N_4978,N_4927);
nand UO_886 (O_886,N_4935,N_4946);
nor UO_887 (O_887,N_4920,N_4981);
and UO_888 (O_888,N_4997,N_4931);
xor UO_889 (O_889,N_4939,N_4917);
nor UO_890 (O_890,N_4993,N_4984);
nand UO_891 (O_891,N_4932,N_4992);
nor UO_892 (O_892,N_4912,N_4954);
nand UO_893 (O_893,N_4922,N_4909);
and UO_894 (O_894,N_4906,N_4954);
or UO_895 (O_895,N_4955,N_4935);
and UO_896 (O_896,N_4952,N_4962);
xor UO_897 (O_897,N_4944,N_4911);
xor UO_898 (O_898,N_4907,N_4908);
nand UO_899 (O_899,N_4957,N_4930);
and UO_900 (O_900,N_4934,N_4912);
nand UO_901 (O_901,N_4943,N_4979);
nor UO_902 (O_902,N_4930,N_4992);
and UO_903 (O_903,N_4919,N_4977);
nand UO_904 (O_904,N_4917,N_4948);
or UO_905 (O_905,N_4930,N_4933);
nand UO_906 (O_906,N_4978,N_4948);
nand UO_907 (O_907,N_4910,N_4967);
nor UO_908 (O_908,N_4920,N_4950);
or UO_909 (O_909,N_4996,N_4940);
or UO_910 (O_910,N_4946,N_4963);
and UO_911 (O_911,N_4996,N_4947);
nand UO_912 (O_912,N_4904,N_4939);
nor UO_913 (O_913,N_4988,N_4915);
nand UO_914 (O_914,N_4971,N_4942);
or UO_915 (O_915,N_4974,N_4953);
or UO_916 (O_916,N_4923,N_4935);
nor UO_917 (O_917,N_4972,N_4901);
or UO_918 (O_918,N_4966,N_4971);
or UO_919 (O_919,N_4906,N_4978);
xor UO_920 (O_920,N_4901,N_4966);
or UO_921 (O_921,N_4985,N_4958);
nand UO_922 (O_922,N_4914,N_4918);
and UO_923 (O_923,N_4955,N_4961);
nor UO_924 (O_924,N_4933,N_4935);
or UO_925 (O_925,N_4929,N_4940);
xor UO_926 (O_926,N_4962,N_4970);
xnor UO_927 (O_927,N_4934,N_4922);
and UO_928 (O_928,N_4977,N_4933);
or UO_929 (O_929,N_4951,N_4923);
nand UO_930 (O_930,N_4988,N_4930);
nor UO_931 (O_931,N_4941,N_4900);
xor UO_932 (O_932,N_4985,N_4906);
nor UO_933 (O_933,N_4948,N_4960);
nor UO_934 (O_934,N_4959,N_4942);
nand UO_935 (O_935,N_4990,N_4918);
nand UO_936 (O_936,N_4921,N_4969);
nor UO_937 (O_937,N_4982,N_4972);
nor UO_938 (O_938,N_4954,N_4945);
and UO_939 (O_939,N_4941,N_4963);
nor UO_940 (O_940,N_4979,N_4949);
and UO_941 (O_941,N_4915,N_4901);
nand UO_942 (O_942,N_4947,N_4936);
nor UO_943 (O_943,N_4937,N_4916);
and UO_944 (O_944,N_4974,N_4963);
or UO_945 (O_945,N_4950,N_4931);
xnor UO_946 (O_946,N_4933,N_4922);
nand UO_947 (O_947,N_4913,N_4903);
nand UO_948 (O_948,N_4972,N_4938);
xor UO_949 (O_949,N_4956,N_4957);
nand UO_950 (O_950,N_4928,N_4923);
or UO_951 (O_951,N_4922,N_4903);
xnor UO_952 (O_952,N_4904,N_4900);
nand UO_953 (O_953,N_4955,N_4980);
nor UO_954 (O_954,N_4955,N_4959);
nor UO_955 (O_955,N_4945,N_4964);
or UO_956 (O_956,N_4937,N_4935);
and UO_957 (O_957,N_4955,N_4905);
nor UO_958 (O_958,N_4940,N_4947);
or UO_959 (O_959,N_4910,N_4985);
nor UO_960 (O_960,N_4929,N_4963);
nor UO_961 (O_961,N_4901,N_4962);
nor UO_962 (O_962,N_4978,N_4950);
xnor UO_963 (O_963,N_4942,N_4943);
nor UO_964 (O_964,N_4977,N_4931);
nand UO_965 (O_965,N_4969,N_4985);
nand UO_966 (O_966,N_4900,N_4927);
or UO_967 (O_967,N_4978,N_4934);
nand UO_968 (O_968,N_4930,N_4923);
xnor UO_969 (O_969,N_4936,N_4962);
nand UO_970 (O_970,N_4934,N_4955);
xnor UO_971 (O_971,N_4965,N_4901);
nand UO_972 (O_972,N_4987,N_4912);
nor UO_973 (O_973,N_4960,N_4959);
nor UO_974 (O_974,N_4943,N_4903);
nor UO_975 (O_975,N_4944,N_4918);
xnor UO_976 (O_976,N_4946,N_4924);
and UO_977 (O_977,N_4973,N_4914);
xor UO_978 (O_978,N_4988,N_4946);
and UO_979 (O_979,N_4902,N_4946);
and UO_980 (O_980,N_4954,N_4973);
or UO_981 (O_981,N_4978,N_4998);
or UO_982 (O_982,N_4995,N_4920);
nand UO_983 (O_983,N_4905,N_4979);
or UO_984 (O_984,N_4960,N_4907);
or UO_985 (O_985,N_4921,N_4935);
and UO_986 (O_986,N_4926,N_4961);
nand UO_987 (O_987,N_4932,N_4993);
nand UO_988 (O_988,N_4924,N_4980);
and UO_989 (O_989,N_4972,N_4962);
xnor UO_990 (O_990,N_4910,N_4945);
nor UO_991 (O_991,N_4917,N_4920);
or UO_992 (O_992,N_4929,N_4951);
and UO_993 (O_993,N_4978,N_4930);
nor UO_994 (O_994,N_4928,N_4972);
nor UO_995 (O_995,N_4999,N_4981);
xor UO_996 (O_996,N_4920,N_4921);
nand UO_997 (O_997,N_4932,N_4938);
and UO_998 (O_998,N_4905,N_4969);
and UO_999 (O_999,N_4969,N_4948);
endmodule