module basic_750_5000_1000_50_levels_1xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
xnor U0 (N_0,In_706,In_311);
and U1 (N_1,In_699,In_423);
or U2 (N_2,In_263,In_581);
nand U3 (N_3,In_521,In_181);
or U4 (N_4,In_590,In_55);
and U5 (N_5,In_541,In_461);
nor U6 (N_6,In_632,In_663);
nor U7 (N_7,In_719,In_738);
nand U8 (N_8,In_450,In_379);
nor U9 (N_9,In_582,In_146);
nor U10 (N_10,In_748,In_315);
nor U11 (N_11,In_256,In_71);
nor U12 (N_12,In_275,In_444);
nand U13 (N_13,In_395,In_64);
nor U14 (N_14,In_287,In_208);
or U15 (N_15,In_668,In_333);
nor U16 (N_16,In_204,In_222);
and U17 (N_17,In_407,In_231);
nor U18 (N_18,In_303,In_614);
nor U19 (N_19,In_368,In_485);
nand U20 (N_20,In_118,In_726);
and U21 (N_21,In_587,In_735);
and U22 (N_22,In_631,In_0);
nand U23 (N_23,In_202,In_106);
nand U24 (N_24,In_563,In_459);
nand U25 (N_25,In_388,In_438);
nor U26 (N_26,In_649,In_361);
nand U27 (N_27,In_504,In_480);
or U28 (N_28,In_416,In_651);
nor U29 (N_29,In_434,In_348);
nand U30 (N_30,In_321,In_548);
nor U31 (N_31,In_397,In_694);
nand U32 (N_32,In_575,In_137);
nand U33 (N_33,In_286,In_13);
nor U34 (N_34,In_210,In_441);
nor U35 (N_35,In_383,In_598);
nor U36 (N_36,In_377,In_96);
nand U37 (N_37,In_712,In_661);
nor U38 (N_38,In_620,In_662);
nand U39 (N_39,In_513,In_595);
and U40 (N_40,In_469,In_299);
nand U41 (N_41,In_338,In_10);
or U42 (N_42,In_544,In_401);
nor U43 (N_43,In_33,In_746);
nand U44 (N_44,In_345,In_269);
nand U45 (N_45,In_696,In_253);
nor U46 (N_46,In_515,In_678);
nor U47 (N_47,In_390,In_260);
nand U48 (N_48,In_81,In_335);
nor U49 (N_49,In_145,In_46);
nor U50 (N_50,In_105,In_221);
or U51 (N_51,In_178,In_498);
nand U52 (N_52,In_346,In_182);
or U53 (N_53,In_683,In_215);
nor U54 (N_54,In_610,In_101);
nor U55 (N_55,In_670,In_41);
and U56 (N_56,In_56,In_98);
and U57 (N_57,In_418,In_657);
nor U58 (N_58,In_642,In_23);
nand U59 (N_59,In_391,In_396);
nand U60 (N_60,In_337,In_91);
nand U61 (N_61,In_555,In_659);
and U62 (N_62,In_262,In_163);
or U63 (N_63,In_705,In_51);
nand U64 (N_64,In_453,In_591);
or U65 (N_65,In_609,In_433);
nand U66 (N_66,In_367,In_325);
nor U67 (N_67,In_95,In_148);
and U68 (N_68,In_162,In_568);
nand U69 (N_69,In_8,In_490);
and U70 (N_70,In_271,In_314);
or U71 (N_71,In_213,In_429);
and U72 (N_72,In_186,In_627);
or U73 (N_73,In_421,In_7);
and U74 (N_74,In_528,In_704);
and U75 (N_75,In_280,In_261);
nor U76 (N_76,In_184,In_736);
nor U77 (N_77,In_608,In_681);
and U78 (N_78,In_349,In_107);
and U79 (N_79,In_402,In_328);
nand U80 (N_80,In_18,In_359);
or U81 (N_81,In_20,In_722);
nand U82 (N_82,In_266,In_482);
and U83 (N_83,In_339,In_693);
and U84 (N_84,In_87,In_400);
or U85 (N_85,In_296,In_411);
or U86 (N_86,In_16,In_237);
or U87 (N_87,In_239,In_422);
nand U88 (N_88,In_243,In_641);
and U89 (N_89,In_537,In_47);
xnor U90 (N_90,In_473,In_656);
nand U91 (N_91,In_257,In_652);
and U92 (N_92,In_268,In_218);
and U93 (N_93,In_398,In_102);
nor U94 (N_94,In_448,In_604);
or U95 (N_95,In_153,In_113);
nor U96 (N_96,In_110,In_192);
nand U97 (N_97,In_284,In_82);
or U98 (N_98,In_466,In_464);
xnor U99 (N_99,In_564,In_512);
nand U100 (N_100,In_35,In_516);
or U101 (N_101,In_496,In_507);
xnor U102 (N_102,In_252,In_530);
nand U103 (N_103,In_617,In_574);
nor U104 (N_104,In_517,N_44);
or U105 (N_105,In_440,In_19);
nor U106 (N_106,In_612,N_88);
nor U107 (N_107,In_535,In_130);
nor U108 (N_108,In_191,N_0);
or U109 (N_109,In_447,N_74);
nor U110 (N_110,In_38,In_320);
and U111 (N_111,In_616,In_393);
and U112 (N_112,In_144,In_281);
and U113 (N_113,In_352,In_723);
nor U114 (N_114,In_242,In_37);
nand U115 (N_115,In_588,In_212);
or U116 (N_116,In_224,In_539);
and U117 (N_117,In_427,In_131);
or U118 (N_118,In_700,In_86);
nor U119 (N_119,N_21,In_749);
nand U120 (N_120,In_625,In_417);
and U121 (N_121,In_549,In_59);
nor U122 (N_122,In_29,In_295);
and U123 (N_123,In_351,In_54);
or U124 (N_124,In_120,In_386);
or U125 (N_125,In_36,In_119);
and U126 (N_126,In_501,In_665);
and U127 (N_127,In_394,In_578);
nor U128 (N_128,In_254,N_49);
or U129 (N_129,In_527,In_139);
and U130 (N_130,In_474,In_565);
and U131 (N_131,In_621,In_207);
nand U132 (N_132,In_72,In_688);
and U133 (N_133,In_514,In_2);
or U134 (N_134,In_274,In_430);
nor U135 (N_135,In_716,In_660);
nand U136 (N_136,In_276,In_741);
and U137 (N_137,In_292,In_463);
and U138 (N_138,In_158,In_554);
nand U139 (N_139,In_135,In_682);
and U140 (N_140,In_166,In_97);
nor U141 (N_141,In_586,In_371);
or U142 (N_142,In_70,In_489);
and U143 (N_143,In_109,In_691);
nand U144 (N_144,N_91,N_28);
and U145 (N_145,In_518,In_99);
or U146 (N_146,In_606,In_698);
and U147 (N_147,In_572,In_15);
nor U148 (N_148,N_84,In_194);
and U149 (N_149,In_701,In_420);
nand U150 (N_150,In_6,In_225);
or U151 (N_151,In_585,In_45);
or U152 (N_152,In_509,In_354);
nor U153 (N_153,In_477,In_172);
or U154 (N_154,In_249,In_357);
and U155 (N_155,In_643,In_344);
or U156 (N_156,In_745,In_143);
nor U157 (N_157,In_532,N_99);
nor U158 (N_158,N_63,N_9);
nor U159 (N_159,In_493,In_471);
nor U160 (N_160,In_577,N_57);
nand U161 (N_161,In_410,In_687);
nand U162 (N_162,In_714,In_63);
and U163 (N_163,In_123,In_251);
and U164 (N_164,In_510,In_80);
nand U165 (N_165,In_245,In_435);
nor U166 (N_166,In_319,In_503);
nand U167 (N_167,In_707,In_330);
or U168 (N_168,In_511,In_39);
nor U169 (N_169,In_27,In_446);
and U170 (N_170,In_155,In_169);
or U171 (N_171,N_39,In_179);
nor U172 (N_172,In_298,In_497);
nor U173 (N_173,In_232,In_68);
nor U174 (N_174,In_538,In_385);
nand U175 (N_175,In_556,In_236);
or U176 (N_176,In_347,N_41);
or U177 (N_177,In_52,In_133);
xor U178 (N_178,In_671,In_138);
nor U179 (N_179,In_93,N_30);
nand U180 (N_180,In_605,In_200);
or U181 (N_181,N_45,In_432);
and U182 (N_182,In_533,In_536);
nand U183 (N_183,N_47,In_654);
or U184 (N_184,N_7,In_358);
nor U185 (N_185,In_28,In_710);
nand U186 (N_186,In_505,N_69);
or U187 (N_187,In_404,N_6);
nor U188 (N_188,In_522,In_740);
or U189 (N_189,In_553,In_487);
and U190 (N_190,In_676,In_645);
or U191 (N_191,In_278,In_409);
and U192 (N_192,N_38,In_32);
nor U193 (N_193,In_680,In_175);
and U194 (N_194,In_437,In_206);
or U195 (N_195,In_89,In_664);
and U196 (N_196,In_531,In_164);
or U197 (N_197,In_452,In_326);
nor U198 (N_198,N_92,In_729);
nand U199 (N_199,In_331,In_114);
or U200 (N_200,In_579,N_188);
and U201 (N_201,N_148,In_1);
or U202 (N_202,In_50,N_153);
nand U203 (N_203,In_301,In_62);
or U204 (N_204,In_14,N_97);
nor U205 (N_205,In_695,In_336);
nand U206 (N_206,In_195,In_626);
or U207 (N_207,N_197,In_742);
nand U208 (N_208,In_403,In_499);
xor U209 (N_209,In_647,In_264);
and U210 (N_210,N_124,In_566);
or U211 (N_211,N_105,In_26);
nor U212 (N_212,In_159,N_145);
and U213 (N_213,In_711,N_120);
or U214 (N_214,In_188,In_183);
nor U215 (N_215,N_166,In_355);
nand U216 (N_216,N_118,In_732);
or U217 (N_217,In_546,In_140);
or U218 (N_218,N_24,In_177);
nor U219 (N_219,N_36,In_61);
and U220 (N_220,In_628,N_131);
nand U221 (N_221,N_146,In_132);
nor U222 (N_222,N_196,In_115);
or U223 (N_223,In_77,N_158);
and U224 (N_224,In_378,N_50);
xor U225 (N_225,N_156,N_85);
nand U226 (N_226,In_289,In_74);
nor U227 (N_227,In_112,In_279);
or U228 (N_228,In_273,N_35);
nor U229 (N_229,In_350,In_679);
and U230 (N_230,In_34,In_734);
or U231 (N_231,N_154,In_715);
or U232 (N_232,In_88,In_288);
and U233 (N_233,In_644,In_247);
and U234 (N_234,N_14,In_265);
nor U235 (N_235,In_633,In_58);
or U236 (N_236,In_483,In_443);
and U237 (N_237,N_1,N_51);
nand U238 (N_238,In_241,In_316);
nand U239 (N_239,N_139,N_187);
nand U240 (N_240,In_436,N_182);
nand U241 (N_241,In_309,N_185);
or U242 (N_242,In_545,N_109);
and U243 (N_243,N_104,In_669);
nor U244 (N_244,In_743,In_601);
nor U245 (N_245,In_117,In_467);
or U246 (N_246,In_76,N_167);
nor U247 (N_247,In_53,In_342);
or U248 (N_248,In_160,N_161);
nand U249 (N_249,N_168,In_233);
and U250 (N_250,In_561,In_214);
nand U251 (N_251,In_454,N_195);
and U252 (N_252,In_307,In_363);
and U253 (N_253,N_180,In_650);
or U254 (N_254,N_67,In_703);
or U255 (N_255,N_133,N_172);
nor U256 (N_256,In_376,In_629);
nand U257 (N_257,In_709,In_424);
nand U258 (N_258,N_94,In_580);
nand U259 (N_259,In_686,In_25);
nor U260 (N_260,N_140,In_306);
nand U261 (N_261,In_460,In_674);
and U262 (N_262,In_730,In_111);
nor U263 (N_263,In_685,N_58);
or U264 (N_264,In_476,In_108);
or U265 (N_265,In_360,N_198);
or U266 (N_266,In_92,In_619);
nand U267 (N_267,In_57,N_117);
nand U268 (N_268,N_129,In_67);
nand U269 (N_269,N_113,N_165);
or U270 (N_270,In_189,In_180);
or U271 (N_271,In_468,In_744);
nand U272 (N_272,In_380,N_40);
nand U273 (N_273,In_285,In_211);
nor U274 (N_274,In_121,N_80);
nor U275 (N_275,In_557,N_46);
nor U276 (N_276,In_79,In_250);
and U277 (N_277,N_181,In_203);
nor U278 (N_278,In_12,In_584);
nor U279 (N_279,N_29,N_27);
or U280 (N_280,In_638,In_141);
or U281 (N_281,N_83,In_603);
or U282 (N_282,In_73,In_151);
or U283 (N_283,In_428,In_727);
nor U284 (N_284,N_81,In_611);
and U285 (N_285,In_646,N_60);
and U286 (N_286,N_56,In_724);
nand U287 (N_287,N_8,In_282);
nand U288 (N_288,N_141,N_98);
or U289 (N_289,N_25,N_134);
nor U290 (N_290,In_653,In_547);
and U291 (N_291,N_71,N_11);
nor U292 (N_292,In_370,N_16);
nor U293 (N_293,N_76,In_90);
and U294 (N_294,N_137,In_502);
or U295 (N_295,In_85,In_475);
xnor U296 (N_296,In_323,In_83);
nand U297 (N_297,In_365,In_472);
nor U298 (N_298,In_374,In_419);
nor U299 (N_299,In_602,N_171);
nor U300 (N_300,In_562,N_86);
nand U301 (N_301,In_217,N_123);
and U302 (N_302,In_353,N_192);
and U303 (N_303,In_43,In_341);
and U304 (N_304,N_163,N_136);
nand U305 (N_305,In_640,N_82);
or U306 (N_306,N_240,In_75);
nand U307 (N_307,In_465,In_228);
nand U308 (N_308,In_220,In_542);
nor U309 (N_309,In_666,N_62);
nor U310 (N_310,N_110,N_194);
and U311 (N_311,N_255,In_226);
and U312 (N_312,N_103,In_31);
and U313 (N_313,In_318,N_270);
nor U314 (N_314,N_13,N_273);
and U315 (N_315,In_550,In_291);
and U316 (N_316,In_94,N_100);
and U317 (N_317,In_387,In_30);
and U318 (N_318,N_252,N_249);
or U319 (N_319,In_731,N_253);
or U320 (N_320,In_40,N_48);
and U321 (N_321,N_132,In_322);
or U322 (N_322,N_298,In_142);
and U323 (N_323,N_201,N_234);
or U324 (N_324,In_634,N_257);
nand U325 (N_325,In_702,N_17);
nor U326 (N_326,In_607,In_240);
and U327 (N_327,N_89,N_66);
and U328 (N_328,In_488,In_630);
nor U329 (N_329,In_364,In_571);
or U330 (N_330,N_26,N_111);
or U331 (N_331,In_413,N_152);
or U332 (N_332,N_242,N_101);
and U333 (N_333,In_576,N_55);
nand U334 (N_334,In_495,N_200);
and U335 (N_335,In_399,N_293);
or U336 (N_336,In_462,N_233);
nor U337 (N_337,In_11,In_149);
and U338 (N_338,In_150,N_119);
nor U339 (N_339,N_149,In_270);
nor U340 (N_340,N_176,N_73);
and U341 (N_341,In_372,In_412);
and U342 (N_342,In_343,N_268);
nor U343 (N_343,N_169,N_157);
and U344 (N_344,In_733,In_718);
or U345 (N_345,N_170,In_21);
or U346 (N_346,In_84,In_312);
and U347 (N_347,N_70,N_178);
nand U348 (N_348,N_212,N_90);
and U349 (N_349,In_229,In_558);
nor U350 (N_350,In_272,In_324);
and U351 (N_351,In_508,In_523);
nor U352 (N_352,N_217,N_205);
nand U353 (N_353,In_543,N_262);
nor U354 (N_354,N_292,N_228);
nand U355 (N_355,In_613,In_304);
or U356 (N_356,In_478,N_155);
and U357 (N_357,In_173,In_171);
nor U358 (N_358,N_238,In_49);
and U359 (N_359,In_449,In_725);
nand U360 (N_360,N_230,In_655);
and U361 (N_361,N_202,In_238);
and U362 (N_362,N_210,N_175);
nor U363 (N_363,N_229,In_219);
and U364 (N_364,In_290,In_414);
nor U365 (N_365,In_300,N_289);
and U366 (N_366,In_672,In_161);
nor U367 (N_367,N_236,In_246);
or U368 (N_368,In_277,In_3);
nor U369 (N_369,N_75,In_332);
and U370 (N_370,N_115,N_79);
and U371 (N_371,In_293,In_305);
nand U372 (N_372,N_121,In_78);
nand U373 (N_373,In_494,In_524);
or U374 (N_374,N_125,In_392);
nand U375 (N_375,N_280,N_281);
or U376 (N_376,N_43,In_259);
nor U377 (N_377,In_570,N_199);
nor U378 (N_378,In_5,In_356);
nor U379 (N_379,N_226,In_381);
nand U380 (N_380,In_308,In_244);
or U381 (N_381,N_204,N_183);
nor U382 (N_382,In_116,N_128);
and U383 (N_383,In_22,N_61);
and U384 (N_384,In_129,In_622);
nor U385 (N_385,N_15,In_185);
or U386 (N_386,In_136,In_66);
nand U387 (N_387,In_205,N_247);
nor U388 (N_388,N_122,N_297);
or U389 (N_389,N_151,In_567);
or U390 (N_390,N_34,In_534);
nand U391 (N_391,In_248,In_190);
nand U392 (N_392,In_167,N_162);
and U393 (N_393,N_108,In_431);
and U394 (N_394,In_60,In_624);
and U395 (N_395,In_594,N_211);
or U396 (N_396,In_481,In_648);
or U397 (N_397,N_18,N_215);
or U398 (N_398,In_201,In_593);
and U399 (N_399,In_708,N_4);
nor U400 (N_400,N_224,N_312);
or U401 (N_401,N_106,N_317);
nor U402 (N_402,In_17,In_442);
nand U403 (N_403,N_283,N_335);
nor U404 (N_404,N_279,N_184);
or U405 (N_405,In_728,In_405);
or U406 (N_406,N_87,N_397);
nand U407 (N_407,N_239,N_348);
xnor U408 (N_408,In_334,In_170);
and U409 (N_409,In_426,N_254);
or U410 (N_410,N_301,N_150);
or U411 (N_411,N_364,N_302);
and U412 (N_412,N_33,N_322);
and U413 (N_413,N_223,In_589);
nor U414 (N_414,In_599,N_393);
nor U415 (N_415,N_388,N_386);
nor U416 (N_416,In_552,N_263);
nand U417 (N_417,N_275,In_445);
nor U418 (N_418,In_526,N_160);
nand U419 (N_419,In_124,N_107);
or U420 (N_420,N_313,N_306);
nor U421 (N_421,N_272,N_59);
nand U422 (N_422,N_295,N_357);
nor U423 (N_423,N_339,N_307);
or U424 (N_424,N_328,In_470);
nand U425 (N_425,In_637,N_334);
nor U426 (N_426,In_455,N_315);
nor U427 (N_427,N_367,N_112);
nor U428 (N_428,N_353,N_12);
and U429 (N_429,In_618,N_218);
nor U430 (N_430,N_330,N_299);
or U431 (N_431,N_95,In_313);
nand U432 (N_432,In_600,In_174);
nand U433 (N_433,In_500,N_383);
and U434 (N_434,In_255,In_747);
xnor U435 (N_435,N_189,In_366);
nor U436 (N_436,N_277,N_379);
or U437 (N_437,N_395,N_311);
nand U438 (N_438,In_415,In_152);
or U439 (N_439,In_48,In_597);
nand U440 (N_440,N_102,In_187);
or U441 (N_441,In_491,In_327);
and U442 (N_442,N_159,In_44);
nor U443 (N_443,In_283,N_333);
nand U444 (N_444,In_223,In_689);
or U445 (N_445,N_237,N_243);
nor U446 (N_446,In_439,N_220);
and U447 (N_447,N_193,In_739);
or U448 (N_448,In_165,N_314);
and U449 (N_449,N_331,N_389);
or U450 (N_450,N_22,In_134);
nor U451 (N_451,N_37,N_68);
nand U452 (N_452,N_374,N_207);
xor U453 (N_453,N_93,In_690);
and U454 (N_454,N_2,In_122);
and U455 (N_455,N_227,In_596);
or U456 (N_456,N_221,In_677);
nor U457 (N_457,In_559,N_271);
nor U458 (N_458,In_569,In_451);
nand U459 (N_459,N_250,N_274);
and U460 (N_460,N_241,N_355);
or U461 (N_461,N_208,In_636);
nor U462 (N_462,In_198,In_127);
nand U463 (N_463,N_341,N_318);
nand U464 (N_464,N_349,N_360);
or U465 (N_465,N_179,N_376);
nand U466 (N_466,N_394,N_219);
nand U467 (N_467,In_721,N_251);
nand U468 (N_468,In_329,N_351);
and U469 (N_469,In_147,In_667);
and U470 (N_470,N_248,In_103);
or U471 (N_471,N_303,N_350);
nor U472 (N_472,In_294,N_373);
or U473 (N_473,In_4,In_484);
or U474 (N_474,N_372,N_365);
nor U475 (N_475,N_391,N_324);
nor U476 (N_476,N_377,N_147);
nand U477 (N_477,In_128,In_551);
or U478 (N_478,N_356,N_143);
or U479 (N_479,N_256,N_231);
and U480 (N_480,N_296,N_177);
or U481 (N_481,N_269,N_266);
or U482 (N_482,In_373,N_327);
nor U483 (N_483,In_227,In_486);
nor U484 (N_484,N_368,In_267);
and U485 (N_485,N_309,N_130);
and U486 (N_486,N_378,N_282);
and U487 (N_487,N_325,N_232);
or U488 (N_488,N_78,In_458);
and U489 (N_489,N_338,N_114);
or U490 (N_490,In_382,In_197);
nand U491 (N_491,N_290,N_343);
or U492 (N_492,N_265,N_291);
or U493 (N_493,In_456,N_213);
and U494 (N_494,N_332,In_24);
nor U495 (N_495,In_375,In_492);
nand U496 (N_496,In_408,N_278);
nor U497 (N_497,In_302,N_387);
and U498 (N_498,N_305,In_635);
nand U499 (N_499,N_244,N_5);
or U500 (N_500,N_418,N_408);
nand U501 (N_501,N_401,N_412);
nand U502 (N_502,N_415,N_403);
nand U503 (N_503,In_9,N_435);
and U504 (N_504,N_96,N_382);
nor U505 (N_505,N_116,N_428);
nor U506 (N_506,N_450,In_168);
or U507 (N_507,N_42,N_261);
or U508 (N_508,N_20,N_260);
and U509 (N_509,N_246,N_484);
nor U510 (N_510,N_362,N_422);
nand U511 (N_511,N_441,N_476);
or U512 (N_512,N_451,N_380);
nor U513 (N_513,N_358,N_459);
or U514 (N_514,N_354,N_416);
nand U515 (N_515,In_583,In_525);
or U516 (N_516,N_498,N_430);
nand U517 (N_517,N_321,N_225);
or U518 (N_518,N_398,In_615);
nor U519 (N_519,N_77,N_493);
or U520 (N_520,In_310,N_319);
or U521 (N_521,N_497,N_467);
nand U522 (N_522,In_234,N_65);
nor U523 (N_523,N_456,N_471);
nand U524 (N_524,N_320,N_491);
nor U525 (N_525,N_359,N_53);
nand U526 (N_526,N_442,N_481);
nand U527 (N_527,N_490,In_230);
nor U528 (N_528,N_209,N_431);
or U529 (N_529,N_72,In_209);
and U530 (N_530,N_344,In_479);
and U531 (N_531,In_216,N_345);
and U532 (N_532,N_138,N_433);
nand U533 (N_533,N_477,N_417);
or U534 (N_534,In_156,N_499);
and U535 (N_535,N_144,In_69);
and U536 (N_536,N_457,In_713);
or U537 (N_537,N_323,N_52);
nand U538 (N_538,N_142,In_125);
and U539 (N_539,N_173,In_457);
and U540 (N_540,N_494,N_402);
nand U541 (N_541,N_361,N_485);
nor U542 (N_542,In_369,N_429);
and U543 (N_543,N_288,N_326);
or U544 (N_544,N_448,N_424);
nand U545 (N_545,N_342,N_206);
nand U546 (N_546,N_347,N_437);
nor U547 (N_547,N_258,N_474);
nand U548 (N_548,In_100,In_529);
nand U549 (N_549,N_411,N_407);
nand U550 (N_550,N_3,N_190);
or U551 (N_551,In_717,N_245);
nor U552 (N_552,N_458,In_675);
or U553 (N_553,N_370,N_473);
nor U554 (N_554,N_443,N_464);
and U555 (N_555,In_639,N_495);
and U556 (N_556,In_519,N_409);
nor U557 (N_557,In_154,N_284);
and U558 (N_558,N_135,In_196);
nor U559 (N_559,In_592,N_423);
or U560 (N_560,In_697,N_436);
nand U561 (N_561,N_316,N_465);
and U562 (N_562,N_216,In_126);
nand U563 (N_563,N_304,In_235);
nand U564 (N_564,In_623,In_658);
nor U565 (N_565,N_414,N_308);
and U566 (N_566,In_199,N_492);
nand U567 (N_567,N_427,N_445);
or U568 (N_568,N_23,N_426);
or U569 (N_569,N_405,In_425);
and U570 (N_570,N_438,N_384);
or U571 (N_571,N_466,In_673);
nand U572 (N_572,N_410,N_419);
or U573 (N_573,N_329,N_340);
and U574 (N_574,N_310,N_214);
and U575 (N_575,N_287,N_32);
nor U576 (N_576,N_267,N_406);
nor U577 (N_577,N_432,N_276);
nor U578 (N_578,N_186,N_174);
or U579 (N_579,In_104,N_449);
or U580 (N_580,N_390,N_126);
nand U581 (N_581,N_396,N_453);
and U582 (N_582,N_454,N_480);
or U583 (N_583,N_337,N_294);
nor U584 (N_584,N_420,In_340);
or U585 (N_585,N_468,N_375);
or U586 (N_586,N_352,N_444);
or U587 (N_587,N_203,N_164);
or U588 (N_588,N_439,In_720);
nand U589 (N_589,N_235,N_447);
or U590 (N_590,N_483,N_434);
nand U591 (N_591,N_300,N_404);
nor U592 (N_592,In_540,N_19);
nor U593 (N_593,In_193,N_496);
and U594 (N_594,N_222,N_472);
and U595 (N_595,N_475,N_463);
nor U596 (N_596,In_176,N_421);
nor U597 (N_597,N_286,N_455);
or U598 (N_598,In_384,N_127);
nand U599 (N_599,N_191,N_489);
nor U600 (N_600,N_574,N_577);
and U601 (N_601,N_371,N_583);
or U602 (N_602,In_520,N_509);
nand U603 (N_603,N_599,N_580);
nor U604 (N_604,N_576,N_536);
nor U605 (N_605,N_558,N_488);
and U606 (N_606,N_595,N_529);
nor U607 (N_607,N_392,N_446);
nand U608 (N_608,N_522,N_578);
nor U609 (N_609,N_64,N_561);
nor U610 (N_610,N_533,N_542);
and U611 (N_611,N_10,In_573);
and U612 (N_612,N_508,N_545);
nor U613 (N_613,N_546,N_518);
or U614 (N_614,N_535,N_461);
nand U615 (N_615,N_552,N_506);
nor U616 (N_616,N_523,N_385);
nor U617 (N_617,N_31,N_596);
and U618 (N_618,In_42,N_512);
xnor U619 (N_619,In_692,N_482);
and U620 (N_620,N_589,N_564);
nor U621 (N_621,N_400,In_362);
and U622 (N_622,N_515,N_530);
nand U623 (N_623,In_684,N_539);
nand U624 (N_624,N_514,N_503);
nor U625 (N_625,N_579,N_513);
or U626 (N_626,N_592,N_588);
nor U627 (N_627,N_548,N_547);
and U628 (N_628,N_469,In_65);
or U629 (N_629,N_525,N_336);
or U630 (N_630,N_487,N_590);
and U631 (N_631,N_366,N_584);
or U632 (N_632,N_502,N_516);
nand U633 (N_633,N_550,N_381);
nand U634 (N_634,N_532,N_527);
or U635 (N_635,N_544,N_537);
nor U636 (N_636,N_568,N_534);
and U637 (N_637,N_586,N_565);
nor U638 (N_638,N_553,N_582);
or U639 (N_639,N_470,N_399);
nor U640 (N_640,In_737,N_264);
or U641 (N_641,N_585,N_440);
and U642 (N_642,N_505,N_521);
xnor U643 (N_643,In_389,N_540);
nor U644 (N_644,N_507,N_541);
and U645 (N_645,N_519,N_581);
or U646 (N_646,N_598,N_478);
nor U647 (N_647,N_500,N_549);
or U648 (N_648,N_369,In_317);
or U649 (N_649,N_538,N_593);
nor U650 (N_650,N_425,N_560);
nor U651 (N_651,N_413,N_555);
or U652 (N_652,N_572,N_526);
nand U653 (N_653,N_524,N_566);
nor U654 (N_654,N_511,N_452);
and U655 (N_655,N_554,N_570);
nand U656 (N_656,N_543,N_556);
nor U657 (N_657,N_259,N_462);
and U658 (N_658,N_363,In_406);
or U659 (N_659,N_531,N_575);
or U660 (N_660,N_479,N_567);
and U661 (N_661,N_460,N_551);
nor U662 (N_662,N_591,N_285);
nand U663 (N_663,In_506,N_563);
or U664 (N_664,N_510,N_571);
or U665 (N_665,N_486,N_557);
and U666 (N_666,N_54,N_504);
and U667 (N_667,N_501,N_594);
nand U668 (N_668,N_573,N_559);
and U669 (N_669,N_562,N_517);
or U670 (N_670,N_587,N_597);
or U671 (N_671,N_346,In_560);
and U672 (N_672,N_528,In_157);
and U673 (N_673,N_520,In_258);
nor U674 (N_674,N_569,In_297);
nand U675 (N_675,In_684,N_259);
and U676 (N_676,N_520,N_586);
and U677 (N_677,N_526,N_569);
or U678 (N_678,N_548,N_591);
or U679 (N_679,N_425,N_385);
and U680 (N_680,N_578,N_594);
nand U681 (N_681,N_509,N_527);
and U682 (N_682,N_542,N_399);
nand U683 (N_683,N_573,N_563);
nand U684 (N_684,N_539,N_536);
nor U685 (N_685,N_381,N_517);
or U686 (N_686,N_564,N_54);
or U687 (N_687,N_392,N_525);
nand U688 (N_688,N_569,N_543);
or U689 (N_689,N_530,In_406);
or U690 (N_690,N_578,N_392);
and U691 (N_691,In_297,N_487);
xnor U692 (N_692,N_518,N_535);
nand U693 (N_693,N_478,N_461);
nor U694 (N_694,N_594,N_587);
and U695 (N_695,N_392,N_590);
or U696 (N_696,N_582,N_363);
and U697 (N_697,N_547,N_553);
nand U698 (N_698,In_297,N_505);
or U699 (N_699,N_578,N_513);
nor U700 (N_700,N_642,N_677);
nand U701 (N_701,N_616,N_669);
or U702 (N_702,N_637,N_639);
nand U703 (N_703,N_696,N_673);
nor U704 (N_704,N_623,N_627);
nand U705 (N_705,N_601,N_688);
or U706 (N_706,N_657,N_604);
or U707 (N_707,N_603,N_681);
or U708 (N_708,N_615,N_647);
and U709 (N_709,N_694,N_634);
or U710 (N_710,N_670,N_633);
nor U711 (N_711,N_625,N_624);
and U712 (N_712,N_687,N_632);
and U713 (N_713,N_679,N_619);
or U714 (N_714,N_658,N_664);
and U715 (N_715,N_644,N_651);
nand U716 (N_716,N_646,N_665);
nand U717 (N_717,N_661,N_611);
and U718 (N_718,N_649,N_675);
nor U719 (N_719,N_684,N_691);
and U720 (N_720,N_607,N_635);
nor U721 (N_721,N_693,N_683);
or U722 (N_722,N_648,N_671);
or U723 (N_723,N_645,N_695);
and U724 (N_724,N_667,N_660);
or U725 (N_725,N_600,N_656);
and U726 (N_726,N_638,N_653);
and U727 (N_727,N_608,N_622);
or U728 (N_728,N_609,N_655);
and U729 (N_729,N_663,N_666);
nor U730 (N_730,N_641,N_640);
or U731 (N_731,N_668,N_650);
or U732 (N_732,N_636,N_685);
or U733 (N_733,N_617,N_620);
nor U734 (N_734,N_626,N_606);
nand U735 (N_735,N_631,N_613);
nor U736 (N_736,N_662,N_698);
or U737 (N_737,N_630,N_674);
nand U738 (N_738,N_699,N_680);
or U739 (N_739,N_628,N_629);
nand U740 (N_740,N_612,N_697);
or U741 (N_741,N_672,N_614);
and U742 (N_742,N_654,N_689);
or U743 (N_743,N_682,N_692);
nand U744 (N_744,N_621,N_659);
nand U745 (N_745,N_618,N_652);
nand U746 (N_746,N_686,N_678);
nor U747 (N_747,N_605,N_610);
nor U748 (N_748,N_643,N_690);
or U749 (N_749,N_602,N_676);
nand U750 (N_750,N_683,N_660);
or U751 (N_751,N_680,N_613);
or U752 (N_752,N_632,N_685);
and U753 (N_753,N_643,N_680);
and U754 (N_754,N_694,N_690);
nand U755 (N_755,N_618,N_616);
or U756 (N_756,N_664,N_676);
or U757 (N_757,N_600,N_648);
nand U758 (N_758,N_667,N_675);
or U759 (N_759,N_685,N_613);
or U760 (N_760,N_699,N_636);
or U761 (N_761,N_675,N_658);
and U762 (N_762,N_639,N_683);
and U763 (N_763,N_656,N_650);
nor U764 (N_764,N_694,N_655);
nand U765 (N_765,N_659,N_669);
and U766 (N_766,N_698,N_666);
and U767 (N_767,N_680,N_688);
or U768 (N_768,N_608,N_666);
nand U769 (N_769,N_662,N_607);
nand U770 (N_770,N_619,N_613);
nor U771 (N_771,N_668,N_695);
or U772 (N_772,N_638,N_672);
and U773 (N_773,N_620,N_664);
nand U774 (N_774,N_616,N_634);
or U775 (N_775,N_670,N_644);
xor U776 (N_776,N_644,N_693);
nand U777 (N_777,N_619,N_612);
or U778 (N_778,N_658,N_622);
nor U779 (N_779,N_662,N_676);
and U780 (N_780,N_624,N_621);
nand U781 (N_781,N_662,N_642);
nor U782 (N_782,N_629,N_677);
and U783 (N_783,N_690,N_618);
nor U784 (N_784,N_611,N_601);
nand U785 (N_785,N_676,N_630);
nand U786 (N_786,N_626,N_611);
and U787 (N_787,N_635,N_615);
nand U788 (N_788,N_662,N_601);
and U789 (N_789,N_636,N_633);
and U790 (N_790,N_696,N_694);
nor U791 (N_791,N_683,N_618);
or U792 (N_792,N_694,N_695);
nand U793 (N_793,N_669,N_640);
and U794 (N_794,N_614,N_651);
nor U795 (N_795,N_673,N_636);
or U796 (N_796,N_679,N_628);
nand U797 (N_797,N_692,N_651);
nor U798 (N_798,N_602,N_690);
nand U799 (N_799,N_689,N_611);
and U800 (N_800,N_758,N_795);
and U801 (N_801,N_722,N_748);
and U802 (N_802,N_723,N_773);
and U803 (N_803,N_753,N_712);
nand U804 (N_804,N_741,N_793);
nand U805 (N_805,N_703,N_751);
nor U806 (N_806,N_791,N_755);
nor U807 (N_807,N_768,N_769);
or U808 (N_808,N_767,N_745);
nor U809 (N_809,N_777,N_772);
and U810 (N_810,N_770,N_775);
nand U811 (N_811,N_744,N_711);
nor U812 (N_812,N_771,N_766);
and U813 (N_813,N_797,N_798);
nand U814 (N_814,N_713,N_796);
or U815 (N_815,N_729,N_765);
and U816 (N_816,N_757,N_760);
nor U817 (N_817,N_727,N_756);
or U818 (N_818,N_776,N_794);
nand U819 (N_819,N_761,N_708);
nand U820 (N_820,N_759,N_732);
or U821 (N_821,N_785,N_763);
or U822 (N_822,N_743,N_783);
nor U823 (N_823,N_738,N_782);
and U824 (N_824,N_715,N_799);
or U825 (N_825,N_700,N_705);
or U826 (N_826,N_790,N_709);
nand U827 (N_827,N_707,N_778);
nor U828 (N_828,N_792,N_725);
and U829 (N_829,N_704,N_742);
or U830 (N_830,N_702,N_784);
nor U831 (N_831,N_749,N_726);
or U832 (N_832,N_746,N_733);
nand U833 (N_833,N_714,N_734);
nand U834 (N_834,N_780,N_728);
nor U835 (N_835,N_739,N_706);
or U836 (N_836,N_720,N_710);
nand U837 (N_837,N_718,N_736);
nor U838 (N_838,N_779,N_781);
or U839 (N_839,N_754,N_787);
and U840 (N_840,N_762,N_724);
nor U841 (N_841,N_701,N_716);
and U842 (N_842,N_788,N_750);
or U843 (N_843,N_789,N_730);
nand U844 (N_844,N_717,N_737);
nor U845 (N_845,N_735,N_786);
or U846 (N_846,N_764,N_719);
nand U847 (N_847,N_721,N_740);
nand U848 (N_848,N_774,N_747);
nor U849 (N_849,N_731,N_752);
or U850 (N_850,N_773,N_736);
or U851 (N_851,N_774,N_711);
or U852 (N_852,N_743,N_763);
or U853 (N_853,N_753,N_779);
nand U854 (N_854,N_725,N_731);
or U855 (N_855,N_766,N_712);
nand U856 (N_856,N_700,N_786);
nand U857 (N_857,N_731,N_729);
nand U858 (N_858,N_765,N_739);
or U859 (N_859,N_705,N_718);
or U860 (N_860,N_738,N_723);
and U861 (N_861,N_790,N_748);
nand U862 (N_862,N_796,N_721);
and U863 (N_863,N_781,N_761);
or U864 (N_864,N_762,N_758);
nor U865 (N_865,N_710,N_751);
nand U866 (N_866,N_786,N_741);
and U867 (N_867,N_707,N_757);
or U868 (N_868,N_713,N_777);
and U869 (N_869,N_768,N_747);
nand U870 (N_870,N_716,N_795);
nand U871 (N_871,N_751,N_747);
or U872 (N_872,N_716,N_727);
nor U873 (N_873,N_760,N_776);
nor U874 (N_874,N_746,N_755);
or U875 (N_875,N_786,N_747);
xnor U876 (N_876,N_710,N_790);
and U877 (N_877,N_771,N_789);
nand U878 (N_878,N_756,N_799);
nand U879 (N_879,N_793,N_745);
or U880 (N_880,N_776,N_791);
and U881 (N_881,N_701,N_798);
nand U882 (N_882,N_755,N_723);
or U883 (N_883,N_748,N_725);
nand U884 (N_884,N_743,N_706);
nand U885 (N_885,N_792,N_712);
or U886 (N_886,N_743,N_769);
or U887 (N_887,N_778,N_753);
nor U888 (N_888,N_703,N_723);
or U889 (N_889,N_787,N_742);
nor U890 (N_890,N_728,N_750);
or U891 (N_891,N_741,N_712);
or U892 (N_892,N_714,N_703);
and U893 (N_893,N_777,N_726);
or U894 (N_894,N_776,N_702);
or U895 (N_895,N_724,N_760);
nand U896 (N_896,N_723,N_785);
and U897 (N_897,N_754,N_776);
or U898 (N_898,N_720,N_745);
or U899 (N_899,N_736,N_770);
and U900 (N_900,N_864,N_815);
and U901 (N_901,N_802,N_884);
or U902 (N_902,N_896,N_804);
nand U903 (N_903,N_865,N_863);
and U904 (N_904,N_891,N_876);
and U905 (N_905,N_885,N_827);
nor U906 (N_906,N_856,N_899);
nand U907 (N_907,N_845,N_844);
nand U908 (N_908,N_855,N_897);
or U909 (N_909,N_886,N_812);
or U910 (N_910,N_837,N_866);
or U911 (N_911,N_862,N_859);
nand U912 (N_912,N_880,N_850);
and U913 (N_913,N_882,N_825);
or U914 (N_914,N_873,N_824);
or U915 (N_915,N_887,N_807);
nor U916 (N_916,N_822,N_817);
nor U917 (N_917,N_861,N_877);
or U918 (N_918,N_895,N_839);
and U919 (N_919,N_803,N_819);
or U920 (N_920,N_820,N_869);
nand U921 (N_921,N_872,N_801);
or U922 (N_922,N_893,N_806);
or U923 (N_923,N_874,N_835);
or U924 (N_924,N_846,N_854);
and U925 (N_925,N_883,N_871);
nor U926 (N_926,N_878,N_879);
or U927 (N_927,N_805,N_889);
or U928 (N_928,N_830,N_860);
nand U929 (N_929,N_832,N_800);
xnor U930 (N_930,N_823,N_842);
nand U931 (N_931,N_849,N_831);
or U932 (N_932,N_852,N_834);
and U933 (N_933,N_843,N_828);
or U934 (N_934,N_810,N_847);
or U935 (N_935,N_868,N_841);
and U936 (N_936,N_813,N_840);
or U937 (N_937,N_858,N_826);
or U938 (N_938,N_811,N_818);
nor U939 (N_939,N_836,N_821);
or U940 (N_940,N_851,N_870);
and U941 (N_941,N_814,N_892);
nand U942 (N_942,N_881,N_867);
and U943 (N_943,N_898,N_829);
nor U944 (N_944,N_853,N_888);
or U945 (N_945,N_816,N_838);
or U946 (N_946,N_848,N_894);
or U947 (N_947,N_833,N_890);
nor U948 (N_948,N_875,N_857);
nand U949 (N_949,N_808,N_809);
nand U950 (N_950,N_893,N_872);
or U951 (N_951,N_874,N_868);
or U952 (N_952,N_864,N_898);
nand U953 (N_953,N_850,N_846);
or U954 (N_954,N_880,N_831);
or U955 (N_955,N_829,N_809);
and U956 (N_956,N_813,N_819);
or U957 (N_957,N_804,N_803);
and U958 (N_958,N_889,N_809);
nand U959 (N_959,N_865,N_833);
and U960 (N_960,N_858,N_811);
nor U961 (N_961,N_836,N_833);
nor U962 (N_962,N_843,N_861);
nand U963 (N_963,N_835,N_832);
nand U964 (N_964,N_889,N_871);
nand U965 (N_965,N_824,N_802);
or U966 (N_966,N_806,N_811);
and U967 (N_967,N_886,N_871);
and U968 (N_968,N_889,N_895);
nand U969 (N_969,N_801,N_899);
nand U970 (N_970,N_871,N_816);
nor U971 (N_971,N_855,N_800);
and U972 (N_972,N_818,N_880);
and U973 (N_973,N_849,N_875);
and U974 (N_974,N_846,N_887);
nor U975 (N_975,N_873,N_898);
nor U976 (N_976,N_895,N_888);
and U977 (N_977,N_849,N_838);
nor U978 (N_978,N_868,N_806);
nand U979 (N_979,N_848,N_811);
nand U980 (N_980,N_848,N_818);
and U981 (N_981,N_865,N_899);
and U982 (N_982,N_863,N_810);
or U983 (N_983,N_850,N_833);
nor U984 (N_984,N_809,N_890);
and U985 (N_985,N_809,N_896);
and U986 (N_986,N_825,N_807);
nand U987 (N_987,N_842,N_839);
and U988 (N_988,N_804,N_816);
or U989 (N_989,N_820,N_895);
and U990 (N_990,N_879,N_806);
nor U991 (N_991,N_883,N_898);
nand U992 (N_992,N_879,N_851);
or U993 (N_993,N_816,N_805);
nor U994 (N_994,N_855,N_867);
nand U995 (N_995,N_881,N_876);
xnor U996 (N_996,N_894,N_841);
nand U997 (N_997,N_828,N_855);
nand U998 (N_998,N_810,N_899);
nor U999 (N_999,N_852,N_889);
and U1000 (N_1000,N_902,N_907);
or U1001 (N_1001,N_933,N_909);
or U1002 (N_1002,N_991,N_924);
or U1003 (N_1003,N_986,N_937);
or U1004 (N_1004,N_927,N_957);
or U1005 (N_1005,N_940,N_956);
and U1006 (N_1006,N_970,N_915);
or U1007 (N_1007,N_900,N_979);
and U1008 (N_1008,N_994,N_992);
or U1009 (N_1009,N_976,N_982);
or U1010 (N_1010,N_950,N_995);
and U1011 (N_1011,N_938,N_960);
and U1012 (N_1012,N_987,N_906);
or U1013 (N_1013,N_905,N_965);
nor U1014 (N_1014,N_972,N_908);
nor U1015 (N_1015,N_952,N_920);
nand U1016 (N_1016,N_939,N_984);
and U1017 (N_1017,N_934,N_928);
or U1018 (N_1018,N_935,N_945);
nor U1019 (N_1019,N_917,N_904);
nor U1020 (N_1020,N_923,N_962);
nor U1021 (N_1021,N_903,N_998);
nand U1022 (N_1022,N_975,N_990);
nor U1023 (N_1023,N_914,N_931);
nor U1024 (N_1024,N_974,N_969);
or U1025 (N_1025,N_989,N_951);
nor U1026 (N_1026,N_997,N_948);
or U1027 (N_1027,N_921,N_958);
or U1028 (N_1028,N_966,N_959);
or U1029 (N_1029,N_913,N_942);
nor U1030 (N_1030,N_941,N_947);
and U1031 (N_1031,N_973,N_911);
or U1032 (N_1032,N_955,N_949);
or U1033 (N_1033,N_912,N_930);
nor U1034 (N_1034,N_918,N_932);
nand U1035 (N_1035,N_944,N_985);
nor U1036 (N_1036,N_981,N_916);
nor U1037 (N_1037,N_925,N_954);
nor U1038 (N_1038,N_971,N_983);
nor U1039 (N_1039,N_929,N_996);
nor U1040 (N_1040,N_964,N_910);
or U1041 (N_1041,N_993,N_968);
or U1042 (N_1042,N_901,N_953);
and U1043 (N_1043,N_978,N_946);
nand U1044 (N_1044,N_926,N_943);
or U1045 (N_1045,N_988,N_967);
or U1046 (N_1046,N_977,N_961);
nand U1047 (N_1047,N_922,N_936);
nand U1048 (N_1048,N_919,N_963);
and U1049 (N_1049,N_999,N_980);
and U1050 (N_1050,N_966,N_937);
nand U1051 (N_1051,N_943,N_976);
nor U1052 (N_1052,N_920,N_900);
and U1053 (N_1053,N_902,N_911);
and U1054 (N_1054,N_925,N_928);
nor U1055 (N_1055,N_982,N_934);
nor U1056 (N_1056,N_931,N_921);
and U1057 (N_1057,N_963,N_948);
and U1058 (N_1058,N_983,N_905);
or U1059 (N_1059,N_942,N_947);
nand U1060 (N_1060,N_962,N_924);
and U1061 (N_1061,N_945,N_953);
nand U1062 (N_1062,N_933,N_940);
nand U1063 (N_1063,N_979,N_994);
and U1064 (N_1064,N_988,N_987);
nand U1065 (N_1065,N_952,N_954);
and U1066 (N_1066,N_904,N_928);
nand U1067 (N_1067,N_996,N_957);
or U1068 (N_1068,N_980,N_998);
nor U1069 (N_1069,N_919,N_904);
and U1070 (N_1070,N_985,N_912);
and U1071 (N_1071,N_960,N_904);
or U1072 (N_1072,N_991,N_925);
nor U1073 (N_1073,N_947,N_940);
nor U1074 (N_1074,N_934,N_909);
and U1075 (N_1075,N_923,N_908);
or U1076 (N_1076,N_952,N_959);
and U1077 (N_1077,N_944,N_922);
nor U1078 (N_1078,N_963,N_927);
or U1079 (N_1079,N_980,N_918);
nand U1080 (N_1080,N_951,N_965);
or U1081 (N_1081,N_926,N_938);
nand U1082 (N_1082,N_958,N_949);
or U1083 (N_1083,N_945,N_970);
or U1084 (N_1084,N_979,N_949);
nand U1085 (N_1085,N_902,N_975);
nand U1086 (N_1086,N_914,N_938);
or U1087 (N_1087,N_952,N_974);
xor U1088 (N_1088,N_963,N_921);
nor U1089 (N_1089,N_905,N_923);
or U1090 (N_1090,N_907,N_988);
or U1091 (N_1091,N_925,N_972);
nand U1092 (N_1092,N_978,N_986);
and U1093 (N_1093,N_954,N_902);
nor U1094 (N_1094,N_906,N_972);
nor U1095 (N_1095,N_999,N_944);
and U1096 (N_1096,N_998,N_982);
nor U1097 (N_1097,N_954,N_943);
or U1098 (N_1098,N_953,N_995);
or U1099 (N_1099,N_936,N_988);
or U1100 (N_1100,N_1011,N_1010);
and U1101 (N_1101,N_1069,N_1065);
nor U1102 (N_1102,N_1080,N_1027);
nor U1103 (N_1103,N_1034,N_1070);
nor U1104 (N_1104,N_1087,N_1074);
xnor U1105 (N_1105,N_1063,N_1092);
or U1106 (N_1106,N_1035,N_1022);
nor U1107 (N_1107,N_1006,N_1021);
nor U1108 (N_1108,N_1054,N_1061);
and U1109 (N_1109,N_1019,N_1044);
nor U1110 (N_1110,N_1057,N_1008);
nand U1111 (N_1111,N_1051,N_1085);
nand U1112 (N_1112,N_1047,N_1068);
or U1113 (N_1113,N_1023,N_1050);
or U1114 (N_1114,N_1058,N_1028);
nand U1115 (N_1115,N_1096,N_1090);
and U1116 (N_1116,N_1098,N_1072);
and U1117 (N_1117,N_1009,N_1083);
and U1118 (N_1118,N_1071,N_1039);
or U1119 (N_1119,N_1030,N_1045);
and U1120 (N_1120,N_1055,N_1097);
nor U1121 (N_1121,N_1040,N_1077);
nand U1122 (N_1122,N_1079,N_1020);
nor U1123 (N_1123,N_1015,N_1060);
or U1124 (N_1124,N_1095,N_1052);
and U1125 (N_1125,N_1046,N_1002);
nand U1126 (N_1126,N_1024,N_1073);
or U1127 (N_1127,N_1048,N_1016);
or U1128 (N_1128,N_1056,N_1053);
and U1129 (N_1129,N_1025,N_1033);
nor U1130 (N_1130,N_1000,N_1005);
nor U1131 (N_1131,N_1031,N_1084);
nor U1132 (N_1132,N_1099,N_1088);
nand U1133 (N_1133,N_1094,N_1091);
and U1134 (N_1134,N_1013,N_1036);
and U1135 (N_1135,N_1067,N_1012);
and U1136 (N_1136,N_1059,N_1081);
or U1137 (N_1137,N_1066,N_1093);
nand U1138 (N_1138,N_1037,N_1018);
or U1139 (N_1139,N_1078,N_1001);
or U1140 (N_1140,N_1043,N_1026);
nor U1141 (N_1141,N_1004,N_1029);
nor U1142 (N_1142,N_1032,N_1014);
nand U1143 (N_1143,N_1041,N_1089);
and U1144 (N_1144,N_1049,N_1076);
nor U1145 (N_1145,N_1062,N_1038);
and U1146 (N_1146,N_1042,N_1086);
nor U1147 (N_1147,N_1003,N_1075);
and U1148 (N_1148,N_1007,N_1082);
or U1149 (N_1149,N_1017,N_1064);
nor U1150 (N_1150,N_1062,N_1079);
nor U1151 (N_1151,N_1034,N_1079);
nor U1152 (N_1152,N_1059,N_1022);
or U1153 (N_1153,N_1012,N_1048);
or U1154 (N_1154,N_1075,N_1090);
and U1155 (N_1155,N_1009,N_1058);
nor U1156 (N_1156,N_1027,N_1077);
nand U1157 (N_1157,N_1098,N_1000);
or U1158 (N_1158,N_1039,N_1035);
or U1159 (N_1159,N_1074,N_1065);
nor U1160 (N_1160,N_1080,N_1075);
nand U1161 (N_1161,N_1099,N_1031);
nor U1162 (N_1162,N_1047,N_1017);
nand U1163 (N_1163,N_1066,N_1004);
nor U1164 (N_1164,N_1087,N_1004);
and U1165 (N_1165,N_1042,N_1026);
nand U1166 (N_1166,N_1003,N_1091);
xnor U1167 (N_1167,N_1047,N_1009);
xor U1168 (N_1168,N_1035,N_1068);
nor U1169 (N_1169,N_1092,N_1040);
nand U1170 (N_1170,N_1023,N_1020);
or U1171 (N_1171,N_1021,N_1061);
nor U1172 (N_1172,N_1075,N_1060);
and U1173 (N_1173,N_1056,N_1011);
nor U1174 (N_1174,N_1094,N_1028);
nor U1175 (N_1175,N_1064,N_1031);
nor U1176 (N_1176,N_1005,N_1097);
nand U1177 (N_1177,N_1098,N_1071);
nand U1178 (N_1178,N_1069,N_1077);
nand U1179 (N_1179,N_1049,N_1097);
nor U1180 (N_1180,N_1039,N_1094);
nor U1181 (N_1181,N_1033,N_1024);
nor U1182 (N_1182,N_1049,N_1060);
or U1183 (N_1183,N_1001,N_1055);
nand U1184 (N_1184,N_1037,N_1071);
and U1185 (N_1185,N_1091,N_1048);
nand U1186 (N_1186,N_1007,N_1092);
nor U1187 (N_1187,N_1045,N_1027);
nor U1188 (N_1188,N_1046,N_1089);
nor U1189 (N_1189,N_1033,N_1081);
nand U1190 (N_1190,N_1059,N_1069);
or U1191 (N_1191,N_1055,N_1096);
xnor U1192 (N_1192,N_1034,N_1016);
nand U1193 (N_1193,N_1043,N_1030);
xor U1194 (N_1194,N_1046,N_1076);
and U1195 (N_1195,N_1023,N_1088);
and U1196 (N_1196,N_1029,N_1098);
nand U1197 (N_1197,N_1045,N_1086);
or U1198 (N_1198,N_1064,N_1048);
nand U1199 (N_1199,N_1006,N_1044);
and U1200 (N_1200,N_1158,N_1154);
and U1201 (N_1201,N_1117,N_1100);
or U1202 (N_1202,N_1155,N_1127);
nor U1203 (N_1203,N_1136,N_1142);
or U1204 (N_1204,N_1163,N_1134);
and U1205 (N_1205,N_1166,N_1102);
and U1206 (N_1206,N_1173,N_1153);
nand U1207 (N_1207,N_1108,N_1109);
and U1208 (N_1208,N_1171,N_1185);
nand U1209 (N_1209,N_1144,N_1156);
and U1210 (N_1210,N_1149,N_1174);
or U1211 (N_1211,N_1133,N_1119);
or U1212 (N_1212,N_1105,N_1141);
nand U1213 (N_1213,N_1101,N_1161);
or U1214 (N_1214,N_1182,N_1172);
and U1215 (N_1215,N_1115,N_1194);
or U1216 (N_1216,N_1186,N_1184);
nand U1217 (N_1217,N_1125,N_1188);
and U1218 (N_1218,N_1162,N_1151);
nor U1219 (N_1219,N_1130,N_1169);
or U1220 (N_1220,N_1140,N_1179);
and U1221 (N_1221,N_1116,N_1180);
nor U1222 (N_1222,N_1160,N_1196);
and U1223 (N_1223,N_1177,N_1112);
nor U1224 (N_1224,N_1139,N_1195);
and U1225 (N_1225,N_1168,N_1110);
nor U1226 (N_1226,N_1175,N_1170);
xor U1227 (N_1227,N_1164,N_1145);
and U1228 (N_1228,N_1126,N_1189);
nand U1229 (N_1229,N_1143,N_1192);
and U1230 (N_1230,N_1114,N_1198);
and U1231 (N_1231,N_1178,N_1121);
and U1232 (N_1232,N_1118,N_1111);
nand U1233 (N_1233,N_1106,N_1138);
or U1234 (N_1234,N_1124,N_1167);
and U1235 (N_1235,N_1122,N_1128);
nor U1236 (N_1236,N_1135,N_1152);
nand U1237 (N_1237,N_1190,N_1157);
and U1238 (N_1238,N_1131,N_1103);
nor U1239 (N_1239,N_1146,N_1199);
and U1240 (N_1240,N_1129,N_1123);
nor U1241 (N_1241,N_1107,N_1183);
and U1242 (N_1242,N_1148,N_1193);
or U1243 (N_1243,N_1181,N_1176);
or U1244 (N_1244,N_1187,N_1120);
and U1245 (N_1245,N_1104,N_1113);
or U1246 (N_1246,N_1165,N_1159);
and U1247 (N_1247,N_1147,N_1150);
or U1248 (N_1248,N_1132,N_1191);
and U1249 (N_1249,N_1197,N_1137);
or U1250 (N_1250,N_1137,N_1133);
nor U1251 (N_1251,N_1113,N_1194);
or U1252 (N_1252,N_1138,N_1128);
or U1253 (N_1253,N_1136,N_1107);
and U1254 (N_1254,N_1138,N_1192);
xnor U1255 (N_1255,N_1159,N_1151);
or U1256 (N_1256,N_1158,N_1189);
nand U1257 (N_1257,N_1114,N_1167);
and U1258 (N_1258,N_1142,N_1128);
nand U1259 (N_1259,N_1194,N_1193);
or U1260 (N_1260,N_1181,N_1150);
nor U1261 (N_1261,N_1156,N_1195);
nand U1262 (N_1262,N_1169,N_1105);
nand U1263 (N_1263,N_1103,N_1106);
and U1264 (N_1264,N_1187,N_1178);
nor U1265 (N_1265,N_1145,N_1109);
nor U1266 (N_1266,N_1139,N_1174);
nor U1267 (N_1267,N_1166,N_1172);
and U1268 (N_1268,N_1107,N_1167);
and U1269 (N_1269,N_1143,N_1159);
or U1270 (N_1270,N_1123,N_1150);
and U1271 (N_1271,N_1194,N_1114);
or U1272 (N_1272,N_1196,N_1133);
nand U1273 (N_1273,N_1178,N_1125);
nor U1274 (N_1274,N_1134,N_1149);
nand U1275 (N_1275,N_1165,N_1174);
nor U1276 (N_1276,N_1141,N_1144);
or U1277 (N_1277,N_1100,N_1104);
nand U1278 (N_1278,N_1140,N_1158);
nor U1279 (N_1279,N_1159,N_1174);
nand U1280 (N_1280,N_1187,N_1175);
nand U1281 (N_1281,N_1164,N_1115);
or U1282 (N_1282,N_1131,N_1112);
nand U1283 (N_1283,N_1137,N_1126);
and U1284 (N_1284,N_1142,N_1137);
nand U1285 (N_1285,N_1141,N_1112);
and U1286 (N_1286,N_1111,N_1180);
and U1287 (N_1287,N_1184,N_1138);
or U1288 (N_1288,N_1106,N_1198);
nand U1289 (N_1289,N_1183,N_1157);
nor U1290 (N_1290,N_1126,N_1144);
or U1291 (N_1291,N_1193,N_1178);
nand U1292 (N_1292,N_1103,N_1198);
and U1293 (N_1293,N_1144,N_1114);
or U1294 (N_1294,N_1101,N_1107);
and U1295 (N_1295,N_1139,N_1150);
or U1296 (N_1296,N_1183,N_1116);
nand U1297 (N_1297,N_1137,N_1145);
and U1298 (N_1298,N_1126,N_1135);
nand U1299 (N_1299,N_1113,N_1188);
nor U1300 (N_1300,N_1290,N_1225);
or U1301 (N_1301,N_1200,N_1236);
and U1302 (N_1302,N_1251,N_1237);
nor U1303 (N_1303,N_1280,N_1209);
nor U1304 (N_1304,N_1202,N_1205);
nor U1305 (N_1305,N_1277,N_1232);
nor U1306 (N_1306,N_1293,N_1210);
or U1307 (N_1307,N_1204,N_1283);
and U1308 (N_1308,N_1261,N_1250);
and U1309 (N_1309,N_1230,N_1292);
nand U1310 (N_1310,N_1273,N_1276);
nor U1311 (N_1311,N_1270,N_1275);
or U1312 (N_1312,N_1278,N_1258);
or U1313 (N_1313,N_1221,N_1226);
or U1314 (N_1314,N_1219,N_1244);
and U1315 (N_1315,N_1255,N_1285);
or U1316 (N_1316,N_1214,N_1242);
and U1317 (N_1317,N_1218,N_1207);
xor U1318 (N_1318,N_1266,N_1298);
nor U1319 (N_1319,N_1297,N_1281);
or U1320 (N_1320,N_1247,N_1238);
nand U1321 (N_1321,N_1227,N_1216);
or U1322 (N_1322,N_1256,N_1233);
or U1323 (N_1323,N_1265,N_1267);
or U1324 (N_1324,N_1253,N_1262);
or U1325 (N_1325,N_1222,N_1268);
nand U1326 (N_1326,N_1257,N_1284);
or U1327 (N_1327,N_1211,N_1246);
nor U1328 (N_1328,N_1282,N_1288);
nand U1329 (N_1329,N_1274,N_1264);
or U1330 (N_1330,N_1259,N_1206);
nand U1331 (N_1331,N_1239,N_1252);
and U1332 (N_1332,N_1243,N_1271);
and U1333 (N_1333,N_1208,N_1229);
or U1334 (N_1334,N_1215,N_1217);
nand U1335 (N_1335,N_1201,N_1279);
and U1336 (N_1336,N_1287,N_1223);
or U1337 (N_1337,N_1289,N_1294);
xnor U1338 (N_1338,N_1254,N_1241);
nor U1339 (N_1339,N_1245,N_1235);
nand U1340 (N_1340,N_1269,N_1234);
nor U1341 (N_1341,N_1213,N_1260);
and U1342 (N_1342,N_1296,N_1240);
or U1343 (N_1343,N_1224,N_1220);
nand U1344 (N_1344,N_1263,N_1228);
nor U1345 (N_1345,N_1248,N_1299);
or U1346 (N_1346,N_1231,N_1249);
or U1347 (N_1347,N_1286,N_1203);
nor U1348 (N_1348,N_1291,N_1295);
nand U1349 (N_1349,N_1212,N_1272);
nor U1350 (N_1350,N_1278,N_1214);
nor U1351 (N_1351,N_1255,N_1243);
nor U1352 (N_1352,N_1219,N_1238);
or U1353 (N_1353,N_1204,N_1223);
nand U1354 (N_1354,N_1296,N_1260);
nand U1355 (N_1355,N_1223,N_1298);
nor U1356 (N_1356,N_1255,N_1250);
nand U1357 (N_1357,N_1255,N_1284);
or U1358 (N_1358,N_1222,N_1283);
and U1359 (N_1359,N_1228,N_1246);
nor U1360 (N_1360,N_1292,N_1261);
nor U1361 (N_1361,N_1254,N_1201);
nor U1362 (N_1362,N_1268,N_1249);
nand U1363 (N_1363,N_1214,N_1282);
and U1364 (N_1364,N_1230,N_1218);
xor U1365 (N_1365,N_1278,N_1281);
and U1366 (N_1366,N_1245,N_1208);
or U1367 (N_1367,N_1252,N_1299);
nand U1368 (N_1368,N_1215,N_1229);
or U1369 (N_1369,N_1233,N_1257);
nor U1370 (N_1370,N_1215,N_1228);
or U1371 (N_1371,N_1268,N_1245);
nor U1372 (N_1372,N_1216,N_1283);
nor U1373 (N_1373,N_1204,N_1208);
nand U1374 (N_1374,N_1269,N_1243);
nor U1375 (N_1375,N_1233,N_1260);
nor U1376 (N_1376,N_1211,N_1221);
nor U1377 (N_1377,N_1204,N_1269);
nor U1378 (N_1378,N_1278,N_1260);
or U1379 (N_1379,N_1229,N_1241);
and U1380 (N_1380,N_1285,N_1204);
or U1381 (N_1381,N_1258,N_1234);
nor U1382 (N_1382,N_1283,N_1229);
nand U1383 (N_1383,N_1221,N_1202);
nand U1384 (N_1384,N_1247,N_1281);
or U1385 (N_1385,N_1285,N_1296);
nand U1386 (N_1386,N_1261,N_1283);
or U1387 (N_1387,N_1268,N_1267);
and U1388 (N_1388,N_1210,N_1264);
nand U1389 (N_1389,N_1220,N_1247);
or U1390 (N_1390,N_1223,N_1254);
nand U1391 (N_1391,N_1230,N_1280);
nand U1392 (N_1392,N_1226,N_1214);
or U1393 (N_1393,N_1219,N_1292);
and U1394 (N_1394,N_1245,N_1279);
nor U1395 (N_1395,N_1225,N_1283);
and U1396 (N_1396,N_1266,N_1237);
nand U1397 (N_1397,N_1246,N_1240);
nor U1398 (N_1398,N_1204,N_1256);
nor U1399 (N_1399,N_1232,N_1252);
and U1400 (N_1400,N_1377,N_1354);
nor U1401 (N_1401,N_1326,N_1349);
nand U1402 (N_1402,N_1308,N_1321);
nand U1403 (N_1403,N_1388,N_1368);
or U1404 (N_1404,N_1323,N_1322);
nand U1405 (N_1405,N_1391,N_1339);
or U1406 (N_1406,N_1305,N_1307);
and U1407 (N_1407,N_1387,N_1373);
and U1408 (N_1408,N_1312,N_1378);
nor U1409 (N_1409,N_1301,N_1356);
nand U1410 (N_1410,N_1313,N_1398);
nor U1411 (N_1411,N_1332,N_1304);
or U1412 (N_1412,N_1362,N_1360);
nand U1413 (N_1413,N_1314,N_1336);
and U1414 (N_1414,N_1340,N_1309);
or U1415 (N_1415,N_1343,N_1371);
nand U1416 (N_1416,N_1350,N_1366);
or U1417 (N_1417,N_1382,N_1365);
nor U1418 (N_1418,N_1345,N_1393);
nand U1419 (N_1419,N_1300,N_1310);
nor U1420 (N_1420,N_1324,N_1311);
and U1421 (N_1421,N_1338,N_1306);
and U1422 (N_1422,N_1347,N_1399);
or U1423 (N_1423,N_1315,N_1341);
nor U1424 (N_1424,N_1372,N_1329);
nor U1425 (N_1425,N_1337,N_1318);
nor U1426 (N_1426,N_1374,N_1328);
or U1427 (N_1427,N_1359,N_1394);
or U1428 (N_1428,N_1361,N_1316);
or U1429 (N_1429,N_1381,N_1385);
nand U1430 (N_1430,N_1327,N_1370);
and U1431 (N_1431,N_1302,N_1335);
and U1432 (N_1432,N_1351,N_1389);
or U1433 (N_1433,N_1379,N_1348);
nand U1434 (N_1434,N_1363,N_1396);
or U1435 (N_1435,N_1320,N_1319);
nor U1436 (N_1436,N_1303,N_1353);
or U1437 (N_1437,N_1397,N_1380);
nor U1438 (N_1438,N_1357,N_1358);
nor U1439 (N_1439,N_1383,N_1331);
nand U1440 (N_1440,N_1375,N_1395);
or U1441 (N_1441,N_1392,N_1342);
or U1442 (N_1442,N_1352,N_1367);
or U1443 (N_1443,N_1325,N_1390);
xnor U1444 (N_1444,N_1369,N_1355);
nand U1445 (N_1445,N_1384,N_1333);
and U1446 (N_1446,N_1330,N_1344);
and U1447 (N_1447,N_1334,N_1376);
or U1448 (N_1448,N_1386,N_1317);
or U1449 (N_1449,N_1346,N_1364);
xor U1450 (N_1450,N_1331,N_1325);
or U1451 (N_1451,N_1393,N_1315);
and U1452 (N_1452,N_1361,N_1363);
or U1453 (N_1453,N_1304,N_1303);
nor U1454 (N_1454,N_1339,N_1309);
and U1455 (N_1455,N_1361,N_1365);
or U1456 (N_1456,N_1390,N_1349);
and U1457 (N_1457,N_1375,N_1391);
nand U1458 (N_1458,N_1376,N_1352);
xor U1459 (N_1459,N_1353,N_1398);
nand U1460 (N_1460,N_1354,N_1345);
nand U1461 (N_1461,N_1352,N_1387);
nor U1462 (N_1462,N_1376,N_1375);
nor U1463 (N_1463,N_1397,N_1324);
nor U1464 (N_1464,N_1320,N_1374);
nand U1465 (N_1465,N_1392,N_1312);
nand U1466 (N_1466,N_1343,N_1351);
and U1467 (N_1467,N_1302,N_1324);
and U1468 (N_1468,N_1330,N_1378);
nand U1469 (N_1469,N_1387,N_1315);
or U1470 (N_1470,N_1372,N_1321);
nand U1471 (N_1471,N_1323,N_1315);
nor U1472 (N_1472,N_1384,N_1363);
nand U1473 (N_1473,N_1350,N_1349);
and U1474 (N_1474,N_1395,N_1316);
and U1475 (N_1475,N_1329,N_1380);
nor U1476 (N_1476,N_1353,N_1332);
nand U1477 (N_1477,N_1386,N_1349);
or U1478 (N_1478,N_1339,N_1351);
and U1479 (N_1479,N_1379,N_1315);
nand U1480 (N_1480,N_1328,N_1329);
or U1481 (N_1481,N_1399,N_1336);
and U1482 (N_1482,N_1355,N_1352);
or U1483 (N_1483,N_1369,N_1341);
nand U1484 (N_1484,N_1327,N_1313);
nand U1485 (N_1485,N_1335,N_1325);
nand U1486 (N_1486,N_1398,N_1357);
or U1487 (N_1487,N_1340,N_1372);
nor U1488 (N_1488,N_1309,N_1335);
or U1489 (N_1489,N_1312,N_1348);
or U1490 (N_1490,N_1381,N_1366);
and U1491 (N_1491,N_1318,N_1324);
nand U1492 (N_1492,N_1362,N_1311);
nor U1493 (N_1493,N_1373,N_1318);
nand U1494 (N_1494,N_1370,N_1311);
and U1495 (N_1495,N_1354,N_1384);
or U1496 (N_1496,N_1301,N_1381);
nand U1497 (N_1497,N_1342,N_1303);
nor U1498 (N_1498,N_1311,N_1394);
nor U1499 (N_1499,N_1349,N_1344);
or U1500 (N_1500,N_1440,N_1468);
and U1501 (N_1501,N_1403,N_1431);
nand U1502 (N_1502,N_1402,N_1474);
and U1503 (N_1503,N_1497,N_1444);
or U1504 (N_1504,N_1467,N_1439);
or U1505 (N_1505,N_1461,N_1421);
nand U1506 (N_1506,N_1416,N_1406);
nor U1507 (N_1507,N_1481,N_1405);
or U1508 (N_1508,N_1414,N_1466);
or U1509 (N_1509,N_1407,N_1453);
xor U1510 (N_1510,N_1408,N_1464);
and U1511 (N_1511,N_1483,N_1463);
and U1512 (N_1512,N_1425,N_1470);
and U1513 (N_1513,N_1426,N_1465);
or U1514 (N_1514,N_1434,N_1415);
and U1515 (N_1515,N_1418,N_1457);
nand U1516 (N_1516,N_1489,N_1485);
nor U1517 (N_1517,N_1496,N_1451);
nand U1518 (N_1518,N_1411,N_1455);
nand U1519 (N_1519,N_1495,N_1480);
xnor U1520 (N_1520,N_1456,N_1429);
and U1521 (N_1521,N_1460,N_1428);
and U1522 (N_1522,N_1424,N_1417);
nand U1523 (N_1523,N_1433,N_1454);
nor U1524 (N_1524,N_1449,N_1458);
nor U1525 (N_1525,N_1488,N_1410);
and U1526 (N_1526,N_1423,N_1413);
nand U1527 (N_1527,N_1445,N_1427);
nand U1528 (N_1528,N_1404,N_1492);
nor U1529 (N_1529,N_1437,N_1435);
nor U1530 (N_1530,N_1475,N_1487);
nand U1531 (N_1531,N_1401,N_1438);
or U1532 (N_1532,N_1452,N_1420);
and U1533 (N_1533,N_1471,N_1441);
nor U1534 (N_1534,N_1478,N_1409);
nor U1535 (N_1535,N_1446,N_1422);
nand U1536 (N_1536,N_1493,N_1447);
nand U1537 (N_1537,N_1476,N_1450);
nand U1538 (N_1538,N_1400,N_1430);
and U1539 (N_1539,N_1419,N_1479);
nor U1540 (N_1540,N_1486,N_1490);
or U1541 (N_1541,N_1448,N_1462);
and U1542 (N_1542,N_1494,N_1459);
nor U1543 (N_1543,N_1491,N_1473);
nor U1544 (N_1544,N_1484,N_1472);
and U1545 (N_1545,N_1498,N_1443);
and U1546 (N_1546,N_1477,N_1436);
nor U1547 (N_1547,N_1442,N_1482);
nor U1548 (N_1548,N_1469,N_1499);
nand U1549 (N_1549,N_1412,N_1432);
and U1550 (N_1550,N_1498,N_1450);
and U1551 (N_1551,N_1460,N_1430);
nand U1552 (N_1552,N_1468,N_1402);
or U1553 (N_1553,N_1473,N_1435);
and U1554 (N_1554,N_1443,N_1458);
and U1555 (N_1555,N_1461,N_1493);
nand U1556 (N_1556,N_1467,N_1423);
nor U1557 (N_1557,N_1416,N_1423);
nand U1558 (N_1558,N_1496,N_1403);
and U1559 (N_1559,N_1425,N_1479);
or U1560 (N_1560,N_1434,N_1410);
or U1561 (N_1561,N_1415,N_1402);
nor U1562 (N_1562,N_1419,N_1433);
and U1563 (N_1563,N_1482,N_1493);
nand U1564 (N_1564,N_1401,N_1453);
or U1565 (N_1565,N_1450,N_1491);
and U1566 (N_1566,N_1420,N_1403);
or U1567 (N_1567,N_1479,N_1455);
nand U1568 (N_1568,N_1425,N_1492);
nor U1569 (N_1569,N_1458,N_1488);
and U1570 (N_1570,N_1430,N_1408);
nor U1571 (N_1571,N_1444,N_1481);
nor U1572 (N_1572,N_1478,N_1447);
nor U1573 (N_1573,N_1494,N_1425);
nor U1574 (N_1574,N_1434,N_1411);
or U1575 (N_1575,N_1458,N_1401);
nand U1576 (N_1576,N_1471,N_1409);
and U1577 (N_1577,N_1452,N_1403);
nor U1578 (N_1578,N_1446,N_1443);
nor U1579 (N_1579,N_1420,N_1467);
or U1580 (N_1580,N_1444,N_1403);
nor U1581 (N_1581,N_1451,N_1460);
or U1582 (N_1582,N_1450,N_1475);
or U1583 (N_1583,N_1496,N_1407);
or U1584 (N_1584,N_1416,N_1463);
or U1585 (N_1585,N_1412,N_1489);
nand U1586 (N_1586,N_1448,N_1452);
nand U1587 (N_1587,N_1455,N_1413);
and U1588 (N_1588,N_1471,N_1415);
nand U1589 (N_1589,N_1484,N_1432);
or U1590 (N_1590,N_1439,N_1457);
nand U1591 (N_1591,N_1406,N_1420);
nand U1592 (N_1592,N_1443,N_1495);
nor U1593 (N_1593,N_1446,N_1441);
nand U1594 (N_1594,N_1402,N_1457);
nor U1595 (N_1595,N_1409,N_1474);
and U1596 (N_1596,N_1439,N_1483);
and U1597 (N_1597,N_1457,N_1446);
nand U1598 (N_1598,N_1404,N_1401);
or U1599 (N_1599,N_1410,N_1469);
nand U1600 (N_1600,N_1532,N_1561);
or U1601 (N_1601,N_1544,N_1579);
and U1602 (N_1602,N_1599,N_1553);
nor U1603 (N_1603,N_1535,N_1550);
or U1604 (N_1604,N_1570,N_1513);
or U1605 (N_1605,N_1564,N_1514);
nand U1606 (N_1606,N_1523,N_1530);
nor U1607 (N_1607,N_1571,N_1567);
nor U1608 (N_1608,N_1554,N_1538);
or U1609 (N_1609,N_1506,N_1569);
nand U1610 (N_1610,N_1528,N_1578);
nand U1611 (N_1611,N_1568,N_1508);
nor U1612 (N_1612,N_1542,N_1598);
nor U1613 (N_1613,N_1541,N_1588);
nor U1614 (N_1614,N_1500,N_1504);
and U1615 (N_1615,N_1520,N_1595);
nor U1616 (N_1616,N_1531,N_1587);
nor U1617 (N_1617,N_1533,N_1549);
nand U1618 (N_1618,N_1505,N_1556);
nand U1619 (N_1619,N_1518,N_1548);
nor U1620 (N_1620,N_1512,N_1558);
and U1621 (N_1621,N_1591,N_1502);
or U1622 (N_1622,N_1540,N_1522);
nand U1623 (N_1623,N_1584,N_1575);
or U1624 (N_1624,N_1524,N_1526);
or U1625 (N_1625,N_1593,N_1586);
nand U1626 (N_1626,N_1583,N_1589);
nand U1627 (N_1627,N_1510,N_1527);
nor U1628 (N_1628,N_1534,N_1557);
and U1629 (N_1629,N_1515,N_1577);
nand U1630 (N_1630,N_1501,N_1511);
nor U1631 (N_1631,N_1594,N_1573);
or U1632 (N_1632,N_1536,N_1572);
nor U1633 (N_1633,N_1529,N_1507);
nor U1634 (N_1634,N_1516,N_1563);
nor U1635 (N_1635,N_1547,N_1509);
and U1636 (N_1636,N_1585,N_1517);
nor U1637 (N_1637,N_1580,N_1581);
or U1638 (N_1638,N_1560,N_1546);
and U1639 (N_1639,N_1582,N_1539);
and U1640 (N_1640,N_1555,N_1525);
or U1641 (N_1641,N_1543,N_1596);
nor U1642 (N_1642,N_1576,N_1537);
and U1643 (N_1643,N_1551,N_1566);
or U1644 (N_1644,N_1521,N_1592);
nand U1645 (N_1645,N_1552,N_1565);
nor U1646 (N_1646,N_1597,N_1559);
or U1647 (N_1647,N_1519,N_1545);
or U1648 (N_1648,N_1590,N_1503);
or U1649 (N_1649,N_1574,N_1562);
and U1650 (N_1650,N_1566,N_1540);
nand U1651 (N_1651,N_1515,N_1576);
nor U1652 (N_1652,N_1582,N_1505);
or U1653 (N_1653,N_1527,N_1591);
and U1654 (N_1654,N_1542,N_1509);
and U1655 (N_1655,N_1588,N_1594);
or U1656 (N_1656,N_1578,N_1576);
nand U1657 (N_1657,N_1571,N_1505);
or U1658 (N_1658,N_1507,N_1510);
and U1659 (N_1659,N_1508,N_1517);
or U1660 (N_1660,N_1536,N_1511);
nor U1661 (N_1661,N_1520,N_1509);
nor U1662 (N_1662,N_1545,N_1517);
nor U1663 (N_1663,N_1578,N_1596);
nand U1664 (N_1664,N_1504,N_1520);
nor U1665 (N_1665,N_1579,N_1543);
or U1666 (N_1666,N_1515,N_1543);
nor U1667 (N_1667,N_1591,N_1522);
or U1668 (N_1668,N_1582,N_1590);
or U1669 (N_1669,N_1512,N_1503);
or U1670 (N_1670,N_1512,N_1505);
nand U1671 (N_1671,N_1579,N_1511);
or U1672 (N_1672,N_1565,N_1550);
nor U1673 (N_1673,N_1591,N_1559);
or U1674 (N_1674,N_1587,N_1539);
nor U1675 (N_1675,N_1556,N_1595);
nor U1676 (N_1676,N_1583,N_1523);
or U1677 (N_1677,N_1572,N_1560);
nor U1678 (N_1678,N_1524,N_1557);
nor U1679 (N_1679,N_1532,N_1535);
or U1680 (N_1680,N_1503,N_1586);
or U1681 (N_1681,N_1538,N_1542);
nand U1682 (N_1682,N_1579,N_1576);
nand U1683 (N_1683,N_1503,N_1545);
or U1684 (N_1684,N_1538,N_1548);
and U1685 (N_1685,N_1552,N_1595);
nand U1686 (N_1686,N_1554,N_1567);
nand U1687 (N_1687,N_1539,N_1510);
or U1688 (N_1688,N_1503,N_1582);
or U1689 (N_1689,N_1547,N_1552);
or U1690 (N_1690,N_1552,N_1571);
nand U1691 (N_1691,N_1572,N_1577);
nand U1692 (N_1692,N_1593,N_1534);
nor U1693 (N_1693,N_1513,N_1502);
and U1694 (N_1694,N_1587,N_1598);
and U1695 (N_1695,N_1513,N_1527);
nand U1696 (N_1696,N_1598,N_1572);
nor U1697 (N_1697,N_1564,N_1560);
or U1698 (N_1698,N_1565,N_1573);
or U1699 (N_1699,N_1541,N_1502);
nor U1700 (N_1700,N_1682,N_1690);
and U1701 (N_1701,N_1635,N_1683);
nor U1702 (N_1702,N_1643,N_1652);
and U1703 (N_1703,N_1674,N_1638);
nor U1704 (N_1704,N_1624,N_1697);
nand U1705 (N_1705,N_1678,N_1650);
xnor U1706 (N_1706,N_1689,N_1601);
and U1707 (N_1707,N_1636,N_1691);
nand U1708 (N_1708,N_1603,N_1628);
nor U1709 (N_1709,N_1669,N_1633);
and U1710 (N_1710,N_1607,N_1618);
and U1711 (N_1711,N_1660,N_1639);
nand U1712 (N_1712,N_1613,N_1694);
nor U1713 (N_1713,N_1688,N_1699);
or U1714 (N_1714,N_1680,N_1667);
and U1715 (N_1715,N_1696,N_1631);
or U1716 (N_1716,N_1646,N_1671);
and U1717 (N_1717,N_1645,N_1640);
or U1718 (N_1718,N_1614,N_1644);
nand U1719 (N_1719,N_1679,N_1661);
nand U1720 (N_1720,N_1658,N_1654);
nand U1721 (N_1721,N_1606,N_1656);
or U1722 (N_1722,N_1622,N_1626);
nor U1723 (N_1723,N_1670,N_1609);
and U1724 (N_1724,N_1625,N_1685);
nand U1725 (N_1725,N_1637,N_1634);
or U1726 (N_1726,N_1630,N_1611);
nand U1727 (N_1727,N_1672,N_1649);
nand U1728 (N_1728,N_1627,N_1632);
nor U1729 (N_1729,N_1657,N_1653);
and U1730 (N_1730,N_1648,N_1647);
and U1731 (N_1731,N_1687,N_1681);
nor U1732 (N_1732,N_1620,N_1695);
nand U1733 (N_1733,N_1668,N_1673);
nand U1734 (N_1734,N_1662,N_1604);
or U1735 (N_1735,N_1608,N_1686);
nand U1736 (N_1736,N_1623,N_1664);
nand U1737 (N_1737,N_1602,N_1677);
or U1738 (N_1738,N_1666,N_1663);
and U1739 (N_1739,N_1641,N_1612);
nor U1740 (N_1740,N_1651,N_1621);
nor U1741 (N_1741,N_1610,N_1659);
nor U1742 (N_1742,N_1665,N_1617);
nand U1743 (N_1743,N_1684,N_1642);
or U1744 (N_1744,N_1605,N_1693);
and U1745 (N_1745,N_1615,N_1616);
nor U1746 (N_1746,N_1698,N_1619);
and U1747 (N_1747,N_1629,N_1675);
and U1748 (N_1748,N_1655,N_1676);
nor U1749 (N_1749,N_1600,N_1692);
nand U1750 (N_1750,N_1625,N_1681);
nor U1751 (N_1751,N_1676,N_1636);
and U1752 (N_1752,N_1650,N_1627);
and U1753 (N_1753,N_1676,N_1669);
or U1754 (N_1754,N_1697,N_1611);
nand U1755 (N_1755,N_1648,N_1683);
or U1756 (N_1756,N_1624,N_1649);
and U1757 (N_1757,N_1644,N_1666);
or U1758 (N_1758,N_1654,N_1693);
nand U1759 (N_1759,N_1673,N_1613);
or U1760 (N_1760,N_1659,N_1615);
or U1761 (N_1761,N_1602,N_1695);
and U1762 (N_1762,N_1641,N_1625);
and U1763 (N_1763,N_1675,N_1678);
and U1764 (N_1764,N_1672,N_1643);
nand U1765 (N_1765,N_1618,N_1681);
nor U1766 (N_1766,N_1663,N_1635);
or U1767 (N_1767,N_1619,N_1659);
nand U1768 (N_1768,N_1663,N_1645);
nor U1769 (N_1769,N_1636,N_1690);
and U1770 (N_1770,N_1607,N_1660);
or U1771 (N_1771,N_1696,N_1690);
nand U1772 (N_1772,N_1639,N_1695);
or U1773 (N_1773,N_1677,N_1630);
or U1774 (N_1774,N_1648,N_1696);
and U1775 (N_1775,N_1636,N_1624);
nor U1776 (N_1776,N_1638,N_1608);
or U1777 (N_1777,N_1641,N_1672);
and U1778 (N_1778,N_1612,N_1682);
nand U1779 (N_1779,N_1616,N_1680);
nor U1780 (N_1780,N_1683,N_1661);
xor U1781 (N_1781,N_1661,N_1692);
nor U1782 (N_1782,N_1665,N_1609);
nor U1783 (N_1783,N_1619,N_1634);
or U1784 (N_1784,N_1648,N_1687);
or U1785 (N_1785,N_1614,N_1657);
nor U1786 (N_1786,N_1672,N_1658);
nor U1787 (N_1787,N_1680,N_1626);
nor U1788 (N_1788,N_1624,N_1681);
nor U1789 (N_1789,N_1614,N_1645);
nand U1790 (N_1790,N_1632,N_1623);
nor U1791 (N_1791,N_1650,N_1606);
nor U1792 (N_1792,N_1605,N_1677);
nor U1793 (N_1793,N_1671,N_1612);
and U1794 (N_1794,N_1685,N_1648);
or U1795 (N_1795,N_1672,N_1670);
nand U1796 (N_1796,N_1608,N_1641);
or U1797 (N_1797,N_1699,N_1651);
or U1798 (N_1798,N_1607,N_1666);
nor U1799 (N_1799,N_1645,N_1690);
nor U1800 (N_1800,N_1765,N_1755);
and U1801 (N_1801,N_1797,N_1773);
nand U1802 (N_1802,N_1770,N_1766);
nand U1803 (N_1803,N_1751,N_1743);
nand U1804 (N_1804,N_1706,N_1729);
or U1805 (N_1805,N_1772,N_1753);
or U1806 (N_1806,N_1715,N_1747);
or U1807 (N_1807,N_1708,N_1784);
nand U1808 (N_1808,N_1754,N_1709);
and U1809 (N_1809,N_1793,N_1734);
nor U1810 (N_1810,N_1722,N_1710);
nand U1811 (N_1811,N_1796,N_1767);
and U1812 (N_1812,N_1732,N_1738);
or U1813 (N_1813,N_1771,N_1787);
or U1814 (N_1814,N_1701,N_1728);
or U1815 (N_1815,N_1759,N_1752);
and U1816 (N_1816,N_1758,N_1739);
nor U1817 (N_1817,N_1720,N_1749);
and U1818 (N_1818,N_1727,N_1768);
xor U1819 (N_1819,N_1724,N_1774);
nand U1820 (N_1820,N_1792,N_1776);
nor U1821 (N_1821,N_1726,N_1760);
nand U1822 (N_1822,N_1712,N_1780);
nand U1823 (N_1823,N_1775,N_1781);
xor U1824 (N_1824,N_1764,N_1741);
nor U1825 (N_1825,N_1769,N_1745);
nor U1826 (N_1826,N_1795,N_1799);
nor U1827 (N_1827,N_1779,N_1782);
and U1828 (N_1828,N_1786,N_1721);
nand U1829 (N_1829,N_1704,N_1746);
or U1830 (N_1830,N_1756,N_1783);
nand U1831 (N_1831,N_1716,N_1735);
and U1832 (N_1832,N_1757,N_1762);
nor U1833 (N_1833,N_1744,N_1778);
nor U1834 (N_1834,N_1717,N_1703);
nor U1835 (N_1835,N_1702,N_1740);
nor U1836 (N_1836,N_1790,N_1718);
and U1837 (N_1837,N_1798,N_1723);
and U1838 (N_1838,N_1748,N_1777);
or U1839 (N_1839,N_1750,N_1788);
nand U1840 (N_1840,N_1730,N_1791);
nor U1841 (N_1841,N_1763,N_1785);
xor U1842 (N_1842,N_1737,N_1719);
nor U1843 (N_1843,N_1714,N_1700);
nor U1844 (N_1844,N_1794,N_1789);
or U1845 (N_1845,N_1707,N_1725);
or U1846 (N_1846,N_1761,N_1731);
nand U1847 (N_1847,N_1733,N_1742);
nand U1848 (N_1848,N_1711,N_1736);
and U1849 (N_1849,N_1713,N_1705);
nand U1850 (N_1850,N_1708,N_1727);
and U1851 (N_1851,N_1790,N_1708);
and U1852 (N_1852,N_1723,N_1791);
nand U1853 (N_1853,N_1797,N_1790);
nor U1854 (N_1854,N_1700,N_1713);
nand U1855 (N_1855,N_1770,N_1748);
or U1856 (N_1856,N_1774,N_1705);
and U1857 (N_1857,N_1733,N_1724);
and U1858 (N_1858,N_1790,N_1719);
and U1859 (N_1859,N_1787,N_1737);
or U1860 (N_1860,N_1743,N_1745);
and U1861 (N_1861,N_1701,N_1743);
or U1862 (N_1862,N_1711,N_1778);
and U1863 (N_1863,N_1761,N_1795);
or U1864 (N_1864,N_1781,N_1714);
or U1865 (N_1865,N_1781,N_1774);
and U1866 (N_1866,N_1716,N_1721);
nand U1867 (N_1867,N_1790,N_1780);
or U1868 (N_1868,N_1775,N_1771);
nand U1869 (N_1869,N_1713,N_1755);
nor U1870 (N_1870,N_1729,N_1740);
nor U1871 (N_1871,N_1746,N_1785);
and U1872 (N_1872,N_1771,N_1776);
and U1873 (N_1873,N_1704,N_1723);
and U1874 (N_1874,N_1742,N_1725);
nor U1875 (N_1875,N_1755,N_1747);
nor U1876 (N_1876,N_1769,N_1732);
nor U1877 (N_1877,N_1753,N_1721);
nor U1878 (N_1878,N_1708,N_1715);
nor U1879 (N_1879,N_1771,N_1793);
or U1880 (N_1880,N_1727,N_1742);
or U1881 (N_1881,N_1747,N_1757);
or U1882 (N_1882,N_1715,N_1742);
nor U1883 (N_1883,N_1727,N_1714);
nand U1884 (N_1884,N_1730,N_1787);
nor U1885 (N_1885,N_1777,N_1714);
nand U1886 (N_1886,N_1755,N_1742);
nor U1887 (N_1887,N_1723,N_1731);
and U1888 (N_1888,N_1784,N_1798);
or U1889 (N_1889,N_1742,N_1744);
nand U1890 (N_1890,N_1784,N_1700);
or U1891 (N_1891,N_1717,N_1743);
nand U1892 (N_1892,N_1716,N_1747);
nand U1893 (N_1893,N_1750,N_1735);
nand U1894 (N_1894,N_1754,N_1748);
and U1895 (N_1895,N_1714,N_1769);
nand U1896 (N_1896,N_1795,N_1703);
nand U1897 (N_1897,N_1787,N_1721);
nand U1898 (N_1898,N_1734,N_1732);
and U1899 (N_1899,N_1782,N_1728);
xor U1900 (N_1900,N_1864,N_1883);
and U1901 (N_1901,N_1811,N_1809);
nor U1902 (N_1902,N_1893,N_1837);
nor U1903 (N_1903,N_1822,N_1807);
nand U1904 (N_1904,N_1801,N_1812);
nor U1905 (N_1905,N_1895,N_1834);
nand U1906 (N_1906,N_1850,N_1823);
nand U1907 (N_1907,N_1863,N_1886);
nand U1908 (N_1908,N_1856,N_1844);
nor U1909 (N_1909,N_1871,N_1820);
nor U1910 (N_1910,N_1840,N_1876);
or U1911 (N_1911,N_1877,N_1880);
nor U1912 (N_1912,N_1814,N_1838);
nor U1913 (N_1913,N_1860,N_1831);
nor U1914 (N_1914,N_1867,N_1832);
nor U1915 (N_1915,N_1841,N_1824);
nand U1916 (N_1916,N_1804,N_1842);
or U1917 (N_1917,N_1874,N_1819);
and U1918 (N_1918,N_1887,N_1805);
or U1919 (N_1919,N_1894,N_1869);
nand U1920 (N_1920,N_1833,N_1881);
nand U1921 (N_1921,N_1828,N_1866);
and U1922 (N_1922,N_1810,N_1843);
or U1923 (N_1923,N_1897,N_1854);
nor U1924 (N_1924,N_1846,N_1839);
nand U1925 (N_1925,N_1890,N_1862);
or U1926 (N_1926,N_1879,N_1885);
nand U1927 (N_1927,N_1891,N_1821);
or U1928 (N_1928,N_1870,N_1813);
or U1929 (N_1929,N_1889,N_1829);
nor U1930 (N_1930,N_1835,N_1892);
nor U1931 (N_1931,N_1899,N_1848);
nor U1932 (N_1932,N_1800,N_1827);
and U1933 (N_1933,N_1888,N_1808);
nor U1934 (N_1934,N_1836,N_1817);
and U1935 (N_1935,N_1857,N_1875);
nand U1936 (N_1936,N_1847,N_1868);
and U1937 (N_1937,N_1882,N_1859);
nor U1938 (N_1938,N_1802,N_1849);
nand U1939 (N_1939,N_1896,N_1873);
nand U1940 (N_1940,N_1872,N_1825);
nand U1941 (N_1941,N_1803,N_1852);
and U1942 (N_1942,N_1826,N_1806);
or U1943 (N_1943,N_1816,N_1858);
and U1944 (N_1944,N_1851,N_1818);
nand U1945 (N_1945,N_1861,N_1878);
nand U1946 (N_1946,N_1865,N_1853);
nor U1947 (N_1947,N_1884,N_1830);
nand U1948 (N_1948,N_1845,N_1815);
or U1949 (N_1949,N_1898,N_1855);
nand U1950 (N_1950,N_1834,N_1881);
nor U1951 (N_1951,N_1889,N_1864);
or U1952 (N_1952,N_1869,N_1879);
nor U1953 (N_1953,N_1899,N_1825);
and U1954 (N_1954,N_1886,N_1828);
nand U1955 (N_1955,N_1800,N_1860);
or U1956 (N_1956,N_1831,N_1870);
and U1957 (N_1957,N_1861,N_1889);
or U1958 (N_1958,N_1851,N_1830);
nor U1959 (N_1959,N_1807,N_1856);
or U1960 (N_1960,N_1817,N_1840);
or U1961 (N_1961,N_1822,N_1894);
or U1962 (N_1962,N_1808,N_1825);
nor U1963 (N_1963,N_1871,N_1882);
and U1964 (N_1964,N_1894,N_1855);
nor U1965 (N_1965,N_1821,N_1806);
nor U1966 (N_1966,N_1846,N_1826);
nor U1967 (N_1967,N_1846,N_1884);
nand U1968 (N_1968,N_1809,N_1805);
or U1969 (N_1969,N_1829,N_1872);
nand U1970 (N_1970,N_1889,N_1847);
nand U1971 (N_1971,N_1815,N_1892);
nand U1972 (N_1972,N_1893,N_1845);
or U1973 (N_1973,N_1893,N_1812);
nor U1974 (N_1974,N_1833,N_1810);
or U1975 (N_1975,N_1824,N_1828);
or U1976 (N_1976,N_1878,N_1810);
and U1977 (N_1977,N_1890,N_1838);
and U1978 (N_1978,N_1864,N_1887);
or U1979 (N_1979,N_1892,N_1811);
nor U1980 (N_1980,N_1824,N_1821);
nor U1981 (N_1981,N_1884,N_1856);
nand U1982 (N_1982,N_1876,N_1894);
nor U1983 (N_1983,N_1844,N_1819);
nand U1984 (N_1984,N_1839,N_1845);
and U1985 (N_1985,N_1894,N_1810);
or U1986 (N_1986,N_1801,N_1858);
or U1987 (N_1987,N_1873,N_1801);
and U1988 (N_1988,N_1892,N_1870);
nand U1989 (N_1989,N_1811,N_1856);
and U1990 (N_1990,N_1878,N_1884);
nand U1991 (N_1991,N_1896,N_1867);
nor U1992 (N_1992,N_1897,N_1862);
nand U1993 (N_1993,N_1804,N_1828);
or U1994 (N_1994,N_1821,N_1838);
and U1995 (N_1995,N_1882,N_1875);
or U1996 (N_1996,N_1824,N_1857);
and U1997 (N_1997,N_1845,N_1878);
nand U1998 (N_1998,N_1865,N_1861);
and U1999 (N_1999,N_1889,N_1806);
and U2000 (N_2000,N_1941,N_1914);
or U2001 (N_2001,N_1935,N_1982);
or U2002 (N_2002,N_1952,N_1938);
or U2003 (N_2003,N_1943,N_1984);
nand U2004 (N_2004,N_1964,N_1910);
nor U2005 (N_2005,N_1936,N_1996);
or U2006 (N_2006,N_1993,N_1921);
or U2007 (N_2007,N_1928,N_1909);
nand U2008 (N_2008,N_1908,N_1973);
and U2009 (N_2009,N_1981,N_1934);
nor U2010 (N_2010,N_1916,N_1995);
or U2011 (N_2011,N_1951,N_1991);
nand U2012 (N_2012,N_1968,N_1923);
or U2013 (N_2013,N_1912,N_1937);
nor U2014 (N_2014,N_1927,N_1966);
nor U2015 (N_2015,N_1930,N_1929);
nor U2016 (N_2016,N_1940,N_1925);
and U2017 (N_2017,N_1974,N_1922);
and U2018 (N_2018,N_1945,N_1946);
or U2019 (N_2019,N_1975,N_1917);
nand U2020 (N_2020,N_1944,N_1939);
nand U2021 (N_2021,N_1972,N_1915);
or U2022 (N_2022,N_1997,N_1901);
and U2023 (N_2023,N_1920,N_1989);
and U2024 (N_2024,N_1947,N_1977);
or U2025 (N_2025,N_1978,N_1988);
nand U2026 (N_2026,N_1924,N_1953);
and U2027 (N_2027,N_1942,N_1956);
and U2028 (N_2028,N_1959,N_1933);
nor U2029 (N_2029,N_1954,N_1987);
nor U2030 (N_2030,N_1986,N_1961);
xor U2031 (N_2031,N_1949,N_1963);
and U2032 (N_2032,N_1970,N_1960);
or U2033 (N_2033,N_1980,N_1950);
nor U2034 (N_2034,N_1976,N_1992);
or U2035 (N_2035,N_1932,N_1955);
or U2036 (N_2036,N_1999,N_1903);
nand U2037 (N_2037,N_1958,N_1919);
and U2038 (N_2038,N_1983,N_1931);
and U2039 (N_2039,N_1979,N_1971);
nand U2040 (N_2040,N_1998,N_1913);
nor U2041 (N_2041,N_1967,N_1905);
nand U2042 (N_2042,N_1900,N_1906);
or U2043 (N_2043,N_1990,N_1904);
and U2044 (N_2044,N_1926,N_1965);
nand U2045 (N_2045,N_1911,N_1994);
and U2046 (N_2046,N_1985,N_1962);
nand U2047 (N_2047,N_1969,N_1907);
and U2048 (N_2048,N_1948,N_1957);
or U2049 (N_2049,N_1902,N_1918);
nand U2050 (N_2050,N_1941,N_1901);
nor U2051 (N_2051,N_1965,N_1935);
nor U2052 (N_2052,N_1937,N_1953);
nand U2053 (N_2053,N_1923,N_1917);
nand U2054 (N_2054,N_1920,N_1986);
or U2055 (N_2055,N_1991,N_1936);
and U2056 (N_2056,N_1959,N_1998);
or U2057 (N_2057,N_1948,N_1965);
or U2058 (N_2058,N_1961,N_1946);
nand U2059 (N_2059,N_1974,N_1918);
nor U2060 (N_2060,N_1997,N_1928);
nor U2061 (N_2061,N_1933,N_1925);
and U2062 (N_2062,N_1972,N_1984);
nor U2063 (N_2063,N_1965,N_1980);
nand U2064 (N_2064,N_1963,N_1929);
and U2065 (N_2065,N_1907,N_1919);
or U2066 (N_2066,N_1946,N_1964);
or U2067 (N_2067,N_1923,N_1959);
and U2068 (N_2068,N_1982,N_1923);
nor U2069 (N_2069,N_1983,N_1922);
and U2070 (N_2070,N_1982,N_1941);
and U2071 (N_2071,N_1968,N_1943);
nand U2072 (N_2072,N_1965,N_1944);
and U2073 (N_2073,N_1986,N_1942);
and U2074 (N_2074,N_1957,N_1970);
and U2075 (N_2075,N_1979,N_1907);
nand U2076 (N_2076,N_1915,N_1994);
nand U2077 (N_2077,N_1969,N_1947);
and U2078 (N_2078,N_1956,N_1901);
nor U2079 (N_2079,N_1982,N_1961);
nand U2080 (N_2080,N_1977,N_1990);
or U2081 (N_2081,N_1985,N_1901);
nand U2082 (N_2082,N_1932,N_1928);
nand U2083 (N_2083,N_1959,N_1930);
nor U2084 (N_2084,N_1962,N_1964);
and U2085 (N_2085,N_1908,N_1943);
or U2086 (N_2086,N_1930,N_1984);
nand U2087 (N_2087,N_1963,N_1935);
nor U2088 (N_2088,N_1927,N_1929);
nand U2089 (N_2089,N_1962,N_1926);
nor U2090 (N_2090,N_1990,N_1937);
nor U2091 (N_2091,N_1981,N_1972);
nand U2092 (N_2092,N_1933,N_1943);
and U2093 (N_2093,N_1952,N_1994);
nor U2094 (N_2094,N_1911,N_1952);
nor U2095 (N_2095,N_1998,N_1943);
nand U2096 (N_2096,N_1913,N_1918);
or U2097 (N_2097,N_1965,N_1956);
or U2098 (N_2098,N_1954,N_1964);
nand U2099 (N_2099,N_1915,N_1903);
or U2100 (N_2100,N_2001,N_2089);
nand U2101 (N_2101,N_2022,N_2087);
nor U2102 (N_2102,N_2030,N_2073);
or U2103 (N_2103,N_2036,N_2086);
and U2104 (N_2104,N_2035,N_2034);
and U2105 (N_2105,N_2096,N_2027);
and U2106 (N_2106,N_2000,N_2011);
or U2107 (N_2107,N_2052,N_2049);
and U2108 (N_2108,N_2041,N_2032);
nor U2109 (N_2109,N_2066,N_2021);
and U2110 (N_2110,N_2048,N_2084);
nor U2111 (N_2111,N_2031,N_2044);
nand U2112 (N_2112,N_2069,N_2024);
or U2113 (N_2113,N_2046,N_2054);
nand U2114 (N_2114,N_2014,N_2010);
nor U2115 (N_2115,N_2016,N_2023);
or U2116 (N_2116,N_2051,N_2009);
nand U2117 (N_2117,N_2047,N_2078);
and U2118 (N_2118,N_2040,N_2002);
nor U2119 (N_2119,N_2062,N_2063);
nand U2120 (N_2120,N_2098,N_2017);
nor U2121 (N_2121,N_2072,N_2042);
nand U2122 (N_2122,N_2037,N_2043);
or U2123 (N_2123,N_2094,N_2003);
or U2124 (N_2124,N_2095,N_2065);
nand U2125 (N_2125,N_2053,N_2033);
or U2126 (N_2126,N_2081,N_2056);
or U2127 (N_2127,N_2064,N_2079);
and U2128 (N_2128,N_2055,N_2008);
or U2129 (N_2129,N_2071,N_2020);
nand U2130 (N_2130,N_2088,N_2007);
nand U2131 (N_2131,N_2090,N_2059);
nor U2132 (N_2132,N_2074,N_2038);
nor U2133 (N_2133,N_2082,N_2099);
nand U2134 (N_2134,N_2025,N_2068);
and U2135 (N_2135,N_2019,N_2092);
nand U2136 (N_2136,N_2039,N_2075);
nor U2137 (N_2137,N_2026,N_2060);
or U2138 (N_2138,N_2045,N_2006);
or U2139 (N_2139,N_2097,N_2076);
and U2140 (N_2140,N_2004,N_2029);
nor U2141 (N_2141,N_2067,N_2012);
nand U2142 (N_2142,N_2077,N_2061);
nand U2143 (N_2143,N_2091,N_2058);
nand U2144 (N_2144,N_2015,N_2028);
nand U2145 (N_2145,N_2093,N_2085);
and U2146 (N_2146,N_2005,N_2070);
and U2147 (N_2147,N_2057,N_2018);
and U2148 (N_2148,N_2083,N_2013);
nand U2149 (N_2149,N_2050,N_2080);
and U2150 (N_2150,N_2053,N_2000);
or U2151 (N_2151,N_2049,N_2078);
nand U2152 (N_2152,N_2088,N_2017);
or U2153 (N_2153,N_2072,N_2016);
or U2154 (N_2154,N_2008,N_2096);
nand U2155 (N_2155,N_2004,N_2016);
and U2156 (N_2156,N_2006,N_2000);
and U2157 (N_2157,N_2036,N_2023);
nor U2158 (N_2158,N_2058,N_2017);
xnor U2159 (N_2159,N_2069,N_2020);
or U2160 (N_2160,N_2061,N_2027);
and U2161 (N_2161,N_2003,N_2005);
nand U2162 (N_2162,N_2091,N_2087);
and U2163 (N_2163,N_2029,N_2045);
and U2164 (N_2164,N_2004,N_2062);
nor U2165 (N_2165,N_2044,N_2057);
nor U2166 (N_2166,N_2034,N_2073);
nand U2167 (N_2167,N_2026,N_2076);
or U2168 (N_2168,N_2093,N_2084);
nor U2169 (N_2169,N_2060,N_2007);
nand U2170 (N_2170,N_2054,N_2086);
and U2171 (N_2171,N_2084,N_2028);
and U2172 (N_2172,N_2047,N_2023);
nor U2173 (N_2173,N_2037,N_2071);
or U2174 (N_2174,N_2062,N_2098);
and U2175 (N_2175,N_2059,N_2097);
or U2176 (N_2176,N_2097,N_2019);
nor U2177 (N_2177,N_2091,N_2071);
nand U2178 (N_2178,N_2001,N_2041);
nand U2179 (N_2179,N_2033,N_2008);
nor U2180 (N_2180,N_2088,N_2060);
and U2181 (N_2181,N_2080,N_2055);
or U2182 (N_2182,N_2084,N_2021);
or U2183 (N_2183,N_2067,N_2022);
or U2184 (N_2184,N_2027,N_2010);
or U2185 (N_2185,N_2060,N_2019);
nand U2186 (N_2186,N_2035,N_2058);
nor U2187 (N_2187,N_2000,N_2071);
nor U2188 (N_2188,N_2030,N_2072);
or U2189 (N_2189,N_2017,N_2025);
nand U2190 (N_2190,N_2051,N_2056);
or U2191 (N_2191,N_2070,N_2079);
nor U2192 (N_2192,N_2017,N_2037);
and U2193 (N_2193,N_2029,N_2008);
nor U2194 (N_2194,N_2030,N_2021);
nand U2195 (N_2195,N_2058,N_2085);
or U2196 (N_2196,N_2017,N_2053);
or U2197 (N_2197,N_2044,N_2084);
and U2198 (N_2198,N_2056,N_2040);
nand U2199 (N_2199,N_2003,N_2039);
nand U2200 (N_2200,N_2144,N_2147);
nand U2201 (N_2201,N_2118,N_2179);
and U2202 (N_2202,N_2199,N_2172);
nor U2203 (N_2203,N_2191,N_2173);
and U2204 (N_2204,N_2153,N_2194);
or U2205 (N_2205,N_2115,N_2138);
or U2206 (N_2206,N_2142,N_2193);
and U2207 (N_2207,N_2160,N_2148);
nor U2208 (N_2208,N_2110,N_2152);
nor U2209 (N_2209,N_2109,N_2143);
nor U2210 (N_2210,N_2105,N_2124);
nor U2211 (N_2211,N_2184,N_2111);
nand U2212 (N_2212,N_2154,N_2121);
or U2213 (N_2213,N_2103,N_2188);
or U2214 (N_2214,N_2185,N_2134);
nand U2215 (N_2215,N_2159,N_2132);
and U2216 (N_2216,N_2125,N_2137);
and U2217 (N_2217,N_2180,N_2139);
or U2218 (N_2218,N_2129,N_2100);
nor U2219 (N_2219,N_2119,N_2146);
nor U2220 (N_2220,N_2196,N_2130);
or U2221 (N_2221,N_2128,N_2106);
nor U2222 (N_2222,N_2187,N_2101);
and U2223 (N_2223,N_2150,N_2116);
or U2224 (N_2224,N_2169,N_2113);
nor U2225 (N_2225,N_2177,N_2151);
nand U2226 (N_2226,N_2165,N_2197);
nor U2227 (N_2227,N_2135,N_2190);
or U2228 (N_2228,N_2123,N_2104);
and U2229 (N_2229,N_2126,N_2161);
nor U2230 (N_2230,N_2186,N_2107);
nand U2231 (N_2231,N_2192,N_2181);
or U2232 (N_2232,N_2195,N_2183);
and U2233 (N_2233,N_2163,N_2170);
nand U2234 (N_2234,N_2158,N_2171);
or U2235 (N_2235,N_2108,N_2198);
nor U2236 (N_2236,N_2189,N_2176);
nand U2237 (N_2237,N_2168,N_2122);
nor U2238 (N_2238,N_2102,N_2114);
nand U2239 (N_2239,N_2178,N_2164);
nand U2240 (N_2240,N_2162,N_2166);
nor U2241 (N_2241,N_2117,N_2131);
nor U2242 (N_2242,N_2127,N_2112);
xor U2243 (N_2243,N_2136,N_2175);
nand U2244 (N_2244,N_2133,N_2145);
nor U2245 (N_2245,N_2182,N_2155);
nor U2246 (N_2246,N_2156,N_2157);
and U2247 (N_2247,N_2140,N_2141);
nor U2248 (N_2248,N_2120,N_2174);
and U2249 (N_2249,N_2167,N_2149);
and U2250 (N_2250,N_2135,N_2123);
nand U2251 (N_2251,N_2194,N_2156);
or U2252 (N_2252,N_2123,N_2142);
nand U2253 (N_2253,N_2134,N_2125);
and U2254 (N_2254,N_2103,N_2154);
and U2255 (N_2255,N_2136,N_2182);
nor U2256 (N_2256,N_2145,N_2115);
and U2257 (N_2257,N_2100,N_2128);
nand U2258 (N_2258,N_2188,N_2184);
and U2259 (N_2259,N_2107,N_2184);
nor U2260 (N_2260,N_2197,N_2179);
and U2261 (N_2261,N_2197,N_2133);
and U2262 (N_2262,N_2184,N_2138);
nand U2263 (N_2263,N_2116,N_2158);
nor U2264 (N_2264,N_2110,N_2138);
or U2265 (N_2265,N_2194,N_2178);
nand U2266 (N_2266,N_2192,N_2186);
and U2267 (N_2267,N_2129,N_2116);
nand U2268 (N_2268,N_2176,N_2187);
nand U2269 (N_2269,N_2106,N_2155);
and U2270 (N_2270,N_2154,N_2122);
and U2271 (N_2271,N_2124,N_2100);
or U2272 (N_2272,N_2140,N_2161);
nand U2273 (N_2273,N_2102,N_2136);
and U2274 (N_2274,N_2139,N_2131);
nand U2275 (N_2275,N_2182,N_2107);
nand U2276 (N_2276,N_2189,N_2132);
nor U2277 (N_2277,N_2168,N_2105);
nor U2278 (N_2278,N_2129,N_2106);
nand U2279 (N_2279,N_2196,N_2184);
nand U2280 (N_2280,N_2101,N_2136);
and U2281 (N_2281,N_2130,N_2183);
nor U2282 (N_2282,N_2182,N_2180);
and U2283 (N_2283,N_2146,N_2195);
xor U2284 (N_2284,N_2109,N_2141);
nor U2285 (N_2285,N_2103,N_2146);
nand U2286 (N_2286,N_2172,N_2191);
nand U2287 (N_2287,N_2142,N_2113);
or U2288 (N_2288,N_2125,N_2128);
or U2289 (N_2289,N_2189,N_2192);
nor U2290 (N_2290,N_2100,N_2133);
nor U2291 (N_2291,N_2182,N_2138);
or U2292 (N_2292,N_2100,N_2157);
and U2293 (N_2293,N_2117,N_2193);
nor U2294 (N_2294,N_2159,N_2164);
nor U2295 (N_2295,N_2184,N_2135);
nor U2296 (N_2296,N_2141,N_2108);
or U2297 (N_2297,N_2190,N_2159);
nand U2298 (N_2298,N_2118,N_2119);
or U2299 (N_2299,N_2133,N_2144);
or U2300 (N_2300,N_2214,N_2259);
or U2301 (N_2301,N_2200,N_2257);
or U2302 (N_2302,N_2203,N_2206);
or U2303 (N_2303,N_2281,N_2225);
nor U2304 (N_2304,N_2204,N_2285);
nor U2305 (N_2305,N_2222,N_2266);
and U2306 (N_2306,N_2273,N_2243);
nor U2307 (N_2307,N_2210,N_2253);
or U2308 (N_2308,N_2224,N_2230);
or U2309 (N_2309,N_2209,N_2233);
nand U2310 (N_2310,N_2249,N_2292);
and U2311 (N_2311,N_2289,N_2239);
and U2312 (N_2312,N_2265,N_2201);
or U2313 (N_2313,N_2254,N_2279);
or U2314 (N_2314,N_2264,N_2271);
or U2315 (N_2315,N_2255,N_2241);
or U2316 (N_2316,N_2238,N_2261);
xor U2317 (N_2317,N_2234,N_2226);
nand U2318 (N_2318,N_2220,N_2227);
and U2319 (N_2319,N_2297,N_2256);
and U2320 (N_2320,N_2216,N_2269);
nor U2321 (N_2321,N_2237,N_2283);
or U2322 (N_2322,N_2250,N_2231);
nand U2323 (N_2323,N_2208,N_2267);
and U2324 (N_2324,N_2282,N_2258);
nor U2325 (N_2325,N_2221,N_2240);
nor U2326 (N_2326,N_2290,N_2235);
nor U2327 (N_2327,N_2280,N_2244);
nand U2328 (N_2328,N_2268,N_2278);
nor U2329 (N_2329,N_2270,N_2218);
nand U2330 (N_2330,N_2223,N_2291);
or U2331 (N_2331,N_2217,N_2288);
nor U2332 (N_2332,N_2274,N_2276);
and U2333 (N_2333,N_2245,N_2262);
or U2334 (N_2334,N_2251,N_2205);
nand U2335 (N_2335,N_2207,N_2293);
and U2336 (N_2336,N_2284,N_2248);
nand U2337 (N_2337,N_2298,N_2286);
nand U2338 (N_2338,N_2242,N_2219);
or U2339 (N_2339,N_2232,N_2263);
nor U2340 (N_2340,N_2215,N_2211);
and U2341 (N_2341,N_2246,N_2229);
or U2342 (N_2342,N_2213,N_2294);
and U2343 (N_2343,N_2202,N_2212);
or U2344 (N_2344,N_2275,N_2287);
and U2345 (N_2345,N_2247,N_2272);
nor U2346 (N_2346,N_2277,N_2228);
nor U2347 (N_2347,N_2236,N_2260);
nor U2348 (N_2348,N_2252,N_2296);
or U2349 (N_2349,N_2299,N_2295);
or U2350 (N_2350,N_2298,N_2238);
nand U2351 (N_2351,N_2296,N_2208);
or U2352 (N_2352,N_2201,N_2228);
nand U2353 (N_2353,N_2219,N_2218);
and U2354 (N_2354,N_2213,N_2244);
nor U2355 (N_2355,N_2228,N_2293);
xor U2356 (N_2356,N_2286,N_2261);
nand U2357 (N_2357,N_2225,N_2235);
or U2358 (N_2358,N_2289,N_2260);
nor U2359 (N_2359,N_2211,N_2263);
nand U2360 (N_2360,N_2239,N_2274);
or U2361 (N_2361,N_2208,N_2299);
nor U2362 (N_2362,N_2284,N_2252);
and U2363 (N_2363,N_2250,N_2215);
or U2364 (N_2364,N_2298,N_2256);
xnor U2365 (N_2365,N_2219,N_2226);
and U2366 (N_2366,N_2219,N_2236);
nand U2367 (N_2367,N_2268,N_2233);
and U2368 (N_2368,N_2291,N_2220);
or U2369 (N_2369,N_2241,N_2226);
nor U2370 (N_2370,N_2257,N_2223);
nor U2371 (N_2371,N_2274,N_2296);
nand U2372 (N_2372,N_2256,N_2264);
or U2373 (N_2373,N_2246,N_2239);
and U2374 (N_2374,N_2293,N_2248);
nor U2375 (N_2375,N_2212,N_2236);
or U2376 (N_2376,N_2263,N_2279);
or U2377 (N_2377,N_2259,N_2250);
nor U2378 (N_2378,N_2297,N_2215);
and U2379 (N_2379,N_2287,N_2241);
and U2380 (N_2380,N_2239,N_2280);
or U2381 (N_2381,N_2216,N_2285);
or U2382 (N_2382,N_2237,N_2241);
or U2383 (N_2383,N_2229,N_2286);
nor U2384 (N_2384,N_2269,N_2286);
nand U2385 (N_2385,N_2298,N_2222);
nor U2386 (N_2386,N_2218,N_2202);
and U2387 (N_2387,N_2235,N_2271);
and U2388 (N_2388,N_2262,N_2243);
or U2389 (N_2389,N_2281,N_2290);
nand U2390 (N_2390,N_2293,N_2282);
or U2391 (N_2391,N_2209,N_2247);
and U2392 (N_2392,N_2258,N_2259);
and U2393 (N_2393,N_2260,N_2224);
or U2394 (N_2394,N_2288,N_2228);
and U2395 (N_2395,N_2200,N_2201);
nor U2396 (N_2396,N_2203,N_2265);
or U2397 (N_2397,N_2246,N_2213);
nor U2398 (N_2398,N_2245,N_2288);
nor U2399 (N_2399,N_2256,N_2208);
and U2400 (N_2400,N_2337,N_2347);
or U2401 (N_2401,N_2346,N_2342);
or U2402 (N_2402,N_2389,N_2390);
and U2403 (N_2403,N_2334,N_2303);
nand U2404 (N_2404,N_2375,N_2357);
nor U2405 (N_2405,N_2398,N_2333);
nand U2406 (N_2406,N_2376,N_2354);
nor U2407 (N_2407,N_2345,N_2332);
and U2408 (N_2408,N_2322,N_2309);
nand U2409 (N_2409,N_2329,N_2349);
and U2410 (N_2410,N_2340,N_2310);
nand U2411 (N_2411,N_2391,N_2317);
or U2412 (N_2412,N_2331,N_2328);
or U2413 (N_2413,N_2348,N_2314);
or U2414 (N_2414,N_2387,N_2311);
or U2415 (N_2415,N_2397,N_2304);
and U2416 (N_2416,N_2306,N_2338);
or U2417 (N_2417,N_2301,N_2393);
nand U2418 (N_2418,N_2350,N_2369);
nor U2419 (N_2419,N_2382,N_2365);
nand U2420 (N_2420,N_2377,N_2330);
nor U2421 (N_2421,N_2355,N_2313);
and U2422 (N_2422,N_2308,N_2305);
and U2423 (N_2423,N_2378,N_2363);
nor U2424 (N_2424,N_2362,N_2385);
and U2425 (N_2425,N_2392,N_2388);
and U2426 (N_2426,N_2370,N_2379);
nand U2427 (N_2427,N_2352,N_2384);
nand U2428 (N_2428,N_2373,N_2315);
or U2429 (N_2429,N_2320,N_2321);
or U2430 (N_2430,N_2364,N_2386);
or U2431 (N_2431,N_2316,N_2318);
or U2432 (N_2432,N_2399,N_2383);
and U2433 (N_2433,N_2371,N_2374);
and U2434 (N_2434,N_2323,N_2396);
or U2435 (N_2435,N_2351,N_2336);
and U2436 (N_2436,N_2339,N_2344);
and U2437 (N_2437,N_2326,N_2394);
nand U2438 (N_2438,N_2325,N_2312);
or U2439 (N_2439,N_2324,N_2327);
nand U2440 (N_2440,N_2307,N_2341);
and U2441 (N_2441,N_2300,N_2335);
or U2442 (N_2442,N_2358,N_2395);
or U2443 (N_2443,N_2372,N_2319);
nand U2444 (N_2444,N_2353,N_2368);
nor U2445 (N_2445,N_2343,N_2381);
and U2446 (N_2446,N_2380,N_2359);
nand U2447 (N_2447,N_2360,N_2356);
or U2448 (N_2448,N_2361,N_2367);
nand U2449 (N_2449,N_2302,N_2366);
and U2450 (N_2450,N_2328,N_2323);
nor U2451 (N_2451,N_2319,N_2395);
and U2452 (N_2452,N_2389,N_2347);
nand U2453 (N_2453,N_2346,N_2336);
and U2454 (N_2454,N_2338,N_2368);
and U2455 (N_2455,N_2320,N_2351);
nand U2456 (N_2456,N_2316,N_2305);
and U2457 (N_2457,N_2311,N_2337);
and U2458 (N_2458,N_2352,N_2371);
nand U2459 (N_2459,N_2342,N_2378);
nor U2460 (N_2460,N_2334,N_2369);
or U2461 (N_2461,N_2319,N_2327);
nor U2462 (N_2462,N_2324,N_2369);
or U2463 (N_2463,N_2376,N_2391);
or U2464 (N_2464,N_2348,N_2347);
or U2465 (N_2465,N_2365,N_2354);
nor U2466 (N_2466,N_2318,N_2319);
nand U2467 (N_2467,N_2359,N_2376);
nor U2468 (N_2468,N_2347,N_2357);
and U2469 (N_2469,N_2309,N_2311);
nor U2470 (N_2470,N_2341,N_2375);
and U2471 (N_2471,N_2312,N_2338);
and U2472 (N_2472,N_2318,N_2360);
nand U2473 (N_2473,N_2313,N_2373);
nand U2474 (N_2474,N_2387,N_2313);
or U2475 (N_2475,N_2314,N_2319);
and U2476 (N_2476,N_2370,N_2386);
or U2477 (N_2477,N_2386,N_2339);
or U2478 (N_2478,N_2326,N_2334);
and U2479 (N_2479,N_2361,N_2327);
nor U2480 (N_2480,N_2353,N_2324);
nand U2481 (N_2481,N_2365,N_2380);
or U2482 (N_2482,N_2399,N_2336);
and U2483 (N_2483,N_2315,N_2385);
or U2484 (N_2484,N_2323,N_2390);
and U2485 (N_2485,N_2327,N_2370);
and U2486 (N_2486,N_2322,N_2380);
and U2487 (N_2487,N_2362,N_2331);
nor U2488 (N_2488,N_2376,N_2394);
nor U2489 (N_2489,N_2326,N_2330);
nor U2490 (N_2490,N_2374,N_2313);
nand U2491 (N_2491,N_2362,N_2300);
or U2492 (N_2492,N_2372,N_2359);
nand U2493 (N_2493,N_2301,N_2304);
nor U2494 (N_2494,N_2307,N_2343);
or U2495 (N_2495,N_2376,N_2355);
nand U2496 (N_2496,N_2307,N_2346);
and U2497 (N_2497,N_2395,N_2348);
or U2498 (N_2498,N_2342,N_2325);
nand U2499 (N_2499,N_2388,N_2374);
xnor U2500 (N_2500,N_2429,N_2420);
nor U2501 (N_2501,N_2403,N_2497);
nor U2502 (N_2502,N_2470,N_2437);
or U2503 (N_2503,N_2453,N_2442);
and U2504 (N_2504,N_2484,N_2400);
nand U2505 (N_2505,N_2485,N_2406);
or U2506 (N_2506,N_2401,N_2443);
nor U2507 (N_2507,N_2446,N_2412);
nor U2508 (N_2508,N_2488,N_2436);
or U2509 (N_2509,N_2433,N_2483);
nor U2510 (N_2510,N_2478,N_2471);
or U2511 (N_2511,N_2460,N_2418);
nand U2512 (N_2512,N_2447,N_2431);
and U2513 (N_2513,N_2410,N_2480);
and U2514 (N_2514,N_2454,N_2452);
and U2515 (N_2515,N_2439,N_2432);
and U2516 (N_2516,N_2494,N_2416);
or U2517 (N_2517,N_2413,N_2472);
and U2518 (N_2518,N_2440,N_2493);
and U2519 (N_2519,N_2456,N_2459);
or U2520 (N_2520,N_2487,N_2491);
nand U2521 (N_2521,N_2404,N_2495);
or U2522 (N_2522,N_2457,N_2444);
or U2523 (N_2523,N_2402,N_2496);
nor U2524 (N_2524,N_2417,N_2421);
or U2525 (N_2525,N_2423,N_2408);
nand U2526 (N_2526,N_2481,N_2474);
or U2527 (N_2527,N_2490,N_2489);
and U2528 (N_2528,N_2424,N_2426);
or U2529 (N_2529,N_2448,N_2435);
and U2530 (N_2530,N_2441,N_2407);
xnor U2531 (N_2531,N_2427,N_2461);
nor U2532 (N_2532,N_2415,N_2438);
or U2533 (N_2533,N_2473,N_2468);
or U2534 (N_2534,N_2422,N_2405);
and U2535 (N_2535,N_2451,N_2498);
nand U2536 (N_2536,N_2411,N_2499);
nor U2537 (N_2537,N_2469,N_2467);
nand U2538 (N_2538,N_2477,N_2464);
xnor U2539 (N_2539,N_2428,N_2445);
nand U2540 (N_2540,N_2463,N_2425);
nor U2541 (N_2541,N_2458,N_2462);
and U2542 (N_2542,N_2476,N_2455);
and U2543 (N_2543,N_2486,N_2450);
nand U2544 (N_2544,N_2430,N_2434);
nand U2545 (N_2545,N_2409,N_2492);
nand U2546 (N_2546,N_2419,N_2465);
and U2547 (N_2547,N_2482,N_2466);
or U2548 (N_2548,N_2414,N_2449);
nor U2549 (N_2549,N_2475,N_2479);
and U2550 (N_2550,N_2417,N_2485);
and U2551 (N_2551,N_2476,N_2474);
nand U2552 (N_2552,N_2404,N_2455);
xor U2553 (N_2553,N_2456,N_2449);
nand U2554 (N_2554,N_2451,N_2497);
or U2555 (N_2555,N_2485,N_2451);
or U2556 (N_2556,N_2441,N_2495);
nand U2557 (N_2557,N_2429,N_2402);
nor U2558 (N_2558,N_2418,N_2498);
nor U2559 (N_2559,N_2411,N_2417);
nand U2560 (N_2560,N_2493,N_2405);
and U2561 (N_2561,N_2460,N_2478);
and U2562 (N_2562,N_2422,N_2450);
nand U2563 (N_2563,N_2453,N_2466);
or U2564 (N_2564,N_2461,N_2426);
nor U2565 (N_2565,N_2487,N_2443);
nor U2566 (N_2566,N_2429,N_2426);
nor U2567 (N_2567,N_2408,N_2414);
nor U2568 (N_2568,N_2406,N_2409);
nor U2569 (N_2569,N_2421,N_2414);
or U2570 (N_2570,N_2426,N_2434);
nor U2571 (N_2571,N_2450,N_2476);
and U2572 (N_2572,N_2451,N_2442);
and U2573 (N_2573,N_2420,N_2468);
nand U2574 (N_2574,N_2445,N_2487);
nand U2575 (N_2575,N_2433,N_2469);
or U2576 (N_2576,N_2473,N_2425);
nor U2577 (N_2577,N_2421,N_2465);
nand U2578 (N_2578,N_2480,N_2402);
nor U2579 (N_2579,N_2478,N_2498);
and U2580 (N_2580,N_2422,N_2499);
nand U2581 (N_2581,N_2401,N_2475);
or U2582 (N_2582,N_2485,N_2407);
nand U2583 (N_2583,N_2494,N_2484);
or U2584 (N_2584,N_2456,N_2430);
nand U2585 (N_2585,N_2406,N_2488);
nand U2586 (N_2586,N_2485,N_2476);
nand U2587 (N_2587,N_2410,N_2429);
or U2588 (N_2588,N_2428,N_2444);
nor U2589 (N_2589,N_2461,N_2463);
nor U2590 (N_2590,N_2404,N_2492);
nor U2591 (N_2591,N_2456,N_2428);
nand U2592 (N_2592,N_2446,N_2490);
nand U2593 (N_2593,N_2432,N_2456);
and U2594 (N_2594,N_2405,N_2440);
nand U2595 (N_2595,N_2481,N_2493);
nor U2596 (N_2596,N_2480,N_2467);
nor U2597 (N_2597,N_2443,N_2469);
nor U2598 (N_2598,N_2441,N_2467);
or U2599 (N_2599,N_2479,N_2464);
nor U2600 (N_2600,N_2582,N_2502);
and U2601 (N_2601,N_2508,N_2537);
and U2602 (N_2602,N_2594,N_2542);
nor U2603 (N_2603,N_2538,N_2506);
nor U2604 (N_2604,N_2597,N_2523);
nand U2605 (N_2605,N_2522,N_2509);
or U2606 (N_2606,N_2570,N_2578);
and U2607 (N_2607,N_2500,N_2531);
nor U2608 (N_2608,N_2534,N_2564);
and U2609 (N_2609,N_2555,N_2526);
nor U2610 (N_2610,N_2579,N_2584);
and U2611 (N_2611,N_2596,N_2574);
and U2612 (N_2612,N_2503,N_2533);
nor U2613 (N_2613,N_2581,N_2572);
nor U2614 (N_2614,N_2529,N_2539);
nor U2615 (N_2615,N_2525,N_2515);
nor U2616 (N_2616,N_2549,N_2552);
and U2617 (N_2617,N_2507,N_2575);
nand U2618 (N_2618,N_2532,N_2599);
xor U2619 (N_2619,N_2545,N_2544);
nand U2620 (N_2620,N_2505,N_2521);
nand U2621 (N_2621,N_2547,N_2530);
or U2622 (N_2622,N_2556,N_2577);
and U2623 (N_2623,N_2518,N_2541);
and U2624 (N_2624,N_2548,N_2565);
nor U2625 (N_2625,N_2569,N_2519);
or U2626 (N_2626,N_2504,N_2517);
and U2627 (N_2627,N_2559,N_2540);
nand U2628 (N_2628,N_2510,N_2592);
and U2629 (N_2629,N_2591,N_2593);
or U2630 (N_2630,N_2554,N_2524);
nand U2631 (N_2631,N_2520,N_2590);
nor U2632 (N_2632,N_2511,N_2560);
nand U2633 (N_2633,N_2589,N_2586);
nor U2634 (N_2634,N_2571,N_2573);
nand U2635 (N_2635,N_2513,N_2535);
or U2636 (N_2636,N_2576,N_2566);
nor U2637 (N_2637,N_2543,N_2512);
nand U2638 (N_2638,N_2514,N_2588);
or U2639 (N_2639,N_2580,N_2501);
and U2640 (N_2640,N_2546,N_2558);
or U2641 (N_2641,N_2528,N_2553);
nand U2642 (N_2642,N_2595,N_2562);
nor U2643 (N_2643,N_2587,N_2557);
and U2644 (N_2644,N_2568,N_2536);
or U2645 (N_2645,N_2561,N_2585);
nand U2646 (N_2646,N_2583,N_2516);
and U2647 (N_2647,N_2551,N_2527);
or U2648 (N_2648,N_2563,N_2550);
nand U2649 (N_2649,N_2567,N_2598);
and U2650 (N_2650,N_2555,N_2508);
and U2651 (N_2651,N_2558,N_2503);
nor U2652 (N_2652,N_2529,N_2596);
nor U2653 (N_2653,N_2531,N_2529);
and U2654 (N_2654,N_2586,N_2500);
nand U2655 (N_2655,N_2553,N_2583);
or U2656 (N_2656,N_2534,N_2540);
nor U2657 (N_2657,N_2513,N_2537);
or U2658 (N_2658,N_2557,N_2558);
nand U2659 (N_2659,N_2545,N_2569);
or U2660 (N_2660,N_2559,N_2590);
nor U2661 (N_2661,N_2509,N_2534);
and U2662 (N_2662,N_2595,N_2596);
nand U2663 (N_2663,N_2511,N_2585);
and U2664 (N_2664,N_2597,N_2500);
nor U2665 (N_2665,N_2514,N_2567);
nand U2666 (N_2666,N_2556,N_2546);
or U2667 (N_2667,N_2561,N_2531);
and U2668 (N_2668,N_2596,N_2585);
or U2669 (N_2669,N_2589,N_2541);
nand U2670 (N_2670,N_2537,N_2583);
nor U2671 (N_2671,N_2554,N_2578);
nand U2672 (N_2672,N_2524,N_2581);
and U2673 (N_2673,N_2502,N_2504);
or U2674 (N_2674,N_2541,N_2579);
or U2675 (N_2675,N_2566,N_2589);
and U2676 (N_2676,N_2503,N_2525);
or U2677 (N_2677,N_2598,N_2538);
or U2678 (N_2678,N_2549,N_2531);
and U2679 (N_2679,N_2552,N_2502);
nand U2680 (N_2680,N_2597,N_2513);
or U2681 (N_2681,N_2544,N_2540);
and U2682 (N_2682,N_2515,N_2571);
or U2683 (N_2683,N_2551,N_2566);
and U2684 (N_2684,N_2550,N_2519);
nor U2685 (N_2685,N_2519,N_2585);
nor U2686 (N_2686,N_2515,N_2548);
nor U2687 (N_2687,N_2524,N_2541);
or U2688 (N_2688,N_2578,N_2566);
nor U2689 (N_2689,N_2511,N_2574);
nor U2690 (N_2690,N_2503,N_2597);
or U2691 (N_2691,N_2580,N_2550);
nor U2692 (N_2692,N_2547,N_2560);
nand U2693 (N_2693,N_2528,N_2511);
nor U2694 (N_2694,N_2564,N_2527);
or U2695 (N_2695,N_2591,N_2521);
xnor U2696 (N_2696,N_2541,N_2506);
nand U2697 (N_2697,N_2506,N_2546);
and U2698 (N_2698,N_2597,N_2587);
or U2699 (N_2699,N_2562,N_2569);
nor U2700 (N_2700,N_2673,N_2656);
nor U2701 (N_2701,N_2628,N_2691);
and U2702 (N_2702,N_2668,N_2614);
nand U2703 (N_2703,N_2616,N_2658);
and U2704 (N_2704,N_2625,N_2686);
and U2705 (N_2705,N_2603,N_2694);
nor U2706 (N_2706,N_2698,N_2605);
or U2707 (N_2707,N_2657,N_2695);
and U2708 (N_2708,N_2693,N_2647);
or U2709 (N_2709,N_2672,N_2635);
or U2710 (N_2710,N_2680,N_2654);
nor U2711 (N_2711,N_2643,N_2671);
or U2712 (N_2712,N_2630,N_2662);
nor U2713 (N_2713,N_2642,N_2663);
or U2714 (N_2714,N_2632,N_2624);
or U2715 (N_2715,N_2627,N_2638);
nor U2716 (N_2716,N_2622,N_2633);
nor U2717 (N_2717,N_2689,N_2655);
and U2718 (N_2718,N_2629,N_2634);
nand U2719 (N_2719,N_2651,N_2631);
nand U2720 (N_2720,N_2697,N_2612);
and U2721 (N_2721,N_2692,N_2652);
xor U2722 (N_2722,N_2676,N_2661);
or U2723 (N_2723,N_2608,N_2636);
nand U2724 (N_2724,N_2682,N_2675);
and U2725 (N_2725,N_2665,N_2641);
nor U2726 (N_2726,N_2621,N_2650);
or U2727 (N_2727,N_2681,N_2610);
nor U2728 (N_2728,N_2602,N_2670);
and U2729 (N_2729,N_2617,N_2639);
and U2730 (N_2730,N_2677,N_2645);
or U2731 (N_2731,N_2601,N_2688);
nor U2732 (N_2732,N_2646,N_2678);
nand U2733 (N_2733,N_2685,N_2637);
nand U2734 (N_2734,N_2619,N_2623);
nand U2735 (N_2735,N_2611,N_2644);
nand U2736 (N_2736,N_2600,N_2667);
and U2737 (N_2737,N_2613,N_2609);
nand U2738 (N_2738,N_2687,N_2648);
and U2739 (N_2739,N_2607,N_2684);
and U2740 (N_2740,N_2683,N_2696);
nand U2741 (N_2741,N_2659,N_2679);
nor U2742 (N_2742,N_2653,N_2615);
nand U2743 (N_2743,N_2664,N_2666);
nand U2744 (N_2744,N_2618,N_2674);
nor U2745 (N_2745,N_2606,N_2690);
and U2746 (N_2746,N_2699,N_2640);
or U2747 (N_2747,N_2649,N_2626);
or U2748 (N_2748,N_2660,N_2604);
and U2749 (N_2749,N_2620,N_2669);
nand U2750 (N_2750,N_2666,N_2640);
or U2751 (N_2751,N_2643,N_2661);
xor U2752 (N_2752,N_2666,N_2613);
and U2753 (N_2753,N_2690,N_2626);
or U2754 (N_2754,N_2632,N_2677);
and U2755 (N_2755,N_2684,N_2609);
nor U2756 (N_2756,N_2629,N_2652);
and U2757 (N_2757,N_2662,N_2679);
or U2758 (N_2758,N_2629,N_2648);
or U2759 (N_2759,N_2668,N_2604);
nor U2760 (N_2760,N_2608,N_2603);
nor U2761 (N_2761,N_2633,N_2615);
or U2762 (N_2762,N_2692,N_2685);
and U2763 (N_2763,N_2626,N_2688);
nand U2764 (N_2764,N_2660,N_2641);
or U2765 (N_2765,N_2656,N_2611);
or U2766 (N_2766,N_2645,N_2628);
nand U2767 (N_2767,N_2699,N_2613);
and U2768 (N_2768,N_2605,N_2609);
nor U2769 (N_2769,N_2683,N_2611);
nand U2770 (N_2770,N_2682,N_2692);
nor U2771 (N_2771,N_2633,N_2629);
and U2772 (N_2772,N_2650,N_2614);
nor U2773 (N_2773,N_2667,N_2692);
nand U2774 (N_2774,N_2605,N_2614);
nor U2775 (N_2775,N_2623,N_2637);
and U2776 (N_2776,N_2692,N_2608);
nand U2777 (N_2777,N_2605,N_2656);
nand U2778 (N_2778,N_2671,N_2642);
and U2779 (N_2779,N_2645,N_2614);
and U2780 (N_2780,N_2612,N_2672);
or U2781 (N_2781,N_2610,N_2669);
or U2782 (N_2782,N_2636,N_2600);
or U2783 (N_2783,N_2680,N_2665);
nand U2784 (N_2784,N_2642,N_2678);
and U2785 (N_2785,N_2612,N_2632);
nand U2786 (N_2786,N_2618,N_2628);
nand U2787 (N_2787,N_2655,N_2662);
or U2788 (N_2788,N_2614,N_2693);
nand U2789 (N_2789,N_2662,N_2699);
and U2790 (N_2790,N_2675,N_2661);
nand U2791 (N_2791,N_2628,N_2621);
and U2792 (N_2792,N_2690,N_2607);
and U2793 (N_2793,N_2603,N_2688);
nor U2794 (N_2794,N_2648,N_2607);
nand U2795 (N_2795,N_2679,N_2621);
and U2796 (N_2796,N_2698,N_2676);
nor U2797 (N_2797,N_2669,N_2639);
nor U2798 (N_2798,N_2652,N_2699);
nand U2799 (N_2799,N_2680,N_2640);
or U2800 (N_2800,N_2768,N_2793);
or U2801 (N_2801,N_2746,N_2778);
nor U2802 (N_2802,N_2710,N_2734);
or U2803 (N_2803,N_2733,N_2716);
nand U2804 (N_2804,N_2706,N_2774);
nor U2805 (N_2805,N_2757,N_2713);
or U2806 (N_2806,N_2766,N_2748);
or U2807 (N_2807,N_2782,N_2705);
and U2808 (N_2808,N_2790,N_2724);
and U2809 (N_2809,N_2781,N_2744);
or U2810 (N_2810,N_2798,N_2747);
or U2811 (N_2811,N_2789,N_2738);
or U2812 (N_2812,N_2785,N_2786);
or U2813 (N_2813,N_2772,N_2714);
or U2814 (N_2814,N_2775,N_2735);
nor U2815 (N_2815,N_2795,N_2721);
nand U2816 (N_2816,N_2730,N_2729);
nand U2817 (N_2817,N_2737,N_2777);
and U2818 (N_2818,N_2756,N_2771);
or U2819 (N_2819,N_2788,N_2723);
and U2820 (N_2820,N_2743,N_2740);
or U2821 (N_2821,N_2722,N_2769);
nor U2822 (N_2822,N_2752,N_2755);
or U2823 (N_2823,N_2712,N_2751);
and U2824 (N_2824,N_2701,N_2763);
and U2825 (N_2825,N_2754,N_2742);
nand U2826 (N_2826,N_2728,N_2796);
or U2827 (N_2827,N_2709,N_2741);
or U2828 (N_2828,N_2779,N_2726);
nor U2829 (N_2829,N_2764,N_2773);
or U2830 (N_2830,N_2765,N_2739);
nand U2831 (N_2831,N_2753,N_2718);
nor U2832 (N_2832,N_2715,N_2792);
and U2833 (N_2833,N_2731,N_2704);
and U2834 (N_2834,N_2791,N_2784);
or U2835 (N_2835,N_2711,N_2708);
and U2836 (N_2836,N_2727,N_2780);
nand U2837 (N_2837,N_2725,N_2749);
and U2838 (N_2838,N_2720,N_2736);
or U2839 (N_2839,N_2783,N_2745);
or U2840 (N_2840,N_2797,N_2707);
and U2841 (N_2841,N_2717,N_2702);
or U2842 (N_2842,N_2770,N_2762);
or U2843 (N_2843,N_2758,N_2794);
nand U2844 (N_2844,N_2799,N_2787);
and U2845 (N_2845,N_2776,N_2750);
nor U2846 (N_2846,N_2759,N_2761);
or U2847 (N_2847,N_2703,N_2760);
or U2848 (N_2848,N_2700,N_2719);
and U2849 (N_2849,N_2767,N_2732);
or U2850 (N_2850,N_2796,N_2750);
nand U2851 (N_2851,N_2730,N_2769);
or U2852 (N_2852,N_2745,N_2786);
nand U2853 (N_2853,N_2744,N_2703);
xor U2854 (N_2854,N_2742,N_2772);
or U2855 (N_2855,N_2776,N_2795);
nor U2856 (N_2856,N_2735,N_2774);
and U2857 (N_2857,N_2738,N_2742);
nand U2858 (N_2858,N_2792,N_2725);
nor U2859 (N_2859,N_2775,N_2705);
or U2860 (N_2860,N_2737,N_2735);
nand U2861 (N_2861,N_2732,N_2720);
and U2862 (N_2862,N_2796,N_2775);
nor U2863 (N_2863,N_2766,N_2736);
nand U2864 (N_2864,N_2784,N_2782);
or U2865 (N_2865,N_2788,N_2730);
nand U2866 (N_2866,N_2716,N_2774);
or U2867 (N_2867,N_2787,N_2776);
and U2868 (N_2868,N_2729,N_2710);
nor U2869 (N_2869,N_2761,N_2730);
or U2870 (N_2870,N_2797,N_2724);
or U2871 (N_2871,N_2735,N_2768);
nand U2872 (N_2872,N_2715,N_2709);
nor U2873 (N_2873,N_2779,N_2704);
or U2874 (N_2874,N_2746,N_2751);
and U2875 (N_2875,N_2757,N_2774);
or U2876 (N_2876,N_2757,N_2746);
and U2877 (N_2877,N_2799,N_2731);
nor U2878 (N_2878,N_2780,N_2753);
or U2879 (N_2879,N_2761,N_2725);
nor U2880 (N_2880,N_2790,N_2708);
nor U2881 (N_2881,N_2732,N_2737);
or U2882 (N_2882,N_2787,N_2739);
nor U2883 (N_2883,N_2796,N_2791);
nor U2884 (N_2884,N_2761,N_2763);
nand U2885 (N_2885,N_2790,N_2705);
or U2886 (N_2886,N_2709,N_2732);
nand U2887 (N_2887,N_2771,N_2798);
and U2888 (N_2888,N_2727,N_2787);
nand U2889 (N_2889,N_2749,N_2760);
nand U2890 (N_2890,N_2789,N_2776);
or U2891 (N_2891,N_2708,N_2760);
nand U2892 (N_2892,N_2768,N_2713);
and U2893 (N_2893,N_2746,N_2735);
nand U2894 (N_2894,N_2707,N_2750);
nor U2895 (N_2895,N_2777,N_2752);
nor U2896 (N_2896,N_2723,N_2746);
or U2897 (N_2897,N_2708,N_2755);
or U2898 (N_2898,N_2733,N_2782);
or U2899 (N_2899,N_2748,N_2768);
or U2900 (N_2900,N_2855,N_2874);
nor U2901 (N_2901,N_2892,N_2867);
or U2902 (N_2902,N_2841,N_2873);
and U2903 (N_2903,N_2898,N_2881);
or U2904 (N_2904,N_2831,N_2857);
and U2905 (N_2905,N_2800,N_2801);
and U2906 (N_2906,N_2828,N_2820);
nand U2907 (N_2907,N_2851,N_2880);
nand U2908 (N_2908,N_2882,N_2824);
nand U2909 (N_2909,N_2884,N_2807);
or U2910 (N_2910,N_2812,N_2823);
and U2911 (N_2911,N_2848,N_2822);
nand U2912 (N_2912,N_2809,N_2891);
or U2913 (N_2913,N_2849,N_2839);
or U2914 (N_2914,N_2886,N_2834);
or U2915 (N_2915,N_2866,N_2803);
nand U2916 (N_2916,N_2846,N_2897);
or U2917 (N_2917,N_2890,N_2810);
and U2918 (N_2918,N_2861,N_2816);
and U2919 (N_2919,N_2832,N_2889);
nor U2920 (N_2920,N_2885,N_2863);
nand U2921 (N_2921,N_2888,N_2872);
nor U2922 (N_2922,N_2856,N_2879);
and U2923 (N_2923,N_2876,N_2843);
or U2924 (N_2924,N_2877,N_2821);
and U2925 (N_2925,N_2847,N_2804);
or U2926 (N_2926,N_2852,N_2826);
nand U2927 (N_2927,N_2887,N_2858);
nor U2928 (N_2928,N_2835,N_2806);
or U2929 (N_2929,N_2811,N_2883);
nand U2930 (N_2930,N_2854,N_2860);
nand U2931 (N_2931,N_2838,N_2825);
or U2932 (N_2932,N_2836,N_2895);
nand U2933 (N_2933,N_2865,N_2894);
nand U2934 (N_2934,N_2837,N_2845);
or U2935 (N_2935,N_2813,N_2868);
or U2936 (N_2936,N_2859,N_2869);
and U2937 (N_2937,N_2896,N_2805);
nand U2938 (N_2938,N_2842,N_2864);
or U2939 (N_2939,N_2850,N_2870);
or U2940 (N_2940,N_2814,N_2802);
and U2941 (N_2941,N_2862,N_2827);
or U2942 (N_2942,N_2871,N_2899);
and U2943 (N_2943,N_2844,N_2819);
nand U2944 (N_2944,N_2878,N_2893);
nand U2945 (N_2945,N_2875,N_2808);
and U2946 (N_2946,N_2817,N_2833);
and U2947 (N_2947,N_2830,N_2840);
nand U2948 (N_2948,N_2829,N_2853);
and U2949 (N_2949,N_2815,N_2818);
and U2950 (N_2950,N_2804,N_2841);
or U2951 (N_2951,N_2874,N_2863);
and U2952 (N_2952,N_2880,N_2803);
nor U2953 (N_2953,N_2893,N_2809);
nand U2954 (N_2954,N_2819,N_2846);
nor U2955 (N_2955,N_2866,N_2885);
nand U2956 (N_2956,N_2860,N_2870);
and U2957 (N_2957,N_2879,N_2819);
nand U2958 (N_2958,N_2833,N_2804);
nand U2959 (N_2959,N_2868,N_2879);
and U2960 (N_2960,N_2813,N_2820);
nor U2961 (N_2961,N_2893,N_2867);
or U2962 (N_2962,N_2886,N_2880);
and U2963 (N_2963,N_2889,N_2838);
nand U2964 (N_2964,N_2842,N_2867);
nand U2965 (N_2965,N_2858,N_2850);
nand U2966 (N_2966,N_2821,N_2891);
nand U2967 (N_2967,N_2874,N_2809);
nand U2968 (N_2968,N_2837,N_2834);
and U2969 (N_2969,N_2866,N_2873);
and U2970 (N_2970,N_2810,N_2858);
nor U2971 (N_2971,N_2875,N_2812);
nand U2972 (N_2972,N_2861,N_2897);
nand U2973 (N_2973,N_2880,N_2857);
and U2974 (N_2974,N_2853,N_2828);
or U2975 (N_2975,N_2843,N_2863);
nand U2976 (N_2976,N_2856,N_2887);
or U2977 (N_2977,N_2875,N_2872);
nor U2978 (N_2978,N_2836,N_2829);
or U2979 (N_2979,N_2837,N_2894);
nand U2980 (N_2980,N_2875,N_2834);
nor U2981 (N_2981,N_2864,N_2839);
or U2982 (N_2982,N_2848,N_2841);
and U2983 (N_2983,N_2802,N_2888);
nand U2984 (N_2984,N_2841,N_2876);
nor U2985 (N_2985,N_2826,N_2853);
nand U2986 (N_2986,N_2813,N_2836);
or U2987 (N_2987,N_2843,N_2848);
nor U2988 (N_2988,N_2843,N_2889);
nand U2989 (N_2989,N_2833,N_2819);
nand U2990 (N_2990,N_2879,N_2837);
nor U2991 (N_2991,N_2878,N_2829);
nand U2992 (N_2992,N_2828,N_2838);
and U2993 (N_2993,N_2866,N_2816);
or U2994 (N_2994,N_2808,N_2842);
and U2995 (N_2995,N_2843,N_2839);
or U2996 (N_2996,N_2871,N_2800);
nand U2997 (N_2997,N_2887,N_2803);
and U2998 (N_2998,N_2848,N_2813);
nor U2999 (N_2999,N_2875,N_2848);
xor U3000 (N_3000,N_2961,N_2995);
nand U3001 (N_3001,N_2932,N_2965);
nand U3002 (N_3002,N_2944,N_2933);
nor U3003 (N_3003,N_2978,N_2927);
nor U3004 (N_3004,N_2900,N_2953);
nand U3005 (N_3005,N_2955,N_2967);
or U3006 (N_3006,N_2983,N_2913);
and U3007 (N_3007,N_2974,N_2909);
nand U3008 (N_3008,N_2972,N_2993);
nor U3009 (N_3009,N_2941,N_2911);
nand U3010 (N_3010,N_2942,N_2916);
and U3011 (N_3011,N_2922,N_2960);
nand U3012 (N_3012,N_2997,N_2976);
and U3013 (N_3013,N_2924,N_2903);
and U3014 (N_3014,N_2986,N_2954);
or U3015 (N_3015,N_2988,N_2969);
or U3016 (N_3016,N_2950,N_2930);
and U3017 (N_3017,N_2977,N_2946);
nand U3018 (N_3018,N_2964,N_2984);
or U3019 (N_3019,N_2994,N_2951);
nor U3020 (N_3020,N_2999,N_2952);
or U3021 (N_3021,N_2996,N_2973);
nor U3022 (N_3022,N_2912,N_2902);
and U3023 (N_3023,N_2938,N_2989);
or U3024 (N_3024,N_2985,N_2963);
or U3025 (N_3025,N_2925,N_2982);
nand U3026 (N_3026,N_2956,N_2905);
nor U3027 (N_3027,N_2923,N_2998);
nand U3028 (N_3028,N_2931,N_2948);
or U3029 (N_3029,N_2962,N_2940);
or U3030 (N_3030,N_2975,N_2980);
nand U3031 (N_3031,N_2908,N_2991);
nor U3032 (N_3032,N_2917,N_2920);
nand U3033 (N_3033,N_2929,N_2958);
nor U3034 (N_3034,N_2981,N_2915);
and U3035 (N_3035,N_2939,N_2918);
or U3036 (N_3036,N_2992,N_2987);
nor U3037 (N_3037,N_2959,N_2926);
and U3038 (N_3038,N_2949,N_2914);
or U3039 (N_3039,N_2945,N_2936);
or U3040 (N_3040,N_2947,N_2901);
and U3041 (N_3041,N_2935,N_2943);
or U3042 (N_3042,N_2990,N_2928);
and U3043 (N_3043,N_2906,N_2971);
nand U3044 (N_3044,N_2919,N_2934);
nand U3045 (N_3045,N_2910,N_2921);
nand U3046 (N_3046,N_2957,N_2979);
and U3047 (N_3047,N_2907,N_2966);
nor U3048 (N_3048,N_2937,N_2904);
nand U3049 (N_3049,N_2968,N_2970);
or U3050 (N_3050,N_2980,N_2983);
nand U3051 (N_3051,N_2975,N_2905);
nor U3052 (N_3052,N_2978,N_2982);
and U3053 (N_3053,N_2925,N_2901);
and U3054 (N_3054,N_2977,N_2950);
nand U3055 (N_3055,N_2948,N_2957);
nor U3056 (N_3056,N_2967,N_2988);
and U3057 (N_3057,N_2938,N_2984);
or U3058 (N_3058,N_2980,N_2966);
or U3059 (N_3059,N_2930,N_2985);
nand U3060 (N_3060,N_2946,N_2911);
nand U3061 (N_3061,N_2914,N_2976);
nor U3062 (N_3062,N_2962,N_2974);
nand U3063 (N_3063,N_2962,N_2994);
and U3064 (N_3064,N_2910,N_2977);
nor U3065 (N_3065,N_2914,N_2992);
nor U3066 (N_3066,N_2984,N_2982);
nand U3067 (N_3067,N_2993,N_2983);
nand U3068 (N_3068,N_2928,N_2977);
nand U3069 (N_3069,N_2973,N_2959);
and U3070 (N_3070,N_2982,N_2926);
nand U3071 (N_3071,N_2900,N_2971);
or U3072 (N_3072,N_2995,N_2976);
nand U3073 (N_3073,N_2901,N_2999);
or U3074 (N_3074,N_2980,N_2969);
and U3075 (N_3075,N_2949,N_2916);
and U3076 (N_3076,N_2970,N_2929);
and U3077 (N_3077,N_2958,N_2942);
or U3078 (N_3078,N_2966,N_2906);
xnor U3079 (N_3079,N_2990,N_2932);
nor U3080 (N_3080,N_2951,N_2976);
nand U3081 (N_3081,N_2915,N_2964);
nor U3082 (N_3082,N_2979,N_2941);
and U3083 (N_3083,N_2995,N_2968);
nand U3084 (N_3084,N_2955,N_2932);
or U3085 (N_3085,N_2955,N_2992);
and U3086 (N_3086,N_2955,N_2920);
or U3087 (N_3087,N_2959,N_2984);
and U3088 (N_3088,N_2962,N_2946);
or U3089 (N_3089,N_2999,N_2921);
nand U3090 (N_3090,N_2941,N_2926);
nand U3091 (N_3091,N_2979,N_2901);
nand U3092 (N_3092,N_2966,N_2956);
or U3093 (N_3093,N_2907,N_2969);
or U3094 (N_3094,N_2986,N_2971);
and U3095 (N_3095,N_2969,N_2912);
and U3096 (N_3096,N_2934,N_2973);
nor U3097 (N_3097,N_2961,N_2913);
nand U3098 (N_3098,N_2949,N_2942);
or U3099 (N_3099,N_2901,N_2932);
or U3100 (N_3100,N_3034,N_3005);
or U3101 (N_3101,N_3013,N_3086);
nand U3102 (N_3102,N_3066,N_3074);
nor U3103 (N_3103,N_3068,N_3004);
nand U3104 (N_3104,N_3098,N_3085);
and U3105 (N_3105,N_3011,N_3076);
nand U3106 (N_3106,N_3019,N_3055);
or U3107 (N_3107,N_3094,N_3042);
and U3108 (N_3108,N_3012,N_3031);
or U3109 (N_3109,N_3099,N_3010);
nand U3110 (N_3110,N_3060,N_3033);
xor U3111 (N_3111,N_3078,N_3093);
nand U3112 (N_3112,N_3038,N_3015);
or U3113 (N_3113,N_3039,N_3067);
nand U3114 (N_3114,N_3045,N_3018);
and U3115 (N_3115,N_3046,N_3023);
nand U3116 (N_3116,N_3024,N_3059);
and U3117 (N_3117,N_3002,N_3030);
or U3118 (N_3118,N_3043,N_3069);
nand U3119 (N_3119,N_3006,N_3063);
or U3120 (N_3120,N_3057,N_3079);
nand U3121 (N_3121,N_3020,N_3083);
or U3122 (N_3122,N_3044,N_3021);
nand U3123 (N_3123,N_3064,N_3029);
nor U3124 (N_3124,N_3014,N_3070);
nand U3125 (N_3125,N_3054,N_3016);
and U3126 (N_3126,N_3095,N_3065);
nand U3127 (N_3127,N_3050,N_3071);
nand U3128 (N_3128,N_3058,N_3062);
and U3129 (N_3129,N_3061,N_3035);
and U3130 (N_3130,N_3049,N_3072);
nor U3131 (N_3131,N_3032,N_3022);
nor U3132 (N_3132,N_3053,N_3082);
nor U3133 (N_3133,N_3056,N_3077);
nand U3134 (N_3134,N_3037,N_3026);
nor U3135 (N_3135,N_3001,N_3040);
or U3136 (N_3136,N_3091,N_3089);
nand U3137 (N_3137,N_3025,N_3047);
nand U3138 (N_3138,N_3097,N_3000);
or U3139 (N_3139,N_3084,N_3096);
or U3140 (N_3140,N_3087,N_3041);
nand U3141 (N_3141,N_3009,N_3027);
nand U3142 (N_3142,N_3028,N_3075);
nor U3143 (N_3143,N_3008,N_3092);
or U3144 (N_3144,N_3052,N_3081);
or U3145 (N_3145,N_3051,N_3003);
or U3146 (N_3146,N_3017,N_3048);
nor U3147 (N_3147,N_3088,N_3090);
and U3148 (N_3148,N_3080,N_3073);
and U3149 (N_3149,N_3036,N_3007);
nand U3150 (N_3150,N_3015,N_3059);
nor U3151 (N_3151,N_3062,N_3077);
and U3152 (N_3152,N_3087,N_3020);
nand U3153 (N_3153,N_3045,N_3076);
and U3154 (N_3154,N_3054,N_3034);
nand U3155 (N_3155,N_3074,N_3057);
nor U3156 (N_3156,N_3082,N_3003);
nand U3157 (N_3157,N_3095,N_3081);
and U3158 (N_3158,N_3020,N_3019);
or U3159 (N_3159,N_3082,N_3058);
or U3160 (N_3160,N_3019,N_3047);
and U3161 (N_3161,N_3069,N_3001);
nor U3162 (N_3162,N_3081,N_3058);
and U3163 (N_3163,N_3001,N_3078);
nor U3164 (N_3164,N_3057,N_3063);
nor U3165 (N_3165,N_3042,N_3085);
and U3166 (N_3166,N_3016,N_3000);
or U3167 (N_3167,N_3014,N_3097);
and U3168 (N_3168,N_3071,N_3090);
or U3169 (N_3169,N_3003,N_3062);
nor U3170 (N_3170,N_3052,N_3062);
nand U3171 (N_3171,N_3023,N_3043);
nand U3172 (N_3172,N_3072,N_3059);
nor U3173 (N_3173,N_3099,N_3023);
nor U3174 (N_3174,N_3092,N_3053);
or U3175 (N_3175,N_3010,N_3026);
and U3176 (N_3176,N_3098,N_3066);
and U3177 (N_3177,N_3091,N_3031);
nand U3178 (N_3178,N_3095,N_3035);
nor U3179 (N_3179,N_3073,N_3056);
or U3180 (N_3180,N_3027,N_3021);
and U3181 (N_3181,N_3009,N_3020);
nand U3182 (N_3182,N_3024,N_3043);
nand U3183 (N_3183,N_3018,N_3008);
or U3184 (N_3184,N_3027,N_3006);
and U3185 (N_3185,N_3042,N_3050);
nor U3186 (N_3186,N_3058,N_3017);
nand U3187 (N_3187,N_3087,N_3054);
xor U3188 (N_3188,N_3030,N_3020);
or U3189 (N_3189,N_3074,N_3096);
and U3190 (N_3190,N_3045,N_3043);
and U3191 (N_3191,N_3031,N_3065);
or U3192 (N_3192,N_3035,N_3031);
and U3193 (N_3193,N_3052,N_3013);
and U3194 (N_3194,N_3008,N_3010);
nor U3195 (N_3195,N_3083,N_3044);
nand U3196 (N_3196,N_3088,N_3093);
nand U3197 (N_3197,N_3098,N_3054);
nor U3198 (N_3198,N_3036,N_3004);
nand U3199 (N_3199,N_3001,N_3034);
nor U3200 (N_3200,N_3138,N_3152);
nand U3201 (N_3201,N_3117,N_3125);
nor U3202 (N_3202,N_3180,N_3173);
and U3203 (N_3203,N_3136,N_3153);
or U3204 (N_3204,N_3184,N_3189);
and U3205 (N_3205,N_3120,N_3103);
and U3206 (N_3206,N_3134,N_3116);
nand U3207 (N_3207,N_3150,N_3127);
and U3208 (N_3208,N_3106,N_3176);
nor U3209 (N_3209,N_3161,N_3121);
or U3210 (N_3210,N_3147,N_3157);
nand U3211 (N_3211,N_3118,N_3177);
nor U3212 (N_3212,N_3172,N_3178);
or U3213 (N_3213,N_3114,N_3197);
nor U3214 (N_3214,N_3196,N_3193);
or U3215 (N_3215,N_3139,N_3160);
or U3216 (N_3216,N_3146,N_3145);
xnor U3217 (N_3217,N_3144,N_3175);
nor U3218 (N_3218,N_3123,N_3105);
nand U3219 (N_3219,N_3100,N_3128);
nand U3220 (N_3220,N_3191,N_3170);
nor U3221 (N_3221,N_3101,N_3190);
and U3222 (N_3222,N_3158,N_3129);
or U3223 (N_3223,N_3186,N_3102);
and U3224 (N_3224,N_3142,N_3133);
nor U3225 (N_3225,N_3122,N_3166);
nor U3226 (N_3226,N_3104,N_3135);
and U3227 (N_3227,N_3188,N_3163);
and U3228 (N_3228,N_3115,N_3185);
nand U3229 (N_3229,N_3155,N_3165);
xor U3230 (N_3230,N_3143,N_3167);
and U3231 (N_3231,N_3194,N_3171);
nor U3232 (N_3232,N_3164,N_3109);
or U3233 (N_3233,N_3149,N_3110);
or U3234 (N_3234,N_3169,N_3124);
nand U3235 (N_3235,N_3154,N_3199);
nand U3236 (N_3236,N_3187,N_3198);
nand U3237 (N_3237,N_3126,N_3168);
nor U3238 (N_3238,N_3130,N_3132);
nor U3239 (N_3239,N_3162,N_3108);
or U3240 (N_3240,N_3140,N_3111);
and U3241 (N_3241,N_3107,N_3174);
or U3242 (N_3242,N_3151,N_3141);
and U3243 (N_3243,N_3195,N_3113);
or U3244 (N_3244,N_3159,N_3131);
nand U3245 (N_3245,N_3179,N_3183);
nor U3246 (N_3246,N_3137,N_3192);
or U3247 (N_3247,N_3119,N_3182);
and U3248 (N_3248,N_3112,N_3156);
nor U3249 (N_3249,N_3148,N_3181);
and U3250 (N_3250,N_3163,N_3118);
and U3251 (N_3251,N_3133,N_3110);
nor U3252 (N_3252,N_3162,N_3110);
nor U3253 (N_3253,N_3109,N_3165);
and U3254 (N_3254,N_3191,N_3134);
and U3255 (N_3255,N_3147,N_3152);
and U3256 (N_3256,N_3156,N_3185);
or U3257 (N_3257,N_3145,N_3175);
nand U3258 (N_3258,N_3114,N_3132);
nand U3259 (N_3259,N_3177,N_3100);
and U3260 (N_3260,N_3196,N_3136);
and U3261 (N_3261,N_3161,N_3154);
or U3262 (N_3262,N_3133,N_3107);
and U3263 (N_3263,N_3185,N_3124);
nor U3264 (N_3264,N_3187,N_3190);
or U3265 (N_3265,N_3154,N_3140);
or U3266 (N_3266,N_3149,N_3101);
and U3267 (N_3267,N_3174,N_3122);
or U3268 (N_3268,N_3125,N_3134);
and U3269 (N_3269,N_3176,N_3180);
or U3270 (N_3270,N_3126,N_3195);
nor U3271 (N_3271,N_3131,N_3147);
nor U3272 (N_3272,N_3143,N_3125);
nor U3273 (N_3273,N_3163,N_3126);
nand U3274 (N_3274,N_3178,N_3141);
nand U3275 (N_3275,N_3179,N_3156);
or U3276 (N_3276,N_3181,N_3173);
nand U3277 (N_3277,N_3105,N_3109);
or U3278 (N_3278,N_3109,N_3108);
and U3279 (N_3279,N_3105,N_3107);
nor U3280 (N_3280,N_3199,N_3156);
nand U3281 (N_3281,N_3138,N_3158);
and U3282 (N_3282,N_3190,N_3164);
xnor U3283 (N_3283,N_3112,N_3129);
nor U3284 (N_3284,N_3167,N_3151);
nand U3285 (N_3285,N_3168,N_3198);
nor U3286 (N_3286,N_3195,N_3144);
nand U3287 (N_3287,N_3161,N_3173);
nand U3288 (N_3288,N_3197,N_3133);
nor U3289 (N_3289,N_3150,N_3185);
nand U3290 (N_3290,N_3106,N_3199);
nand U3291 (N_3291,N_3113,N_3142);
or U3292 (N_3292,N_3159,N_3116);
nor U3293 (N_3293,N_3118,N_3120);
and U3294 (N_3294,N_3194,N_3114);
or U3295 (N_3295,N_3171,N_3188);
nor U3296 (N_3296,N_3192,N_3151);
nand U3297 (N_3297,N_3143,N_3183);
or U3298 (N_3298,N_3128,N_3162);
or U3299 (N_3299,N_3162,N_3132);
and U3300 (N_3300,N_3254,N_3237);
nand U3301 (N_3301,N_3200,N_3243);
nand U3302 (N_3302,N_3290,N_3259);
and U3303 (N_3303,N_3224,N_3249);
nand U3304 (N_3304,N_3280,N_3268);
nand U3305 (N_3305,N_3281,N_3272);
or U3306 (N_3306,N_3239,N_3267);
or U3307 (N_3307,N_3291,N_3212);
and U3308 (N_3308,N_3238,N_3274);
and U3309 (N_3309,N_3270,N_3222);
nand U3310 (N_3310,N_3248,N_3256);
or U3311 (N_3311,N_3209,N_3247);
or U3312 (N_3312,N_3282,N_3217);
and U3313 (N_3313,N_3206,N_3275);
or U3314 (N_3314,N_3246,N_3271);
and U3315 (N_3315,N_3225,N_3263);
nand U3316 (N_3316,N_3219,N_3210);
or U3317 (N_3317,N_3295,N_3203);
or U3318 (N_3318,N_3218,N_3264);
and U3319 (N_3319,N_3273,N_3227);
or U3320 (N_3320,N_3229,N_3296);
or U3321 (N_3321,N_3231,N_3284);
nor U3322 (N_3322,N_3255,N_3214);
nor U3323 (N_3323,N_3278,N_3265);
or U3324 (N_3324,N_3204,N_3208);
nor U3325 (N_3325,N_3213,N_3201);
or U3326 (N_3326,N_3245,N_3244);
nand U3327 (N_3327,N_3223,N_3215);
or U3328 (N_3328,N_3207,N_3252);
or U3329 (N_3329,N_3298,N_3286);
or U3330 (N_3330,N_3294,N_3220);
or U3331 (N_3331,N_3299,N_3289);
nand U3332 (N_3332,N_3240,N_3283);
nand U3333 (N_3333,N_3234,N_3293);
nand U3334 (N_3334,N_3262,N_3230);
nor U3335 (N_3335,N_3276,N_3288);
nor U3336 (N_3336,N_3253,N_3285);
or U3337 (N_3337,N_3251,N_3287);
nor U3338 (N_3338,N_3261,N_3258);
nor U3339 (N_3339,N_3242,N_3277);
or U3340 (N_3340,N_3233,N_3216);
nor U3341 (N_3341,N_3235,N_3297);
nor U3342 (N_3342,N_3236,N_3257);
or U3343 (N_3343,N_3221,N_3226);
nand U3344 (N_3344,N_3241,N_3211);
or U3345 (N_3345,N_3260,N_3202);
nand U3346 (N_3346,N_3266,N_3232);
nand U3347 (N_3347,N_3250,N_3292);
nand U3348 (N_3348,N_3205,N_3279);
nor U3349 (N_3349,N_3269,N_3228);
or U3350 (N_3350,N_3271,N_3214);
or U3351 (N_3351,N_3222,N_3205);
nand U3352 (N_3352,N_3246,N_3249);
and U3353 (N_3353,N_3248,N_3241);
and U3354 (N_3354,N_3221,N_3253);
and U3355 (N_3355,N_3279,N_3270);
nor U3356 (N_3356,N_3260,N_3290);
nand U3357 (N_3357,N_3289,N_3215);
nor U3358 (N_3358,N_3247,N_3213);
and U3359 (N_3359,N_3210,N_3294);
or U3360 (N_3360,N_3270,N_3248);
and U3361 (N_3361,N_3204,N_3238);
nor U3362 (N_3362,N_3241,N_3247);
and U3363 (N_3363,N_3287,N_3289);
nand U3364 (N_3364,N_3202,N_3266);
or U3365 (N_3365,N_3296,N_3258);
or U3366 (N_3366,N_3259,N_3210);
nor U3367 (N_3367,N_3281,N_3229);
or U3368 (N_3368,N_3251,N_3231);
and U3369 (N_3369,N_3267,N_3278);
and U3370 (N_3370,N_3289,N_3231);
nand U3371 (N_3371,N_3244,N_3229);
nor U3372 (N_3372,N_3256,N_3217);
nor U3373 (N_3373,N_3218,N_3288);
and U3374 (N_3374,N_3208,N_3246);
nand U3375 (N_3375,N_3282,N_3229);
nand U3376 (N_3376,N_3256,N_3291);
nand U3377 (N_3377,N_3247,N_3264);
nand U3378 (N_3378,N_3291,N_3273);
or U3379 (N_3379,N_3260,N_3255);
and U3380 (N_3380,N_3216,N_3275);
and U3381 (N_3381,N_3204,N_3207);
and U3382 (N_3382,N_3228,N_3244);
or U3383 (N_3383,N_3257,N_3242);
nand U3384 (N_3384,N_3239,N_3249);
or U3385 (N_3385,N_3230,N_3226);
nand U3386 (N_3386,N_3285,N_3272);
or U3387 (N_3387,N_3282,N_3259);
and U3388 (N_3388,N_3283,N_3218);
nand U3389 (N_3389,N_3267,N_3210);
nand U3390 (N_3390,N_3257,N_3239);
nor U3391 (N_3391,N_3214,N_3228);
nand U3392 (N_3392,N_3232,N_3200);
or U3393 (N_3393,N_3298,N_3221);
nand U3394 (N_3394,N_3222,N_3223);
xor U3395 (N_3395,N_3229,N_3264);
nor U3396 (N_3396,N_3295,N_3241);
and U3397 (N_3397,N_3231,N_3227);
and U3398 (N_3398,N_3243,N_3250);
nor U3399 (N_3399,N_3246,N_3205);
nand U3400 (N_3400,N_3358,N_3378);
and U3401 (N_3401,N_3368,N_3305);
or U3402 (N_3402,N_3392,N_3387);
nor U3403 (N_3403,N_3383,N_3343);
or U3404 (N_3404,N_3374,N_3382);
and U3405 (N_3405,N_3316,N_3340);
nor U3406 (N_3406,N_3385,N_3350);
and U3407 (N_3407,N_3345,N_3328);
and U3408 (N_3408,N_3335,N_3363);
nor U3409 (N_3409,N_3307,N_3362);
nand U3410 (N_3410,N_3331,N_3320);
nor U3411 (N_3411,N_3390,N_3351);
and U3412 (N_3412,N_3356,N_3309);
and U3413 (N_3413,N_3377,N_3315);
or U3414 (N_3414,N_3355,N_3376);
nor U3415 (N_3415,N_3318,N_3354);
or U3416 (N_3416,N_3391,N_3344);
and U3417 (N_3417,N_3301,N_3373);
nand U3418 (N_3418,N_3333,N_3346);
nand U3419 (N_3419,N_3394,N_3341);
or U3420 (N_3420,N_3388,N_3325);
nand U3421 (N_3421,N_3338,N_3369);
and U3422 (N_3422,N_3396,N_3398);
and U3423 (N_3423,N_3366,N_3360);
nor U3424 (N_3424,N_3397,N_3399);
and U3425 (N_3425,N_3321,N_3303);
or U3426 (N_3426,N_3319,N_3372);
or U3427 (N_3427,N_3330,N_3389);
or U3428 (N_3428,N_3370,N_3302);
or U3429 (N_3429,N_3314,N_3326);
nor U3430 (N_3430,N_3365,N_3347);
or U3431 (N_3431,N_3312,N_3395);
nor U3432 (N_3432,N_3322,N_3332);
nand U3433 (N_3433,N_3349,N_3381);
and U3434 (N_3434,N_3342,N_3329);
or U3435 (N_3435,N_3323,N_3384);
nor U3436 (N_3436,N_3337,N_3334);
and U3437 (N_3437,N_3304,N_3380);
nand U3438 (N_3438,N_3300,N_3313);
nor U3439 (N_3439,N_3367,N_3359);
nand U3440 (N_3440,N_3352,N_3306);
nor U3441 (N_3441,N_3375,N_3364);
nand U3442 (N_3442,N_3327,N_3308);
nand U3443 (N_3443,N_3310,N_3386);
nor U3444 (N_3444,N_3353,N_3348);
nor U3445 (N_3445,N_3339,N_3379);
nand U3446 (N_3446,N_3317,N_3357);
nor U3447 (N_3447,N_3324,N_3371);
nor U3448 (N_3448,N_3336,N_3361);
nor U3449 (N_3449,N_3393,N_3311);
nand U3450 (N_3450,N_3386,N_3335);
nor U3451 (N_3451,N_3390,N_3310);
nor U3452 (N_3452,N_3312,N_3316);
and U3453 (N_3453,N_3392,N_3314);
nor U3454 (N_3454,N_3378,N_3362);
and U3455 (N_3455,N_3302,N_3335);
nor U3456 (N_3456,N_3307,N_3327);
and U3457 (N_3457,N_3347,N_3303);
nor U3458 (N_3458,N_3378,N_3328);
or U3459 (N_3459,N_3352,N_3387);
or U3460 (N_3460,N_3331,N_3374);
nand U3461 (N_3461,N_3380,N_3301);
nor U3462 (N_3462,N_3300,N_3302);
or U3463 (N_3463,N_3395,N_3382);
nor U3464 (N_3464,N_3380,N_3308);
nor U3465 (N_3465,N_3387,N_3358);
xnor U3466 (N_3466,N_3333,N_3398);
nand U3467 (N_3467,N_3355,N_3330);
nand U3468 (N_3468,N_3371,N_3306);
nand U3469 (N_3469,N_3387,N_3340);
nor U3470 (N_3470,N_3366,N_3386);
or U3471 (N_3471,N_3339,N_3373);
nand U3472 (N_3472,N_3339,N_3380);
nand U3473 (N_3473,N_3397,N_3300);
or U3474 (N_3474,N_3364,N_3395);
or U3475 (N_3475,N_3390,N_3345);
or U3476 (N_3476,N_3356,N_3373);
and U3477 (N_3477,N_3380,N_3376);
nand U3478 (N_3478,N_3356,N_3371);
and U3479 (N_3479,N_3320,N_3311);
and U3480 (N_3480,N_3343,N_3344);
nor U3481 (N_3481,N_3347,N_3372);
nand U3482 (N_3482,N_3333,N_3312);
and U3483 (N_3483,N_3386,N_3340);
and U3484 (N_3484,N_3314,N_3391);
and U3485 (N_3485,N_3323,N_3379);
or U3486 (N_3486,N_3387,N_3330);
nor U3487 (N_3487,N_3313,N_3341);
or U3488 (N_3488,N_3390,N_3301);
and U3489 (N_3489,N_3367,N_3313);
and U3490 (N_3490,N_3345,N_3342);
nor U3491 (N_3491,N_3342,N_3307);
nor U3492 (N_3492,N_3395,N_3372);
nor U3493 (N_3493,N_3351,N_3352);
and U3494 (N_3494,N_3307,N_3393);
and U3495 (N_3495,N_3380,N_3309);
or U3496 (N_3496,N_3328,N_3386);
nand U3497 (N_3497,N_3308,N_3314);
nand U3498 (N_3498,N_3309,N_3332);
or U3499 (N_3499,N_3303,N_3311);
or U3500 (N_3500,N_3489,N_3408);
and U3501 (N_3501,N_3417,N_3420);
nor U3502 (N_3502,N_3481,N_3453);
nand U3503 (N_3503,N_3442,N_3452);
nand U3504 (N_3504,N_3477,N_3409);
or U3505 (N_3505,N_3414,N_3410);
nand U3506 (N_3506,N_3493,N_3441);
or U3507 (N_3507,N_3475,N_3439);
and U3508 (N_3508,N_3478,N_3425);
or U3509 (N_3509,N_3415,N_3461);
and U3510 (N_3510,N_3451,N_3492);
nor U3511 (N_3511,N_3440,N_3449);
nor U3512 (N_3512,N_3497,N_3406);
or U3513 (N_3513,N_3433,N_3476);
or U3514 (N_3514,N_3418,N_3459);
nand U3515 (N_3515,N_3494,N_3443);
or U3516 (N_3516,N_3486,N_3404);
nor U3517 (N_3517,N_3436,N_3483);
nand U3518 (N_3518,N_3469,N_3479);
nor U3519 (N_3519,N_3407,N_3456);
nand U3520 (N_3520,N_3444,N_3402);
or U3521 (N_3521,N_3472,N_3465);
and U3522 (N_3522,N_3445,N_3467);
nor U3523 (N_3523,N_3499,N_3419);
nand U3524 (N_3524,N_3470,N_3413);
or U3525 (N_3525,N_3498,N_3460);
nand U3526 (N_3526,N_3482,N_3448);
nand U3527 (N_3527,N_3463,N_3428);
nor U3528 (N_3528,N_3487,N_3496);
or U3529 (N_3529,N_3454,N_3416);
or U3530 (N_3530,N_3430,N_3466);
or U3531 (N_3531,N_3495,N_3403);
or U3532 (N_3532,N_3429,N_3423);
or U3533 (N_3533,N_3484,N_3491);
and U3534 (N_3534,N_3488,N_3411);
or U3535 (N_3535,N_3450,N_3474);
or U3536 (N_3536,N_3455,N_3412);
nor U3537 (N_3537,N_3434,N_3485);
nor U3538 (N_3538,N_3421,N_3401);
and U3539 (N_3539,N_3473,N_3405);
nor U3540 (N_3540,N_3446,N_3424);
nor U3541 (N_3541,N_3464,N_3426);
nor U3542 (N_3542,N_3422,N_3447);
or U3543 (N_3543,N_3400,N_3471);
nor U3544 (N_3544,N_3438,N_3427);
and U3545 (N_3545,N_3432,N_3437);
nand U3546 (N_3546,N_3490,N_3458);
nand U3547 (N_3547,N_3431,N_3480);
nor U3548 (N_3548,N_3462,N_3435);
xnor U3549 (N_3549,N_3457,N_3468);
nor U3550 (N_3550,N_3463,N_3417);
or U3551 (N_3551,N_3477,N_3406);
nand U3552 (N_3552,N_3457,N_3491);
nor U3553 (N_3553,N_3488,N_3434);
nand U3554 (N_3554,N_3403,N_3481);
or U3555 (N_3555,N_3481,N_3462);
or U3556 (N_3556,N_3493,N_3492);
or U3557 (N_3557,N_3456,N_3418);
or U3558 (N_3558,N_3419,N_3433);
nor U3559 (N_3559,N_3429,N_3499);
nor U3560 (N_3560,N_3401,N_3407);
and U3561 (N_3561,N_3446,N_3451);
or U3562 (N_3562,N_3413,N_3473);
nand U3563 (N_3563,N_3495,N_3447);
nor U3564 (N_3564,N_3476,N_3419);
nand U3565 (N_3565,N_3443,N_3424);
nor U3566 (N_3566,N_3455,N_3408);
and U3567 (N_3567,N_3403,N_3433);
nand U3568 (N_3568,N_3488,N_3485);
and U3569 (N_3569,N_3499,N_3435);
nand U3570 (N_3570,N_3434,N_3476);
or U3571 (N_3571,N_3454,N_3407);
nand U3572 (N_3572,N_3444,N_3419);
nand U3573 (N_3573,N_3439,N_3413);
xnor U3574 (N_3574,N_3459,N_3405);
or U3575 (N_3575,N_3420,N_3458);
nand U3576 (N_3576,N_3406,N_3496);
or U3577 (N_3577,N_3483,N_3435);
or U3578 (N_3578,N_3444,N_3407);
or U3579 (N_3579,N_3441,N_3420);
or U3580 (N_3580,N_3409,N_3418);
nand U3581 (N_3581,N_3471,N_3443);
nand U3582 (N_3582,N_3410,N_3452);
nor U3583 (N_3583,N_3406,N_3433);
nor U3584 (N_3584,N_3477,N_3481);
nor U3585 (N_3585,N_3447,N_3451);
and U3586 (N_3586,N_3452,N_3496);
nor U3587 (N_3587,N_3439,N_3468);
or U3588 (N_3588,N_3468,N_3428);
and U3589 (N_3589,N_3498,N_3413);
and U3590 (N_3590,N_3456,N_3419);
nand U3591 (N_3591,N_3403,N_3490);
or U3592 (N_3592,N_3491,N_3414);
or U3593 (N_3593,N_3426,N_3445);
or U3594 (N_3594,N_3451,N_3474);
and U3595 (N_3595,N_3427,N_3402);
and U3596 (N_3596,N_3408,N_3412);
and U3597 (N_3597,N_3459,N_3472);
nand U3598 (N_3598,N_3461,N_3454);
nor U3599 (N_3599,N_3429,N_3468);
nor U3600 (N_3600,N_3523,N_3537);
nor U3601 (N_3601,N_3574,N_3563);
and U3602 (N_3602,N_3578,N_3550);
nand U3603 (N_3603,N_3579,N_3510);
nor U3604 (N_3604,N_3532,N_3519);
nand U3605 (N_3605,N_3561,N_3595);
nor U3606 (N_3606,N_3572,N_3560);
or U3607 (N_3607,N_3546,N_3525);
nor U3608 (N_3608,N_3568,N_3514);
and U3609 (N_3609,N_3590,N_3538);
or U3610 (N_3610,N_3554,N_3599);
xnor U3611 (N_3611,N_3577,N_3556);
nand U3612 (N_3612,N_3586,N_3508);
nand U3613 (N_3613,N_3503,N_3516);
and U3614 (N_3614,N_3582,N_3583);
nor U3615 (N_3615,N_3594,N_3593);
nand U3616 (N_3616,N_3526,N_3536);
nor U3617 (N_3617,N_3559,N_3562);
nand U3618 (N_3618,N_3543,N_3547);
and U3619 (N_3619,N_3545,N_3581);
or U3620 (N_3620,N_3597,N_3548);
nand U3621 (N_3621,N_3587,N_3544);
nand U3622 (N_3622,N_3501,N_3517);
and U3623 (N_3623,N_3535,N_3521);
nor U3624 (N_3624,N_3551,N_3592);
or U3625 (N_3625,N_3540,N_3558);
or U3626 (N_3626,N_3552,N_3515);
or U3627 (N_3627,N_3570,N_3585);
nand U3628 (N_3628,N_3530,N_3541);
or U3629 (N_3629,N_3512,N_3507);
nor U3630 (N_3630,N_3518,N_3520);
or U3631 (N_3631,N_3505,N_3534);
or U3632 (N_3632,N_3500,N_3513);
nand U3633 (N_3633,N_3566,N_3549);
and U3634 (N_3634,N_3567,N_3504);
nand U3635 (N_3635,N_3531,N_3527);
nand U3636 (N_3636,N_3596,N_3509);
nor U3637 (N_3637,N_3529,N_3557);
or U3638 (N_3638,N_3598,N_3506);
or U3639 (N_3639,N_3576,N_3571);
nor U3640 (N_3640,N_3589,N_3588);
and U3641 (N_3641,N_3533,N_3580);
nor U3642 (N_3642,N_3575,N_3555);
and U3643 (N_3643,N_3528,N_3591);
and U3644 (N_3644,N_3565,N_3553);
and U3645 (N_3645,N_3502,N_3542);
nor U3646 (N_3646,N_3573,N_3564);
or U3647 (N_3647,N_3524,N_3569);
or U3648 (N_3648,N_3584,N_3522);
nand U3649 (N_3649,N_3539,N_3511);
or U3650 (N_3650,N_3524,N_3550);
and U3651 (N_3651,N_3548,N_3598);
and U3652 (N_3652,N_3576,N_3588);
nand U3653 (N_3653,N_3512,N_3599);
or U3654 (N_3654,N_3533,N_3555);
and U3655 (N_3655,N_3545,N_3507);
or U3656 (N_3656,N_3573,N_3596);
nor U3657 (N_3657,N_3579,N_3553);
nand U3658 (N_3658,N_3522,N_3541);
and U3659 (N_3659,N_3559,N_3569);
or U3660 (N_3660,N_3524,N_3566);
nor U3661 (N_3661,N_3530,N_3543);
nor U3662 (N_3662,N_3536,N_3523);
and U3663 (N_3663,N_3508,N_3552);
nor U3664 (N_3664,N_3573,N_3558);
nand U3665 (N_3665,N_3556,N_3512);
and U3666 (N_3666,N_3503,N_3563);
and U3667 (N_3667,N_3521,N_3548);
nor U3668 (N_3668,N_3537,N_3575);
and U3669 (N_3669,N_3520,N_3547);
nand U3670 (N_3670,N_3547,N_3556);
or U3671 (N_3671,N_3584,N_3579);
or U3672 (N_3672,N_3579,N_3508);
nor U3673 (N_3673,N_3567,N_3512);
nor U3674 (N_3674,N_3575,N_3598);
or U3675 (N_3675,N_3572,N_3500);
and U3676 (N_3676,N_3519,N_3571);
or U3677 (N_3677,N_3578,N_3565);
and U3678 (N_3678,N_3526,N_3565);
or U3679 (N_3679,N_3509,N_3541);
nor U3680 (N_3680,N_3560,N_3503);
or U3681 (N_3681,N_3512,N_3536);
nand U3682 (N_3682,N_3546,N_3588);
nand U3683 (N_3683,N_3581,N_3522);
and U3684 (N_3684,N_3533,N_3514);
and U3685 (N_3685,N_3513,N_3535);
nand U3686 (N_3686,N_3539,N_3581);
or U3687 (N_3687,N_3533,N_3553);
and U3688 (N_3688,N_3581,N_3537);
or U3689 (N_3689,N_3571,N_3589);
and U3690 (N_3690,N_3589,N_3509);
nor U3691 (N_3691,N_3549,N_3552);
or U3692 (N_3692,N_3581,N_3513);
nor U3693 (N_3693,N_3578,N_3586);
nand U3694 (N_3694,N_3532,N_3549);
nand U3695 (N_3695,N_3597,N_3525);
or U3696 (N_3696,N_3512,N_3550);
and U3697 (N_3697,N_3516,N_3589);
nor U3698 (N_3698,N_3524,N_3548);
nand U3699 (N_3699,N_3582,N_3570);
nor U3700 (N_3700,N_3645,N_3688);
nand U3701 (N_3701,N_3671,N_3646);
and U3702 (N_3702,N_3693,N_3629);
nand U3703 (N_3703,N_3638,N_3689);
nand U3704 (N_3704,N_3642,N_3618);
nor U3705 (N_3705,N_3648,N_3686);
and U3706 (N_3706,N_3613,N_3655);
nor U3707 (N_3707,N_3600,N_3603);
or U3708 (N_3708,N_3609,N_3652);
and U3709 (N_3709,N_3679,N_3683);
or U3710 (N_3710,N_3614,N_3665);
nand U3711 (N_3711,N_3658,N_3624);
or U3712 (N_3712,N_3611,N_3685);
and U3713 (N_3713,N_3699,N_3634);
nor U3714 (N_3714,N_3656,N_3695);
nand U3715 (N_3715,N_3664,N_3670);
and U3716 (N_3716,N_3615,N_3650);
nand U3717 (N_3717,N_3625,N_3639);
or U3718 (N_3718,N_3607,N_3660);
nor U3719 (N_3719,N_3631,N_3636);
nor U3720 (N_3720,N_3681,N_3617);
nor U3721 (N_3721,N_3675,N_3677);
nand U3722 (N_3722,N_3654,N_3657);
or U3723 (N_3723,N_3649,N_3626);
nand U3724 (N_3724,N_3651,N_3643);
and U3725 (N_3725,N_3687,N_3667);
and U3726 (N_3726,N_3659,N_3640);
and U3727 (N_3727,N_3672,N_3663);
nor U3728 (N_3728,N_3608,N_3682);
or U3729 (N_3729,N_3661,N_3633);
or U3730 (N_3730,N_3684,N_3630);
or U3731 (N_3731,N_3662,N_3653);
nor U3732 (N_3732,N_3698,N_3666);
or U3733 (N_3733,N_3604,N_3623);
and U3734 (N_3734,N_3669,N_3612);
and U3735 (N_3735,N_3637,N_3647);
nand U3736 (N_3736,N_3619,N_3602);
or U3737 (N_3737,N_3691,N_3641);
nand U3738 (N_3738,N_3605,N_3610);
or U3739 (N_3739,N_3644,N_3635);
or U3740 (N_3740,N_3680,N_3616);
and U3741 (N_3741,N_3694,N_3676);
or U3742 (N_3742,N_3621,N_3601);
nand U3743 (N_3743,N_3620,N_3606);
and U3744 (N_3744,N_3628,N_3673);
or U3745 (N_3745,N_3692,N_3697);
nor U3746 (N_3746,N_3622,N_3627);
nor U3747 (N_3747,N_3678,N_3632);
nor U3748 (N_3748,N_3696,N_3690);
nor U3749 (N_3749,N_3668,N_3674);
or U3750 (N_3750,N_3696,N_3647);
nand U3751 (N_3751,N_3631,N_3648);
nor U3752 (N_3752,N_3606,N_3607);
and U3753 (N_3753,N_3679,N_3632);
nor U3754 (N_3754,N_3676,N_3639);
nand U3755 (N_3755,N_3621,N_3636);
and U3756 (N_3756,N_3665,N_3624);
nand U3757 (N_3757,N_3628,N_3661);
and U3758 (N_3758,N_3689,N_3678);
nand U3759 (N_3759,N_3683,N_3670);
nand U3760 (N_3760,N_3646,N_3697);
and U3761 (N_3761,N_3669,N_3618);
and U3762 (N_3762,N_3663,N_3611);
and U3763 (N_3763,N_3678,N_3663);
nor U3764 (N_3764,N_3647,N_3602);
and U3765 (N_3765,N_3681,N_3620);
and U3766 (N_3766,N_3642,N_3613);
nand U3767 (N_3767,N_3679,N_3649);
or U3768 (N_3768,N_3605,N_3666);
and U3769 (N_3769,N_3641,N_3648);
nand U3770 (N_3770,N_3694,N_3668);
nor U3771 (N_3771,N_3654,N_3692);
or U3772 (N_3772,N_3678,N_3668);
nand U3773 (N_3773,N_3674,N_3691);
or U3774 (N_3774,N_3652,N_3630);
nor U3775 (N_3775,N_3692,N_3620);
nor U3776 (N_3776,N_3642,N_3696);
nand U3777 (N_3777,N_3660,N_3649);
nand U3778 (N_3778,N_3607,N_3619);
and U3779 (N_3779,N_3659,N_3631);
nand U3780 (N_3780,N_3620,N_3693);
nand U3781 (N_3781,N_3625,N_3693);
or U3782 (N_3782,N_3627,N_3602);
nand U3783 (N_3783,N_3681,N_3676);
or U3784 (N_3784,N_3667,N_3693);
or U3785 (N_3785,N_3623,N_3695);
nor U3786 (N_3786,N_3650,N_3610);
or U3787 (N_3787,N_3653,N_3605);
and U3788 (N_3788,N_3609,N_3658);
and U3789 (N_3789,N_3618,N_3628);
or U3790 (N_3790,N_3673,N_3622);
xor U3791 (N_3791,N_3650,N_3673);
nor U3792 (N_3792,N_3696,N_3628);
or U3793 (N_3793,N_3626,N_3601);
nand U3794 (N_3794,N_3619,N_3699);
nand U3795 (N_3795,N_3663,N_3634);
nor U3796 (N_3796,N_3678,N_3669);
or U3797 (N_3797,N_3658,N_3688);
and U3798 (N_3798,N_3686,N_3657);
nand U3799 (N_3799,N_3640,N_3695);
nand U3800 (N_3800,N_3710,N_3729);
nor U3801 (N_3801,N_3789,N_3785);
and U3802 (N_3802,N_3700,N_3754);
and U3803 (N_3803,N_3798,N_3747);
nand U3804 (N_3804,N_3757,N_3712);
or U3805 (N_3805,N_3759,N_3771);
or U3806 (N_3806,N_3704,N_3733);
or U3807 (N_3807,N_3774,N_3701);
nor U3808 (N_3808,N_3781,N_3705);
or U3809 (N_3809,N_3715,N_3752);
nor U3810 (N_3810,N_3763,N_3751);
nor U3811 (N_3811,N_3796,N_3743);
nand U3812 (N_3812,N_3760,N_3740);
nand U3813 (N_3813,N_3790,N_3711);
and U3814 (N_3814,N_3797,N_3703);
nor U3815 (N_3815,N_3719,N_3721);
nand U3816 (N_3816,N_3714,N_3764);
nor U3817 (N_3817,N_3769,N_3748);
and U3818 (N_3818,N_3720,N_3728);
and U3819 (N_3819,N_3723,N_3762);
nand U3820 (N_3820,N_3707,N_3742);
nor U3821 (N_3821,N_3775,N_3745);
nor U3822 (N_3822,N_3734,N_3727);
and U3823 (N_3823,N_3713,N_3792);
or U3824 (N_3824,N_3708,N_3716);
nand U3825 (N_3825,N_3766,N_3791);
and U3826 (N_3826,N_3765,N_3772);
or U3827 (N_3827,N_3722,N_3788);
or U3828 (N_3828,N_3753,N_3709);
or U3829 (N_3829,N_3736,N_3777);
nor U3830 (N_3830,N_3768,N_3718);
or U3831 (N_3831,N_3776,N_3756);
or U3832 (N_3832,N_3724,N_3758);
and U3833 (N_3833,N_3735,N_3778);
nor U3834 (N_3834,N_3755,N_3786);
and U3835 (N_3835,N_3725,N_3702);
nor U3836 (N_3836,N_3773,N_3738);
nor U3837 (N_3837,N_3750,N_3741);
nand U3838 (N_3838,N_3739,N_3737);
or U3839 (N_3839,N_3749,N_3780);
or U3840 (N_3840,N_3793,N_3794);
nand U3841 (N_3841,N_3726,N_3746);
or U3842 (N_3842,N_3799,N_3783);
and U3843 (N_3843,N_3732,N_3779);
nand U3844 (N_3844,N_3787,N_3782);
or U3845 (N_3845,N_3744,N_3795);
or U3846 (N_3846,N_3784,N_3730);
nor U3847 (N_3847,N_3761,N_3770);
and U3848 (N_3848,N_3706,N_3767);
or U3849 (N_3849,N_3731,N_3717);
nor U3850 (N_3850,N_3748,N_3702);
nand U3851 (N_3851,N_3706,N_3719);
nand U3852 (N_3852,N_3704,N_3776);
nor U3853 (N_3853,N_3748,N_3792);
or U3854 (N_3854,N_3790,N_3723);
nand U3855 (N_3855,N_3774,N_3770);
nor U3856 (N_3856,N_3794,N_3703);
nor U3857 (N_3857,N_3768,N_3745);
nor U3858 (N_3858,N_3746,N_3776);
nor U3859 (N_3859,N_3786,N_3720);
or U3860 (N_3860,N_3749,N_3706);
nor U3861 (N_3861,N_3716,N_3744);
and U3862 (N_3862,N_3769,N_3781);
nor U3863 (N_3863,N_3736,N_3759);
or U3864 (N_3864,N_3783,N_3727);
nor U3865 (N_3865,N_3766,N_3788);
nand U3866 (N_3866,N_3771,N_3716);
or U3867 (N_3867,N_3713,N_3759);
nor U3868 (N_3868,N_3757,N_3721);
or U3869 (N_3869,N_3733,N_3768);
and U3870 (N_3870,N_3768,N_3781);
nor U3871 (N_3871,N_3765,N_3799);
nand U3872 (N_3872,N_3744,N_3736);
and U3873 (N_3873,N_3711,N_3756);
nor U3874 (N_3874,N_3740,N_3765);
nor U3875 (N_3875,N_3737,N_3749);
or U3876 (N_3876,N_3787,N_3790);
nand U3877 (N_3877,N_3723,N_3721);
xnor U3878 (N_3878,N_3702,N_3712);
xor U3879 (N_3879,N_3717,N_3702);
or U3880 (N_3880,N_3798,N_3731);
and U3881 (N_3881,N_3762,N_3732);
nor U3882 (N_3882,N_3791,N_3735);
or U3883 (N_3883,N_3799,N_3791);
xnor U3884 (N_3884,N_3745,N_3777);
and U3885 (N_3885,N_3793,N_3764);
nand U3886 (N_3886,N_3717,N_3728);
and U3887 (N_3887,N_3765,N_3756);
nor U3888 (N_3888,N_3792,N_3701);
nand U3889 (N_3889,N_3778,N_3766);
nand U3890 (N_3890,N_3724,N_3735);
nor U3891 (N_3891,N_3723,N_3768);
nor U3892 (N_3892,N_3740,N_3751);
and U3893 (N_3893,N_3745,N_3772);
and U3894 (N_3894,N_3749,N_3761);
nor U3895 (N_3895,N_3702,N_3795);
or U3896 (N_3896,N_3746,N_3793);
nor U3897 (N_3897,N_3762,N_3704);
nand U3898 (N_3898,N_3718,N_3783);
nand U3899 (N_3899,N_3766,N_3762);
nor U3900 (N_3900,N_3842,N_3876);
nor U3901 (N_3901,N_3894,N_3847);
nand U3902 (N_3902,N_3803,N_3885);
and U3903 (N_3903,N_3836,N_3857);
nor U3904 (N_3904,N_3888,N_3851);
or U3905 (N_3905,N_3804,N_3812);
nand U3906 (N_3906,N_3811,N_3897);
or U3907 (N_3907,N_3878,N_3867);
and U3908 (N_3908,N_3840,N_3866);
nor U3909 (N_3909,N_3835,N_3854);
nand U3910 (N_3910,N_3871,N_3898);
nor U3911 (N_3911,N_3831,N_3814);
nor U3912 (N_3912,N_3880,N_3865);
and U3913 (N_3913,N_3853,N_3829);
nor U3914 (N_3914,N_3859,N_3822);
xor U3915 (N_3915,N_3891,N_3849);
and U3916 (N_3916,N_3877,N_3802);
nor U3917 (N_3917,N_3801,N_3852);
or U3918 (N_3918,N_3868,N_3850);
nand U3919 (N_3919,N_3846,N_3809);
nand U3920 (N_3920,N_3856,N_3848);
nor U3921 (N_3921,N_3820,N_3834);
nand U3922 (N_3922,N_3887,N_3832);
and U3923 (N_3923,N_3821,N_3874);
or U3924 (N_3924,N_3861,N_3870);
nand U3925 (N_3925,N_3889,N_3813);
or U3926 (N_3926,N_3893,N_3863);
and U3927 (N_3927,N_3819,N_3862);
nand U3928 (N_3928,N_3839,N_3841);
and U3929 (N_3929,N_3872,N_3825);
and U3930 (N_3930,N_3899,N_3830);
nor U3931 (N_3931,N_3828,N_3858);
nand U3932 (N_3932,N_3805,N_3807);
and U3933 (N_3933,N_3808,N_3843);
nor U3934 (N_3934,N_3884,N_3806);
nand U3935 (N_3935,N_3833,N_3810);
nor U3936 (N_3936,N_3881,N_3815);
nand U3937 (N_3937,N_3879,N_3864);
nand U3938 (N_3938,N_3855,N_3890);
nand U3939 (N_3939,N_3860,N_3800);
or U3940 (N_3940,N_3869,N_3817);
nand U3941 (N_3941,N_3886,N_3895);
and U3942 (N_3942,N_3882,N_3896);
or U3943 (N_3943,N_3837,N_3827);
nand U3944 (N_3944,N_3823,N_3818);
and U3945 (N_3945,N_3824,N_3838);
and U3946 (N_3946,N_3875,N_3892);
nor U3947 (N_3947,N_3826,N_3816);
or U3948 (N_3948,N_3844,N_3873);
or U3949 (N_3949,N_3883,N_3845);
nor U3950 (N_3950,N_3823,N_3890);
nor U3951 (N_3951,N_3834,N_3871);
nor U3952 (N_3952,N_3840,N_3810);
and U3953 (N_3953,N_3837,N_3814);
nand U3954 (N_3954,N_3855,N_3842);
and U3955 (N_3955,N_3859,N_3890);
nor U3956 (N_3956,N_3894,N_3843);
xor U3957 (N_3957,N_3851,N_3850);
or U3958 (N_3958,N_3821,N_3859);
or U3959 (N_3959,N_3856,N_3837);
nor U3960 (N_3960,N_3852,N_3891);
nand U3961 (N_3961,N_3840,N_3816);
or U3962 (N_3962,N_3843,N_3823);
and U3963 (N_3963,N_3837,N_3875);
nor U3964 (N_3964,N_3859,N_3816);
or U3965 (N_3965,N_3840,N_3870);
and U3966 (N_3966,N_3859,N_3864);
nand U3967 (N_3967,N_3848,N_3876);
nand U3968 (N_3968,N_3895,N_3864);
and U3969 (N_3969,N_3871,N_3883);
nor U3970 (N_3970,N_3826,N_3899);
or U3971 (N_3971,N_3872,N_3881);
and U3972 (N_3972,N_3853,N_3880);
nand U3973 (N_3973,N_3851,N_3827);
nand U3974 (N_3974,N_3801,N_3818);
xnor U3975 (N_3975,N_3866,N_3839);
nor U3976 (N_3976,N_3828,N_3862);
and U3977 (N_3977,N_3815,N_3851);
or U3978 (N_3978,N_3838,N_3839);
nor U3979 (N_3979,N_3850,N_3877);
nor U3980 (N_3980,N_3871,N_3875);
or U3981 (N_3981,N_3800,N_3868);
or U3982 (N_3982,N_3861,N_3890);
nor U3983 (N_3983,N_3876,N_3853);
nor U3984 (N_3984,N_3899,N_3867);
nor U3985 (N_3985,N_3815,N_3835);
nor U3986 (N_3986,N_3851,N_3876);
nand U3987 (N_3987,N_3818,N_3832);
nand U3988 (N_3988,N_3858,N_3851);
nand U3989 (N_3989,N_3881,N_3878);
or U3990 (N_3990,N_3868,N_3825);
nor U3991 (N_3991,N_3849,N_3877);
or U3992 (N_3992,N_3893,N_3869);
and U3993 (N_3993,N_3801,N_3841);
or U3994 (N_3994,N_3892,N_3820);
nand U3995 (N_3995,N_3897,N_3873);
and U3996 (N_3996,N_3873,N_3889);
nor U3997 (N_3997,N_3855,N_3899);
nor U3998 (N_3998,N_3815,N_3869);
nor U3999 (N_3999,N_3881,N_3873);
and U4000 (N_4000,N_3993,N_3950);
nand U4001 (N_4001,N_3926,N_3935);
nor U4002 (N_4002,N_3998,N_3949);
nor U4003 (N_4003,N_3985,N_3932);
nor U4004 (N_4004,N_3909,N_3994);
or U4005 (N_4005,N_3918,N_3944);
nand U4006 (N_4006,N_3900,N_3999);
nor U4007 (N_4007,N_3964,N_3948);
and U4008 (N_4008,N_3924,N_3981);
and U4009 (N_4009,N_3960,N_3952);
nor U4010 (N_4010,N_3934,N_3906);
nor U4011 (N_4011,N_3951,N_3915);
or U4012 (N_4012,N_3989,N_3992);
nor U4013 (N_4013,N_3930,N_3961);
nand U4014 (N_4014,N_3931,N_3954);
nor U4015 (N_4015,N_3958,N_3920);
nand U4016 (N_4016,N_3955,N_3916);
and U4017 (N_4017,N_3974,N_3956);
and U4018 (N_4018,N_3902,N_3953);
nor U4019 (N_4019,N_3904,N_3969);
and U4020 (N_4020,N_3907,N_3959);
nand U4021 (N_4021,N_3984,N_3982);
nand U4022 (N_4022,N_3928,N_3991);
nor U4023 (N_4023,N_3923,N_3990);
nor U4024 (N_4024,N_3977,N_3936);
or U4025 (N_4025,N_3967,N_3925);
nand U4026 (N_4026,N_3940,N_3913);
or U4027 (N_4027,N_3976,N_3914);
and U4028 (N_4028,N_3903,N_3997);
nor U4029 (N_4029,N_3927,N_3996);
or U4030 (N_4030,N_3922,N_3975);
nor U4031 (N_4031,N_3946,N_3968);
or U4032 (N_4032,N_3901,N_3987);
and U4033 (N_4033,N_3917,N_3980);
and U4034 (N_4034,N_3911,N_3986);
nor U4035 (N_4035,N_3965,N_3937);
and U4036 (N_4036,N_3962,N_3963);
nor U4037 (N_4037,N_3910,N_3957);
and U4038 (N_4038,N_3971,N_3943);
xor U4039 (N_4039,N_3947,N_3938);
nand U4040 (N_4040,N_3983,N_3905);
and U4041 (N_4041,N_3970,N_3929);
nor U4042 (N_4042,N_3919,N_3933);
and U4043 (N_4043,N_3988,N_3966);
and U4044 (N_4044,N_3945,N_3939);
nor U4045 (N_4045,N_3942,N_3941);
nand U4046 (N_4046,N_3973,N_3908);
and U4047 (N_4047,N_3912,N_3995);
nand U4048 (N_4048,N_3979,N_3978);
nand U4049 (N_4049,N_3972,N_3921);
nand U4050 (N_4050,N_3953,N_3913);
nor U4051 (N_4051,N_3937,N_3971);
nand U4052 (N_4052,N_3973,N_3917);
nand U4053 (N_4053,N_3931,N_3912);
nand U4054 (N_4054,N_3974,N_3978);
and U4055 (N_4055,N_3994,N_3965);
or U4056 (N_4056,N_3915,N_3920);
nand U4057 (N_4057,N_3929,N_3975);
or U4058 (N_4058,N_3984,N_3926);
or U4059 (N_4059,N_3986,N_3949);
nor U4060 (N_4060,N_3901,N_3928);
and U4061 (N_4061,N_3949,N_3907);
nand U4062 (N_4062,N_3946,N_3966);
and U4063 (N_4063,N_3913,N_3990);
nor U4064 (N_4064,N_3903,N_3912);
nor U4065 (N_4065,N_3920,N_3979);
and U4066 (N_4066,N_3954,N_3984);
nor U4067 (N_4067,N_3976,N_3965);
or U4068 (N_4068,N_3904,N_3992);
nor U4069 (N_4069,N_3989,N_3948);
nor U4070 (N_4070,N_3995,N_3972);
nand U4071 (N_4071,N_3921,N_3997);
nand U4072 (N_4072,N_3958,N_3961);
nand U4073 (N_4073,N_3977,N_3989);
and U4074 (N_4074,N_3929,N_3996);
and U4075 (N_4075,N_3940,N_3968);
nor U4076 (N_4076,N_3912,N_3979);
nor U4077 (N_4077,N_3960,N_3945);
and U4078 (N_4078,N_3934,N_3990);
nor U4079 (N_4079,N_3960,N_3923);
and U4080 (N_4080,N_3997,N_3943);
or U4081 (N_4081,N_3905,N_3991);
nand U4082 (N_4082,N_3911,N_3936);
nor U4083 (N_4083,N_3995,N_3945);
or U4084 (N_4084,N_3979,N_3974);
and U4085 (N_4085,N_3905,N_3915);
nand U4086 (N_4086,N_3935,N_3946);
nor U4087 (N_4087,N_3960,N_3934);
nor U4088 (N_4088,N_3997,N_3901);
nor U4089 (N_4089,N_3968,N_3939);
nand U4090 (N_4090,N_3965,N_3911);
nand U4091 (N_4091,N_3931,N_3983);
and U4092 (N_4092,N_3947,N_3997);
or U4093 (N_4093,N_3970,N_3955);
or U4094 (N_4094,N_3927,N_3988);
and U4095 (N_4095,N_3941,N_3956);
and U4096 (N_4096,N_3993,N_3910);
nand U4097 (N_4097,N_3912,N_3948);
nor U4098 (N_4098,N_3923,N_3928);
nor U4099 (N_4099,N_3917,N_3984);
or U4100 (N_4100,N_4032,N_4069);
nand U4101 (N_4101,N_4041,N_4010);
nor U4102 (N_4102,N_4071,N_4058);
nand U4103 (N_4103,N_4019,N_4080);
nor U4104 (N_4104,N_4089,N_4060);
nor U4105 (N_4105,N_4022,N_4084);
and U4106 (N_4106,N_4024,N_4059);
nand U4107 (N_4107,N_4067,N_4087);
nand U4108 (N_4108,N_4012,N_4030);
or U4109 (N_4109,N_4051,N_4001);
nor U4110 (N_4110,N_4074,N_4063);
and U4111 (N_4111,N_4085,N_4025);
or U4112 (N_4112,N_4002,N_4064);
and U4113 (N_4113,N_4053,N_4004);
nand U4114 (N_4114,N_4011,N_4061);
nand U4115 (N_4115,N_4018,N_4016);
nor U4116 (N_4116,N_4037,N_4076);
and U4117 (N_4117,N_4055,N_4014);
nand U4118 (N_4118,N_4082,N_4013);
nor U4119 (N_4119,N_4054,N_4027);
or U4120 (N_4120,N_4044,N_4007);
nor U4121 (N_4121,N_4094,N_4034);
nand U4122 (N_4122,N_4042,N_4021);
and U4123 (N_4123,N_4046,N_4068);
and U4124 (N_4124,N_4088,N_4056);
nor U4125 (N_4125,N_4073,N_4003);
nand U4126 (N_4126,N_4083,N_4049);
nand U4127 (N_4127,N_4052,N_4048);
xnor U4128 (N_4128,N_4065,N_4006);
nand U4129 (N_4129,N_4008,N_4079);
nor U4130 (N_4130,N_4072,N_4029);
nor U4131 (N_4131,N_4036,N_4099);
nand U4132 (N_4132,N_4081,N_4028);
and U4133 (N_4133,N_4095,N_4026);
nor U4134 (N_4134,N_4020,N_4050);
nor U4135 (N_4135,N_4077,N_4045);
and U4136 (N_4136,N_4035,N_4038);
or U4137 (N_4137,N_4009,N_4057);
and U4138 (N_4138,N_4043,N_4023);
and U4139 (N_4139,N_4031,N_4078);
and U4140 (N_4140,N_4098,N_4005);
nor U4141 (N_4141,N_4097,N_4015);
and U4142 (N_4142,N_4017,N_4086);
nor U4143 (N_4143,N_4075,N_4090);
and U4144 (N_4144,N_4070,N_4040);
or U4145 (N_4145,N_4093,N_4062);
nor U4146 (N_4146,N_4033,N_4039);
or U4147 (N_4147,N_4096,N_4000);
or U4148 (N_4148,N_4092,N_4047);
nor U4149 (N_4149,N_4091,N_4066);
or U4150 (N_4150,N_4057,N_4084);
nor U4151 (N_4151,N_4026,N_4051);
or U4152 (N_4152,N_4072,N_4094);
and U4153 (N_4153,N_4002,N_4058);
nand U4154 (N_4154,N_4029,N_4002);
nor U4155 (N_4155,N_4024,N_4087);
nor U4156 (N_4156,N_4015,N_4044);
and U4157 (N_4157,N_4025,N_4054);
and U4158 (N_4158,N_4017,N_4060);
nor U4159 (N_4159,N_4027,N_4029);
and U4160 (N_4160,N_4004,N_4092);
nor U4161 (N_4161,N_4062,N_4064);
and U4162 (N_4162,N_4065,N_4023);
or U4163 (N_4163,N_4017,N_4002);
nor U4164 (N_4164,N_4076,N_4077);
or U4165 (N_4165,N_4015,N_4092);
nor U4166 (N_4166,N_4004,N_4022);
nor U4167 (N_4167,N_4018,N_4079);
nand U4168 (N_4168,N_4092,N_4029);
nand U4169 (N_4169,N_4030,N_4079);
or U4170 (N_4170,N_4012,N_4032);
nand U4171 (N_4171,N_4092,N_4067);
nand U4172 (N_4172,N_4072,N_4011);
and U4173 (N_4173,N_4056,N_4019);
and U4174 (N_4174,N_4004,N_4032);
nor U4175 (N_4175,N_4032,N_4083);
or U4176 (N_4176,N_4075,N_4044);
or U4177 (N_4177,N_4060,N_4015);
nand U4178 (N_4178,N_4058,N_4090);
nand U4179 (N_4179,N_4020,N_4051);
nand U4180 (N_4180,N_4011,N_4008);
or U4181 (N_4181,N_4028,N_4080);
nand U4182 (N_4182,N_4079,N_4092);
nor U4183 (N_4183,N_4014,N_4062);
nand U4184 (N_4184,N_4029,N_4070);
nor U4185 (N_4185,N_4077,N_4094);
or U4186 (N_4186,N_4074,N_4008);
nor U4187 (N_4187,N_4084,N_4068);
and U4188 (N_4188,N_4000,N_4081);
and U4189 (N_4189,N_4044,N_4085);
nor U4190 (N_4190,N_4001,N_4006);
and U4191 (N_4191,N_4000,N_4013);
nand U4192 (N_4192,N_4088,N_4070);
or U4193 (N_4193,N_4034,N_4005);
nand U4194 (N_4194,N_4051,N_4049);
and U4195 (N_4195,N_4063,N_4085);
or U4196 (N_4196,N_4063,N_4008);
nand U4197 (N_4197,N_4058,N_4093);
nand U4198 (N_4198,N_4088,N_4041);
and U4199 (N_4199,N_4023,N_4007);
and U4200 (N_4200,N_4137,N_4121);
nand U4201 (N_4201,N_4140,N_4103);
or U4202 (N_4202,N_4179,N_4172);
and U4203 (N_4203,N_4186,N_4170);
nand U4204 (N_4204,N_4136,N_4129);
nor U4205 (N_4205,N_4183,N_4181);
nand U4206 (N_4206,N_4162,N_4128);
and U4207 (N_4207,N_4138,N_4143);
nand U4208 (N_4208,N_4104,N_4106);
nor U4209 (N_4209,N_4149,N_4130);
nand U4210 (N_4210,N_4173,N_4175);
nor U4211 (N_4211,N_4192,N_4180);
nor U4212 (N_4212,N_4188,N_4124);
and U4213 (N_4213,N_4101,N_4161);
or U4214 (N_4214,N_4108,N_4195);
or U4215 (N_4215,N_4182,N_4166);
nand U4216 (N_4216,N_4145,N_4132);
nor U4217 (N_4217,N_4157,N_4159);
nand U4218 (N_4218,N_4113,N_4153);
or U4219 (N_4219,N_4174,N_4123);
nor U4220 (N_4220,N_4142,N_4135);
nand U4221 (N_4221,N_4100,N_4118);
and U4222 (N_4222,N_4111,N_4178);
nor U4223 (N_4223,N_4165,N_4158);
and U4224 (N_4224,N_4126,N_4120);
nand U4225 (N_4225,N_4107,N_4169);
nand U4226 (N_4226,N_4148,N_4134);
nor U4227 (N_4227,N_4154,N_4171);
and U4228 (N_4228,N_4125,N_4190);
and U4229 (N_4229,N_4168,N_4109);
nor U4230 (N_4230,N_4133,N_4102);
nor U4231 (N_4231,N_4176,N_4114);
or U4232 (N_4232,N_4117,N_4150);
or U4233 (N_4233,N_4131,N_4147);
and U4234 (N_4234,N_4184,N_4191);
nand U4235 (N_4235,N_4196,N_4199);
and U4236 (N_4236,N_4163,N_4160);
nand U4237 (N_4237,N_4156,N_4167);
nor U4238 (N_4238,N_4112,N_4164);
and U4239 (N_4239,N_4139,N_4151);
or U4240 (N_4240,N_4105,N_4116);
or U4241 (N_4241,N_4127,N_4115);
nand U4242 (N_4242,N_4197,N_4152);
and U4243 (N_4243,N_4119,N_4185);
nand U4244 (N_4244,N_4189,N_4141);
or U4245 (N_4245,N_4122,N_4198);
and U4246 (N_4246,N_4194,N_4144);
and U4247 (N_4247,N_4110,N_4146);
nand U4248 (N_4248,N_4155,N_4193);
or U4249 (N_4249,N_4177,N_4187);
and U4250 (N_4250,N_4101,N_4117);
and U4251 (N_4251,N_4185,N_4165);
or U4252 (N_4252,N_4149,N_4191);
nor U4253 (N_4253,N_4193,N_4150);
and U4254 (N_4254,N_4149,N_4150);
nand U4255 (N_4255,N_4199,N_4193);
or U4256 (N_4256,N_4174,N_4176);
and U4257 (N_4257,N_4131,N_4151);
or U4258 (N_4258,N_4196,N_4110);
and U4259 (N_4259,N_4130,N_4119);
nor U4260 (N_4260,N_4166,N_4177);
and U4261 (N_4261,N_4101,N_4104);
or U4262 (N_4262,N_4153,N_4114);
and U4263 (N_4263,N_4150,N_4130);
nor U4264 (N_4264,N_4135,N_4163);
nor U4265 (N_4265,N_4102,N_4189);
nor U4266 (N_4266,N_4116,N_4160);
or U4267 (N_4267,N_4161,N_4120);
nor U4268 (N_4268,N_4174,N_4148);
nand U4269 (N_4269,N_4199,N_4139);
or U4270 (N_4270,N_4199,N_4121);
nand U4271 (N_4271,N_4172,N_4105);
nor U4272 (N_4272,N_4174,N_4155);
or U4273 (N_4273,N_4105,N_4156);
nand U4274 (N_4274,N_4132,N_4143);
and U4275 (N_4275,N_4132,N_4144);
nand U4276 (N_4276,N_4122,N_4180);
nor U4277 (N_4277,N_4119,N_4153);
nor U4278 (N_4278,N_4196,N_4109);
and U4279 (N_4279,N_4130,N_4179);
nand U4280 (N_4280,N_4105,N_4142);
xnor U4281 (N_4281,N_4131,N_4129);
and U4282 (N_4282,N_4132,N_4122);
or U4283 (N_4283,N_4120,N_4194);
nand U4284 (N_4284,N_4168,N_4149);
and U4285 (N_4285,N_4193,N_4156);
and U4286 (N_4286,N_4185,N_4182);
nand U4287 (N_4287,N_4136,N_4103);
and U4288 (N_4288,N_4164,N_4195);
and U4289 (N_4289,N_4194,N_4143);
nor U4290 (N_4290,N_4135,N_4128);
nand U4291 (N_4291,N_4135,N_4130);
nand U4292 (N_4292,N_4181,N_4177);
nor U4293 (N_4293,N_4112,N_4138);
or U4294 (N_4294,N_4185,N_4173);
nand U4295 (N_4295,N_4116,N_4159);
nand U4296 (N_4296,N_4167,N_4199);
nor U4297 (N_4297,N_4139,N_4177);
or U4298 (N_4298,N_4193,N_4113);
xnor U4299 (N_4299,N_4111,N_4123);
and U4300 (N_4300,N_4213,N_4258);
or U4301 (N_4301,N_4204,N_4293);
nor U4302 (N_4302,N_4264,N_4208);
and U4303 (N_4303,N_4248,N_4242);
or U4304 (N_4304,N_4239,N_4270);
nand U4305 (N_4305,N_4294,N_4206);
and U4306 (N_4306,N_4202,N_4275);
nand U4307 (N_4307,N_4254,N_4238);
or U4308 (N_4308,N_4255,N_4233);
nand U4309 (N_4309,N_4219,N_4227);
nor U4310 (N_4310,N_4297,N_4291);
and U4311 (N_4311,N_4234,N_4220);
xnor U4312 (N_4312,N_4201,N_4262);
nand U4313 (N_4313,N_4261,N_4205);
nand U4314 (N_4314,N_4276,N_4250);
or U4315 (N_4315,N_4232,N_4237);
and U4316 (N_4316,N_4229,N_4221);
and U4317 (N_4317,N_4286,N_4226);
nor U4318 (N_4318,N_4245,N_4282);
and U4319 (N_4319,N_4216,N_4296);
and U4320 (N_4320,N_4247,N_4284);
xnor U4321 (N_4321,N_4260,N_4299);
and U4322 (N_4322,N_4278,N_4223);
nand U4323 (N_4323,N_4289,N_4225);
or U4324 (N_4324,N_4235,N_4280);
or U4325 (N_4325,N_4253,N_4271);
and U4326 (N_4326,N_4277,N_4298);
or U4327 (N_4327,N_4222,N_4285);
or U4328 (N_4328,N_4288,N_4281);
and U4329 (N_4329,N_4266,N_4265);
nor U4330 (N_4330,N_4292,N_4267);
and U4331 (N_4331,N_4215,N_4203);
or U4332 (N_4332,N_4273,N_4274);
and U4333 (N_4333,N_4257,N_4210);
nand U4334 (N_4334,N_4207,N_4246);
nand U4335 (N_4335,N_4295,N_4251);
and U4336 (N_4336,N_4211,N_4252);
nand U4337 (N_4337,N_4230,N_4200);
and U4338 (N_4338,N_4256,N_4224);
or U4339 (N_4339,N_4269,N_4217);
and U4340 (N_4340,N_4249,N_4290);
and U4341 (N_4341,N_4283,N_4214);
nand U4342 (N_4342,N_4231,N_4272);
and U4343 (N_4343,N_4236,N_4244);
nor U4344 (N_4344,N_4218,N_4243);
nand U4345 (N_4345,N_4228,N_4212);
or U4346 (N_4346,N_4263,N_4279);
nor U4347 (N_4347,N_4209,N_4259);
and U4348 (N_4348,N_4268,N_4287);
nand U4349 (N_4349,N_4240,N_4241);
nor U4350 (N_4350,N_4288,N_4217);
nand U4351 (N_4351,N_4284,N_4281);
nor U4352 (N_4352,N_4277,N_4206);
or U4353 (N_4353,N_4287,N_4265);
or U4354 (N_4354,N_4206,N_4230);
nor U4355 (N_4355,N_4273,N_4248);
or U4356 (N_4356,N_4278,N_4221);
or U4357 (N_4357,N_4251,N_4270);
or U4358 (N_4358,N_4295,N_4204);
xnor U4359 (N_4359,N_4276,N_4268);
or U4360 (N_4360,N_4213,N_4277);
nand U4361 (N_4361,N_4219,N_4233);
nor U4362 (N_4362,N_4201,N_4267);
and U4363 (N_4363,N_4209,N_4265);
or U4364 (N_4364,N_4230,N_4225);
nand U4365 (N_4365,N_4226,N_4261);
or U4366 (N_4366,N_4254,N_4216);
nor U4367 (N_4367,N_4239,N_4269);
or U4368 (N_4368,N_4272,N_4238);
nor U4369 (N_4369,N_4261,N_4276);
and U4370 (N_4370,N_4291,N_4236);
nand U4371 (N_4371,N_4230,N_4274);
and U4372 (N_4372,N_4230,N_4282);
and U4373 (N_4373,N_4292,N_4268);
or U4374 (N_4374,N_4242,N_4218);
or U4375 (N_4375,N_4249,N_4284);
nor U4376 (N_4376,N_4205,N_4241);
and U4377 (N_4377,N_4258,N_4271);
and U4378 (N_4378,N_4210,N_4277);
or U4379 (N_4379,N_4218,N_4239);
nand U4380 (N_4380,N_4229,N_4286);
or U4381 (N_4381,N_4260,N_4251);
nor U4382 (N_4382,N_4231,N_4236);
or U4383 (N_4383,N_4255,N_4253);
nand U4384 (N_4384,N_4268,N_4206);
and U4385 (N_4385,N_4289,N_4236);
or U4386 (N_4386,N_4239,N_4282);
or U4387 (N_4387,N_4240,N_4201);
or U4388 (N_4388,N_4284,N_4251);
or U4389 (N_4389,N_4232,N_4263);
or U4390 (N_4390,N_4292,N_4269);
or U4391 (N_4391,N_4241,N_4266);
and U4392 (N_4392,N_4231,N_4257);
nand U4393 (N_4393,N_4225,N_4282);
or U4394 (N_4394,N_4293,N_4224);
or U4395 (N_4395,N_4281,N_4290);
nor U4396 (N_4396,N_4222,N_4276);
and U4397 (N_4397,N_4245,N_4274);
nand U4398 (N_4398,N_4286,N_4292);
and U4399 (N_4399,N_4290,N_4244);
nand U4400 (N_4400,N_4341,N_4386);
nor U4401 (N_4401,N_4337,N_4324);
nor U4402 (N_4402,N_4390,N_4330);
nor U4403 (N_4403,N_4392,N_4328);
or U4404 (N_4404,N_4394,N_4355);
or U4405 (N_4405,N_4387,N_4314);
or U4406 (N_4406,N_4320,N_4385);
nor U4407 (N_4407,N_4393,N_4353);
nand U4408 (N_4408,N_4371,N_4308);
nor U4409 (N_4409,N_4348,N_4366);
nand U4410 (N_4410,N_4309,N_4399);
nor U4411 (N_4411,N_4327,N_4360);
and U4412 (N_4412,N_4322,N_4323);
or U4413 (N_4413,N_4333,N_4347);
and U4414 (N_4414,N_4375,N_4344);
xor U4415 (N_4415,N_4326,N_4365);
nor U4416 (N_4416,N_4357,N_4319);
nand U4417 (N_4417,N_4305,N_4313);
or U4418 (N_4418,N_4363,N_4332);
nor U4419 (N_4419,N_4389,N_4346);
nor U4420 (N_4420,N_4339,N_4372);
nand U4421 (N_4421,N_4345,N_4310);
or U4422 (N_4422,N_4349,N_4398);
nor U4423 (N_4423,N_4343,N_4376);
nand U4424 (N_4424,N_4378,N_4359);
nand U4425 (N_4425,N_4354,N_4334);
or U4426 (N_4426,N_4311,N_4396);
or U4427 (N_4427,N_4361,N_4374);
nor U4428 (N_4428,N_4367,N_4300);
or U4429 (N_4429,N_4342,N_4397);
and U4430 (N_4430,N_4307,N_4350);
or U4431 (N_4431,N_4381,N_4336);
nor U4432 (N_4432,N_4368,N_4321);
or U4433 (N_4433,N_4306,N_4329);
or U4434 (N_4434,N_4395,N_4391);
nor U4435 (N_4435,N_4304,N_4317);
and U4436 (N_4436,N_4351,N_4370);
and U4437 (N_4437,N_4318,N_4362);
nand U4438 (N_4438,N_4316,N_4301);
or U4439 (N_4439,N_4356,N_4377);
nand U4440 (N_4440,N_4302,N_4340);
nand U4441 (N_4441,N_4384,N_4373);
or U4442 (N_4442,N_4315,N_4369);
or U4443 (N_4443,N_4380,N_4338);
and U4444 (N_4444,N_4358,N_4388);
nand U4445 (N_4445,N_4325,N_4364);
or U4446 (N_4446,N_4383,N_4303);
and U4447 (N_4447,N_4379,N_4352);
nor U4448 (N_4448,N_4331,N_4382);
nand U4449 (N_4449,N_4335,N_4312);
nand U4450 (N_4450,N_4399,N_4315);
nor U4451 (N_4451,N_4327,N_4392);
xor U4452 (N_4452,N_4336,N_4377);
or U4453 (N_4453,N_4373,N_4335);
and U4454 (N_4454,N_4307,N_4382);
and U4455 (N_4455,N_4399,N_4325);
and U4456 (N_4456,N_4364,N_4324);
nand U4457 (N_4457,N_4369,N_4334);
nor U4458 (N_4458,N_4364,N_4326);
nor U4459 (N_4459,N_4338,N_4397);
nor U4460 (N_4460,N_4387,N_4339);
and U4461 (N_4461,N_4312,N_4377);
nor U4462 (N_4462,N_4362,N_4349);
and U4463 (N_4463,N_4389,N_4327);
nor U4464 (N_4464,N_4347,N_4317);
nor U4465 (N_4465,N_4366,N_4352);
or U4466 (N_4466,N_4367,N_4316);
or U4467 (N_4467,N_4326,N_4331);
nor U4468 (N_4468,N_4378,N_4329);
nand U4469 (N_4469,N_4321,N_4352);
and U4470 (N_4470,N_4309,N_4322);
nand U4471 (N_4471,N_4359,N_4343);
or U4472 (N_4472,N_4375,N_4358);
nand U4473 (N_4473,N_4384,N_4327);
nor U4474 (N_4474,N_4346,N_4353);
nor U4475 (N_4475,N_4392,N_4330);
or U4476 (N_4476,N_4357,N_4317);
nor U4477 (N_4477,N_4323,N_4306);
nand U4478 (N_4478,N_4373,N_4300);
nand U4479 (N_4479,N_4349,N_4304);
and U4480 (N_4480,N_4305,N_4319);
nor U4481 (N_4481,N_4377,N_4326);
or U4482 (N_4482,N_4397,N_4316);
and U4483 (N_4483,N_4357,N_4391);
or U4484 (N_4484,N_4324,N_4382);
nand U4485 (N_4485,N_4308,N_4342);
nor U4486 (N_4486,N_4350,N_4347);
and U4487 (N_4487,N_4308,N_4384);
nor U4488 (N_4488,N_4395,N_4325);
nor U4489 (N_4489,N_4359,N_4321);
nor U4490 (N_4490,N_4367,N_4394);
nand U4491 (N_4491,N_4364,N_4358);
or U4492 (N_4492,N_4318,N_4303);
or U4493 (N_4493,N_4366,N_4329);
or U4494 (N_4494,N_4300,N_4392);
nand U4495 (N_4495,N_4344,N_4322);
nand U4496 (N_4496,N_4399,N_4337);
nor U4497 (N_4497,N_4367,N_4315);
or U4498 (N_4498,N_4384,N_4389);
nor U4499 (N_4499,N_4361,N_4354);
nor U4500 (N_4500,N_4451,N_4444);
nor U4501 (N_4501,N_4426,N_4434);
nor U4502 (N_4502,N_4424,N_4453);
and U4503 (N_4503,N_4496,N_4448);
and U4504 (N_4504,N_4464,N_4410);
nor U4505 (N_4505,N_4477,N_4482);
nand U4506 (N_4506,N_4435,N_4468);
and U4507 (N_4507,N_4474,N_4483);
or U4508 (N_4508,N_4432,N_4416);
nor U4509 (N_4509,N_4462,N_4429);
or U4510 (N_4510,N_4454,N_4459);
or U4511 (N_4511,N_4420,N_4460);
and U4512 (N_4512,N_4438,N_4415);
and U4513 (N_4513,N_4422,N_4463);
or U4514 (N_4514,N_4405,N_4437);
nand U4515 (N_4515,N_4430,N_4495);
or U4516 (N_4516,N_4473,N_4469);
or U4517 (N_4517,N_4498,N_4466);
nand U4518 (N_4518,N_4404,N_4445);
or U4519 (N_4519,N_4493,N_4476);
nand U4520 (N_4520,N_4492,N_4490);
or U4521 (N_4521,N_4414,N_4479);
nor U4522 (N_4522,N_4409,N_4488);
or U4523 (N_4523,N_4400,N_4470);
nor U4524 (N_4524,N_4455,N_4408);
nor U4525 (N_4525,N_4442,N_4478);
and U4526 (N_4526,N_4457,N_4497);
nand U4527 (N_4527,N_4428,N_4458);
nand U4528 (N_4528,N_4494,N_4402);
and U4529 (N_4529,N_4401,N_4487);
nand U4530 (N_4530,N_4418,N_4436);
and U4531 (N_4531,N_4431,N_4417);
nand U4532 (N_4532,N_4439,N_4461);
nand U4533 (N_4533,N_4412,N_4449);
and U4534 (N_4534,N_4440,N_4407);
nand U4535 (N_4535,N_4465,N_4433);
nand U4536 (N_4536,N_4489,N_4456);
nor U4537 (N_4537,N_4472,N_4481);
nand U4538 (N_4538,N_4421,N_4475);
and U4539 (N_4539,N_4441,N_4425);
or U4540 (N_4540,N_4485,N_4467);
nand U4541 (N_4541,N_4446,N_4480);
or U4542 (N_4542,N_4411,N_4484);
nand U4543 (N_4543,N_4471,N_4403);
nand U4544 (N_4544,N_4413,N_4443);
nor U4545 (N_4545,N_4419,N_4450);
or U4546 (N_4546,N_4499,N_4423);
and U4547 (N_4547,N_4491,N_4452);
nand U4548 (N_4548,N_4486,N_4406);
and U4549 (N_4549,N_4447,N_4427);
and U4550 (N_4550,N_4464,N_4475);
nand U4551 (N_4551,N_4465,N_4477);
nor U4552 (N_4552,N_4416,N_4425);
and U4553 (N_4553,N_4459,N_4445);
nand U4554 (N_4554,N_4461,N_4433);
nand U4555 (N_4555,N_4462,N_4438);
nand U4556 (N_4556,N_4436,N_4481);
nand U4557 (N_4557,N_4482,N_4467);
and U4558 (N_4558,N_4401,N_4443);
or U4559 (N_4559,N_4490,N_4443);
and U4560 (N_4560,N_4409,N_4479);
nor U4561 (N_4561,N_4445,N_4402);
nor U4562 (N_4562,N_4479,N_4449);
nor U4563 (N_4563,N_4414,N_4402);
nor U4564 (N_4564,N_4418,N_4450);
nand U4565 (N_4565,N_4489,N_4406);
nand U4566 (N_4566,N_4417,N_4426);
or U4567 (N_4567,N_4407,N_4424);
nand U4568 (N_4568,N_4481,N_4484);
nor U4569 (N_4569,N_4426,N_4429);
and U4570 (N_4570,N_4410,N_4422);
and U4571 (N_4571,N_4490,N_4419);
and U4572 (N_4572,N_4446,N_4431);
nand U4573 (N_4573,N_4445,N_4493);
and U4574 (N_4574,N_4460,N_4434);
or U4575 (N_4575,N_4415,N_4441);
or U4576 (N_4576,N_4491,N_4442);
nand U4577 (N_4577,N_4402,N_4456);
nand U4578 (N_4578,N_4488,N_4456);
and U4579 (N_4579,N_4432,N_4464);
and U4580 (N_4580,N_4468,N_4466);
nand U4581 (N_4581,N_4427,N_4412);
or U4582 (N_4582,N_4476,N_4431);
nor U4583 (N_4583,N_4408,N_4474);
nor U4584 (N_4584,N_4461,N_4483);
or U4585 (N_4585,N_4464,N_4460);
or U4586 (N_4586,N_4459,N_4463);
and U4587 (N_4587,N_4412,N_4471);
or U4588 (N_4588,N_4490,N_4456);
nor U4589 (N_4589,N_4483,N_4429);
or U4590 (N_4590,N_4410,N_4497);
and U4591 (N_4591,N_4413,N_4475);
nand U4592 (N_4592,N_4419,N_4449);
nand U4593 (N_4593,N_4449,N_4463);
nand U4594 (N_4594,N_4456,N_4494);
and U4595 (N_4595,N_4407,N_4405);
or U4596 (N_4596,N_4499,N_4422);
nor U4597 (N_4597,N_4485,N_4481);
or U4598 (N_4598,N_4447,N_4469);
or U4599 (N_4599,N_4476,N_4442);
nand U4600 (N_4600,N_4561,N_4580);
and U4601 (N_4601,N_4514,N_4520);
or U4602 (N_4602,N_4597,N_4509);
or U4603 (N_4603,N_4559,N_4502);
nor U4604 (N_4604,N_4510,N_4578);
and U4605 (N_4605,N_4550,N_4579);
or U4606 (N_4606,N_4567,N_4554);
and U4607 (N_4607,N_4591,N_4583);
and U4608 (N_4608,N_4584,N_4596);
nor U4609 (N_4609,N_4589,N_4588);
and U4610 (N_4610,N_4531,N_4568);
or U4611 (N_4611,N_4537,N_4529);
nor U4612 (N_4612,N_4595,N_4574);
nand U4613 (N_4613,N_4534,N_4562);
and U4614 (N_4614,N_4540,N_4507);
nor U4615 (N_4615,N_4586,N_4513);
nor U4616 (N_4616,N_4528,N_4503);
and U4617 (N_4617,N_4522,N_4500);
and U4618 (N_4618,N_4530,N_4519);
nor U4619 (N_4619,N_4599,N_4587);
or U4620 (N_4620,N_4524,N_4523);
nor U4621 (N_4621,N_4598,N_4552);
and U4622 (N_4622,N_4585,N_4556);
and U4623 (N_4623,N_4539,N_4551);
and U4624 (N_4624,N_4563,N_4506);
and U4625 (N_4625,N_4504,N_4581);
or U4626 (N_4626,N_4549,N_4511);
and U4627 (N_4627,N_4515,N_4570);
or U4628 (N_4628,N_4516,N_4541);
nand U4629 (N_4629,N_4590,N_4548);
and U4630 (N_4630,N_4536,N_4555);
nand U4631 (N_4631,N_4512,N_4593);
and U4632 (N_4632,N_4582,N_4518);
and U4633 (N_4633,N_4572,N_4560);
nand U4634 (N_4634,N_4538,N_4517);
nand U4635 (N_4635,N_4571,N_4576);
or U4636 (N_4636,N_4532,N_4533);
and U4637 (N_4637,N_4594,N_4592);
nor U4638 (N_4638,N_4545,N_4525);
and U4639 (N_4639,N_4577,N_4526);
nand U4640 (N_4640,N_4547,N_4564);
nor U4641 (N_4641,N_4573,N_4557);
or U4642 (N_4642,N_4535,N_4543);
or U4643 (N_4643,N_4508,N_4569);
nand U4644 (N_4644,N_4553,N_4505);
or U4645 (N_4645,N_4565,N_4558);
and U4646 (N_4646,N_4566,N_4546);
or U4647 (N_4647,N_4501,N_4575);
nand U4648 (N_4648,N_4521,N_4542);
and U4649 (N_4649,N_4527,N_4544);
nor U4650 (N_4650,N_4568,N_4565);
nand U4651 (N_4651,N_4556,N_4584);
nand U4652 (N_4652,N_4512,N_4587);
or U4653 (N_4653,N_4575,N_4545);
nand U4654 (N_4654,N_4533,N_4564);
nand U4655 (N_4655,N_4527,N_4536);
nor U4656 (N_4656,N_4599,N_4523);
or U4657 (N_4657,N_4575,N_4551);
nor U4658 (N_4658,N_4512,N_4581);
nand U4659 (N_4659,N_4534,N_4588);
and U4660 (N_4660,N_4509,N_4527);
nor U4661 (N_4661,N_4525,N_4527);
nor U4662 (N_4662,N_4504,N_4549);
or U4663 (N_4663,N_4579,N_4518);
or U4664 (N_4664,N_4594,N_4510);
nor U4665 (N_4665,N_4555,N_4507);
or U4666 (N_4666,N_4511,N_4584);
and U4667 (N_4667,N_4517,N_4533);
and U4668 (N_4668,N_4562,N_4541);
or U4669 (N_4669,N_4596,N_4512);
nor U4670 (N_4670,N_4564,N_4559);
or U4671 (N_4671,N_4589,N_4553);
nor U4672 (N_4672,N_4503,N_4535);
nor U4673 (N_4673,N_4557,N_4539);
and U4674 (N_4674,N_4549,N_4518);
nand U4675 (N_4675,N_4514,N_4578);
and U4676 (N_4676,N_4536,N_4587);
and U4677 (N_4677,N_4566,N_4592);
nor U4678 (N_4678,N_4567,N_4540);
nand U4679 (N_4679,N_4550,N_4573);
or U4680 (N_4680,N_4585,N_4598);
or U4681 (N_4681,N_4586,N_4529);
nor U4682 (N_4682,N_4573,N_4597);
nand U4683 (N_4683,N_4526,N_4561);
and U4684 (N_4684,N_4548,N_4596);
nand U4685 (N_4685,N_4553,N_4510);
or U4686 (N_4686,N_4522,N_4590);
nor U4687 (N_4687,N_4546,N_4533);
and U4688 (N_4688,N_4560,N_4512);
or U4689 (N_4689,N_4599,N_4566);
and U4690 (N_4690,N_4503,N_4551);
and U4691 (N_4691,N_4565,N_4515);
or U4692 (N_4692,N_4560,N_4597);
and U4693 (N_4693,N_4552,N_4505);
nand U4694 (N_4694,N_4582,N_4589);
nor U4695 (N_4695,N_4539,N_4534);
or U4696 (N_4696,N_4556,N_4583);
nor U4697 (N_4697,N_4584,N_4559);
or U4698 (N_4698,N_4541,N_4519);
nor U4699 (N_4699,N_4538,N_4502);
and U4700 (N_4700,N_4649,N_4682);
and U4701 (N_4701,N_4636,N_4610);
and U4702 (N_4702,N_4643,N_4639);
or U4703 (N_4703,N_4657,N_4613);
and U4704 (N_4704,N_4601,N_4672);
nor U4705 (N_4705,N_4680,N_4681);
or U4706 (N_4706,N_4624,N_4616);
or U4707 (N_4707,N_4602,N_4664);
and U4708 (N_4708,N_4607,N_4663);
nor U4709 (N_4709,N_4658,N_4692);
nand U4710 (N_4710,N_4650,N_4683);
nor U4711 (N_4711,N_4696,N_4697);
nand U4712 (N_4712,N_4675,N_4678);
nor U4713 (N_4713,N_4644,N_4641);
and U4714 (N_4714,N_4669,N_4611);
and U4715 (N_4715,N_4634,N_4653);
and U4716 (N_4716,N_4606,N_4654);
nor U4717 (N_4717,N_4630,N_4620);
or U4718 (N_4718,N_4638,N_4684);
and U4719 (N_4719,N_4688,N_4659);
or U4720 (N_4720,N_4642,N_4617);
nand U4721 (N_4721,N_4637,N_4686);
or U4722 (N_4722,N_4671,N_4646);
nand U4723 (N_4723,N_4615,N_4604);
nor U4724 (N_4724,N_4619,N_4618);
nor U4725 (N_4725,N_4623,N_4679);
and U4726 (N_4726,N_4687,N_4640);
nand U4727 (N_4727,N_4628,N_4677);
nand U4728 (N_4728,N_4690,N_4661);
and U4729 (N_4729,N_4629,N_4689);
nor U4730 (N_4730,N_4633,N_4621);
nor U4731 (N_4731,N_4648,N_4691);
nor U4732 (N_4732,N_4625,N_4656);
and U4733 (N_4733,N_4647,N_4673);
nor U4734 (N_4734,N_4603,N_4614);
nor U4735 (N_4735,N_4627,N_4631);
nand U4736 (N_4736,N_4676,N_4668);
or U4737 (N_4737,N_4670,N_4695);
nand U4738 (N_4738,N_4600,N_4665);
and U4739 (N_4739,N_4632,N_4605);
nor U4740 (N_4740,N_4622,N_4645);
and U4741 (N_4741,N_4608,N_4694);
or U4742 (N_4742,N_4674,N_4626);
nand U4743 (N_4743,N_4693,N_4667);
and U4744 (N_4744,N_4651,N_4699);
nor U4745 (N_4745,N_4698,N_4685);
nand U4746 (N_4746,N_4666,N_4609);
nand U4747 (N_4747,N_4635,N_4660);
nor U4748 (N_4748,N_4655,N_4652);
nand U4749 (N_4749,N_4612,N_4662);
nor U4750 (N_4750,N_4657,N_4614);
or U4751 (N_4751,N_4667,N_4637);
and U4752 (N_4752,N_4687,N_4622);
and U4753 (N_4753,N_4668,N_4616);
nand U4754 (N_4754,N_4667,N_4654);
and U4755 (N_4755,N_4619,N_4656);
nand U4756 (N_4756,N_4666,N_4632);
nor U4757 (N_4757,N_4640,N_4692);
and U4758 (N_4758,N_4636,N_4681);
and U4759 (N_4759,N_4608,N_4659);
or U4760 (N_4760,N_4678,N_4691);
and U4761 (N_4761,N_4616,N_4680);
nor U4762 (N_4762,N_4660,N_4611);
or U4763 (N_4763,N_4618,N_4662);
and U4764 (N_4764,N_4678,N_4644);
and U4765 (N_4765,N_4632,N_4616);
nor U4766 (N_4766,N_4657,N_4655);
or U4767 (N_4767,N_4601,N_4690);
nor U4768 (N_4768,N_4633,N_4627);
xnor U4769 (N_4769,N_4651,N_4670);
nor U4770 (N_4770,N_4611,N_4681);
nand U4771 (N_4771,N_4638,N_4690);
nand U4772 (N_4772,N_4678,N_4613);
or U4773 (N_4773,N_4682,N_4645);
or U4774 (N_4774,N_4682,N_4692);
nor U4775 (N_4775,N_4663,N_4608);
or U4776 (N_4776,N_4632,N_4687);
and U4777 (N_4777,N_4644,N_4602);
and U4778 (N_4778,N_4610,N_4634);
nor U4779 (N_4779,N_4611,N_4613);
nand U4780 (N_4780,N_4694,N_4640);
or U4781 (N_4781,N_4658,N_4652);
nand U4782 (N_4782,N_4617,N_4619);
nand U4783 (N_4783,N_4687,N_4637);
nor U4784 (N_4784,N_4687,N_4633);
nor U4785 (N_4785,N_4634,N_4651);
and U4786 (N_4786,N_4679,N_4680);
and U4787 (N_4787,N_4618,N_4633);
nand U4788 (N_4788,N_4611,N_4684);
or U4789 (N_4789,N_4617,N_4640);
nand U4790 (N_4790,N_4697,N_4623);
and U4791 (N_4791,N_4618,N_4654);
and U4792 (N_4792,N_4651,N_4623);
and U4793 (N_4793,N_4685,N_4622);
and U4794 (N_4794,N_4659,N_4625);
and U4795 (N_4795,N_4658,N_4622);
xor U4796 (N_4796,N_4684,N_4649);
nand U4797 (N_4797,N_4625,N_4623);
nand U4798 (N_4798,N_4653,N_4662);
or U4799 (N_4799,N_4686,N_4690);
nand U4800 (N_4800,N_4740,N_4748);
and U4801 (N_4801,N_4704,N_4737);
or U4802 (N_4802,N_4725,N_4756);
nand U4803 (N_4803,N_4713,N_4750);
nand U4804 (N_4804,N_4724,N_4799);
nand U4805 (N_4805,N_4709,N_4783);
nand U4806 (N_4806,N_4720,N_4702);
and U4807 (N_4807,N_4771,N_4790);
nor U4808 (N_4808,N_4743,N_4739);
nor U4809 (N_4809,N_4787,N_4782);
or U4810 (N_4810,N_4732,N_4745);
or U4811 (N_4811,N_4716,N_4744);
nor U4812 (N_4812,N_4770,N_4728);
nor U4813 (N_4813,N_4736,N_4717);
nand U4814 (N_4814,N_4764,N_4701);
and U4815 (N_4815,N_4793,N_4761);
nor U4816 (N_4816,N_4779,N_4747);
or U4817 (N_4817,N_4773,N_4746);
and U4818 (N_4818,N_4797,N_4796);
or U4819 (N_4819,N_4772,N_4703);
or U4820 (N_4820,N_4731,N_4735);
or U4821 (N_4821,N_4763,N_4733);
or U4822 (N_4822,N_4721,N_4784);
nor U4823 (N_4823,N_4705,N_4708);
or U4824 (N_4824,N_4751,N_4727);
xor U4825 (N_4825,N_4741,N_4700);
nor U4826 (N_4826,N_4719,N_4730);
nor U4827 (N_4827,N_4752,N_4765);
nor U4828 (N_4828,N_4707,N_4769);
nor U4829 (N_4829,N_4785,N_4798);
or U4830 (N_4830,N_4723,N_4759);
and U4831 (N_4831,N_4762,N_4795);
nand U4832 (N_4832,N_4714,N_4757);
and U4833 (N_4833,N_4767,N_4766);
nor U4834 (N_4834,N_4791,N_4753);
nand U4835 (N_4835,N_4775,N_4768);
nand U4836 (N_4836,N_4754,N_4780);
nor U4837 (N_4837,N_4722,N_4776);
nor U4838 (N_4838,N_4760,N_4742);
or U4839 (N_4839,N_4758,N_4711);
nor U4840 (N_4840,N_4710,N_4755);
and U4841 (N_4841,N_4794,N_4777);
nand U4842 (N_4842,N_4706,N_4738);
or U4843 (N_4843,N_4774,N_4726);
or U4844 (N_4844,N_4786,N_4749);
nor U4845 (N_4845,N_4729,N_4718);
nor U4846 (N_4846,N_4778,N_4715);
nand U4847 (N_4847,N_4734,N_4792);
nand U4848 (N_4848,N_4712,N_4789);
or U4849 (N_4849,N_4781,N_4788);
and U4850 (N_4850,N_4710,N_4760);
nor U4851 (N_4851,N_4797,N_4721);
nor U4852 (N_4852,N_4724,N_4745);
nor U4853 (N_4853,N_4763,N_4799);
or U4854 (N_4854,N_4702,N_4712);
and U4855 (N_4855,N_4738,N_4732);
nor U4856 (N_4856,N_4739,N_4715);
and U4857 (N_4857,N_4725,N_4705);
nand U4858 (N_4858,N_4703,N_4796);
or U4859 (N_4859,N_4772,N_4779);
or U4860 (N_4860,N_4756,N_4787);
or U4861 (N_4861,N_4724,N_4782);
or U4862 (N_4862,N_4709,N_4710);
nand U4863 (N_4863,N_4731,N_4726);
nor U4864 (N_4864,N_4717,N_4796);
nand U4865 (N_4865,N_4706,N_4793);
nor U4866 (N_4866,N_4717,N_4773);
or U4867 (N_4867,N_4797,N_4799);
nor U4868 (N_4868,N_4762,N_4723);
nor U4869 (N_4869,N_4750,N_4736);
nand U4870 (N_4870,N_4769,N_4723);
nand U4871 (N_4871,N_4762,N_4709);
xnor U4872 (N_4872,N_4743,N_4700);
nor U4873 (N_4873,N_4712,N_4717);
and U4874 (N_4874,N_4741,N_4725);
nand U4875 (N_4875,N_4702,N_4741);
or U4876 (N_4876,N_4782,N_4774);
and U4877 (N_4877,N_4775,N_4786);
or U4878 (N_4878,N_4755,N_4746);
nand U4879 (N_4879,N_4789,N_4769);
or U4880 (N_4880,N_4706,N_4724);
and U4881 (N_4881,N_4754,N_4755);
nand U4882 (N_4882,N_4719,N_4771);
or U4883 (N_4883,N_4765,N_4725);
nand U4884 (N_4884,N_4792,N_4785);
nor U4885 (N_4885,N_4791,N_4790);
or U4886 (N_4886,N_4765,N_4747);
nor U4887 (N_4887,N_4746,N_4757);
nor U4888 (N_4888,N_4729,N_4792);
or U4889 (N_4889,N_4785,N_4774);
nand U4890 (N_4890,N_4781,N_4716);
nand U4891 (N_4891,N_4734,N_4752);
nor U4892 (N_4892,N_4799,N_4744);
and U4893 (N_4893,N_4779,N_4746);
and U4894 (N_4894,N_4787,N_4714);
or U4895 (N_4895,N_4724,N_4757);
and U4896 (N_4896,N_4735,N_4740);
nor U4897 (N_4897,N_4797,N_4715);
nand U4898 (N_4898,N_4745,N_4785);
nand U4899 (N_4899,N_4704,N_4741);
nor U4900 (N_4900,N_4885,N_4827);
nor U4901 (N_4901,N_4871,N_4877);
and U4902 (N_4902,N_4860,N_4895);
nand U4903 (N_4903,N_4800,N_4846);
nor U4904 (N_4904,N_4893,N_4808);
or U4905 (N_4905,N_4812,N_4855);
nor U4906 (N_4906,N_4844,N_4876);
nand U4907 (N_4907,N_4829,N_4823);
and U4908 (N_4908,N_4804,N_4863);
and U4909 (N_4909,N_4867,N_4887);
or U4910 (N_4910,N_4879,N_4825);
or U4911 (N_4911,N_4837,N_4824);
or U4912 (N_4912,N_4842,N_4833);
or U4913 (N_4913,N_4890,N_4814);
nor U4914 (N_4914,N_4849,N_4832);
nor U4915 (N_4915,N_4852,N_4898);
and U4916 (N_4916,N_4811,N_4892);
and U4917 (N_4917,N_4858,N_4801);
or U4918 (N_4918,N_4822,N_4816);
nand U4919 (N_4919,N_4856,N_4859);
nand U4920 (N_4920,N_4884,N_4882);
nand U4921 (N_4921,N_4853,N_4865);
and U4922 (N_4922,N_4805,N_4843);
nand U4923 (N_4923,N_4813,N_4869);
nand U4924 (N_4924,N_4820,N_4840);
nand U4925 (N_4925,N_4841,N_4817);
and U4926 (N_4926,N_4838,N_4897);
or U4927 (N_4927,N_4815,N_4866);
nand U4928 (N_4928,N_4810,N_4880);
nor U4929 (N_4929,N_4899,N_4872);
or U4930 (N_4930,N_4870,N_4881);
and U4931 (N_4931,N_4836,N_4839);
or U4932 (N_4932,N_4828,N_4864);
and U4933 (N_4933,N_4862,N_4894);
and U4934 (N_4934,N_4873,N_4851);
nor U4935 (N_4935,N_4826,N_4857);
nor U4936 (N_4936,N_4889,N_4821);
or U4937 (N_4937,N_4802,N_4886);
and U4938 (N_4938,N_4809,N_4834);
nand U4939 (N_4939,N_4831,N_4818);
or U4940 (N_4940,N_4819,N_4847);
nand U4941 (N_4941,N_4803,N_4874);
nor U4942 (N_4942,N_4891,N_4878);
nor U4943 (N_4943,N_4883,N_4806);
or U4944 (N_4944,N_4896,N_4868);
nand U4945 (N_4945,N_4861,N_4830);
nand U4946 (N_4946,N_4835,N_4850);
and U4947 (N_4947,N_4888,N_4848);
or U4948 (N_4948,N_4854,N_4845);
nor U4949 (N_4949,N_4875,N_4807);
nor U4950 (N_4950,N_4862,N_4821);
or U4951 (N_4951,N_4856,N_4809);
nand U4952 (N_4952,N_4800,N_4853);
or U4953 (N_4953,N_4803,N_4815);
or U4954 (N_4954,N_4828,N_4880);
nand U4955 (N_4955,N_4811,N_4832);
nand U4956 (N_4956,N_4837,N_4817);
and U4957 (N_4957,N_4801,N_4816);
or U4958 (N_4958,N_4821,N_4863);
nor U4959 (N_4959,N_4897,N_4861);
nand U4960 (N_4960,N_4891,N_4869);
nor U4961 (N_4961,N_4887,N_4816);
or U4962 (N_4962,N_4888,N_4829);
and U4963 (N_4963,N_4837,N_4890);
nor U4964 (N_4964,N_4860,N_4846);
nand U4965 (N_4965,N_4879,N_4876);
nor U4966 (N_4966,N_4898,N_4839);
nand U4967 (N_4967,N_4866,N_4810);
or U4968 (N_4968,N_4895,N_4863);
nand U4969 (N_4969,N_4854,N_4890);
and U4970 (N_4970,N_4883,N_4821);
and U4971 (N_4971,N_4850,N_4843);
or U4972 (N_4972,N_4821,N_4835);
and U4973 (N_4973,N_4832,N_4837);
or U4974 (N_4974,N_4847,N_4852);
nand U4975 (N_4975,N_4804,N_4848);
and U4976 (N_4976,N_4848,N_4829);
and U4977 (N_4977,N_4871,N_4851);
nand U4978 (N_4978,N_4876,N_4828);
nor U4979 (N_4979,N_4881,N_4827);
and U4980 (N_4980,N_4830,N_4845);
or U4981 (N_4981,N_4829,N_4867);
and U4982 (N_4982,N_4810,N_4820);
nand U4983 (N_4983,N_4877,N_4814);
and U4984 (N_4984,N_4893,N_4848);
nor U4985 (N_4985,N_4806,N_4822);
nand U4986 (N_4986,N_4890,N_4849);
and U4987 (N_4987,N_4828,N_4899);
nand U4988 (N_4988,N_4896,N_4889);
or U4989 (N_4989,N_4829,N_4885);
nor U4990 (N_4990,N_4831,N_4829);
and U4991 (N_4991,N_4827,N_4819);
nand U4992 (N_4992,N_4863,N_4823);
nand U4993 (N_4993,N_4857,N_4874);
and U4994 (N_4994,N_4896,N_4803);
or U4995 (N_4995,N_4856,N_4865);
or U4996 (N_4996,N_4861,N_4807);
and U4997 (N_4997,N_4848,N_4815);
nor U4998 (N_4998,N_4843,N_4880);
nor U4999 (N_4999,N_4812,N_4890);
and UO_0 (O_0,N_4991,N_4918);
or UO_1 (O_1,N_4988,N_4930);
nand UO_2 (O_2,N_4999,N_4974);
nor UO_3 (O_3,N_4969,N_4990);
or UO_4 (O_4,N_4929,N_4943);
and UO_5 (O_5,N_4959,N_4958);
and UO_6 (O_6,N_4992,N_4912);
and UO_7 (O_7,N_4942,N_4956);
nand UO_8 (O_8,N_4997,N_4901);
nor UO_9 (O_9,N_4920,N_4963);
and UO_10 (O_10,N_4994,N_4961);
nor UO_11 (O_11,N_4916,N_4939);
nor UO_12 (O_12,N_4950,N_4944);
nand UO_13 (O_13,N_4902,N_4975);
nand UO_14 (O_14,N_4906,N_4970);
nor UO_15 (O_15,N_4957,N_4907);
nor UO_16 (O_16,N_4953,N_4936);
nor UO_17 (O_17,N_4979,N_4987);
nand UO_18 (O_18,N_4993,N_4968);
or UO_19 (O_19,N_4985,N_4927);
nor UO_20 (O_20,N_4980,N_4911);
nor UO_21 (O_21,N_4984,N_4982);
and UO_22 (O_22,N_4938,N_4995);
or UO_23 (O_23,N_4903,N_4908);
or UO_24 (O_24,N_4983,N_4913);
or UO_25 (O_25,N_4949,N_4910);
and UO_26 (O_26,N_4955,N_4914);
nor UO_27 (O_27,N_4946,N_4945);
and UO_28 (O_28,N_4931,N_4965);
or UO_29 (O_29,N_4934,N_4998);
nand UO_30 (O_30,N_4923,N_4917);
or UO_31 (O_31,N_4952,N_4926);
and UO_32 (O_32,N_4937,N_4954);
and UO_33 (O_33,N_4922,N_4977);
nor UO_34 (O_34,N_4935,N_4941);
nand UO_35 (O_35,N_4971,N_4921);
or UO_36 (O_36,N_4948,N_4904);
or UO_37 (O_37,N_4919,N_4976);
nor UO_38 (O_38,N_4915,N_4940);
nor UO_39 (O_39,N_4900,N_4964);
nand UO_40 (O_40,N_4947,N_4932);
and UO_41 (O_41,N_4973,N_4933);
nor UO_42 (O_42,N_4951,N_4962);
or UO_43 (O_43,N_4905,N_4960);
nand UO_44 (O_44,N_4981,N_4978);
or UO_45 (O_45,N_4989,N_4996);
or UO_46 (O_46,N_4972,N_4924);
or UO_47 (O_47,N_4986,N_4909);
nor UO_48 (O_48,N_4928,N_4966);
nor UO_49 (O_49,N_4967,N_4925);
nor UO_50 (O_50,N_4957,N_4997);
or UO_51 (O_51,N_4936,N_4990);
or UO_52 (O_52,N_4974,N_4976);
nor UO_53 (O_53,N_4938,N_4965);
nor UO_54 (O_54,N_4976,N_4963);
nand UO_55 (O_55,N_4930,N_4902);
and UO_56 (O_56,N_4938,N_4941);
nand UO_57 (O_57,N_4968,N_4954);
or UO_58 (O_58,N_4935,N_4904);
or UO_59 (O_59,N_4991,N_4946);
nor UO_60 (O_60,N_4936,N_4987);
and UO_61 (O_61,N_4994,N_4956);
nand UO_62 (O_62,N_4954,N_4911);
nor UO_63 (O_63,N_4927,N_4977);
nand UO_64 (O_64,N_4979,N_4972);
or UO_65 (O_65,N_4909,N_4990);
nor UO_66 (O_66,N_4987,N_4993);
and UO_67 (O_67,N_4946,N_4921);
nor UO_68 (O_68,N_4951,N_4932);
nand UO_69 (O_69,N_4982,N_4926);
nor UO_70 (O_70,N_4952,N_4944);
nand UO_71 (O_71,N_4994,N_4931);
and UO_72 (O_72,N_4907,N_4932);
nor UO_73 (O_73,N_4967,N_4991);
nor UO_74 (O_74,N_4919,N_4914);
xnor UO_75 (O_75,N_4957,N_4928);
nor UO_76 (O_76,N_4975,N_4980);
or UO_77 (O_77,N_4913,N_4979);
and UO_78 (O_78,N_4964,N_4920);
and UO_79 (O_79,N_4926,N_4939);
nor UO_80 (O_80,N_4949,N_4973);
and UO_81 (O_81,N_4997,N_4941);
or UO_82 (O_82,N_4987,N_4914);
or UO_83 (O_83,N_4946,N_4958);
and UO_84 (O_84,N_4987,N_4980);
nor UO_85 (O_85,N_4985,N_4929);
nand UO_86 (O_86,N_4919,N_4913);
or UO_87 (O_87,N_4958,N_4964);
nand UO_88 (O_88,N_4928,N_4942);
and UO_89 (O_89,N_4919,N_4920);
and UO_90 (O_90,N_4950,N_4905);
or UO_91 (O_91,N_4979,N_4918);
nand UO_92 (O_92,N_4930,N_4924);
or UO_93 (O_93,N_4942,N_4959);
nand UO_94 (O_94,N_4902,N_4971);
and UO_95 (O_95,N_4914,N_4915);
nor UO_96 (O_96,N_4982,N_4975);
nor UO_97 (O_97,N_4966,N_4910);
nand UO_98 (O_98,N_4955,N_4900);
or UO_99 (O_99,N_4980,N_4955);
or UO_100 (O_100,N_4908,N_4953);
nor UO_101 (O_101,N_4925,N_4959);
and UO_102 (O_102,N_4909,N_4941);
or UO_103 (O_103,N_4905,N_4902);
and UO_104 (O_104,N_4996,N_4965);
and UO_105 (O_105,N_4940,N_4988);
or UO_106 (O_106,N_4916,N_4915);
nor UO_107 (O_107,N_4990,N_4997);
or UO_108 (O_108,N_4970,N_4923);
or UO_109 (O_109,N_4964,N_4901);
nor UO_110 (O_110,N_4971,N_4931);
nand UO_111 (O_111,N_4990,N_4915);
and UO_112 (O_112,N_4921,N_4935);
nor UO_113 (O_113,N_4925,N_4998);
and UO_114 (O_114,N_4958,N_4986);
nor UO_115 (O_115,N_4994,N_4919);
nand UO_116 (O_116,N_4905,N_4918);
nor UO_117 (O_117,N_4906,N_4902);
nor UO_118 (O_118,N_4934,N_4943);
nand UO_119 (O_119,N_4946,N_4942);
or UO_120 (O_120,N_4965,N_4995);
and UO_121 (O_121,N_4979,N_4948);
or UO_122 (O_122,N_4964,N_4906);
nand UO_123 (O_123,N_4967,N_4972);
or UO_124 (O_124,N_4990,N_4979);
nor UO_125 (O_125,N_4936,N_4926);
or UO_126 (O_126,N_4949,N_4996);
nor UO_127 (O_127,N_4983,N_4923);
nor UO_128 (O_128,N_4933,N_4905);
nor UO_129 (O_129,N_4916,N_4940);
and UO_130 (O_130,N_4991,N_4919);
nor UO_131 (O_131,N_4912,N_4941);
and UO_132 (O_132,N_4922,N_4920);
nand UO_133 (O_133,N_4930,N_4986);
and UO_134 (O_134,N_4993,N_4903);
nand UO_135 (O_135,N_4928,N_4931);
nor UO_136 (O_136,N_4966,N_4912);
and UO_137 (O_137,N_4986,N_4980);
or UO_138 (O_138,N_4980,N_4984);
nand UO_139 (O_139,N_4959,N_4926);
nand UO_140 (O_140,N_4942,N_4902);
or UO_141 (O_141,N_4946,N_4931);
and UO_142 (O_142,N_4996,N_4925);
xnor UO_143 (O_143,N_4905,N_4921);
and UO_144 (O_144,N_4982,N_4970);
or UO_145 (O_145,N_4904,N_4926);
nand UO_146 (O_146,N_4915,N_4907);
nand UO_147 (O_147,N_4940,N_4997);
nand UO_148 (O_148,N_4983,N_4990);
or UO_149 (O_149,N_4972,N_4990);
nor UO_150 (O_150,N_4982,N_4928);
or UO_151 (O_151,N_4912,N_4987);
and UO_152 (O_152,N_4915,N_4999);
and UO_153 (O_153,N_4999,N_4929);
or UO_154 (O_154,N_4948,N_4943);
nor UO_155 (O_155,N_4966,N_4996);
nand UO_156 (O_156,N_4946,N_4979);
or UO_157 (O_157,N_4991,N_4968);
nand UO_158 (O_158,N_4993,N_4905);
or UO_159 (O_159,N_4964,N_4965);
nand UO_160 (O_160,N_4999,N_4925);
nor UO_161 (O_161,N_4989,N_4959);
and UO_162 (O_162,N_4981,N_4934);
nor UO_163 (O_163,N_4996,N_4959);
or UO_164 (O_164,N_4984,N_4939);
and UO_165 (O_165,N_4978,N_4977);
or UO_166 (O_166,N_4945,N_4967);
nand UO_167 (O_167,N_4991,N_4941);
or UO_168 (O_168,N_4954,N_4918);
nor UO_169 (O_169,N_4965,N_4946);
nor UO_170 (O_170,N_4983,N_4927);
and UO_171 (O_171,N_4955,N_4938);
nand UO_172 (O_172,N_4981,N_4941);
or UO_173 (O_173,N_4987,N_4904);
and UO_174 (O_174,N_4900,N_4996);
or UO_175 (O_175,N_4942,N_4905);
and UO_176 (O_176,N_4997,N_4911);
nand UO_177 (O_177,N_4916,N_4953);
and UO_178 (O_178,N_4982,N_4987);
and UO_179 (O_179,N_4924,N_4905);
nand UO_180 (O_180,N_4978,N_4959);
or UO_181 (O_181,N_4921,N_4963);
or UO_182 (O_182,N_4980,N_4970);
nor UO_183 (O_183,N_4925,N_4909);
and UO_184 (O_184,N_4959,N_4973);
or UO_185 (O_185,N_4923,N_4904);
or UO_186 (O_186,N_4929,N_4972);
and UO_187 (O_187,N_4997,N_4924);
or UO_188 (O_188,N_4924,N_4970);
nor UO_189 (O_189,N_4958,N_4915);
or UO_190 (O_190,N_4973,N_4991);
nand UO_191 (O_191,N_4952,N_4969);
or UO_192 (O_192,N_4932,N_4999);
and UO_193 (O_193,N_4911,N_4991);
nor UO_194 (O_194,N_4971,N_4910);
nand UO_195 (O_195,N_4909,N_4997);
nor UO_196 (O_196,N_4972,N_4976);
nand UO_197 (O_197,N_4928,N_4993);
and UO_198 (O_198,N_4963,N_4900);
nor UO_199 (O_199,N_4953,N_4919);
or UO_200 (O_200,N_4939,N_4907);
and UO_201 (O_201,N_4982,N_4978);
or UO_202 (O_202,N_4968,N_4950);
nand UO_203 (O_203,N_4921,N_4998);
xor UO_204 (O_204,N_4979,N_4949);
nor UO_205 (O_205,N_4944,N_4943);
nor UO_206 (O_206,N_4928,N_4930);
nand UO_207 (O_207,N_4907,N_4998);
and UO_208 (O_208,N_4982,N_4946);
or UO_209 (O_209,N_4947,N_4993);
or UO_210 (O_210,N_4997,N_4982);
and UO_211 (O_211,N_4944,N_4954);
nand UO_212 (O_212,N_4952,N_4989);
nor UO_213 (O_213,N_4989,N_4904);
and UO_214 (O_214,N_4909,N_4955);
and UO_215 (O_215,N_4900,N_4946);
nand UO_216 (O_216,N_4906,N_4981);
or UO_217 (O_217,N_4995,N_4934);
nand UO_218 (O_218,N_4919,N_4931);
nor UO_219 (O_219,N_4977,N_4905);
or UO_220 (O_220,N_4989,N_4910);
nand UO_221 (O_221,N_4920,N_4948);
and UO_222 (O_222,N_4957,N_4999);
nand UO_223 (O_223,N_4916,N_4961);
nand UO_224 (O_224,N_4949,N_4938);
and UO_225 (O_225,N_4901,N_4914);
and UO_226 (O_226,N_4988,N_4924);
nor UO_227 (O_227,N_4920,N_4914);
nor UO_228 (O_228,N_4954,N_4949);
or UO_229 (O_229,N_4970,N_4908);
or UO_230 (O_230,N_4925,N_4910);
nand UO_231 (O_231,N_4957,N_4918);
nand UO_232 (O_232,N_4903,N_4911);
nand UO_233 (O_233,N_4982,N_4945);
and UO_234 (O_234,N_4954,N_4973);
and UO_235 (O_235,N_4902,N_4908);
nand UO_236 (O_236,N_4996,N_4921);
and UO_237 (O_237,N_4952,N_4930);
or UO_238 (O_238,N_4943,N_4976);
nand UO_239 (O_239,N_4975,N_4904);
nand UO_240 (O_240,N_4970,N_4946);
nor UO_241 (O_241,N_4958,N_4910);
nor UO_242 (O_242,N_4965,N_4993);
or UO_243 (O_243,N_4999,N_4997);
nor UO_244 (O_244,N_4986,N_4933);
nor UO_245 (O_245,N_4903,N_4996);
or UO_246 (O_246,N_4921,N_4976);
and UO_247 (O_247,N_4950,N_4918);
and UO_248 (O_248,N_4936,N_4966);
nor UO_249 (O_249,N_4958,N_4948);
nand UO_250 (O_250,N_4922,N_4930);
and UO_251 (O_251,N_4978,N_4906);
xor UO_252 (O_252,N_4989,N_4997);
nor UO_253 (O_253,N_4987,N_4952);
and UO_254 (O_254,N_4979,N_4966);
or UO_255 (O_255,N_4952,N_4951);
and UO_256 (O_256,N_4972,N_4938);
and UO_257 (O_257,N_4949,N_4930);
and UO_258 (O_258,N_4995,N_4931);
nand UO_259 (O_259,N_4956,N_4925);
and UO_260 (O_260,N_4969,N_4920);
or UO_261 (O_261,N_4963,N_4966);
nor UO_262 (O_262,N_4983,N_4974);
nand UO_263 (O_263,N_4913,N_4912);
or UO_264 (O_264,N_4926,N_4965);
nor UO_265 (O_265,N_4934,N_4950);
and UO_266 (O_266,N_4992,N_4953);
or UO_267 (O_267,N_4970,N_4936);
nor UO_268 (O_268,N_4959,N_4998);
and UO_269 (O_269,N_4995,N_4990);
and UO_270 (O_270,N_4941,N_4944);
and UO_271 (O_271,N_4958,N_4967);
or UO_272 (O_272,N_4904,N_4985);
or UO_273 (O_273,N_4991,N_4985);
nor UO_274 (O_274,N_4902,N_4910);
nand UO_275 (O_275,N_4990,N_4974);
nand UO_276 (O_276,N_4905,N_4947);
or UO_277 (O_277,N_4983,N_4997);
and UO_278 (O_278,N_4904,N_4945);
or UO_279 (O_279,N_4908,N_4992);
nor UO_280 (O_280,N_4930,N_4906);
or UO_281 (O_281,N_4940,N_4966);
nor UO_282 (O_282,N_4940,N_4926);
nand UO_283 (O_283,N_4930,N_4926);
or UO_284 (O_284,N_4961,N_4978);
or UO_285 (O_285,N_4959,N_4993);
or UO_286 (O_286,N_4935,N_4973);
or UO_287 (O_287,N_4943,N_4945);
or UO_288 (O_288,N_4955,N_4969);
nor UO_289 (O_289,N_4960,N_4930);
nor UO_290 (O_290,N_4939,N_4981);
nand UO_291 (O_291,N_4908,N_4976);
or UO_292 (O_292,N_4945,N_4912);
or UO_293 (O_293,N_4990,N_4941);
nand UO_294 (O_294,N_4936,N_4937);
nand UO_295 (O_295,N_4917,N_4913);
or UO_296 (O_296,N_4900,N_4925);
nand UO_297 (O_297,N_4984,N_4900);
or UO_298 (O_298,N_4946,N_4987);
nand UO_299 (O_299,N_4999,N_4901);
or UO_300 (O_300,N_4945,N_4953);
and UO_301 (O_301,N_4959,N_4951);
nand UO_302 (O_302,N_4913,N_4916);
or UO_303 (O_303,N_4950,N_4949);
or UO_304 (O_304,N_4936,N_4956);
nand UO_305 (O_305,N_4926,N_4948);
nor UO_306 (O_306,N_4991,N_4960);
or UO_307 (O_307,N_4960,N_4947);
xor UO_308 (O_308,N_4952,N_4901);
or UO_309 (O_309,N_4999,N_4917);
or UO_310 (O_310,N_4900,N_4942);
nand UO_311 (O_311,N_4974,N_4948);
and UO_312 (O_312,N_4951,N_4999);
nor UO_313 (O_313,N_4905,N_4994);
nand UO_314 (O_314,N_4965,N_4921);
nor UO_315 (O_315,N_4947,N_4913);
nand UO_316 (O_316,N_4907,N_4917);
nand UO_317 (O_317,N_4911,N_4970);
and UO_318 (O_318,N_4998,N_4946);
nor UO_319 (O_319,N_4954,N_4962);
nand UO_320 (O_320,N_4941,N_4965);
nor UO_321 (O_321,N_4928,N_4919);
and UO_322 (O_322,N_4941,N_4946);
nand UO_323 (O_323,N_4929,N_4954);
nand UO_324 (O_324,N_4999,N_4960);
and UO_325 (O_325,N_4911,N_4956);
nor UO_326 (O_326,N_4943,N_4922);
and UO_327 (O_327,N_4972,N_4952);
or UO_328 (O_328,N_4947,N_4956);
or UO_329 (O_329,N_4989,N_4980);
nor UO_330 (O_330,N_4947,N_4912);
nand UO_331 (O_331,N_4924,N_4931);
nand UO_332 (O_332,N_4966,N_4952);
and UO_333 (O_333,N_4967,N_4992);
nand UO_334 (O_334,N_4971,N_4957);
nor UO_335 (O_335,N_4994,N_4930);
nor UO_336 (O_336,N_4979,N_4902);
and UO_337 (O_337,N_4928,N_4911);
nand UO_338 (O_338,N_4956,N_4907);
nand UO_339 (O_339,N_4928,N_4940);
and UO_340 (O_340,N_4913,N_4971);
and UO_341 (O_341,N_4903,N_4970);
and UO_342 (O_342,N_4995,N_4948);
and UO_343 (O_343,N_4967,N_4960);
or UO_344 (O_344,N_4913,N_4900);
nor UO_345 (O_345,N_4904,N_4972);
nor UO_346 (O_346,N_4945,N_4989);
or UO_347 (O_347,N_4958,N_4935);
and UO_348 (O_348,N_4986,N_4988);
nor UO_349 (O_349,N_4951,N_4998);
or UO_350 (O_350,N_4906,N_4997);
nand UO_351 (O_351,N_4929,N_4915);
and UO_352 (O_352,N_4965,N_4939);
or UO_353 (O_353,N_4927,N_4938);
nand UO_354 (O_354,N_4922,N_4923);
and UO_355 (O_355,N_4939,N_4944);
xnor UO_356 (O_356,N_4915,N_4964);
or UO_357 (O_357,N_4986,N_4995);
and UO_358 (O_358,N_4921,N_4930);
nor UO_359 (O_359,N_4993,N_4973);
nor UO_360 (O_360,N_4996,N_4992);
nand UO_361 (O_361,N_4939,N_4948);
nand UO_362 (O_362,N_4953,N_4949);
or UO_363 (O_363,N_4958,N_4975);
nor UO_364 (O_364,N_4980,N_4967);
and UO_365 (O_365,N_4932,N_4968);
or UO_366 (O_366,N_4946,N_4966);
and UO_367 (O_367,N_4904,N_4966);
nand UO_368 (O_368,N_4941,N_4970);
nand UO_369 (O_369,N_4949,N_4969);
nor UO_370 (O_370,N_4996,N_4945);
or UO_371 (O_371,N_4947,N_4930);
nand UO_372 (O_372,N_4981,N_4904);
and UO_373 (O_373,N_4970,N_4991);
nor UO_374 (O_374,N_4940,N_4990);
or UO_375 (O_375,N_4912,N_4978);
and UO_376 (O_376,N_4989,N_4926);
nor UO_377 (O_377,N_4920,N_4917);
nand UO_378 (O_378,N_4915,N_4920);
and UO_379 (O_379,N_4903,N_4945);
or UO_380 (O_380,N_4905,N_4901);
nand UO_381 (O_381,N_4940,N_4976);
nor UO_382 (O_382,N_4978,N_4952);
or UO_383 (O_383,N_4984,N_4968);
nor UO_384 (O_384,N_4936,N_4962);
nand UO_385 (O_385,N_4961,N_4999);
or UO_386 (O_386,N_4925,N_4997);
and UO_387 (O_387,N_4933,N_4971);
nand UO_388 (O_388,N_4999,N_4904);
or UO_389 (O_389,N_4907,N_4965);
and UO_390 (O_390,N_4910,N_4930);
nor UO_391 (O_391,N_4985,N_4992);
nor UO_392 (O_392,N_4911,N_4906);
nand UO_393 (O_393,N_4960,N_4954);
and UO_394 (O_394,N_4914,N_4908);
nand UO_395 (O_395,N_4923,N_4933);
xor UO_396 (O_396,N_4998,N_4960);
nor UO_397 (O_397,N_4925,N_4912);
nor UO_398 (O_398,N_4962,N_4923);
xnor UO_399 (O_399,N_4973,N_4906);
nand UO_400 (O_400,N_4923,N_4979);
nand UO_401 (O_401,N_4938,N_4997);
and UO_402 (O_402,N_4957,N_4931);
nand UO_403 (O_403,N_4971,N_4904);
nor UO_404 (O_404,N_4969,N_4925);
and UO_405 (O_405,N_4920,N_4977);
nand UO_406 (O_406,N_4998,N_4949);
nand UO_407 (O_407,N_4920,N_4916);
nor UO_408 (O_408,N_4962,N_4965);
or UO_409 (O_409,N_4926,N_4990);
nand UO_410 (O_410,N_4927,N_4996);
nand UO_411 (O_411,N_4934,N_4965);
nand UO_412 (O_412,N_4998,N_4932);
nor UO_413 (O_413,N_4973,N_4932);
or UO_414 (O_414,N_4977,N_4993);
or UO_415 (O_415,N_4968,N_4974);
or UO_416 (O_416,N_4917,N_4947);
nand UO_417 (O_417,N_4958,N_4911);
and UO_418 (O_418,N_4957,N_4908);
and UO_419 (O_419,N_4987,N_4991);
nor UO_420 (O_420,N_4952,N_4924);
nand UO_421 (O_421,N_4995,N_4909);
or UO_422 (O_422,N_4929,N_4982);
and UO_423 (O_423,N_4927,N_4940);
nor UO_424 (O_424,N_4906,N_4992);
nand UO_425 (O_425,N_4923,N_4941);
nor UO_426 (O_426,N_4956,N_4905);
nand UO_427 (O_427,N_4913,N_4960);
nand UO_428 (O_428,N_4972,N_4957);
or UO_429 (O_429,N_4932,N_4925);
nor UO_430 (O_430,N_4912,N_4934);
nand UO_431 (O_431,N_4910,N_4953);
or UO_432 (O_432,N_4901,N_4911);
and UO_433 (O_433,N_4906,N_4972);
and UO_434 (O_434,N_4910,N_4923);
nand UO_435 (O_435,N_4952,N_4932);
and UO_436 (O_436,N_4957,N_4914);
and UO_437 (O_437,N_4908,N_4935);
nor UO_438 (O_438,N_4925,N_4960);
or UO_439 (O_439,N_4966,N_4961);
or UO_440 (O_440,N_4967,N_4995);
or UO_441 (O_441,N_4918,N_4937);
and UO_442 (O_442,N_4977,N_4956);
and UO_443 (O_443,N_4988,N_4933);
nand UO_444 (O_444,N_4911,N_4961);
nand UO_445 (O_445,N_4905,N_4900);
and UO_446 (O_446,N_4962,N_4944);
nand UO_447 (O_447,N_4970,N_4967);
nor UO_448 (O_448,N_4979,N_4991);
and UO_449 (O_449,N_4944,N_4916);
nor UO_450 (O_450,N_4922,N_4968);
or UO_451 (O_451,N_4946,N_4944);
and UO_452 (O_452,N_4957,N_4923);
nand UO_453 (O_453,N_4922,N_4904);
nand UO_454 (O_454,N_4978,N_4939);
nand UO_455 (O_455,N_4933,N_4951);
and UO_456 (O_456,N_4900,N_4981);
and UO_457 (O_457,N_4921,N_4952);
nand UO_458 (O_458,N_4912,N_4997);
nand UO_459 (O_459,N_4979,N_4994);
and UO_460 (O_460,N_4922,N_4919);
nand UO_461 (O_461,N_4903,N_4913);
xnor UO_462 (O_462,N_4936,N_4996);
nor UO_463 (O_463,N_4900,N_4965);
and UO_464 (O_464,N_4981,N_4976);
and UO_465 (O_465,N_4975,N_4908);
nor UO_466 (O_466,N_4993,N_4920);
nor UO_467 (O_467,N_4912,N_4938);
and UO_468 (O_468,N_4944,N_4989);
or UO_469 (O_469,N_4992,N_4955);
or UO_470 (O_470,N_4915,N_4998);
nor UO_471 (O_471,N_4937,N_4947);
or UO_472 (O_472,N_4956,N_4986);
nand UO_473 (O_473,N_4910,N_4941);
nand UO_474 (O_474,N_4976,N_4932);
nor UO_475 (O_475,N_4976,N_4993);
and UO_476 (O_476,N_4902,N_4901);
xnor UO_477 (O_477,N_4961,N_4912);
nor UO_478 (O_478,N_4969,N_4940);
and UO_479 (O_479,N_4968,N_4918);
or UO_480 (O_480,N_4902,N_4935);
or UO_481 (O_481,N_4943,N_4931);
and UO_482 (O_482,N_4918,N_4942);
or UO_483 (O_483,N_4925,N_4905);
or UO_484 (O_484,N_4971,N_4942);
nor UO_485 (O_485,N_4923,N_4989);
nand UO_486 (O_486,N_4951,N_4901);
nor UO_487 (O_487,N_4943,N_4952);
nand UO_488 (O_488,N_4909,N_4956);
and UO_489 (O_489,N_4954,N_4902);
nand UO_490 (O_490,N_4923,N_4931);
nor UO_491 (O_491,N_4955,N_4978);
nand UO_492 (O_492,N_4918,N_4909);
nor UO_493 (O_493,N_4950,N_4936);
nor UO_494 (O_494,N_4982,N_4902);
and UO_495 (O_495,N_4960,N_4922);
nand UO_496 (O_496,N_4964,N_4935);
and UO_497 (O_497,N_4905,N_4996);
or UO_498 (O_498,N_4947,N_4948);
and UO_499 (O_499,N_4931,N_4930);
and UO_500 (O_500,N_4948,N_4906);
and UO_501 (O_501,N_4964,N_4954);
and UO_502 (O_502,N_4908,N_4964);
and UO_503 (O_503,N_4923,N_4993);
and UO_504 (O_504,N_4925,N_4987);
nand UO_505 (O_505,N_4905,N_4991);
nor UO_506 (O_506,N_4945,N_4963);
or UO_507 (O_507,N_4910,N_4901);
or UO_508 (O_508,N_4960,N_4958);
nand UO_509 (O_509,N_4992,N_4994);
nand UO_510 (O_510,N_4937,N_4929);
or UO_511 (O_511,N_4983,N_4940);
nand UO_512 (O_512,N_4951,N_4956);
or UO_513 (O_513,N_4927,N_4916);
and UO_514 (O_514,N_4955,N_4993);
and UO_515 (O_515,N_4947,N_4967);
nor UO_516 (O_516,N_4909,N_4991);
or UO_517 (O_517,N_4991,N_4996);
and UO_518 (O_518,N_4993,N_4992);
nor UO_519 (O_519,N_4932,N_4978);
nand UO_520 (O_520,N_4930,N_4942);
and UO_521 (O_521,N_4947,N_4970);
nor UO_522 (O_522,N_4950,N_4945);
nor UO_523 (O_523,N_4965,N_4913);
nor UO_524 (O_524,N_4986,N_4950);
or UO_525 (O_525,N_4977,N_4968);
and UO_526 (O_526,N_4999,N_4972);
or UO_527 (O_527,N_4993,N_4943);
or UO_528 (O_528,N_4929,N_4953);
and UO_529 (O_529,N_4935,N_4929);
and UO_530 (O_530,N_4928,N_4913);
or UO_531 (O_531,N_4989,N_4947);
nor UO_532 (O_532,N_4935,N_4910);
nor UO_533 (O_533,N_4927,N_4937);
nand UO_534 (O_534,N_4927,N_4967);
nand UO_535 (O_535,N_4990,N_4900);
nand UO_536 (O_536,N_4936,N_4910);
nand UO_537 (O_537,N_4944,N_4923);
nor UO_538 (O_538,N_4974,N_4975);
or UO_539 (O_539,N_4926,N_4996);
nand UO_540 (O_540,N_4945,N_4983);
or UO_541 (O_541,N_4933,N_4942);
and UO_542 (O_542,N_4940,N_4996);
or UO_543 (O_543,N_4998,N_4953);
nand UO_544 (O_544,N_4990,N_4967);
nor UO_545 (O_545,N_4977,N_4932);
and UO_546 (O_546,N_4979,N_4962);
nand UO_547 (O_547,N_4902,N_4928);
and UO_548 (O_548,N_4961,N_4931);
nor UO_549 (O_549,N_4940,N_4945);
nor UO_550 (O_550,N_4976,N_4918);
or UO_551 (O_551,N_4924,N_4939);
or UO_552 (O_552,N_4933,N_4987);
and UO_553 (O_553,N_4998,N_4928);
and UO_554 (O_554,N_4999,N_4941);
nand UO_555 (O_555,N_4936,N_4982);
nor UO_556 (O_556,N_4950,N_4966);
and UO_557 (O_557,N_4911,N_4993);
and UO_558 (O_558,N_4946,N_4968);
nand UO_559 (O_559,N_4907,N_4912);
and UO_560 (O_560,N_4939,N_4992);
or UO_561 (O_561,N_4944,N_4958);
nand UO_562 (O_562,N_4941,N_4950);
or UO_563 (O_563,N_4906,N_4996);
nand UO_564 (O_564,N_4938,N_4998);
nor UO_565 (O_565,N_4934,N_4991);
nor UO_566 (O_566,N_4914,N_4900);
and UO_567 (O_567,N_4927,N_4972);
and UO_568 (O_568,N_4962,N_4976);
and UO_569 (O_569,N_4989,N_4999);
nand UO_570 (O_570,N_4907,N_4931);
nand UO_571 (O_571,N_4905,N_4930);
xor UO_572 (O_572,N_4999,N_4981);
nand UO_573 (O_573,N_4993,N_4950);
or UO_574 (O_574,N_4930,N_4935);
nand UO_575 (O_575,N_4991,N_4964);
or UO_576 (O_576,N_4928,N_4901);
or UO_577 (O_577,N_4921,N_4908);
or UO_578 (O_578,N_4929,N_4942);
nor UO_579 (O_579,N_4967,N_4966);
or UO_580 (O_580,N_4958,N_4924);
nor UO_581 (O_581,N_4930,N_4944);
or UO_582 (O_582,N_4997,N_4910);
and UO_583 (O_583,N_4933,N_4925);
nor UO_584 (O_584,N_4942,N_4920);
and UO_585 (O_585,N_4946,N_4925);
nand UO_586 (O_586,N_4930,N_4998);
or UO_587 (O_587,N_4982,N_4923);
or UO_588 (O_588,N_4992,N_4981);
nand UO_589 (O_589,N_4915,N_4973);
or UO_590 (O_590,N_4922,N_4952);
or UO_591 (O_591,N_4947,N_4976);
nand UO_592 (O_592,N_4987,N_4900);
nor UO_593 (O_593,N_4918,N_4952);
and UO_594 (O_594,N_4931,N_4996);
nor UO_595 (O_595,N_4936,N_4932);
nor UO_596 (O_596,N_4997,N_4936);
or UO_597 (O_597,N_4986,N_4920);
and UO_598 (O_598,N_4937,N_4945);
or UO_599 (O_599,N_4950,N_4997);
and UO_600 (O_600,N_4986,N_4948);
nand UO_601 (O_601,N_4986,N_4993);
and UO_602 (O_602,N_4985,N_4957);
or UO_603 (O_603,N_4967,N_4986);
and UO_604 (O_604,N_4995,N_4944);
nor UO_605 (O_605,N_4971,N_4987);
or UO_606 (O_606,N_4966,N_4938);
nor UO_607 (O_607,N_4966,N_4905);
nand UO_608 (O_608,N_4999,N_4906);
or UO_609 (O_609,N_4935,N_4946);
or UO_610 (O_610,N_4930,N_4948);
and UO_611 (O_611,N_4934,N_4986);
nor UO_612 (O_612,N_4994,N_4921);
and UO_613 (O_613,N_4995,N_4975);
and UO_614 (O_614,N_4937,N_4941);
nor UO_615 (O_615,N_4939,N_4943);
nor UO_616 (O_616,N_4994,N_4960);
and UO_617 (O_617,N_4906,N_4982);
nor UO_618 (O_618,N_4923,N_4996);
nand UO_619 (O_619,N_4977,N_4992);
or UO_620 (O_620,N_4972,N_4959);
and UO_621 (O_621,N_4953,N_4948);
nand UO_622 (O_622,N_4929,N_4958);
nor UO_623 (O_623,N_4956,N_4962);
and UO_624 (O_624,N_4935,N_4955);
or UO_625 (O_625,N_4941,N_4960);
and UO_626 (O_626,N_4916,N_4948);
nand UO_627 (O_627,N_4912,N_4914);
nor UO_628 (O_628,N_4918,N_4906);
or UO_629 (O_629,N_4977,N_4933);
or UO_630 (O_630,N_4948,N_4942);
and UO_631 (O_631,N_4925,N_4923);
or UO_632 (O_632,N_4979,N_4934);
or UO_633 (O_633,N_4910,N_4988);
nor UO_634 (O_634,N_4917,N_4971);
or UO_635 (O_635,N_4975,N_4927);
or UO_636 (O_636,N_4967,N_4944);
or UO_637 (O_637,N_4979,N_4974);
and UO_638 (O_638,N_4994,N_4917);
nor UO_639 (O_639,N_4969,N_4903);
or UO_640 (O_640,N_4927,N_4962);
and UO_641 (O_641,N_4986,N_4987);
and UO_642 (O_642,N_4965,N_4933);
or UO_643 (O_643,N_4935,N_4967);
or UO_644 (O_644,N_4940,N_4949);
nand UO_645 (O_645,N_4984,N_4927);
nor UO_646 (O_646,N_4982,N_4992);
and UO_647 (O_647,N_4901,N_4944);
or UO_648 (O_648,N_4929,N_4917);
nor UO_649 (O_649,N_4977,N_4944);
nor UO_650 (O_650,N_4975,N_4965);
and UO_651 (O_651,N_4924,N_4998);
nor UO_652 (O_652,N_4981,N_4972);
and UO_653 (O_653,N_4979,N_4999);
and UO_654 (O_654,N_4983,N_4905);
nor UO_655 (O_655,N_4967,N_4929);
and UO_656 (O_656,N_4907,N_4964);
and UO_657 (O_657,N_4972,N_4998);
or UO_658 (O_658,N_4911,N_4960);
and UO_659 (O_659,N_4942,N_4931);
nor UO_660 (O_660,N_4901,N_4946);
or UO_661 (O_661,N_4942,N_4995);
or UO_662 (O_662,N_4983,N_4937);
or UO_663 (O_663,N_4950,N_4969);
and UO_664 (O_664,N_4983,N_4910);
nand UO_665 (O_665,N_4937,N_4987);
or UO_666 (O_666,N_4969,N_4986);
nor UO_667 (O_667,N_4911,N_4973);
or UO_668 (O_668,N_4939,N_4977);
nand UO_669 (O_669,N_4980,N_4925);
nor UO_670 (O_670,N_4914,N_4974);
and UO_671 (O_671,N_4970,N_4918);
or UO_672 (O_672,N_4902,N_4963);
nand UO_673 (O_673,N_4987,N_4940);
nor UO_674 (O_674,N_4994,N_4942);
or UO_675 (O_675,N_4982,N_4990);
and UO_676 (O_676,N_4970,N_4939);
nand UO_677 (O_677,N_4992,N_4917);
nor UO_678 (O_678,N_4915,N_4962);
nor UO_679 (O_679,N_4955,N_4999);
nand UO_680 (O_680,N_4955,N_4923);
or UO_681 (O_681,N_4912,N_4932);
nand UO_682 (O_682,N_4990,N_4980);
nand UO_683 (O_683,N_4919,N_4904);
or UO_684 (O_684,N_4950,N_4984);
and UO_685 (O_685,N_4999,N_4982);
or UO_686 (O_686,N_4937,N_4905);
nor UO_687 (O_687,N_4953,N_4931);
nand UO_688 (O_688,N_4910,N_4911);
and UO_689 (O_689,N_4941,N_4939);
or UO_690 (O_690,N_4969,N_4931);
nor UO_691 (O_691,N_4995,N_4989);
nand UO_692 (O_692,N_4954,N_4994);
nand UO_693 (O_693,N_4902,N_4923);
and UO_694 (O_694,N_4943,N_4991);
or UO_695 (O_695,N_4908,N_4973);
nor UO_696 (O_696,N_4958,N_4982);
or UO_697 (O_697,N_4941,N_4966);
xnor UO_698 (O_698,N_4957,N_4994);
nor UO_699 (O_699,N_4936,N_4933);
or UO_700 (O_700,N_4932,N_4904);
nand UO_701 (O_701,N_4990,N_4999);
nand UO_702 (O_702,N_4905,N_4910);
nor UO_703 (O_703,N_4951,N_4964);
nand UO_704 (O_704,N_4952,N_4970);
or UO_705 (O_705,N_4945,N_4969);
nor UO_706 (O_706,N_4991,N_4924);
nand UO_707 (O_707,N_4911,N_4925);
nor UO_708 (O_708,N_4978,N_4902);
nand UO_709 (O_709,N_4932,N_4960);
and UO_710 (O_710,N_4944,N_4927);
and UO_711 (O_711,N_4991,N_4998);
nor UO_712 (O_712,N_4987,N_4998);
nor UO_713 (O_713,N_4952,N_4903);
nor UO_714 (O_714,N_4922,N_4961);
and UO_715 (O_715,N_4928,N_4933);
nor UO_716 (O_716,N_4912,N_4929);
or UO_717 (O_717,N_4930,N_4987);
nand UO_718 (O_718,N_4961,N_4930);
or UO_719 (O_719,N_4977,N_4900);
nand UO_720 (O_720,N_4955,N_4966);
or UO_721 (O_721,N_4946,N_4972);
nor UO_722 (O_722,N_4976,N_4906);
nor UO_723 (O_723,N_4983,N_4960);
nand UO_724 (O_724,N_4996,N_4975);
and UO_725 (O_725,N_4980,N_4971);
and UO_726 (O_726,N_4950,N_4989);
nor UO_727 (O_727,N_4955,N_4944);
nor UO_728 (O_728,N_4905,N_4969);
nor UO_729 (O_729,N_4966,N_4960);
or UO_730 (O_730,N_4919,N_4988);
nor UO_731 (O_731,N_4924,N_4951);
and UO_732 (O_732,N_4986,N_4964);
or UO_733 (O_733,N_4965,N_4909);
nand UO_734 (O_734,N_4979,N_4908);
nor UO_735 (O_735,N_4982,N_4967);
or UO_736 (O_736,N_4978,N_4909);
nand UO_737 (O_737,N_4950,N_4922);
or UO_738 (O_738,N_4911,N_4994);
and UO_739 (O_739,N_4941,N_4969);
or UO_740 (O_740,N_4908,N_4967);
nor UO_741 (O_741,N_4912,N_4943);
and UO_742 (O_742,N_4909,N_4971);
and UO_743 (O_743,N_4975,N_4986);
and UO_744 (O_744,N_4900,N_4948);
nand UO_745 (O_745,N_4945,N_4935);
nand UO_746 (O_746,N_4950,N_4970);
and UO_747 (O_747,N_4970,N_4977);
and UO_748 (O_748,N_4927,N_4917);
or UO_749 (O_749,N_4918,N_4958);
nand UO_750 (O_750,N_4952,N_4958);
nor UO_751 (O_751,N_4962,N_4933);
or UO_752 (O_752,N_4924,N_4935);
nand UO_753 (O_753,N_4935,N_4983);
nor UO_754 (O_754,N_4978,N_4995);
or UO_755 (O_755,N_4966,N_4915);
nor UO_756 (O_756,N_4989,N_4902);
or UO_757 (O_757,N_4942,N_4952);
nand UO_758 (O_758,N_4903,N_4959);
xor UO_759 (O_759,N_4986,N_4951);
xor UO_760 (O_760,N_4922,N_4932);
or UO_761 (O_761,N_4934,N_4988);
or UO_762 (O_762,N_4947,N_4996);
or UO_763 (O_763,N_4919,N_4942);
nand UO_764 (O_764,N_4996,N_4962);
nor UO_765 (O_765,N_4948,N_4981);
nand UO_766 (O_766,N_4910,N_4979);
and UO_767 (O_767,N_4992,N_4902);
nand UO_768 (O_768,N_4903,N_4947);
nand UO_769 (O_769,N_4927,N_4988);
nor UO_770 (O_770,N_4972,N_4920);
nor UO_771 (O_771,N_4997,N_4918);
nand UO_772 (O_772,N_4904,N_4939);
or UO_773 (O_773,N_4904,N_4988);
or UO_774 (O_774,N_4996,N_4980);
xor UO_775 (O_775,N_4980,N_4981);
or UO_776 (O_776,N_4924,N_4979);
and UO_777 (O_777,N_4991,N_4957);
nand UO_778 (O_778,N_4945,N_4991);
or UO_779 (O_779,N_4912,N_4917);
or UO_780 (O_780,N_4971,N_4958);
and UO_781 (O_781,N_4929,N_4923);
xor UO_782 (O_782,N_4903,N_4975);
nor UO_783 (O_783,N_4938,N_4971);
nor UO_784 (O_784,N_4912,N_4982);
nand UO_785 (O_785,N_4997,N_4915);
nand UO_786 (O_786,N_4970,N_4996);
or UO_787 (O_787,N_4900,N_4967);
nand UO_788 (O_788,N_4914,N_4972);
or UO_789 (O_789,N_4942,N_4947);
or UO_790 (O_790,N_4904,N_4908);
or UO_791 (O_791,N_4907,N_4992);
nand UO_792 (O_792,N_4926,N_4942);
nand UO_793 (O_793,N_4999,N_4958);
nor UO_794 (O_794,N_4922,N_4937);
nand UO_795 (O_795,N_4924,N_4964);
or UO_796 (O_796,N_4902,N_4996);
nand UO_797 (O_797,N_4974,N_4959);
nor UO_798 (O_798,N_4970,N_4926);
nand UO_799 (O_799,N_4971,N_4990);
or UO_800 (O_800,N_4923,N_4940);
and UO_801 (O_801,N_4928,N_4996);
and UO_802 (O_802,N_4949,N_4985);
nand UO_803 (O_803,N_4958,N_4934);
nor UO_804 (O_804,N_4925,N_4962);
and UO_805 (O_805,N_4943,N_4969);
and UO_806 (O_806,N_4980,N_4928);
nor UO_807 (O_807,N_4999,N_4968);
or UO_808 (O_808,N_4929,N_4977);
and UO_809 (O_809,N_4919,N_4944);
nand UO_810 (O_810,N_4953,N_4902);
nor UO_811 (O_811,N_4976,N_4951);
nor UO_812 (O_812,N_4932,N_4994);
and UO_813 (O_813,N_4937,N_4925);
nand UO_814 (O_814,N_4968,N_4928);
and UO_815 (O_815,N_4995,N_4902);
nand UO_816 (O_816,N_4915,N_4950);
nor UO_817 (O_817,N_4956,N_4967);
and UO_818 (O_818,N_4949,N_4936);
or UO_819 (O_819,N_4990,N_4916);
or UO_820 (O_820,N_4988,N_4950);
or UO_821 (O_821,N_4966,N_4927);
or UO_822 (O_822,N_4916,N_4925);
or UO_823 (O_823,N_4927,N_4943);
nand UO_824 (O_824,N_4967,N_4902);
and UO_825 (O_825,N_4916,N_4967);
and UO_826 (O_826,N_4915,N_4980);
nor UO_827 (O_827,N_4960,N_4986);
nor UO_828 (O_828,N_4945,N_4998);
nand UO_829 (O_829,N_4965,N_4977);
and UO_830 (O_830,N_4984,N_4985);
nor UO_831 (O_831,N_4925,N_4904);
nor UO_832 (O_832,N_4947,N_4936);
nand UO_833 (O_833,N_4919,N_4957);
and UO_834 (O_834,N_4908,N_4966);
or UO_835 (O_835,N_4970,N_4973);
and UO_836 (O_836,N_4958,N_4961);
nand UO_837 (O_837,N_4989,N_4948);
or UO_838 (O_838,N_4918,N_4962);
nand UO_839 (O_839,N_4962,N_4992);
or UO_840 (O_840,N_4964,N_4975);
or UO_841 (O_841,N_4969,N_4989);
nor UO_842 (O_842,N_4949,N_4989);
nand UO_843 (O_843,N_4996,N_4993);
or UO_844 (O_844,N_4925,N_4942);
nor UO_845 (O_845,N_4910,N_4965);
and UO_846 (O_846,N_4907,N_4988);
nor UO_847 (O_847,N_4990,N_4987);
nand UO_848 (O_848,N_4950,N_4932);
nand UO_849 (O_849,N_4981,N_4932);
or UO_850 (O_850,N_4988,N_4941);
nand UO_851 (O_851,N_4982,N_4914);
or UO_852 (O_852,N_4979,N_4982);
and UO_853 (O_853,N_4966,N_4994);
nor UO_854 (O_854,N_4939,N_4983);
nor UO_855 (O_855,N_4967,N_4948);
and UO_856 (O_856,N_4909,N_4908);
nand UO_857 (O_857,N_4931,N_4936);
and UO_858 (O_858,N_4957,N_4992);
and UO_859 (O_859,N_4984,N_4960);
and UO_860 (O_860,N_4928,N_4958);
or UO_861 (O_861,N_4901,N_4977);
nand UO_862 (O_862,N_4918,N_4987);
and UO_863 (O_863,N_4973,N_4947);
or UO_864 (O_864,N_4963,N_4958);
nor UO_865 (O_865,N_4953,N_4980);
nor UO_866 (O_866,N_4969,N_4917);
or UO_867 (O_867,N_4986,N_4984);
nand UO_868 (O_868,N_4993,N_4989);
nand UO_869 (O_869,N_4965,N_4994);
and UO_870 (O_870,N_4980,N_4995);
and UO_871 (O_871,N_4988,N_4901);
or UO_872 (O_872,N_4960,N_4924);
nand UO_873 (O_873,N_4959,N_4971);
or UO_874 (O_874,N_4950,N_4979);
and UO_875 (O_875,N_4934,N_4932);
and UO_876 (O_876,N_4939,N_4999);
nand UO_877 (O_877,N_4926,N_4973);
or UO_878 (O_878,N_4963,N_4983);
nand UO_879 (O_879,N_4909,N_4933);
nand UO_880 (O_880,N_4938,N_4954);
nor UO_881 (O_881,N_4901,N_4993);
nand UO_882 (O_882,N_4944,N_4921);
nor UO_883 (O_883,N_4974,N_4981);
and UO_884 (O_884,N_4922,N_4966);
or UO_885 (O_885,N_4943,N_4900);
nand UO_886 (O_886,N_4992,N_4923);
nand UO_887 (O_887,N_4936,N_4902);
or UO_888 (O_888,N_4967,N_4976);
nor UO_889 (O_889,N_4931,N_4977);
or UO_890 (O_890,N_4909,N_4983);
nand UO_891 (O_891,N_4979,N_4917);
nor UO_892 (O_892,N_4950,N_4953);
and UO_893 (O_893,N_4978,N_4927);
and UO_894 (O_894,N_4953,N_4918);
nand UO_895 (O_895,N_4998,N_4906);
or UO_896 (O_896,N_4977,N_4980);
and UO_897 (O_897,N_4948,N_4918);
nand UO_898 (O_898,N_4937,N_4902);
nand UO_899 (O_899,N_4987,N_4975);
nor UO_900 (O_900,N_4926,N_4955);
nand UO_901 (O_901,N_4976,N_4933);
nand UO_902 (O_902,N_4961,N_4918);
nand UO_903 (O_903,N_4921,N_4949);
or UO_904 (O_904,N_4955,N_4910);
nor UO_905 (O_905,N_4954,N_4920);
or UO_906 (O_906,N_4914,N_4956);
and UO_907 (O_907,N_4967,N_4924);
nand UO_908 (O_908,N_4923,N_4907);
or UO_909 (O_909,N_4989,N_4960);
or UO_910 (O_910,N_4949,N_4971);
nor UO_911 (O_911,N_4981,N_4961);
or UO_912 (O_912,N_4946,N_4922);
nor UO_913 (O_913,N_4929,N_4957);
nand UO_914 (O_914,N_4948,N_4977);
nand UO_915 (O_915,N_4904,N_4953);
nor UO_916 (O_916,N_4925,N_4995);
or UO_917 (O_917,N_4952,N_4986);
nor UO_918 (O_918,N_4960,N_4916);
nor UO_919 (O_919,N_4901,N_4926);
nor UO_920 (O_920,N_4954,N_4905);
nand UO_921 (O_921,N_4939,N_4998);
and UO_922 (O_922,N_4983,N_4914);
nand UO_923 (O_923,N_4951,N_4938);
nor UO_924 (O_924,N_4951,N_4980);
nand UO_925 (O_925,N_4907,N_4948);
or UO_926 (O_926,N_4918,N_4917);
nand UO_927 (O_927,N_4976,N_4924);
nand UO_928 (O_928,N_4931,N_4976);
and UO_929 (O_929,N_4945,N_4933);
nand UO_930 (O_930,N_4993,N_4907);
or UO_931 (O_931,N_4995,N_4920);
nand UO_932 (O_932,N_4948,N_4994);
nand UO_933 (O_933,N_4981,N_4928);
nor UO_934 (O_934,N_4923,N_4945);
nand UO_935 (O_935,N_4955,N_4928);
nand UO_936 (O_936,N_4934,N_4928);
or UO_937 (O_937,N_4959,N_4985);
and UO_938 (O_938,N_4983,N_4976);
or UO_939 (O_939,N_4967,N_4978);
nor UO_940 (O_940,N_4961,N_4977);
or UO_941 (O_941,N_4918,N_4931);
or UO_942 (O_942,N_4980,N_4939);
nand UO_943 (O_943,N_4969,N_4924);
nand UO_944 (O_944,N_4947,N_4985);
nor UO_945 (O_945,N_4984,N_4943);
or UO_946 (O_946,N_4994,N_4927);
nor UO_947 (O_947,N_4990,N_4945);
nand UO_948 (O_948,N_4986,N_4976);
and UO_949 (O_949,N_4912,N_4952);
nor UO_950 (O_950,N_4997,N_4931);
nand UO_951 (O_951,N_4964,N_4992);
or UO_952 (O_952,N_4992,N_4931);
nor UO_953 (O_953,N_4988,N_4951);
and UO_954 (O_954,N_4910,N_4994);
or UO_955 (O_955,N_4966,N_4985);
or UO_956 (O_956,N_4937,N_4990);
nand UO_957 (O_957,N_4902,N_4993);
and UO_958 (O_958,N_4962,N_4999);
or UO_959 (O_959,N_4958,N_4981);
and UO_960 (O_960,N_4931,N_4970);
nand UO_961 (O_961,N_4941,N_4901);
nor UO_962 (O_962,N_4947,N_4925);
or UO_963 (O_963,N_4948,N_4917);
nand UO_964 (O_964,N_4982,N_4913);
and UO_965 (O_965,N_4944,N_4932);
nand UO_966 (O_966,N_4949,N_4900);
or UO_967 (O_967,N_4901,N_4976);
nand UO_968 (O_968,N_4998,N_4943);
nand UO_969 (O_969,N_4923,N_4906);
and UO_970 (O_970,N_4934,N_4983);
or UO_971 (O_971,N_4907,N_4978);
nor UO_972 (O_972,N_4904,N_4978);
or UO_973 (O_973,N_4942,N_4911);
or UO_974 (O_974,N_4913,N_4985);
nor UO_975 (O_975,N_4950,N_4907);
and UO_976 (O_976,N_4963,N_4922);
and UO_977 (O_977,N_4940,N_4956);
and UO_978 (O_978,N_4985,N_4962);
or UO_979 (O_979,N_4962,N_4977);
and UO_980 (O_980,N_4910,N_4928);
nand UO_981 (O_981,N_4935,N_4907);
nor UO_982 (O_982,N_4989,N_4931);
and UO_983 (O_983,N_4902,N_4950);
nand UO_984 (O_984,N_4953,N_4909);
and UO_985 (O_985,N_4942,N_4954);
or UO_986 (O_986,N_4961,N_4990);
and UO_987 (O_987,N_4984,N_4988);
nand UO_988 (O_988,N_4932,N_4987);
nor UO_989 (O_989,N_4939,N_4919);
nor UO_990 (O_990,N_4997,N_4933);
and UO_991 (O_991,N_4995,N_4947);
nor UO_992 (O_992,N_4955,N_4972);
nand UO_993 (O_993,N_4929,N_4995);
or UO_994 (O_994,N_4924,N_4925);
or UO_995 (O_995,N_4995,N_4954);
nand UO_996 (O_996,N_4940,N_4900);
nand UO_997 (O_997,N_4903,N_4921);
and UO_998 (O_998,N_4973,N_4957);
or UO_999 (O_999,N_4982,N_4976);
endmodule