module basic_500_3000_500_40_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_200,In_416);
nor U1 (N_1,In_226,In_456);
or U2 (N_2,In_453,In_219);
nand U3 (N_3,In_38,In_155);
or U4 (N_4,In_498,In_477);
or U5 (N_5,In_344,In_339);
and U6 (N_6,In_111,In_83);
nor U7 (N_7,In_136,In_444);
or U8 (N_8,In_249,In_142);
or U9 (N_9,In_326,In_228);
and U10 (N_10,In_215,In_399);
and U11 (N_11,In_189,In_379);
and U12 (N_12,In_359,In_352);
or U13 (N_13,In_293,In_295);
xnor U14 (N_14,In_311,In_66);
nand U15 (N_15,In_166,In_121);
and U16 (N_16,In_402,In_482);
or U17 (N_17,In_6,In_169);
and U18 (N_18,In_92,In_120);
or U19 (N_19,In_467,In_139);
or U20 (N_20,In_350,In_179);
and U21 (N_21,In_408,In_97);
or U22 (N_22,In_99,In_318);
and U23 (N_23,In_167,In_255);
xnor U24 (N_24,In_263,In_476);
or U25 (N_25,In_440,In_17);
or U26 (N_26,In_433,In_390);
and U27 (N_27,In_406,In_48);
nor U28 (N_28,In_144,In_306);
or U29 (N_29,In_42,In_397);
and U30 (N_30,In_487,In_108);
and U31 (N_31,In_439,In_22);
nand U32 (N_32,In_158,In_472);
xnor U33 (N_33,In_53,In_71);
nor U34 (N_34,In_239,In_63);
or U35 (N_35,In_361,In_259);
and U36 (N_36,In_58,In_109);
nand U37 (N_37,In_0,In_330);
nand U38 (N_38,In_128,In_74);
nand U39 (N_39,In_199,In_130);
nand U40 (N_40,In_65,In_165);
nor U41 (N_41,In_320,In_377);
nand U42 (N_42,In_140,In_192);
nand U43 (N_43,In_395,In_428);
or U44 (N_44,In_355,In_91);
and U45 (N_45,In_151,In_314);
nand U46 (N_46,In_378,In_281);
nor U47 (N_47,In_368,In_25);
or U48 (N_48,In_322,In_360);
or U49 (N_49,In_59,In_298);
nor U50 (N_50,In_449,In_491);
nor U51 (N_51,In_362,In_429);
or U52 (N_52,In_105,In_160);
or U53 (N_53,In_224,In_60);
nor U54 (N_54,In_329,In_427);
and U55 (N_55,In_405,In_264);
and U56 (N_56,In_177,In_44);
and U57 (N_57,In_431,In_82);
and U58 (N_58,In_371,In_443);
xnor U59 (N_59,In_323,In_162);
nor U60 (N_60,In_212,In_117);
xor U61 (N_61,In_262,In_244);
and U62 (N_62,In_183,In_240);
nand U63 (N_63,In_430,In_208);
or U64 (N_64,In_229,In_287);
and U65 (N_65,In_29,In_37);
or U66 (N_66,In_21,In_277);
nor U67 (N_67,In_119,In_319);
and U68 (N_68,In_210,In_247);
and U69 (N_69,In_424,In_363);
nor U70 (N_70,In_204,In_354);
and U71 (N_71,In_332,In_389);
nand U72 (N_72,In_253,In_450);
and U73 (N_73,In_129,In_358);
xor U74 (N_74,In_468,In_241);
nor U75 (N_75,In_297,In_296);
or U76 (N_76,In_370,In_180);
or U77 (N_77,In_112,In_341);
and U78 (N_78,In_470,N_58);
nand U79 (N_79,In_9,In_267);
nand U80 (N_80,In_385,In_150);
or U81 (N_81,In_205,In_118);
nand U82 (N_82,In_421,In_134);
and U83 (N_83,N_31,In_410);
xnor U84 (N_84,N_14,N_71);
nor U85 (N_85,In_356,In_43);
and U86 (N_86,In_452,In_24);
nand U87 (N_87,In_492,In_373);
xor U88 (N_88,In_475,In_245);
or U89 (N_89,In_81,In_425);
and U90 (N_90,N_37,In_233);
nand U91 (N_91,N_74,In_79);
nand U92 (N_92,In_11,In_309);
or U93 (N_93,In_214,N_4);
nor U94 (N_94,In_87,In_412);
nor U95 (N_95,N_16,In_176);
and U96 (N_96,In_266,In_488);
xor U97 (N_97,N_24,In_174);
or U98 (N_98,N_72,In_156);
xor U99 (N_99,In_13,In_55);
nor U100 (N_100,In_54,In_102);
nand U101 (N_101,In_455,In_321);
nor U102 (N_102,In_481,In_451);
nand U103 (N_103,N_21,N_1);
or U104 (N_104,In_380,N_35);
nor U105 (N_105,In_432,In_294);
and U106 (N_106,In_232,In_497);
and U107 (N_107,In_8,In_260);
nand U108 (N_108,N_3,In_300);
nor U109 (N_109,In_152,N_68);
xor U110 (N_110,In_195,N_0);
and U111 (N_111,In_357,In_334);
nor U112 (N_112,In_122,In_178);
nor U113 (N_113,In_285,In_434);
nand U114 (N_114,In_51,In_206);
nand U115 (N_115,In_252,N_61);
nand U116 (N_116,In_175,In_374);
or U117 (N_117,In_459,In_191);
xnor U118 (N_118,In_442,In_248);
or U119 (N_119,In_254,In_190);
and U120 (N_120,In_69,In_127);
nand U121 (N_121,In_203,In_324);
or U122 (N_122,N_36,In_448);
or U123 (N_123,In_35,In_84);
or U124 (N_124,In_495,In_85);
nor U125 (N_125,In_230,In_317);
nor U126 (N_126,In_251,In_426);
xnor U127 (N_127,In_49,In_225);
nand U128 (N_128,In_499,In_146);
or U129 (N_129,In_202,In_496);
or U130 (N_130,In_172,In_145);
or U131 (N_131,In_479,In_327);
nor U132 (N_132,In_26,In_164);
or U133 (N_133,In_315,In_486);
nor U134 (N_134,In_336,In_394);
nand U135 (N_135,In_471,In_286);
nand U136 (N_136,In_170,In_305);
or U137 (N_137,In_473,N_66);
or U138 (N_138,N_12,In_391);
nand U139 (N_139,N_53,In_265);
nor U140 (N_140,In_269,N_64);
nand U141 (N_141,In_2,In_104);
and U142 (N_142,In_422,In_173);
nand U143 (N_143,In_159,In_365);
and U144 (N_144,N_52,In_367);
xnor U145 (N_145,In_77,N_19);
nand U146 (N_146,N_7,In_388);
and U147 (N_147,In_52,In_36);
and U148 (N_148,In_168,In_401);
xnor U149 (N_149,In_282,N_10);
nor U150 (N_150,In_125,In_141);
and U151 (N_151,In_96,In_4);
xnor U152 (N_152,In_88,In_438);
or U153 (N_153,In_218,In_40);
nor U154 (N_154,N_75,N_138);
and U155 (N_155,In_147,In_484);
and U156 (N_156,N_85,In_46);
nor U157 (N_157,In_15,In_221);
nand U158 (N_158,N_69,N_121);
nand U159 (N_159,In_485,N_45);
and U160 (N_160,N_63,N_57);
nor U161 (N_161,In_338,In_86);
and U162 (N_162,In_135,N_77);
and U163 (N_163,In_236,N_43);
nor U164 (N_164,In_103,N_82);
nand U165 (N_165,In_291,N_5);
xor U166 (N_166,N_131,In_364);
or U167 (N_167,In_303,In_19);
or U168 (N_168,In_101,In_187);
or U169 (N_169,In_369,N_41);
or U170 (N_170,In_123,In_268);
nor U171 (N_171,N_100,N_144);
or U172 (N_172,In_20,In_131);
and U173 (N_173,In_217,In_474);
nor U174 (N_174,In_447,N_46);
and U175 (N_175,In_478,In_489);
or U176 (N_176,In_256,N_129);
xor U177 (N_177,In_372,N_112);
and U178 (N_178,N_29,In_290);
or U179 (N_179,N_11,N_38);
nor U180 (N_180,In_308,In_93);
nand U181 (N_181,N_143,In_325);
and U182 (N_182,In_400,In_387);
nand U183 (N_183,In_494,N_70);
or U184 (N_184,In_28,N_107);
nand U185 (N_185,In_14,In_386);
and U186 (N_186,In_465,In_301);
nand U187 (N_187,N_39,N_104);
nand U188 (N_188,In_279,N_106);
nand U189 (N_189,N_9,N_92);
nor U190 (N_190,In_89,In_348);
nand U191 (N_191,In_64,N_98);
xor U192 (N_192,In_246,In_132);
and U193 (N_193,In_415,In_220);
and U194 (N_194,N_113,In_148);
and U195 (N_195,N_108,In_67);
nand U196 (N_196,N_67,In_154);
and U197 (N_197,In_39,N_27);
or U198 (N_198,In_342,In_61);
and U199 (N_199,In_107,In_292);
or U200 (N_200,In_276,In_95);
nor U201 (N_201,N_90,N_116);
nand U202 (N_202,In_331,In_198);
or U203 (N_203,N_51,In_403);
or U204 (N_204,N_60,In_345);
and U205 (N_205,N_125,In_445);
nand U206 (N_206,In_437,In_454);
and U207 (N_207,N_49,In_222);
nand U208 (N_208,In_157,N_149);
nand U209 (N_209,In_413,In_392);
or U210 (N_210,In_273,In_261);
xnor U211 (N_211,N_91,N_79);
nor U212 (N_212,In_31,In_423);
nand U213 (N_213,In_181,In_258);
nor U214 (N_214,In_68,N_62);
nor U215 (N_215,In_409,N_2);
xnor U216 (N_216,N_54,In_435);
nor U217 (N_217,N_132,In_76);
nand U218 (N_218,N_147,N_118);
xor U219 (N_219,In_126,In_124);
nor U220 (N_220,N_15,In_113);
or U221 (N_221,N_23,In_404);
and U222 (N_222,In_275,In_312);
and U223 (N_223,N_33,N_50);
nor U224 (N_224,In_419,N_42);
nand U225 (N_225,N_181,In_223);
or U226 (N_226,In_393,N_169);
or U227 (N_227,In_70,In_185);
or U228 (N_228,N_22,In_90);
xnor U229 (N_229,N_219,N_222);
nand U230 (N_230,In_384,N_223);
and U231 (N_231,N_95,N_28);
xnor U232 (N_232,In_75,N_93);
nand U233 (N_233,In_464,In_231);
and U234 (N_234,N_44,In_271);
and U235 (N_235,N_142,In_243);
xnor U236 (N_236,N_190,In_80);
or U237 (N_237,N_220,In_196);
or U238 (N_238,N_154,In_62);
and U239 (N_239,In_283,In_349);
nand U240 (N_240,In_33,N_188);
nand U241 (N_241,In_73,In_313);
or U242 (N_242,N_160,In_493);
nand U243 (N_243,N_99,In_272);
or U244 (N_244,In_184,In_34);
nand U245 (N_245,N_172,In_110);
or U246 (N_246,N_195,In_418);
nor U247 (N_247,N_101,N_193);
and U248 (N_248,In_227,N_161);
nor U249 (N_249,In_396,N_192);
or U250 (N_250,N_207,N_141);
nand U251 (N_251,N_212,N_55);
and U252 (N_252,N_133,N_215);
and U253 (N_253,N_156,In_299);
or U254 (N_254,In_375,In_420);
xnor U255 (N_255,In_257,N_196);
and U256 (N_256,In_337,In_436);
or U257 (N_257,N_174,N_189);
nand U258 (N_258,In_138,N_206);
and U259 (N_259,N_185,N_165);
nor U260 (N_260,N_56,In_161);
nor U261 (N_261,In_56,In_289);
nor U262 (N_262,N_202,N_86);
nor U263 (N_263,N_30,In_483);
nor U264 (N_264,N_199,In_316);
and U265 (N_265,N_48,N_32);
nand U266 (N_266,N_187,In_366);
nor U267 (N_267,N_153,In_16);
nor U268 (N_268,N_217,In_284);
xor U269 (N_269,N_216,N_155);
xor U270 (N_270,N_73,N_123);
xnor U271 (N_271,In_333,In_12);
or U272 (N_272,In_351,N_186);
or U273 (N_273,N_211,N_105);
and U274 (N_274,N_115,N_8);
nor U275 (N_275,In_188,In_194);
nor U276 (N_276,In_57,N_183);
nand U277 (N_277,In_328,N_184);
or U278 (N_278,In_201,In_411);
and U279 (N_279,N_148,In_250);
nand U280 (N_280,In_376,N_159);
or U281 (N_281,N_168,In_417);
and U282 (N_282,N_162,In_30);
and U283 (N_283,In_462,In_398);
or U284 (N_284,N_170,In_274);
or U285 (N_285,In_280,In_211);
nand U286 (N_286,N_109,N_18);
or U287 (N_287,N_25,N_146);
nand U288 (N_288,In_458,N_114);
or U289 (N_289,In_463,N_103);
nand U290 (N_290,In_98,In_45);
or U291 (N_291,In_213,N_150);
and U292 (N_292,In_461,N_175);
nand U293 (N_293,In_480,In_114);
nor U294 (N_294,N_47,N_179);
or U295 (N_295,N_164,In_27);
and U296 (N_296,N_81,N_145);
nand U297 (N_297,In_94,N_124);
nor U298 (N_298,N_40,N_180);
and U299 (N_299,N_191,N_102);
and U300 (N_300,N_97,In_143);
nor U301 (N_301,N_285,N_229);
or U302 (N_302,In_182,N_279);
xor U303 (N_303,N_271,In_381);
and U304 (N_304,N_203,N_194);
nor U305 (N_305,N_6,N_96);
nor U306 (N_306,N_259,N_126);
nand U307 (N_307,N_287,N_260);
and U308 (N_308,In_441,N_237);
and U309 (N_309,In_346,N_83);
or U310 (N_310,N_134,N_252);
nand U311 (N_311,N_228,N_230);
and U312 (N_312,In_207,In_353);
nor U313 (N_313,N_238,N_200);
nor U314 (N_314,N_110,N_78);
nor U315 (N_315,N_264,N_34);
xor U316 (N_316,N_111,N_163);
nor U317 (N_317,N_17,In_78);
nor U318 (N_318,In_23,N_282);
or U319 (N_319,In_304,N_139);
xor U320 (N_320,In_234,N_177);
and U321 (N_321,N_234,N_270);
or U322 (N_322,N_299,N_210);
or U323 (N_323,In_133,In_446);
and U324 (N_324,N_89,In_469);
xnor U325 (N_325,N_233,N_209);
nor U326 (N_326,N_136,In_193);
nand U327 (N_327,N_262,N_280);
or U328 (N_328,In_238,N_213);
and U329 (N_329,N_135,N_128);
nor U330 (N_330,N_88,N_13);
nand U331 (N_331,In_50,In_197);
nor U332 (N_332,N_140,N_295);
and U333 (N_333,In_3,N_267);
or U334 (N_334,N_269,N_65);
nand U335 (N_335,N_275,N_218);
nor U336 (N_336,N_243,N_281);
or U337 (N_337,In_163,N_20);
nor U338 (N_338,N_253,In_47);
xor U339 (N_339,N_261,In_343);
and U340 (N_340,N_152,In_5);
or U341 (N_341,In_335,In_115);
or U342 (N_342,In_237,N_289);
or U343 (N_343,In_288,In_307);
and U344 (N_344,N_257,N_266);
or U345 (N_345,N_130,N_122);
nor U346 (N_346,In_7,In_10);
nor U347 (N_347,N_176,N_278);
nor U348 (N_348,N_80,N_297);
or U349 (N_349,N_208,In_32);
nor U350 (N_350,In_347,N_221);
nand U351 (N_351,N_178,N_248);
nor U352 (N_352,N_250,In_466);
nand U353 (N_353,N_294,N_205);
xnor U354 (N_354,N_227,N_249);
and U355 (N_355,N_242,In_186);
nor U356 (N_356,N_268,N_226);
or U357 (N_357,N_265,In_414);
and U358 (N_358,N_277,N_76);
nand U359 (N_359,N_235,N_231);
nor U360 (N_360,In_490,N_236);
nor U361 (N_361,N_84,N_263);
xor U362 (N_362,In_382,In_457);
nor U363 (N_363,N_166,N_288);
or U364 (N_364,In_137,In_383);
nand U365 (N_365,N_284,N_225);
xor U366 (N_366,N_151,N_232);
nor U367 (N_367,N_201,In_149);
nand U368 (N_368,In_242,N_120);
nor U369 (N_369,N_198,N_296);
xor U370 (N_370,In_209,N_167);
or U371 (N_371,N_182,N_239);
and U372 (N_372,N_276,N_256);
nor U373 (N_373,N_117,N_26);
and U374 (N_374,N_283,In_340);
nor U375 (N_375,N_247,N_127);
and U376 (N_376,N_246,N_347);
nand U377 (N_377,N_366,In_310);
nor U378 (N_378,N_292,N_358);
xor U379 (N_379,N_300,N_274);
nand U380 (N_380,N_311,N_309);
or U381 (N_381,N_371,N_312);
and U382 (N_382,N_330,N_331);
and U383 (N_383,N_369,N_272);
nand U384 (N_384,N_338,N_362);
nand U385 (N_385,N_350,N_316);
or U386 (N_386,N_351,In_1);
nor U387 (N_387,N_334,N_204);
nand U388 (N_388,N_214,N_304);
or U389 (N_389,N_329,N_359);
nor U390 (N_390,N_322,N_245);
xor U391 (N_391,N_372,N_321);
and U392 (N_392,N_290,N_361);
nor U393 (N_393,N_87,N_326);
nor U394 (N_394,N_332,N_333);
or U395 (N_395,N_293,N_306);
xor U396 (N_396,N_314,N_119);
and U397 (N_397,N_173,N_258);
or U398 (N_398,N_313,In_116);
nor U399 (N_399,N_224,N_303);
nand U400 (N_400,In_153,In_216);
and U401 (N_401,N_318,N_373);
nand U402 (N_402,N_357,N_251);
or U403 (N_403,In_106,N_368);
nand U404 (N_404,N_370,In_18);
or U405 (N_405,N_345,N_374);
nand U406 (N_406,N_336,N_360);
nand U407 (N_407,N_328,In_460);
or U408 (N_408,N_348,N_137);
nor U409 (N_409,N_291,N_254);
nand U410 (N_410,In_100,N_353);
xor U411 (N_411,N_324,N_341);
nand U412 (N_412,N_244,N_327);
or U413 (N_413,N_302,N_157);
and U414 (N_414,N_356,N_339);
nor U415 (N_415,N_363,In_302);
xnor U416 (N_416,N_241,In_72);
nand U417 (N_417,N_342,N_367);
nand U418 (N_418,In_407,N_337);
nor U419 (N_419,In_171,N_171);
and U420 (N_420,In_235,N_197);
or U421 (N_421,N_307,N_301);
nor U422 (N_422,N_317,N_335);
and U423 (N_423,In_41,N_325);
or U424 (N_424,N_94,N_310);
or U425 (N_425,N_308,N_355);
or U426 (N_426,N_340,N_346);
nand U427 (N_427,In_278,N_365);
xnor U428 (N_428,N_352,N_323);
or U429 (N_429,N_349,N_59);
or U430 (N_430,N_158,N_240);
nand U431 (N_431,In_270,N_298);
xnor U432 (N_432,N_305,N_273);
nor U433 (N_433,N_319,N_286);
or U434 (N_434,N_364,N_343);
or U435 (N_435,N_255,N_344);
and U436 (N_436,N_315,N_354);
and U437 (N_437,N_320,N_303);
nand U438 (N_438,N_251,N_367);
and U439 (N_439,N_247,N_333);
and U440 (N_440,N_240,N_59);
or U441 (N_441,N_244,N_307);
xnor U442 (N_442,N_292,N_255);
nor U443 (N_443,N_274,In_270);
or U444 (N_444,N_312,N_359);
nor U445 (N_445,N_321,N_325);
nand U446 (N_446,N_347,N_171);
and U447 (N_447,N_308,N_137);
nand U448 (N_448,In_407,N_331);
and U449 (N_449,N_254,N_342);
or U450 (N_450,N_394,N_396);
or U451 (N_451,N_433,N_399);
and U452 (N_452,N_384,N_431);
and U453 (N_453,N_402,N_424);
and U454 (N_454,N_391,N_422);
nand U455 (N_455,N_395,N_436);
nand U456 (N_456,N_388,N_447);
and U457 (N_457,N_393,N_430);
and U458 (N_458,N_442,N_387);
and U459 (N_459,N_380,N_412);
nand U460 (N_460,N_385,N_437);
nand U461 (N_461,N_416,N_443);
nor U462 (N_462,N_407,N_413);
or U463 (N_463,N_409,N_420);
nand U464 (N_464,N_401,N_434);
or U465 (N_465,N_421,N_445);
and U466 (N_466,N_432,N_418);
or U467 (N_467,N_446,N_379);
nand U468 (N_468,N_405,N_441);
and U469 (N_469,N_398,N_435);
nand U470 (N_470,N_392,N_414);
and U471 (N_471,N_415,N_417);
nor U472 (N_472,N_444,N_438);
nor U473 (N_473,N_448,N_429);
or U474 (N_474,N_377,N_404);
xor U475 (N_475,N_419,N_386);
nor U476 (N_476,N_411,N_449);
nand U477 (N_477,N_423,N_390);
xnor U478 (N_478,N_400,N_375);
nor U479 (N_479,N_378,N_406);
nor U480 (N_480,N_428,N_426);
and U481 (N_481,N_425,N_383);
and U482 (N_482,N_427,N_440);
and U483 (N_483,N_376,N_397);
and U484 (N_484,N_410,N_408);
nor U485 (N_485,N_403,N_381);
nand U486 (N_486,N_389,N_382);
and U487 (N_487,N_439,N_421);
nand U488 (N_488,N_386,N_389);
or U489 (N_489,N_438,N_422);
nor U490 (N_490,N_424,N_425);
nor U491 (N_491,N_416,N_377);
nor U492 (N_492,N_423,N_409);
or U493 (N_493,N_428,N_424);
xnor U494 (N_494,N_383,N_423);
nand U495 (N_495,N_438,N_418);
nor U496 (N_496,N_389,N_421);
xor U497 (N_497,N_383,N_419);
nand U498 (N_498,N_390,N_396);
nor U499 (N_499,N_426,N_430);
xor U500 (N_500,N_395,N_430);
nand U501 (N_501,N_446,N_449);
xnor U502 (N_502,N_400,N_379);
and U503 (N_503,N_417,N_444);
or U504 (N_504,N_437,N_449);
and U505 (N_505,N_429,N_433);
and U506 (N_506,N_395,N_384);
and U507 (N_507,N_405,N_391);
nand U508 (N_508,N_377,N_413);
xor U509 (N_509,N_447,N_415);
nand U510 (N_510,N_423,N_429);
nor U511 (N_511,N_418,N_379);
nor U512 (N_512,N_399,N_397);
or U513 (N_513,N_422,N_405);
and U514 (N_514,N_416,N_417);
and U515 (N_515,N_439,N_441);
xnor U516 (N_516,N_430,N_434);
nand U517 (N_517,N_408,N_448);
nor U518 (N_518,N_442,N_430);
and U519 (N_519,N_380,N_393);
and U520 (N_520,N_419,N_438);
or U521 (N_521,N_435,N_427);
or U522 (N_522,N_396,N_433);
nand U523 (N_523,N_427,N_418);
nand U524 (N_524,N_394,N_432);
xnor U525 (N_525,N_507,N_499);
nand U526 (N_526,N_472,N_479);
and U527 (N_527,N_469,N_503);
and U528 (N_528,N_463,N_504);
and U529 (N_529,N_518,N_495);
or U530 (N_530,N_462,N_466);
or U531 (N_531,N_467,N_522);
or U532 (N_532,N_454,N_509);
and U533 (N_533,N_490,N_451);
nor U534 (N_534,N_452,N_457);
nor U535 (N_535,N_482,N_506);
and U536 (N_536,N_481,N_465);
nor U537 (N_537,N_480,N_510);
or U538 (N_538,N_513,N_470);
nor U539 (N_539,N_502,N_515);
and U540 (N_540,N_520,N_468);
nand U541 (N_541,N_521,N_488);
and U542 (N_542,N_475,N_471);
nor U543 (N_543,N_459,N_456);
and U544 (N_544,N_516,N_501);
or U545 (N_545,N_476,N_455);
and U546 (N_546,N_460,N_492);
nand U547 (N_547,N_489,N_500);
nand U548 (N_548,N_493,N_523);
nor U549 (N_549,N_483,N_458);
or U550 (N_550,N_519,N_496);
nor U551 (N_551,N_494,N_491);
or U552 (N_552,N_524,N_485);
or U553 (N_553,N_473,N_464);
nand U554 (N_554,N_508,N_514);
and U555 (N_555,N_505,N_450);
or U556 (N_556,N_497,N_474);
nor U557 (N_557,N_478,N_453);
nor U558 (N_558,N_486,N_511);
and U559 (N_559,N_484,N_477);
nor U560 (N_560,N_498,N_461);
and U561 (N_561,N_512,N_517);
nand U562 (N_562,N_487,N_464);
and U563 (N_563,N_504,N_464);
nand U564 (N_564,N_514,N_505);
nand U565 (N_565,N_482,N_454);
or U566 (N_566,N_454,N_498);
or U567 (N_567,N_498,N_506);
or U568 (N_568,N_480,N_475);
and U569 (N_569,N_465,N_508);
nor U570 (N_570,N_502,N_521);
nor U571 (N_571,N_509,N_517);
nor U572 (N_572,N_481,N_503);
and U573 (N_573,N_456,N_505);
or U574 (N_574,N_460,N_500);
nor U575 (N_575,N_517,N_481);
and U576 (N_576,N_517,N_467);
xor U577 (N_577,N_496,N_516);
xnor U578 (N_578,N_471,N_488);
and U579 (N_579,N_457,N_516);
xor U580 (N_580,N_459,N_500);
nor U581 (N_581,N_471,N_490);
or U582 (N_582,N_517,N_471);
and U583 (N_583,N_468,N_504);
nand U584 (N_584,N_461,N_451);
nor U585 (N_585,N_497,N_471);
and U586 (N_586,N_491,N_511);
xnor U587 (N_587,N_455,N_451);
and U588 (N_588,N_511,N_476);
xor U589 (N_589,N_476,N_510);
or U590 (N_590,N_467,N_476);
or U591 (N_591,N_494,N_518);
nand U592 (N_592,N_472,N_492);
nor U593 (N_593,N_515,N_463);
nor U594 (N_594,N_520,N_469);
nand U595 (N_595,N_459,N_484);
nor U596 (N_596,N_462,N_510);
nand U597 (N_597,N_474,N_450);
nor U598 (N_598,N_474,N_462);
nor U599 (N_599,N_490,N_456);
nor U600 (N_600,N_534,N_548);
or U601 (N_601,N_561,N_567);
nor U602 (N_602,N_588,N_595);
or U603 (N_603,N_525,N_569);
or U604 (N_604,N_560,N_555);
nor U605 (N_605,N_593,N_584);
nand U606 (N_606,N_591,N_592);
nor U607 (N_607,N_558,N_598);
nor U608 (N_608,N_532,N_559);
nand U609 (N_609,N_544,N_570);
nand U610 (N_610,N_550,N_541);
or U611 (N_611,N_554,N_576);
xnor U612 (N_612,N_585,N_538);
nand U613 (N_613,N_553,N_527);
nor U614 (N_614,N_552,N_589);
nor U615 (N_615,N_542,N_529);
nor U616 (N_616,N_531,N_545);
nor U617 (N_617,N_571,N_535);
or U618 (N_618,N_547,N_574);
and U619 (N_619,N_594,N_581);
nor U620 (N_620,N_580,N_572);
and U621 (N_621,N_590,N_546);
xnor U622 (N_622,N_562,N_573);
or U623 (N_623,N_556,N_533);
or U624 (N_624,N_596,N_579);
and U625 (N_625,N_549,N_597);
and U626 (N_626,N_566,N_575);
and U627 (N_627,N_563,N_539);
xor U628 (N_628,N_586,N_557);
nand U629 (N_629,N_537,N_583);
or U630 (N_630,N_564,N_551);
xnor U631 (N_631,N_565,N_582);
or U632 (N_632,N_568,N_578);
xnor U633 (N_633,N_577,N_528);
nor U634 (N_634,N_540,N_530);
nor U635 (N_635,N_536,N_543);
or U636 (N_636,N_599,N_587);
nand U637 (N_637,N_526,N_551);
and U638 (N_638,N_568,N_583);
and U639 (N_639,N_535,N_578);
and U640 (N_640,N_543,N_591);
or U641 (N_641,N_543,N_559);
nor U642 (N_642,N_543,N_561);
and U643 (N_643,N_556,N_528);
and U644 (N_644,N_553,N_526);
or U645 (N_645,N_554,N_542);
nand U646 (N_646,N_578,N_585);
nor U647 (N_647,N_588,N_593);
or U648 (N_648,N_599,N_567);
nand U649 (N_649,N_556,N_552);
nand U650 (N_650,N_599,N_591);
nand U651 (N_651,N_565,N_563);
or U652 (N_652,N_581,N_545);
and U653 (N_653,N_557,N_593);
xor U654 (N_654,N_565,N_568);
xnor U655 (N_655,N_543,N_554);
and U656 (N_656,N_594,N_595);
nand U657 (N_657,N_541,N_599);
and U658 (N_658,N_581,N_579);
nand U659 (N_659,N_552,N_587);
and U660 (N_660,N_569,N_528);
and U661 (N_661,N_581,N_591);
nor U662 (N_662,N_551,N_544);
and U663 (N_663,N_532,N_542);
or U664 (N_664,N_582,N_586);
or U665 (N_665,N_539,N_542);
xor U666 (N_666,N_568,N_591);
nand U667 (N_667,N_530,N_568);
and U668 (N_668,N_578,N_550);
or U669 (N_669,N_596,N_599);
and U670 (N_670,N_539,N_577);
or U671 (N_671,N_546,N_579);
or U672 (N_672,N_547,N_596);
nand U673 (N_673,N_543,N_599);
nor U674 (N_674,N_528,N_597);
nor U675 (N_675,N_673,N_620);
nor U676 (N_676,N_649,N_627);
xnor U677 (N_677,N_672,N_664);
xor U678 (N_678,N_657,N_624);
and U679 (N_679,N_658,N_643);
and U680 (N_680,N_631,N_670);
xnor U681 (N_681,N_663,N_648);
nand U682 (N_682,N_636,N_638);
or U683 (N_683,N_661,N_633);
nand U684 (N_684,N_611,N_634);
nor U685 (N_685,N_622,N_618);
nor U686 (N_686,N_612,N_667);
and U687 (N_687,N_652,N_603);
nor U688 (N_688,N_602,N_637);
or U689 (N_689,N_669,N_639);
nor U690 (N_690,N_647,N_646);
or U691 (N_691,N_644,N_665);
nor U692 (N_692,N_621,N_614);
and U693 (N_693,N_645,N_660);
and U694 (N_694,N_616,N_626);
and U695 (N_695,N_600,N_662);
xor U696 (N_696,N_608,N_651);
nand U697 (N_697,N_604,N_605);
and U698 (N_698,N_655,N_607);
nor U699 (N_699,N_628,N_668);
or U700 (N_700,N_601,N_617);
nor U701 (N_701,N_606,N_659);
and U702 (N_702,N_619,N_615);
nor U703 (N_703,N_623,N_630);
nand U704 (N_704,N_610,N_629);
nand U705 (N_705,N_656,N_635);
or U706 (N_706,N_613,N_671);
and U707 (N_707,N_653,N_650);
nand U708 (N_708,N_632,N_654);
xor U709 (N_709,N_640,N_666);
nor U710 (N_710,N_609,N_625);
nand U711 (N_711,N_642,N_674);
or U712 (N_712,N_641,N_646);
and U713 (N_713,N_656,N_643);
and U714 (N_714,N_652,N_642);
xor U715 (N_715,N_667,N_611);
xor U716 (N_716,N_620,N_621);
nor U717 (N_717,N_623,N_640);
and U718 (N_718,N_608,N_610);
and U719 (N_719,N_656,N_613);
and U720 (N_720,N_605,N_668);
or U721 (N_721,N_616,N_661);
or U722 (N_722,N_648,N_668);
nor U723 (N_723,N_609,N_624);
nor U724 (N_724,N_646,N_649);
nand U725 (N_725,N_637,N_611);
nor U726 (N_726,N_650,N_611);
nand U727 (N_727,N_625,N_635);
nand U728 (N_728,N_664,N_660);
nand U729 (N_729,N_640,N_647);
and U730 (N_730,N_622,N_674);
and U731 (N_731,N_646,N_644);
nor U732 (N_732,N_658,N_617);
xor U733 (N_733,N_653,N_662);
and U734 (N_734,N_627,N_624);
or U735 (N_735,N_624,N_632);
nor U736 (N_736,N_623,N_666);
xnor U737 (N_737,N_657,N_625);
nor U738 (N_738,N_619,N_647);
nand U739 (N_739,N_605,N_606);
nor U740 (N_740,N_617,N_608);
and U741 (N_741,N_601,N_644);
nand U742 (N_742,N_659,N_612);
nand U743 (N_743,N_625,N_634);
nor U744 (N_744,N_651,N_660);
nand U745 (N_745,N_629,N_631);
or U746 (N_746,N_617,N_624);
and U747 (N_747,N_654,N_650);
and U748 (N_748,N_600,N_648);
nand U749 (N_749,N_657,N_660);
xnor U750 (N_750,N_707,N_687);
or U751 (N_751,N_680,N_689);
nor U752 (N_752,N_745,N_729);
and U753 (N_753,N_688,N_739);
nand U754 (N_754,N_695,N_719);
nand U755 (N_755,N_749,N_701);
or U756 (N_756,N_735,N_691);
and U757 (N_757,N_681,N_734);
nor U758 (N_758,N_737,N_736);
nor U759 (N_759,N_704,N_682);
or U760 (N_760,N_706,N_710);
or U761 (N_761,N_692,N_693);
nor U762 (N_762,N_726,N_709);
and U763 (N_763,N_713,N_700);
nor U764 (N_764,N_702,N_724);
xor U765 (N_765,N_711,N_699);
and U766 (N_766,N_722,N_714);
nor U767 (N_767,N_712,N_723);
or U768 (N_768,N_677,N_697);
and U769 (N_769,N_747,N_679);
or U770 (N_770,N_738,N_744);
or U771 (N_771,N_740,N_733);
nand U772 (N_772,N_715,N_708);
nand U773 (N_773,N_731,N_684);
and U774 (N_774,N_720,N_732);
and U775 (N_775,N_685,N_675);
or U776 (N_776,N_746,N_718);
xor U777 (N_777,N_743,N_748);
and U778 (N_778,N_683,N_742);
nand U779 (N_779,N_727,N_690);
nor U780 (N_780,N_741,N_705);
or U781 (N_781,N_717,N_696);
nor U782 (N_782,N_716,N_728);
or U783 (N_783,N_678,N_698);
or U784 (N_784,N_703,N_725);
xor U785 (N_785,N_721,N_694);
nand U786 (N_786,N_730,N_676);
nor U787 (N_787,N_686,N_709);
nand U788 (N_788,N_704,N_715);
nand U789 (N_789,N_690,N_700);
and U790 (N_790,N_742,N_715);
and U791 (N_791,N_730,N_702);
nor U792 (N_792,N_748,N_691);
or U793 (N_793,N_740,N_718);
xnor U794 (N_794,N_718,N_703);
or U795 (N_795,N_747,N_697);
xnor U796 (N_796,N_729,N_736);
and U797 (N_797,N_728,N_711);
or U798 (N_798,N_726,N_696);
and U799 (N_799,N_745,N_721);
and U800 (N_800,N_727,N_716);
and U801 (N_801,N_695,N_694);
nor U802 (N_802,N_688,N_720);
nor U803 (N_803,N_705,N_745);
nor U804 (N_804,N_720,N_707);
nor U805 (N_805,N_692,N_724);
nor U806 (N_806,N_710,N_735);
nor U807 (N_807,N_677,N_736);
nand U808 (N_808,N_681,N_740);
and U809 (N_809,N_736,N_728);
xnor U810 (N_810,N_683,N_675);
and U811 (N_811,N_715,N_746);
or U812 (N_812,N_722,N_736);
nor U813 (N_813,N_705,N_687);
and U814 (N_814,N_743,N_732);
and U815 (N_815,N_739,N_705);
nand U816 (N_816,N_688,N_693);
nand U817 (N_817,N_735,N_717);
and U818 (N_818,N_677,N_711);
and U819 (N_819,N_689,N_687);
and U820 (N_820,N_707,N_739);
xnor U821 (N_821,N_694,N_696);
nand U822 (N_822,N_737,N_744);
and U823 (N_823,N_676,N_722);
xnor U824 (N_824,N_731,N_694);
nand U825 (N_825,N_763,N_783);
nor U826 (N_826,N_775,N_789);
nand U827 (N_827,N_768,N_757);
or U828 (N_828,N_762,N_777);
nand U829 (N_829,N_770,N_755);
and U830 (N_830,N_803,N_812);
nand U831 (N_831,N_815,N_772);
nand U832 (N_832,N_754,N_822);
nor U833 (N_833,N_778,N_794);
or U834 (N_834,N_819,N_786);
and U835 (N_835,N_771,N_751);
nor U836 (N_836,N_816,N_792);
nor U837 (N_837,N_773,N_799);
or U838 (N_838,N_769,N_824);
nand U839 (N_839,N_809,N_796);
and U840 (N_840,N_761,N_805);
or U841 (N_841,N_808,N_823);
and U842 (N_842,N_767,N_804);
or U843 (N_843,N_756,N_780);
nand U844 (N_844,N_797,N_793);
nand U845 (N_845,N_784,N_806);
and U846 (N_846,N_782,N_764);
or U847 (N_847,N_750,N_774);
and U848 (N_848,N_788,N_791);
xnor U849 (N_849,N_811,N_807);
or U850 (N_850,N_787,N_765);
nand U851 (N_851,N_802,N_821);
xor U852 (N_852,N_785,N_760);
and U853 (N_853,N_801,N_820);
nand U854 (N_854,N_766,N_752);
or U855 (N_855,N_818,N_753);
nor U856 (N_856,N_813,N_779);
or U857 (N_857,N_758,N_776);
or U858 (N_858,N_759,N_814);
xor U859 (N_859,N_810,N_817);
and U860 (N_860,N_781,N_800);
nor U861 (N_861,N_790,N_795);
nor U862 (N_862,N_798,N_757);
nand U863 (N_863,N_816,N_811);
nand U864 (N_864,N_777,N_792);
nor U865 (N_865,N_758,N_753);
and U866 (N_866,N_807,N_762);
nand U867 (N_867,N_766,N_807);
nand U868 (N_868,N_799,N_791);
or U869 (N_869,N_755,N_776);
and U870 (N_870,N_756,N_797);
nor U871 (N_871,N_787,N_774);
nand U872 (N_872,N_784,N_762);
nor U873 (N_873,N_777,N_795);
nand U874 (N_874,N_815,N_789);
xnor U875 (N_875,N_795,N_802);
nand U876 (N_876,N_798,N_820);
or U877 (N_877,N_823,N_758);
nand U878 (N_878,N_791,N_793);
nor U879 (N_879,N_785,N_755);
or U880 (N_880,N_807,N_754);
or U881 (N_881,N_780,N_817);
xnor U882 (N_882,N_786,N_794);
xnor U883 (N_883,N_764,N_790);
nand U884 (N_884,N_752,N_759);
or U885 (N_885,N_766,N_790);
and U886 (N_886,N_818,N_752);
nand U887 (N_887,N_777,N_816);
or U888 (N_888,N_773,N_775);
or U889 (N_889,N_796,N_752);
or U890 (N_890,N_762,N_817);
nand U891 (N_891,N_806,N_759);
xor U892 (N_892,N_770,N_809);
nand U893 (N_893,N_789,N_755);
and U894 (N_894,N_788,N_818);
or U895 (N_895,N_774,N_757);
nand U896 (N_896,N_810,N_796);
nand U897 (N_897,N_808,N_779);
xor U898 (N_898,N_764,N_820);
and U899 (N_899,N_786,N_752);
xor U900 (N_900,N_874,N_889);
or U901 (N_901,N_851,N_843);
and U902 (N_902,N_826,N_865);
nor U903 (N_903,N_844,N_846);
and U904 (N_904,N_892,N_880);
and U905 (N_905,N_841,N_842);
nand U906 (N_906,N_863,N_868);
nand U907 (N_907,N_876,N_878);
nand U908 (N_908,N_891,N_887);
nand U909 (N_909,N_879,N_831);
nor U910 (N_910,N_828,N_838);
nor U911 (N_911,N_853,N_836);
nor U912 (N_912,N_855,N_886);
nor U913 (N_913,N_896,N_833);
or U914 (N_914,N_840,N_864);
or U915 (N_915,N_884,N_872);
and U916 (N_916,N_885,N_895);
nor U917 (N_917,N_845,N_849);
or U918 (N_918,N_860,N_852);
nand U919 (N_919,N_847,N_862);
nand U920 (N_920,N_888,N_870);
or U921 (N_921,N_899,N_827);
xor U922 (N_922,N_873,N_871);
nand U923 (N_923,N_839,N_848);
or U924 (N_924,N_825,N_875);
and U925 (N_925,N_856,N_854);
nor U926 (N_926,N_894,N_861);
nand U927 (N_927,N_832,N_893);
xor U928 (N_928,N_897,N_837);
or U929 (N_929,N_857,N_834);
or U930 (N_930,N_858,N_829);
nor U931 (N_931,N_859,N_850);
or U932 (N_932,N_883,N_877);
or U933 (N_933,N_882,N_830);
xor U934 (N_934,N_898,N_869);
nor U935 (N_935,N_867,N_881);
nor U936 (N_936,N_866,N_835);
and U937 (N_937,N_890,N_855);
nand U938 (N_938,N_880,N_889);
or U939 (N_939,N_874,N_846);
nor U940 (N_940,N_850,N_828);
or U941 (N_941,N_845,N_825);
or U942 (N_942,N_839,N_876);
nor U943 (N_943,N_874,N_895);
nand U944 (N_944,N_826,N_837);
or U945 (N_945,N_849,N_882);
or U946 (N_946,N_878,N_880);
nand U947 (N_947,N_888,N_898);
nand U948 (N_948,N_850,N_865);
or U949 (N_949,N_862,N_829);
or U950 (N_950,N_832,N_829);
nand U951 (N_951,N_898,N_830);
nand U952 (N_952,N_869,N_884);
and U953 (N_953,N_826,N_860);
and U954 (N_954,N_860,N_830);
and U955 (N_955,N_849,N_874);
nor U956 (N_956,N_852,N_858);
and U957 (N_957,N_898,N_838);
and U958 (N_958,N_847,N_891);
nor U959 (N_959,N_887,N_894);
or U960 (N_960,N_860,N_867);
and U961 (N_961,N_828,N_856);
or U962 (N_962,N_863,N_859);
or U963 (N_963,N_847,N_845);
and U964 (N_964,N_826,N_845);
or U965 (N_965,N_887,N_836);
nand U966 (N_966,N_843,N_869);
nor U967 (N_967,N_865,N_868);
and U968 (N_968,N_853,N_892);
and U969 (N_969,N_857,N_878);
nand U970 (N_970,N_840,N_888);
or U971 (N_971,N_843,N_889);
nand U972 (N_972,N_877,N_851);
and U973 (N_973,N_897,N_827);
nor U974 (N_974,N_857,N_866);
nand U975 (N_975,N_947,N_941);
and U976 (N_976,N_902,N_956);
and U977 (N_977,N_948,N_952);
xor U978 (N_978,N_970,N_960);
nor U979 (N_979,N_910,N_922);
nor U980 (N_980,N_958,N_973);
xnor U981 (N_981,N_927,N_966);
nand U982 (N_982,N_968,N_946);
nor U983 (N_983,N_919,N_962);
nor U984 (N_984,N_943,N_934);
and U985 (N_985,N_906,N_912);
and U986 (N_986,N_913,N_911);
xor U987 (N_987,N_901,N_971);
nor U988 (N_988,N_949,N_917);
and U989 (N_989,N_925,N_903);
and U990 (N_990,N_939,N_933);
or U991 (N_991,N_929,N_921);
or U992 (N_992,N_918,N_936);
and U993 (N_993,N_967,N_950);
nand U994 (N_994,N_905,N_965);
nand U995 (N_995,N_969,N_961);
nor U996 (N_996,N_932,N_915);
xor U997 (N_997,N_937,N_924);
or U998 (N_998,N_951,N_909);
nand U999 (N_999,N_955,N_974);
nand U1000 (N_1000,N_963,N_908);
or U1001 (N_1001,N_928,N_935);
or U1002 (N_1002,N_940,N_953);
nor U1003 (N_1003,N_938,N_900);
nor U1004 (N_1004,N_904,N_923);
nand U1005 (N_1005,N_944,N_945);
or U1006 (N_1006,N_926,N_942);
xor U1007 (N_1007,N_931,N_920);
or U1008 (N_1008,N_914,N_916);
xnor U1009 (N_1009,N_954,N_957);
or U1010 (N_1010,N_972,N_907);
or U1011 (N_1011,N_959,N_930);
and U1012 (N_1012,N_964,N_905);
nor U1013 (N_1013,N_907,N_927);
nor U1014 (N_1014,N_940,N_968);
xnor U1015 (N_1015,N_928,N_952);
nor U1016 (N_1016,N_946,N_922);
and U1017 (N_1017,N_918,N_965);
and U1018 (N_1018,N_917,N_936);
and U1019 (N_1019,N_911,N_948);
and U1020 (N_1020,N_913,N_953);
nand U1021 (N_1021,N_970,N_941);
nand U1022 (N_1022,N_940,N_957);
and U1023 (N_1023,N_920,N_941);
nand U1024 (N_1024,N_930,N_974);
nand U1025 (N_1025,N_954,N_935);
and U1026 (N_1026,N_919,N_963);
nand U1027 (N_1027,N_904,N_903);
nand U1028 (N_1028,N_923,N_959);
and U1029 (N_1029,N_902,N_921);
and U1030 (N_1030,N_947,N_902);
and U1031 (N_1031,N_962,N_906);
and U1032 (N_1032,N_970,N_910);
and U1033 (N_1033,N_961,N_941);
nand U1034 (N_1034,N_953,N_973);
nand U1035 (N_1035,N_913,N_964);
xor U1036 (N_1036,N_964,N_925);
nand U1037 (N_1037,N_965,N_945);
nor U1038 (N_1038,N_957,N_921);
and U1039 (N_1039,N_905,N_974);
nand U1040 (N_1040,N_928,N_917);
or U1041 (N_1041,N_974,N_932);
or U1042 (N_1042,N_957,N_958);
nand U1043 (N_1043,N_955,N_967);
xnor U1044 (N_1044,N_966,N_914);
nor U1045 (N_1045,N_907,N_963);
nand U1046 (N_1046,N_917,N_966);
nand U1047 (N_1047,N_937,N_960);
or U1048 (N_1048,N_905,N_931);
nand U1049 (N_1049,N_900,N_936);
or U1050 (N_1050,N_1031,N_989);
xnor U1051 (N_1051,N_1047,N_991);
and U1052 (N_1052,N_1000,N_1011);
or U1053 (N_1053,N_995,N_977);
nand U1054 (N_1054,N_1032,N_1009);
and U1055 (N_1055,N_1008,N_987);
and U1056 (N_1056,N_1029,N_1001);
and U1057 (N_1057,N_1045,N_1004);
and U1058 (N_1058,N_979,N_1048);
or U1059 (N_1059,N_988,N_993);
nand U1060 (N_1060,N_1043,N_1013);
nand U1061 (N_1061,N_990,N_997);
xor U1062 (N_1062,N_1046,N_1010);
nor U1063 (N_1063,N_1018,N_1002);
nand U1064 (N_1064,N_1007,N_1020);
or U1065 (N_1065,N_1019,N_1014);
nand U1066 (N_1066,N_1036,N_1025);
xor U1067 (N_1067,N_1016,N_1049);
or U1068 (N_1068,N_980,N_1037);
nor U1069 (N_1069,N_1023,N_975);
and U1070 (N_1070,N_978,N_1006);
xor U1071 (N_1071,N_1035,N_982);
or U1072 (N_1072,N_981,N_1039);
nor U1073 (N_1073,N_976,N_1003);
and U1074 (N_1074,N_1028,N_1044);
and U1075 (N_1075,N_1026,N_999);
nor U1076 (N_1076,N_1017,N_986);
and U1077 (N_1077,N_1021,N_1015);
and U1078 (N_1078,N_1042,N_1022);
nand U1079 (N_1079,N_1041,N_1005);
and U1080 (N_1080,N_992,N_985);
xor U1081 (N_1081,N_1030,N_983);
and U1082 (N_1082,N_984,N_1012);
nand U1083 (N_1083,N_996,N_994);
nand U1084 (N_1084,N_1027,N_998);
or U1085 (N_1085,N_1040,N_1024);
nor U1086 (N_1086,N_1034,N_1033);
xor U1087 (N_1087,N_1038,N_981);
and U1088 (N_1088,N_985,N_997);
nand U1089 (N_1089,N_1027,N_987);
nor U1090 (N_1090,N_983,N_1003);
and U1091 (N_1091,N_1023,N_1014);
nor U1092 (N_1092,N_976,N_1010);
and U1093 (N_1093,N_1014,N_1028);
and U1094 (N_1094,N_999,N_1038);
or U1095 (N_1095,N_999,N_976);
nand U1096 (N_1096,N_994,N_998);
or U1097 (N_1097,N_1005,N_996);
nor U1098 (N_1098,N_979,N_1046);
nand U1099 (N_1099,N_1013,N_987);
and U1100 (N_1100,N_1002,N_987);
and U1101 (N_1101,N_989,N_981);
or U1102 (N_1102,N_997,N_1043);
and U1103 (N_1103,N_1028,N_1023);
nor U1104 (N_1104,N_1014,N_1041);
nand U1105 (N_1105,N_1027,N_1030);
or U1106 (N_1106,N_1020,N_1048);
or U1107 (N_1107,N_989,N_1005);
or U1108 (N_1108,N_1043,N_985);
and U1109 (N_1109,N_1007,N_995);
nor U1110 (N_1110,N_977,N_1009);
nand U1111 (N_1111,N_1048,N_1028);
nand U1112 (N_1112,N_1022,N_977);
or U1113 (N_1113,N_1021,N_989);
or U1114 (N_1114,N_975,N_1043);
or U1115 (N_1115,N_999,N_1042);
or U1116 (N_1116,N_987,N_1023);
or U1117 (N_1117,N_1017,N_1015);
and U1118 (N_1118,N_991,N_997);
or U1119 (N_1119,N_978,N_1011);
and U1120 (N_1120,N_993,N_1034);
and U1121 (N_1121,N_1015,N_1006);
or U1122 (N_1122,N_1033,N_1036);
nor U1123 (N_1123,N_998,N_984);
nand U1124 (N_1124,N_1014,N_1022);
xor U1125 (N_1125,N_1110,N_1084);
nand U1126 (N_1126,N_1093,N_1087);
and U1127 (N_1127,N_1109,N_1073);
or U1128 (N_1128,N_1060,N_1094);
nand U1129 (N_1129,N_1052,N_1072);
or U1130 (N_1130,N_1064,N_1116);
nand U1131 (N_1131,N_1117,N_1054);
or U1132 (N_1132,N_1097,N_1083);
nor U1133 (N_1133,N_1112,N_1068);
or U1134 (N_1134,N_1067,N_1078);
or U1135 (N_1135,N_1124,N_1086);
or U1136 (N_1136,N_1096,N_1113);
nand U1137 (N_1137,N_1085,N_1115);
nor U1138 (N_1138,N_1062,N_1051);
xnor U1139 (N_1139,N_1061,N_1100);
nand U1140 (N_1140,N_1079,N_1099);
and U1141 (N_1141,N_1050,N_1111);
and U1142 (N_1142,N_1059,N_1122);
and U1143 (N_1143,N_1121,N_1082);
nand U1144 (N_1144,N_1095,N_1090);
nor U1145 (N_1145,N_1066,N_1055);
or U1146 (N_1146,N_1091,N_1070);
nor U1147 (N_1147,N_1089,N_1080);
nor U1148 (N_1148,N_1071,N_1119);
and U1149 (N_1149,N_1105,N_1120);
nand U1150 (N_1150,N_1081,N_1053);
nand U1151 (N_1151,N_1074,N_1114);
or U1152 (N_1152,N_1107,N_1103);
xor U1153 (N_1153,N_1063,N_1088);
nor U1154 (N_1154,N_1108,N_1058);
or U1155 (N_1155,N_1077,N_1104);
or U1156 (N_1156,N_1123,N_1056);
nor U1157 (N_1157,N_1069,N_1092);
nand U1158 (N_1158,N_1098,N_1075);
or U1159 (N_1159,N_1101,N_1065);
nor U1160 (N_1160,N_1106,N_1076);
nor U1161 (N_1161,N_1057,N_1118);
or U1162 (N_1162,N_1102,N_1119);
nand U1163 (N_1163,N_1103,N_1100);
and U1164 (N_1164,N_1091,N_1123);
or U1165 (N_1165,N_1122,N_1112);
or U1166 (N_1166,N_1060,N_1091);
or U1167 (N_1167,N_1060,N_1120);
and U1168 (N_1168,N_1096,N_1097);
nand U1169 (N_1169,N_1051,N_1093);
or U1170 (N_1170,N_1122,N_1053);
nor U1171 (N_1171,N_1097,N_1092);
and U1172 (N_1172,N_1110,N_1114);
and U1173 (N_1173,N_1082,N_1061);
and U1174 (N_1174,N_1096,N_1120);
nand U1175 (N_1175,N_1058,N_1083);
and U1176 (N_1176,N_1097,N_1098);
nand U1177 (N_1177,N_1122,N_1096);
nand U1178 (N_1178,N_1094,N_1077);
or U1179 (N_1179,N_1115,N_1100);
or U1180 (N_1180,N_1110,N_1088);
nand U1181 (N_1181,N_1069,N_1054);
nand U1182 (N_1182,N_1083,N_1109);
nor U1183 (N_1183,N_1087,N_1071);
nor U1184 (N_1184,N_1094,N_1116);
xnor U1185 (N_1185,N_1068,N_1065);
xor U1186 (N_1186,N_1119,N_1090);
nor U1187 (N_1187,N_1078,N_1108);
nor U1188 (N_1188,N_1087,N_1073);
nor U1189 (N_1189,N_1067,N_1094);
or U1190 (N_1190,N_1050,N_1085);
or U1191 (N_1191,N_1095,N_1052);
xor U1192 (N_1192,N_1099,N_1052);
or U1193 (N_1193,N_1106,N_1101);
nor U1194 (N_1194,N_1110,N_1082);
or U1195 (N_1195,N_1102,N_1053);
nand U1196 (N_1196,N_1071,N_1124);
and U1197 (N_1197,N_1108,N_1116);
xnor U1198 (N_1198,N_1053,N_1096);
and U1199 (N_1199,N_1097,N_1072);
xor U1200 (N_1200,N_1142,N_1166);
nand U1201 (N_1201,N_1181,N_1196);
or U1202 (N_1202,N_1186,N_1163);
and U1203 (N_1203,N_1136,N_1133);
or U1204 (N_1204,N_1141,N_1169);
nor U1205 (N_1205,N_1183,N_1127);
xor U1206 (N_1206,N_1187,N_1158);
nand U1207 (N_1207,N_1179,N_1138);
xor U1208 (N_1208,N_1125,N_1156);
nand U1209 (N_1209,N_1168,N_1197);
nor U1210 (N_1210,N_1162,N_1155);
and U1211 (N_1211,N_1149,N_1152);
and U1212 (N_1212,N_1148,N_1131);
and U1213 (N_1213,N_1170,N_1199);
nor U1214 (N_1214,N_1134,N_1180);
nor U1215 (N_1215,N_1151,N_1190);
nor U1216 (N_1216,N_1154,N_1178);
nor U1217 (N_1217,N_1137,N_1126);
nor U1218 (N_1218,N_1146,N_1157);
or U1219 (N_1219,N_1159,N_1174);
nand U1220 (N_1220,N_1182,N_1191);
and U1221 (N_1221,N_1195,N_1192);
or U1222 (N_1222,N_1171,N_1164);
and U1223 (N_1223,N_1167,N_1130);
nand U1224 (N_1224,N_1143,N_1176);
nand U1225 (N_1225,N_1194,N_1135);
or U1226 (N_1226,N_1175,N_1153);
and U1227 (N_1227,N_1189,N_1188);
and U1228 (N_1228,N_1139,N_1165);
or U1229 (N_1229,N_1129,N_1144);
and U1230 (N_1230,N_1184,N_1128);
nor U1231 (N_1231,N_1160,N_1172);
and U1232 (N_1232,N_1185,N_1198);
nand U1233 (N_1233,N_1193,N_1173);
and U1234 (N_1234,N_1177,N_1145);
nand U1235 (N_1235,N_1140,N_1132);
nand U1236 (N_1236,N_1150,N_1147);
xnor U1237 (N_1237,N_1161,N_1135);
nand U1238 (N_1238,N_1177,N_1182);
nand U1239 (N_1239,N_1133,N_1150);
nor U1240 (N_1240,N_1125,N_1151);
nand U1241 (N_1241,N_1148,N_1132);
and U1242 (N_1242,N_1156,N_1134);
nand U1243 (N_1243,N_1191,N_1174);
or U1244 (N_1244,N_1170,N_1180);
and U1245 (N_1245,N_1133,N_1197);
or U1246 (N_1246,N_1180,N_1126);
and U1247 (N_1247,N_1192,N_1168);
or U1248 (N_1248,N_1150,N_1125);
xnor U1249 (N_1249,N_1131,N_1184);
nor U1250 (N_1250,N_1143,N_1151);
nor U1251 (N_1251,N_1137,N_1125);
xor U1252 (N_1252,N_1169,N_1162);
nand U1253 (N_1253,N_1149,N_1143);
nor U1254 (N_1254,N_1165,N_1194);
nor U1255 (N_1255,N_1155,N_1125);
xnor U1256 (N_1256,N_1135,N_1158);
or U1257 (N_1257,N_1189,N_1178);
nand U1258 (N_1258,N_1175,N_1143);
or U1259 (N_1259,N_1166,N_1189);
nand U1260 (N_1260,N_1189,N_1195);
nand U1261 (N_1261,N_1146,N_1148);
nand U1262 (N_1262,N_1171,N_1132);
or U1263 (N_1263,N_1157,N_1162);
nor U1264 (N_1264,N_1186,N_1191);
nand U1265 (N_1265,N_1191,N_1189);
nand U1266 (N_1266,N_1195,N_1188);
and U1267 (N_1267,N_1156,N_1159);
nor U1268 (N_1268,N_1182,N_1173);
nand U1269 (N_1269,N_1132,N_1150);
or U1270 (N_1270,N_1159,N_1135);
nor U1271 (N_1271,N_1142,N_1198);
or U1272 (N_1272,N_1194,N_1158);
nor U1273 (N_1273,N_1196,N_1171);
nor U1274 (N_1274,N_1143,N_1147);
xnor U1275 (N_1275,N_1262,N_1215);
nor U1276 (N_1276,N_1230,N_1201);
nand U1277 (N_1277,N_1257,N_1225);
or U1278 (N_1278,N_1213,N_1269);
and U1279 (N_1279,N_1202,N_1273);
nor U1280 (N_1280,N_1245,N_1204);
and U1281 (N_1281,N_1247,N_1263);
and U1282 (N_1282,N_1268,N_1242);
and U1283 (N_1283,N_1233,N_1224);
nor U1284 (N_1284,N_1229,N_1218);
and U1285 (N_1285,N_1255,N_1252);
xor U1286 (N_1286,N_1207,N_1236);
and U1287 (N_1287,N_1265,N_1241);
and U1288 (N_1288,N_1240,N_1228);
and U1289 (N_1289,N_1217,N_1259);
nor U1290 (N_1290,N_1272,N_1219);
nand U1291 (N_1291,N_1254,N_1231);
or U1292 (N_1292,N_1211,N_1221);
nor U1293 (N_1293,N_1212,N_1237);
or U1294 (N_1294,N_1239,N_1235);
nand U1295 (N_1295,N_1206,N_1249);
nand U1296 (N_1296,N_1210,N_1208);
nand U1297 (N_1297,N_1243,N_1261);
or U1298 (N_1298,N_1227,N_1223);
and U1299 (N_1299,N_1222,N_1220);
nand U1300 (N_1300,N_1209,N_1246);
or U1301 (N_1301,N_1232,N_1214);
and U1302 (N_1302,N_1258,N_1226);
nor U1303 (N_1303,N_1200,N_1248);
or U1304 (N_1304,N_1264,N_1251);
nand U1305 (N_1305,N_1203,N_1274);
nor U1306 (N_1306,N_1234,N_1266);
and U1307 (N_1307,N_1256,N_1253);
nand U1308 (N_1308,N_1250,N_1271);
nand U1309 (N_1309,N_1260,N_1238);
nor U1310 (N_1310,N_1267,N_1205);
or U1311 (N_1311,N_1244,N_1216);
and U1312 (N_1312,N_1270,N_1228);
nand U1313 (N_1313,N_1220,N_1273);
nand U1314 (N_1314,N_1238,N_1237);
nand U1315 (N_1315,N_1243,N_1217);
or U1316 (N_1316,N_1241,N_1217);
nand U1317 (N_1317,N_1265,N_1217);
nand U1318 (N_1318,N_1249,N_1251);
nor U1319 (N_1319,N_1220,N_1200);
or U1320 (N_1320,N_1233,N_1207);
xnor U1321 (N_1321,N_1243,N_1254);
and U1322 (N_1322,N_1201,N_1271);
nand U1323 (N_1323,N_1210,N_1204);
and U1324 (N_1324,N_1212,N_1244);
nor U1325 (N_1325,N_1221,N_1267);
and U1326 (N_1326,N_1255,N_1262);
and U1327 (N_1327,N_1204,N_1235);
and U1328 (N_1328,N_1222,N_1208);
or U1329 (N_1329,N_1240,N_1265);
nand U1330 (N_1330,N_1207,N_1214);
and U1331 (N_1331,N_1228,N_1216);
and U1332 (N_1332,N_1271,N_1219);
or U1333 (N_1333,N_1208,N_1229);
nand U1334 (N_1334,N_1249,N_1272);
nor U1335 (N_1335,N_1249,N_1264);
nand U1336 (N_1336,N_1274,N_1214);
xnor U1337 (N_1337,N_1234,N_1219);
or U1338 (N_1338,N_1267,N_1273);
and U1339 (N_1339,N_1208,N_1214);
nand U1340 (N_1340,N_1201,N_1251);
nor U1341 (N_1341,N_1213,N_1246);
xor U1342 (N_1342,N_1252,N_1218);
xnor U1343 (N_1343,N_1207,N_1218);
or U1344 (N_1344,N_1216,N_1267);
or U1345 (N_1345,N_1265,N_1272);
nor U1346 (N_1346,N_1219,N_1257);
and U1347 (N_1347,N_1244,N_1271);
or U1348 (N_1348,N_1235,N_1268);
or U1349 (N_1349,N_1233,N_1205);
or U1350 (N_1350,N_1298,N_1277);
xor U1351 (N_1351,N_1322,N_1307);
or U1352 (N_1352,N_1343,N_1332);
or U1353 (N_1353,N_1313,N_1284);
and U1354 (N_1354,N_1331,N_1334);
xor U1355 (N_1355,N_1301,N_1296);
nor U1356 (N_1356,N_1336,N_1325);
nor U1357 (N_1357,N_1326,N_1339);
and U1358 (N_1358,N_1308,N_1299);
or U1359 (N_1359,N_1291,N_1303);
and U1360 (N_1360,N_1321,N_1323);
or U1361 (N_1361,N_1305,N_1278);
nor U1362 (N_1362,N_1285,N_1335);
nor U1363 (N_1363,N_1314,N_1318);
or U1364 (N_1364,N_1311,N_1283);
nand U1365 (N_1365,N_1310,N_1287);
nand U1366 (N_1366,N_1293,N_1337);
or U1367 (N_1367,N_1348,N_1294);
nor U1368 (N_1368,N_1304,N_1324);
or U1369 (N_1369,N_1279,N_1342);
nand U1370 (N_1370,N_1317,N_1276);
and U1371 (N_1371,N_1281,N_1290);
nor U1372 (N_1372,N_1292,N_1297);
nand U1373 (N_1373,N_1328,N_1302);
nor U1374 (N_1374,N_1333,N_1347);
nor U1375 (N_1375,N_1275,N_1288);
nor U1376 (N_1376,N_1286,N_1320);
or U1377 (N_1377,N_1300,N_1341);
or U1378 (N_1378,N_1346,N_1344);
xor U1379 (N_1379,N_1349,N_1295);
nand U1380 (N_1380,N_1282,N_1309);
or U1381 (N_1381,N_1306,N_1312);
nand U1382 (N_1382,N_1315,N_1316);
or U1383 (N_1383,N_1330,N_1338);
xnor U1384 (N_1384,N_1327,N_1340);
nor U1385 (N_1385,N_1345,N_1280);
nor U1386 (N_1386,N_1289,N_1319);
nand U1387 (N_1387,N_1329,N_1315);
nor U1388 (N_1388,N_1322,N_1319);
nor U1389 (N_1389,N_1321,N_1290);
nand U1390 (N_1390,N_1303,N_1346);
nand U1391 (N_1391,N_1325,N_1321);
and U1392 (N_1392,N_1305,N_1308);
and U1393 (N_1393,N_1289,N_1301);
or U1394 (N_1394,N_1332,N_1276);
xnor U1395 (N_1395,N_1316,N_1275);
xor U1396 (N_1396,N_1321,N_1281);
nand U1397 (N_1397,N_1299,N_1340);
xor U1398 (N_1398,N_1330,N_1346);
and U1399 (N_1399,N_1333,N_1313);
nand U1400 (N_1400,N_1280,N_1278);
nand U1401 (N_1401,N_1329,N_1299);
or U1402 (N_1402,N_1321,N_1329);
and U1403 (N_1403,N_1293,N_1347);
xor U1404 (N_1404,N_1301,N_1308);
nand U1405 (N_1405,N_1322,N_1345);
nor U1406 (N_1406,N_1335,N_1300);
and U1407 (N_1407,N_1340,N_1308);
nor U1408 (N_1408,N_1275,N_1304);
nor U1409 (N_1409,N_1325,N_1280);
and U1410 (N_1410,N_1336,N_1323);
xor U1411 (N_1411,N_1287,N_1328);
and U1412 (N_1412,N_1277,N_1279);
and U1413 (N_1413,N_1347,N_1341);
or U1414 (N_1414,N_1322,N_1320);
and U1415 (N_1415,N_1287,N_1321);
or U1416 (N_1416,N_1304,N_1279);
and U1417 (N_1417,N_1283,N_1333);
nor U1418 (N_1418,N_1293,N_1285);
nor U1419 (N_1419,N_1276,N_1343);
or U1420 (N_1420,N_1316,N_1319);
nand U1421 (N_1421,N_1303,N_1304);
nand U1422 (N_1422,N_1287,N_1312);
nor U1423 (N_1423,N_1303,N_1281);
nand U1424 (N_1424,N_1320,N_1278);
nor U1425 (N_1425,N_1415,N_1379);
or U1426 (N_1426,N_1371,N_1413);
nand U1427 (N_1427,N_1376,N_1384);
nor U1428 (N_1428,N_1419,N_1357);
and U1429 (N_1429,N_1402,N_1411);
nor U1430 (N_1430,N_1410,N_1351);
nand U1431 (N_1431,N_1404,N_1380);
xor U1432 (N_1432,N_1355,N_1403);
nor U1433 (N_1433,N_1414,N_1409);
and U1434 (N_1434,N_1375,N_1383);
and U1435 (N_1435,N_1396,N_1363);
or U1436 (N_1436,N_1420,N_1372);
or U1437 (N_1437,N_1378,N_1377);
and U1438 (N_1438,N_1386,N_1400);
nor U1439 (N_1439,N_1350,N_1417);
and U1440 (N_1440,N_1381,N_1401);
nor U1441 (N_1441,N_1398,N_1391);
xnor U1442 (N_1442,N_1359,N_1389);
or U1443 (N_1443,N_1397,N_1388);
nand U1444 (N_1444,N_1390,N_1360);
nand U1445 (N_1445,N_1422,N_1385);
nor U1446 (N_1446,N_1423,N_1424);
or U1447 (N_1447,N_1356,N_1364);
or U1448 (N_1448,N_1374,N_1366);
and U1449 (N_1449,N_1392,N_1408);
xnor U1450 (N_1450,N_1393,N_1368);
nand U1451 (N_1451,N_1405,N_1387);
or U1452 (N_1452,N_1367,N_1362);
nor U1453 (N_1453,N_1358,N_1370);
nor U1454 (N_1454,N_1418,N_1399);
xor U1455 (N_1455,N_1395,N_1394);
and U1456 (N_1456,N_1416,N_1353);
or U1457 (N_1457,N_1412,N_1354);
nor U1458 (N_1458,N_1407,N_1365);
nor U1459 (N_1459,N_1352,N_1421);
and U1460 (N_1460,N_1369,N_1382);
xnor U1461 (N_1461,N_1406,N_1373);
nand U1462 (N_1462,N_1361,N_1357);
nand U1463 (N_1463,N_1389,N_1410);
nor U1464 (N_1464,N_1373,N_1381);
and U1465 (N_1465,N_1411,N_1364);
nand U1466 (N_1466,N_1421,N_1355);
nand U1467 (N_1467,N_1363,N_1397);
nand U1468 (N_1468,N_1390,N_1380);
or U1469 (N_1469,N_1369,N_1410);
and U1470 (N_1470,N_1356,N_1415);
or U1471 (N_1471,N_1401,N_1359);
nor U1472 (N_1472,N_1406,N_1401);
nand U1473 (N_1473,N_1422,N_1374);
nor U1474 (N_1474,N_1410,N_1352);
and U1475 (N_1475,N_1389,N_1356);
or U1476 (N_1476,N_1359,N_1417);
xnor U1477 (N_1477,N_1417,N_1377);
xnor U1478 (N_1478,N_1422,N_1421);
or U1479 (N_1479,N_1356,N_1369);
or U1480 (N_1480,N_1392,N_1394);
or U1481 (N_1481,N_1384,N_1367);
nor U1482 (N_1482,N_1403,N_1406);
and U1483 (N_1483,N_1357,N_1402);
or U1484 (N_1484,N_1409,N_1379);
nor U1485 (N_1485,N_1366,N_1361);
nor U1486 (N_1486,N_1406,N_1355);
nand U1487 (N_1487,N_1371,N_1388);
or U1488 (N_1488,N_1396,N_1368);
xnor U1489 (N_1489,N_1379,N_1414);
nor U1490 (N_1490,N_1359,N_1352);
nand U1491 (N_1491,N_1367,N_1403);
and U1492 (N_1492,N_1396,N_1392);
and U1493 (N_1493,N_1397,N_1414);
xnor U1494 (N_1494,N_1398,N_1418);
nor U1495 (N_1495,N_1410,N_1395);
nor U1496 (N_1496,N_1357,N_1371);
and U1497 (N_1497,N_1422,N_1412);
nor U1498 (N_1498,N_1397,N_1382);
or U1499 (N_1499,N_1404,N_1372);
nand U1500 (N_1500,N_1435,N_1459);
xnor U1501 (N_1501,N_1464,N_1476);
nor U1502 (N_1502,N_1499,N_1439);
xnor U1503 (N_1503,N_1460,N_1454);
nor U1504 (N_1504,N_1457,N_1442);
and U1505 (N_1505,N_1462,N_1467);
nand U1506 (N_1506,N_1471,N_1481);
or U1507 (N_1507,N_1474,N_1492);
xor U1508 (N_1508,N_1430,N_1445);
and U1509 (N_1509,N_1441,N_1437);
or U1510 (N_1510,N_1478,N_1427);
or U1511 (N_1511,N_1485,N_1472);
nor U1512 (N_1512,N_1477,N_1479);
nand U1513 (N_1513,N_1487,N_1433);
nor U1514 (N_1514,N_1444,N_1469);
or U1515 (N_1515,N_1465,N_1451);
nor U1516 (N_1516,N_1496,N_1486);
or U1517 (N_1517,N_1426,N_1483);
nand U1518 (N_1518,N_1428,N_1431);
or U1519 (N_1519,N_1473,N_1468);
and U1520 (N_1520,N_1434,N_1443);
and U1521 (N_1521,N_1440,N_1489);
nor U1522 (N_1522,N_1497,N_1436);
nor U1523 (N_1523,N_1455,N_1466);
nor U1524 (N_1524,N_1495,N_1425);
xnor U1525 (N_1525,N_1447,N_1463);
and U1526 (N_1526,N_1498,N_1452);
nand U1527 (N_1527,N_1429,N_1484);
or U1528 (N_1528,N_1458,N_1491);
nor U1529 (N_1529,N_1448,N_1482);
and U1530 (N_1530,N_1480,N_1453);
nand U1531 (N_1531,N_1432,N_1449);
and U1532 (N_1532,N_1450,N_1475);
nor U1533 (N_1533,N_1456,N_1461);
or U1534 (N_1534,N_1490,N_1493);
xor U1535 (N_1535,N_1470,N_1494);
nor U1536 (N_1536,N_1446,N_1438);
xor U1537 (N_1537,N_1488,N_1444);
nor U1538 (N_1538,N_1467,N_1450);
xor U1539 (N_1539,N_1428,N_1467);
and U1540 (N_1540,N_1488,N_1451);
nand U1541 (N_1541,N_1487,N_1441);
nand U1542 (N_1542,N_1446,N_1437);
or U1543 (N_1543,N_1465,N_1471);
or U1544 (N_1544,N_1463,N_1494);
nand U1545 (N_1545,N_1466,N_1476);
and U1546 (N_1546,N_1492,N_1445);
nor U1547 (N_1547,N_1442,N_1447);
nor U1548 (N_1548,N_1494,N_1428);
nor U1549 (N_1549,N_1442,N_1453);
or U1550 (N_1550,N_1469,N_1459);
nand U1551 (N_1551,N_1425,N_1463);
nor U1552 (N_1552,N_1459,N_1489);
nor U1553 (N_1553,N_1451,N_1493);
nand U1554 (N_1554,N_1499,N_1431);
nor U1555 (N_1555,N_1498,N_1493);
nor U1556 (N_1556,N_1473,N_1427);
xnor U1557 (N_1557,N_1433,N_1438);
nand U1558 (N_1558,N_1442,N_1434);
nor U1559 (N_1559,N_1494,N_1480);
or U1560 (N_1560,N_1497,N_1442);
or U1561 (N_1561,N_1460,N_1455);
or U1562 (N_1562,N_1461,N_1442);
nand U1563 (N_1563,N_1447,N_1426);
nor U1564 (N_1564,N_1450,N_1485);
or U1565 (N_1565,N_1440,N_1453);
nand U1566 (N_1566,N_1454,N_1496);
nand U1567 (N_1567,N_1433,N_1472);
nor U1568 (N_1568,N_1438,N_1462);
and U1569 (N_1569,N_1430,N_1467);
nor U1570 (N_1570,N_1432,N_1435);
nor U1571 (N_1571,N_1458,N_1478);
or U1572 (N_1572,N_1433,N_1460);
xnor U1573 (N_1573,N_1469,N_1489);
or U1574 (N_1574,N_1483,N_1467);
nand U1575 (N_1575,N_1570,N_1558);
nor U1576 (N_1576,N_1537,N_1524);
nor U1577 (N_1577,N_1518,N_1571);
or U1578 (N_1578,N_1526,N_1555);
xnor U1579 (N_1579,N_1511,N_1540);
or U1580 (N_1580,N_1547,N_1504);
nand U1581 (N_1581,N_1501,N_1534);
nor U1582 (N_1582,N_1564,N_1567);
xor U1583 (N_1583,N_1559,N_1573);
xnor U1584 (N_1584,N_1549,N_1538);
or U1585 (N_1585,N_1508,N_1502);
nand U1586 (N_1586,N_1568,N_1513);
and U1587 (N_1587,N_1531,N_1550);
and U1588 (N_1588,N_1546,N_1522);
nand U1589 (N_1589,N_1542,N_1553);
nor U1590 (N_1590,N_1565,N_1519);
nor U1591 (N_1591,N_1528,N_1532);
nor U1592 (N_1592,N_1566,N_1520);
nor U1593 (N_1593,N_1512,N_1561);
or U1594 (N_1594,N_1507,N_1505);
nand U1595 (N_1595,N_1574,N_1517);
and U1596 (N_1596,N_1544,N_1533);
nor U1597 (N_1597,N_1509,N_1530);
nor U1598 (N_1598,N_1521,N_1557);
xnor U1599 (N_1599,N_1503,N_1523);
and U1600 (N_1600,N_1539,N_1548);
and U1601 (N_1601,N_1536,N_1551);
nand U1602 (N_1602,N_1525,N_1560);
nor U1603 (N_1603,N_1500,N_1563);
and U1604 (N_1604,N_1527,N_1515);
xnor U1605 (N_1605,N_1529,N_1541);
nand U1606 (N_1606,N_1569,N_1510);
nor U1607 (N_1607,N_1552,N_1556);
nor U1608 (N_1608,N_1545,N_1543);
and U1609 (N_1609,N_1562,N_1516);
nand U1610 (N_1610,N_1572,N_1506);
or U1611 (N_1611,N_1554,N_1514);
and U1612 (N_1612,N_1535,N_1552);
and U1613 (N_1613,N_1562,N_1502);
or U1614 (N_1614,N_1501,N_1543);
xor U1615 (N_1615,N_1539,N_1574);
nand U1616 (N_1616,N_1537,N_1502);
nor U1617 (N_1617,N_1531,N_1538);
or U1618 (N_1618,N_1528,N_1573);
nor U1619 (N_1619,N_1549,N_1531);
nor U1620 (N_1620,N_1537,N_1539);
nand U1621 (N_1621,N_1500,N_1536);
xnor U1622 (N_1622,N_1542,N_1514);
nor U1623 (N_1623,N_1545,N_1541);
nor U1624 (N_1624,N_1502,N_1554);
or U1625 (N_1625,N_1505,N_1510);
xnor U1626 (N_1626,N_1537,N_1559);
or U1627 (N_1627,N_1536,N_1505);
nor U1628 (N_1628,N_1519,N_1556);
or U1629 (N_1629,N_1574,N_1566);
nor U1630 (N_1630,N_1570,N_1568);
nor U1631 (N_1631,N_1573,N_1534);
or U1632 (N_1632,N_1574,N_1546);
nor U1633 (N_1633,N_1565,N_1548);
and U1634 (N_1634,N_1558,N_1510);
nand U1635 (N_1635,N_1532,N_1510);
nand U1636 (N_1636,N_1548,N_1536);
nor U1637 (N_1637,N_1501,N_1540);
xnor U1638 (N_1638,N_1521,N_1503);
nor U1639 (N_1639,N_1502,N_1572);
nor U1640 (N_1640,N_1510,N_1506);
nor U1641 (N_1641,N_1566,N_1511);
and U1642 (N_1642,N_1557,N_1520);
nor U1643 (N_1643,N_1502,N_1530);
and U1644 (N_1644,N_1507,N_1500);
and U1645 (N_1645,N_1538,N_1566);
and U1646 (N_1646,N_1505,N_1530);
nand U1647 (N_1647,N_1514,N_1568);
xnor U1648 (N_1648,N_1570,N_1500);
nor U1649 (N_1649,N_1541,N_1564);
and U1650 (N_1650,N_1613,N_1642);
nand U1651 (N_1651,N_1628,N_1601);
xor U1652 (N_1652,N_1609,N_1584);
and U1653 (N_1653,N_1643,N_1637);
and U1654 (N_1654,N_1624,N_1585);
nand U1655 (N_1655,N_1579,N_1644);
nand U1656 (N_1656,N_1626,N_1620);
and U1657 (N_1657,N_1600,N_1612);
or U1658 (N_1658,N_1615,N_1616);
or U1659 (N_1659,N_1593,N_1608);
and U1660 (N_1660,N_1583,N_1621);
nand U1661 (N_1661,N_1614,N_1631);
nor U1662 (N_1662,N_1599,N_1580);
nor U1663 (N_1663,N_1596,N_1581);
and U1664 (N_1664,N_1623,N_1597);
or U1665 (N_1665,N_1617,N_1606);
or U1666 (N_1666,N_1632,N_1587);
nor U1667 (N_1667,N_1594,N_1634);
or U1668 (N_1668,N_1638,N_1635);
and U1669 (N_1669,N_1611,N_1598);
and U1670 (N_1670,N_1619,N_1639);
nand U1671 (N_1671,N_1592,N_1618);
nand U1672 (N_1672,N_1627,N_1603);
or U1673 (N_1673,N_1640,N_1646);
nand U1674 (N_1674,N_1589,N_1625);
or U1675 (N_1675,N_1622,N_1647);
and U1676 (N_1676,N_1582,N_1586);
or U1677 (N_1677,N_1576,N_1578);
nor U1678 (N_1678,N_1575,N_1648);
or U1679 (N_1679,N_1633,N_1610);
nand U1680 (N_1680,N_1595,N_1636);
or U1681 (N_1681,N_1588,N_1645);
or U1682 (N_1682,N_1649,N_1604);
nand U1683 (N_1683,N_1629,N_1607);
and U1684 (N_1684,N_1590,N_1630);
and U1685 (N_1685,N_1605,N_1602);
or U1686 (N_1686,N_1577,N_1641);
and U1687 (N_1687,N_1591,N_1639);
and U1688 (N_1688,N_1629,N_1638);
nor U1689 (N_1689,N_1625,N_1607);
and U1690 (N_1690,N_1600,N_1617);
nor U1691 (N_1691,N_1645,N_1623);
nor U1692 (N_1692,N_1637,N_1617);
and U1693 (N_1693,N_1626,N_1601);
and U1694 (N_1694,N_1620,N_1621);
nand U1695 (N_1695,N_1638,N_1583);
nand U1696 (N_1696,N_1621,N_1642);
xor U1697 (N_1697,N_1606,N_1640);
and U1698 (N_1698,N_1610,N_1617);
nor U1699 (N_1699,N_1599,N_1584);
or U1700 (N_1700,N_1593,N_1595);
and U1701 (N_1701,N_1587,N_1592);
and U1702 (N_1702,N_1575,N_1642);
nor U1703 (N_1703,N_1635,N_1595);
nor U1704 (N_1704,N_1607,N_1603);
nand U1705 (N_1705,N_1596,N_1588);
nand U1706 (N_1706,N_1628,N_1577);
nor U1707 (N_1707,N_1636,N_1586);
nor U1708 (N_1708,N_1578,N_1648);
nor U1709 (N_1709,N_1639,N_1626);
or U1710 (N_1710,N_1601,N_1642);
or U1711 (N_1711,N_1594,N_1584);
nand U1712 (N_1712,N_1590,N_1611);
nand U1713 (N_1713,N_1629,N_1604);
or U1714 (N_1714,N_1645,N_1596);
and U1715 (N_1715,N_1585,N_1584);
and U1716 (N_1716,N_1585,N_1593);
nand U1717 (N_1717,N_1604,N_1625);
or U1718 (N_1718,N_1646,N_1612);
and U1719 (N_1719,N_1610,N_1645);
or U1720 (N_1720,N_1602,N_1581);
nand U1721 (N_1721,N_1613,N_1601);
and U1722 (N_1722,N_1627,N_1639);
nor U1723 (N_1723,N_1594,N_1590);
or U1724 (N_1724,N_1604,N_1607);
and U1725 (N_1725,N_1692,N_1695);
nor U1726 (N_1726,N_1654,N_1705);
and U1727 (N_1727,N_1703,N_1661);
nand U1728 (N_1728,N_1655,N_1702);
or U1729 (N_1729,N_1677,N_1665);
nand U1730 (N_1730,N_1681,N_1672);
nor U1731 (N_1731,N_1685,N_1678);
nor U1732 (N_1732,N_1673,N_1658);
nor U1733 (N_1733,N_1667,N_1724);
or U1734 (N_1734,N_1675,N_1723);
and U1735 (N_1735,N_1686,N_1704);
nor U1736 (N_1736,N_1669,N_1699);
and U1737 (N_1737,N_1722,N_1683);
or U1738 (N_1738,N_1684,N_1663);
xor U1739 (N_1739,N_1657,N_1662);
and U1740 (N_1740,N_1698,N_1690);
xnor U1741 (N_1741,N_1714,N_1660);
or U1742 (N_1742,N_1694,N_1720);
nand U1743 (N_1743,N_1652,N_1712);
nand U1744 (N_1744,N_1713,N_1680);
and U1745 (N_1745,N_1691,N_1659);
nand U1746 (N_1746,N_1711,N_1679);
or U1747 (N_1747,N_1671,N_1689);
nor U1748 (N_1748,N_1664,N_1651);
nand U1749 (N_1749,N_1650,N_1670);
nand U1750 (N_1750,N_1697,N_1674);
nor U1751 (N_1751,N_1676,N_1696);
and U1752 (N_1752,N_1706,N_1687);
xor U1753 (N_1753,N_1701,N_1688);
and U1754 (N_1754,N_1708,N_1656);
or U1755 (N_1755,N_1707,N_1716);
nand U1756 (N_1756,N_1653,N_1721);
or U1757 (N_1757,N_1682,N_1668);
or U1758 (N_1758,N_1700,N_1709);
or U1759 (N_1759,N_1666,N_1717);
xnor U1760 (N_1760,N_1710,N_1693);
or U1761 (N_1761,N_1715,N_1718);
nor U1762 (N_1762,N_1719,N_1724);
xnor U1763 (N_1763,N_1706,N_1691);
xor U1764 (N_1764,N_1674,N_1655);
nand U1765 (N_1765,N_1716,N_1658);
xor U1766 (N_1766,N_1652,N_1664);
and U1767 (N_1767,N_1712,N_1688);
nand U1768 (N_1768,N_1712,N_1665);
nand U1769 (N_1769,N_1685,N_1658);
nor U1770 (N_1770,N_1650,N_1683);
and U1771 (N_1771,N_1654,N_1717);
nor U1772 (N_1772,N_1667,N_1723);
and U1773 (N_1773,N_1669,N_1655);
and U1774 (N_1774,N_1714,N_1689);
or U1775 (N_1775,N_1693,N_1688);
nor U1776 (N_1776,N_1681,N_1650);
nand U1777 (N_1777,N_1721,N_1720);
or U1778 (N_1778,N_1669,N_1720);
nand U1779 (N_1779,N_1717,N_1724);
and U1780 (N_1780,N_1692,N_1667);
xnor U1781 (N_1781,N_1691,N_1686);
nor U1782 (N_1782,N_1721,N_1667);
nor U1783 (N_1783,N_1668,N_1698);
or U1784 (N_1784,N_1676,N_1674);
or U1785 (N_1785,N_1699,N_1671);
nand U1786 (N_1786,N_1696,N_1681);
or U1787 (N_1787,N_1661,N_1722);
or U1788 (N_1788,N_1692,N_1700);
and U1789 (N_1789,N_1669,N_1717);
or U1790 (N_1790,N_1719,N_1665);
nand U1791 (N_1791,N_1671,N_1723);
and U1792 (N_1792,N_1659,N_1710);
nor U1793 (N_1793,N_1699,N_1723);
nor U1794 (N_1794,N_1673,N_1698);
xor U1795 (N_1795,N_1706,N_1679);
nor U1796 (N_1796,N_1651,N_1724);
or U1797 (N_1797,N_1720,N_1674);
and U1798 (N_1798,N_1722,N_1651);
and U1799 (N_1799,N_1690,N_1691);
nand U1800 (N_1800,N_1733,N_1778);
or U1801 (N_1801,N_1793,N_1760);
nand U1802 (N_1802,N_1731,N_1757);
nand U1803 (N_1803,N_1725,N_1748);
nor U1804 (N_1804,N_1734,N_1795);
nor U1805 (N_1805,N_1736,N_1764);
and U1806 (N_1806,N_1744,N_1729);
and U1807 (N_1807,N_1763,N_1745);
nor U1808 (N_1808,N_1772,N_1771);
or U1809 (N_1809,N_1730,N_1762);
xor U1810 (N_1810,N_1759,N_1726);
nand U1811 (N_1811,N_1781,N_1796);
nand U1812 (N_1812,N_1773,N_1798);
and U1813 (N_1813,N_1766,N_1755);
nor U1814 (N_1814,N_1783,N_1784);
nand U1815 (N_1815,N_1782,N_1740);
nor U1816 (N_1816,N_1758,N_1732);
nand U1817 (N_1817,N_1727,N_1747);
nand U1818 (N_1818,N_1742,N_1797);
nor U1819 (N_1819,N_1787,N_1767);
or U1820 (N_1820,N_1749,N_1738);
and U1821 (N_1821,N_1791,N_1756);
and U1822 (N_1822,N_1753,N_1739);
nand U1823 (N_1823,N_1786,N_1754);
nor U1824 (N_1824,N_1777,N_1789);
or U1825 (N_1825,N_1728,N_1735);
nor U1826 (N_1826,N_1746,N_1765);
and U1827 (N_1827,N_1743,N_1741);
nand U1828 (N_1828,N_1790,N_1792);
and U1829 (N_1829,N_1770,N_1785);
and U1830 (N_1830,N_1794,N_1750);
and U1831 (N_1831,N_1799,N_1776);
nand U1832 (N_1832,N_1768,N_1751);
or U1833 (N_1833,N_1769,N_1775);
and U1834 (N_1834,N_1780,N_1774);
xor U1835 (N_1835,N_1737,N_1752);
nor U1836 (N_1836,N_1788,N_1761);
or U1837 (N_1837,N_1779,N_1760);
nor U1838 (N_1838,N_1729,N_1730);
nand U1839 (N_1839,N_1777,N_1781);
nand U1840 (N_1840,N_1750,N_1749);
nand U1841 (N_1841,N_1778,N_1768);
nand U1842 (N_1842,N_1774,N_1797);
xnor U1843 (N_1843,N_1748,N_1784);
nand U1844 (N_1844,N_1744,N_1759);
nor U1845 (N_1845,N_1764,N_1776);
nor U1846 (N_1846,N_1732,N_1737);
nor U1847 (N_1847,N_1769,N_1799);
nand U1848 (N_1848,N_1764,N_1766);
xnor U1849 (N_1849,N_1738,N_1785);
and U1850 (N_1850,N_1761,N_1736);
and U1851 (N_1851,N_1742,N_1766);
nand U1852 (N_1852,N_1791,N_1743);
nand U1853 (N_1853,N_1760,N_1764);
nor U1854 (N_1854,N_1763,N_1774);
nor U1855 (N_1855,N_1726,N_1755);
or U1856 (N_1856,N_1774,N_1771);
and U1857 (N_1857,N_1786,N_1739);
or U1858 (N_1858,N_1750,N_1760);
or U1859 (N_1859,N_1791,N_1739);
and U1860 (N_1860,N_1771,N_1745);
or U1861 (N_1861,N_1798,N_1748);
xor U1862 (N_1862,N_1776,N_1771);
and U1863 (N_1863,N_1785,N_1745);
or U1864 (N_1864,N_1748,N_1778);
nor U1865 (N_1865,N_1779,N_1773);
nand U1866 (N_1866,N_1745,N_1755);
nand U1867 (N_1867,N_1751,N_1732);
or U1868 (N_1868,N_1731,N_1785);
nor U1869 (N_1869,N_1746,N_1738);
or U1870 (N_1870,N_1771,N_1783);
xnor U1871 (N_1871,N_1733,N_1749);
nand U1872 (N_1872,N_1767,N_1765);
and U1873 (N_1873,N_1731,N_1736);
nor U1874 (N_1874,N_1748,N_1794);
and U1875 (N_1875,N_1825,N_1858);
nand U1876 (N_1876,N_1869,N_1817);
nor U1877 (N_1877,N_1826,N_1863);
nand U1878 (N_1878,N_1846,N_1840);
and U1879 (N_1879,N_1850,N_1832);
nand U1880 (N_1880,N_1874,N_1865);
nand U1881 (N_1881,N_1824,N_1864);
and U1882 (N_1882,N_1813,N_1815);
and U1883 (N_1883,N_1816,N_1828);
or U1884 (N_1884,N_1802,N_1812);
nand U1885 (N_1885,N_1857,N_1800);
and U1886 (N_1886,N_1809,N_1873);
nand U1887 (N_1887,N_1862,N_1849);
xnor U1888 (N_1888,N_1829,N_1838);
nand U1889 (N_1889,N_1867,N_1835);
and U1890 (N_1890,N_1856,N_1806);
and U1891 (N_1891,N_1855,N_1811);
and U1892 (N_1892,N_1861,N_1804);
and U1893 (N_1893,N_1851,N_1836);
nand U1894 (N_1894,N_1827,N_1848);
nor U1895 (N_1895,N_1833,N_1843);
or U1896 (N_1896,N_1868,N_1818);
nor U1897 (N_1897,N_1810,N_1820);
nand U1898 (N_1898,N_1866,N_1844);
nand U1899 (N_1899,N_1805,N_1814);
nor U1900 (N_1900,N_1837,N_1872);
nand U1901 (N_1901,N_1847,N_1808);
nand U1902 (N_1902,N_1807,N_1845);
nor U1903 (N_1903,N_1803,N_1852);
xor U1904 (N_1904,N_1853,N_1860);
nand U1905 (N_1905,N_1819,N_1859);
and U1906 (N_1906,N_1841,N_1871);
and U1907 (N_1907,N_1823,N_1834);
nor U1908 (N_1908,N_1870,N_1830);
and U1909 (N_1909,N_1822,N_1854);
nand U1910 (N_1910,N_1839,N_1821);
nand U1911 (N_1911,N_1801,N_1831);
and U1912 (N_1912,N_1842,N_1859);
nand U1913 (N_1913,N_1869,N_1810);
and U1914 (N_1914,N_1802,N_1820);
nor U1915 (N_1915,N_1820,N_1873);
and U1916 (N_1916,N_1813,N_1873);
nor U1917 (N_1917,N_1804,N_1860);
nand U1918 (N_1918,N_1804,N_1864);
nand U1919 (N_1919,N_1868,N_1861);
nor U1920 (N_1920,N_1865,N_1822);
nand U1921 (N_1921,N_1845,N_1819);
nor U1922 (N_1922,N_1825,N_1874);
xor U1923 (N_1923,N_1834,N_1849);
and U1924 (N_1924,N_1814,N_1804);
nor U1925 (N_1925,N_1847,N_1837);
or U1926 (N_1926,N_1862,N_1848);
or U1927 (N_1927,N_1845,N_1835);
and U1928 (N_1928,N_1810,N_1802);
and U1929 (N_1929,N_1854,N_1812);
or U1930 (N_1930,N_1828,N_1826);
or U1931 (N_1931,N_1859,N_1850);
nor U1932 (N_1932,N_1833,N_1821);
nand U1933 (N_1933,N_1869,N_1838);
or U1934 (N_1934,N_1864,N_1818);
or U1935 (N_1935,N_1839,N_1828);
and U1936 (N_1936,N_1807,N_1804);
nor U1937 (N_1937,N_1827,N_1858);
nor U1938 (N_1938,N_1845,N_1867);
and U1939 (N_1939,N_1800,N_1817);
or U1940 (N_1940,N_1808,N_1812);
and U1941 (N_1941,N_1809,N_1844);
nor U1942 (N_1942,N_1802,N_1860);
or U1943 (N_1943,N_1874,N_1861);
xnor U1944 (N_1944,N_1866,N_1822);
nor U1945 (N_1945,N_1864,N_1853);
and U1946 (N_1946,N_1864,N_1846);
xnor U1947 (N_1947,N_1840,N_1863);
xor U1948 (N_1948,N_1867,N_1836);
or U1949 (N_1949,N_1851,N_1809);
and U1950 (N_1950,N_1894,N_1938);
and U1951 (N_1951,N_1905,N_1944);
nand U1952 (N_1952,N_1902,N_1877);
nor U1953 (N_1953,N_1925,N_1935);
or U1954 (N_1954,N_1879,N_1886);
or U1955 (N_1955,N_1949,N_1904);
nor U1956 (N_1956,N_1932,N_1890);
nand U1957 (N_1957,N_1926,N_1931);
or U1958 (N_1958,N_1878,N_1948);
nor U1959 (N_1959,N_1939,N_1891);
nor U1960 (N_1960,N_1896,N_1934);
xor U1961 (N_1961,N_1919,N_1895);
nor U1962 (N_1962,N_1882,N_1947);
or U1963 (N_1963,N_1916,N_1912);
nor U1964 (N_1964,N_1881,N_1900);
nand U1965 (N_1965,N_1918,N_1883);
and U1966 (N_1966,N_1880,N_1897);
and U1967 (N_1967,N_1941,N_1910);
nor U1968 (N_1968,N_1913,N_1914);
nand U1969 (N_1969,N_1887,N_1917);
nor U1970 (N_1970,N_1923,N_1922);
nand U1971 (N_1971,N_1940,N_1936);
nor U1972 (N_1972,N_1898,N_1911);
nand U1973 (N_1973,N_1893,N_1892);
nor U1974 (N_1974,N_1933,N_1901);
nor U1975 (N_1975,N_1908,N_1937);
nand U1976 (N_1976,N_1942,N_1876);
and U1977 (N_1977,N_1885,N_1884);
nand U1978 (N_1978,N_1920,N_1915);
nor U1979 (N_1979,N_1899,N_1903);
nor U1980 (N_1980,N_1909,N_1945);
nand U1981 (N_1981,N_1875,N_1907);
or U1982 (N_1982,N_1928,N_1906);
or U1983 (N_1983,N_1888,N_1889);
and U1984 (N_1984,N_1924,N_1946);
xnor U1985 (N_1985,N_1921,N_1943);
nand U1986 (N_1986,N_1929,N_1927);
and U1987 (N_1987,N_1930,N_1913);
nand U1988 (N_1988,N_1902,N_1926);
nand U1989 (N_1989,N_1927,N_1883);
nor U1990 (N_1990,N_1937,N_1935);
xor U1991 (N_1991,N_1875,N_1942);
and U1992 (N_1992,N_1924,N_1879);
xor U1993 (N_1993,N_1921,N_1900);
nor U1994 (N_1994,N_1895,N_1947);
nand U1995 (N_1995,N_1920,N_1882);
nand U1996 (N_1996,N_1903,N_1913);
nand U1997 (N_1997,N_1949,N_1916);
or U1998 (N_1998,N_1938,N_1939);
xor U1999 (N_1999,N_1883,N_1891);
nor U2000 (N_2000,N_1939,N_1906);
and U2001 (N_2001,N_1912,N_1875);
nor U2002 (N_2002,N_1942,N_1897);
or U2003 (N_2003,N_1938,N_1921);
nor U2004 (N_2004,N_1927,N_1919);
nand U2005 (N_2005,N_1902,N_1886);
or U2006 (N_2006,N_1908,N_1882);
or U2007 (N_2007,N_1943,N_1897);
and U2008 (N_2008,N_1946,N_1942);
or U2009 (N_2009,N_1943,N_1898);
xor U2010 (N_2010,N_1946,N_1907);
nand U2011 (N_2011,N_1898,N_1920);
nand U2012 (N_2012,N_1905,N_1901);
or U2013 (N_2013,N_1936,N_1948);
xnor U2014 (N_2014,N_1935,N_1880);
nor U2015 (N_2015,N_1933,N_1936);
nor U2016 (N_2016,N_1935,N_1895);
nor U2017 (N_2017,N_1897,N_1886);
or U2018 (N_2018,N_1883,N_1947);
and U2019 (N_2019,N_1928,N_1877);
nand U2020 (N_2020,N_1926,N_1949);
or U2021 (N_2021,N_1898,N_1949);
nor U2022 (N_2022,N_1904,N_1899);
nand U2023 (N_2023,N_1884,N_1923);
xnor U2024 (N_2024,N_1887,N_1877);
nor U2025 (N_2025,N_2024,N_1970);
and U2026 (N_2026,N_1958,N_1951);
and U2027 (N_2027,N_1953,N_1990);
xnor U2028 (N_2028,N_1974,N_1980);
or U2029 (N_2029,N_1978,N_1979);
nor U2030 (N_2030,N_1999,N_1998);
xnor U2031 (N_2031,N_1956,N_1960);
and U2032 (N_2032,N_2003,N_1969);
xor U2033 (N_2033,N_1977,N_1972);
and U2034 (N_2034,N_2012,N_2021);
xor U2035 (N_2035,N_1997,N_1963);
and U2036 (N_2036,N_2019,N_2007);
xor U2037 (N_2037,N_1959,N_2014);
xor U2038 (N_2038,N_1986,N_1996);
nor U2039 (N_2039,N_2017,N_2005);
nand U2040 (N_2040,N_1966,N_1985);
nand U2041 (N_2041,N_1961,N_1991);
xnor U2042 (N_2042,N_2018,N_2016);
and U2043 (N_2043,N_1962,N_1994);
or U2044 (N_2044,N_1989,N_1976);
nor U2045 (N_2045,N_2015,N_2013);
or U2046 (N_2046,N_2010,N_1995);
or U2047 (N_2047,N_2004,N_2000);
and U2048 (N_2048,N_2011,N_2008);
xor U2049 (N_2049,N_1950,N_1971);
or U2050 (N_2050,N_1992,N_1954);
nor U2051 (N_2051,N_1981,N_1968);
xor U2052 (N_2052,N_1984,N_1993);
and U2053 (N_2053,N_1965,N_1975);
nor U2054 (N_2054,N_2023,N_1988);
nand U2055 (N_2055,N_2009,N_1952);
nor U2056 (N_2056,N_1957,N_1955);
nand U2057 (N_2057,N_1987,N_2006);
xnor U2058 (N_2058,N_2001,N_2002);
nand U2059 (N_2059,N_2022,N_1983);
nor U2060 (N_2060,N_1973,N_1964);
xnor U2061 (N_2061,N_1967,N_1982);
nand U2062 (N_2062,N_2020,N_1974);
and U2063 (N_2063,N_1971,N_1958);
and U2064 (N_2064,N_1954,N_1972);
nor U2065 (N_2065,N_2001,N_2013);
nand U2066 (N_2066,N_2007,N_2001);
nor U2067 (N_2067,N_1962,N_1970);
or U2068 (N_2068,N_1956,N_1992);
or U2069 (N_2069,N_2001,N_1968);
xnor U2070 (N_2070,N_1976,N_2024);
and U2071 (N_2071,N_2012,N_1964);
and U2072 (N_2072,N_1997,N_1973);
nor U2073 (N_2073,N_1984,N_1954);
nand U2074 (N_2074,N_1972,N_2011);
nand U2075 (N_2075,N_1974,N_2011);
nor U2076 (N_2076,N_1980,N_2019);
nand U2077 (N_2077,N_2004,N_1993);
xor U2078 (N_2078,N_1987,N_1983);
xnor U2079 (N_2079,N_1963,N_2010);
and U2080 (N_2080,N_1983,N_2003);
nand U2081 (N_2081,N_1965,N_1997);
and U2082 (N_2082,N_1960,N_2007);
and U2083 (N_2083,N_1999,N_2011);
and U2084 (N_2084,N_1952,N_1984);
and U2085 (N_2085,N_1978,N_1991);
nor U2086 (N_2086,N_1989,N_2021);
and U2087 (N_2087,N_1987,N_1999);
and U2088 (N_2088,N_2020,N_1994);
or U2089 (N_2089,N_1989,N_1971);
and U2090 (N_2090,N_1993,N_1977);
nand U2091 (N_2091,N_2011,N_2010);
and U2092 (N_2092,N_2008,N_1997);
or U2093 (N_2093,N_1978,N_2012);
or U2094 (N_2094,N_1988,N_1984);
and U2095 (N_2095,N_1952,N_1976);
or U2096 (N_2096,N_2015,N_2008);
or U2097 (N_2097,N_1956,N_1950);
or U2098 (N_2098,N_2013,N_2018);
xnor U2099 (N_2099,N_1978,N_1981);
and U2100 (N_2100,N_2059,N_2070);
nand U2101 (N_2101,N_2079,N_2078);
nand U2102 (N_2102,N_2082,N_2095);
nand U2103 (N_2103,N_2034,N_2049);
or U2104 (N_2104,N_2098,N_2029);
or U2105 (N_2105,N_2047,N_2061);
and U2106 (N_2106,N_2035,N_2076);
and U2107 (N_2107,N_2064,N_2072);
or U2108 (N_2108,N_2068,N_2092);
nand U2109 (N_2109,N_2037,N_2045);
nor U2110 (N_2110,N_2032,N_2054);
and U2111 (N_2111,N_2067,N_2027);
or U2112 (N_2112,N_2093,N_2089);
and U2113 (N_2113,N_2058,N_2066);
nand U2114 (N_2114,N_2087,N_2084);
or U2115 (N_2115,N_2083,N_2099);
xnor U2116 (N_2116,N_2086,N_2056);
or U2117 (N_2117,N_2030,N_2055);
nand U2118 (N_2118,N_2060,N_2065);
nor U2119 (N_2119,N_2036,N_2080);
nor U2120 (N_2120,N_2085,N_2042);
xor U2121 (N_2121,N_2028,N_2025);
and U2122 (N_2122,N_2040,N_2094);
and U2123 (N_2123,N_2075,N_2091);
nand U2124 (N_2124,N_2053,N_2026);
or U2125 (N_2125,N_2044,N_2074);
nor U2126 (N_2126,N_2088,N_2063);
and U2127 (N_2127,N_2077,N_2033);
and U2128 (N_2128,N_2097,N_2051);
and U2129 (N_2129,N_2071,N_2073);
nor U2130 (N_2130,N_2081,N_2043);
nand U2131 (N_2131,N_2031,N_2069);
nor U2132 (N_2132,N_2039,N_2046);
nand U2133 (N_2133,N_2090,N_2052);
nor U2134 (N_2134,N_2038,N_2041);
nor U2135 (N_2135,N_2096,N_2050);
or U2136 (N_2136,N_2062,N_2048);
or U2137 (N_2137,N_2057,N_2070);
and U2138 (N_2138,N_2043,N_2091);
nor U2139 (N_2139,N_2043,N_2073);
nor U2140 (N_2140,N_2048,N_2033);
and U2141 (N_2141,N_2088,N_2067);
nand U2142 (N_2142,N_2036,N_2055);
nand U2143 (N_2143,N_2035,N_2063);
nand U2144 (N_2144,N_2083,N_2046);
or U2145 (N_2145,N_2077,N_2072);
and U2146 (N_2146,N_2078,N_2080);
nand U2147 (N_2147,N_2065,N_2078);
and U2148 (N_2148,N_2091,N_2085);
or U2149 (N_2149,N_2088,N_2037);
or U2150 (N_2150,N_2037,N_2065);
or U2151 (N_2151,N_2097,N_2083);
nor U2152 (N_2152,N_2074,N_2057);
and U2153 (N_2153,N_2037,N_2027);
or U2154 (N_2154,N_2076,N_2061);
and U2155 (N_2155,N_2056,N_2029);
or U2156 (N_2156,N_2029,N_2067);
nand U2157 (N_2157,N_2059,N_2035);
or U2158 (N_2158,N_2037,N_2079);
nor U2159 (N_2159,N_2093,N_2045);
xnor U2160 (N_2160,N_2025,N_2060);
or U2161 (N_2161,N_2079,N_2076);
nor U2162 (N_2162,N_2075,N_2029);
or U2163 (N_2163,N_2031,N_2071);
or U2164 (N_2164,N_2039,N_2082);
nor U2165 (N_2165,N_2099,N_2061);
nand U2166 (N_2166,N_2040,N_2056);
nand U2167 (N_2167,N_2029,N_2078);
nor U2168 (N_2168,N_2077,N_2027);
and U2169 (N_2169,N_2086,N_2036);
nand U2170 (N_2170,N_2068,N_2032);
and U2171 (N_2171,N_2050,N_2039);
and U2172 (N_2172,N_2095,N_2076);
xor U2173 (N_2173,N_2097,N_2092);
or U2174 (N_2174,N_2047,N_2065);
nand U2175 (N_2175,N_2168,N_2166);
and U2176 (N_2176,N_2108,N_2136);
nor U2177 (N_2177,N_2118,N_2172);
xnor U2178 (N_2178,N_2115,N_2127);
and U2179 (N_2179,N_2155,N_2116);
nor U2180 (N_2180,N_2154,N_2117);
xor U2181 (N_2181,N_2124,N_2107);
and U2182 (N_2182,N_2125,N_2169);
and U2183 (N_2183,N_2164,N_2132);
and U2184 (N_2184,N_2129,N_2149);
and U2185 (N_2185,N_2148,N_2141);
nand U2186 (N_2186,N_2126,N_2156);
or U2187 (N_2187,N_2103,N_2174);
nor U2188 (N_2188,N_2133,N_2111);
and U2189 (N_2189,N_2145,N_2113);
nand U2190 (N_2190,N_2173,N_2144);
xor U2191 (N_2191,N_2160,N_2146);
nand U2192 (N_2192,N_2162,N_2139);
nor U2193 (N_2193,N_2143,N_2142);
nand U2194 (N_2194,N_2120,N_2106);
or U2195 (N_2195,N_2128,N_2147);
and U2196 (N_2196,N_2135,N_2151);
nor U2197 (N_2197,N_2170,N_2140);
or U2198 (N_2198,N_2153,N_2130);
nor U2199 (N_2199,N_2102,N_2123);
and U2200 (N_2200,N_2157,N_2110);
xnor U2201 (N_2201,N_2112,N_2161);
nand U2202 (N_2202,N_2158,N_2104);
nand U2203 (N_2203,N_2137,N_2109);
and U2204 (N_2204,N_2114,N_2150);
nand U2205 (N_2205,N_2101,N_2121);
or U2206 (N_2206,N_2131,N_2152);
and U2207 (N_2207,N_2134,N_2119);
or U2208 (N_2208,N_2167,N_2138);
nor U2209 (N_2209,N_2105,N_2171);
nand U2210 (N_2210,N_2165,N_2163);
nor U2211 (N_2211,N_2100,N_2159);
nor U2212 (N_2212,N_2122,N_2129);
nor U2213 (N_2213,N_2124,N_2163);
and U2214 (N_2214,N_2114,N_2141);
and U2215 (N_2215,N_2105,N_2106);
and U2216 (N_2216,N_2174,N_2134);
or U2217 (N_2217,N_2115,N_2158);
and U2218 (N_2218,N_2153,N_2158);
or U2219 (N_2219,N_2163,N_2100);
or U2220 (N_2220,N_2166,N_2134);
and U2221 (N_2221,N_2135,N_2122);
nand U2222 (N_2222,N_2171,N_2114);
and U2223 (N_2223,N_2173,N_2133);
and U2224 (N_2224,N_2167,N_2139);
xnor U2225 (N_2225,N_2129,N_2164);
and U2226 (N_2226,N_2172,N_2140);
and U2227 (N_2227,N_2124,N_2137);
nor U2228 (N_2228,N_2124,N_2134);
and U2229 (N_2229,N_2141,N_2125);
and U2230 (N_2230,N_2118,N_2159);
nand U2231 (N_2231,N_2137,N_2166);
nor U2232 (N_2232,N_2122,N_2132);
and U2233 (N_2233,N_2151,N_2136);
and U2234 (N_2234,N_2121,N_2120);
nor U2235 (N_2235,N_2110,N_2163);
and U2236 (N_2236,N_2147,N_2172);
xor U2237 (N_2237,N_2131,N_2169);
nand U2238 (N_2238,N_2132,N_2100);
or U2239 (N_2239,N_2105,N_2165);
or U2240 (N_2240,N_2164,N_2144);
xnor U2241 (N_2241,N_2144,N_2138);
nor U2242 (N_2242,N_2119,N_2115);
xor U2243 (N_2243,N_2150,N_2107);
or U2244 (N_2244,N_2104,N_2149);
nor U2245 (N_2245,N_2145,N_2148);
xor U2246 (N_2246,N_2145,N_2165);
and U2247 (N_2247,N_2158,N_2118);
nand U2248 (N_2248,N_2126,N_2167);
or U2249 (N_2249,N_2157,N_2109);
nor U2250 (N_2250,N_2228,N_2209);
nor U2251 (N_2251,N_2212,N_2224);
nand U2252 (N_2252,N_2179,N_2177);
nor U2253 (N_2253,N_2241,N_2186);
nand U2254 (N_2254,N_2200,N_2227);
xnor U2255 (N_2255,N_2182,N_2226);
or U2256 (N_2256,N_2229,N_2244);
nand U2257 (N_2257,N_2237,N_2240);
and U2258 (N_2258,N_2183,N_2184);
or U2259 (N_2259,N_2232,N_2203);
and U2260 (N_2260,N_2198,N_2202);
and U2261 (N_2261,N_2195,N_2234);
nand U2262 (N_2262,N_2180,N_2216);
and U2263 (N_2263,N_2235,N_2213);
nand U2264 (N_2264,N_2219,N_2178);
nor U2265 (N_2265,N_2205,N_2221);
nor U2266 (N_2266,N_2242,N_2194);
nor U2267 (N_2267,N_2233,N_2220);
and U2268 (N_2268,N_2238,N_2181);
and U2269 (N_2269,N_2231,N_2239);
nor U2270 (N_2270,N_2225,N_2197);
nor U2271 (N_2271,N_2185,N_2176);
or U2272 (N_2272,N_2223,N_2210);
or U2273 (N_2273,N_2214,N_2199);
nor U2274 (N_2274,N_2222,N_2245);
nor U2275 (N_2275,N_2175,N_2192);
nand U2276 (N_2276,N_2201,N_2188);
nand U2277 (N_2277,N_2196,N_2215);
or U2278 (N_2278,N_2190,N_2230);
nand U2279 (N_2279,N_2247,N_2236);
nor U2280 (N_2280,N_2243,N_2217);
or U2281 (N_2281,N_2249,N_2187);
and U2282 (N_2282,N_2207,N_2189);
and U2283 (N_2283,N_2248,N_2191);
or U2284 (N_2284,N_2208,N_2204);
nor U2285 (N_2285,N_2246,N_2211);
nand U2286 (N_2286,N_2206,N_2193);
xor U2287 (N_2287,N_2218,N_2249);
and U2288 (N_2288,N_2218,N_2229);
xor U2289 (N_2289,N_2233,N_2198);
and U2290 (N_2290,N_2243,N_2221);
nor U2291 (N_2291,N_2178,N_2194);
or U2292 (N_2292,N_2239,N_2210);
nand U2293 (N_2293,N_2181,N_2219);
xor U2294 (N_2294,N_2189,N_2211);
nand U2295 (N_2295,N_2234,N_2194);
xor U2296 (N_2296,N_2213,N_2185);
and U2297 (N_2297,N_2195,N_2196);
or U2298 (N_2298,N_2225,N_2217);
and U2299 (N_2299,N_2238,N_2212);
nor U2300 (N_2300,N_2216,N_2200);
nand U2301 (N_2301,N_2243,N_2180);
nand U2302 (N_2302,N_2213,N_2236);
nand U2303 (N_2303,N_2220,N_2184);
and U2304 (N_2304,N_2196,N_2184);
nor U2305 (N_2305,N_2215,N_2214);
or U2306 (N_2306,N_2217,N_2240);
nand U2307 (N_2307,N_2247,N_2222);
or U2308 (N_2308,N_2189,N_2244);
or U2309 (N_2309,N_2187,N_2182);
nand U2310 (N_2310,N_2205,N_2185);
xor U2311 (N_2311,N_2206,N_2240);
nand U2312 (N_2312,N_2203,N_2215);
nor U2313 (N_2313,N_2194,N_2203);
xnor U2314 (N_2314,N_2241,N_2225);
xnor U2315 (N_2315,N_2189,N_2246);
nand U2316 (N_2316,N_2187,N_2226);
nor U2317 (N_2317,N_2209,N_2185);
nor U2318 (N_2318,N_2195,N_2219);
or U2319 (N_2319,N_2189,N_2243);
nor U2320 (N_2320,N_2244,N_2221);
or U2321 (N_2321,N_2193,N_2228);
xnor U2322 (N_2322,N_2211,N_2245);
nor U2323 (N_2323,N_2191,N_2197);
or U2324 (N_2324,N_2203,N_2199);
and U2325 (N_2325,N_2267,N_2323);
nand U2326 (N_2326,N_2278,N_2263);
nand U2327 (N_2327,N_2298,N_2307);
xor U2328 (N_2328,N_2276,N_2320);
nand U2329 (N_2329,N_2308,N_2288);
or U2330 (N_2330,N_2268,N_2314);
nand U2331 (N_2331,N_2275,N_2277);
or U2332 (N_2332,N_2262,N_2319);
or U2333 (N_2333,N_2261,N_2271);
nor U2334 (N_2334,N_2272,N_2291);
nor U2335 (N_2335,N_2257,N_2282);
nand U2336 (N_2336,N_2252,N_2316);
and U2337 (N_2337,N_2259,N_2281);
and U2338 (N_2338,N_2300,N_2250);
and U2339 (N_2339,N_2321,N_2254);
nand U2340 (N_2340,N_2292,N_2301);
nand U2341 (N_2341,N_2309,N_2286);
or U2342 (N_2342,N_2284,N_2310);
nor U2343 (N_2343,N_2273,N_2280);
xnor U2344 (N_2344,N_2260,N_2285);
and U2345 (N_2345,N_2304,N_2306);
or U2346 (N_2346,N_2303,N_2322);
nand U2347 (N_2347,N_2269,N_2256);
and U2348 (N_2348,N_2253,N_2274);
xor U2349 (N_2349,N_2299,N_2294);
nand U2350 (N_2350,N_2290,N_2305);
or U2351 (N_2351,N_2311,N_2324);
or U2352 (N_2352,N_2317,N_2279);
nor U2353 (N_2353,N_2270,N_2266);
nor U2354 (N_2354,N_2265,N_2255);
xnor U2355 (N_2355,N_2312,N_2251);
nand U2356 (N_2356,N_2258,N_2293);
nor U2357 (N_2357,N_2318,N_2295);
or U2358 (N_2358,N_2264,N_2296);
nand U2359 (N_2359,N_2302,N_2283);
nand U2360 (N_2360,N_2313,N_2289);
xor U2361 (N_2361,N_2315,N_2297);
and U2362 (N_2362,N_2287,N_2290);
or U2363 (N_2363,N_2265,N_2260);
and U2364 (N_2364,N_2285,N_2261);
nor U2365 (N_2365,N_2299,N_2319);
or U2366 (N_2366,N_2281,N_2300);
nor U2367 (N_2367,N_2306,N_2280);
nor U2368 (N_2368,N_2289,N_2292);
and U2369 (N_2369,N_2288,N_2312);
xnor U2370 (N_2370,N_2295,N_2308);
nor U2371 (N_2371,N_2286,N_2319);
nor U2372 (N_2372,N_2264,N_2265);
or U2373 (N_2373,N_2273,N_2302);
nor U2374 (N_2374,N_2250,N_2274);
or U2375 (N_2375,N_2313,N_2295);
and U2376 (N_2376,N_2324,N_2310);
and U2377 (N_2377,N_2309,N_2312);
nand U2378 (N_2378,N_2288,N_2305);
or U2379 (N_2379,N_2322,N_2281);
nand U2380 (N_2380,N_2252,N_2287);
nand U2381 (N_2381,N_2299,N_2312);
nor U2382 (N_2382,N_2297,N_2269);
nand U2383 (N_2383,N_2311,N_2317);
nand U2384 (N_2384,N_2315,N_2287);
nand U2385 (N_2385,N_2257,N_2320);
nor U2386 (N_2386,N_2311,N_2277);
nor U2387 (N_2387,N_2300,N_2302);
and U2388 (N_2388,N_2277,N_2269);
nand U2389 (N_2389,N_2297,N_2305);
nand U2390 (N_2390,N_2322,N_2301);
nand U2391 (N_2391,N_2294,N_2275);
nor U2392 (N_2392,N_2286,N_2280);
xnor U2393 (N_2393,N_2281,N_2262);
nand U2394 (N_2394,N_2259,N_2322);
xnor U2395 (N_2395,N_2309,N_2310);
nand U2396 (N_2396,N_2277,N_2253);
and U2397 (N_2397,N_2271,N_2288);
xor U2398 (N_2398,N_2314,N_2305);
nor U2399 (N_2399,N_2303,N_2277);
nand U2400 (N_2400,N_2362,N_2382);
or U2401 (N_2401,N_2343,N_2365);
or U2402 (N_2402,N_2374,N_2330);
or U2403 (N_2403,N_2370,N_2334);
or U2404 (N_2404,N_2375,N_2331);
nor U2405 (N_2405,N_2391,N_2350);
xnor U2406 (N_2406,N_2371,N_2329);
and U2407 (N_2407,N_2372,N_2361);
xor U2408 (N_2408,N_2363,N_2342);
and U2409 (N_2409,N_2393,N_2351);
nand U2410 (N_2410,N_2373,N_2390);
and U2411 (N_2411,N_2385,N_2392);
or U2412 (N_2412,N_2366,N_2388);
xnor U2413 (N_2413,N_2358,N_2356);
xnor U2414 (N_2414,N_2338,N_2367);
nor U2415 (N_2415,N_2387,N_2341);
and U2416 (N_2416,N_2359,N_2339);
and U2417 (N_2417,N_2354,N_2369);
and U2418 (N_2418,N_2325,N_2353);
nor U2419 (N_2419,N_2397,N_2333);
nand U2420 (N_2420,N_2386,N_2376);
and U2421 (N_2421,N_2360,N_2368);
or U2422 (N_2422,N_2337,N_2344);
nand U2423 (N_2423,N_2346,N_2377);
nand U2424 (N_2424,N_2380,N_2335);
nand U2425 (N_2425,N_2357,N_2399);
and U2426 (N_2426,N_2383,N_2355);
nor U2427 (N_2427,N_2332,N_2395);
nand U2428 (N_2428,N_2396,N_2347);
nand U2429 (N_2429,N_2381,N_2398);
xor U2430 (N_2430,N_2348,N_2378);
and U2431 (N_2431,N_2384,N_2364);
nand U2432 (N_2432,N_2327,N_2340);
nand U2433 (N_2433,N_2352,N_2328);
and U2434 (N_2434,N_2326,N_2394);
xnor U2435 (N_2435,N_2345,N_2389);
or U2436 (N_2436,N_2379,N_2336);
or U2437 (N_2437,N_2349,N_2356);
and U2438 (N_2438,N_2365,N_2361);
and U2439 (N_2439,N_2338,N_2361);
nand U2440 (N_2440,N_2354,N_2340);
and U2441 (N_2441,N_2388,N_2395);
nor U2442 (N_2442,N_2347,N_2363);
or U2443 (N_2443,N_2358,N_2363);
and U2444 (N_2444,N_2349,N_2354);
nor U2445 (N_2445,N_2398,N_2328);
and U2446 (N_2446,N_2338,N_2327);
or U2447 (N_2447,N_2381,N_2388);
or U2448 (N_2448,N_2350,N_2373);
xnor U2449 (N_2449,N_2349,N_2350);
nor U2450 (N_2450,N_2348,N_2343);
nor U2451 (N_2451,N_2391,N_2345);
or U2452 (N_2452,N_2397,N_2334);
and U2453 (N_2453,N_2359,N_2325);
or U2454 (N_2454,N_2359,N_2374);
or U2455 (N_2455,N_2362,N_2337);
or U2456 (N_2456,N_2371,N_2352);
or U2457 (N_2457,N_2356,N_2331);
nand U2458 (N_2458,N_2339,N_2364);
or U2459 (N_2459,N_2376,N_2380);
and U2460 (N_2460,N_2360,N_2330);
and U2461 (N_2461,N_2354,N_2362);
nand U2462 (N_2462,N_2365,N_2386);
or U2463 (N_2463,N_2370,N_2344);
xnor U2464 (N_2464,N_2337,N_2336);
nand U2465 (N_2465,N_2378,N_2346);
and U2466 (N_2466,N_2356,N_2341);
nand U2467 (N_2467,N_2379,N_2337);
nand U2468 (N_2468,N_2351,N_2352);
or U2469 (N_2469,N_2359,N_2392);
or U2470 (N_2470,N_2344,N_2396);
and U2471 (N_2471,N_2389,N_2387);
and U2472 (N_2472,N_2383,N_2398);
and U2473 (N_2473,N_2363,N_2372);
nand U2474 (N_2474,N_2380,N_2374);
or U2475 (N_2475,N_2462,N_2436);
xor U2476 (N_2476,N_2467,N_2411);
and U2477 (N_2477,N_2458,N_2430);
and U2478 (N_2478,N_2423,N_2419);
nor U2479 (N_2479,N_2473,N_2457);
or U2480 (N_2480,N_2474,N_2422);
nand U2481 (N_2481,N_2460,N_2447);
nand U2482 (N_2482,N_2409,N_2412);
or U2483 (N_2483,N_2463,N_2407);
and U2484 (N_2484,N_2414,N_2421);
nor U2485 (N_2485,N_2404,N_2410);
nand U2486 (N_2486,N_2459,N_2429);
nor U2487 (N_2487,N_2431,N_2468);
and U2488 (N_2488,N_2442,N_2453);
and U2489 (N_2489,N_2413,N_2452);
nor U2490 (N_2490,N_2441,N_2425);
nor U2491 (N_2491,N_2433,N_2440);
and U2492 (N_2492,N_2466,N_2444);
and U2493 (N_2493,N_2432,N_2405);
nand U2494 (N_2494,N_2445,N_2456);
nor U2495 (N_2495,N_2449,N_2408);
nor U2496 (N_2496,N_2434,N_2446);
nand U2497 (N_2497,N_2426,N_2471);
and U2498 (N_2498,N_2427,N_2435);
or U2499 (N_2499,N_2437,N_2400);
nand U2500 (N_2500,N_2401,N_2428);
or U2501 (N_2501,N_2406,N_2438);
or U2502 (N_2502,N_2464,N_2415);
nand U2503 (N_2503,N_2451,N_2424);
nand U2504 (N_2504,N_2461,N_2418);
nor U2505 (N_2505,N_2465,N_2416);
and U2506 (N_2506,N_2455,N_2469);
or U2507 (N_2507,N_2448,N_2402);
nor U2508 (N_2508,N_2443,N_2439);
and U2509 (N_2509,N_2420,N_2454);
nor U2510 (N_2510,N_2403,N_2450);
nand U2511 (N_2511,N_2472,N_2417);
xnor U2512 (N_2512,N_2470,N_2434);
nand U2513 (N_2513,N_2447,N_2435);
nand U2514 (N_2514,N_2441,N_2455);
and U2515 (N_2515,N_2411,N_2459);
nor U2516 (N_2516,N_2471,N_2419);
or U2517 (N_2517,N_2465,N_2456);
or U2518 (N_2518,N_2474,N_2420);
nor U2519 (N_2519,N_2400,N_2446);
nand U2520 (N_2520,N_2412,N_2421);
or U2521 (N_2521,N_2434,N_2438);
or U2522 (N_2522,N_2461,N_2413);
nand U2523 (N_2523,N_2452,N_2440);
and U2524 (N_2524,N_2445,N_2474);
xor U2525 (N_2525,N_2454,N_2406);
nor U2526 (N_2526,N_2423,N_2428);
or U2527 (N_2527,N_2464,N_2447);
xor U2528 (N_2528,N_2410,N_2435);
nor U2529 (N_2529,N_2411,N_2413);
nor U2530 (N_2530,N_2445,N_2410);
and U2531 (N_2531,N_2443,N_2474);
xor U2532 (N_2532,N_2426,N_2469);
or U2533 (N_2533,N_2406,N_2412);
nor U2534 (N_2534,N_2465,N_2453);
or U2535 (N_2535,N_2438,N_2442);
nand U2536 (N_2536,N_2460,N_2440);
nand U2537 (N_2537,N_2438,N_2473);
nand U2538 (N_2538,N_2409,N_2451);
nor U2539 (N_2539,N_2469,N_2425);
xnor U2540 (N_2540,N_2467,N_2422);
nand U2541 (N_2541,N_2473,N_2401);
and U2542 (N_2542,N_2435,N_2461);
nand U2543 (N_2543,N_2431,N_2418);
or U2544 (N_2544,N_2430,N_2433);
and U2545 (N_2545,N_2419,N_2429);
and U2546 (N_2546,N_2466,N_2443);
nand U2547 (N_2547,N_2415,N_2471);
nor U2548 (N_2548,N_2442,N_2409);
or U2549 (N_2549,N_2453,N_2407);
and U2550 (N_2550,N_2502,N_2527);
xnor U2551 (N_2551,N_2477,N_2530);
and U2552 (N_2552,N_2488,N_2478);
and U2553 (N_2553,N_2521,N_2543);
and U2554 (N_2554,N_2520,N_2494);
or U2555 (N_2555,N_2490,N_2500);
xnor U2556 (N_2556,N_2522,N_2508);
and U2557 (N_2557,N_2542,N_2546);
nand U2558 (N_2558,N_2504,N_2495);
and U2559 (N_2559,N_2525,N_2512);
or U2560 (N_2560,N_2485,N_2541);
nor U2561 (N_2561,N_2513,N_2532);
nor U2562 (N_2562,N_2540,N_2524);
and U2563 (N_2563,N_2515,N_2492);
nor U2564 (N_2564,N_2534,N_2538);
or U2565 (N_2565,N_2548,N_2511);
nor U2566 (N_2566,N_2505,N_2531);
xor U2567 (N_2567,N_2482,N_2487);
xnor U2568 (N_2568,N_2518,N_2483);
nand U2569 (N_2569,N_2498,N_2509);
nor U2570 (N_2570,N_2537,N_2529);
nor U2571 (N_2571,N_2503,N_2517);
and U2572 (N_2572,N_2536,N_2523);
and U2573 (N_2573,N_2549,N_2519);
or U2574 (N_2574,N_2499,N_2489);
and U2575 (N_2575,N_2496,N_2475);
and U2576 (N_2576,N_2486,N_2497);
xor U2577 (N_2577,N_2547,N_2476);
nor U2578 (N_2578,N_2507,N_2526);
and U2579 (N_2579,N_2479,N_2493);
and U2580 (N_2580,N_2544,N_2535);
or U2581 (N_2581,N_2484,N_2501);
or U2582 (N_2582,N_2528,N_2481);
or U2583 (N_2583,N_2506,N_2545);
and U2584 (N_2584,N_2539,N_2491);
xor U2585 (N_2585,N_2514,N_2516);
nor U2586 (N_2586,N_2510,N_2533);
xor U2587 (N_2587,N_2480,N_2487);
or U2588 (N_2588,N_2538,N_2476);
xnor U2589 (N_2589,N_2512,N_2538);
or U2590 (N_2590,N_2484,N_2522);
or U2591 (N_2591,N_2476,N_2537);
xor U2592 (N_2592,N_2526,N_2511);
nand U2593 (N_2593,N_2499,N_2515);
or U2594 (N_2594,N_2489,N_2530);
or U2595 (N_2595,N_2482,N_2526);
nor U2596 (N_2596,N_2500,N_2505);
or U2597 (N_2597,N_2490,N_2527);
and U2598 (N_2598,N_2540,N_2541);
xnor U2599 (N_2599,N_2498,N_2548);
or U2600 (N_2600,N_2486,N_2539);
nand U2601 (N_2601,N_2540,N_2520);
and U2602 (N_2602,N_2477,N_2544);
nand U2603 (N_2603,N_2510,N_2512);
and U2604 (N_2604,N_2536,N_2519);
nand U2605 (N_2605,N_2511,N_2494);
or U2606 (N_2606,N_2532,N_2494);
nand U2607 (N_2607,N_2490,N_2501);
and U2608 (N_2608,N_2539,N_2501);
nand U2609 (N_2609,N_2526,N_2537);
or U2610 (N_2610,N_2486,N_2546);
nand U2611 (N_2611,N_2542,N_2544);
nand U2612 (N_2612,N_2512,N_2496);
nand U2613 (N_2613,N_2508,N_2483);
or U2614 (N_2614,N_2545,N_2497);
nor U2615 (N_2615,N_2513,N_2515);
and U2616 (N_2616,N_2530,N_2490);
xor U2617 (N_2617,N_2520,N_2504);
nand U2618 (N_2618,N_2537,N_2518);
nand U2619 (N_2619,N_2482,N_2536);
and U2620 (N_2620,N_2515,N_2527);
nand U2621 (N_2621,N_2527,N_2482);
or U2622 (N_2622,N_2524,N_2537);
and U2623 (N_2623,N_2493,N_2514);
nand U2624 (N_2624,N_2484,N_2521);
or U2625 (N_2625,N_2600,N_2568);
xnor U2626 (N_2626,N_2599,N_2608);
or U2627 (N_2627,N_2578,N_2611);
and U2628 (N_2628,N_2587,N_2595);
nor U2629 (N_2629,N_2607,N_2584);
nor U2630 (N_2630,N_2603,N_2616);
nor U2631 (N_2631,N_2555,N_2550);
nand U2632 (N_2632,N_2570,N_2601);
nand U2633 (N_2633,N_2619,N_2604);
nor U2634 (N_2634,N_2623,N_2561);
or U2635 (N_2635,N_2614,N_2588);
nor U2636 (N_2636,N_2581,N_2559);
nand U2637 (N_2637,N_2572,N_2577);
and U2638 (N_2638,N_2609,N_2560);
or U2639 (N_2639,N_2593,N_2569);
and U2640 (N_2640,N_2602,N_2576);
and U2641 (N_2641,N_2566,N_2554);
nand U2642 (N_2642,N_2624,N_2563);
and U2643 (N_2643,N_2598,N_2567);
or U2644 (N_2644,N_2586,N_2589);
nand U2645 (N_2645,N_2610,N_2556);
nand U2646 (N_2646,N_2592,N_2596);
nand U2647 (N_2647,N_2612,N_2562);
xnor U2648 (N_2648,N_2594,N_2553);
nor U2649 (N_2649,N_2565,N_2597);
nor U2650 (N_2650,N_2574,N_2585);
nor U2651 (N_2651,N_2620,N_2605);
and U2652 (N_2652,N_2615,N_2571);
nand U2653 (N_2653,N_2580,N_2613);
nor U2654 (N_2654,N_2575,N_2583);
nand U2655 (N_2655,N_2622,N_2582);
nor U2656 (N_2656,N_2552,N_2618);
nor U2657 (N_2657,N_2591,N_2606);
xnor U2658 (N_2658,N_2557,N_2551);
and U2659 (N_2659,N_2564,N_2558);
and U2660 (N_2660,N_2621,N_2617);
or U2661 (N_2661,N_2590,N_2579);
nor U2662 (N_2662,N_2573,N_2557);
and U2663 (N_2663,N_2618,N_2554);
nor U2664 (N_2664,N_2596,N_2572);
nand U2665 (N_2665,N_2599,N_2601);
nand U2666 (N_2666,N_2612,N_2570);
and U2667 (N_2667,N_2566,N_2570);
and U2668 (N_2668,N_2600,N_2589);
nor U2669 (N_2669,N_2608,N_2593);
and U2670 (N_2670,N_2594,N_2566);
or U2671 (N_2671,N_2555,N_2598);
nor U2672 (N_2672,N_2593,N_2580);
and U2673 (N_2673,N_2620,N_2587);
nor U2674 (N_2674,N_2619,N_2595);
or U2675 (N_2675,N_2559,N_2605);
nor U2676 (N_2676,N_2596,N_2560);
and U2677 (N_2677,N_2561,N_2585);
or U2678 (N_2678,N_2593,N_2614);
and U2679 (N_2679,N_2598,N_2620);
or U2680 (N_2680,N_2591,N_2616);
and U2681 (N_2681,N_2618,N_2617);
and U2682 (N_2682,N_2623,N_2612);
and U2683 (N_2683,N_2592,N_2607);
or U2684 (N_2684,N_2551,N_2615);
xnor U2685 (N_2685,N_2551,N_2560);
and U2686 (N_2686,N_2612,N_2617);
nor U2687 (N_2687,N_2570,N_2583);
xor U2688 (N_2688,N_2571,N_2584);
nor U2689 (N_2689,N_2557,N_2622);
xor U2690 (N_2690,N_2624,N_2576);
and U2691 (N_2691,N_2614,N_2616);
xnor U2692 (N_2692,N_2563,N_2615);
or U2693 (N_2693,N_2611,N_2566);
nand U2694 (N_2694,N_2591,N_2570);
and U2695 (N_2695,N_2566,N_2562);
and U2696 (N_2696,N_2569,N_2615);
or U2697 (N_2697,N_2586,N_2560);
nand U2698 (N_2698,N_2555,N_2587);
and U2699 (N_2699,N_2608,N_2611);
nand U2700 (N_2700,N_2647,N_2695);
nor U2701 (N_2701,N_2666,N_2678);
or U2702 (N_2702,N_2649,N_2657);
nor U2703 (N_2703,N_2694,N_2697);
nor U2704 (N_2704,N_2665,N_2641);
and U2705 (N_2705,N_2662,N_2639);
nor U2706 (N_2706,N_2638,N_2683);
nor U2707 (N_2707,N_2632,N_2655);
and U2708 (N_2708,N_2661,N_2684);
nand U2709 (N_2709,N_2630,N_2698);
nand U2710 (N_2710,N_2672,N_2680);
nand U2711 (N_2711,N_2664,N_2692);
or U2712 (N_2712,N_2636,N_2675);
or U2713 (N_2713,N_2663,N_2681);
nand U2714 (N_2714,N_2643,N_2656);
and U2715 (N_2715,N_2627,N_2640);
nor U2716 (N_2716,N_2693,N_2644);
or U2717 (N_2717,N_2654,N_2634);
nand U2718 (N_2718,N_2648,N_2676);
nor U2719 (N_2719,N_2645,N_2690);
nand U2720 (N_2720,N_2699,N_2631);
nand U2721 (N_2721,N_2671,N_2646);
nand U2722 (N_2722,N_2625,N_2670);
or U2723 (N_2723,N_2653,N_2650);
nand U2724 (N_2724,N_2677,N_2685);
and U2725 (N_2725,N_2687,N_2682);
nand U2726 (N_2726,N_2691,N_2674);
or U2727 (N_2727,N_2673,N_2633);
and U2728 (N_2728,N_2629,N_2637);
or U2729 (N_2729,N_2688,N_2626);
nor U2730 (N_2730,N_2679,N_2668);
and U2731 (N_2731,N_2686,N_2658);
or U2732 (N_2732,N_2628,N_2660);
nor U2733 (N_2733,N_2652,N_2651);
nand U2734 (N_2734,N_2667,N_2642);
nand U2735 (N_2735,N_2689,N_2669);
nand U2736 (N_2736,N_2635,N_2659);
nor U2737 (N_2737,N_2696,N_2628);
or U2738 (N_2738,N_2674,N_2659);
xnor U2739 (N_2739,N_2688,N_2631);
nor U2740 (N_2740,N_2680,N_2645);
or U2741 (N_2741,N_2642,N_2645);
nor U2742 (N_2742,N_2650,N_2638);
nor U2743 (N_2743,N_2694,N_2638);
nor U2744 (N_2744,N_2687,N_2653);
or U2745 (N_2745,N_2672,N_2645);
and U2746 (N_2746,N_2628,N_2647);
nor U2747 (N_2747,N_2693,N_2660);
and U2748 (N_2748,N_2699,N_2638);
nand U2749 (N_2749,N_2690,N_2648);
nor U2750 (N_2750,N_2649,N_2673);
nor U2751 (N_2751,N_2649,N_2626);
and U2752 (N_2752,N_2673,N_2691);
and U2753 (N_2753,N_2675,N_2692);
xnor U2754 (N_2754,N_2671,N_2669);
nor U2755 (N_2755,N_2696,N_2656);
nand U2756 (N_2756,N_2652,N_2654);
xor U2757 (N_2757,N_2686,N_2677);
xnor U2758 (N_2758,N_2638,N_2630);
nor U2759 (N_2759,N_2678,N_2656);
nor U2760 (N_2760,N_2672,N_2635);
nor U2761 (N_2761,N_2670,N_2630);
or U2762 (N_2762,N_2634,N_2684);
nor U2763 (N_2763,N_2675,N_2689);
or U2764 (N_2764,N_2632,N_2646);
nor U2765 (N_2765,N_2635,N_2628);
and U2766 (N_2766,N_2637,N_2698);
and U2767 (N_2767,N_2671,N_2639);
or U2768 (N_2768,N_2650,N_2631);
nor U2769 (N_2769,N_2688,N_2690);
or U2770 (N_2770,N_2670,N_2689);
and U2771 (N_2771,N_2669,N_2655);
and U2772 (N_2772,N_2634,N_2635);
nor U2773 (N_2773,N_2675,N_2674);
and U2774 (N_2774,N_2633,N_2637);
nand U2775 (N_2775,N_2750,N_2748);
nand U2776 (N_2776,N_2742,N_2700);
xnor U2777 (N_2777,N_2724,N_2763);
and U2778 (N_2778,N_2768,N_2772);
nor U2779 (N_2779,N_2721,N_2729);
nand U2780 (N_2780,N_2752,N_2734);
nand U2781 (N_2781,N_2701,N_2757);
or U2782 (N_2782,N_2755,N_2764);
or U2783 (N_2783,N_2727,N_2759);
xnor U2784 (N_2784,N_2740,N_2716);
and U2785 (N_2785,N_2710,N_2719);
nor U2786 (N_2786,N_2723,N_2746);
nand U2787 (N_2787,N_2713,N_2725);
xnor U2788 (N_2788,N_2744,N_2743);
nand U2789 (N_2789,N_2753,N_2739);
or U2790 (N_2790,N_2704,N_2766);
xnor U2791 (N_2791,N_2761,N_2718);
nor U2792 (N_2792,N_2765,N_2745);
or U2793 (N_2793,N_2741,N_2703);
and U2794 (N_2794,N_2767,N_2774);
and U2795 (N_2795,N_2756,N_2712);
or U2796 (N_2796,N_2715,N_2747);
nand U2797 (N_2797,N_2708,N_2762);
nand U2798 (N_2798,N_2730,N_2737);
nor U2799 (N_2799,N_2769,N_2702);
and U2800 (N_2800,N_2733,N_2770);
nand U2801 (N_2801,N_2760,N_2705);
and U2802 (N_2802,N_2726,N_2735);
and U2803 (N_2803,N_2717,N_2706);
and U2804 (N_2804,N_2738,N_2758);
or U2805 (N_2805,N_2714,N_2732);
nor U2806 (N_2806,N_2707,N_2736);
nor U2807 (N_2807,N_2751,N_2773);
and U2808 (N_2808,N_2754,N_2720);
and U2809 (N_2809,N_2728,N_2731);
xnor U2810 (N_2810,N_2749,N_2709);
nor U2811 (N_2811,N_2711,N_2722);
nand U2812 (N_2812,N_2771,N_2766);
nor U2813 (N_2813,N_2702,N_2746);
nor U2814 (N_2814,N_2714,N_2763);
nand U2815 (N_2815,N_2732,N_2771);
or U2816 (N_2816,N_2769,N_2728);
nand U2817 (N_2817,N_2740,N_2764);
xor U2818 (N_2818,N_2737,N_2722);
or U2819 (N_2819,N_2725,N_2768);
and U2820 (N_2820,N_2715,N_2701);
nand U2821 (N_2821,N_2743,N_2724);
or U2822 (N_2822,N_2737,N_2761);
xnor U2823 (N_2823,N_2717,N_2700);
nand U2824 (N_2824,N_2758,N_2746);
or U2825 (N_2825,N_2762,N_2767);
nor U2826 (N_2826,N_2709,N_2759);
nand U2827 (N_2827,N_2763,N_2756);
nor U2828 (N_2828,N_2739,N_2705);
nor U2829 (N_2829,N_2755,N_2753);
or U2830 (N_2830,N_2765,N_2730);
or U2831 (N_2831,N_2765,N_2735);
and U2832 (N_2832,N_2728,N_2713);
xnor U2833 (N_2833,N_2741,N_2767);
nor U2834 (N_2834,N_2748,N_2753);
xor U2835 (N_2835,N_2760,N_2709);
nor U2836 (N_2836,N_2710,N_2707);
nor U2837 (N_2837,N_2730,N_2768);
nand U2838 (N_2838,N_2717,N_2727);
or U2839 (N_2839,N_2714,N_2760);
nor U2840 (N_2840,N_2711,N_2719);
nand U2841 (N_2841,N_2771,N_2700);
or U2842 (N_2842,N_2726,N_2737);
or U2843 (N_2843,N_2759,N_2752);
nor U2844 (N_2844,N_2761,N_2706);
and U2845 (N_2845,N_2758,N_2743);
nand U2846 (N_2846,N_2714,N_2704);
nand U2847 (N_2847,N_2736,N_2730);
and U2848 (N_2848,N_2773,N_2770);
or U2849 (N_2849,N_2769,N_2735);
or U2850 (N_2850,N_2825,N_2847);
and U2851 (N_2851,N_2790,N_2776);
nand U2852 (N_2852,N_2791,N_2814);
and U2853 (N_2853,N_2834,N_2832);
or U2854 (N_2854,N_2837,N_2812);
xor U2855 (N_2855,N_2793,N_2817);
xnor U2856 (N_2856,N_2818,N_2795);
nand U2857 (N_2857,N_2836,N_2798);
nand U2858 (N_2858,N_2816,N_2811);
nand U2859 (N_2859,N_2796,N_2806);
and U2860 (N_2860,N_2820,N_2801);
nand U2861 (N_2861,N_2815,N_2823);
and U2862 (N_2862,N_2848,N_2786);
nand U2863 (N_2863,N_2810,N_2829);
nor U2864 (N_2864,N_2808,N_2822);
and U2865 (N_2865,N_2846,N_2794);
nand U2866 (N_2866,N_2835,N_2777);
nor U2867 (N_2867,N_2805,N_2804);
nor U2868 (N_2868,N_2803,N_2792);
nor U2869 (N_2869,N_2783,N_2824);
nand U2870 (N_2870,N_2826,N_2841);
and U2871 (N_2871,N_2785,N_2845);
nand U2872 (N_2872,N_2800,N_2797);
xnor U2873 (N_2873,N_2839,N_2802);
nor U2874 (N_2874,N_2781,N_2840);
or U2875 (N_2875,N_2844,N_2821);
nor U2876 (N_2876,N_2779,N_2828);
or U2877 (N_2877,N_2838,N_2827);
and U2878 (N_2878,N_2849,N_2775);
xnor U2879 (N_2879,N_2782,N_2830);
or U2880 (N_2880,N_2788,N_2809);
nor U2881 (N_2881,N_2819,N_2807);
xnor U2882 (N_2882,N_2780,N_2833);
nand U2883 (N_2883,N_2799,N_2789);
and U2884 (N_2884,N_2778,N_2842);
or U2885 (N_2885,N_2843,N_2813);
nor U2886 (N_2886,N_2784,N_2787);
nand U2887 (N_2887,N_2831,N_2778);
and U2888 (N_2888,N_2795,N_2784);
xnor U2889 (N_2889,N_2814,N_2830);
or U2890 (N_2890,N_2775,N_2802);
nand U2891 (N_2891,N_2818,N_2830);
or U2892 (N_2892,N_2829,N_2830);
nor U2893 (N_2893,N_2814,N_2781);
nand U2894 (N_2894,N_2821,N_2843);
or U2895 (N_2895,N_2846,N_2822);
nand U2896 (N_2896,N_2810,N_2826);
or U2897 (N_2897,N_2793,N_2845);
or U2898 (N_2898,N_2787,N_2804);
nor U2899 (N_2899,N_2778,N_2836);
and U2900 (N_2900,N_2813,N_2808);
xor U2901 (N_2901,N_2825,N_2839);
or U2902 (N_2902,N_2797,N_2798);
nor U2903 (N_2903,N_2801,N_2786);
xor U2904 (N_2904,N_2783,N_2782);
or U2905 (N_2905,N_2823,N_2797);
nand U2906 (N_2906,N_2843,N_2785);
and U2907 (N_2907,N_2821,N_2792);
nor U2908 (N_2908,N_2776,N_2819);
nor U2909 (N_2909,N_2792,N_2784);
nand U2910 (N_2910,N_2839,N_2791);
and U2911 (N_2911,N_2786,N_2785);
or U2912 (N_2912,N_2842,N_2817);
nor U2913 (N_2913,N_2780,N_2785);
or U2914 (N_2914,N_2783,N_2800);
xor U2915 (N_2915,N_2799,N_2783);
or U2916 (N_2916,N_2844,N_2796);
and U2917 (N_2917,N_2778,N_2815);
nor U2918 (N_2918,N_2831,N_2797);
and U2919 (N_2919,N_2827,N_2793);
and U2920 (N_2920,N_2784,N_2798);
nor U2921 (N_2921,N_2786,N_2793);
nand U2922 (N_2922,N_2829,N_2846);
nor U2923 (N_2923,N_2824,N_2790);
nor U2924 (N_2924,N_2816,N_2795);
or U2925 (N_2925,N_2875,N_2868);
or U2926 (N_2926,N_2900,N_2889);
nor U2927 (N_2927,N_2879,N_2865);
or U2928 (N_2928,N_2901,N_2924);
nor U2929 (N_2929,N_2867,N_2921);
or U2930 (N_2930,N_2859,N_2919);
or U2931 (N_2931,N_2886,N_2861);
or U2932 (N_2932,N_2896,N_2855);
nand U2933 (N_2933,N_2862,N_2856);
nand U2934 (N_2934,N_2918,N_2878);
nand U2935 (N_2935,N_2897,N_2884);
nor U2936 (N_2936,N_2908,N_2905);
or U2937 (N_2937,N_2866,N_2903);
and U2938 (N_2938,N_2910,N_2888);
nor U2939 (N_2939,N_2850,N_2871);
or U2940 (N_2940,N_2858,N_2857);
and U2941 (N_2941,N_2920,N_2887);
nor U2942 (N_2942,N_2869,N_2902);
nor U2943 (N_2943,N_2882,N_2874);
or U2944 (N_2944,N_2881,N_2851);
nand U2945 (N_2945,N_2890,N_2907);
xor U2946 (N_2946,N_2863,N_2877);
xor U2947 (N_2947,N_2894,N_2912);
and U2948 (N_2948,N_2909,N_2898);
nand U2949 (N_2949,N_2899,N_2883);
nand U2950 (N_2950,N_2891,N_2904);
xnor U2951 (N_2951,N_2892,N_2852);
nor U2952 (N_2952,N_2911,N_2876);
nand U2953 (N_2953,N_2915,N_2893);
or U2954 (N_2954,N_2922,N_2885);
and U2955 (N_2955,N_2870,N_2923);
nand U2956 (N_2956,N_2906,N_2895);
nand U2957 (N_2957,N_2880,N_2872);
nor U2958 (N_2958,N_2860,N_2917);
and U2959 (N_2959,N_2873,N_2854);
nand U2960 (N_2960,N_2913,N_2916);
and U2961 (N_2961,N_2914,N_2853);
nor U2962 (N_2962,N_2864,N_2877);
or U2963 (N_2963,N_2924,N_2917);
and U2964 (N_2964,N_2909,N_2907);
or U2965 (N_2965,N_2890,N_2862);
nor U2966 (N_2966,N_2888,N_2893);
xor U2967 (N_2967,N_2886,N_2866);
nor U2968 (N_2968,N_2855,N_2892);
or U2969 (N_2969,N_2886,N_2888);
nand U2970 (N_2970,N_2906,N_2864);
and U2971 (N_2971,N_2865,N_2855);
or U2972 (N_2972,N_2882,N_2910);
or U2973 (N_2973,N_2914,N_2885);
nor U2974 (N_2974,N_2858,N_2868);
or U2975 (N_2975,N_2909,N_2905);
or U2976 (N_2976,N_2915,N_2865);
xnor U2977 (N_2977,N_2918,N_2862);
nand U2978 (N_2978,N_2888,N_2878);
or U2979 (N_2979,N_2855,N_2918);
and U2980 (N_2980,N_2881,N_2910);
nor U2981 (N_2981,N_2906,N_2851);
and U2982 (N_2982,N_2881,N_2852);
and U2983 (N_2983,N_2871,N_2906);
or U2984 (N_2984,N_2908,N_2861);
nand U2985 (N_2985,N_2878,N_2850);
or U2986 (N_2986,N_2873,N_2871);
nand U2987 (N_2987,N_2885,N_2862);
or U2988 (N_2988,N_2861,N_2890);
nor U2989 (N_2989,N_2867,N_2875);
nand U2990 (N_2990,N_2880,N_2913);
nor U2991 (N_2991,N_2903,N_2913);
and U2992 (N_2992,N_2867,N_2882);
and U2993 (N_2993,N_2910,N_2859);
nand U2994 (N_2994,N_2867,N_2865);
and U2995 (N_2995,N_2850,N_2865);
or U2996 (N_2996,N_2915,N_2884);
and U2997 (N_2997,N_2870,N_2861);
and U2998 (N_2998,N_2853,N_2886);
and U2999 (N_2999,N_2885,N_2852);
nor UO_0 (O_0,N_2969,N_2934);
nand UO_1 (O_1,N_2988,N_2997);
xor UO_2 (O_2,N_2970,N_2957);
nand UO_3 (O_3,N_2942,N_2925);
nand UO_4 (O_4,N_2978,N_2975);
or UO_5 (O_5,N_2939,N_2982);
or UO_6 (O_6,N_2960,N_2929);
xor UO_7 (O_7,N_2987,N_2961);
or UO_8 (O_8,N_2967,N_2945);
or UO_9 (O_9,N_2986,N_2973);
or UO_10 (O_10,N_2938,N_2956);
xnor UO_11 (O_11,N_2971,N_2936);
nand UO_12 (O_12,N_2963,N_2980);
or UO_13 (O_13,N_2994,N_2955);
nor UO_14 (O_14,N_2993,N_2996);
or UO_15 (O_15,N_2947,N_2984);
or UO_16 (O_16,N_2990,N_2941);
or UO_17 (O_17,N_2979,N_2946);
nor UO_18 (O_18,N_2930,N_2940);
or UO_19 (O_19,N_2974,N_2972);
nor UO_20 (O_20,N_2926,N_2943);
nor UO_21 (O_21,N_2981,N_2995);
nor UO_22 (O_22,N_2966,N_2935);
nand UO_23 (O_23,N_2983,N_2999);
or UO_24 (O_24,N_2948,N_2944);
or UO_25 (O_25,N_2954,N_2992);
and UO_26 (O_26,N_2931,N_2965);
and UO_27 (O_27,N_2958,N_2950);
nand UO_28 (O_28,N_2953,N_2959);
xnor UO_29 (O_29,N_2952,N_2977);
nor UO_30 (O_30,N_2968,N_2976);
and UO_31 (O_31,N_2937,N_2998);
xnor UO_32 (O_32,N_2962,N_2927);
or UO_33 (O_33,N_2951,N_2932);
nor UO_34 (O_34,N_2949,N_2985);
nand UO_35 (O_35,N_2933,N_2928);
nor UO_36 (O_36,N_2991,N_2989);
and UO_37 (O_37,N_2964,N_2931);
or UO_38 (O_38,N_2958,N_2938);
or UO_39 (O_39,N_2960,N_2967);
nor UO_40 (O_40,N_2966,N_2941);
and UO_41 (O_41,N_2967,N_2974);
nand UO_42 (O_42,N_2956,N_2986);
or UO_43 (O_43,N_2928,N_2952);
or UO_44 (O_44,N_2951,N_2990);
or UO_45 (O_45,N_2997,N_2994);
nor UO_46 (O_46,N_2960,N_2980);
nand UO_47 (O_47,N_2929,N_2966);
and UO_48 (O_48,N_2949,N_2981);
nor UO_49 (O_49,N_2960,N_2985);
nor UO_50 (O_50,N_2982,N_2966);
xnor UO_51 (O_51,N_2996,N_2936);
and UO_52 (O_52,N_2969,N_2972);
and UO_53 (O_53,N_2930,N_2982);
or UO_54 (O_54,N_2964,N_2982);
nand UO_55 (O_55,N_2985,N_2988);
and UO_56 (O_56,N_2993,N_2990);
or UO_57 (O_57,N_2998,N_2952);
or UO_58 (O_58,N_2959,N_2962);
nand UO_59 (O_59,N_2984,N_2982);
nand UO_60 (O_60,N_2960,N_2999);
and UO_61 (O_61,N_2970,N_2986);
nor UO_62 (O_62,N_2970,N_2998);
or UO_63 (O_63,N_2940,N_2976);
nand UO_64 (O_64,N_2936,N_2945);
and UO_65 (O_65,N_2969,N_2971);
nor UO_66 (O_66,N_2938,N_2934);
nand UO_67 (O_67,N_2938,N_2970);
and UO_68 (O_68,N_2929,N_2931);
nor UO_69 (O_69,N_2951,N_2976);
nor UO_70 (O_70,N_2992,N_2931);
and UO_71 (O_71,N_2963,N_2931);
xor UO_72 (O_72,N_2930,N_2949);
and UO_73 (O_73,N_2931,N_2981);
nor UO_74 (O_74,N_2937,N_2969);
or UO_75 (O_75,N_2967,N_2938);
nor UO_76 (O_76,N_2966,N_2990);
nor UO_77 (O_77,N_2934,N_2968);
xnor UO_78 (O_78,N_2985,N_2945);
and UO_79 (O_79,N_2990,N_2976);
or UO_80 (O_80,N_2949,N_2934);
nand UO_81 (O_81,N_2964,N_2972);
or UO_82 (O_82,N_2948,N_2981);
nand UO_83 (O_83,N_2937,N_2982);
nor UO_84 (O_84,N_2967,N_2951);
nor UO_85 (O_85,N_2925,N_2965);
nor UO_86 (O_86,N_2932,N_2967);
and UO_87 (O_87,N_2931,N_2982);
xor UO_88 (O_88,N_2956,N_2958);
nor UO_89 (O_89,N_2950,N_2944);
nor UO_90 (O_90,N_2925,N_2986);
nor UO_91 (O_91,N_2997,N_2986);
or UO_92 (O_92,N_2985,N_2986);
nand UO_93 (O_93,N_2928,N_2959);
and UO_94 (O_94,N_2932,N_2988);
nor UO_95 (O_95,N_2961,N_2933);
nand UO_96 (O_96,N_2956,N_2979);
and UO_97 (O_97,N_2951,N_2991);
nor UO_98 (O_98,N_2993,N_2937);
nor UO_99 (O_99,N_2950,N_2947);
or UO_100 (O_100,N_2947,N_2981);
nand UO_101 (O_101,N_2992,N_2978);
and UO_102 (O_102,N_2998,N_2966);
and UO_103 (O_103,N_2976,N_2994);
and UO_104 (O_104,N_2928,N_2993);
nand UO_105 (O_105,N_2948,N_2958);
and UO_106 (O_106,N_2945,N_2949);
and UO_107 (O_107,N_2962,N_2992);
nor UO_108 (O_108,N_2970,N_2988);
nor UO_109 (O_109,N_2986,N_2942);
xnor UO_110 (O_110,N_2926,N_2925);
nand UO_111 (O_111,N_2965,N_2996);
and UO_112 (O_112,N_2968,N_2971);
or UO_113 (O_113,N_2955,N_2971);
nand UO_114 (O_114,N_2987,N_2968);
and UO_115 (O_115,N_2946,N_2966);
or UO_116 (O_116,N_2928,N_2989);
nor UO_117 (O_117,N_2980,N_2932);
or UO_118 (O_118,N_2949,N_2975);
xor UO_119 (O_119,N_2926,N_2969);
or UO_120 (O_120,N_2992,N_2930);
nand UO_121 (O_121,N_2995,N_2931);
nand UO_122 (O_122,N_2972,N_2999);
or UO_123 (O_123,N_2953,N_2937);
and UO_124 (O_124,N_2947,N_2940);
nor UO_125 (O_125,N_2936,N_2955);
or UO_126 (O_126,N_2925,N_2947);
and UO_127 (O_127,N_2954,N_2925);
nor UO_128 (O_128,N_2944,N_2956);
or UO_129 (O_129,N_2927,N_2998);
or UO_130 (O_130,N_2938,N_2973);
and UO_131 (O_131,N_2970,N_2979);
xor UO_132 (O_132,N_2940,N_2954);
xor UO_133 (O_133,N_2978,N_2948);
or UO_134 (O_134,N_2970,N_2927);
or UO_135 (O_135,N_2957,N_2963);
nand UO_136 (O_136,N_2986,N_2933);
or UO_137 (O_137,N_2950,N_2936);
and UO_138 (O_138,N_2966,N_2962);
nand UO_139 (O_139,N_2935,N_2958);
or UO_140 (O_140,N_2937,N_2951);
nor UO_141 (O_141,N_2994,N_2938);
and UO_142 (O_142,N_2973,N_2992);
or UO_143 (O_143,N_2951,N_2952);
xnor UO_144 (O_144,N_2997,N_2926);
nor UO_145 (O_145,N_2944,N_2994);
and UO_146 (O_146,N_2995,N_2945);
or UO_147 (O_147,N_2925,N_2997);
or UO_148 (O_148,N_2964,N_2944);
nor UO_149 (O_149,N_2958,N_2975);
or UO_150 (O_150,N_2988,N_2956);
and UO_151 (O_151,N_2959,N_2990);
and UO_152 (O_152,N_2957,N_2962);
and UO_153 (O_153,N_2968,N_2931);
xnor UO_154 (O_154,N_2997,N_2950);
nor UO_155 (O_155,N_2982,N_2991);
or UO_156 (O_156,N_2986,N_2979);
xnor UO_157 (O_157,N_2948,N_2970);
or UO_158 (O_158,N_2986,N_2949);
nand UO_159 (O_159,N_2944,N_2925);
xor UO_160 (O_160,N_2926,N_2993);
and UO_161 (O_161,N_2980,N_2979);
nand UO_162 (O_162,N_2998,N_2925);
and UO_163 (O_163,N_2969,N_2941);
nor UO_164 (O_164,N_2957,N_2932);
and UO_165 (O_165,N_2964,N_2975);
and UO_166 (O_166,N_2987,N_2954);
nand UO_167 (O_167,N_2943,N_2959);
nor UO_168 (O_168,N_2979,N_2939);
and UO_169 (O_169,N_2980,N_2983);
and UO_170 (O_170,N_2990,N_2942);
xor UO_171 (O_171,N_2952,N_2993);
nand UO_172 (O_172,N_2997,N_2965);
nand UO_173 (O_173,N_2994,N_2927);
nand UO_174 (O_174,N_2997,N_2970);
or UO_175 (O_175,N_2974,N_2994);
nor UO_176 (O_176,N_2954,N_2999);
nor UO_177 (O_177,N_2945,N_2933);
and UO_178 (O_178,N_2956,N_2950);
or UO_179 (O_179,N_2969,N_2957);
and UO_180 (O_180,N_2956,N_2987);
and UO_181 (O_181,N_2931,N_2955);
and UO_182 (O_182,N_2963,N_2997);
or UO_183 (O_183,N_2965,N_2951);
and UO_184 (O_184,N_2974,N_2953);
or UO_185 (O_185,N_2947,N_2993);
nor UO_186 (O_186,N_2968,N_2975);
nand UO_187 (O_187,N_2957,N_2927);
nor UO_188 (O_188,N_2988,N_2946);
nor UO_189 (O_189,N_2984,N_2983);
or UO_190 (O_190,N_2943,N_2945);
nand UO_191 (O_191,N_2930,N_2934);
and UO_192 (O_192,N_2964,N_2984);
nor UO_193 (O_193,N_2958,N_2992);
or UO_194 (O_194,N_2931,N_2938);
nand UO_195 (O_195,N_2939,N_2998);
or UO_196 (O_196,N_2934,N_2983);
nor UO_197 (O_197,N_2947,N_2988);
or UO_198 (O_198,N_2949,N_2997);
and UO_199 (O_199,N_2941,N_2991);
nor UO_200 (O_200,N_2964,N_2978);
nand UO_201 (O_201,N_2929,N_2972);
and UO_202 (O_202,N_2945,N_2932);
nand UO_203 (O_203,N_2950,N_2926);
nand UO_204 (O_204,N_2974,N_2980);
nand UO_205 (O_205,N_2945,N_2962);
or UO_206 (O_206,N_2993,N_2992);
xnor UO_207 (O_207,N_2992,N_2939);
or UO_208 (O_208,N_2943,N_2996);
xnor UO_209 (O_209,N_2978,N_2958);
nor UO_210 (O_210,N_2956,N_2984);
nand UO_211 (O_211,N_2980,N_2981);
nand UO_212 (O_212,N_2962,N_2953);
or UO_213 (O_213,N_2995,N_2956);
or UO_214 (O_214,N_2982,N_2935);
and UO_215 (O_215,N_2963,N_2967);
and UO_216 (O_216,N_2992,N_2934);
nor UO_217 (O_217,N_2999,N_2992);
nor UO_218 (O_218,N_2970,N_2960);
nor UO_219 (O_219,N_2977,N_2989);
nor UO_220 (O_220,N_2983,N_2979);
or UO_221 (O_221,N_2996,N_2977);
nor UO_222 (O_222,N_2974,N_2942);
nand UO_223 (O_223,N_2980,N_2948);
and UO_224 (O_224,N_2932,N_2955);
or UO_225 (O_225,N_2955,N_2973);
or UO_226 (O_226,N_2977,N_2925);
and UO_227 (O_227,N_2943,N_2971);
nand UO_228 (O_228,N_2955,N_2949);
nor UO_229 (O_229,N_2933,N_2925);
nand UO_230 (O_230,N_2983,N_2932);
nor UO_231 (O_231,N_2968,N_2933);
nand UO_232 (O_232,N_2998,N_2938);
nor UO_233 (O_233,N_2990,N_2984);
and UO_234 (O_234,N_2993,N_2934);
or UO_235 (O_235,N_2977,N_2981);
and UO_236 (O_236,N_2929,N_2938);
or UO_237 (O_237,N_2994,N_2936);
xnor UO_238 (O_238,N_2972,N_2939);
nand UO_239 (O_239,N_2944,N_2933);
xor UO_240 (O_240,N_2950,N_2977);
or UO_241 (O_241,N_2929,N_2940);
or UO_242 (O_242,N_2962,N_2958);
xnor UO_243 (O_243,N_2926,N_2937);
nand UO_244 (O_244,N_2932,N_2943);
nor UO_245 (O_245,N_2947,N_2983);
nand UO_246 (O_246,N_2989,N_2933);
xnor UO_247 (O_247,N_2985,N_2983);
or UO_248 (O_248,N_2982,N_2956);
and UO_249 (O_249,N_2942,N_2928);
or UO_250 (O_250,N_2934,N_2962);
nor UO_251 (O_251,N_2994,N_2958);
nor UO_252 (O_252,N_2935,N_2937);
or UO_253 (O_253,N_2960,N_2975);
xor UO_254 (O_254,N_2999,N_2974);
and UO_255 (O_255,N_2985,N_2978);
xnor UO_256 (O_256,N_2948,N_2952);
or UO_257 (O_257,N_2960,N_2938);
or UO_258 (O_258,N_2936,N_2970);
xor UO_259 (O_259,N_2962,N_2967);
or UO_260 (O_260,N_2982,N_2977);
nand UO_261 (O_261,N_2966,N_2948);
or UO_262 (O_262,N_2932,N_2935);
nand UO_263 (O_263,N_2964,N_2949);
nor UO_264 (O_264,N_2959,N_2946);
nor UO_265 (O_265,N_2955,N_2975);
and UO_266 (O_266,N_2958,N_2933);
and UO_267 (O_267,N_2933,N_2969);
and UO_268 (O_268,N_2957,N_2964);
nor UO_269 (O_269,N_2985,N_2968);
nor UO_270 (O_270,N_2942,N_2952);
and UO_271 (O_271,N_2985,N_2926);
or UO_272 (O_272,N_2950,N_2954);
nor UO_273 (O_273,N_2987,N_2959);
nand UO_274 (O_274,N_2926,N_2994);
nand UO_275 (O_275,N_2971,N_2967);
and UO_276 (O_276,N_2938,N_2926);
or UO_277 (O_277,N_2999,N_2950);
nor UO_278 (O_278,N_2980,N_2947);
nand UO_279 (O_279,N_2968,N_2990);
nand UO_280 (O_280,N_2953,N_2965);
or UO_281 (O_281,N_2967,N_2980);
nor UO_282 (O_282,N_2946,N_2934);
nand UO_283 (O_283,N_2981,N_2930);
nand UO_284 (O_284,N_2954,N_2930);
nand UO_285 (O_285,N_2929,N_2934);
or UO_286 (O_286,N_2988,N_2987);
and UO_287 (O_287,N_2978,N_2938);
and UO_288 (O_288,N_2988,N_2929);
nand UO_289 (O_289,N_2925,N_2940);
and UO_290 (O_290,N_2972,N_2976);
and UO_291 (O_291,N_2965,N_2949);
or UO_292 (O_292,N_2970,N_2993);
nand UO_293 (O_293,N_2967,N_2925);
and UO_294 (O_294,N_2961,N_2966);
and UO_295 (O_295,N_2994,N_2967);
and UO_296 (O_296,N_2939,N_2965);
or UO_297 (O_297,N_2996,N_2963);
nor UO_298 (O_298,N_2928,N_2991);
or UO_299 (O_299,N_2966,N_2996);
nand UO_300 (O_300,N_2950,N_2935);
nor UO_301 (O_301,N_2938,N_2939);
nand UO_302 (O_302,N_2994,N_2999);
and UO_303 (O_303,N_2957,N_2954);
xor UO_304 (O_304,N_2928,N_2999);
or UO_305 (O_305,N_2972,N_2959);
nor UO_306 (O_306,N_2945,N_2968);
xor UO_307 (O_307,N_2977,N_2972);
nand UO_308 (O_308,N_2980,N_2968);
or UO_309 (O_309,N_2994,N_2986);
or UO_310 (O_310,N_2968,N_2925);
and UO_311 (O_311,N_2997,N_2983);
or UO_312 (O_312,N_2935,N_2925);
nand UO_313 (O_313,N_2937,N_2956);
nand UO_314 (O_314,N_2942,N_2936);
xnor UO_315 (O_315,N_2954,N_2972);
or UO_316 (O_316,N_2929,N_2990);
nand UO_317 (O_317,N_2971,N_2944);
or UO_318 (O_318,N_2926,N_2955);
nand UO_319 (O_319,N_2970,N_2974);
nor UO_320 (O_320,N_2951,N_2964);
nor UO_321 (O_321,N_2932,N_2997);
xnor UO_322 (O_322,N_2978,N_2926);
xnor UO_323 (O_323,N_2966,N_2944);
and UO_324 (O_324,N_2977,N_2995);
or UO_325 (O_325,N_2956,N_2930);
and UO_326 (O_326,N_2961,N_2951);
nand UO_327 (O_327,N_2941,N_2949);
and UO_328 (O_328,N_2939,N_2945);
nor UO_329 (O_329,N_2979,N_2982);
nor UO_330 (O_330,N_2939,N_2980);
and UO_331 (O_331,N_2947,N_2971);
nand UO_332 (O_332,N_2941,N_2937);
xor UO_333 (O_333,N_2984,N_2930);
nor UO_334 (O_334,N_2932,N_2954);
and UO_335 (O_335,N_2943,N_2942);
or UO_336 (O_336,N_2988,N_2953);
nand UO_337 (O_337,N_2975,N_2944);
xor UO_338 (O_338,N_2926,N_2942);
nand UO_339 (O_339,N_2954,N_2933);
xnor UO_340 (O_340,N_2984,N_2962);
nand UO_341 (O_341,N_2942,N_2950);
nand UO_342 (O_342,N_2965,N_2988);
and UO_343 (O_343,N_2927,N_2932);
xor UO_344 (O_344,N_2967,N_2996);
nand UO_345 (O_345,N_2963,N_2984);
xnor UO_346 (O_346,N_2972,N_2991);
xor UO_347 (O_347,N_2944,N_2983);
and UO_348 (O_348,N_2991,N_2957);
nor UO_349 (O_349,N_2977,N_2956);
nor UO_350 (O_350,N_2981,N_2976);
nand UO_351 (O_351,N_2927,N_2984);
nand UO_352 (O_352,N_2954,N_2976);
and UO_353 (O_353,N_2998,N_2929);
nor UO_354 (O_354,N_2989,N_2942);
and UO_355 (O_355,N_2997,N_2991);
xnor UO_356 (O_356,N_2977,N_2944);
and UO_357 (O_357,N_2976,N_2998);
nor UO_358 (O_358,N_2931,N_2962);
and UO_359 (O_359,N_2963,N_2932);
and UO_360 (O_360,N_2940,N_2972);
nor UO_361 (O_361,N_2936,N_2986);
or UO_362 (O_362,N_2959,N_2929);
or UO_363 (O_363,N_2936,N_2982);
nor UO_364 (O_364,N_2939,N_2936);
and UO_365 (O_365,N_2926,N_2980);
and UO_366 (O_366,N_2999,N_2959);
and UO_367 (O_367,N_2946,N_2991);
or UO_368 (O_368,N_2949,N_2976);
or UO_369 (O_369,N_2987,N_2986);
or UO_370 (O_370,N_2989,N_2992);
or UO_371 (O_371,N_2978,N_2986);
and UO_372 (O_372,N_2977,N_2949);
and UO_373 (O_373,N_2935,N_2968);
nand UO_374 (O_374,N_2965,N_2935);
and UO_375 (O_375,N_2954,N_2998);
nor UO_376 (O_376,N_2947,N_2977);
nand UO_377 (O_377,N_2968,N_2955);
xor UO_378 (O_378,N_2976,N_2993);
nand UO_379 (O_379,N_2991,N_2993);
nor UO_380 (O_380,N_2946,N_2944);
nand UO_381 (O_381,N_2997,N_2960);
and UO_382 (O_382,N_2947,N_2938);
xnor UO_383 (O_383,N_2948,N_2999);
nand UO_384 (O_384,N_2940,N_2983);
xnor UO_385 (O_385,N_2973,N_2993);
nor UO_386 (O_386,N_2985,N_2959);
xor UO_387 (O_387,N_2937,N_2947);
and UO_388 (O_388,N_2994,N_2946);
and UO_389 (O_389,N_2967,N_2987);
nand UO_390 (O_390,N_2941,N_2945);
nor UO_391 (O_391,N_2996,N_2952);
or UO_392 (O_392,N_2933,N_2972);
nand UO_393 (O_393,N_2985,N_2938);
or UO_394 (O_394,N_2941,N_2993);
or UO_395 (O_395,N_2987,N_2936);
xnor UO_396 (O_396,N_2964,N_2952);
and UO_397 (O_397,N_2990,N_2973);
nand UO_398 (O_398,N_2925,N_2985);
nand UO_399 (O_399,N_2957,N_2986);
or UO_400 (O_400,N_2945,N_2975);
and UO_401 (O_401,N_2937,N_2946);
or UO_402 (O_402,N_2941,N_2952);
or UO_403 (O_403,N_2943,N_2972);
nor UO_404 (O_404,N_2947,N_2929);
nand UO_405 (O_405,N_2933,N_2975);
nand UO_406 (O_406,N_2941,N_2979);
nand UO_407 (O_407,N_2982,N_2961);
and UO_408 (O_408,N_2926,N_2968);
nand UO_409 (O_409,N_2983,N_2969);
nand UO_410 (O_410,N_2987,N_2980);
or UO_411 (O_411,N_2938,N_2935);
xor UO_412 (O_412,N_2925,N_2956);
xor UO_413 (O_413,N_2965,N_2967);
xor UO_414 (O_414,N_2956,N_2967);
or UO_415 (O_415,N_2961,N_2958);
nor UO_416 (O_416,N_2948,N_2976);
nand UO_417 (O_417,N_2940,N_2969);
nor UO_418 (O_418,N_2991,N_2956);
nor UO_419 (O_419,N_2931,N_2941);
or UO_420 (O_420,N_2928,N_2980);
and UO_421 (O_421,N_2968,N_2948);
and UO_422 (O_422,N_2967,N_2931);
and UO_423 (O_423,N_2963,N_2977);
and UO_424 (O_424,N_2995,N_2940);
nand UO_425 (O_425,N_2932,N_2986);
nand UO_426 (O_426,N_2958,N_2993);
or UO_427 (O_427,N_2977,N_2941);
or UO_428 (O_428,N_2959,N_2971);
or UO_429 (O_429,N_2978,N_2984);
nor UO_430 (O_430,N_2941,N_2978);
nor UO_431 (O_431,N_2978,N_2965);
and UO_432 (O_432,N_2935,N_2990);
or UO_433 (O_433,N_2970,N_2994);
and UO_434 (O_434,N_2931,N_2926);
or UO_435 (O_435,N_2933,N_2936);
nor UO_436 (O_436,N_2967,N_2958);
or UO_437 (O_437,N_2970,N_2949);
nor UO_438 (O_438,N_2940,N_2982);
nor UO_439 (O_439,N_2997,N_2982);
and UO_440 (O_440,N_2993,N_2983);
nor UO_441 (O_441,N_2968,N_2998);
or UO_442 (O_442,N_2992,N_2983);
nand UO_443 (O_443,N_2952,N_2962);
nor UO_444 (O_444,N_2941,N_2942);
nor UO_445 (O_445,N_2966,N_2936);
nand UO_446 (O_446,N_2944,N_2974);
or UO_447 (O_447,N_2961,N_2931);
or UO_448 (O_448,N_2933,N_2943);
and UO_449 (O_449,N_2963,N_2969);
or UO_450 (O_450,N_2927,N_2947);
or UO_451 (O_451,N_2929,N_2930);
or UO_452 (O_452,N_2986,N_2999);
xor UO_453 (O_453,N_2929,N_2935);
or UO_454 (O_454,N_2991,N_2977);
or UO_455 (O_455,N_2987,N_2997);
nand UO_456 (O_456,N_2980,N_2953);
or UO_457 (O_457,N_2978,N_2990);
and UO_458 (O_458,N_2954,N_2986);
nand UO_459 (O_459,N_2968,N_2941);
or UO_460 (O_460,N_2942,N_2927);
or UO_461 (O_461,N_2978,N_2936);
and UO_462 (O_462,N_2939,N_2934);
nand UO_463 (O_463,N_2947,N_2964);
xor UO_464 (O_464,N_2993,N_2953);
nand UO_465 (O_465,N_2970,N_2969);
or UO_466 (O_466,N_2974,N_2946);
nor UO_467 (O_467,N_2974,N_2992);
nor UO_468 (O_468,N_2942,N_2937);
and UO_469 (O_469,N_2969,N_2960);
or UO_470 (O_470,N_2961,N_2999);
nand UO_471 (O_471,N_2964,N_2961);
nand UO_472 (O_472,N_2992,N_2967);
and UO_473 (O_473,N_2947,N_2958);
or UO_474 (O_474,N_2928,N_2981);
or UO_475 (O_475,N_2934,N_2926);
and UO_476 (O_476,N_2997,N_2945);
and UO_477 (O_477,N_2962,N_2978);
nand UO_478 (O_478,N_2948,N_2995);
or UO_479 (O_479,N_2993,N_2949);
nand UO_480 (O_480,N_2952,N_2944);
nand UO_481 (O_481,N_2929,N_2968);
and UO_482 (O_482,N_2963,N_2990);
nand UO_483 (O_483,N_2952,N_2963);
nor UO_484 (O_484,N_2972,N_2936);
xnor UO_485 (O_485,N_2978,N_2953);
and UO_486 (O_486,N_2930,N_2965);
nand UO_487 (O_487,N_2931,N_2999);
nor UO_488 (O_488,N_2985,N_2993);
and UO_489 (O_489,N_2953,N_2957);
or UO_490 (O_490,N_2932,N_2992);
nand UO_491 (O_491,N_2987,N_2930);
and UO_492 (O_492,N_2940,N_2938);
xor UO_493 (O_493,N_2933,N_2957);
or UO_494 (O_494,N_2979,N_2925);
or UO_495 (O_495,N_2963,N_2988);
nor UO_496 (O_496,N_2944,N_2969);
and UO_497 (O_497,N_2943,N_2953);
nor UO_498 (O_498,N_2977,N_2976);
xor UO_499 (O_499,N_2951,N_2974);
endmodule