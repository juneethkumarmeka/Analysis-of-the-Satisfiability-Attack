module basic_500_3000_500_5_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_265,In_247);
and U1 (N_1,In_81,In_25);
and U2 (N_2,In_214,In_143);
nor U3 (N_3,In_170,In_173);
or U4 (N_4,In_116,In_200);
nand U5 (N_5,In_105,In_24);
or U6 (N_6,In_49,In_102);
xnor U7 (N_7,In_227,In_103);
nor U8 (N_8,In_15,In_231);
nor U9 (N_9,In_230,In_184);
and U10 (N_10,In_325,In_219);
xnor U11 (N_11,In_248,In_8);
xnor U12 (N_12,In_235,In_221);
and U13 (N_13,In_346,In_62);
and U14 (N_14,In_146,In_109);
and U15 (N_15,In_56,In_157);
or U16 (N_16,In_381,In_349);
nor U17 (N_17,In_107,In_236);
and U18 (N_18,In_17,In_437);
nor U19 (N_19,In_30,In_337);
and U20 (N_20,In_194,In_254);
or U21 (N_21,In_487,In_176);
nand U22 (N_22,In_322,In_493);
xnor U23 (N_23,In_417,In_71);
or U24 (N_24,In_87,In_376);
nand U25 (N_25,In_270,In_141);
and U26 (N_26,In_338,In_388);
xor U27 (N_27,In_140,In_326);
and U28 (N_28,In_51,In_447);
and U29 (N_29,In_492,In_308);
nor U30 (N_30,In_422,In_138);
and U31 (N_31,In_432,In_153);
nand U32 (N_32,In_411,In_54);
nor U33 (N_33,In_11,In_131);
or U34 (N_34,In_22,In_180);
nor U35 (N_35,In_104,In_307);
and U36 (N_36,In_208,In_150);
xnor U37 (N_37,In_452,In_21);
nor U38 (N_38,In_53,In_499);
xor U39 (N_39,In_202,In_234);
or U40 (N_40,In_66,In_498);
and U41 (N_41,In_398,In_240);
or U42 (N_42,In_204,In_195);
nand U43 (N_43,In_471,In_354);
nand U44 (N_44,In_98,In_186);
xnor U45 (N_45,In_343,In_435);
xor U46 (N_46,In_413,In_275);
nand U47 (N_47,In_50,In_122);
or U48 (N_48,In_332,In_392);
nand U49 (N_49,In_191,In_478);
or U50 (N_50,In_277,In_205);
nor U51 (N_51,In_7,In_249);
or U52 (N_52,In_427,In_237);
or U53 (N_53,In_433,In_134);
xor U54 (N_54,In_160,In_100);
xor U55 (N_55,In_166,In_375);
or U56 (N_56,In_189,In_360);
and U57 (N_57,In_350,In_266);
nor U58 (N_58,In_335,In_142);
or U59 (N_59,In_94,In_224);
or U60 (N_60,In_255,In_488);
nand U61 (N_61,In_60,In_286);
or U62 (N_62,In_276,In_319);
or U63 (N_63,In_111,In_347);
xor U64 (N_64,In_260,In_355);
and U65 (N_65,In_179,In_279);
xnor U66 (N_66,In_35,In_4);
or U67 (N_67,In_79,In_465);
nor U68 (N_68,In_440,In_190);
nand U69 (N_69,In_232,In_34);
nor U70 (N_70,In_419,In_164);
and U71 (N_71,In_161,In_269);
or U72 (N_72,In_412,In_245);
nand U73 (N_73,In_1,In_321);
and U74 (N_74,In_213,In_48);
and U75 (N_75,In_373,In_222);
nor U76 (N_76,In_272,In_379);
nand U77 (N_77,In_424,In_409);
and U78 (N_78,In_284,In_340);
nand U79 (N_79,In_348,In_241);
nand U80 (N_80,In_421,In_434);
and U81 (N_81,In_387,In_470);
nor U82 (N_82,In_152,In_239);
nand U83 (N_83,In_108,In_121);
and U84 (N_84,In_3,In_271);
or U85 (N_85,In_77,In_117);
or U86 (N_86,In_404,In_262);
nor U87 (N_87,In_395,In_252);
nor U88 (N_88,In_97,In_410);
and U89 (N_89,In_414,In_13);
and U90 (N_90,In_257,In_210);
nand U91 (N_91,In_75,In_386);
or U92 (N_92,In_26,In_137);
nor U93 (N_93,In_162,In_455);
xnor U94 (N_94,In_441,In_463);
nor U95 (N_95,In_420,In_84);
and U96 (N_96,In_206,In_460);
xnor U97 (N_97,In_361,In_293);
nand U98 (N_98,In_494,In_2);
xor U99 (N_99,In_85,In_74);
nand U100 (N_100,In_144,In_370);
and U101 (N_101,In_211,In_55);
nor U102 (N_102,In_451,In_393);
and U103 (N_103,In_172,In_442);
and U104 (N_104,In_182,In_342);
nand U105 (N_105,In_52,In_174);
nand U106 (N_106,In_242,In_453);
nor U107 (N_107,In_120,In_401);
nor U108 (N_108,In_96,In_132);
and U109 (N_109,In_139,In_358);
nor U110 (N_110,In_44,In_19);
nor U111 (N_111,In_9,In_45);
nor U112 (N_112,In_16,In_368);
or U113 (N_113,In_443,In_93);
xor U114 (N_114,In_264,In_273);
and U115 (N_115,In_253,In_391);
or U116 (N_116,In_445,In_278);
nand U117 (N_117,In_47,In_333);
nor U118 (N_118,In_438,In_446);
nor U119 (N_119,In_396,In_155);
and U120 (N_120,In_197,In_285);
and U121 (N_121,In_251,In_261);
nand U122 (N_122,In_67,In_145);
or U123 (N_123,In_481,In_83);
and U124 (N_124,In_130,In_405);
or U125 (N_125,In_5,In_14);
nor U126 (N_126,In_151,In_324);
and U127 (N_127,In_316,In_95);
nor U128 (N_128,In_135,In_426);
nor U129 (N_129,In_268,In_218);
xor U130 (N_130,In_159,In_344);
nand U131 (N_131,In_362,In_397);
or U132 (N_132,In_439,In_294);
nand U133 (N_133,In_418,In_46);
xnor U134 (N_134,In_288,In_178);
nor U135 (N_135,In_124,In_456);
or U136 (N_136,In_486,In_147);
nand U137 (N_137,In_225,In_385);
nor U138 (N_138,In_450,In_416);
xor U139 (N_139,In_383,In_181);
xor U140 (N_140,In_497,In_199);
or U141 (N_141,In_323,In_298);
nand U142 (N_142,In_462,In_136);
or U143 (N_143,In_457,In_374);
or U144 (N_144,In_317,In_198);
xor U145 (N_145,In_65,In_78);
or U146 (N_146,In_101,In_299);
nand U147 (N_147,In_472,In_246);
xnor U148 (N_148,In_58,In_171);
or U149 (N_149,In_430,In_436);
or U150 (N_150,In_495,In_28);
nor U151 (N_151,In_402,In_390);
or U152 (N_152,In_351,In_209);
xnor U153 (N_153,In_356,In_454);
xnor U154 (N_154,In_37,In_314);
xnor U155 (N_155,In_244,In_267);
and U156 (N_156,In_399,In_217);
nand U157 (N_157,In_90,In_88);
nand U158 (N_158,In_490,In_468);
and U159 (N_159,In_309,In_106);
nor U160 (N_160,In_310,In_18);
or U161 (N_161,In_280,In_43);
and U162 (N_162,In_377,In_489);
xor U163 (N_163,In_364,In_91);
nor U164 (N_164,In_320,In_315);
and U165 (N_165,In_301,In_133);
nor U166 (N_166,In_201,In_367);
and U167 (N_167,In_41,In_148);
or U168 (N_168,In_313,In_287);
nand U169 (N_169,In_86,In_305);
nor U170 (N_170,In_281,In_473);
nand U171 (N_171,In_223,In_233);
nand U172 (N_172,In_425,In_363);
nor U173 (N_173,In_192,In_467);
xor U174 (N_174,In_295,In_482);
xor U175 (N_175,In_458,In_196);
nand U176 (N_176,In_39,In_479);
nand U177 (N_177,In_291,In_114);
or U178 (N_178,In_0,In_444);
xnor U179 (N_179,In_431,In_183);
xor U180 (N_180,In_448,In_68);
and U181 (N_181,In_274,In_384);
xnor U182 (N_182,In_359,In_289);
nor U183 (N_183,In_353,In_331);
nor U184 (N_184,In_163,In_403);
or U185 (N_185,In_327,In_345);
or U186 (N_186,In_318,In_123);
and U187 (N_187,In_169,In_483);
and U188 (N_188,In_57,In_449);
and U189 (N_189,In_27,In_423);
nor U190 (N_190,In_302,In_70);
xnor U191 (N_191,In_12,In_259);
nand U192 (N_192,In_283,In_29);
or U193 (N_193,In_177,In_193);
xor U194 (N_194,In_389,In_466);
or U195 (N_195,In_113,In_36);
nor U196 (N_196,In_185,In_484);
xnor U197 (N_197,In_330,In_115);
xor U198 (N_198,In_175,In_10);
xor U199 (N_199,In_336,In_207);
or U200 (N_200,In_69,In_406);
or U201 (N_201,In_352,In_304);
and U202 (N_202,In_394,In_334);
and U203 (N_203,In_328,In_258);
nand U204 (N_204,In_119,In_464);
xor U205 (N_205,In_42,In_256);
xnor U206 (N_206,In_64,In_33);
xnor U207 (N_207,In_480,In_127);
xnor U208 (N_208,In_6,In_282);
nand U209 (N_209,In_187,In_149);
or U210 (N_210,In_168,In_429);
or U211 (N_211,In_372,In_20);
and U212 (N_212,In_38,In_371);
nor U213 (N_213,In_165,In_80);
and U214 (N_214,In_167,In_408);
or U215 (N_215,In_357,In_112);
or U216 (N_216,In_92,In_243);
and U217 (N_217,In_110,In_188);
xor U218 (N_218,In_329,In_128);
nor U219 (N_219,In_99,In_476);
or U220 (N_220,In_126,In_250);
and U221 (N_221,In_306,In_461);
and U222 (N_222,In_73,In_303);
nand U223 (N_223,In_215,In_365);
nand U224 (N_224,In_382,In_311);
nand U225 (N_225,In_40,In_31);
nand U226 (N_226,In_300,In_89);
and U227 (N_227,In_415,In_459);
xnor U228 (N_228,In_292,In_263);
or U229 (N_229,In_228,In_474);
nand U230 (N_230,In_59,In_216);
nand U231 (N_231,In_220,In_61);
or U232 (N_232,In_496,In_297);
nand U233 (N_233,In_341,In_290);
nand U234 (N_234,In_63,In_339);
and U235 (N_235,In_428,In_118);
nor U236 (N_236,In_312,In_380);
or U237 (N_237,In_76,In_477);
and U238 (N_238,In_156,In_229);
nor U239 (N_239,In_400,In_158);
nand U240 (N_240,In_82,In_32);
nor U241 (N_241,In_366,In_369);
xor U242 (N_242,In_475,In_296);
and U243 (N_243,In_407,In_72);
nor U244 (N_244,In_378,In_469);
or U245 (N_245,In_129,In_125);
or U246 (N_246,In_154,In_226);
nor U247 (N_247,In_485,In_491);
nand U248 (N_248,In_203,In_23);
nor U249 (N_249,In_238,In_212);
and U250 (N_250,In_177,In_434);
or U251 (N_251,In_360,In_487);
nor U252 (N_252,In_471,In_162);
and U253 (N_253,In_28,In_471);
nor U254 (N_254,In_334,In_293);
nor U255 (N_255,In_477,In_231);
nor U256 (N_256,In_470,In_4);
nand U257 (N_257,In_367,In_289);
xor U258 (N_258,In_210,In_37);
xor U259 (N_259,In_370,In_99);
nor U260 (N_260,In_457,In_461);
nand U261 (N_261,In_51,In_358);
and U262 (N_262,In_368,In_476);
and U263 (N_263,In_171,In_165);
nand U264 (N_264,In_70,In_105);
xor U265 (N_265,In_441,In_261);
nor U266 (N_266,In_197,In_114);
and U267 (N_267,In_279,In_159);
or U268 (N_268,In_94,In_446);
nor U269 (N_269,In_157,In_19);
and U270 (N_270,In_263,In_490);
and U271 (N_271,In_325,In_323);
nand U272 (N_272,In_231,In_126);
and U273 (N_273,In_156,In_432);
or U274 (N_274,In_379,In_13);
and U275 (N_275,In_465,In_63);
and U276 (N_276,In_7,In_36);
nand U277 (N_277,In_257,In_296);
nand U278 (N_278,In_240,In_365);
or U279 (N_279,In_161,In_93);
xnor U280 (N_280,In_328,In_224);
and U281 (N_281,In_185,In_149);
nor U282 (N_282,In_219,In_450);
and U283 (N_283,In_352,In_177);
or U284 (N_284,In_81,In_51);
nor U285 (N_285,In_470,In_354);
or U286 (N_286,In_184,In_237);
nor U287 (N_287,In_404,In_336);
or U288 (N_288,In_111,In_309);
nor U289 (N_289,In_91,In_24);
nand U290 (N_290,In_220,In_30);
or U291 (N_291,In_71,In_409);
xnor U292 (N_292,In_64,In_67);
and U293 (N_293,In_128,In_440);
or U294 (N_294,In_193,In_70);
and U295 (N_295,In_170,In_385);
or U296 (N_296,In_391,In_288);
nand U297 (N_297,In_475,In_424);
xor U298 (N_298,In_276,In_235);
nand U299 (N_299,In_408,In_96);
or U300 (N_300,In_317,In_341);
xnor U301 (N_301,In_186,In_141);
nand U302 (N_302,In_88,In_487);
and U303 (N_303,In_499,In_169);
nand U304 (N_304,In_488,In_430);
nor U305 (N_305,In_164,In_469);
or U306 (N_306,In_60,In_159);
nor U307 (N_307,In_88,In_22);
xnor U308 (N_308,In_281,In_341);
nand U309 (N_309,In_288,In_159);
nand U310 (N_310,In_35,In_452);
nand U311 (N_311,In_213,In_202);
xnor U312 (N_312,In_240,In_261);
or U313 (N_313,In_160,In_215);
nor U314 (N_314,In_183,In_258);
nand U315 (N_315,In_335,In_12);
or U316 (N_316,In_496,In_84);
nor U317 (N_317,In_107,In_225);
xor U318 (N_318,In_25,In_340);
xor U319 (N_319,In_155,In_351);
xnor U320 (N_320,In_359,In_429);
and U321 (N_321,In_364,In_210);
xor U322 (N_322,In_80,In_206);
and U323 (N_323,In_138,In_200);
and U324 (N_324,In_126,In_208);
nand U325 (N_325,In_240,In_320);
nor U326 (N_326,In_242,In_456);
xnor U327 (N_327,In_128,In_35);
nor U328 (N_328,In_147,In_45);
nor U329 (N_329,In_83,In_164);
xnor U330 (N_330,In_25,In_479);
xor U331 (N_331,In_42,In_337);
and U332 (N_332,In_406,In_485);
and U333 (N_333,In_294,In_13);
nor U334 (N_334,In_484,In_335);
nand U335 (N_335,In_469,In_158);
nor U336 (N_336,In_463,In_377);
nand U337 (N_337,In_300,In_127);
nand U338 (N_338,In_24,In_117);
nand U339 (N_339,In_69,In_263);
nor U340 (N_340,In_477,In_106);
xor U341 (N_341,In_404,In_99);
nand U342 (N_342,In_360,In_134);
and U343 (N_343,In_488,In_461);
nand U344 (N_344,In_455,In_87);
nand U345 (N_345,In_214,In_481);
or U346 (N_346,In_355,In_282);
and U347 (N_347,In_329,In_28);
nor U348 (N_348,In_323,In_300);
and U349 (N_349,In_126,In_443);
or U350 (N_350,In_277,In_395);
or U351 (N_351,In_4,In_288);
nand U352 (N_352,In_95,In_259);
and U353 (N_353,In_236,In_171);
nor U354 (N_354,In_26,In_428);
nor U355 (N_355,In_126,In_289);
or U356 (N_356,In_76,In_326);
or U357 (N_357,In_255,In_240);
or U358 (N_358,In_27,In_338);
and U359 (N_359,In_313,In_253);
or U360 (N_360,In_451,In_484);
or U361 (N_361,In_378,In_255);
and U362 (N_362,In_323,In_136);
or U363 (N_363,In_199,In_180);
xnor U364 (N_364,In_77,In_12);
nand U365 (N_365,In_182,In_265);
and U366 (N_366,In_380,In_268);
nand U367 (N_367,In_256,In_352);
or U368 (N_368,In_334,In_144);
nand U369 (N_369,In_150,In_406);
or U370 (N_370,In_317,In_353);
or U371 (N_371,In_94,In_368);
xor U372 (N_372,In_440,In_62);
nor U373 (N_373,In_141,In_253);
xor U374 (N_374,In_51,In_406);
or U375 (N_375,In_261,In_338);
or U376 (N_376,In_426,In_82);
xnor U377 (N_377,In_452,In_115);
xnor U378 (N_378,In_349,In_496);
or U379 (N_379,In_359,In_93);
and U380 (N_380,In_365,In_361);
nand U381 (N_381,In_56,In_215);
and U382 (N_382,In_184,In_191);
nor U383 (N_383,In_261,In_88);
xnor U384 (N_384,In_451,In_247);
or U385 (N_385,In_235,In_424);
nor U386 (N_386,In_282,In_158);
nand U387 (N_387,In_57,In_448);
nor U388 (N_388,In_185,In_360);
or U389 (N_389,In_170,In_357);
nand U390 (N_390,In_245,In_160);
xnor U391 (N_391,In_389,In_475);
and U392 (N_392,In_322,In_175);
or U393 (N_393,In_233,In_399);
nand U394 (N_394,In_61,In_314);
or U395 (N_395,In_493,In_34);
xnor U396 (N_396,In_349,In_71);
and U397 (N_397,In_235,In_392);
nor U398 (N_398,In_423,In_331);
and U399 (N_399,In_229,In_93);
xor U400 (N_400,In_488,In_138);
nor U401 (N_401,In_438,In_112);
nand U402 (N_402,In_421,In_316);
and U403 (N_403,In_239,In_267);
nand U404 (N_404,In_467,In_102);
and U405 (N_405,In_72,In_21);
xnor U406 (N_406,In_496,In_363);
and U407 (N_407,In_270,In_259);
nand U408 (N_408,In_155,In_73);
xnor U409 (N_409,In_265,In_343);
or U410 (N_410,In_477,In_99);
nor U411 (N_411,In_421,In_419);
and U412 (N_412,In_60,In_150);
and U413 (N_413,In_423,In_435);
and U414 (N_414,In_292,In_420);
nand U415 (N_415,In_199,In_249);
and U416 (N_416,In_468,In_119);
nand U417 (N_417,In_410,In_473);
xor U418 (N_418,In_483,In_11);
and U419 (N_419,In_278,In_473);
and U420 (N_420,In_499,In_124);
xnor U421 (N_421,In_264,In_8);
nor U422 (N_422,In_313,In_449);
xor U423 (N_423,In_207,In_108);
nand U424 (N_424,In_45,In_65);
nand U425 (N_425,In_411,In_403);
xor U426 (N_426,In_53,In_282);
nor U427 (N_427,In_242,In_163);
or U428 (N_428,In_476,In_132);
nor U429 (N_429,In_371,In_134);
xnor U430 (N_430,In_158,In_314);
nor U431 (N_431,In_246,In_125);
nand U432 (N_432,In_370,In_60);
or U433 (N_433,In_214,In_109);
and U434 (N_434,In_283,In_86);
and U435 (N_435,In_453,In_298);
nor U436 (N_436,In_213,In_179);
nor U437 (N_437,In_247,In_322);
and U438 (N_438,In_312,In_232);
nor U439 (N_439,In_491,In_108);
nand U440 (N_440,In_166,In_348);
and U441 (N_441,In_464,In_187);
nand U442 (N_442,In_396,In_71);
nand U443 (N_443,In_169,In_63);
and U444 (N_444,In_195,In_122);
or U445 (N_445,In_284,In_215);
nor U446 (N_446,In_273,In_326);
and U447 (N_447,In_20,In_318);
nor U448 (N_448,In_37,In_454);
xor U449 (N_449,In_496,In_95);
xnor U450 (N_450,In_28,In_117);
and U451 (N_451,In_293,In_363);
and U452 (N_452,In_71,In_490);
and U453 (N_453,In_486,In_303);
nor U454 (N_454,In_268,In_265);
nand U455 (N_455,In_489,In_12);
nor U456 (N_456,In_83,In_475);
and U457 (N_457,In_270,In_189);
xnor U458 (N_458,In_382,In_393);
or U459 (N_459,In_43,In_30);
xnor U460 (N_460,In_402,In_149);
or U461 (N_461,In_192,In_426);
nand U462 (N_462,In_406,In_275);
xnor U463 (N_463,In_254,In_231);
nor U464 (N_464,In_345,In_94);
and U465 (N_465,In_13,In_295);
nor U466 (N_466,In_251,In_192);
nand U467 (N_467,In_64,In_127);
and U468 (N_468,In_160,In_113);
xor U469 (N_469,In_21,In_156);
or U470 (N_470,In_72,In_14);
or U471 (N_471,In_474,In_343);
nand U472 (N_472,In_182,In_336);
nand U473 (N_473,In_395,In_332);
nand U474 (N_474,In_467,In_291);
xnor U475 (N_475,In_77,In_456);
nand U476 (N_476,In_150,In_105);
and U477 (N_477,In_151,In_371);
and U478 (N_478,In_102,In_269);
or U479 (N_479,In_330,In_302);
nand U480 (N_480,In_230,In_126);
xnor U481 (N_481,In_211,In_104);
and U482 (N_482,In_350,In_481);
nor U483 (N_483,In_102,In_370);
xnor U484 (N_484,In_360,In_202);
xnor U485 (N_485,In_59,In_484);
xnor U486 (N_486,In_481,In_62);
xnor U487 (N_487,In_63,In_326);
nand U488 (N_488,In_139,In_286);
nor U489 (N_489,In_219,In_455);
and U490 (N_490,In_64,In_261);
xnor U491 (N_491,In_115,In_234);
xor U492 (N_492,In_23,In_411);
nand U493 (N_493,In_209,In_311);
and U494 (N_494,In_308,In_413);
and U495 (N_495,In_190,In_246);
or U496 (N_496,In_78,In_218);
xor U497 (N_497,In_52,In_29);
nor U498 (N_498,In_462,In_159);
nand U499 (N_499,In_109,In_477);
and U500 (N_500,In_175,In_335);
nand U501 (N_501,In_224,In_415);
nand U502 (N_502,In_193,In_142);
and U503 (N_503,In_318,In_79);
or U504 (N_504,In_258,In_419);
and U505 (N_505,In_153,In_203);
or U506 (N_506,In_134,In_335);
nand U507 (N_507,In_448,In_274);
nor U508 (N_508,In_152,In_229);
nand U509 (N_509,In_21,In_232);
nor U510 (N_510,In_73,In_181);
and U511 (N_511,In_412,In_106);
nand U512 (N_512,In_75,In_155);
nand U513 (N_513,In_212,In_425);
and U514 (N_514,In_199,In_426);
and U515 (N_515,In_372,In_314);
xnor U516 (N_516,In_260,In_320);
and U517 (N_517,In_268,In_77);
or U518 (N_518,In_235,In_395);
or U519 (N_519,In_62,In_245);
nor U520 (N_520,In_83,In_283);
nor U521 (N_521,In_382,In_245);
xor U522 (N_522,In_82,In_209);
nor U523 (N_523,In_467,In_464);
nor U524 (N_524,In_27,In_201);
or U525 (N_525,In_69,In_59);
xor U526 (N_526,In_339,In_345);
nand U527 (N_527,In_416,In_58);
nand U528 (N_528,In_455,In_164);
xor U529 (N_529,In_247,In_414);
nor U530 (N_530,In_384,In_308);
nand U531 (N_531,In_376,In_215);
nand U532 (N_532,In_1,In_325);
xnor U533 (N_533,In_87,In_320);
and U534 (N_534,In_489,In_417);
and U535 (N_535,In_355,In_119);
and U536 (N_536,In_395,In_151);
and U537 (N_537,In_244,In_413);
nand U538 (N_538,In_246,In_485);
or U539 (N_539,In_25,In_182);
xor U540 (N_540,In_285,In_463);
nand U541 (N_541,In_445,In_15);
nor U542 (N_542,In_44,In_355);
xnor U543 (N_543,In_92,In_447);
and U544 (N_544,In_230,In_433);
nand U545 (N_545,In_447,In_78);
or U546 (N_546,In_374,In_99);
nand U547 (N_547,In_235,In_412);
and U548 (N_548,In_468,In_446);
nand U549 (N_549,In_383,In_224);
nand U550 (N_550,In_142,In_178);
nand U551 (N_551,In_255,In_146);
and U552 (N_552,In_317,In_131);
and U553 (N_553,In_290,In_156);
nor U554 (N_554,In_398,In_171);
nand U555 (N_555,In_198,In_1);
or U556 (N_556,In_153,In_455);
and U557 (N_557,In_201,In_439);
nor U558 (N_558,In_190,In_450);
nor U559 (N_559,In_217,In_426);
xor U560 (N_560,In_99,In_80);
nand U561 (N_561,In_46,In_269);
nand U562 (N_562,In_12,In_432);
or U563 (N_563,In_357,In_403);
xor U564 (N_564,In_240,In_338);
nand U565 (N_565,In_323,In_386);
nand U566 (N_566,In_120,In_128);
nor U567 (N_567,In_132,In_338);
or U568 (N_568,In_288,In_130);
and U569 (N_569,In_251,In_277);
nor U570 (N_570,In_226,In_187);
nand U571 (N_571,In_493,In_211);
nand U572 (N_572,In_273,In_403);
xnor U573 (N_573,In_291,In_157);
nand U574 (N_574,In_434,In_153);
xnor U575 (N_575,In_301,In_466);
and U576 (N_576,In_272,In_121);
xnor U577 (N_577,In_202,In_398);
or U578 (N_578,In_374,In_359);
or U579 (N_579,In_366,In_383);
nor U580 (N_580,In_106,In_328);
nand U581 (N_581,In_30,In_302);
nand U582 (N_582,In_83,In_77);
xnor U583 (N_583,In_226,In_111);
nand U584 (N_584,In_82,In_323);
nor U585 (N_585,In_379,In_388);
nor U586 (N_586,In_17,In_414);
xnor U587 (N_587,In_293,In_31);
nor U588 (N_588,In_436,In_228);
or U589 (N_589,In_257,In_183);
xor U590 (N_590,In_10,In_243);
nand U591 (N_591,In_280,In_328);
nand U592 (N_592,In_473,In_194);
nand U593 (N_593,In_383,In_390);
and U594 (N_594,In_420,In_210);
xor U595 (N_595,In_126,In_74);
and U596 (N_596,In_345,In_265);
nand U597 (N_597,In_83,In_479);
nand U598 (N_598,In_173,In_157);
or U599 (N_599,In_434,In_342);
or U600 (N_600,N_93,N_469);
and U601 (N_601,N_351,N_12);
or U602 (N_602,N_532,N_171);
nor U603 (N_603,N_26,N_394);
and U604 (N_604,N_598,N_110);
xnor U605 (N_605,N_238,N_11);
or U606 (N_606,N_432,N_275);
xnor U607 (N_607,N_262,N_95);
xnor U608 (N_608,N_311,N_373);
xor U609 (N_609,N_267,N_553);
xor U610 (N_610,N_511,N_249);
and U611 (N_611,N_59,N_575);
nor U612 (N_612,N_470,N_542);
and U613 (N_613,N_263,N_415);
nor U614 (N_614,N_458,N_335);
nand U615 (N_615,N_259,N_569);
and U616 (N_616,N_465,N_295);
or U617 (N_617,N_80,N_428);
and U618 (N_618,N_481,N_228);
xor U619 (N_619,N_418,N_375);
nand U620 (N_620,N_65,N_552);
xnor U621 (N_621,N_515,N_451);
xnor U622 (N_622,N_279,N_277);
or U623 (N_623,N_152,N_136);
and U624 (N_624,N_529,N_500);
nand U625 (N_625,N_298,N_597);
nand U626 (N_626,N_146,N_468);
nor U627 (N_627,N_27,N_54);
or U628 (N_628,N_138,N_240);
and U629 (N_629,N_91,N_567);
xor U630 (N_630,N_79,N_431);
nor U631 (N_631,N_245,N_10);
nor U632 (N_632,N_61,N_524);
nor U633 (N_633,N_301,N_292);
and U634 (N_634,N_272,N_304);
xnor U635 (N_635,N_227,N_549);
or U636 (N_636,N_509,N_480);
xnor U637 (N_637,N_105,N_398);
or U638 (N_638,N_571,N_250);
nand U639 (N_639,N_131,N_260);
or U640 (N_640,N_495,N_8);
xor U641 (N_641,N_362,N_220);
and U642 (N_642,N_577,N_324);
nor U643 (N_643,N_380,N_315);
nand U644 (N_644,N_134,N_24);
xor U645 (N_645,N_63,N_452);
nor U646 (N_646,N_256,N_303);
and U647 (N_647,N_169,N_76);
xnor U648 (N_648,N_180,N_165);
nand U649 (N_649,N_416,N_159);
xor U650 (N_650,N_290,N_425);
nand U651 (N_651,N_233,N_563);
xnor U652 (N_652,N_251,N_235);
and U653 (N_653,N_118,N_18);
or U654 (N_654,N_411,N_525);
nor U655 (N_655,N_196,N_331);
nor U656 (N_656,N_217,N_148);
nand U657 (N_657,N_121,N_13);
nand U658 (N_658,N_551,N_51);
or U659 (N_659,N_475,N_439);
nor U660 (N_660,N_316,N_401);
and U661 (N_661,N_589,N_482);
nor U662 (N_662,N_184,N_536);
nor U663 (N_663,N_47,N_492);
nor U664 (N_664,N_281,N_278);
or U665 (N_665,N_269,N_357);
nand U666 (N_666,N_581,N_572);
nor U667 (N_667,N_463,N_62);
nand U668 (N_668,N_173,N_69);
and U669 (N_669,N_58,N_285);
xnor U670 (N_670,N_160,N_122);
and U671 (N_671,N_81,N_3);
and U672 (N_672,N_503,N_406);
nand U673 (N_673,N_20,N_135);
or U674 (N_674,N_109,N_177);
nor U675 (N_675,N_53,N_502);
nand U676 (N_676,N_6,N_283);
xnor U677 (N_677,N_385,N_528);
nor U678 (N_678,N_161,N_151);
xnor U679 (N_679,N_442,N_370);
nand U680 (N_680,N_195,N_381);
nor U681 (N_681,N_38,N_188);
nor U682 (N_682,N_302,N_293);
xnor U683 (N_683,N_57,N_353);
and U684 (N_684,N_545,N_207);
nand U685 (N_685,N_43,N_543);
nand U686 (N_686,N_547,N_143);
nor U687 (N_687,N_319,N_198);
or U688 (N_688,N_371,N_55);
and U689 (N_689,N_450,N_126);
or U690 (N_690,N_153,N_533);
nand U691 (N_691,N_423,N_133);
nand U692 (N_692,N_505,N_102);
xor U693 (N_693,N_211,N_328);
nor U694 (N_694,N_424,N_30);
and U695 (N_695,N_87,N_554);
nand U696 (N_696,N_99,N_265);
and U697 (N_697,N_237,N_300);
or U698 (N_698,N_535,N_590);
and U699 (N_699,N_336,N_224);
xor U700 (N_700,N_125,N_352);
nand U701 (N_701,N_60,N_580);
or U702 (N_702,N_129,N_197);
and U703 (N_703,N_550,N_253);
and U704 (N_704,N_71,N_314);
or U705 (N_705,N_430,N_241);
xnor U706 (N_706,N_408,N_268);
and U707 (N_707,N_142,N_141);
nor U708 (N_708,N_313,N_578);
xor U709 (N_709,N_513,N_579);
nor U710 (N_710,N_203,N_409);
and U711 (N_711,N_527,N_599);
and U712 (N_712,N_396,N_541);
nor U713 (N_713,N_212,N_378);
nor U714 (N_714,N_46,N_417);
nor U715 (N_715,N_364,N_489);
nand U716 (N_716,N_360,N_507);
nor U717 (N_717,N_116,N_44);
nor U718 (N_718,N_181,N_391);
xor U719 (N_719,N_257,N_86);
nor U720 (N_720,N_484,N_150);
xnor U721 (N_721,N_98,N_178);
or U722 (N_722,N_37,N_232);
xnor U723 (N_723,N_462,N_548);
xor U724 (N_724,N_83,N_214);
or U725 (N_725,N_100,N_382);
and U726 (N_726,N_588,N_326);
and U727 (N_727,N_390,N_128);
nor U728 (N_728,N_544,N_174);
xnor U729 (N_729,N_296,N_478);
or U730 (N_730,N_299,N_591);
and U731 (N_731,N_49,N_570);
nor U732 (N_732,N_139,N_137);
and U733 (N_733,N_132,N_187);
xor U734 (N_734,N_555,N_208);
nor U735 (N_735,N_321,N_106);
xor U736 (N_736,N_255,N_246);
nor U737 (N_737,N_466,N_271);
nand U738 (N_738,N_216,N_377);
xnor U739 (N_739,N_127,N_77);
or U740 (N_740,N_52,N_234);
nor U741 (N_741,N_23,N_446);
and U742 (N_742,N_222,N_89);
nand U743 (N_743,N_88,N_460);
and U744 (N_744,N_114,N_70);
xnor U745 (N_745,N_501,N_297);
and U746 (N_746,N_154,N_506);
xnor U747 (N_747,N_386,N_383);
nand U748 (N_748,N_596,N_252);
or U749 (N_749,N_123,N_202);
nand U750 (N_750,N_166,N_183);
nor U751 (N_751,N_68,N_107);
nor U752 (N_752,N_103,N_341);
xnor U753 (N_753,N_45,N_270);
or U754 (N_754,N_434,N_147);
and U755 (N_755,N_537,N_453);
nor U756 (N_756,N_587,N_340);
nor U757 (N_757,N_4,N_429);
nand U758 (N_758,N_402,N_2);
xor U759 (N_759,N_582,N_444);
nand U760 (N_760,N_437,N_16);
nor U761 (N_761,N_163,N_339);
and U762 (N_762,N_50,N_117);
and U763 (N_763,N_155,N_476);
nor U764 (N_764,N_226,N_318);
and U765 (N_765,N_498,N_193);
and U766 (N_766,N_0,N_574);
and U767 (N_767,N_28,N_200);
or U768 (N_768,N_307,N_162);
or U769 (N_769,N_464,N_194);
nand U770 (N_770,N_40,N_517);
xnor U771 (N_771,N_397,N_504);
and U772 (N_772,N_519,N_204);
nand U773 (N_773,N_365,N_546);
xor U774 (N_774,N_101,N_461);
and U775 (N_775,N_113,N_244);
nand U776 (N_776,N_170,N_308);
and U777 (N_777,N_440,N_286);
xnor U778 (N_778,N_231,N_329);
nor U779 (N_779,N_477,N_119);
xor U780 (N_780,N_447,N_562);
nand U781 (N_781,N_449,N_540);
and U782 (N_782,N_454,N_175);
and U783 (N_783,N_90,N_97);
and U784 (N_784,N_512,N_564);
nand U785 (N_785,N_355,N_156);
and U786 (N_786,N_510,N_74);
or U787 (N_787,N_73,N_345);
nand U788 (N_788,N_348,N_48);
xor U789 (N_789,N_309,N_322);
and U790 (N_790,N_158,N_347);
or U791 (N_791,N_523,N_585);
nand U792 (N_792,N_349,N_25);
nor U793 (N_793,N_221,N_145);
xor U794 (N_794,N_435,N_514);
and U795 (N_795,N_559,N_539);
xor U796 (N_796,N_333,N_530);
xnor U797 (N_797,N_414,N_491);
and U798 (N_798,N_366,N_82);
nor U799 (N_799,N_236,N_115);
xor U800 (N_800,N_291,N_108);
xor U801 (N_801,N_258,N_508);
or U802 (N_802,N_359,N_376);
nor U803 (N_803,N_32,N_242);
xor U804 (N_804,N_39,N_337);
and U805 (N_805,N_457,N_199);
nor U806 (N_806,N_410,N_254);
and U807 (N_807,N_179,N_42);
nand U808 (N_808,N_521,N_284);
xor U809 (N_809,N_384,N_310);
or U810 (N_810,N_276,N_164);
nand U811 (N_811,N_593,N_22);
xor U812 (N_812,N_210,N_558);
nand U813 (N_813,N_312,N_342);
and U814 (N_814,N_334,N_248);
nor U815 (N_815,N_534,N_443);
or U816 (N_816,N_361,N_92);
xor U817 (N_817,N_219,N_294);
nor U818 (N_818,N_413,N_7);
xnor U819 (N_819,N_420,N_407);
or U820 (N_820,N_393,N_280);
nor U821 (N_821,N_190,N_191);
and U822 (N_822,N_455,N_531);
nor U823 (N_823,N_387,N_483);
xor U824 (N_824,N_516,N_392);
and U825 (N_825,N_273,N_111);
xor U826 (N_826,N_186,N_405);
nand U827 (N_827,N_168,N_239);
nand U828 (N_828,N_56,N_568);
and U829 (N_829,N_485,N_592);
and U830 (N_830,N_72,N_419);
or U831 (N_831,N_488,N_206);
nand U832 (N_832,N_427,N_167);
nor U833 (N_833,N_225,N_5);
nand U834 (N_834,N_64,N_560);
or U835 (N_835,N_354,N_379);
and U836 (N_836,N_34,N_472);
nor U837 (N_837,N_343,N_209);
nand U838 (N_838,N_306,N_474);
or U839 (N_839,N_467,N_487);
nor U840 (N_840,N_33,N_67);
xnor U841 (N_841,N_94,N_338);
and U842 (N_842,N_104,N_403);
or U843 (N_843,N_584,N_213);
xor U844 (N_844,N_448,N_75);
xnor U845 (N_845,N_243,N_586);
nand U846 (N_846,N_85,N_29);
nor U847 (N_847,N_266,N_96);
or U848 (N_848,N_325,N_287);
or U849 (N_849,N_288,N_486);
xnor U850 (N_850,N_399,N_182);
nor U851 (N_851,N_422,N_566);
or U852 (N_852,N_526,N_573);
nor U853 (N_853,N_176,N_323);
xor U854 (N_854,N_412,N_201);
nand U855 (N_855,N_493,N_31);
and U856 (N_856,N_556,N_445);
and U857 (N_857,N_66,N_14);
or U858 (N_858,N_389,N_395);
xnor U859 (N_859,N_330,N_400);
xnor U860 (N_860,N_594,N_78);
nor U861 (N_861,N_595,N_230);
xnor U862 (N_862,N_149,N_356);
nand U863 (N_863,N_144,N_35);
and U864 (N_864,N_350,N_368);
xnor U865 (N_865,N_218,N_473);
and U866 (N_866,N_441,N_479);
nor U867 (N_867,N_15,N_459);
xnor U868 (N_868,N_520,N_19);
nand U869 (N_869,N_84,N_332);
xor U870 (N_870,N_565,N_433);
or U871 (N_871,N_426,N_367);
nand U872 (N_872,N_305,N_9);
nand U873 (N_873,N_456,N_358);
and U874 (N_874,N_499,N_436);
nor U875 (N_875,N_557,N_229);
nor U876 (N_876,N_247,N_497);
or U877 (N_877,N_327,N_124);
xor U878 (N_878,N_374,N_185);
and U879 (N_879,N_112,N_496);
or U880 (N_880,N_189,N_421);
and U881 (N_881,N_471,N_369);
xnor U882 (N_882,N_21,N_494);
xor U883 (N_883,N_261,N_538);
or U884 (N_884,N_172,N_41);
xnor U885 (N_885,N_215,N_317);
xnor U886 (N_886,N_518,N_264);
or U887 (N_887,N_522,N_192);
xnor U888 (N_888,N_157,N_130);
nor U889 (N_889,N_583,N_346);
nor U890 (N_890,N_223,N_1);
or U891 (N_891,N_404,N_388);
and U892 (N_892,N_36,N_363);
nor U893 (N_893,N_274,N_282);
nor U894 (N_894,N_490,N_17);
nor U895 (N_895,N_140,N_561);
xnor U896 (N_896,N_576,N_438);
and U897 (N_897,N_205,N_320);
nand U898 (N_898,N_120,N_344);
or U899 (N_899,N_372,N_289);
xnor U900 (N_900,N_261,N_376);
xnor U901 (N_901,N_443,N_182);
nor U902 (N_902,N_496,N_473);
and U903 (N_903,N_369,N_197);
nand U904 (N_904,N_588,N_456);
xor U905 (N_905,N_555,N_521);
and U906 (N_906,N_288,N_591);
and U907 (N_907,N_326,N_141);
xnor U908 (N_908,N_449,N_59);
and U909 (N_909,N_438,N_407);
or U910 (N_910,N_370,N_403);
or U911 (N_911,N_159,N_109);
and U912 (N_912,N_533,N_387);
nand U913 (N_913,N_179,N_572);
nor U914 (N_914,N_438,N_86);
xnor U915 (N_915,N_279,N_174);
nand U916 (N_916,N_480,N_228);
nor U917 (N_917,N_458,N_279);
xor U918 (N_918,N_388,N_236);
nand U919 (N_919,N_464,N_554);
and U920 (N_920,N_469,N_138);
or U921 (N_921,N_482,N_338);
and U922 (N_922,N_426,N_101);
nand U923 (N_923,N_129,N_74);
nor U924 (N_924,N_390,N_93);
nor U925 (N_925,N_247,N_418);
and U926 (N_926,N_398,N_306);
and U927 (N_927,N_593,N_494);
nand U928 (N_928,N_249,N_115);
nor U929 (N_929,N_245,N_86);
or U930 (N_930,N_538,N_339);
nand U931 (N_931,N_410,N_261);
nor U932 (N_932,N_423,N_593);
nor U933 (N_933,N_179,N_505);
xnor U934 (N_934,N_152,N_232);
nor U935 (N_935,N_103,N_144);
or U936 (N_936,N_11,N_568);
and U937 (N_937,N_48,N_373);
nor U938 (N_938,N_243,N_196);
xnor U939 (N_939,N_359,N_181);
nor U940 (N_940,N_91,N_514);
and U941 (N_941,N_518,N_437);
or U942 (N_942,N_571,N_178);
and U943 (N_943,N_232,N_486);
nor U944 (N_944,N_594,N_102);
or U945 (N_945,N_538,N_232);
nand U946 (N_946,N_112,N_89);
xor U947 (N_947,N_185,N_483);
xor U948 (N_948,N_373,N_555);
nor U949 (N_949,N_571,N_130);
nand U950 (N_950,N_428,N_70);
nor U951 (N_951,N_255,N_367);
nor U952 (N_952,N_68,N_467);
nor U953 (N_953,N_532,N_95);
or U954 (N_954,N_526,N_431);
and U955 (N_955,N_594,N_320);
and U956 (N_956,N_547,N_568);
and U957 (N_957,N_578,N_571);
and U958 (N_958,N_414,N_464);
nor U959 (N_959,N_313,N_555);
nor U960 (N_960,N_12,N_101);
nor U961 (N_961,N_298,N_545);
or U962 (N_962,N_215,N_483);
nor U963 (N_963,N_452,N_349);
nor U964 (N_964,N_336,N_143);
nand U965 (N_965,N_477,N_480);
and U966 (N_966,N_223,N_545);
nand U967 (N_967,N_432,N_17);
nand U968 (N_968,N_183,N_20);
or U969 (N_969,N_95,N_281);
nor U970 (N_970,N_510,N_272);
xor U971 (N_971,N_326,N_483);
xor U972 (N_972,N_32,N_108);
xor U973 (N_973,N_257,N_295);
nor U974 (N_974,N_145,N_96);
and U975 (N_975,N_345,N_467);
nand U976 (N_976,N_305,N_206);
xor U977 (N_977,N_408,N_386);
or U978 (N_978,N_596,N_540);
and U979 (N_979,N_373,N_198);
and U980 (N_980,N_343,N_337);
nand U981 (N_981,N_166,N_272);
and U982 (N_982,N_149,N_223);
xor U983 (N_983,N_317,N_493);
nand U984 (N_984,N_570,N_511);
nor U985 (N_985,N_86,N_505);
nand U986 (N_986,N_241,N_404);
nor U987 (N_987,N_37,N_214);
nor U988 (N_988,N_398,N_11);
or U989 (N_989,N_283,N_398);
or U990 (N_990,N_215,N_511);
xor U991 (N_991,N_12,N_384);
nor U992 (N_992,N_394,N_497);
nand U993 (N_993,N_437,N_405);
nor U994 (N_994,N_450,N_547);
xnor U995 (N_995,N_331,N_451);
nand U996 (N_996,N_112,N_272);
nor U997 (N_997,N_551,N_131);
or U998 (N_998,N_476,N_142);
nor U999 (N_999,N_585,N_459);
and U1000 (N_1000,N_573,N_12);
xnor U1001 (N_1001,N_209,N_450);
xor U1002 (N_1002,N_174,N_439);
or U1003 (N_1003,N_556,N_592);
and U1004 (N_1004,N_155,N_567);
and U1005 (N_1005,N_0,N_169);
nor U1006 (N_1006,N_465,N_101);
and U1007 (N_1007,N_72,N_294);
and U1008 (N_1008,N_227,N_183);
xnor U1009 (N_1009,N_313,N_151);
or U1010 (N_1010,N_190,N_229);
xor U1011 (N_1011,N_542,N_546);
or U1012 (N_1012,N_300,N_594);
nand U1013 (N_1013,N_464,N_63);
or U1014 (N_1014,N_333,N_219);
and U1015 (N_1015,N_348,N_227);
and U1016 (N_1016,N_547,N_582);
and U1017 (N_1017,N_133,N_176);
nand U1018 (N_1018,N_465,N_517);
nand U1019 (N_1019,N_276,N_357);
and U1020 (N_1020,N_289,N_36);
xor U1021 (N_1021,N_382,N_279);
nor U1022 (N_1022,N_134,N_462);
nor U1023 (N_1023,N_409,N_350);
nor U1024 (N_1024,N_492,N_529);
xor U1025 (N_1025,N_290,N_516);
nor U1026 (N_1026,N_244,N_371);
xor U1027 (N_1027,N_224,N_488);
nor U1028 (N_1028,N_105,N_171);
or U1029 (N_1029,N_584,N_59);
nor U1030 (N_1030,N_152,N_403);
or U1031 (N_1031,N_385,N_282);
and U1032 (N_1032,N_254,N_137);
nand U1033 (N_1033,N_38,N_584);
or U1034 (N_1034,N_424,N_38);
or U1035 (N_1035,N_119,N_227);
xnor U1036 (N_1036,N_590,N_127);
nand U1037 (N_1037,N_394,N_19);
xnor U1038 (N_1038,N_447,N_30);
nand U1039 (N_1039,N_65,N_515);
nand U1040 (N_1040,N_304,N_421);
or U1041 (N_1041,N_310,N_589);
nor U1042 (N_1042,N_530,N_346);
nor U1043 (N_1043,N_94,N_29);
and U1044 (N_1044,N_389,N_578);
xor U1045 (N_1045,N_522,N_450);
and U1046 (N_1046,N_384,N_43);
nor U1047 (N_1047,N_558,N_320);
nor U1048 (N_1048,N_446,N_553);
nor U1049 (N_1049,N_85,N_127);
nand U1050 (N_1050,N_23,N_293);
nand U1051 (N_1051,N_109,N_304);
xor U1052 (N_1052,N_230,N_269);
and U1053 (N_1053,N_470,N_362);
or U1054 (N_1054,N_561,N_525);
and U1055 (N_1055,N_96,N_512);
nand U1056 (N_1056,N_21,N_13);
xnor U1057 (N_1057,N_384,N_588);
or U1058 (N_1058,N_415,N_428);
xor U1059 (N_1059,N_495,N_384);
xnor U1060 (N_1060,N_241,N_131);
nor U1061 (N_1061,N_143,N_149);
nand U1062 (N_1062,N_202,N_32);
nand U1063 (N_1063,N_383,N_211);
xor U1064 (N_1064,N_417,N_290);
xnor U1065 (N_1065,N_88,N_42);
nor U1066 (N_1066,N_319,N_190);
nor U1067 (N_1067,N_203,N_425);
xor U1068 (N_1068,N_468,N_258);
nor U1069 (N_1069,N_512,N_364);
nor U1070 (N_1070,N_167,N_178);
nor U1071 (N_1071,N_164,N_292);
xnor U1072 (N_1072,N_270,N_542);
nor U1073 (N_1073,N_69,N_272);
xor U1074 (N_1074,N_339,N_269);
xnor U1075 (N_1075,N_193,N_449);
nor U1076 (N_1076,N_295,N_399);
and U1077 (N_1077,N_282,N_125);
nand U1078 (N_1078,N_593,N_293);
xor U1079 (N_1079,N_503,N_432);
or U1080 (N_1080,N_321,N_52);
xnor U1081 (N_1081,N_197,N_469);
nand U1082 (N_1082,N_215,N_515);
nor U1083 (N_1083,N_488,N_231);
nor U1084 (N_1084,N_372,N_197);
nand U1085 (N_1085,N_479,N_490);
nor U1086 (N_1086,N_187,N_55);
xnor U1087 (N_1087,N_115,N_547);
or U1088 (N_1088,N_149,N_448);
xnor U1089 (N_1089,N_528,N_78);
and U1090 (N_1090,N_449,N_230);
nand U1091 (N_1091,N_318,N_525);
nand U1092 (N_1092,N_142,N_371);
xor U1093 (N_1093,N_222,N_538);
nand U1094 (N_1094,N_461,N_153);
nand U1095 (N_1095,N_26,N_481);
and U1096 (N_1096,N_553,N_576);
and U1097 (N_1097,N_412,N_316);
and U1098 (N_1098,N_379,N_217);
nand U1099 (N_1099,N_292,N_592);
xor U1100 (N_1100,N_587,N_588);
and U1101 (N_1101,N_529,N_69);
or U1102 (N_1102,N_306,N_285);
nand U1103 (N_1103,N_340,N_331);
and U1104 (N_1104,N_573,N_462);
nand U1105 (N_1105,N_224,N_400);
xnor U1106 (N_1106,N_582,N_312);
and U1107 (N_1107,N_282,N_307);
and U1108 (N_1108,N_235,N_41);
and U1109 (N_1109,N_599,N_75);
and U1110 (N_1110,N_495,N_598);
nor U1111 (N_1111,N_127,N_267);
nor U1112 (N_1112,N_381,N_525);
nor U1113 (N_1113,N_595,N_224);
xor U1114 (N_1114,N_482,N_143);
and U1115 (N_1115,N_480,N_287);
and U1116 (N_1116,N_429,N_115);
and U1117 (N_1117,N_558,N_377);
nand U1118 (N_1118,N_502,N_404);
nor U1119 (N_1119,N_520,N_470);
xnor U1120 (N_1120,N_473,N_171);
and U1121 (N_1121,N_398,N_324);
nor U1122 (N_1122,N_180,N_502);
xor U1123 (N_1123,N_563,N_387);
or U1124 (N_1124,N_368,N_77);
or U1125 (N_1125,N_84,N_325);
nor U1126 (N_1126,N_9,N_203);
or U1127 (N_1127,N_463,N_113);
and U1128 (N_1128,N_375,N_356);
nor U1129 (N_1129,N_447,N_438);
xnor U1130 (N_1130,N_323,N_68);
nor U1131 (N_1131,N_156,N_87);
or U1132 (N_1132,N_524,N_484);
and U1133 (N_1133,N_25,N_458);
nand U1134 (N_1134,N_429,N_93);
and U1135 (N_1135,N_408,N_489);
nor U1136 (N_1136,N_456,N_486);
or U1137 (N_1137,N_496,N_435);
or U1138 (N_1138,N_447,N_279);
nor U1139 (N_1139,N_410,N_185);
and U1140 (N_1140,N_405,N_263);
nor U1141 (N_1141,N_448,N_115);
nor U1142 (N_1142,N_298,N_310);
nand U1143 (N_1143,N_465,N_46);
and U1144 (N_1144,N_297,N_507);
xnor U1145 (N_1145,N_192,N_373);
nor U1146 (N_1146,N_41,N_104);
nand U1147 (N_1147,N_584,N_279);
and U1148 (N_1148,N_259,N_5);
and U1149 (N_1149,N_282,N_505);
or U1150 (N_1150,N_540,N_371);
and U1151 (N_1151,N_252,N_487);
and U1152 (N_1152,N_560,N_39);
nand U1153 (N_1153,N_471,N_136);
or U1154 (N_1154,N_354,N_189);
or U1155 (N_1155,N_222,N_128);
and U1156 (N_1156,N_251,N_321);
or U1157 (N_1157,N_63,N_447);
or U1158 (N_1158,N_253,N_233);
nor U1159 (N_1159,N_97,N_198);
xor U1160 (N_1160,N_426,N_117);
or U1161 (N_1161,N_374,N_174);
or U1162 (N_1162,N_148,N_140);
nand U1163 (N_1163,N_428,N_282);
or U1164 (N_1164,N_516,N_515);
or U1165 (N_1165,N_118,N_183);
nor U1166 (N_1166,N_130,N_163);
xor U1167 (N_1167,N_387,N_554);
nand U1168 (N_1168,N_223,N_406);
or U1169 (N_1169,N_118,N_522);
xor U1170 (N_1170,N_203,N_371);
nor U1171 (N_1171,N_404,N_332);
nand U1172 (N_1172,N_47,N_451);
and U1173 (N_1173,N_88,N_367);
nand U1174 (N_1174,N_493,N_532);
xnor U1175 (N_1175,N_521,N_125);
nor U1176 (N_1176,N_240,N_140);
nand U1177 (N_1177,N_290,N_355);
and U1178 (N_1178,N_441,N_423);
nor U1179 (N_1179,N_189,N_324);
nand U1180 (N_1180,N_432,N_123);
xnor U1181 (N_1181,N_353,N_121);
and U1182 (N_1182,N_159,N_553);
and U1183 (N_1183,N_546,N_419);
and U1184 (N_1184,N_480,N_410);
nand U1185 (N_1185,N_227,N_31);
nand U1186 (N_1186,N_594,N_33);
nor U1187 (N_1187,N_276,N_519);
nand U1188 (N_1188,N_270,N_49);
or U1189 (N_1189,N_428,N_1);
nand U1190 (N_1190,N_255,N_423);
and U1191 (N_1191,N_249,N_526);
nand U1192 (N_1192,N_87,N_478);
and U1193 (N_1193,N_178,N_441);
nor U1194 (N_1194,N_226,N_24);
nand U1195 (N_1195,N_218,N_349);
nor U1196 (N_1196,N_259,N_37);
or U1197 (N_1197,N_140,N_23);
nand U1198 (N_1198,N_93,N_97);
or U1199 (N_1199,N_213,N_264);
nand U1200 (N_1200,N_1130,N_1029);
xnor U1201 (N_1201,N_645,N_909);
and U1202 (N_1202,N_819,N_1093);
and U1203 (N_1203,N_991,N_1118);
nand U1204 (N_1204,N_693,N_1014);
or U1205 (N_1205,N_1179,N_706);
xnor U1206 (N_1206,N_671,N_803);
nand U1207 (N_1207,N_1018,N_1135);
xnor U1208 (N_1208,N_1160,N_964);
or U1209 (N_1209,N_1182,N_990);
nor U1210 (N_1210,N_683,N_949);
or U1211 (N_1211,N_732,N_710);
nor U1212 (N_1212,N_777,N_1131);
and U1213 (N_1213,N_1086,N_845);
or U1214 (N_1214,N_751,N_979);
nor U1215 (N_1215,N_1180,N_602);
or U1216 (N_1216,N_1147,N_832);
nand U1217 (N_1217,N_878,N_656);
xor U1218 (N_1218,N_1146,N_1003);
and U1219 (N_1219,N_755,N_1006);
nor U1220 (N_1220,N_1149,N_1079);
or U1221 (N_1221,N_824,N_858);
nand U1222 (N_1222,N_676,N_1030);
nor U1223 (N_1223,N_677,N_1171);
and U1224 (N_1224,N_1110,N_806);
xor U1225 (N_1225,N_1032,N_1158);
xnor U1226 (N_1226,N_700,N_1067);
nor U1227 (N_1227,N_1038,N_1096);
and U1228 (N_1228,N_735,N_932);
nand U1229 (N_1229,N_925,N_1043);
xor U1230 (N_1230,N_881,N_1150);
or U1231 (N_1231,N_969,N_892);
and U1232 (N_1232,N_943,N_885);
nor U1233 (N_1233,N_609,N_601);
nor U1234 (N_1234,N_811,N_1066);
and U1235 (N_1235,N_813,N_708);
and U1236 (N_1236,N_864,N_744);
nor U1237 (N_1237,N_1152,N_940);
and U1238 (N_1238,N_955,N_1101);
and U1239 (N_1239,N_821,N_1194);
or U1240 (N_1240,N_1049,N_1021);
nor U1241 (N_1241,N_768,N_971);
or U1242 (N_1242,N_1071,N_1092);
and U1243 (N_1243,N_673,N_1129);
nor U1244 (N_1244,N_884,N_1088);
xnor U1245 (N_1245,N_801,N_668);
or U1246 (N_1246,N_996,N_1002);
and U1247 (N_1247,N_1060,N_1157);
nand U1248 (N_1248,N_626,N_1120);
nand U1249 (N_1249,N_1119,N_654);
nand U1250 (N_1250,N_1124,N_770);
xnor U1251 (N_1251,N_665,N_787);
nand U1252 (N_1252,N_703,N_818);
xor U1253 (N_1253,N_915,N_1056);
or U1254 (N_1254,N_1022,N_728);
nand U1255 (N_1255,N_793,N_946);
nand U1256 (N_1256,N_653,N_678);
or U1257 (N_1257,N_953,N_775);
or U1258 (N_1258,N_675,N_1132);
xnor U1259 (N_1259,N_786,N_958);
nand U1260 (N_1260,N_906,N_1186);
nand U1261 (N_1261,N_1185,N_1191);
or U1262 (N_1262,N_758,N_869);
nor U1263 (N_1263,N_760,N_887);
nor U1264 (N_1264,N_666,N_746);
or U1265 (N_1265,N_1197,N_967);
xor U1266 (N_1266,N_743,N_1063);
nand U1267 (N_1267,N_600,N_895);
nand U1268 (N_1268,N_960,N_757);
nand U1269 (N_1269,N_618,N_1000);
or U1270 (N_1270,N_1122,N_822);
nand U1271 (N_1271,N_937,N_855);
or U1272 (N_1272,N_748,N_800);
nor U1273 (N_1273,N_1062,N_672);
and U1274 (N_1274,N_817,N_1076);
or U1275 (N_1275,N_712,N_1047);
and U1276 (N_1276,N_1069,N_759);
nor U1277 (N_1277,N_641,N_1137);
and U1278 (N_1278,N_891,N_688);
or U1279 (N_1279,N_919,N_1104);
nor U1280 (N_1280,N_898,N_1077);
and U1281 (N_1281,N_805,N_719);
xor U1282 (N_1282,N_1184,N_608);
xor U1283 (N_1283,N_1116,N_985);
nand U1284 (N_1284,N_938,N_1070);
or U1285 (N_1285,N_1164,N_779);
nor U1286 (N_1286,N_1126,N_970);
or U1287 (N_1287,N_997,N_773);
or U1288 (N_1288,N_1143,N_731);
nand U1289 (N_1289,N_788,N_603);
nor U1290 (N_1290,N_1098,N_1177);
and U1291 (N_1291,N_689,N_650);
or U1292 (N_1292,N_918,N_947);
and U1293 (N_1293,N_1153,N_908);
xor U1294 (N_1294,N_738,N_716);
and U1295 (N_1295,N_942,N_655);
xnor U1296 (N_1296,N_1169,N_747);
nand U1297 (N_1297,N_802,N_863);
xnor U1298 (N_1298,N_1145,N_880);
xor U1299 (N_1299,N_717,N_1199);
or U1300 (N_1300,N_722,N_781);
and U1301 (N_1301,N_823,N_890);
xnor U1302 (N_1302,N_630,N_922);
xnor U1303 (N_1303,N_988,N_1019);
nand U1304 (N_1304,N_1100,N_927);
nand U1305 (N_1305,N_1161,N_1073);
and U1306 (N_1306,N_771,N_1105);
nand U1307 (N_1307,N_1007,N_715);
xor U1308 (N_1308,N_1040,N_923);
nand U1309 (N_1309,N_691,N_935);
and U1310 (N_1310,N_1141,N_726);
xor U1311 (N_1311,N_669,N_1046);
or U1312 (N_1312,N_622,N_707);
or U1313 (N_1313,N_1136,N_632);
xnor U1314 (N_1314,N_934,N_1176);
xnor U1315 (N_1315,N_658,N_612);
nor U1316 (N_1316,N_635,N_861);
nor U1317 (N_1317,N_931,N_692);
nand U1318 (N_1318,N_1192,N_1111);
nand U1319 (N_1319,N_705,N_701);
and U1320 (N_1320,N_981,N_1151);
nand U1321 (N_1321,N_1080,N_1178);
nor U1322 (N_1322,N_910,N_648);
and U1323 (N_1323,N_1121,N_1005);
or U1324 (N_1324,N_896,N_664);
and U1325 (N_1325,N_784,N_1193);
and U1326 (N_1326,N_1095,N_999);
or U1327 (N_1327,N_611,N_815);
nand U1328 (N_1328,N_1154,N_926);
nand U1329 (N_1329,N_1196,N_627);
xor U1330 (N_1330,N_961,N_634);
nor U1331 (N_1331,N_1175,N_972);
or U1332 (N_1332,N_734,N_889);
or U1333 (N_1333,N_1008,N_619);
nor U1334 (N_1334,N_902,N_974);
or U1335 (N_1335,N_742,N_977);
nor U1336 (N_1336,N_1195,N_750);
nand U1337 (N_1337,N_986,N_862);
nor U1338 (N_1338,N_745,N_844);
and U1339 (N_1339,N_852,N_762);
or U1340 (N_1340,N_761,N_1091);
or U1341 (N_1341,N_637,N_903);
nor U1342 (N_1342,N_1159,N_694);
nor U1343 (N_1343,N_1036,N_1011);
nand U1344 (N_1344,N_737,N_936);
xor U1345 (N_1345,N_1156,N_1050);
xor U1346 (N_1346,N_767,N_829);
and U1347 (N_1347,N_605,N_980);
nand U1348 (N_1348,N_956,N_739);
and U1349 (N_1349,N_962,N_992);
nor U1350 (N_1350,N_1134,N_1107);
and U1351 (N_1351,N_789,N_1103);
or U1352 (N_1352,N_644,N_686);
nand U1353 (N_1353,N_831,N_749);
nand U1354 (N_1354,N_838,N_752);
or U1355 (N_1355,N_1045,N_1081);
xor U1356 (N_1356,N_1125,N_973);
nand U1357 (N_1357,N_1028,N_839);
or U1358 (N_1358,N_1140,N_1115);
nand U1359 (N_1359,N_670,N_1189);
or U1360 (N_1360,N_1017,N_1012);
and U1361 (N_1361,N_944,N_1106);
nand U1362 (N_1362,N_1139,N_901);
nand U1363 (N_1363,N_649,N_888);
nor U1364 (N_1364,N_1170,N_1138);
and U1365 (N_1365,N_776,N_1167);
xor U1366 (N_1366,N_850,N_924);
and U1367 (N_1367,N_1001,N_1072);
or U1368 (N_1368,N_948,N_772);
nand U1369 (N_1369,N_1168,N_639);
xnor U1370 (N_1370,N_659,N_1031);
and U1371 (N_1371,N_636,N_867);
nand U1372 (N_1372,N_640,N_975);
and U1373 (N_1373,N_1037,N_965);
xnor U1374 (N_1374,N_921,N_812);
and U1375 (N_1375,N_778,N_1155);
or U1376 (N_1376,N_904,N_856);
xor U1377 (N_1377,N_785,N_667);
nor U1378 (N_1378,N_780,N_685);
nor U1379 (N_1379,N_1054,N_623);
nand U1380 (N_1380,N_769,N_872);
and U1381 (N_1381,N_916,N_621);
nand U1382 (N_1382,N_870,N_998);
or U1383 (N_1383,N_913,N_941);
or U1384 (N_1384,N_729,N_854);
nor U1385 (N_1385,N_723,N_1048);
nor U1386 (N_1386,N_905,N_957);
nor U1387 (N_1387,N_709,N_741);
nand U1388 (N_1388,N_1165,N_1035);
xnor U1389 (N_1389,N_687,N_1113);
nor U1390 (N_1390,N_1004,N_804);
xnor U1391 (N_1391,N_994,N_1112);
and U1392 (N_1392,N_1042,N_836);
nor U1393 (N_1393,N_1065,N_1166);
or U1394 (N_1394,N_657,N_1033);
or U1395 (N_1395,N_899,N_933);
and U1396 (N_1396,N_756,N_1057);
nand U1397 (N_1397,N_1144,N_851);
and U1398 (N_1398,N_826,N_846);
xnor U1399 (N_1399,N_978,N_849);
nand U1400 (N_1400,N_827,N_1068);
nor U1401 (N_1401,N_727,N_914);
xnor U1402 (N_1402,N_625,N_1023);
xor U1403 (N_1403,N_848,N_1198);
or U1404 (N_1404,N_711,N_753);
nand U1405 (N_1405,N_929,N_763);
or U1406 (N_1406,N_920,N_610);
nand U1407 (N_1407,N_840,N_794);
or U1408 (N_1408,N_1085,N_930);
xnor U1409 (N_1409,N_764,N_606);
and U1410 (N_1410,N_1055,N_1114);
and U1411 (N_1411,N_865,N_681);
xnor U1412 (N_1412,N_843,N_1020);
and U1413 (N_1413,N_871,N_917);
or U1414 (N_1414,N_1190,N_1034);
nor U1415 (N_1415,N_882,N_911);
and U1416 (N_1416,N_809,N_1010);
nand U1417 (N_1417,N_983,N_718);
and U1418 (N_1418,N_1097,N_1075);
nor U1419 (N_1419,N_945,N_893);
and U1420 (N_1420,N_1024,N_987);
nor U1421 (N_1421,N_682,N_1009);
nand U1422 (N_1422,N_690,N_950);
xor U1423 (N_1423,N_680,N_993);
or U1424 (N_1424,N_959,N_995);
nor U1425 (N_1425,N_754,N_695);
xnor U1426 (N_1426,N_820,N_631);
nor U1427 (N_1427,N_1083,N_1026);
nand U1428 (N_1428,N_835,N_642);
and U1429 (N_1429,N_797,N_873);
nand U1430 (N_1430,N_816,N_1074);
nor U1431 (N_1431,N_853,N_799);
xnor U1432 (N_1432,N_1123,N_963);
or U1433 (N_1433,N_783,N_1162);
and U1434 (N_1434,N_1084,N_720);
nand U1435 (N_1435,N_798,N_828);
nand U1436 (N_1436,N_875,N_1053);
and U1437 (N_1437,N_679,N_1025);
and U1438 (N_1438,N_1087,N_662);
or U1439 (N_1439,N_646,N_1041);
nor U1440 (N_1440,N_814,N_968);
nor U1441 (N_1441,N_808,N_982);
nor U1442 (N_1442,N_837,N_833);
nand U1443 (N_1443,N_1173,N_841);
nand U1444 (N_1444,N_614,N_766);
nor U1445 (N_1445,N_647,N_790);
xor U1446 (N_1446,N_886,N_696);
nand U1447 (N_1447,N_1109,N_733);
or U1448 (N_1448,N_730,N_651);
nor U1449 (N_1449,N_1148,N_661);
xnor U1450 (N_1450,N_1188,N_1044);
or U1451 (N_1451,N_1102,N_1133);
xnor U1452 (N_1452,N_1174,N_866);
xnor U1453 (N_1453,N_714,N_663);
xnor U1454 (N_1454,N_795,N_652);
nor U1455 (N_1455,N_1090,N_697);
nor U1456 (N_1456,N_604,N_713);
or U1457 (N_1457,N_907,N_616);
nand U1458 (N_1458,N_1108,N_633);
nand U1459 (N_1459,N_1027,N_1127);
and U1460 (N_1460,N_1183,N_825);
xnor U1461 (N_1461,N_1059,N_900);
and U1462 (N_1462,N_954,N_1016);
nor U1463 (N_1463,N_912,N_740);
nor U1464 (N_1464,N_859,N_660);
or U1465 (N_1465,N_704,N_834);
nor U1466 (N_1466,N_1117,N_1064);
nor U1467 (N_1467,N_1082,N_868);
or U1468 (N_1468,N_1099,N_807);
xor U1469 (N_1469,N_879,N_928);
nor U1470 (N_1470,N_952,N_684);
xnor U1471 (N_1471,N_620,N_725);
and U1472 (N_1472,N_874,N_847);
or U1473 (N_1473,N_613,N_699);
and U1474 (N_1474,N_883,N_894);
and U1475 (N_1475,N_1187,N_966);
xor U1476 (N_1476,N_1051,N_774);
or U1477 (N_1477,N_615,N_951);
xor U1478 (N_1478,N_842,N_830);
nor U1479 (N_1479,N_796,N_1039);
nand U1480 (N_1480,N_1094,N_724);
and U1481 (N_1481,N_698,N_1013);
nor U1482 (N_1482,N_860,N_810);
and U1483 (N_1483,N_876,N_702);
and U1484 (N_1484,N_765,N_1163);
nand U1485 (N_1485,N_1015,N_617);
or U1486 (N_1486,N_791,N_857);
nor U1487 (N_1487,N_607,N_721);
xor U1488 (N_1488,N_792,N_1128);
nor U1489 (N_1489,N_976,N_877);
nand U1490 (N_1490,N_782,N_1078);
nor U1491 (N_1491,N_674,N_939);
nor U1492 (N_1492,N_643,N_1061);
xnor U1493 (N_1493,N_1052,N_629);
xor U1494 (N_1494,N_1172,N_1181);
nor U1495 (N_1495,N_628,N_638);
nand U1496 (N_1496,N_624,N_1058);
nand U1497 (N_1497,N_989,N_1142);
xnor U1498 (N_1498,N_984,N_1089);
and U1499 (N_1499,N_897,N_736);
or U1500 (N_1500,N_966,N_647);
or U1501 (N_1501,N_998,N_837);
xnor U1502 (N_1502,N_837,N_605);
or U1503 (N_1503,N_1139,N_681);
xor U1504 (N_1504,N_815,N_624);
nor U1505 (N_1505,N_1007,N_1049);
or U1506 (N_1506,N_1162,N_806);
and U1507 (N_1507,N_1091,N_1145);
nor U1508 (N_1508,N_1031,N_955);
nor U1509 (N_1509,N_793,N_1103);
xnor U1510 (N_1510,N_674,N_1005);
nor U1511 (N_1511,N_1016,N_671);
nand U1512 (N_1512,N_630,N_673);
nand U1513 (N_1513,N_651,N_994);
xnor U1514 (N_1514,N_980,N_674);
xor U1515 (N_1515,N_621,N_1100);
and U1516 (N_1516,N_978,N_1104);
or U1517 (N_1517,N_1044,N_843);
nor U1518 (N_1518,N_1071,N_738);
and U1519 (N_1519,N_629,N_787);
and U1520 (N_1520,N_669,N_890);
and U1521 (N_1521,N_976,N_1017);
or U1522 (N_1522,N_890,N_1146);
and U1523 (N_1523,N_636,N_899);
nor U1524 (N_1524,N_628,N_927);
and U1525 (N_1525,N_1174,N_966);
and U1526 (N_1526,N_907,N_664);
or U1527 (N_1527,N_897,N_742);
nand U1528 (N_1528,N_995,N_776);
xor U1529 (N_1529,N_708,N_893);
nand U1530 (N_1530,N_812,N_739);
nand U1531 (N_1531,N_1087,N_751);
or U1532 (N_1532,N_781,N_709);
and U1533 (N_1533,N_850,N_817);
xor U1534 (N_1534,N_722,N_943);
xor U1535 (N_1535,N_680,N_683);
xnor U1536 (N_1536,N_906,N_853);
or U1537 (N_1537,N_926,N_653);
nand U1538 (N_1538,N_705,N_996);
or U1539 (N_1539,N_651,N_1173);
xor U1540 (N_1540,N_885,N_1138);
or U1541 (N_1541,N_875,N_1028);
nand U1542 (N_1542,N_1050,N_788);
and U1543 (N_1543,N_957,N_840);
or U1544 (N_1544,N_813,N_710);
nor U1545 (N_1545,N_828,N_997);
and U1546 (N_1546,N_1167,N_815);
or U1547 (N_1547,N_1147,N_1073);
nand U1548 (N_1548,N_1019,N_1182);
nand U1549 (N_1549,N_1006,N_916);
xnor U1550 (N_1550,N_690,N_725);
nand U1551 (N_1551,N_869,N_656);
xor U1552 (N_1552,N_1083,N_825);
and U1553 (N_1553,N_1112,N_711);
xnor U1554 (N_1554,N_643,N_1034);
and U1555 (N_1555,N_1026,N_826);
and U1556 (N_1556,N_1145,N_959);
and U1557 (N_1557,N_833,N_778);
and U1558 (N_1558,N_1151,N_603);
nor U1559 (N_1559,N_1059,N_885);
nor U1560 (N_1560,N_724,N_647);
and U1561 (N_1561,N_1154,N_718);
xor U1562 (N_1562,N_662,N_993);
or U1563 (N_1563,N_824,N_671);
nor U1564 (N_1564,N_1115,N_965);
xnor U1565 (N_1565,N_739,N_964);
and U1566 (N_1566,N_748,N_1172);
and U1567 (N_1567,N_693,N_1095);
nand U1568 (N_1568,N_950,N_971);
or U1569 (N_1569,N_690,N_663);
xor U1570 (N_1570,N_806,N_1067);
nand U1571 (N_1571,N_1017,N_963);
xnor U1572 (N_1572,N_1055,N_1101);
or U1573 (N_1573,N_738,N_832);
or U1574 (N_1574,N_664,N_728);
nor U1575 (N_1575,N_1056,N_759);
or U1576 (N_1576,N_860,N_861);
and U1577 (N_1577,N_802,N_766);
nand U1578 (N_1578,N_1078,N_929);
or U1579 (N_1579,N_732,N_958);
and U1580 (N_1580,N_1015,N_1122);
or U1581 (N_1581,N_876,N_1072);
nand U1582 (N_1582,N_923,N_688);
nand U1583 (N_1583,N_794,N_1029);
nor U1584 (N_1584,N_679,N_958);
nand U1585 (N_1585,N_1196,N_852);
xnor U1586 (N_1586,N_677,N_944);
or U1587 (N_1587,N_768,N_903);
and U1588 (N_1588,N_839,N_1018);
or U1589 (N_1589,N_955,N_762);
xnor U1590 (N_1590,N_979,N_702);
or U1591 (N_1591,N_765,N_729);
nor U1592 (N_1592,N_1126,N_1142);
nor U1593 (N_1593,N_700,N_1055);
nor U1594 (N_1594,N_921,N_793);
nor U1595 (N_1595,N_1088,N_1189);
and U1596 (N_1596,N_804,N_1030);
nand U1597 (N_1597,N_1075,N_730);
or U1598 (N_1598,N_994,N_669);
nand U1599 (N_1599,N_978,N_606);
nor U1600 (N_1600,N_1072,N_765);
or U1601 (N_1601,N_1176,N_906);
nand U1602 (N_1602,N_921,N_1055);
or U1603 (N_1603,N_722,N_836);
nor U1604 (N_1604,N_631,N_658);
xor U1605 (N_1605,N_614,N_1035);
and U1606 (N_1606,N_925,N_1192);
or U1607 (N_1607,N_1115,N_820);
or U1608 (N_1608,N_836,N_697);
nor U1609 (N_1609,N_605,N_1131);
nor U1610 (N_1610,N_1027,N_991);
xnor U1611 (N_1611,N_854,N_779);
and U1612 (N_1612,N_1157,N_1095);
xnor U1613 (N_1613,N_680,N_950);
and U1614 (N_1614,N_1154,N_661);
and U1615 (N_1615,N_1137,N_626);
nor U1616 (N_1616,N_832,N_1078);
nand U1617 (N_1617,N_745,N_1156);
and U1618 (N_1618,N_1027,N_1038);
xor U1619 (N_1619,N_719,N_1116);
nor U1620 (N_1620,N_705,N_1012);
nor U1621 (N_1621,N_678,N_639);
and U1622 (N_1622,N_1168,N_901);
nand U1623 (N_1623,N_798,N_769);
and U1624 (N_1624,N_1072,N_993);
xnor U1625 (N_1625,N_1125,N_1064);
xor U1626 (N_1626,N_943,N_625);
and U1627 (N_1627,N_689,N_1062);
nor U1628 (N_1628,N_620,N_894);
and U1629 (N_1629,N_765,N_901);
nor U1630 (N_1630,N_633,N_626);
and U1631 (N_1631,N_1082,N_725);
xnor U1632 (N_1632,N_719,N_817);
and U1633 (N_1633,N_952,N_600);
and U1634 (N_1634,N_678,N_1131);
and U1635 (N_1635,N_1138,N_883);
nand U1636 (N_1636,N_943,N_634);
nor U1637 (N_1637,N_697,N_1113);
and U1638 (N_1638,N_1081,N_843);
or U1639 (N_1639,N_630,N_945);
and U1640 (N_1640,N_785,N_973);
or U1641 (N_1641,N_708,N_953);
nand U1642 (N_1642,N_998,N_815);
xor U1643 (N_1643,N_789,N_1067);
nor U1644 (N_1644,N_808,N_1123);
nor U1645 (N_1645,N_791,N_941);
or U1646 (N_1646,N_821,N_914);
nand U1647 (N_1647,N_1011,N_789);
or U1648 (N_1648,N_969,N_1166);
xnor U1649 (N_1649,N_893,N_872);
and U1650 (N_1650,N_662,N_1125);
or U1651 (N_1651,N_812,N_773);
and U1652 (N_1652,N_698,N_631);
xnor U1653 (N_1653,N_986,N_680);
and U1654 (N_1654,N_888,N_680);
xnor U1655 (N_1655,N_1019,N_982);
nand U1656 (N_1656,N_1183,N_1065);
or U1657 (N_1657,N_837,N_672);
nand U1658 (N_1658,N_1015,N_1043);
and U1659 (N_1659,N_1081,N_654);
or U1660 (N_1660,N_863,N_673);
or U1661 (N_1661,N_1060,N_739);
nor U1662 (N_1662,N_901,N_1017);
or U1663 (N_1663,N_1154,N_979);
or U1664 (N_1664,N_1199,N_1080);
nand U1665 (N_1665,N_780,N_742);
nand U1666 (N_1666,N_622,N_1098);
and U1667 (N_1667,N_838,N_802);
xor U1668 (N_1668,N_887,N_996);
nor U1669 (N_1669,N_834,N_762);
nor U1670 (N_1670,N_752,N_977);
nand U1671 (N_1671,N_1093,N_1151);
or U1672 (N_1672,N_1188,N_991);
nand U1673 (N_1673,N_635,N_626);
nor U1674 (N_1674,N_640,N_1023);
or U1675 (N_1675,N_911,N_822);
or U1676 (N_1676,N_1104,N_655);
and U1677 (N_1677,N_1072,N_1014);
xor U1678 (N_1678,N_609,N_993);
or U1679 (N_1679,N_931,N_1164);
nand U1680 (N_1680,N_943,N_1057);
nor U1681 (N_1681,N_1177,N_1122);
nor U1682 (N_1682,N_1197,N_1093);
xor U1683 (N_1683,N_827,N_691);
and U1684 (N_1684,N_718,N_804);
and U1685 (N_1685,N_655,N_815);
nand U1686 (N_1686,N_1108,N_863);
nand U1687 (N_1687,N_729,N_869);
and U1688 (N_1688,N_911,N_1081);
nor U1689 (N_1689,N_1090,N_1066);
xnor U1690 (N_1690,N_1132,N_758);
and U1691 (N_1691,N_908,N_678);
and U1692 (N_1692,N_1109,N_1092);
nand U1693 (N_1693,N_874,N_776);
nand U1694 (N_1694,N_898,N_776);
nand U1695 (N_1695,N_805,N_652);
nor U1696 (N_1696,N_1159,N_943);
nand U1697 (N_1697,N_1064,N_613);
xnor U1698 (N_1698,N_886,N_686);
nor U1699 (N_1699,N_627,N_724);
xnor U1700 (N_1700,N_647,N_695);
or U1701 (N_1701,N_1093,N_830);
xnor U1702 (N_1702,N_886,N_790);
or U1703 (N_1703,N_714,N_1021);
and U1704 (N_1704,N_809,N_1187);
nor U1705 (N_1705,N_682,N_1084);
and U1706 (N_1706,N_770,N_889);
nand U1707 (N_1707,N_1034,N_789);
and U1708 (N_1708,N_788,N_714);
xor U1709 (N_1709,N_707,N_1123);
and U1710 (N_1710,N_742,N_1053);
nand U1711 (N_1711,N_707,N_1159);
or U1712 (N_1712,N_1058,N_1098);
nor U1713 (N_1713,N_871,N_660);
xnor U1714 (N_1714,N_617,N_1125);
and U1715 (N_1715,N_754,N_1078);
nor U1716 (N_1716,N_761,N_1172);
nor U1717 (N_1717,N_1049,N_640);
or U1718 (N_1718,N_920,N_759);
and U1719 (N_1719,N_712,N_1116);
and U1720 (N_1720,N_770,N_858);
xor U1721 (N_1721,N_613,N_614);
or U1722 (N_1722,N_646,N_777);
and U1723 (N_1723,N_831,N_773);
xnor U1724 (N_1724,N_1176,N_777);
and U1725 (N_1725,N_740,N_725);
and U1726 (N_1726,N_1154,N_619);
or U1727 (N_1727,N_957,N_1161);
or U1728 (N_1728,N_1064,N_1147);
nor U1729 (N_1729,N_1104,N_902);
or U1730 (N_1730,N_944,N_606);
or U1731 (N_1731,N_687,N_756);
or U1732 (N_1732,N_1099,N_967);
or U1733 (N_1733,N_914,N_1016);
or U1734 (N_1734,N_1111,N_831);
nor U1735 (N_1735,N_648,N_1137);
nor U1736 (N_1736,N_1156,N_664);
and U1737 (N_1737,N_652,N_847);
or U1738 (N_1738,N_636,N_1156);
xnor U1739 (N_1739,N_1035,N_878);
nor U1740 (N_1740,N_997,N_731);
nor U1741 (N_1741,N_695,N_1149);
nand U1742 (N_1742,N_1142,N_770);
xor U1743 (N_1743,N_1172,N_1104);
and U1744 (N_1744,N_1017,N_915);
or U1745 (N_1745,N_1181,N_715);
or U1746 (N_1746,N_707,N_602);
or U1747 (N_1747,N_948,N_732);
nand U1748 (N_1748,N_1102,N_713);
nor U1749 (N_1749,N_703,N_685);
nand U1750 (N_1750,N_782,N_1001);
and U1751 (N_1751,N_1029,N_1118);
xor U1752 (N_1752,N_626,N_676);
and U1753 (N_1753,N_828,N_882);
and U1754 (N_1754,N_992,N_964);
nand U1755 (N_1755,N_1030,N_1113);
and U1756 (N_1756,N_783,N_770);
xnor U1757 (N_1757,N_944,N_1114);
or U1758 (N_1758,N_780,N_1075);
nor U1759 (N_1759,N_1078,N_848);
nor U1760 (N_1760,N_1031,N_1019);
and U1761 (N_1761,N_915,N_625);
nand U1762 (N_1762,N_856,N_1064);
or U1763 (N_1763,N_832,N_696);
nor U1764 (N_1764,N_979,N_1066);
xnor U1765 (N_1765,N_723,N_908);
nand U1766 (N_1766,N_687,N_780);
or U1767 (N_1767,N_706,N_752);
xor U1768 (N_1768,N_1068,N_851);
nor U1769 (N_1769,N_1192,N_1095);
nand U1770 (N_1770,N_819,N_806);
nand U1771 (N_1771,N_752,N_693);
nand U1772 (N_1772,N_1037,N_895);
nand U1773 (N_1773,N_1077,N_630);
nand U1774 (N_1774,N_692,N_649);
xor U1775 (N_1775,N_641,N_831);
xor U1776 (N_1776,N_994,N_739);
xor U1777 (N_1777,N_1135,N_910);
and U1778 (N_1778,N_622,N_633);
nand U1779 (N_1779,N_1058,N_771);
or U1780 (N_1780,N_648,N_1001);
nand U1781 (N_1781,N_1178,N_877);
and U1782 (N_1782,N_745,N_621);
nor U1783 (N_1783,N_900,N_656);
xor U1784 (N_1784,N_980,N_1026);
nor U1785 (N_1785,N_1065,N_805);
or U1786 (N_1786,N_979,N_732);
nand U1787 (N_1787,N_1096,N_908);
or U1788 (N_1788,N_1090,N_679);
or U1789 (N_1789,N_831,N_1004);
nand U1790 (N_1790,N_983,N_1118);
nand U1791 (N_1791,N_983,N_1091);
and U1792 (N_1792,N_719,N_1123);
xor U1793 (N_1793,N_1085,N_1160);
nand U1794 (N_1794,N_744,N_620);
nand U1795 (N_1795,N_961,N_1022);
nor U1796 (N_1796,N_1016,N_1018);
nor U1797 (N_1797,N_617,N_994);
or U1798 (N_1798,N_848,N_1122);
or U1799 (N_1799,N_708,N_967);
nand U1800 (N_1800,N_1679,N_1260);
xnor U1801 (N_1801,N_1768,N_1456);
nor U1802 (N_1802,N_1306,N_1254);
and U1803 (N_1803,N_1744,N_1544);
nand U1804 (N_1804,N_1760,N_1675);
or U1805 (N_1805,N_1654,N_1413);
or U1806 (N_1806,N_1496,N_1606);
or U1807 (N_1807,N_1258,N_1738);
nor U1808 (N_1808,N_1766,N_1502);
nand U1809 (N_1809,N_1761,N_1214);
and U1810 (N_1810,N_1390,N_1526);
xnor U1811 (N_1811,N_1696,N_1750);
nor U1812 (N_1812,N_1657,N_1314);
xor U1813 (N_1813,N_1718,N_1685);
nand U1814 (N_1814,N_1200,N_1579);
xnor U1815 (N_1815,N_1333,N_1653);
and U1816 (N_1816,N_1498,N_1722);
and U1817 (N_1817,N_1274,N_1469);
nand U1818 (N_1818,N_1490,N_1512);
or U1819 (N_1819,N_1478,N_1706);
nand U1820 (N_1820,N_1533,N_1743);
or U1821 (N_1821,N_1624,N_1580);
nor U1822 (N_1822,N_1326,N_1302);
nand U1823 (N_1823,N_1610,N_1735);
and U1824 (N_1824,N_1730,N_1499);
xnor U1825 (N_1825,N_1694,N_1228);
nand U1826 (N_1826,N_1466,N_1224);
xnor U1827 (N_1827,N_1692,N_1748);
nand U1828 (N_1828,N_1446,N_1375);
nand U1829 (N_1829,N_1680,N_1351);
xnor U1830 (N_1830,N_1383,N_1355);
nor U1831 (N_1831,N_1441,N_1204);
nor U1832 (N_1832,N_1514,N_1364);
xor U1833 (N_1833,N_1763,N_1263);
or U1834 (N_1834,N_1546,N_1797);
and U1835 (N_1835,N_1251,N_1795);
or U1836 (N_1836,N_1420,N_1434);
nand U1837 (N_1837,N_1290,N_1244);
and U1838 (N_1838,N_1703,N_1242);
nand U1839 (N_1839,N_1739,N_1361);
nor U1840 (N_1840,N_1246,N_1362);
xor U1841 (N_1841,N_1505,N_1749);
or U1842 (N_1842,N_1764,N_1367);
nand U1843 (N_1843,N_1210,N_1597);
and U1844 (N_1844,N_1540,N_1756);
nor U1845 (N_1845,N_1477,N_1377);
and U1846 (N_1846,N_1671,N_1359);
nor U1847 (N_1847,N_1495,N_1527);
or U1848 (N_1848,N_1457,N_1381);
nand U1849 (N_1849,N_1372,N_1796);
and U1850 (N_1850,N_1645,N_1658);
or U1851 (N_1851,N_1423,N_1243);
or U1852 (N_1852,N_1369,N_1465);
nand U1853 (N_1853,N_1269,N_1710);
nor U1854 (N_1854,N_1471,N_1287);
xor U1855 (N_1855,N_1438,N_1531);
nor U1856 (N_1856,N_1614,N_1767);
nand U1857 (N_1857,N_1412,N_1480);
and U1858 (N_1858,N_1568,N_1239);
nand U1859 (N_1859,N_1599,N_1648);
or U1860 (N_1860,N_1617,N_1476);
and U1861 (N_1861,N_1299,N_1389);
xnor U1862 (N_1862,N_1395,N_1538);
nor U1863 (N_1863,N_1222,N_1785);
nor U1864 (N_1864,N_1387,N_1698);
and U1865 (N_1865,N_1406,N_1550);
or U1866 (N_1866,N_1399,N_1668);
and U1867 (N_1867,N_1264,N_1393);
nor U1868 (N_1868,N_1651,N_1319);
and U1869 (N_1869,N_1640,N_1684);
and U1870 (N_1870,N_1325,N_1588);
or U1871 (N_1871,N_1259,N_1691);
nand U1872 (N_1872,N_1549,N_1408);
xnor U1873 (N_1873,N_1601,N_1202);
or U1874 (N_1874,N_1330,N_1635);
and U1875 (N_1875,N_1596,N_1230);
nand U1876 (N_1876,N_1340,N_1252);
xnor U1877 (N_1877,N_1632,N_1708);
nand U1878 (N_1878,N_1545,N_1422);
and U1879 (N_1879,N_1255,N_1225);
nor U1880 (N_1880,N_1537,N_1752);
nor U1881 (N_1881,N_1391,N_1384);
nor U1882 (N_1882,N_1539,N_1575);
nor U1883 (N_1883,N_1425,N_1633);
nand U1884 (N_1884,N_1553,N_1256);
nor U1885 (N_1885,N_1655,N_1517);
and U1886 (N_1886,N_1304,N_1709);
nor U1887 (N_1887,N_1374,N_1247);
nor U1888 (N_1888,N_1707,N_1649);
nor U1889 (N_1889,N_1404,N_1699);
nand U1890 (N_1890,N_1687,N_1778);
nor U1891 (N_1891,N_1672,N_1628);
or U1892 (N_1892,N_1598,N_1379);
nand U1893 (N_1893,N_1564,N_1736);
nor U1894 (N_1894,N_1737,N_1382);
and U1895 (N_1895,N_1573,N_1720);
nand U1896 (N_1896,N_1558,N_1639);
nor U1897 (N_1897,N_1343,N_1682);
or U1898 (N_1898,N_1317,N_1620);
nor U1899 (N_1899,N_1728,N_1449);
and U1900 (N_1900,N_1603,N_1700);
or U1901 (N_1901,N_1556,N_1626);
nand U1902 (N_1902,N_1448,N_1217);
nand U1903 (N_1903,N_1547,N_1392);
and U1904 (N_1904,N_1616,N_1509);
nor U1905 (N_1905,N_1669,N_1534);
nor U1906 (N_1906,N_1370,N_1551);
and U1907 (N_1907,N_1627,N_1543);
or U1908 (N_1908,N_1646,N_1265);
xor U1909 (N_1909,N_1405,N_1461);
and U1910 (N_1910,N_1226,N_1245);
nand U1911 (N_1911,N_1289,N_1332);
and U1912 (N_1912,N_1552,N_1308);
and U1913 (N_1913,N_1294,N_1237);
nor U1914 (N_1914,N_1535,N_1702);
xnor U1915 (N_1915,N_1286,N_1716);
xor U1916 (N_1916,N_1291,N_1773);
xor U1917 (N_1917,N_1410,N_1746);
and U1918 (N_1918,N_1713,N_1634);
nand U1919 (N_1919,N_1631,N_1486);
xor U1920 (N_1920,N_1799,N_1206);
or U1921 (N_1921,N_1316,N_1723);
and U1922 (N_1922,N_1402,N_1777);
and U1923 (N_1923,N_1636,N_1201);
xnor U1924 (N_1924,N_1417,N_1279);
nand U1925 (N_1925,N_1798,N_1510);
or U1926 (N_1926,N_1401,N_1437);
and U1927 (N_1927,N_1674,N_1781);
nand U1928 (N_1928,N_1775,N_1312);
nor U1929 (N_1929,N_1366,N_1789);
nand U1930 (N_1930,N_1611,N_1585);
or U1931 (N_1931,N_1421,N_1725);
nor U1932 (N_1932,N_1350,N_1429);
nand U1933 (N_1933,N_1378,N_1337);
nand U1934 (N_1934,N_1721,N_1492);
and U1935 (N_1935,N_1213,N_1688);
and U1936 (N_1936,N_1285,N_1637);
nor U1937 (N_1937,N_1605,N_1458);
nand U1938 (N_1938,N_1373,N_1270);
nor U1939 (N_1939,N_1705,N_1661);
or U1940 (N_1940,N_1755,N_1557);
or U1941 (N_1941,N_1371,N_1792);
or U1942 (N_1942,N_1347,N_1442);
xor U1943 (N_1943,N_1583,N_1283);
nand U1944 (N_1944,N_1460,N_1276);
nor U1945 (N_1945,N_1528,N_1336);
and U1946 (N_1946,N_1227,N_1307);
or U1947 (N_1947,N_1338,N_1300);
nand U1948 (N_1948,N_1587,N_1677);
xor U1949 (N_1949,N_1334,N_1418);
nor U1950 (N_1950,N_1787,N_1462);
and U1951 (N_1951,N_1426,N_1615);
and U1952 (N_1952,N_1602,N_1318);
or U1953 (N_1953,N_1467,N_1485);
nand U1954 (N_1954,N_1211,N_1443);
or U1955 (N_1955,N_1591,N_1686);
or U1956 (N_1956,N_1650,N_1488);
nand U1957 (N_1957,N_1253,N_1542);
or U1958 (N_1958,N_1428,N_1786);
xor U1959 (N_1959,N_1439,N_1576);
and U1960 (N_1960,N_1560,N_1315);
nand U1961 (N_1961,N_1641,N_1298);
or U1962 (N_1962,N_1363,N_1323);
nand U1963 (N_1963,N_1747,N_1278);
and U1964 (N_1964,N_1681,N_1209);
or U1965 (N_1965,N_1303,N_1695);
or U1966 (N_1966,N_1578,N_1453);
and U1967 (N_1967,N_1335,N_1501);
xnor U1968 (N_1968,N_1345,N_1380);
nor U1969 (N_1969,N_1772,N_1569);
nor U1970 (N_1970,N_1508,N_1562);
and U1971 (N_1971,N_1280,N_1740);
nor U1972 (N_1972,N_1741,N_1652);
and U1973 (N_1973,N_1444,N_1670);
or U1974 (N_1974,N_1475,N_1277);
nor U1975 (N_1975,N_1301,N_1581);
or U1976 (N_1976,N_1563,N_1574);
nand U1977 (N_1977,N_1577,N_1416);
xnor U1978 (N_1978,N_1793,N_1205);
or U1979 (N_1979,N_1288,N_1548);
xor U1980 (N_1980,N_1223,N_1665);
or U1981 (N_1981,N_1500,N_1292);
or U1982 (N_1982,N_1567,N_1296);
or U1983 (N_1983,N_1497,N_1479);
nand U1984 (N_1984,N_1396,N_1436);
xnor U1985 (N_1985,N_1348,N_1493);
and U1986 (N_1986,N_1594,N_1281);
or U1987 (N_1987,N_1663,N_1431);
nor U1988 (N_1988,N_1250,N_1629);
nor U1989 (N_1989,N_1284,N_1731);
xor U1990 (N_1990,N_1595,N_1689);
nor U1991 (N_1991,N_1690,N_1742);
and U1992 (N_1992,N_1241,N_1791);
and U1993 (N_1993,N_1612,N_1782);
or U1994 (N_1994,N_1403,N_1662);
or U1995 (N_1995,N_1275,N_1608);
nand U1996 (N_1996,N_1607,N_1790);
or U1997 (N_1997,N_1236,N_1697);
nand U1998 (N_1998,N_1714,N_1513);
or U1999 (N_1999,N_1229,N_1464);
xor U2000 (N_2000,N_1704,N_1238);
nor U2001 (N_2001,N_1221,N_1729);
nand U2002 (N_2002,N_1765,N_1432);
nand U2003 (N_2003,N_1309,N_1207);
nor U2004 (N_2004,N_1571,N_1232);
nor U2005 (N_2005,N_1613,N_1257);
or U2006 (N_2006,N_1305,N_1523);
or U2007 (N_2007,N_1504,N_1711);
and U2008 (N_2008,N_1667,N_1435);
and U2009 (N_2009,N_1745,N_1582);
xor U2010 (N_2010,N_1656,N_1774);
nor U2011 (N_2011,N_1400,N_1693);
or U2012 (N_2012,N_1430,N_1481);
xnor U2013 (N_2013,N_1419,N_1758);
xor U2014 (N_2014,N_1394,N_1356);
nor U2015 (N_2015,N_1727,N_1724);
and U2016 (N_2016,N_1249,N_1491);
xnor U2017 (N_2017,N_1203,N_1536);
and U2018 (N_2018,N_1503,N_1376);
or U2019 (N_2019,N_1385,N_1218);
or U2020 (N_2020,N_1521,N_1365);
nor U2021 (N_2021,N_1683,N_1516);
xnor U2022 (N_2022,N_1676,N_1463);
nor U2023 (N_2023,N_1311,N_1555);
xnor U2024 (N_2024,N_1342,N_1762);
xnor U2025 (N_2025,N_1433,N_1489);
nor U2026 (N_2026,N_1261,N_1339);
nand U2027 (N_2027,N_1484,N_1644);
nor U2028 (N_2028,N_1518,N_1451);
and U2029 (N_2029,N_1715,N_1212);
and U2030 (N_2030,N_1407,N_1454);
xor U2031 (N_2031,N_1647,N_1638);
or U2032 (N_2032,N_1271,N_1712);
and U2033 (N_2033,N_1566,N_1570);
and U2034 (N_2034,N_1231,N_1630);
or U2035 (N_2035,N_1520,N_1754);
nand U2036 (N_2036,N_1732,N_1532);
nor U2037 (N_2037,N_1625,N_1324);
xor U2038 (N_2038,N_1483,N_1297);
and U2039 (N_2039,N_1388,N_1659);
nand U2040 (N_2040,N_1559,N_1701);
and U2041 (N_2041,N_1589,N_1219);
xnor U2042 (N_2042,N_1515,N_1320);
nand U2043 (N_2043,N_1445,N_1673);
or U2044 (N_2044,N_1240,N_1726);
nor U2045 (N_2045,N_1660,N_1664);
and U2046 (N_2046,N_1235,N_1530);
or U2047 (N_2047,N_1427,N_1776);
and U2048 (N_2048,N_1354,N_1414);
nand U2049 (N_2049,N_1233,N_1440);
nand U2050 (N_2050,N_1592,N_1216);
xor U2051 (N_2051,N_1397,N_1473);
or U2052 (N_2052,N_1352,N_1328);
xor U2053 (N_2053,N_1751,N_1783);
nand U2054 (N_2054,N_1618,N_1220);
and U2055 (N_2055,N_1719,N_1409);
xor U2056 (N_2056,N_1282,N_1621);
nor U2057 (N_2057,N_1368,N_1519);
and U2058 (N_2058,N_1507,N_1353);
xor U2059 (N_2059,N_1215,N_1358);
and U2060 (N_2060,N_1554,N_1262);
nor U2061 (N_2061,N_1310,N_1590);
and U2062 (N_2062,N_1759,N_1529);
nand U2063 (N_2063,N_1619,N_1734);
nor U2064 (N_2064,N_1586,N_1459);
nor U2065 (N_2065,N_1266,N_1494);
or U2066 (N_2066,N_1313,N_1511);
nor U2067 (N_2067,N_1468,N_1522);
xor U2068 (N_2068,N_1349,N_1600);
nor U2069 (N_2069,N_1455,N_1525);
nor U2070 (N_2070,N_1541,N_1572);
or U2071 (N_2071,N_1487,N_1293);
nand U2072 (N_2072,N_1643,N_1561);
nand U2073 (N_2073,N_1565,N_1450);
and U2074 (N_2074,N_1272,N_1360);
and U2075 (N_2075,N_1452,N_1779);
or U2076 (N_2076,N_1678,N_1447);
and U2077 (N_2077,N_1357,N_1474);
nor U2078 (N_2078,N_1733,N_1780);
nor U2079 (N_2079,N_1346,N_1208);
nor U2080 (N_2080,N_1470,N_1482);
and U2081 (N_2081,N_1415,N_1506);
nand U2082 (N_2082,N_1584,N_1472);
xnor U2083 (N_2083,N_1268,N_1341);
nor U2084 (N_2084,N_1788,N_1593);
and U2085 (N_2085,N_1524,N_1769);
nand U2086 (N_2086,N_1295,N_1770);
nand U2087 (N_2087,N_1331,N_1642);
and U2088 (N_2088,N_1604,N_1267);
and U2089 (N_2089,N_1344,N_1321);
and U2090 (N_2090,N_1273,N_1424);
nand U2091 (N_2091,N_1784,N_1771);
xor U2092 (N_2092,N_1622,N_1609);
or U2093 (N_2093,N_1322,N_1327);
nor U2094 (N_2094,N_1757,N_1386);
nand U2095 (N_2095,N_1717,N_1411);
and U2096 (N_2096,N_1666,N_1248);
xnor U2097 (N_2097,N_1398,N_1329);
xor U2098 (N_2098,N_1794,N_1623);
and U2099 (N_2099,N_1234,N_1753);
or U2100 (N_2100,N_1424,N_1366);
and U2101 (N_2101,N_1331,N_1743);
xor U2102 (N_2102,N_1547,N_1357);
xnor U2103 (N_2103,N_1611,N_1660);
nor U2104 (N_2104,N_1575,N_1636);
xnor U2105 (N_2105,N_1753,N_1272);
xnor U2106 (N_2106,N_1231,N_1516);
and U2107 (N_2107,N_1294,N_1212);
nor U2108 (N_2108,N_1214,N_1230);
nand U2109 (N_2109,N_1329,N_1523);
or U2110 (N_2110,N_1319,N_1709);
nor U2111 (N_2111,N_1604,N_1684);
and U2112 (N_2112,N_1548,N_1585);
and U2113 (N_2113,N_1386,N_1788);
and U2114 (N_2114,N_1686,N_1320);
nor U2115 (N_2115,N_1409,N_1569);
nor U2116 (N_2116,N_1312,N_1260);
nor U2117 (N_2117,N_1527,N_1785);
or U2118 (N_2118,N_1483,N_1548);
or U2119 (N_2119,N_1572,N_1526);
xnor U2120 (N_2120,N_1350,N_1660);
and U2121 (N_2121,N_1636,N_1382);
nand U2122 (N_2122,N_1542,N_1681);
xnor U2123 (N_2123,N_1638,N_1675);
nor U2124 (N_2124,N_1396,N_1573);
and U2125 (N_2125,N_1423,N_1416);
or U2126 (N_2126,N_1711,N_1756);
nor U2127 (N_2127,N_1504,N_1654);
nand U2128 (N_2128,N_1249,N_1569);
nor U2129 (N_2129,N_1420,N_1780);
nand U2130 (N_2130,N_1493,N_1290);
or U2131 (N_2131,N_1767,N_1430);
nand U2132 (N_2132,N_1239,N_1547);
and U2133 (N_2133,N_1432,N_1430);
nand U2134 (N_2134,N_1677,N_1788);
or U2135 (N_2135,N_1772,N_1694);
nand U2136 (N_2136,N_1586,N_1544);
nand U2137 (N_2137,N_1310,N_1366);
and U2138 (N_2138,N_1432,N_1502);
and U2139 (N_2139,N_1494,N_1619);
or U2140 (N_2140,N_1332,N_1555);
nand U2141 (N_2141,N_1487,N_1298);
and U2142 (N_2142,N_1363,N_1791);
nor U2143 (N_2143,N_1721,N_1348);
and U2144 (N_2144,N_1323,N_1764);
or U2145 (N_2145,N_1313,N_1623);
and U2146 (N_2146,N_1272,N_1398);
xor U2147 (N_2147,N_1529,N_1262);
or U2148 (N_2148,N_1436,N_1357);
nand U2149 (N_2149,N_1605,N_1274);
nor U2150 (N_2150,N_1797,N_1695);
and U2151 (N_2151,N_1260,N_1721);
or U2152 (N_2152,N_1542,N_1567);
xnor U2153 (N_2153,N_1713,N_1237);
or U2154 (N_2154,N_1300,N_1770);
and U2155 (N_2155,N_1337,N_1379);
or U2156 (N_2156,N_1702,N_1200);
nor U2157 (N_2157,N_1348,N_1725);
and U2158 (N_2158,N_1745,N_1658);
xor U2159 (N_2159,N_1720,N_1431);
xor U2160 (N_2160,N_1485,N_1369);
xnor U2161 (N_2161,N_1383,N_1747);
and U2162 (N_2162,N_1373,N_1201);
nand U2163 (N_2163,N_1285,N_1346);
or U2164 (N_2164,N_1419,N_1240);
nor U2165 (N_2165,N_1764,N_1430);
nor U2166 (N_2166,N_1365,N_1223);
nand U2167 (N_2167,N_1777,N_1578);
and U2168 (N_2168,N_1432,N_1491);
or U2169 (N_2169,N_1721,N_1759);
xor U2170 (N_2170,N_1245,N_1318);
or U2171 (N_2171,N_1458,N_1606);
nand U2172 (N_2172,N_1287,N_1503);
nand U2173 (N_2173,N_1476,N_1363);
xnor U2174 (N_2174,N_1523,N_1258);
xnor U2175 (N_2175,N_1701,N_1263);
xnor U2176 (N_2176,N_1717,N_1403);
nand U2177 (N_2177,N_1353,N_1610);
xnor U2178 (N_2178,N_1379,N_1232);
and U2179 (N_2179,N_1641,N_1538);
and U2180 (N_2180,N_1630,N_1482);
nand U2181 (N_2181,N_1782,N_1727);
and U2182 (N_2182,N_1549,N_1514);
nor U2183 (N_2183,N_1261,N_1269);
or U2184 (N_2184,N_1283,N_1539);
nor U2185 (N_2185,N_1340,N_1482);
nor U2186 (N_2186,N_1741,N_1755);
and U2187 (N_2187,N_1597,N_1209);
nor U2188 (N_2188,N_1776,N_1200);
and U2189 (N_2189,N_1675,N_1558);
xnor U2190 (N_2190,N_1698,N_1349);
or U2191 (N_2191,N_1283,N_1203);
xor U2192 (N_2192,N_1288,N_1687);
nor U2193 (N_2193,N_1434,N_1726);
and U2194 (N_2194,N_1471,N_1427);
and U2195 (N_2195,N_1747,N_1422);
nor U2196 (N_2196,N_1603,N_1715);
xor U2197 (N_2197,N_1418,N_1301);
and U2198 (N_2198,N_1778,N_1232);
or U2199 (N_2199,N_1657,N_1234);
or U2200 (N_2200,N_1500,N_1620);
nor U2201 (N_2201,N_1736,N_1267);
xnor U2202 (N_2202,N_1299,N_1663);
or U2203 (N_2203,N_1288,N_1397);
and U2204 (N_2204,N_1607,N_1696);
and U2205 (N_2205,N_1545,N_1534);
and U2206 (N_2206,N_1670,N_1370);
and U2207 (N_2207,N_1492,N_1561);
nand U2208 (N_2208,N_1642,N_1277);
or U2209 (N_2209,N_1423,N_1549);
or U2210 (N_2210,N_1364,N_1298);
or U2211 (N_2211,N_1763,N_1383);
and U2212 (N_2212,N_1243,N_1631);
and U2213 (N_2213,N_1418,N_1591);
xor U2214 (N_2214,N_1425,N_1270);
or U2215 (N_2215,N_1767,N_1411);
nand U2216 (N_2216,N_1768,N_1306);
nand U2217 (N_2217,N_1272,N_1380);
and U2218 (N_2218,N_1267,N_1317);
nor U2219 (N_2219,N_1217,N_1571);
and U2220 (N_2220,N_1211,N_1681);
or U2221 (N_2221,N_1426,N_1569);
nor U2222 (N_2222,N_1314,N_1200);
and U2223 (N_2223,N_1201,N_1744);
and U2224 (N_2224,N_1444,N_1660);
and U2225 (N_2225,N_1526,N_1581);
nor U2226 (N_2226,N_1210,N_1653);
nand U2227 (N_2227,N_1785,N_1773);
or U2228 (N_2228,N_1706,N_1539);
nand U2229 (N_2229,N_1666,N_1209);
nand U2230 (N_2230,N_1492,N_1248);
nand U2231 (N_2231,N_1491,N_1279);
xor U2232 (N_2232,N_1331,N_1593);
or U2233 (N_2233,N_1509,N_1626);
nand U2234 (N_2234,N_1471,N_1568);
nand U2235 (N_2235,N_1344,N_1785);
nor U2236 (N_2236,N_1649,N_1251);
or U2237 (N_2237,N_1646,N_1606);
and U2238 (N_2238,N_1783,N_1624);
and U2239 (N_2239,N_1531,N_1698);
nand U2240 (N_2240,N_1709,N_1242);
or U2241 (N_2241,N_1393,N_1269);
and U2242 (N_2242,N_1243,N_1460);
or U2243 (N_2243,N_1630,N_1209);
and U2244 (N_2244,N_1434,N_1765);
or U2245 (N_2245,N_1255,N_1618);
nand U2246 (N_2246,N_1200,N_1292);
nor U2247 (N_2247,N_1345,N_1379);
and U2248 (N_2248,N_1489,N_1595);
nor U2249 (N_2249,N_1566,N_1697);
nand U2250 (N_2250,N_1322,N_1764);
and U2251 (N_2251,N_1679,N_1306);
xnor U2252 (N_2252,N_1351,N_1547);
xor U2253 (N_2253,N_1526,N_1594);
or U2254 (N_2254,N_1276,N_1729);
or U2255 (N_2255,N_1210,N_1655);
nor U2256 (N_2256,N_1657,N_1483);
xnor U2257 (N_2257,N_1201,N_1659);
and U2258 (N_2258,N_1448,N_1393);
nand U2259 (N_2259,N_1283,N_1603);
xnor U2260 (N_2260,N_1368,N_1304);
xor U2261 (N_2261,N_1358,N_1310);
nor U2262 (N_2262,N_1789,N_1327);
and U2263 (N_2263,N_1696,N_1772);
or U2264 (N_2264,N_1793,N_1512);
xor U2265 (N_2265,N_1323,N_1255);
and U2266 (N_2266,N_1461,N_1226);
nand U2267 (N_2267,N_1212,N_1685);
nand U2268 (N_2268,N_1312,N_1569);
or U2269 (N_2269,N_1699,N_1555);
nor U2270 (N_2270,N_1322,N_1230);
xor U2271 (N_2271,N_1288,N_1244);
and U2272 (N_2272,N_1248,N_1500);
nor U2273 (N_2273,N_1226,N_1793);
and U2274 (N_2274,N_1502,N_1533);
nor U2275 (N_2275,N_1276,N_1322);
or U2276 (N_2276,N_1673,N_1782);
xor U2277 (N_2277,N_1697,N_1661);
xnor U2278 (N_2278,N_1323,N_1760);
nor U2279 (N_2279,N_1254,N_1250);
xnor U2280 (N_2280,N_1702,N_1752);
nand U2281 (N_2281,N_1787,N_1457);
nand U2282 (N_2282,N_1430,N_1779);
nand U2283 (N_2283,N_1296,N_1554);
and U2284 (N_2284,N_1289,N_1273);
xnor U2285 (N_2285,N_1370,N_1434);
and U2286 (N_2286,N_1341,N_1459);
and U2287 (N_2287,N_1630,N_1530);
nand U2288 (N_2288,N_1633,N_1762);
nand U2289 (N_2289,N_1518,N_1233);
or U2290 (N_2290,N_1794,N_1664);
nand U2291 (N_2291,N_1225,N_1360);
or U2292 (N_2292,N_1650,N_1590);
nor U2293 (N_2293,N_1329,N_1770);
nor U2294 (N_2294,N_1720,N_1650);
or U2295 (N_2295,N_1474,N_1690);
nor U2296 (N_2296,N_1423,N_1756);
and U2297 (N_2297,N_1661,N_1200);
and U2298 (N_2298,N_1710,N_1315);
nand U2299 (N_2299,N_1256,N_1369);
or U2300 (N_2300,N_1281,N_1245);
nand U2301 (N_2301,N_1252,N_1327);
or U2302 (N_2302,N_1716,N_1628);
xor U2303 (N_2303,N_1642,N_1777);
or U2304 (N_2304,N_1304,N_1540);
or U2305 (N_2305,N_1702,N_1240);
or U2306 (N_2306,N_1607,N_1278);
nor U2307 (N_2307,N_1615,N_1262);
nand U2308 (N_2308,N_1400,N_1608);
or U2309 (N_2309,N_1304,N_1665);
or U2310 (N_2310,N_1660,N_1756);
and U2311 (N_2311,N_1262,N_1476);
or U2312 (N_2312,N_1657,N_1371);
xnor U2313 (N_2313,N_1592,N_1680);
xor U2314 (N_2314,N_1518,N_1319);
nor U2315 (N_2315,N_1516,N_1263);
and U2316 (N_2316,N_1764,N_1239);
and U2317 (N_2317,N_1248,N_1372);
and U2318 (N_2318,N_1518,N_1653);
nand U2319 (N_2319,N_1370,N_1368);
nor U2320 (N_2320,N_1531,N_1736);
and U2321 (N_2321,N_1559,N_1526);
nor U2322 (N_2322,N_1311,N_1610);
xnor U2323 (N_2323,N_1338,N_1454);
xor U2324 (N_2324,N_1277,N_1552);
or U2325 (N_2325,N_1336,N_1298);
and U2326 (N_2326,N_1454,N_1300);
nand U2327 (N_2327,N_1653,N_1555);
nand U2328 (N_2328,N_1543,N_1754);
nor U2329 (N_2329,N_1601,N_1582);
or U2330 (N_2330,N_1244,N_1405);
and U2331 (N_2331,N_1263,N_1739);
nor U2332 (N_2332,N_1495,N_1761);
nand U2333 (N_2333,N_1695,N_1264);
nand U2334 (N_2334,N_1383,N_1658);
xnor U2335 (N_2335,N_1763,N_1755);
xor U2336 (N_2336,N_1565,N_1367);
xnor U2337 (N_2337,N_1597,N_1747);
nand U2338 (N_2338,N_1248,N_1482);
nand U2339 (N_2339,N_1778,N_1433);
nor U2340 (N_2340,N_1528,N_1555);
nand U2341 (N_2341,N_1404,N_1580);
or U2342 (N_2342,N_1283,N_1418);
and U2343 (N_2343,N_1406,N_1428);
nand U2344 (N_2344,N_1591,N_1491);
nor U2345 (N_2345,N_1275,N_1250);
or U2346 (N_2346,N_1499,N_1202);
nor U2347 (N_2347,N_1514,N_1529);
or U2348 (N_2348,N_1765,N_1428);
nand U2349 (N_2349,N_1763,N_1285);
nand U2350 (N_2350,N_1266,N_1373);
nor U2351 (N_2351,N_1377,N_1337);
or U2352 (N_2352,N_1618,N_1422);
nand U2353 (N_2353,N_1300,N_1557);
nor U2354 (N_2354,N_1596,N_1298);
xor U2355 (N_2355,N_1724,N_1506);
nor U2356 (N_2356,N_1297,N_1520);
and U2357 (N_2357,N_1712,N_1724);
or U2358 (N_2358,N_1434,N_1226);
and U2359 (N_2359,N_1291,N_1311);
and U2360 (N_2360,N_1685,N_1299);
nand U2361 (N_2361,N_1680,N_1329);
and U2362 (N_2362,N_1331,N_1477);
xor U2363 (N_2363,N_1580,N_1702);
nor U2364 (N_2364,N_1686,N_1484);
nand U2365 (N_2365,N_1600,N_1323);
nand U2366 (N_2366,N_1568,N_1285);
xor U2367 (N_2367,N_1306,N_1605);
or U2368 (N_2368,N_1351,N_1609);
and U2369 (N_2369,N_1219,N_1660);
nand U2370 (N_2370,N_1519,N_1355);
and U2371 (N_2371,N_1459,N_1537);
or U2372 (N_2372,N_1786,N_1737);
or U2373 (N_2373,N_1430,N_1522);
or U2374 (N_2374,N_1220,N_1263);
and U2375 (N_2375,N_1243,N_1660);
or U2376 (N_2376,N_1546,N_1414);
xnor U2377 (N_2377,N_1582,N_1383);
nor U2378 (N_2378,N_1327,N_1560);
or U2379 (N_2379,N_1785,N_1677);
xor U2380 (N_2380,N_1726,N_1533);
and U2381 (N_2381,N_1760,N_1374);
nor U2382 (N_2382,N_1327,N_1540);
or U2383 (N_2383,N_1744,N_1417);
and U2384 (N_2384,N_1546,N_1607);
nor U2385 (N_2385,N_1356,N_1586);
and U2386 (N_2386,N_1514,N_1372);
xor U2387 (N_2387,N_1558,N_1350);
nor U2388 (N_2388,N_1662,N_1441);
xnor U2389 (N_2389,N_1407,N_1236);
nor U2390 (N_2390,N_1795,N_1637);
xor U2391 (N_2391,N_1739,N_1797);
or U2392 (N_2392,N_1316,N_1317);
and U2393 (N_2393,N_1578,N_1523);
and U2394 (N_2394,N_1564,N_1253);
or U2395 (N_2395,N_1768,N_1215);
nand U2396 (N_2396,N_1467,N_1450);
or U2397 (N_2397,N_1312,N_1740);
nand U2398 (N_2398,N_1679,N_1697);
or U2399 (N_2399,N_1733,N_1379);
or U2400 (N_2400,N_1801,N_2039);
and U2401 (N_2401,N_1919,N_2202);
nor U2402 (N_2402,N_1889,N_2393);
nand U2403 (N_2403,N_2106,N_2097);
nand U2404 (N_2404,N_2307,N_1968);
and U2405 (N_2405,N_2129,N_2142);
nor U2406 (N_2406,N_1806,N_1846);
nor U2407 (N_2407,N_1940,N_2086);
xnor U2408 (N_2408,N_2283,N_2174);
nand U2409 (N_2409,N_1861,N_2376);
nor U2410 (N_2410,N_2156,N_2210);
or U2411 (N_2411,N_1969,N_1820);
xnor U2412 (N_2412,N_2367,N_1850);
and U2413 (N_2413,N_1954,N_2115);
nor U2414 (N_2414,N_1922,N_1972);
and U2415 (N_2415,N_1992,N_1994);
and U2416 (N_2416,N_2343,N_1896);
nand U2417 (N_2417,N_2294,N_2073);
or U2418 (N_2418,N_2151,N_2193);
or U2419 (N_2419,N_1865,N_2235);
xor U2420 (N_2420,N_2325,N_2070);
nand U2421 (N_2421,N_2028,N_1811);
nor U2422 (N_2422,N_1895,N_1835);
xor U2423 (N_2423,N_2183,N_1942);
or U2424 (N_2424,N_2079,N_1989);
and U2425 (N_2425,N_1904,N_2279);
and U2426 (N_2426,N_2242,N_2113);
and U2427 (N_2427,N_2114,N_1862);
nor U2428 (N_2428,N_1819,N_1917);
or U2429 (N_2429,N_2365,N_2378);
nor U2430 (N_2430,N_1997,N_2253);
nor U2431 (N_2431,N_2065,N_2381);
nand U2432 (N_2432,N_2020,N_1856);
nand U2433 (N_2433,N_1946,N_1983);
nand U2434 (N_2434,N_2328,N_2177);
or U2435 (N_2435,N_2297,N_2096);
nor U2436 (N_2436,N_2132,N_2387);
nor U2437 (N_2437,N_1974,N_2329);
xor U2438 (N_2438,N_1805,N_2255);
and U2439 (N_2439,N_2000,N_1828);
and U2440 (N_2440,N_1934,N_1993);
xnor U2441 (N_2441,N_2184,N_2155);
nand U2442 (N_2442,N_1888,N_2230);
xnor U2443 (N_2443,N_1851,N_2111);
or U2444 (N_2444,N_2056,N_1981);
or U2445 (N_2445,N_1886,N_2293);
xor U2446 (N_2446,N_2214,N_2045);
xnor U2447 (N_2447,N_1990,N_2093);
and U2448 (N_2448,N_2379,N_1834);
nand U2449 (N_2449,N_2354,N_1925);
or U2450 (N_2450,N_1817,N_2200);
or U2451 (N_2451,N_2290,N_2352);
xnor U2452 (N_2452,N_2292,N_2076);
and U2453 (N_2453,N_1943,N_1843);
nand U2454 (N_2454,N_2391,N_2388);
and U2455 (N_2455,N_2148,N_2122);
xnor U2456 (N_2456,N_1823,N_2143);
nand U2457 (N_2457,N_2116,N_1840);
or U2458 (N_2458,N_2091,N_2336);
nand U2459 (N_2459,N_2057,N_2394);
and U2460 (N_2460,N_2171,N_2252);
xor U2461 (N_2461,N_2008,N_2134);
xor U2462 (N_2462,N_1881,N_2058);
and U2463 (N_2463,N_2326,N_2211);
nor U2464 (N_2464,N_1833,N_2263);
nand U2465 (N_2465,N_1814,N_2044);
xnor U2466 (N_2466,N_2135,N_1855);
nand U2467 (N_2467,N_2082,N_1824);
or U2468 (N_2468,N_2353,N_2147);
and U2469 (N_2469,N_2095,N_2011);
or U2470 (N_2470,N_2267,N_1908);
or U2471 (N_2471,N_1853,N_2346);
and U2472 (N_2472,N_2261,N_1953);
and U2473 (N_2473,N_1829,N_2078);
or U2474 (N_2474,N_1804,N_2306);
and U2475 (N_2475,N_1980,N_2153);
xor U2476 (N_2476,N_2108,N_2101);
and U2477 (N_2477,N_2052,N_1978);
or U2478 (N_2478,N_1952,N_1956);
xnor U2479 (N_2479,N_2257,N_2303);
nor U2480 (N_2480,N_2144,N_1818);
or U2481 (N_2481,N_2218,N_2075);
and U2482 (N_2482,N_2006,N_2339);
and U2483 (N_2483,N_1960,N_1914);
xor U2484 (N_2484,N_1988,N_2236);
or U2485 (N_2485,N_2180,N_1893);
or U2486 (N_2486,N_1808,N_1857);
nor U2487 (N_2487,N_2163,N_2334);
xnor U2488 (N_2488,N_1854,N_1955);
nor U2489 (N_2489,N_2201,N_2223);
nor U2490 (N_2490,N_2015,N_2187);
and U2491 (N_2491,N_2295,N_2398);
and U2492 (N_2492,N_2229,N_1945);
xnor U2493 (N_2493,N_1932,N_2060);
and U2494 (N_2494,N_1849,N_1991);
nor U2495 (N_2495,N_2068,N_1852);
nand U2496 (N_2496,N_2314,N_2222);
nor U2497 (N_2497,N_1891,N_2291);
nor U2498 (N_2498,N_2025,N_1867);
or U2499 (N_2499,N_1836,N_2085);
xnor U2500 (N_2500,N_2347,N_1938);
or U2501 (N_2501,N_2285,N_2231);
nor U2502 (N_2502,N_2001,N_1961);
nor U2503 (N_2503,N_1935,N_2190);
xor U2504 (N_2504,N_2166,N_1839);
nand U2505 (N_2505,N_1929,N_2186);
xor U2506 (N_2506,N_2102,N_2031);
nand U2507 (N_2507,N_2178,N_2162);
nand U2508 (N_2508,N_2004,N_2127);
nor U2509 (N_2509,N_2247,N_2043);
nand U2510 (N_2510,N_1926,N_2133);
xor U2511 (N_2511,N_2207,N_1903);
nor U2512 (N_2512,N_1967,N_2119);
nor U2513 (N_2513,N_2227,N_2337);
and U2514 (N_2514,N_1996,N_1913);
and U2515 (N_2515,N_2040,N_2141);
or U2516 (N_2516,N_2194,N_2249);
xor U2517 (N_2517,N_1832,N_2110);
nor U2518 (N_2518,N_1957,N_1918);
xnor U2519 (N_2519,N_2032,N_2172);
and U2520 (N_2520,N_2185,N_2240);
nor U2521 (N_2521,N_2107,N_2358);
nand U2522 (N_2522,N_2100,N_2021);
nand U2523 (N_2523,N_2118,N_2026);
or U2524 (N_2524,N_2164,N_2150);
xor U2525 (N_2525,N_1951,N_2383);
xor U2526 (N_2526,N_2029,N_2055);
and U2527 (N_2527,N_2274,N_2375);
nand U2528 (N_2528,N_1905,N_2286);
or U2529 (N_2529,N_1920,N_1830);
xor U2530 (N_2530,N_1979,N_1977);
or U2531 (N_2531,N_2179,N_2137);
nor U2532 (N_2532,N_2050,N_2089);
xor U2533 (N_2533,N_2212,N_2309);
xnor U2534 (N_2534,N_2321,N_1927);
or U2535 (N_2535,N_2136,N_2121);
nor U2536 (N_2536,N_2323,N_2077);
and U2537 (N_2537,N_2273,N_2298);
or U2538 (N_2538,N_2198,N_2239);
nor U2539 (N_2539,N_2226,N_1831);
and U2540 (N_2540,N_1890,N_1810);
and U2541 (N_2541,N_1860,N_1950);
xnor U2542 (N_2542,N_2251,N_1882);
nor U2543 (N_2543,N_2099,N_1984);
and U2544 (N_2544,N_2131,N_1916);
nand U2545 (N_2545,N_2259,N_2277);
nor U2546 (N_2546,N_2356,N_2188);
nand U2547 (N_2547,N_1872,N_2370);
and U2548 (N_2548,N_1877,N_1803);
or U2549 (N_2549,N_2244,N_2013);
and U2550 (N_2550,N_2002,N_2299);
and U2551 (N_2551,N_2120,N_1858);
and U2552 (N_2552,N_1887,N_1947);
or U2553 (N_2553,N_2012,N_2192);
xor U2554 (N_2554,N_1987,N_2300);
or U2555 (N_2555,N_2363,N_1902);
xor U2556 (N_2556,N_2359,N_1866);
xnor U2557 (N_2557,N_2302,N_2081);
or U2558 (N_2558,N_2167,N_1973);
and U2559 (N_2559,N_1826,N_2220);
and U2560 (N_2560,N_2175,N_1962);
xor U2561 (N_2561,N_1847,N_2335);
nor U2562 (N_2562,N_2382,N_1821);
nor U2563 (N_2563,N_2272,N_1848);
or U2564 (N_2564,N_2204,N_1875);
or U2565 (N_2565,N_2173,N_1901);
nand U2566 (N_2566,N_2250,N_1964);
nor U2567 (N_2567,N_1883,N_2313);
or U2568 (N_2568,N_1995,N_1939);
nor U2569 (N_2569,N_2003,N_2288);
nand U2570 (N_2570,N_1911,N_1982);
nand U2571 (N_2571,N_2237,N_2130);
nand U2572 (N_2572,N_2312,N_2117);
xor U2573 (N_2573,N_2366,N_2246);
xnor U2574 (N_2574,N_2084,N_1813);
or U2575 (N_2575,N_2215,N_2063);
xor U2576 (N_2576,N_1869,N_2189);
or U2577 (N_2577,N_2203,N_2351);
and U2578 (N_2578,N_2320,N_2152);
nand U2579 (N_2579,N_2361,N_2169);
nand U2580 (N_2580,N_1841,N_1959);
and U2581 (N_2581,N_2276,N_1970);
nand U2582 (N_2582,N_1870,N_2157);
nand U2583 (N_2583,N_1965,N_2331);
nand U2584 (N_2584,N_2260,N_2072);
and U2585 (N_2585,N_2199,N_2030);
and U2586 (N_2586,N_1915,N_1924);
xnor U2587 (N_2587,N_2158,N_2289);
xnor U2588 (N_2588,N_2281,N_1827);
or U2589 (N_2589,N_2344,N_2308);
or U2590 (N_2590,N_1985,N_2083);
nand U2591 (N_2591,N_2282,N_1937);
nor U2592 (N_2592,N_1936,N_2062);
and U2593 (N_2593,N_2245,N_2213);
xor U2594 (N_2594,N_2010,N_2348);
or U2595 (N_2595,N_2064,N_2338);
or U2596 (N_2596,N_1899,N_1859);
and U2597 (N_2597,N_2233,N_2191);
nor U2598 (N_2598,N_1873,N_2048);
or U2599 (N_2599,N_2305,N_2384);
nor U2600 (N_2600,N_1941,N_2268);
nor U2601 (N_2601,N_2316,N_2208);
or U2602 (N_2602,N_2311,N_2265);
and U2603 (N_2603,N_1878,N_2037);
and U2604 (N_2604,N_2080,N_2094);
nand U2605 (N_2605,N_2066,N_2053);
and U2606 (N_2606,N_2389,N_2105);
xnor U2607 (N_2607,N_2264,N_2269);
and U2608 (N_2608,N_1897,N_2266);
or U2609 (N_2609,N_2228,N_2278);
xor U2610 (N_2610,N_2146,N_2019);
and U2611 (N_2611,N_2034,N_2168);
or U2612 (N_2612,N_2350,N_2332);
nand U2613 (N_2613,N_1930,N_1910);
or U2614 (N_2614,N_1907,N_1837);
nor U2615 (N_2615,N_2125,N_2392);
nand U2616 (N_2616,N_2195,N_1909);
nand U2617 (N_2617,N_2275,N_2154);
nand U2618 (N_2618,N_1971,N_2395);
nand U2619 (N_2619,N_1963,N_2219);
nand U2620 (N_2620,N_1809,N_2176);
xor U2621 (N_2621,N_1933,N_2042);
nand U2622 (N_2622,N_2139,N_2197);
nand U2623 (N_2623,N_2254,N_1825);
and U2624 (N_2624,N_1958,N_2377);
and U2625 (N_2625,N_2364,N_1898);
and U2626 (N_2626,N_1966,N_1892);
and U2627 (N_2627,N_2380,N_1906);
and U2628 (N_2628,N_2138,N_2046);
nand U2629 (N_2629,N_2374,N_2196);
nor U2630 (N_2630,N_1949,N_1864);
and U2631 (N_2631,N_2074,N_2386);
or U2632 (N_2632,N_2007,N_2181);
xnor U2633 (N_2633,N_1871,N_2225);
xnor U2634 (N_2634,N_2161,N_2221);
or U2635 (N_2635,N_2396,N_2360);
nand U2636 (N_2636,N_2022,N_2373);
nand U2637 (N_2637,N_1921,N_2310);
or U2638 (N_2638,N_2315,N_2123);
nand U2639 (N_2639,N_1838,N_2397);
and U2640 (N_2640,N_2232,N_2256);
xor U2641 (N_2641,N_1885,N_2069);
nand U2642 (N_2642,N_1998,N_2206);
and U2643 (N_2643,N_2238,N_2126);
nand U2644 (N_2644,N_2330,N_2087);
and U2645 (N_2645,N_2038,N_2271);
and U2646 (N_2646,N_1868,N_1876);
or U2647 (N_2647,N_1822,N_1874);
nor U2648 (N_2648,N_2033,N_2041);
xnor U2649 (N_2649,N_2009,N_1863);
xor U2650 (N_2650,N_2371,N_2390);
xnor U2651 (N_2651,N_2149,N_1802);
and U2652 (N_2652,N_2355,N_2124);
and U2653 (N_2653,N_1880,N_2287);
nor U2654 (N_2654,N_2304,N_2243);
xnor U2655 (N_2655,N_2324,N_2090);
or U2656 (N_2656,N_2322,N_2224);
xor U2657 (N_2657,N_2160,N_2036);
nor U2658 (N_2658,N_2047,N_2284);
xor U2659 (N_2659,N_1912,N_2005);
or U2660 (N_2660,N_2296,N_2399);
xnor U2661 (N_2661,N_2241,N_2280);
or U2662 (N_2662,N_1842,N_2362);
or U2663 (N_2663,N_2349,N_1815);
or U2664 (N_2664,N_2165,N_2112);
or U2665 (N_2665,N_2327,N_1894);
nor U2666 (N_2666,N_2014,N_2301);
nand U2667 (N_2667,N_2018,N_2051);
xor U2668 (N_2668,N_1928,N_2049);
and U2669 (N_2669,N_2061,N_2217);
nor U2670 (N_2670,N_2103,N_1879);
xnor U2671 (N_2671,N_2067,N_2023);
or U2672 (N_2672,N_1923,N_2270);
nand U2673 (N_2673,N_2248,N_2017);
and U2674 (N_2674,N_2109,N_1931);
nor U2675 (N_2675,N_1807,N_2092);
and U2676 (N_2676,N_2140,N_2319);
xor U2677 (N_2677,N_1975,N_1884);
nand U2678 (N_2678,N_2385,N_2128);
xor U2679 (N_2679,N_2357,N_2098);
xor U2680 (N_2680,N_1986,N_2318);
nor U2681 (N_2681,N_2054,N_1948);
or U2682 (N_2682,N_2024,N_2372);
or U2683 (N_2683,N_2368,N_2262);
and U2684 (N_2684,N_1900,N_2170);
xnor U2685 (N_2685,N_2205,N_1816);
nand U2686 (N_2686,N_2340,N_1845);
nor U2687 (N_2687,N_2035,N_2234);
xor U2688 (N_2688,N_1812,N_1999);
xor U2689 (N_2689,N_1844,N_2342);
xnor U2690 (N_2690,N_2345,N_2182);
xor U2691 (N_2691,N_1944,N_2333);
and U2692 (N_2692,N_2369,N_1800);
xnor U2693 (N_2693,N_2027,N_2145);
nand U2694 (N_2694,N_2071,N_2258);
nor U2695 (N_2695,N_1976,N_2159);
or U2696 (N_2696,N_2104,N_2088);
and U2697 (N_2697,N_2016,N_2341);
nor U2698 (N_2698,N_2317,N_2059);
nand U2699 (N_2699,N_2209,N_2216);
nand U2700 (N_2700,N_2105,N_2316);
nor U2701 (N_2701,N_2155,N_1846);
nand U2702 (N_2702,N_2016,N_2070);
nor U2703 (N_2703,N_2168,N_2067);
or U2704 (N_2704,N_2111,N_2301);
and U2705 (N_2705,N_2349,N_1997);
and U2706 (N_2706,N_2379,N_1966);
or U2707 (N_2707,N_2330,N_2077);
nand U2708 (N_2708,N_2036,N_2219);
or U2709 (N_2709,N_1926,N_2177);
nor U2710 (N_2710,N_2392,N_2244);
or U2711 (N_2711,N_2048,N_2070);
nand U2712 (N_2712,N_2028,N_2352);
or U2713 (N_2713,N_1803,N_1843);
nand U2714 (N_2714,N_1817,N_2041);
nand U2715 (N_2715,N_1924,N_2108);
and U2716 (N_2716,N_1814,N_2036);
nor U2717 (N_2717,N_1980,N_2279);
nor U2718 (N_2718,N_2258,N_2291);
xor U2719 (N_2719,N_2054,N_2376);
or U2720 (N_2720,N_1833,N_2341);
nor U2721 (N_2721,N_1854,N_2337);
nor U2722 (N_2722,N_1850,N_2118);
or U2723 (N_2723,N_2243,N_1878);
xor U2724 (N_2724,N_2329,N_2234);
and U2725 (N_2725,N_1805,N_2351);
and U2726 (N_2726,N_2111,N_2399);
or U2727 (N_2727,N_2286,N_2251);
xnor U2728 (N_2728,N_2210,N_1991);
nor U2729 (N_2729,N_1909,N_2029);
and U2730 (N_2730,N_1889,N_2180);
nor U2731 (N_2731,N_1974,N_2282);
or U2732 (N_2732,N_2314,N_2165);
nand U2733 (N_2733,N_2032,N_2025);
and U2734 (N_2734,N_2042,N_2268);
xor U2735 (N_2735,N_1889,N_1853);
xor U2736 (N_2736,N_2044,N_1969);
and U2737 (N_2737,N_1872,N_2109);
and U2738 (N_2738,N_2298,N_1957);
nand U2739 (N_2739,N_2072,N_2077);
xor U2740 (N_2740,N_2118,N_2255);
nor U2741 (N_2741,N_1912,N_2345);
or U2742 (N_2742,N_2395,N_2376);
nand U2743 (N_2743,N_2341,N_2132);
xnor U2744 (N_2744,N_2049,N_2363);
or U2745 (N_2745,N_2363,N_1827);
nor U2746 (N_2746,N_2305,N_2127);
nand U2747 (N_2747,N_2230,N_2233);
xor U2748 (N_2748,N_2307,N_2106);
nor U2749 (N_2749,N_2087,N_2255);
and U2750 (N_2750,N_1871,N_2076);
nand U2751 (N_2751,N_1859,N_2084);
xnor U2752 (N_2752,N_2325,N_2374);
or U2753 (N_2753,N_2000,N_2164);
nor U2754 (N_2754,N_2108,N_2201);
and U2755 (N_2755,N_1911,N_2069);
nor U2756 (N_2756,N_2113,N_1948);
nor U2757 (N_2757,N_2102,N_1866);
nor U2758 (N_2758,N_1822,N_2340);
nor U2759 (N_2759,N_2071,N_2395);
xnor U2760 (N_2760,N_2284,N_2369);
xor U2761 (N_2761,N_2174,N_2226);
xnor U2762 (N_2762,N_2287,N_1815);
nor U2763 (N_2763,N_2213,N_2143);
xnor U2764 (N_2764,N_1810,N_2043);
xnor U2765 (N_2765,N_2031,N_2398);
xor U2766 (N_2766,N_1928,N_1894);
or U2767 (N_2767,N_1939,N_1819);
nand U2768 (N_2768,N_2070,N_2103);
nand U2769 (N_2769,N_2340,N_2209);
nand U2770 (N_2770,N_2381,N_1972);
nand U2771 (N_2771,N_1871,N_2182);
xor U2772 (N_2772,N_2020,N_2317);
nand U2773 (N_2773,N_1917,N_2214);
or U2774 (N_2774,N_2345,N_2375);
nand U2775 (N_2775,N_2391,N_2028);
nor U2776 (N_2776,N_1877,N_2320);
nand U2777 (N_2777,N_2050,N_2362);
xor U2778 (N_2778,N_2350,N_1899);
nand U2779 (N_2779,N_2364,N_1810);
nor U2780 (N_2780,N_2337,N_2050);
nand U2781 (N_2781,N_1985,N_2016);
nand U2782 (N_2782,N_2211,N_2008);
nor U2783 (N_2783,N_2080,N_2273);
nand U2784 (N_2784,N_2286,N_2347);
nand U2785 (N_2785,N_2282,N_2120);
xor U2786 (N_2786,N_2147,N_2120);
xor U2787 (N_2787,N_2099,N_2017);
and U2788 (N_2788,N_1825,N_1836);
xor U2789 (N_2789,N_1815,N_2282);
and U2790 (N_2790,N_2238,N_2267);
xnor U2791 (N_2791,N_1905,N_1998);
nor U2792 (N_2792,N_2173,N_2156);
nand U2793 (N_2793,N_2172,N_1963);
nand U2794 (N_2794,N_2084,N_2253);
xnor U2795 (N_2795,N_2033,N_2109);
or U2796 (N_2796,N_1838,N_2166);
and U2797 (N_2797,N_2044,N_2380);
or U2798 (N_2798,N_2168,N_2236);
nor U2799 (N_2799,N_1933,N_1956);
nor U2800 (N_2800,N_2114,N_1961);
nor U2801 (N_2801,N_1860,N_2329);
nor U2802 (N_2802,N_2134,N_2022);
nor U2803 (N_2803,N_2025,N_2084);
or U2804 (N_2804,N_1974,N_1945);
nor U2805 (N_2805,N_2344,N_1912);
xnor U2806 (N_2806,N_2047,N_2161);
nand U2807 (N_2807,N_2280,N_1884);
xor U2808 (N_2808,N_2345,N_2171);
nand U2809 (N_2809,N_2358,N_2207);
and U2810 (N_2810,N_1803,N_2100);
nand U2811 (N_2811,N_1988,N_1858);
xnor U2812 (N_2812,N_1860,N_1925);
nand U2813 (N_2813,N_1812,N_2214);
and U2814 (N_2814,N_2166,N_2224);
and U2815 (N_2815,N_2361,N_2168);
xor U2816 (N_2816,N_2353,N_2104);
xor U2817 (N_2817,N_1901,N_1985);
or U2818 (N_2818,N_2022,N_1887);
nor U2819 (N_2819,N_2145,N_2032);
xnor U2820 (N_2820,N_1873,N_1966);
nand U2821 (N_2821,N_2356,N_2375);
nand U2822 (N_2822,N_1929,N_2116);
xnor U2823 (N_2823,N_2271,N_1820);
nor U2824 (N_2824,N_2050,N_1997);
and U2825 (N_2825,N_2008,N_1877);
or U2826 (N_2826,N_2099,N_2292);
nand U2827 (N_2827,N_1816,N_1881);
nor U2828 (N_2828,N_2292,N_2200);
xnor U2829 (N_2829,N_2358,N_2317);
nor U2830 (N_2830,N_2249,N_2373);
nor U2831 (N_2831,N_2346,N_2096);
nor U2832 (N_2832,N_1837,N_1969);
xnor U2833 (N_2833,N_1828,N_1805);
nand U2834 (N_2834,N_1822,N_1958);
nor U2835 (N_2835,N_1924,N_2315);
nor U2836 (N_2836,N_1983,N_1896);
xor U2837 (N_2837,N_1992,N_2122);
or U2838 (N_2838,N_2396,N_1901);
or U2839 (N_2839,N_2339,N_1992);
nor U2840 (N_2840,N_1816,N_2316);
xor U2841 (N_2841,N_1965,N_1980);
nor U2842 (N_2842,N_2318,N_1838);
xor U2843 (N_2843,N_2368,N_2163);
xnor U2844 (N_2844,N_1876,N_1933);
xor U2845 (N_2845,N_1996,N_2231);
xnor U2846 (N_2846,N_2216,N_2114);
or U2847 (N_2847,N_2123,N_2227);
xnor U2848 (N_2848,N_2136,N_2069);
xnor U2849 (N_2849,N_2085,N_2306);
or U2850 (N_2850,N_2067,N_2002);
xnor U2851 (N_2851,N_2103,N_2056);
xnor U2852 (N_2852,N_2268,N_1819);
xor U2853 (N_2853,N_1865,N_2055);
xnor U2854 (N_2854,N_2040,N_2337);
nor U2855 (N_2855,N_2092,N_1869);
or U2856 (N_2856,N_2365,N_2359);
or U2857 (N_2857,N_2010,N_1918);
and U2858 (N_2858,N_2143,N_2343);
nor U2859 (N_2859,N_2215,N_2109);
and U2860 (N_2860,N_2175,N_2320);
nor U2861 (N_2861,N_1942,N_2186);
nand U2862 (N_2862,N_1852,N_2397);
or U2863 (N_2863,N_1821,N_1938);
or U2864 (N_2864,N_2228,N_2355);
xnor U2865 (N_2865,N_1942,N_2145);
nand U2866 (N_2866,N_2381,N_2372);
and U2867 (N_2867,N_2113,N_2069);
or U2868 (N_2868,N_2173,N_2335);
or U2869 (N_2869,N_1825,N_2380);
nor U2870 (N_2870,N_2296,N_2363);
nor U2871 (N_2871,N_2203,N_1902);
nand U2872 (N_2872,N_2141,N_1928);
nand U2873 (N_2873,N_2338,N_2013);
xnor U2874 (N_2874,N_2030,N_1852);
nand U2875 (N_2875,N_2319,N_2352);
xor U2876 (N_2876,N_2240,N_1800);
xor U2877 (N_2877,N_2147,N_2221);
nor U2878 (N_2878,N_2000,N_1943);
xor U2879 (N_2879,N_1802,N_2077);
nand U2880 (N_2880,N_2305,N_2273);
nor U2881 (N_2881,N_1854,N_2313);
or U2882 (N_2882,N_2076,N_2065);
nor U2883 (N_2883,N_1999,N_2175);
xnor U2884 (N_2884,N_1805,N_2304);
nor U2885 (N_2885,N_2213,N_2088);
or U2886 (N_2886,N_2294,N_2276);
xor U2887 (N_2887,N_2233,N_2225);
xnor U2888 (N_2888,N_2072,N_1850);
nand U2889 (N_2889,N_2396,N_2282);
or U2890 (N_2890,N_2292,N_2396);
or U2891 (N_2891,N_2397,N_2078);
nand U2892 (N_2892,N_1917,N_1990);
xor U2893 (N_2893,N_2135,N_1872);
and U2894 (N_2894,N_2297,N_1806);
xor U2895 (N_2895,N_2219,N_2334);
and U2896 (N_2896,N_2316,N_2102);
nor U2897 (N_2897,N_1931,N_2388);
and U2898 (N_2898,N_2032,N_2048);
nor U2899 (N_2899,N_1965,N_2350);
and U2900 (N_2900,N_2119,N_2236);
and U2901 (N_2901,N_2081,N_2377);
nand U2902 (N_2902,N_1920,N_2309);
and U2903 (N_2903,N_2272,N_1835);
or U2904 (N_2904,N_1911,N_2205);
xnor U2905 (N_2905,N_2232,N_1981);
nor U2906 (N_2906,N_2009,N_2212);
and U2907 (N_2907,N_1900,N_1983);
nand U2908 (N_2908,N_1931,N_1868);
xor U2909 (N_2909,N_2137,N_1845);
and U2910 (N_2910,N_2220,N_2028);
nor U2911 (N_2911,N_1988,N_1955);
nor U2912 (N_2912,N_2080,N_2145);
nor U2913 (N_2913,N_2252,N_1875);
xor U2914 (N_2914,N_2312,N_2002);
nor U2915 (N_2915,N_1855,N_1947);
nor U2916 (N_2916,N_1853,N_1939);
and U2917 (N_2917,N_2236,N_1902);
nand U2918 (N_2918,N_1885,N_2042);
nand U2919 (N_2919,N_2218,N_2244);
nor U2920 (N_2920,N_2009,N_2251);
nor U2921 (N_2921,N_1919,N_2170);
xor U2922 (N_2922,N_2139,N_1889);
nand U2923 (N_2923,N_1968,N_2376);
nand U2924 (N_2924,N_2339,N_2030);
nand U2925 (N_2925,N_2365,N_2239);
xnor U2926 (N_2926,N_2027,N_1892);
nand U2927 (N_2927,N_2156,N_2032);
xnor U2928 (N_2928,N_1837,N_2006);
or U2929 (N_2929,N_2390,N_2091);
or U2930 (N_2930,N_2173,N_2048);
nor U2931 (N_2931,N_1884,N_2308);
or U2932 (N_2932,N_2254,N_2014);
or U2933 (N_2933,N_1951,N_2050);
nand U2934 (N_2934,N_2127,N_2196);
nor U2935 (N_2935,N_2330,N_2073);
and U2936 (N_2936,N_1875,N_1854);
xnor U2937 (N_2937,N_1983,N_2179);
xnor U2938 (N_2938,N_2113,N_2323);
and U2939 (N_2939,N_2296,N_2227);
nor U2940 (N_2940,N_2111,N_1958);
xor U2941 (N_2941,N_1939,N_2334);
and U2942 (N_2942,N_1968,N_2025);
nand U2943 (N_2943,N_2190,N_1831);
or U2944 (N_2944,N_2270,N_2126);
nor U2945 (N_2945,N_2030,N_1999);
xnor U2946 (N_2946,N_1866,N_2210);
nand U2947 (N_2947,N_1908,N_2341);
and U2948 (N_2948,N_2140,N_2387);
and U2949 (N_2949,N_2038,N_1873);
or U2950 (N_2950,N_2217,N_1951);
and U2951 (N_2951,N_2290,N_2347);
nor U2952 (N_2952,N_1991,N_1803);
or U2953 (N_2953,N_1801,N_2014);
nor U2954 (N_2954,N_2108,N_2235);
or U2955 (N_2955,N_1856,N_2321);
nand U2956 (N_2956,N_2341,N_1987);
nor U2957 (N_2957,N_2234,N_2278);
or U2958 (N_2958,N_2020,N_1893);
nand U2959 (N_2959,N_1853,N_2093);
xor U2960 (N_2960,N_1927,N_2031);
or U2961 (N_2961,N_2171,N_2360);
and U2962 (N_2962,N_1911,N_2306);
and U2963 (N_2963,N_1825,N_1906);
xnor U2964 (N_2964,N_2210,N_1846);
or U2965 (N_2965,N_2138,N_1945);
xnor U2966 (N_2966,N_2359,N_1942);
and U2967 (N_2967,N_2128,N_1876);
nand U2968 (N_2968,N_2092,N_2161);
or U2969 (N_2969,N_1838,N_2099);
and U2970 (N_2970,N_1968,N_2292);
nor U2971 (N_2971,N_2086,N_2350);
and U2972 (N_2972,N_2102,N_2069);
or U2973 (N_2973,N_2313,N_2344);
nand U2974 (N_2974,N_1879,N_2053);
nor U2975 (N_2975,N_1858,N_1996);
nand U2976 (N_2976,N_2090,N_1897);
xnor U2977 (N_2977,N_2164,N_2065);
nor U2978 (N_2978,N_2231,N_1828);
and U2979 (N_2979,N_1866,N_1879);
xnor U2980 (N_2980,N_2139,N_2187);
xnor U2981 (N_2981,N_1843,N_2341);
xor U2982 (N_2982,N_1841,N_1869);
nand U2983 (N_2983,N_2350,N_1981);
or U2984 (N_2984,N_2175,N_2010);
nand U2985 (N_2985,N_1991,N_2171);
and U2986 (N_2986,N_1818,N_2284);
xor U2987 (N_2987,N_1994,N_2355);
nand U2988 (N_2988,N_2323,N_1868);
or U2989 (N_2989,N_2193,N_2098);
or U2990 (N_2990,N_2130,N_2132);
nand U2991 (N_2991,N_2119,N_2303);
nand U2992 (N_2992,N_2304,N_2062);
xor U2993 (N_2993,N_1800,N_2006);
xor U2994 (N_2994,N_2182,N_1868);
or U2995 (N_2995,N_2356,N_1833);
nand U2996 (N_2996,N_2093,N_2179);
nor U2997 (N_2997,N_1978,N_1982);
and U2998 (N_2998,N_2238,N_1829);
and U2999 (N_2999,N_1841,N_2061);
or UO_0 (O_0,N_2430,N_2731);
or UO_1 (O_1,N_2441,N_2432);
nor UO_2 (O_2,N_2952,N_2772);
nor UO_3 (O_3,N_2973,N_2549);
and UO_4 (O_4,N_2898,N_2443);
nand UO_5 (O_5,N_2956,N_2459);
or UO_6 (O_6,N_2594,N_2796);
or UO_7 (O_7,N_2737,N_2483);
and UO_8 (O_8,N_2510,N_2677);
or UO_9 (O_9,N_2636,N_2783);
nand UO_10 (O_10,N_2654,N_2929);
nand UO_11 (O_11,N_2596,N_2774);
xnor UO_12 (O_12,N_2902,N_2975);
nand UO_13 (O_13,N_2908,N_2825);
nor UO_14 (O_14,N_2423,N_2757);
or UO_15 (O_15,N_2684,N_2662);
nor UO_16 (O_16,N_2980,N_2778);
or UO_17 (O_17,N_2450,N_2509);
nor UO_18 (O_18,N_2831,N_2569);
nor UO_19 (O_19,N_2475,N_2574);
and UO_20 (O_20,N_2840,N_2505);
nor UO_21 (O_21,N_2889,N_2890);
nand UO_22 (O_22,N_2528,N_2775);
xnor UO_23 (O_23,N_2713,N_2703);
xnor UO_24 (O_24,N_2769,N_2940);
or UO_25 (O_25,N_2407,N_2927);
or UO_26 (O_26,N_2631,N_2962);
or UO_27 (O_27,N_2697,N_2640);
xor UO_28 (O_28,N_2958,N_2656);
or UO_29 (O_29,N_2595,N_2601);
xnor UO_30 (O_30,N_2708,N_2492);
nand UO_31 (O_31,N_2478,N_2622);
nand UO_32 (O_32,N_2879,N_2758);
and UO_33 (O_33,N_2982,N_2700);
or UO_34 (O_34,N_2672,N_2591);
nand UO_35 (O_35,N_2481,N_2759);
or UO_36 (O_36,N_2981,N_2884);
and UO_37 (O_37,N_2585,N_2638);
nor UO_38 (O_38,N_2909,N_2985);
nand UO_39 (O_39,N_2466,N_2824);
nand UO_40 (O_40,N_2867,N_2634);
or UO_41 (O_41,N_2474,N_2479);
and UO_42 (O_42,N_2959,N_2870);
nand UO_43 (O_43,N_2438,N_2765);
nor UO_44 (O_44,N_2789,N_2935);
xnor UO_45 (O_45,N_2925,N_2923);
and UO_46 (O_46,N_2788,N_2987);
and UO_47 (O_47,N_2428,N_2724);
or UO_48 (O_48,N_2696,N_2426);
and UO_49 (O_49,N_2480,N_2782);
nand UO_50 (O_50,N_2715,N_2946);
and UO_51 (O_51,N_2668,N_2624);
nor UO_52 (O_52,N_2660,N_2705);
and UO_53 (O_53,N_2694,N_2527);
and UO_54 (O_54,N_2750,N_2681);
and UO_55 (O_55,N_2687,N_2873);
nand UO_56 (O_56,N_2515,N_2730);
nor UO_57 (O_57,N_2887,N_2605);
and UO_58 (O_58,N_2673,N_2652);
nand UO_59 (O_59,N_2699,N_2635);
nand UO_60 (O_60,N_2858,N_2588);
nand UO_61 (O_61,N_2462,N_2473);
nor UO_62 (O_62,N_2749,N_2691);
or UO_63 (O_63,N_2553,N_2922);
and UO_64 (O_64,N_2616,N_2732);
and UO_65 (O_65,N_2842,N_2983);
nor UO_66 (O_66,N_2921,N_2989);
and UO_67 (O_67,N_2457,N_2698);
nor UO_68 (O_68,N_2828,N_2690);
xnor UO_69 (O_69,N_2495,N_2997);
xor UO_70 (O_70,N_2550,N_2501);
nor UO_71 (O_71,N_2802,N_2791);
and UO_72 (O_72,N_2875,N_2496);
xor UO_73 (O_73,N_2819,N_2888);
and UO_74 (O_74,N_2785,N_2518);
nor UO_75 (O_75,N_2627,N_2633);
nor UO_76 (O_76,N_2829,N_2904);
nor UO_77 (O_77,N_2598,N_2614);
or UO_78 (O_78,N_2880,N_2512);
and UO_79 (O_79,N_2854,N_2630);
nor UO_80 (O_80,N_2714,N_2972);
xnor UO_81 (O_81,N_2951,N_2948);
nor UO_82 (O_82,N_2744,N_2590);
nor UO_83 (O_83,N_2786,N_2548);
or UO_84 (O_84,N_2811,N_2773);
or UO_85 (O_85,N_2701,N_2801);
nand UO_86 (O_86,N_2628,N_2823);
nor UO_87 (O_87,N_2968,N_2470);
or UO_88 (O_88,N_2816,N_2963);
and UO_89 (O_89,N_2599,N_2657);
nor UO_90 (O_90,N_2612,N_2991);
and UO_91 (O_91,N_2451,N_2799);
nand UO_92 (O_92,N_2860,N_2565);
nor UO_93 (O_93,N_2545,N_2666);
nand UO_94 (O_94,N_2593,N_2996);
or UO_95 (O_95,N_2736,N_2878);
xor UO_96 (O_96,N_2682,N_2709);
and UO_97 (O_97,N_2874,N_2945);
nor UO_98 (O_98,N_2859,N_2846);
nor UO_99 (O_99,N_2755,N_2572);
xnor UO_100 (O_100,N_2544,N_2942);
xor UO_101 (O_101,N_2852,N_2669);
nor UO_102 (O_102,N_2655,N_2770);
xor UO_103 (O_103,N_2833,N_2937);
nand UO_104 (O_104,N_2827,N_2524);
xor UO_105 (O_105,N_2538,N_2924);
or UO_106 (O_106,N_2917,N_2446);
nor UO_107 (O_107,N_2582,N_2517);
or UO_108 (O_108,N_2822,N_2830);
or UO_109 (O_109,N_2651,N_2914);
nor UO_110 (O_110,N_2558,N_2427);
nand UO_111 (O_111,N_2579,N_2583);
or UO_112 (O_112,N_2894,N_2787);
nand UO_113 (O_113,N_2797,N_2485);
xnor UO_114 (O_114,N_2837,N_2866);
or UO_115 (O_115,N_2821,N_2836);
or UO_116 (O_116,N_2847,N_2747);
and UO_117 (O_117,N_2568,N_2776);
nand UO_118 (O_118,N_2621,N_2961);
and UO_119 (O_119,N_2477,N_2977);
nor UO_120 (O_120,N_2564,N_2882);
nor UO_121 (O_121,N_2767,N_2892);
nand UO_122 (O_122,N_2900,N_2577);
nand UO_123 (O_123,N_2853,N_2920);
nand UO_124 (O_124,N_2559,N_2692);
xnor UO_125 (O_125,N_2670,N_2695);
xnor UO_126 (O_126,N_2625,N_2575);
nand UO_127 (O_127,N_2978,N_2536);
nand UO_128 (O_128,N_2886,N_2618);
nor UO_129 (O_129,N_2805,N_2406);
nand UO_130 (O_130,N_2704,N_2442);
nor UO_131 (O_131,N_2916,N_2587);
and UO_132 (O_132,N_2453,N_2606);
nand UO_133 (O_133,N_2994,N_2974);
xnor UO_134 (O_134,N_2885,N_2905);
nor UO_135 (O_135,N_2431,N_2832);
nand UO_136 (O_136,N_2663,N_2611);
nor UO_137 (O_137,N_2642,N_2679);
and UO_138 (O_138,N_2447,N_2607);
nand UO_139 (O_139,N_2800,N_2436);
or UO_140 (O_140,N_2756,N_2792);
or UO_141 (O_141,N_2910,N_2733);
nor UO_142 (O_142,N_2502,N_2530);
xnor UO_143 (O_143,N_2803,N_2561);
and UO_144 (O_144,N_2813,N_2979);
and UO_145 (O_145,N_2895,N_2762);
nor UO_146 (O_146,N_2838,N_2851);
nor UO_147 (O_147,N_2597,N_2417);
or UO_148 (O_148,N_2938,N_2665);
and UO_149 (O_149,N_2600,N_2400);
xnor UO_150 (O_150,N_2988,N_2468);
nand UO_151 (O_151,N_2581,N_2727);
nand UO_152 (O_152,N_2661,N_2723);
nor UO_153 (O_153,N_2926,N_2413);
nand UO_154 (O_154,N_2603,N_2484);
xnor UO_155 (O_155,N_2650,N_2415);
xor UO_156 (O_156,N_2472,N_2465);
or UO_157 (O_157,N_2648,N_2540);
or UO_158 (O_158,N_2418,N_2683);
and UO_159 (O_159,N_2452,N_2491);
xor UO_160 (O_160,N_2421,N_2464);
nor UO_161 (O_161,N_2467,N_2763);
xor UO_162 (O_162,N_2856,N_2516);
xnor UO_163 (O_163,N_2520,N_2716);
and UO_164 (O_164,N_2967,N_2969);
and UO_165 (O_165,N_2779,N_2410);
nor UO_166 (O_166,N_2493,N_2711);
and UO_167 (O_167,N_2918,N_2444);
xor UO_168 (O_168,N_2941,N_2845);
or UO_169 (O_169,N_2498,N_2720);
xor UO_170 (O_170,N_2734,N_2425);
nand UO_171 (O_171,N_2891,N_2604);
nor UO_172 (O_172,N_2643,N_2735);
and UO_173 (O_173,N_2497,N_2482);
or UO_174 (O_174,N_2403,N_2608);
nor UO_175 (O_175,N_2531,N_2993);
nor UO_176 (O_176,N_2613,N_2793);
nor UO_177 (O_177,N_2984,N_2500);
nand UO_178 (O_178,N_2881,N_2998);
or UO_179 (O_179,N_2463,N_2448);
nor UO_180 (O_180,N_2646,N_2855);
or UO_181 (O_181,N_2688,N_2615);
nand UO_182 (O_182,N_2551,N_2740);
or UO_183 (O_183,N_2976,N_2839);
or UO_184 (O_184,N_2843,N_2903);
or UO_185 (O_185,N_2610,N_2434);
and UO_186 (O_186,N_2489,N_2999);
or UO_187 (O_187,N_2835,N_2667);
or UO_188 (O_188,N_2626,N_2990);
nand UO_189 (O_189,N_2766,N_2543);
nor UO_190 (O_190,N_2754,N_2573);
and UO_191 (O_191,N_2523,N_2966);
nand UO_192 (O_192,N_2445,N_2686);
nand UO_193 (O_193,N_2815,N_2764);
and UO_194 (O_194,N_2455,N_2566);
nor UO_195 (O_195,N_2812,N_2893);
or UO_196 (O_196,N_2623,N_2718);
nand UO_197 (O_197,N_2934,N_2586);
nor UO_198 (O_198,N_2671,N_2817);
xor UO_199 (O_199,N_2440,N_2419);
xnor UO_200 (O_200,N_2850,N_2637);
nor UO_201 (O_201,N_2865,N_2971);
nor UO_202 (O_202,N_2741,N_2576);
nand UO_203 (O_203,N_2809,N_2899);
nor UO_204 (O_204,N_2471,N_2957);
or UO_205 (O_205,N_2487,N_2871);
and UO_206 (O_206,N_2726,N_2943);
nor UO_207 (O_207,N_2689,N_2659);
nand UO_208 (O_208,N_2913,N_2532);
xnor UO_209 (O_209,N_2554,N_2702);
or UO_210 (O_210,N_2883,N_2454);
nand UO_211 (O_211,N_2584,N_2546);
and UO_212 (O_212,N_2869,N_2710);
nor UO_213 (O_213,N_2411,N_2868);
xor UO_214 (O_214,N_2513,N_2911);
nand UO_215 (O_215,N_2460,N_2499);
or UO_216 (O_216,N_2742,N_2617);
nand UO_217 (O_217,N_2814,N_2401);
nand UO_218 (O_218,N_2810,N_2632);
or UO_219 (O_219,N_2486,N_2844);
xnor UO_220 (O_220,N_2507,N_2930);
or UO_221 (O_221,N_2685,N_2820);
nor UO_222 (O_222,N_2954,N_2748);
and UO_223 (O_223,N_2589,N_2970);
xor UO_224 (O_224,N_2906,N_2645);
nand UO_225 (O_225,N_2912,N_2907);
and UO_226 (O_226,N_2526,N_2739);
nor UO_227 (O_227,N_2506,N_2490);
xnor UO_228 (O_228,N_2818,N_2519);
and UO_229 (O_229,N_2964,N_2745);
nand UO_230 (O_230,N_2760,N_2944);
or UO_231 (O_231,N_2578,N_2826);
nor UO_232 (O_232,N_2693,N_2547);
and UO_233 (O_233,N_2947,N_2751);
and UO_234 (O_234,N_2919,N_2722);
and UO_235 (O_235,N_2992,N_2539);
or UO_236 (O_236,N_2712,N_2437);
xnor UO_237 (O_237,N_2862,N_2619);
xnor UO_238 (O_238,N_2458,N_2435);
nand UO_239 (O_239,N_2841,N_2402);
nand UO_240 (O_240,N_2795,N_2537);
or UO_241 (O_241,N_2915,N_2707);
nand UO_242 (O_242,N_2488,N_2717);
nor UO_243 (O_243,N_2721,N_2932);
xor UO_244 (O_244,N_2680,N_2780);
nand UO_245 (O_245,N_2794,N_2412);
and UO_246 (O_246,N_2514,N_2525);
and UO_247 (O_247,N_2738,N_2557);
nand UO_248 (O_248,N_2807,N_2609);
nor UO_249 (O_249,N_2602,N_2675);
or UO_250 (O_250,N_2533,N_2469);
nand UO_251 (O_251,N_2535,N_2995);
xnor UO_252 (O_252,N_2728,N_2522);
nand UO_253 (O_253,N_2777,N_2503);
nor UO_254 (O_254,N_2508,N_2872);
nand UO_255 (O_255,N_2567,N_2965);
nand UO_256 (O_256,N_2592,N_2570);
and UO_257 (O_257,N_2706,N_2664);
or UO_258 (O_258,N_2433,N_2541);
or UO_259 (O_259,N_2504,N_2620);
xor UO_260 (O_260,N_2928,N_2939);
or UO_261 (O_261,N_2658,N_2414);
nand UO_262 (O_262,N_2408,N_2950);
nor UO_263 (O_263,N_2529,N_2676);
or UO_264 (O_264,N_2806,N_2580);
nand UO_265 (O_265,N_2953,N_2562);
xor UO_266 (O_266,N_2933,N_2768);
nand UO_267 (O_267,N_2552,N_2429);
xnor UO_268 (O_268,N_2804,N_2897);
nor UO_269 (O_269,N_2864,N_2746);
xnor UO_270 (O_270,N_2729,N_2456);
nand UO_271 (O_271,N_2834,N_2420);
nand UO_272 (O_272,N_2647,N_2639);
or UO_273 (O_273,N_2563,N_2857);
xor UO_274 (O_274,N_2416,N_2405);
nor UO_275 (O_275,N_2808,N_2848);
xor UO_276 (O_276,N_2644,N_2560);
xor UO_277 (O_277,N_2678,N_2877);
or UO_278 (O_278,N_2649,N_2955);
nor UO_279 (O_279,N_2771,N_2461);
or UO_280 (O_280,N_2725,N_2449);
nand UO_281 (O_281,N_2422,N_2743);
xnor UO_282 (O_282,N_2511,N_2931);
or UO_283 (O_283,N_2784,N_2761);
nand UO_284 (O_284,N_2790,N_2542);
nor UO_285 (O_285,N_2753,N_2653);
and UO_286 (O_286,N_2571,N_2936);
nand UO_287 (O_287,N_2409,N_2719);
nor UO_288 (O_288,N_2781,N_2556);
nand UO_289 (O_289,N_2494,N_2521);
and UO_290 (O_290,N_2641,N_2555);
xnor UO_291 (O_291,N_2986,N_2674);
nand UO_292 (O_292,N_2534,N_2752);
xnor UO_293 (O_293,N_2960,N_2798);
nor UO_294 (O_294,N_2896,N_2629);
xnor UO_295 (O_295,N_2849,N_2476);
nand UO_296 (O_296,N_2404,N_2424);
and UO_297 (O_297,N_2876,N_2901);
and UO_298 (O_298,N_2861,N_2949);
and UO_299 (O_299,N_2863,N_2439);
nor UO_300 (O_300,N_2968,N_2643);
and UO_301 (O_301,N_2424,N_2620);
nor UO_302 (O_302,N_2460,N_2808);
and UO_303 (O_303,N_2879,N_2413);
or UO_304 (O_304,N_2919,N_2412);
and UO_305 (O_305,N_2672,N_2995);
nor UO_306 (O_306,N_2442,N_2888);
or UO_307 (O_307,N_2435,N_2751);
nand UO_308 (O_308,N_2521,N_2864);
nor UO_309 (O_309,N_2624,N_2563);
nor UO_310 (O_310,N_2899,N_2404);
nor UO_311 (O_311,N_2838,N_2992);
or UO_312 (O_312,N_2404,N_2907);
nor UO_313 (O_313,N_2570,N_2591);
and UO_314 (O_314,N_2661,N_2883);
xor UO_315 (O_315,N_2404,N_2982);
and UO_316 (O_316,N_2579,N_2751);
and UO_317 (O_317,N_2716,N_2882);
xnor UO_318 (O_318,N_2791,N_2981);
nor UO_319 (O_319,N_2464,N_2920);
nor UO_320 (O_320,N_2809,N_2584);
or UO_321 (O_321,N_2735,N_2707);
nand UO_322 (O_322,N_2443,N_2635);
and UO_323 (O_323,N_2793,N_2932);
nor UO_324 (O_324,N_2404,N_2965);
nor UO_325 (O_325,N_2572,N_2959);
xnor UO_326 (O_326,N_2759,N_2937);
and UO_327 (O_327,N_2773,N_2445);
nand UO_328 (O_328,N_2641,N_2480);
or UO_329 (O_329,N_2495,N_2591);
nand UO_330 (O_330,N_2617,N_2621);
xor UO_331 (O_331,N_2882,N_2441);
nor UO_332 (O_332,N_2834,N_2692);
and UO_333 (O_333,N_2780,N_2950);
xnor UO_334 (O_334,N_2580,N_2609);
and UO_335 (O_335,N_2712,N_2717);
or UO_336 (O_336,N_2697,N_2471);
xnor UO_337 (O_337,N_2617,N_2625);
and UO_338 (O_338,N_2923,N_2984);
and UO_339 (O_339,N_2687,N_2966);
nor UO_340 (O_340,N_2972,N_2614);
nor UO_341 (O_341,N_2487,N_2685);
nor UO_342 (O_342,N_2777,N_2611);
and UO_343 (O_343,N_2710,N_2824);
nor UO_344 (O_344,N_2446,N_2920);
nand UO_345 (O_345,N_2552,N_2545);
and UO_346 (O_346,N_2986,N_2516);
nor UO_347 (O_347,N_2487,N_2810);
or UO_348 (O_348,N_2622,N_2491);
nand UO_349 (O_349,N_2809,N_2587);
nor UO_350 (O_350,N_2808,N_2486);
or UO_351 (O_351,N_2604,N_2900);
and UO_352 (O_352,N_2438,N_2553);
and UO_353 (O_353,N_2602,N_2631);
nand UO_354 (O_354,N_2509,N_2471);
and UO_355 (O_355,N_2597,N_2613);
xor UO_356 (O_356,N_2820,N_2838);
nor UO_357 (O_357,N_2480,N_2619);
nand UO_358 (O_358,N_2490,N_2587);
nand UO_359 (O_359,N_2400,N_2909);
and UO_360 (O_360,N_2840,N_2714);
and UO_361 (O_361,N_2962,N_2541);
nand UO_362 (O_362,N_2802,N_2756);
and UO_363 (O_363,N_2719,N_2780);
xor UO_364 (O_364,N_2686,N_2605);
and UO_365 (O_365,N_2822,N_2618);
or UO_366 (O_366,N_2691,N_2624);
or UO_367 (O_367,N_2450,N_2525);
xnor UO_368 (O_368,N_2569,N_2427);
nand UO_369 (O_369,N_2554,N_2864);
or UO_370 (O_370,N_2612,N_2461);
nor UO_371 (O_371,N_2757,N_2434);
and UO_372 (O_372,N_2445,N_2429);
xor UO_373 (O_373,N_2990,N_2433);
nor UO_374 (O_374,N_2726,N_2686);
and UO_375 (O_375,N_2942,N_2513);
nand UO_376 (O_376,N_2570,N_2540);
and UO_377 (O_377,N_2763,N_2944);
xor UO_378 (O_378,N_2957,N_2972);
nand UO_379 (O_379,N_2776,N_2600);
nor UO_380 (O_380,N_2615,N_2535);
and UO_381 (O_381,N_2628,N_2564);
nor UO_382 (O_382,N_2949,N_2881);
or UO_383 (O_383,N_2613,N_2400);
and UO_384 (O_384,N_2783,N_2558);
or UO_385 (O_385,N_2433,N_2708);
nor UO_386 (O_386,N_2975,N_2489);
nand UO_387 (O_387,N_2878,N_2422);
or UO_388 (O_388,N_2927,N_2555);
or UO_389 (O_389,N_2899,N_2533);
nand UO_390 (O_390,N_2456,N_2523);
nand UO_391 (O_391,N_2578,N_2401);
xnor UO_392 (O_392,N_2469,N_2608);
nand UO_393 (O_393,N_2668,N_2505);
or UO_394 (O_394,N_2485,N_2809);
or UO_395 (O_395,N_2839,N_2613);
and UO_396 (O_396,N_2643,N_2506);
and UO_397 (O_397,N_2591,N_2770);
or UO_398 (O_398,N_2648,N_2794);
xnor UO_399 (O_399,N_2728,N_2550);
nor UO_400 (O_400,N_2979,N_2544);
xnor UO_401 (O_401,N_2415,N_2619);
and UO_402 (O_402,N_2613,N_2600);
or UO_403 (O_403,N_2445,N_2437);
and UO_404 (O_404,N_2401,N_2905);
nand UO_405 (O_405,N_2592,N_2623);
xnor UO_406 (O_406,N_2815,N_2802);
xnor UO_407 (O_407,N_2624,N_2911);
nand UO_408 (O_408,N_2660,N_2507);
nand UO_409 (O_409,N_2813,N_2443);
nor UO_410 (O_410,N_2565,N_2626);
xor UO_411 (O_411,N_2983,N_2940);
nor UO_412 (O_412,N_2401,N_2842);
or UO_413 (O_413,N_2966,N_2791);
xnor UO_414 (O_414,N_2569,N_2584);
and UO_415 (O_415,N_2630,N_2943);
nor UO_416 (O_416,N_2472,N_2480);
nand UO_417 (O_417,N_2917,N_2598);
xnor UO_418 (O_418,N_2777,N_2947);
nand UO_419 (O_419,N_2846,N_2710);
or UO_420 (O_420,N_2486,N_2568);
nor UO_421 (O_421,N_2780,N_2417);
xnor UO_422 (O_422,N_2702,N_2914);
xnor UO_423 (O_423,N_2777,N_2425);
xnor UO_424 (O_424,N_2654,N_2646);
nand UO_425 (O_425,N_2506,N_2445);
xnor UO_426 (O_426,N_2856,N_2980);
or UO_427 (O_427,N_2408,N_2856);
nor UO_428 (O_428,N_2506,N_2418);
and UO_429 (O_429,N_2553,N_2881);
nand UO_430 (O_430,N_2523,N_2554);
xnor UO_431 (O_431,N_2990,N_2505);
nor UO_432 (O_432,N_2702,N_2563);
xor UO_433 (O_433,N_2692,N_2515);
or UO_434 (O_434,N_2544,N_2730);
nand UO_435 (O_435,N_2981,N_2691);
and UO_436 (O_436,N_2860,N_2887);
or UO_437 (O_437,N_2576,N_2676);
or UO_438 (O_438,N_2668,N_2528);
nor UO_439 (O_439,N_2933,N_2975);
xor UO_440 (O_440,N_2946,N_2779);
or UO_441 (O_441,N_2921,N_2476);
nor UO_442 (O_442,N_2435,N_2506);
and UO_443 (O_443,N_2838,N_2955);
nand UO_444 (O_444,N_2743,N_2608);
xnor UO_445 (O_445,N_2730,N_2423);
nand UO_446 (O_446,N_2433,N_2524);
xnor UO_447 (O_447,N_2611,N_2754);
xnor UO_448 (O_448,N_2653,N_2991);
or UO_449 (O_449,N_2762,N_2472);
nand UO_450 (O_450,N_2809,N_2836);
and UO_451 (O_451,N_2770,N_2729);
nand UO_452 (O_452,N_2613,N_2883);
nand UO_453 (O_453,N_2420,N_2734);
or UO_454 (O_454,N_2550,N_2709);
or UO_455 (O_455,N_2408,N_2610);
nor UO_456 (O_456,N_2478,N_2809);
nand UO_457 (O_457,N_2949,N_2723);
or UO_458 (O_458,N_2899,N_2727);
nand UO_459 (O_459,N_2499,N_2742);
nor UO_460 (O_460,N_2810,N_2417);
and UO_461 (O_461,N_2847,N_2665);
and UO_462 (O_462,N_2758,N_2648);
and UO_463 (O_463,N_2579,N_2839);
nor UO_464 (O_464,N_2598,N_2663);
xnor UO_465 (O_465,N_2949,N_2535);
xnor UO_466 (O_466,N_2631,N_2819);
nor UO_467 (O_467,N_2991,N_2486);
xor UO_468 (O_468,N_2457,N_2810);
nand UO_469 (O_469,N_2908,N_2644);
nand UO_470 (O_470,N_2421,N_2528);
or UO_471 (O_471,N_2992,N_2528);
and UO_472 (O_472,N_2848,N_2559);
and UO_473 (O_473,N_2442,N_2884);
nand UO_474 (O_474,N_2565,N_2679);
xor UO_475 (O_475,N_2721,N_2823);
nor UO_476 (O_476,N_2712,N_2810);
nor UO_477 (O_477,N_2959,N_2769);
nand UO_478 (O_478,N_2781,N_2608);
or UO_479 (O_479,N_2676,N_2533);
nor UO_480 (O_480,N_2451,N_2578);
nand UO_481 (O_481,N_2534,N_2615);
nand UO_482 (O_482,N_2631,N_2549);
nand UO_483 (O_483,N_2794,N_2737);
nand UO_484 (O_484,N_2618,N_2758);
or UO_485 (O_485,N_2409,N_2908);
nand UO_486 (O_486,N_2973,N_2750);
nor UO_487 (O_487,N_2951,N_2941);
and UO_488 (O_488,N_2816,N_2912);
or UO_489 (O_489,N_2791,N_2933);
nand UO_490 (O_490,N_2615,N_2608);
and UO_491 (O_491,N_2884,N_2475);
or UO_492 (O_492,N_2812,N_2983);
or UO_493 (O_493,N_2928,N_2925);
and UO_494 (O_494,N_2960,N_2974);
nand UO_495 (O_495,N_2739,N_2705);
xor UO_496 (O_496,N_2468,N_2719);
xnor UO_497 (O_497,N_2495,N_2759);
and UO_498 (O_498,N_2809,N_2907);
nor UO_499 (O_499,N_2954,N_2946);
endmodule