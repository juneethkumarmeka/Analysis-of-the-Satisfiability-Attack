module basic_2000_20000_2500_50_levels_1xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_613,In_1272);
nor U1 (N_1,In_1842,In_1136);
or U2 (N_2,In_720,In_1478);
or U3 (N_3,In_858,In_1578);
nor U4 (N_4,In_1904,In_919);
nor U5 (N_5,In_1969,In_1351);
and U6 (N_6,In_553,In_1252);
or U7 (N_7,In_1838,In_1812);
or U8 (N_8,In_1165,In_1817);
nor U9 (N_9,In_795,In_1556);
nand U10 (N_10,In_1231,In_1859);
nand U11 (N_11,In_305,In_1385);
nor U12 (N_12,In_1721,In_88);
and U13 (N_13,In_95,In_1359);
and U14 (N_14,In_1271,In_859);
nor U15 (N_15,In_307,In_1958);
or U16 (N_16,In_1002,In_1626);
or U17 (N_17,In_1462,In_914);
nor U18 (N_18,In_1083,In_162);
or U19 (N_19,In_59,In_1306);
nor U20 (N_20,In_1387,In_703);
and U21 (N_21,In_632,In_130);
or U22 (N_22,In_997,In_364);
and U23 (N_23,In_1069,In_690);
nor U24 (N_24,In_1996,In_965);
nor U25 (N_25,In_1656,In_878);
nor U26 (N_26,In_836,In_984);
nor U27 (N_27,In_966,In_1919);
and U28 (N_28,In_1939,In_1100);
or U29 (N_29,In_917,In_1960);
nor U30 (N_30,In_1210,In_1161);
or U31 (N_31,In_1664,In_956);
and U32 (N_32,In_758,In_681);
and U33 (N_33,In_55,In_1605);
nand U34 (N_34,In_294,In_346);
nand U35 (N_35,In_1738,In_749);
nand U36 (N_36,In_1752,In_834);
nand U37 (N_37,In_1680,In_1034);
nor U38 (N_38,In_1971,In_715);
or U39 (N_39,In_37,In_1985);
nor U40 (N_40,In_1160,In_92);
nor U41 (N_41,In_134,In_1689);
nand U42 (N_42,In_867,In_281);
or U43 (N_43,In_124,In_838);
nand U44 (N_44,In_1714,In_495);
nand U45 (N_45,In_866,In_1997);
or U46 (N_46,In_136,In_308);
nor U47 (N_47,In_140,In_1800);
nor U48 (N_48,In_1159,In_1312);
or U49 (N_49,In_148,In_1);
nor U50 (N_50,In_893,In_102);
or U51 (N_51,In_145,In_1608);
and U52 (N_52,In_1867,In_1707);
nor U53 (N_53,In_1943,In_1789);
nand U54 (N_54,In_629,In_853);
nor U55 (N_55,In_283,In_454);
xnor U56 (N_56,In_752,In_497);
nor U57 (N_57,In_1585,In_566);
or U58 (N_58,In_706,In_107);
nand U59 (N_59,In_772,In_1023);
nor U60 (N_60,In_119,In_1887);
nor U61 (N_61,In_872,In_0);
nand U62 (N_62,In_1956,In_1729);
and U63 (N_63,In_194,In_252);
or U64 (N_64,In_1910,In_1148);
or U65 (N_65,In_1932,In_328);
or U66 (N_66,In_441,In_1764);
nor U67 (N_67,In_1938,In_774);
nand U68 (N_68,In_1211,In_508);
or U69 (N_69,In_680,In_1001);
nor U70 (N_70,In_266,In_988);
or U71 (N_71,In_773,In_1894);
or U72 (N_72,In_202,In_1056);
and U73 (N_73,In_1831,In_1837);
nand U74 (N_74,In_216,In_1516);
nor U75 (N_75,In_1779,In_1860);
nor U76 (N_76,In_1878,In_763);
and U77 (N_77,In_1039,In_1122);
nor U78 (N_78,In_1114,In_1603);
and U79 (N_79,In_951,In_709);
and U80 (N_80,In_1152,In_707);
nor U81 (N_81,In_1126,In_1518);
or U82 (N_82,In_998,In_556);
nor U83 (N_83,In_1482,In_365);
or U84 (N_84,In_1305,In_1671);
nand U85 (N_85,In_1929,In_1979);
nand U86 (N_86,In_232,In_1639);
nand U87 (N_87,In_837,In_402);
and U88 (N_88,In_1690,In_1710);
nand U89 (N_89,In_577,In_1258);
nor U90 (N_90,In_658,In_527);
and U91 (N_91,In_297,In_846);
nor U92 (N_92,In_980,In_864);
or U93 (N_93,In_849,In_1974);
or U94 (N_94,In_1949,In_1217);
or U95 (N_95,In_383,In_538);
nor U96 (N_96,In_169,In_356);
or U97 (N_97,In_1803,In_950);
and U98 (N_98,In_1830,In_1614);
or U99 (N_99,In_764,In_1374);
nor U100 (N_100,In_381,In_1358);
and U101 (N_101,In_475,In_1437);
or U102 (N_102,In_1247,In_66);
nor U103 (N_103,In_1266,In_1654);
or U104 (N_104,In_1873,In_1469);
and U105 (N_105,In_372,In_334);
and U106 (N_106,In_1570,In_300);
and U107 (N_107,In_1248,In_1554);
or U108 (N_108,In_783,In_1550);
and U109 (N_109,In_712,In_104);
nor U110 (N_110,In_127,In_1401);
nand U111 (N_111,In_560,In_1809);
nand U112 (N_112,In_903,In_871);
nor U113 (N_113,In_228,In_995);
or U114 (N_114,In_1747,In_270);
nor U115 (N_115,In_295,In_367);
nor U116 (N_116,In_762,In_370);
nand U117 (N_117,In_1879,In_807);
nor U118 (N_118,In_1107,In_811);
nor U119 (N_119,In_1262,In_319);
and U120 (N_120,In_357,In_354);
nor U121 (N_121,In_1653,In_682);
nand U122 (N_122,In_1447,In_415);
nand U123 (N_123,In_1806,In_1111);
nor U124 (N_124,In_1998,In_873);
and U125 (N_125,In_1983,In_1142);
nand U126 (N_126,In_510,In_1127);
nor U127 (N_127,In_1383,In_1029);
nand U128 (N_128,In_1991,In_1776);
nor U129 (N_129,In_641,In_1453);
and U130 (N_130,In_474,In_575);
nor U131 (N_131,In_1347,In_458);
or U132 (N_132,In_593,In_1670);
or U133 (N_133,In_278,In_1703);
or U134 (N_134,In_1658,In_1650);
nor U135 (N_135,In_149,In_430);
and U136 (N_136,In_1027,In_1529);
or U137 (N_137,In_1009,In_746);
or U138 (N_138,In_588,In_1396);
nand U139 (N_139,In_1778,In_1203);
and U140 (N_140,In_1790,In_1375);
or U141 (N_141,In_1019,In_1477);
nand U142 (N_142,In_755,In_833);
nand U143 (N_143,In_481,In_1566);
nand U144 (N_144,In_1176,In_516);
and U145 (N_145,In_1087,In_1709);
nand U146 (N_146,In_439,In_1720);
nor U147 (N_147,In_1547,In_1304);
or U148 (N_148,In_1422,In_627);
and U149 (N_149,In_1907,In_1191);
nor U150 (N_150,In_842,In_1851);
and U151 (N_151,In_192,In_1299);
or U152 (N_152,In_1571,In_932);
nand U153 (N_153,In_604,In_960);
and U154 (N_154,In_663,In_1786);
or U155 (N_155,In_1891,In_573);
nand U156 (N_156,In_1818,In_939);
nand U157 (N_157,In_289,In_2);
nor U158 (N_158,In_653,In_1758);
or U159 (N_159,In_431,In_1510);
nand U160 (N_160,In_1535,In_462);
and U161 (N_161,In_455,In_1441);
and U162 (N_162,In_1622,In_111);
nor U163 (N_163,In_1508,In_857);
nand U164 (N_164,In_243,In_794);
nor U165 (N_165,In_994,In_468);
nor U166 (N_166,In_445,In_1874);
or U167 (N_167,In_220,In_193);
nand U168 (N_168,In_689,In_677);
xor U169 (N_169,In_987,In_1538);
nand U170 (N_170,In_1452,In_944);
and U171 (N_171,In_1931,In_1674);
or U172 (N_172,In_234,In_638);
nor U173 (N_173,In_427,In_157);
or U174 (N_174,In_1309,In_1026);
and U175 (N_175,In_963,In_831);
and U176 (N_176,In_1435,In_276);
nor U177 (N_177,In_719,In_159);
nor U178 (N_178,In_760,In_1701);
and U179 (N_179,In_514,In_338);
or U180 (N_180,In_1175,In_1796);
or U181 (N_181,In_302,In_1651);
nand U182 (N_182,In_1143,In_1755);
nand U183 (N_183,In_1320,In_531);
and U184 (N_184,In_579,In_1540);
nand U185 (N_185,In_513,In_1060);
nand U186 (N_186,In_1801,In_105);
or U187 (N_187,In_373,In_1464);
nand U188 (N_188,In_417,In_1303);
and U189 (N_189,In_1468,In_246);
and U190 (N_190,In_470,In_160);
nor U191 (N_191,In_1679,In_1333);
or U192 (N_192,In_606,In_170);
nor U193 (N_193,In_1963,In_517);
xnor U194 (N_194,In_1367,In_1908);
and U195 (N_195,In_961,In_1524);
or U196 (N_196,In_1613,In_1532);
nor U197 (N_197,In_753,In_282);
and U198 (N_198,In_648,In_167);
nand U199 (N_199,In_1757,In_662);
nor U200 (N_200,In_985,In_436);
nand U201 (N_201,In_1986,In_637);
or U202 (N_202,In_110,In_844);
and U203 (N_203,In_459,In_1492);
and U204 (N_204,In_1182,In_896);
nand U205 (N_205,In_444,In_141);
or U206 (N_206,In_1055,In_1025);
and U207 (N_207,In_1989,In_418);
and U208 (N_208,In_1744,In_1461);
and U209 (N_209,In_535,In_1300);
and U210 (N_210,In_1378,In_1393);
and U211 (N_211,In_482,In_1683);
or U212 (N_212,In_804,In_1255);
and U213 (N_213,In_976,In_242);
nand U214 (N_214,In_711,In_1352);
nand U215 (N_215,In_938,In_1233);
nand U216 (N_216,In_313,In_1728);
nand U217 (N_217,In_818,In_473);
and U218 (N_218,In_1037,In_476);
nor U219 (N_219,In_685,In_1768);
nor U220 (N_220,In_1644,In_70);
nor U221 (N_221,In_260,In_983);
or U222 (N_222,In_973,In_683);
nor U223 (N_223,In_256,In_578);
nand U224 (N_224,In_695,In_812);
nor U225 (N_225,In_684,In_123);
nand U226 (N_226,In_1909,In_1414);
or U227 (N_227,In_1253,In_1513);
or U228 (N_228,In_1155,In_1501);
nor U229 (N_229,In_1869,In_1727);
or U230 (N_230,In_608,In_1017);
and U231 (N_231,In_1959,In_1593);
nor U232 (N_232,In_290,In_1350);
nand U233 (N_233,In_1199,In_1973);
or U234 (N_234,In_924,In_1928);
nor U235 (N_235,In_530,In_1844);
nand U236 (N_236,In_740,In_1804);
nand U237 (N_237,In_261,In_977);
nor U238 (N_238,In_1313,In_744);
nand U239 (N_239,In_1207,In_1016);
and U240 (N_240,In_580,In_1681);
nor U241 (N_241,In_541,In_301);
and U242 (N_242,In_499,In_1379);
or U243 (N_243,In_1097,In_840);
and U244 (N_244,In_1224,In_1527);
and U245 (N_245,In_1687,In_1723);
and U246 (N_246,In_1024,In_68);
nor U247 (N_247,In_1074,In_292);
and U248 (N_248,In_1444,In_350);
nor U249 (N_249,In_63,In_910);
or U250 (N_250,In_1657,In_1865);
and U251 (N_251,In_974,In_1490);
nand U252 (N_252,In_1665,In_1712);
nand U253 (N_253,In_955,In_1813);
nor U254 (N_254,In_953,In_723);
nand U255 (N_255,In_1805,In_1449);
xnor U256 (N_256,In_856,In_471);
nand U257 (N_257,In_333,In_404);
nor U258 (N_258,In_1999,In_1408);
nor U259 (N_259,In_1793,In_1440);
or U260 (N_260,In_1648,In_1584);
or U261 (N_261,In_1426,In_562);
nor U262 (N_262,In_224,In_1877);
nand U263 (N_263,In_1495,In_74);
nand U264 (N_264,In_1334,In_787);
nor U265 (N_265,In_756,In_480);
or U266 (N_266,In_1941,In_279);
and U267 (N_267,In_710,In_1256);
nor U268 (N_268,In_751,In_1115);
nor U269 (N_269,In_520,In_1050);
nor U270 (N_270,In_178,In_1412);
or U271 (N_271,In_957,In_633);
nand U272 (N_272,In_1289,In_212);
nor U273 (N_273,In_626,In_1880);
nand U274 (N_274,In_1968,In_1251);
or U275 (N_275,In_750,In_1814);
and U276 (N_276,In_195,In_336);
nor U277 (N_277,In_1295,In_1870);
or U278 (N_278,In_1676,In_948);
or U279 (N_279,In_1118,In_1748);
and U280 (N_280,In_401,In_1641);
and U281 (N_281,In_1771,In_1112);
and U282 (N_282,In_640,In_902);
nand U283 (N_283,In_666,In_1195);
and U284 (N_284,In_203,In_1277);
nor U285 (N_285,In_1609,In_1276);
and U286 (N_286,In_1371,In_1882);
nand U287 (N_287,In_1067,In_1032);
or U288 (N_288,In_156,In_1544);
nand U289 (N_289,In_1265,In_1014);
or U290 (N_290,In_1677,In_1476);
nor U291 (N_291,In_1328,In_398);
nand U292 (N_292,In_971,In_1395);
nor U293 (N_293,In_868,In_1912);
and U294 (N_294,In_1733,In_1153);
nand U295 (N_295,In_1872,In_671);
nor U296 (N_296,In_40,In_574);
nand U297 (N_297,In_1128,In_1763);
nor U298 (N_298,In_355,In_1397);
and U299 (N_299,In_1632,In_726);
nand U300 (N_300,In_748,In_941);
or U301 (N_301,In_236,In_1829);
nor U302 (N_302,In_25,In_549);
nor U303 (N_303,In_1144,In_821);
and U304 (N_304,In_1995,In_1215);
and U305 (N_305,In_1004,In_90);
nand U306 (N_306,In_1560,In_264);
nor U307 (N_307,In_359,In_1784);
nor U308 (N_308,In_805,In_1561);
and U309 (N_309,In_323,In_547);
or U310 (N_310,In_1746,In_879);
nor U311 (N_311,In_808,In_569);
xnor U312 (N_312,In_1848,In_1316);
nor U313 (N_313,In_1293,In_1274);
nand U314 (N_314,In_1332,In_274);
or U315 (N_315,In_1612,In_1052);
or U316 (N_316,In_1214,In_675);
nor U317 (N_317,In_1288,In_1766);
xor U318 (N_318,In_1826,In_506);
or U319 (N_319,In_13,In_1167);
or U320 (N_320,In_1652,In_191);
nor U321 (N_321,In_440,In_979);
and U322 (N_322,In_429,In_1765);
nand U323 (N_323,In_610,In_803);
or U324 (N_324,In_518,In_1028);
nand U325 (N_325,In_1345,In_1698);
nand U326 (N_326,In_1018,In_1607);
and U327 (N_327,In_1530,In_1156);
nor U328 (N_328,In_1811,In_233);
nand U329 (N_329,In_1116,In_1284);
and U330 (N_330,In_1964,In_507);
nand U331 (N_331,In_1278,In_215);
or U332 (N_332,In_767,In_407);
nor U333 (N_333,In_1770,In_806);
nand U334 (N_334,In_1886,In_391);
nor U335 (N_335,In_1285,In_1240);
and U336 (N_336,In_921,In_349);
and U337 (N_337,In_227,In_320);
nor U338 (N_338,In_1740,In_1117);
nand U339 (N_339,In_213,In_1047);
and U340 (N_340,In_1732,In_490);
nor U341 (N_341,In_1166,In_1125);
or U342 (N_342,In_1761,In_643);
or U343 (N_343,In_1405,In_327);
nand U344 (N_344,In_1230,In_413);
or U345 (N_345,In_352,In_1343);
and U346 (N_346,In_396,In_1846);
xor U347 (N_347,In_1536,In_784);
and U348 (N_348,In_27,In_1467);
nor U349 (N_349,In_151,In_1470);
nand U350 (N_350,In_1237,In_489);
and U351 (N_351,In_32,In_1448);
and U352 (N_352,In_542,In_1668);
and U353 (N_353,In_1353,In_1807);
and U354 (N_354,In_933,In_1617);
nand U355 (N_355,In_799,In_713);
and U356 (N_356,In_908,In_1080);
nand U357 (N_357,In_1031,In_434);
nand U358 (N_358,In_1139,In_863);
or U359 (N_359,In_1012,In_511);
or U360 (N_360,In_897,In_649);
and U361 (N_361,In_1413,In_12);
or U362 (N_362,In_990,In_57);
and U363 (N_363,In_1781,In_185);
nand U364 (N_364,In_1390,In_1522);
nor U365 (N_365,In_188,In_565);
xnor U366 (N_366,In_1917,In_1472);
nor U367 (N_367,In_96,In_1586);
xor U368 (N_368,In_888,In_1380);
nand U369 (N_369,In_850,In_1914);
nor U370 (N_370,In_247,In_344);
nor U371 (N_371,In_1219,In_901);
or U372 (N_372,In_1715,In_72);
and U373 (N_373,In_993,In_815);
nand U374 (N_374,In_584,In_991);
nand U375 (N_375,In_539,In_645);
and U376 (N_376,In_1775,In_1824);
nor U377 (N_377,In_285,In_989);
and U378 (N_378,In_1718,In_1488);
nand U379 (N_379,In_1006,In_1298);
and U380 (N_380,In_1895,In_1213);
and U381 (N_381,In_1945,In_909);
nor U382 (N_382,In_1456,In_615);
nor U383 (N_383,In_639,In_887);
nand U384 (N_384,In_718,In_1551);
or U385 (N_385,In_1040,In_56);
nand U386 (N_386,In_1212,In_1466);
nand U387 (N_387,In_1889,In_54);
nand U388 (N_388,In_550,In_1338);
and U389 (N_389,In_1364,In_1699);
nand U390 (N_390,In_26,In_35);
and U391 (N_391,In_17,In_1916);
and U392 (N_392,In_1311,In_464);
nor U393 (N_393,In_1885,In_1283);
or U394 (N_394,In_725,In_730);
nand U395 (N_395,In_1427,In_451);
nor U396 (N_396,In_1317,In_1137);
or U397 (N_397,In_1434,In_1647);
nand U398 (N_398,In_1954,In_347);
nor U399 (N_399,In_1138,In_479);
nand U400 (N_400,In_1777,In_1084);
and U401 (N_401,In_1496,N_376);
or U402 (N_402,In_71,In_1226);
and U403 (N_403,In_722,In_696);
nand U404 (N_404,N_354,In_674);
and U405 (N_405,In_714,In_1043);
and U406 (N_406,N_217,N_159);
nand U407 (N_407,In_1600,In_154);
and U408 (N_408,In_326,In_472);
nand U409 (N_409,N_302,In_403);
nor U410 (N_410,In_1322,In_885);
and U411 (N_411,In_1168,In_612);
or U412 (N_412,In_1753,In_1569);
nor U413 (N_413,In_665,In_654);
nor U414 (N_414,In_727,In_1325);
and U415 (N_415,In_882,In_869);
nor U416 (N_416,In_1319,In_312);
or U417 (N_417,In_655,In_1121);
or U418 (N_418,In_428,In_642);
or U419 (N_419,N_345,In_9);
nand U420 (N_420,In_1920,In_1636);
or U421 (N_421,In_1386,In_1129);
nor U422 (N_422,In_1509,In_1623);
nand U423 (N_423,In_915,In_230);
or U424 (N_424,In_636,In_412);
nand U425 (N_425,In_155,In_1179);
or U426 (N_426,In_830,In_150);
nand U427 (N_427,N_308,In_1596);
nand U428 (N_428,N_141,In_852);
nor U429 (N_429,N_44,In_1227);
or U430 (N_430,In_1988,In_694);
or U431 (N_431,N_242,In_982);
nor U432 (N_432,N_124,In_433);
or U433 (N_433,In_1066,In_1232);
or U434 (N_434,In_1575,N_254);
and U435 (N_435,N_276,In_704);
nor U436 (N_436,In_855,N_88);
nor U437 (N_437,N_148,N_107);
nor U438 (N_438,In_1756,N_115);
xor U439 (N_439,In_1281,In_1433);
and U440 (N_440,N_7,N_203);
nand U441 (N_441,In_44,In_1474);
or U442 (N_442,In_103,N_188);
nor U443 (N_443,N_123,In_442);
nand U444 (N_444,In_1362,In_601);
or U445 (N_445,In_1834,N_119);
nand U446 (N_446,N_191,In_1975);
nor U447 (N_447,In_1287,In_306);
nand U448 (N_448,In_1694,In_30);
nand U449 (N_449,In_1429,In_257);
nor U450 (N_450,N_233,In_238);
or U451 (N_451,N_216,N_67);
or U452 (N_452,In_1512,N_318);
nor U453 (N_453,In_1361,N_282);
nand U454 (N_454,In_620,N_306);
nor U455 (N_455,In_1822,N_176);
nor U456 (N_456,In_1123,In_309);
and U457 (N_457,In_776,In_1105);
nor U458 (N_458,N_287,N_373);
or U459 (N_459,In_981,In_1196);
and U460 (N_460,In_1109,N_359);
or U461 (N_461,In_1344,In_587);
nor U462 (N_462,In_1537,In_291);
nor U463 (N_463,In_1573,In_200);
and U464 (N_464,In_1297,N_362);
and U465 (N_465,In_1141,In_1257);
nor U466 (N_466,In_1135,In_1898);
or U467 (N_467,In_895,N_172);
and U468 (N_468,In_137,N_348);
nand U469 (N_469,In_1836,In_1944);
nand U470 (N_470,In_631,N_315);
or U471 (N_471,In_73,In_1923);
nor U472 (N_472,In_1905,In_1862);
nor U473 (N_473,N_355,In_1079);
nand U474 (N_474,N_383,N_334);
or U475 (N_475,N_270,In_628);
or U476 (N_476,In_1172,N_12);
or U477 (N_477,N_33,N_35);
and U478 (N_478,In_1799,N_155);
nor U479 (N_479,In_1481,In_724);
or U480 (N_480,In_771,In_22);
and U481 (N_481,N_174,N_160);
or U482 (N_482,In_65,In_745);
xnor U483 (N_483,N_136,In_1409);
or U484 (N_484,In_4,In_757);
nand U485 (N_485,In_1645,N_202);
nor U486 (N_486,In_1246,In_387);
or U487 (N_487,In_1268,N_256);
and U488 (N_488,In_1911,In_1145);
nand U489 (N_489,In_362,In_1314);
and U490 (N_490,In_1935,In_1534);
nand U491 (N_491,In_1500,In_699);
nor U492 (N_492,In_206,In_515);
nand U493 (N_493,In_91,N_89);
nor U494 (N_494,N_223,In_1451);
nand U495 (N_495,In_1542,In_721);
and U496 (N_496,In_839,N_31);
or U497 (N_497,In_646,In_847);
nor U498 (N_498,N_184,In_1631);
nor U499 (N_499,In_519,N_139);
or U500 (N_500,N_230,In_822);
or U501 (N_501,In_1235,In_503);
nor U502 (N_502,N_225,In_1339);
nand U503 (N_503,In_1342,N_11);
nand U504 (N_504,In_1130,In_1950);
or U505 (N_505,In_423,In_1013);
and U506 (N_506,In_1792,In_1952);
nor U507 (N_507,In_382,In_147);
or U508 (N_508,In_1331,In_1394);
nor U509 (N_509,N_167,N_154);
and U510 (N_510,In_172,In_1762);
and U511 (N_511,In_358,N_80);
and U512 (N_512,In_432,In_731);
and U513 (N_513,N_322,N_260);
and U514 (N_514,N_163,N_237);
nand U515 (N_515,In_1897,In_1693);
and U516 (N_516,In_778,In_221);
or U517 (N_517,In_1839,N_200);
nor U518 (N_518,N_198,In_884);
or U519 (N_519,In_862,N_5);
nor U520 (N_520,In_1341,In_255);
and U521 (N_521,In_487,In_378);
nand U522 (N_522,In_1169,N_241);
nor U523 (N_523,In_1388,In_1595);
and U524 (N_524,In_196,In_1183);
and U525 (N_525,N_209,In_1853);
or U526 (N_526,In_1722,In_978);
nand U527 (N_527,N_243,In_1154);
nor U528 (N_528,N_331,In_1222);
or U529 (N_529,In_500,N_374);
nand U530 (N_530,N_152,In_813);
and U531 (N_531,In_1627,N_101);
nor U532 (N_532,In_1021,In_265);
or U533 (N_533,In_1091,In_1783);
and U534 (N_534,N_342,In_1881);
nor U535 (N_535,In_734,N_72);
and U536 (N_536,In_935,In_325);
nor U537 (N_537,In_1948,In_874);
and U538 (N_538,N_197,In_996);
and U539 (N_539,N_103,In_1946);
xnor U540 (N_540,N_294,In_99);
nor U541 (N_541,In_1695,N_54);
nor U542 (N_542,In_1925,In_1120);
or U543 (N_543,In_463,N_244);
or U544 (N_544,N_47,In_406);
and U545 (N_545,In_421,N_280);
nor U546 (N_546,In_1625,In_1307);
and U547 (N_547,In_949,In_693);
and U548 (N_548,In_1696,In_1011);
nor U549 (N_549,N_168,In_698);
nand U550 (N_550,In_250,In_1725);
and U551 (N_551,In_85,In_453);
and U552 (N_552,In_1259,N_181);
nand U553 (N_553,In_1164,In_1033);
nand U554 (N_554,In_1022,In_1782);
nor U555 (N_555,In_786,N_114);
nor U556 (N_556,N_73,N_21);
or U557 (N_557,In_741,In_1147);
and U558 (N_558,In_1663,N_236);
nand U559 (N_559,In_1852,N_205);
nand U560 (N_560,In_1220,In_1900);
nand U561 (N_561,N_336,In_735);
or U562 (N_562,N_224,N_218);
nand U563 (N_563,In_1204,In_1146);
and U564 (N_564,In_450,N_96);
and U565 (N_565,In_667,In_1315);
nand U566 (N_566,In_164,In_1106);
or U567 (N_567,N_169,In_1892);
or U568 (N_568,In_1099,In_1735);
or U569 (N_569,In_943,In_1096);
nand U570 (N_570,In_1459,In_791);
nor U571 (N_571,In_1815,In_1808);
or U572 (N_572,In_465,In_118);
or U573 (N_573,In_1957,In_708);
or U574 (N_574,In_634,In_128);
and U575 (N_575,In_1599,In_1921);
nor U576 (N_576,In_1030,In_913);
nand U577 (N_577,In_311,In_819);
nor U578 (N_578,N_235,In_1977);
nand U579 (N_579,In_286,In_1193);
nand U580 (N_580,In_1238,In_1205);
nor U581 (N_581,In_937,N_99);
or U582 (N_582,In_1706,In_1810);
nor U583 (N_583,N_393,N_199);
nor U584 (N_584,In_1086,In_825);
nor U585 (N_585,In_1669,In_1423);
or U586 (N_586,In_174,In_343);
and U587 (N_587,N_229,N_48);
or U588 (N_588,In_371,In_657);
nand U589 (N_589,In_661,N_85);
and U590 (N_590,In_829,N_267);
and U591 (N_591,In_1678,In_1058);
nor U592 (N_592,In_754,In_1590);
or U593 (N_593,In_1719,In_181);
and U594 (N_594,In_1356,In_211);
and U595 (N_595,N_127,In_1321);
or U596 (N_596,In_133,In_165);
and U597 (N_597,In_186,In_737);
and U598 (N_598,In_1545,In_622);
or U599 (N_599,In_82,In_659);
nand U600 (N_600,In_115,N_13);
nor U601 (N_601,In_1875,In_168);
nor U602 (N_602,In_1151,In_229);
nor U603 (N_603,N_185,In_146);
nor U604 (N_604,In_14,N_162);
and U605 (N_605,In_399,In_318);
and U606 (N_606,In_792,In_678);
and U607 (N_607,N_134,In_1454);
and U608 (N_608,In_226,In_385);
nand U609 (N_609,In_1249,In_861);
nand U610 (N_610,In_559,In_1951);
and U611 (N_611,In_1411,In_322);
nor U612 (N_612,In_509,In_1505);
and U613 (N_613,In_1572,N_82);
nor U614 (N_614,In_624,In_1902);
or U615 (N_615,In_251,In_1171);
nor U616 (N_616,In_894,N_108);
and U617 (N_617,In_904,In_324);
or U618 (N_618,In_732,In_144);
nor U619 (N_619,N_333,N_51);
and U620 (N_620,In_525,N_398);
or U621 (N_621,In_5,In_1742);
or U622 (N_622,In_832,N_170);
or U623 (N_623,N_358,In_1794);
or U624 (N_624,In_1324,N_222);
nor U625 (N_625,In_1445,N_189);
nor U626 (N_626,In_1398,In_368);
nand U627 (N_627,In_197,In_1088);
or U628 (N_628,In_1797,N_367);
nand U629 (N_629,In_1736,N_221);
and U630 (N_630,N_219,In_1567);
or U631 (N_631,In_1688,In_1884);
and U632 (N_632,In_1294,In_502);
nor U633 (N_633,In_448,N_397);
or U634 (N_634,In_1533,In_494);
nor U635 (N_635,In_259,In_1857);
xor U636 (N_636,In_687,In_1541);
xor U637 (N_637,N_45,In_1073);
and U638 (N_638,In_1041,In_543);
nand U639 (N_639,In_1984,In_826);
and U640 (N_640,In_798,In_377);
nand U641 (N_641,In_1082,In_83);
and U642 (N_642,In_214,In_1833);
nand U643 (N_643,In_1015,In_876);
nand U644 (N_644,In_1577,In_78);
or U645 (N_645,In_1662,N_328);
or U646 (N_646,In_616,In_1503);
and U647 (N_647,N_86,N_272);
nor U648 (N_648,N_109,N_49);
nor U649 (N_649,In_1292,In_644);
or U650 (N_650,In_449,N_143);
or U651 (N_651,In_1992,N_293);
or U652 (N_652,In_422,In_1225);
and U653 (N_653,In_1749,In_1926);
nor U654 (N_654,In_594,N_271);
nand U655 (N_655,N_138,In_182);
or U656 (N_656,N_93,In_225);
nor U657 (N_657,In_1150,N_351);
nor U658 (N_658,In_1450,In_1876);
or U659 (N_659,N_150,N_375);
and U660 (N_660,In_335,N_281);
or U661 (N_661,N_17,In_733);
nand U662 (N_662,In_728,N_25);
nand U663 (N_663,In_485,In_1937);
or U664 (N_664,In_1188,N_58);
and U665 (N_665,N_180,In_789);
and U666 (N_666,N_356,In_1363);
nand U667 (N_667,In_1587,In_1296);
and U668 (N_668,In_1553,In_1955);
and U669 (N_669,N_196,In_576);
nor U670 (N_670,N_300,N_385);
or U671 (N_671,N_173,N_68);
or U672 (N_672,In_80,In_28);
and U673 (N_673,N_387,N_149);
nand U674 (N_674,N_171,In_1821);
or U675 (N_675,In_814,In_1619);
or U676 (N_676,In_1754,In_625);
or U677 (N_677,In_747,In_208);
or U678 (N_678,In_1318,In_34);
or U679 (N_679,In_1327,In_1399);
nor U680 (N_680,In_331,In_1635);
nor U681 (N_681,In_1443,N_344);
nand U682 (N_682,N_192,In_138);
nand U683 (N_683,In_366,In_1479);
or U684 (N_684,N_59,In_1871);
nor U685 (N_685,In_1489,In_1730);
nand U686 (N_686,In_46,In_1483);
nor U687 (N_687,N_301,N_190);
nand U688 (N_688,In_1198,In_705);
and U689 (N_689,In_1254,N_369);
and U690 (N_690,In_1391,N_105);
nor U691 (N_691,In_1899,In_1369);
and U692 (N_692,In_1863,In_1993);
and U693 (N_693,In_1471,In_962);
nor U694 (N_694,In_337,In_1078);
nand U695 (N_695,In_1200,N_275);
nor U696 (N_696,N_46,In_49);
or U697 (N_697,In_1308,In_1348);
or U698 (N_698,In_533,In_1692);
and U699 (N_699,N_361,In_880);
nor U700 (N_700,In_1242,N_102);
and U701 (N_701,In_304,In_1711);
or U702 (N_702,In_79,N_269);
nand U703 (N_703,In_100,In_1005);
or U704 (N_704,In_339,In_875);
nand U705 (N_705,N_4,In_1475);
and U706 (N_706,N_194,N_36);
nand U707 (N_707,N_38,In_1439);
and U708 (N_708,In_483,In_1181);
nor U709 (N_709,In_512,N_104);
nand U710 (N_710,In_452,In_800);
nand U711 (N_711,In_1346,In_1458);
xnor U712 (N_712,In_936,In_1045);
nand U713 (N_713,In_204,N_90);
or U714 (N_714,In_1402,In_848);
or U715 (N_715,In_1442,In_166);
nand U716 (N_716,In_1774,In_609);
nor U717 (N_717,In_1691,N_394);
nand U718 (N_718,In_1465,N_377);
nor U719 (N_719,In_1847,In_1197);
or U720 (N_720,In_1913,In_701);
and U721 (N_721,In_492,In_1646);
nor U722 (N_722,In_1686,In_1915);
or U723 (N_723,In_1485,N_319);
nor U724 (N_724,In_1134,In_1868);
nor U725 (N_725,In_1245,In_176);
or U726 (N_726,In_860,In_1557);
nand U727 (N_727,In_1549,In_388);
nand U728 (N_728,In_922,N_92);
or U729 (N_729,In_1666,In_883);
xnor U730 (N_730,In_469,N_78);
nand U731 (N_731,In_670,N_158);
and U732 (N_732,In_881,N_352);
or U733 (N_733,In_1404,In_1400);
and U734 (N_734,N_335,In_299);
nand U735 (N_735,In_892,In_1506);
nor U736 (N_736,N_388,N_65);
nand U737 (N_737,In_738,N_147);
or U738 (N_738,N_100,In_1003);
or U739 (N_739,In_1491,In_759);
xnor U740 (N_740,In_900,In_81);
or U741 (N_741,In_590,N_63);
nor U742 (N_742,In_607,In_20);
or U743 (N_743,In_199,In_504);
or U744 (N_744,In_970,In_143);
nor U745 (N_745,In_258,N_379);
nor U746 (N_746,In_1563,N_113);
and U747 (N_747,N_75,In_1773);
or U748 (N_748,N_226,In_69);
nor U749 (N_749,N_204,N_284);
or U750 (N_750,N_240,In_660);
or U751 (N_751,In_614,In_999);
nor U752 (N_752,In_1827,In_198);
or U753 (N_753,In_911,N_137);
nand U754 (N_754,In_1208,In_493);
nand U755 (N_755,In_1376,N_24);
nor U756 (N_756,In_1243,In_114);
or U757 (N_757,N_372,In_552);
and U758 (N_758,In_555,In_108);
or U759 (N_759,In_62,In_48);
nand U760 (N_760,In_1075,N_206);
nor U761 (N_761,In_782,In_563);
nand U762 (N_762,In_218,In_1173);
nor U763 (N_763,In_315,In_1372);
or U764 (N_764,In_1180,In_779);
nor U765 (N_765,In_1970,In_916);
nor U766 (N_766,In_1424,In_1978);
or U767 (N_767,N_118,N_52);
nor U768 (N_768,In_1201,N_215);
nand U769 (N_769,In_1514,In_602);
or U770 (N_770,In_557,In_38);
and U771 (N_771,N_297,In_53);
nor U772 (N_772,N_144,In_61);
nand U773 (N_773,N_391,In_1209);
or U774 (N_774,In_920,In_1724);
or U775 (N_775,N_161,In_769);
or U776 (N_776,In_390,In_183);
or U777 (N_777,In_945,In_1583);
nor U778 (N_778,In_790,N_132);
and U779 (N_779,In_117,N_238);
nand U780 (N_780,In_1640,N_349);
nand U781 (N_781,In_597,In_1972);
or U782 (N_782,In_1930,In_1425);
or U783 (N_783,In_1528,N_37);
nor U784 (N_784,In_1672,In_1062);
or U785 (N_785,In_1734,In_248);
nand U786 (N_786,In_546,In_1684);
and U787 (N_787,In_1832,N_258);
xor U788 (N_788,N_60,N_273);
nor U789 (N_789,In_1618,In_1323);
or U790 (N_790,In_1743,In_1936);
nor U791 (N_791,N_201,In_1499);
or U792 (N_792,N_324,In_820);
and U793 (N_793,In_1068,In_1858);
and U794 (N_794,In_457,In_1103);
nand U795 (N_795,In_1702,In_267);
and U796 (N_796,In_1463,In_1637);
xor U797 (N_797,In_589,In_1381);
and U798 (N_798,In_926,In_1520);
nor U799 (N_799,In_1704,In_877);
and U800 (N_800,N_327,N_630);
and U801 (N_801,N_728,N_628);
or U802 (N_802,N_632,N_557);
or U803 (N_803,In_405,In_1628);
or U804 (N_804,N_317,N_501);
nand U805 (N_805,N_542,In_353);
or U806 (N_806,In_967,In_523);
nor U807 (N_807,N_307,N_684);
and U808 (N_808,In_1697,N_245);
nand U809 (N_809,N_709,In_77);
or U810 (N_810,In_600,In_1008);
xor U811 (N_811,In_1487,In_1629);
nand U812 (N_812,N_321,N_430);
or U813 (N_813,N_178,N_689);
and U814 (N_814,N_476,N_474);
nand U815 (N_815,In_1416,In_51);
or U816 (N_816,In_275,In_36);
or U817 (N_817,In_360,N_637);
nand U818 (N_818,In_1229,N_396);
and U819 (N_819,In_1493,N_529);
nor U820 (N_820,In_1101,N_441);
nor U821 (N_821,In_1841,N_609);
nand U822 (N_822,N_478,N_40);
nand U823 (N_823,In_1194,In_558);
nand U824 (N_824,In_1455,N_432);
nor U825 (N_825,N_541,In_700);
nor U826 (N_826,N_309,N_122);
or U827 (N_827,N_611,In_621);
or U828 (N_828,N_257,N_567);
or U829 (N_829,N_3,N_692);
or U830 (N_830,N_494,In_142);
or U831 (N_831,N_664,In_1250);
nand U832 (N_832,In_122,N_536);
nand U833 (N_833,N_699,N_175);
nor U834 (N_834,N_511,In_1302);
nand U835 (N_835,In_1384,In_262);
and U836 (N_836,In_1990,N_702);
nand U837 (N_837,In_544,In_392);
nor U838 (N_838,N_485,N_489);
or U839 (N_839,In_1177,N_66);
nand U840 (N_840,In_1337,In_298);
xnor U841 (N_841,N_543,In_93);
or U842 (N_842,In_1081,N_695);
nand U843 (N_843,In_1185,N_296);
nor U844 (N_844,In_777,In_567);
and U845 (N_845,In_1054,N_453);
nand U846 (N_846,In_158,N_341);
and U847 (N_847,N_20,In_424);
and U848 (N_848,N_651,In_345);
nor U849 (N_849,In_1890,N_261);
nor U850 (N_850,In_231,N_460);
or U851 (N_851,In_1113,N_10);
nor U852 (N_852,In_1558,In_1038);
nor U853 (N_853,In_1591,N_305);
nor U854 (N_854,In_1419,In_461);
xor U855 (N_855,N_769,In_545);
or U856 (N_856,In_925,In_1849);
nor U857 (N_857,N_610,In_1065);
nand U858 (N_858,N_623,N_568);
and U859 (N_859,In_561,In_425);
and U860 (N_860,N_298,N_440);
or U861 (N_861,In_1349,In_788);
and U862 (N_862,In_420,In_460);
or U863 (N_863,In_1132,N_266);
nor U864 (N_864,N_76,In_688);
nor U865 (N_865,N_130,N_97);
nand U866 (N_866,N_777,N_520);
and U867 (N_867,In_1555,N_427);
and U868 (N_868,N_274,In_184);
and U869 (N_869,N_419,N_177);
or U870 (N_870,In_673,In_964);
nor U871 (N_871,In_1731,In_1700);
and U872 (N_872,N_548,N_771);
nand U873 (N_873,N_762,N_22);
and U874 (N_874,N_481,In_1927);
and U875 (N_875,In_927,N_552);
nand U876 (N_876,N_639,In_1517);
nor U877 (N_877,In_1597,In_201);
nand U878 (N_878,N_550,N_407);
nand U879 (N_879,N_608,In_446);
and U880 (N_880,In_332,N_433);
nand U881 (N_881,N_533,In_384);
nor U882 (N_882,In_1403,In_766);
or U883 (N_883,In_1933,In_1049);
nor U884 (N_884,N_675,In_1750);
nand U885 (N_885,N_129,In_317);
nor U886 (N_886,In_1133,N_744);
or U887 (N_887,N_405,N_773);
nand U888 (N_888,N_793,In_223);
or U889 (N_889,In_1218,N_514);
or U890 (N_890,In_1546,In_1264);
or U891 (N_891,N_500,In_1559);
or U892 (N_892,N_278,In_898);
nor U893 (N_893,N_619,In_33);
and U894 (N_894,N_797,In_86);
nand U895 (N_895,In_817,In_1552);
and U896 (N_896,N_360,N_588);
nand U897 (N_897,N_285,N_116);
and U898 (N_898,N_740,In_443);
nand U899 (N_899,In_1035,In_394);
nand U900 (N_900,N_277,N_451);
and U901 (N_901,N_783,N_579);
or U902 (N_902,N_545,N_710);
nand U903 (N_903,In_1239,N_565);
or U904 (N_904,In_568,In_870);
and U905 (N_905,In_1987,N_730);
nand U906 (N_906,In_1772,N_595);
nor U907 (N_907,In_6,N_18);
nor U908 (N_908,N_694,In_400);
xnor U909 (N_909,In_652,In_1896);
nand U910 (N_910,In_1279,N_787);
and U911 (N_911,N_346,In_379);
or U912 (N_912,In_1787,In_1373);
or U913 (N_913,In_1326,N_16);
nor U914 (N_914,In_435,N_457);
and U915 (N_915,In_1581,N_461);
or U916 (N_916,N_577,N_594);
and U917 (N_917,N_415,N_589);
or U918 (N_918,In_975,N_538);
and U919 (N_919,In_287,N_654);
and U920 (N_920,In_94,In_1357);
and U921 (N_921,N_593,In_179);
nand U922 (N_922,In_426,N_736);
or U923 (N_923,In_1163,N_422);
nor U924 (N_924,In_1594,N_279);
nor U925 (N_925,In_603,In_477);
or U926 (N_926,N_547,N_658);
and U927 (N_927,In_1673,In_761);
or U928 (N_928,In_536,N_570);
and U929 (N_929,N_445,N_350);
and U930 (N_930,In_1053,N_295);
nand U931 (N_931,N_779,N_248);
nor U932 (N_932,In_1745,N_590);
nand U933 (N_933,N_337,N_752);
or U934 (N_934,N_537,N_210);
xnor U935 (N_935,N_128,In_827);
or U936 (N_936,N_84,In_1685);
and U937 (N_937,In_1630,In_1767);
nor U938 (N_938,N_703,In_1267);
nor U939 (N_939,N_796,N_496);
xor U940 (N_940,N_791,N_157);
or U941 (N_941,In_1922,In_906);
nand U942 (N_942,In_717,N_782);
nand U943 (N_943,N_575,N_697);
and U944 (N_944,N_772,N_722);
nor U945 (N_945,N_247,In_173);
nand U946 (N_946,N_553,N_61);
and U947 (N_947,N_698,In_676);
nor U948 (N_948,N_598,In_1966);
nand U949 (N_949,N_580,In_1261);
nor U950 (N_950,N_409,N_723);
nor U951 (N_951,N_381,In_419);
and U952 (N_952,N_564,N_660);
and U953 (N_953,N_551,In_739);
nand U954 (N_954,N_705,In_1504);
or U955 (N_955,N_343,In_237);
nand U956 (N_956,In_816,In_39);
and U957 (N_957,In_912,In_153);
or U958 (N_958,N_420,In_1436);
nand U959 (N_959,In_1845,In_1228);
nand U960 (N_960,N_166,N_512);
nand U961 (N_961,In_928,In_1716);
nand U962 (N_962,In_1523,In_1438);
nand U963 (N_963,N_466,In_1967);
nor U964 (N_964,In_1942,N_386);
or U965 (N_965,In_780,N_532);
and U966 (N_966,In_1791,In_1044);
and U967 (N_967,In_109,In_293);
nand U968 (N_968,N_539,In_106);
or U969 (N_969,N_368,N_663);
and U970 (N_970,In_796,N_390);
or U971 (N_971,N_659,In_113);
nor U972 (N_972,N_592,In_1036);
or U973 (N_973,N_339,N_582);
nor U974 (N_974,In_11,N_437);
nand U975 (N_975,N_428,In_129);
and U976 (N_976,In_1843,N_743);
nor U977 (N_977,N_468,In_187);
and U978 (N_978,N_516,In_1994);
or U979 (N_979,N_574,N_633);
or U980 (N_980,N_497,N_404);
nor U981 (N_981,N_469,N_455);
nand U982 (N_982,N_674,In_89);
or U983 (N_983,In_393,N_125);
and U984 (N_984,In_280,In_271);
or U985 (N_985,N_212,N_213);
and U986 (N_986,In_23,In_1856);
or U987 (N_987,In_376,N_95);
and U988 (N_988,In_582,In_1104);
nand U989 (N_989,N_747,N_600);
nand U990 (N_990,In_1497,In_321);
nand U991 (N_991,N_766,In_1507);
nor U992 (N_992,N_370,N_299);
and U993 (N_993,N_106,N_29);
or U994 (N_994,N_645,In_1961);
nor U995 (N_995,N_556,In_1020);
or U996 (N_996,In_1406,N_449);
nor U997 (N_997,In_522,In_97);
and U998 (N_998,N_259,In_386);
and U999 (N_999,N_688,In_526);
or U1000 (N_1000,N_761,In_1598);
xnor U1001 (N_1001,N_140,N_444);
nor U1002 (N_1002,N_462,N_792);
and U1003 (N_1003,In_743,In_189);
nand U1004 (N_1004,N_701,In_395);
or U1005 (N_1005,In_484,N_392);
or U1006 (N_1006,In_1649,In_1717);
or U1007 (N_1007,In_1511,N_456);
or U1008 (N_1008,In_1965,In_1568);
and U1009 (N_1009,In_1655,N_156);
or U1010 (N_1010,In_581,N_764);
and U1011 (N_1011,N_572,In_1110);
or U1012 (N_1012,N_491,In_716);
nand U1013 (N_1013,In_269,In_1162);
or U1014 (N_1014,N_499,N_490);
or U1015 (N_1015,In_617,N_776);
nand U1016 (N_1016,In_1119,N_83);
nand U1017 (N_1017,N_518,N_502);
and U1018 (N_1018,N_146,N_648);
nand U1019 (N_1019,N_734,N_596);
nand U1020 (N_1020,N_721,N_424);
nor U1021 (N_1021,In_369,N_187);
and U1022 (N_1022,In_284,In_1854);
nor U1023 (N_1023,In_296,N_681);
or U1024 (N_1024,In_363,In_52);
or U1025 (N_1025,N_785,In_907);
nor U1026 (N_1026,In_940,In_132);
or U1027 (N_1027,In_1085,In_586);
nor U1028 (N_1028,In_1428,In_1602);
or U1029 (N_1029,N_513,N_450);
nor U1030 (N_1030,In_1661,N_618);
nand U1031 (N_1031,N_561,N_634);
or U1032 (N_1032,N_683,In_571);
and U1033 (N_1033,N_133,N_412);
nand U1034 (N_1034,In_10,In_21);
and U1035 (N_1035,N_421,In_548);
nor U1036 (N_1036,N_429,In_1270);
and U1037 (N_1037,In_1592,In_31);
nor U1038 (N_1038,In_1864,In_1906);
nor U1039 (N_1039,N_775,In_1093);
or U1040 (N_1040,In_770,N_714);
nor U1041 (N_1041,In_1947,N_642);
nand U1042 (N_1042,In_946,N_434);
or U1043 (N_1043,N_193,In_1751);
nand U1044 (N_1044,N_477,In_954);
and U1045 (N_1045,In_235,In_207);
nor U1046 (N_1046,In_1819,In_277);
nor U1047 (N_1047,N_770,In_534);
and U1048 (N_1048,In_1953,N_715);
and U1049 (N_1049,N_323,N_94);
and U1050 (N_1050,In_1675,In_1515);
or U1051 (N_1051,In_1643,In_618);
nand U1052 (N_1052,In_254,N_458);
or U1053 (N_1053,N_737,In_414);
nor U1054 (N_1054,In_1903,In_905);
and U1055 (N_1055,In_210,N_798);
and U1056 (N_1056,In_1291,N_320);
and U1057 (N_1057,In_84,N_265);
nand U1058 (N_1058,N_232,In_1611);
nor U1059 (N_1059,N_121,N_606);
or U1060 (N_1060,N_696,In_969);
or U1061 (N_1061,In_1667,In_630);
or U1062 (N_1062,In_1051,In_1835);
nand U1063 (N_1063,In_1410,N_41);
or U1064 (N_1064,In_131,N_283);
nand U1065 (N_1065,N_234,N_263);
nor U1066 (N_1066,N_330,In_952);
nand U1067 (N_1067,In_947,N_549);
and U1068 (N_1068,N_347,In_163);
nor U1069 (N_1069,N_371,In_505);
nor U1070 (N_1070,In_1820,In_1360);
or U1071 (N_1071,N_207,N_442);
and U1072 (N_1072,N_262,In_239);
and U1073 (N_1073,In_1202,N_340);
or U1074 (N_1074,In_139,N_253);
nand U1075 (N_1075,In_268,In_7);
or U1076 (N_1076,N_438,In_1883);
nand U1077 (N_1077,N_413,N_656);
or U1078 (N_1078,N_425,N_774);
and U1079 (N_1079,N_43,In_1310);
nand U1080 (N_1080,N_110,N_403);
or U1081 (N_1081,In_1531,N_795);
and U1082 (N_1082,N_290,In_1329);
nand U1083 (N_1083,In_1124,N_691);
nand U1084 (N_1084,N_2,In_1548);
nor U1085 (N_1085,In_496,N_467);
nand U1086 (N_1086,In_1077,N_401);
and U1087 (N_1087,In_272,In_1290);
nor U1088 (N_1088,N_788,N_643);
or U1089 (N_1089,N_599,In_120);
or U1090 (N_1090,N_759,In_1370);
or U1091 (N_1091,N_338,In_361);
and U1092 (N_1092,N_6,N_682);
or U1093 (N_1093,In_75,In_16);
nor U1094 (N_1094,In_1850,N_666);
and U1095 (N_1095,N_585,N_310);
nor U1096 (N_1096,N_416,In_605);
nor U1097 (N_1097,N_495,N_79);
nand U1098 (N_1098,N_249,N_389);
nand U1099 (N_1099,In_58,In_1072);
nand U1100 (N_1100,N_519,N_739);
and U1101 (N_1101,In_986,N_603);
and U1102 (N_1102,In_209,In_554);
and U1103 (N_1103,N_756,N_426);
and U1104 (N_1104,N_754,In_1606);
nand U1105 (N_1105,N_794,N_746);
or U1106 (N_1106,N_601,In_729);
and U1107 (N_1107,N_571,In_1502);
or U1108 (N_1108,N_32,In_1366);
or U1109 (N_1109,N_657,N_690);
nand U1110 (N_1110,N_0,N_704);
nand U1111 (N_1111,N_631,N_26);
and U1112 (N_1112,In_843,N_436);
nand U1113 (N_1113,N_71,In_1076);
or U1114 (N_1114,N_15,In_923);
nand U1115 (N_1115,In_742,In_222);
or U1116 (N_1116,In_532,N_214);
or U1117 (N_1117,N_183,In_1392);
and U1118 (N_1118,N_726,In_314);
nor U1119 (N_1119,In_205,In_498);
nand U1120 (N_1120,N_667,In_1840);
nor U1121 (N_1121,N_733,In_15);
nor U1122 (N_1122,N_484,N_289);
nor U1123 (N_1123,In_1473,N_612);
and U1124 (N_1124,In_1190,In_1158);
xnor U1125 (N_1125,In_1046,In_351);
and U1126 (N_1126,In_1244,In_29);
or U1127 (N_1127,N_126,N_482);
or U1128 (N_1128,N_208,In_521);
nand U1129 (N_1129,In_1260,N_661);
and U1130 (N_1130,In_1389,In_478);
xor U1131 (N_1131,N_607,In_865);
or U1132 (N_1132,In_175,N_57);
nand U1133 (N_1133,N_650,In_466);
nand U1134 (N_1134,In_87,In_672);
and U1135 (N_1135,N_486,N_717);
or U1136 (N_1136,N_363,In_1102);
and U1137 (N_1137,In_1539,N_742);
nor U1138 (N_1138,In_1610,In_1486);
nand U1139 (N_1139,In_171,In_374);
nor U1140 (N_1140,In_664,N_673);
nand U1141 (N_1141,In_1221,N_751);
nand U1142 (N_1142,N_382,In_1760);
and U1143 (N_1143,In_50,N_573);
nor U1144 (N_1144,N_554,N_1);
nor U1145 (N_1145,N_560,In_1336);
nor U1146 (N_1146,N_34,In_958);
or U1147 (N_1147,In_1982,In_1565);
nand U1148 (N_1148,N_69,N_613);
nor U1149 (N_1149,In_619,N_540);
or U1150 (N_1150,In_1726,In_8);
nor U1151 (N_1151,In_1855,In_551);
and U1152 (N_1152,In_1785,N_528);
and U1153 (N_1153,N_786,N_228);
nand U1154 (N_1154,N_732,N_760);
or U1155 (N_1155,N_508,N_70);
nor U1156 (N_1156,N_616,N_19);
xor U1157 (N_1157,In_1330,In_1802);
and U1158 (N_1158,In_570,N_719);
nor U1159 (N_1159,N_448,N_729);
nand U1160 (N_1160,N_42,N_521);
nor U1161 (N_1161,In_1828,N_627);
nand U1162 (N_1162,In_1624,N_636);
nand U1163 (N_1163,N_604,In_1446);
nand U1164 (N_1164,In_528,N_583);
and U1165 (N_1165,In_1981,In_1189);
and U1166 (N_1166,In_1460,In_647);
and U1167 (N_1167,N_559,N_624);
nand U1168 (N_1168,In_1980,In_24);
nor U1169 (N_1169,In_801,In_340);
nand U1170 (N_1170,N_120,N_546);
nor U1171 (N_1171,N_727,N_153);
and U1172 (N_1172,In_1962,In_1186);
nor U1173 (N_1173,In_1739,In_217);
nor U1174 (N_1174,In_416,In_1564);
nand U1175 (N_1175,In_19,N_738);
nor U1176 (N_1176,In_125,In_841);
and U1177 (N_1177,In_1280,N_647);
or U1178 (N_1178,In_253,In_845);
and U1179 (N_1179,In_1071,N_745);
or U1180 (N_1180,N_711,In_375);
nand U1181 (N_1181,N_446,In_76);
nand U1182 (N_1182,In_802,N_165);
nand U1183 (N_1183,In_934,In_177);
or U1184 (N_1184,N_640,N_602);
nand U1185 (N_1185,N_544,In_1355);
xnor U1186 (N_1186,N_748,In_3);
or U1187 (N_1187,In_438,In_245);
nand U1188 (N_1188,In_488,In_1634);
nor U1189 (N_1189,N_765,N_87);
nor U1190 (N_1190,N_220,N_473);
nor U1191 (N_1191,In_43,N_459);
nand U1192 (N_1192,N_584,N_431);
nand U1193 (N_1193,In_1430,In_1140);
nor U1194 (N_1194,N_778,N_378);
nand U1195 (N_1195,In_1089,In_1759);
or U1196 (N_1196,In_1048,N_186);
and U1197 (N_1197,N_758,In_1407);
nor U1198 (N_1198,In_596,N_50);
nand U1199 (N_1199,In_697,In_1263);
and U1200 (N_1200,N_1174,N_973);
nor U1201 (N_1201,N_838,N_839);
or U1202 (N_1202,N_395,N_932);
nand U1203 (N_1203,N_1182,N_1046);
or U1204 (N_1204,In_968,N_1193);
or U1205 (N_1205,In_1234,N_1167);
and U1206 (N_1206,In_1582,N_885);
and U1207 (N_1207,N_1161,In_112);
nand U1208 (N_1208,In_409,N_380);
nand U1209 (N_1209,N_479,N_231);
nor U1210 (N_1210,N_823,N_875);
or U1211 (N_1211,N_904,In_1007);
nor U1212 (N_1212,N_1191,N_641);
nor U1213 (N_1213,N_1151,N_909);
nand U1214 (N_1214,N_685,N_384);
or U1215 (N_1215,N_907,In_1737);
xnor U1216 (N_1216,N_1008,N_1055);
and U1217 (N_1217,N_928,N_881);
nor U1218 (N_1218,N_937,In_1480);
nand U1219 (N_1219,N_1024,In_1431);
nor U1220 (N_1220,N_510,N_1138);
nor U1221 (N_1221,In_486,In_854);
and U1222 (N_1222,N_977,N_969);
or U1223 (N_1223,N_995,N_1089);
or U1224 (N_1224,In_890,N_725);
nand U1225 (N_1225,In_736,In_1708);
xor U1226 (N_1226,N_817,In_529);
or U1227 (N_1227,N_938,N_465);
nand U1228 (N_1228,N_912,N_978);
and U1229 (N_1229,In_611,N_1054);
nor U1230 (N_1230,N_903,N_1118);
nor U1231 (N_1231,In_824,N_1137);
nor U1232 (N_1232,N_563,N_872);
nand U1233 (N_1233,N_913,N_718);
nor U1234 (N_1234,In_456,N_1015);
nand U1235 (N_1235,N_1153,N_1165);
or U1236 (N_1236,N_832,N_1183);
and U1237 (N_1237,N_1132,N_668);
nor U1238 (N_1238,N_845,N_443);
or U1239 (N_1239,N_789,N_1199);
nand U1240 (N_1240,N_811,N_522);
nand U1241 (N_1241,N_77,In_931);
nor U1242 (N_1242,In_1861,N_1068);
nor U1243 (N_1243,In_1519,N_1100);
and U1244 (N_1244,N_578,N_531);
or U1245 (N_1245,N_869,In_691);
or U1246 (N_1246,N_807,N_251);
or U1247 (N_1247,N_1123,N_952);
nor U1248 (N_1248,N_503,N_1041);
nor U1249 (N_1249,N_671,N_264);
or U1250 (N_1250,N_1017,In_389);
nor U1251 (N_1251,In_1340,N_954);
and U1252 (N_1252,In_1976,N_1131);
nor U1253 (N_1253,N_493,In_1579);
and U1254 (N_1254,N_111,N_1000);
or U1255 (N_1255,N_992,N_534);
or U1256 (N_1256,N_239,N_984);
and U1257 (N_1257,N_720,N_861);
or U1258 (N_1258,N_790,N_802);
or U1259 (N_1259,N_53,N_965);
or U1260 (N_1260,N_621,N_860);
and U1261 (N_1261,N_844,N_983);
nor U1262 (N_1262,N_892,N_1079);
and U1263 (N_1263,N_825,In_1417);
nor U1264 (N_1264,N_974,N_927);
nand U1265 (N_1265,N_649,N_142);
and U1266 (N_1266,N_1023,N_955);
nor U1267 (N_1267,In_930,N_506);
nor U1268 (N_1268,N_408,N_439);
nor U1269 (N_1269,N_853,N_1028);
nor U1270 (N_1270,N_1170,N_908);
nand U1271 (N_1271,In_1498,N_1053);
nor U1272 (N_1272,N_492,N_1064);
nor U1273 (N_1273,N_1177,N_741);
nor U1274 (N_1274,In_851,N_498);
nand U1275 (N_1275,N_847,In_1924);
nor U1276 (N_1276,N_255,In_342);
and U1277 (N_1277,In_1059,N_30);
nor U1278 (N_1278,N_399,N_402);
nand U1279 (N_1279,N_286,N_646);
or U1280 (N_1280,N_878,N_1065);
or U1281 (N_1281,N_1043,N_972);
nand U1282 (N_1282,N_406,N_74);
nand U1283 (N_1283,N_1021,N_1013);
nand U1284 (N_1284,N_1194,N_435);
nor U1285 (N_1285,N_1114,In_1788);
nor U1286 (N_1286,N_1172,N_1169);
nand U1287 (N_1287,In_1741,In_635);
and U1288 (N_1288,N_1038,N_924);
nor U1289 (N_1289,N_1142,In_1893);
and U1290 (N_1290,N_957,In_1616);
nand U1291 (N_1291,N_1012,N_195);
nand U1292 (N_1292,N_1075,In_1057);
and U1293 (N_1293,N_1003,N_910);
nor U1294 (N_1294,N_135,N_1102);
and U1295 (N_1295,In_45,N_669);
and U1296 (N_1296,In_918,In_889);
nand U1297 (N_1297,N_1173,N_1081);
nor U1298 (N_1298,In_1064,N_1139);
nor U1299 (N_1299,N_968,N_625);
nand U1300 (N_1300,In_1562,N_1148);
nand U1301 (N_1301,N_930,N_145);
and U1302 (N_1302,In_60,In_1092);
nand U1303 (N_1303,N_808,In_1206);
nand U1304 (N_1304,N_876,N_967);
and U1305 (N_1305,N_164,N_246);
or U1306 (N_1306,In_101,In_408);
nand U1307 (N_1307,N_781,In_1098);
or U1308 (N_1308,N_724,In_823);
nand U1309 (N_1309,In_1236,N_780);
and U1310 (N_1310,N_833,N_1163);
nand U1311 (N_1311,N_605,N_949);
xor U1312 (N_1312,In_1223,N_1022);
and U1313 (N_1313,N_945,In_591);
and U1314 (N_1314,In_447,N_329);
or U1315 (N_1315,N_1044,N_867);
or U1316 (N_1316,N_873,N_530);
nor U1317 (N_1317,In_329,In_1705);
nor U1318 (N_1318,N_919,N_917);
nor U1319 (N_1319,In_524,N_837);
and U1320 (N_1320,N_1002,In_810);
nand U1321 (N_1321,In_623,In_599);
nand U1322 (N_1322,In_1335,In_1090);
nand U1323 (N_1323,In_650,N_475);
nand U1324 (N_1324,N_1036,N_1164);
nor U1325 (N_1325,N_1074,N_1184);
or U1326 (N_1326,N_1066,In_1543);
xor U1327 (N_1327,N_1059,In_64);
or U1328 (N_1328,N_1185,N_679);
or U1329 (N_1329,N_1181,N_472);
or U1330 (N_1330,N_587,In_18);
and U1331 (N_1331,N_898,In_651);
and U1332 (N_1332,N_866,N_418);
and U1333 (N_1333,N_417,N_1005);
and U1334 (N_1334,N_1143,N_812);
nand U1335 (N_1335,N_880,In_781);
nand U1336 (N_1336,N_914,N_735);
nand U1337 (N_1337,N_480,N_1082);
and U1338 (N_1338,In_330,N_943);
or U1339 (N_1339,N_997,In_1042);
or U1340 (N_1340,N_947,N_1067);
nand U1341 (N_1341,N_855,N_81);
nor U1342 (N_1342,N_517,In_564);
nand U1343 (N_1343,N_1127,N_1166);
nand U1344 (N_1344,N_816,N_28);
nor U1345 (N_1345,N_653,N_1061);
and U1346 (N_1346,N_926,In_598);
or U1347 (N_1347,N_980,N_1162);
nand U1348 (N_1348,N_920,In_135);
and U1349 (N_1349,N_931,In_244);
nor U1350 (N_1350,N_98,N_182);
and U1351 (N_1351,N_268,In_572);
nand U1352 (N_1352,N_799,N_828);
and U1353 (N_1353,N_900,N_993);
nand U1354 (N_1354,N_644,N_1031);
and U1355 (N_1355,In_1521,N_1048);
and U1356 (N_1356,N_753,In_1157);
and U1357 (N_1357,N_1150,In_47);
nand U1358 (N_1358,N_996,In_1633);
or U1359 (N_1359,N_452,In_1301);
or U1360 (N_1360,N_1111,N_1032);
nor U1361 (N_1361,N_1176,In_491);
and U1362 (N_1362,N_304,N_941);
nor U1363 (N_1363,N_488,In_1713);
nor U1364 (N_1364,N_1129,N_411);
nor U1365 (N_1365,N_507,In_1269);
nand U1366 (N_1366,N_1035,N_1020);
or U1367 (N_1367,N_1069,N_929);
nand U1368 (N_1368,In_992,N_749);
and U1369 (N_1369,N_535,N_1198);
nand U1370 (N_1370,In_1769,N_767);
or U1371 (N_1371,N_948,N_902);
and U1372 (N_1372,N_483,In_273);
nor U1373 (N_1373,N_874,N_586);
nor U1374 (N_1374,N_999,N_1156);
and U1375 (N_1375,N_1146,N_906);
nand U1376 (N_1376,N_863,N_252);
and U1377 (N_1377,N_1103,N_815);
nor U1378 (N_1378,In_1660,N_1144);
and U1379 (N_1379,N_755,N_615);
xor U1380 (N_1380,N_1042,In_656);
nor U1381 (N_1381,In_152,N_470);
nand U1382 (N_1382,N_708,N_1030);
nand U1383 (N_1383,N_1196,N_865);
nand U1384 (N_1384,N_414,N_505);
nor U1385 (N_1385,N_944,N_1011);
and U1386 (N_1386,N_1107,N_291);
nor U1387 (N_1387,N_971,N_1158);
and U1388 (N_1388,N_1076,N_463);
nand U1389 (N_1389,N_1175,N_312);
and U1390 (N_1390,N_850,In_263);
nor U1391 (N_1391,N_1029,In_809);
and U1392 (N_1392,N_62,N_1094);
nor U1393 (N_1393,In_942,N_1039);
and U1394 (N_1394,In_410,N_1014);
nand U1395 (N_1395,In_190,In_397);
and U1396 (N_1396,N_400,N_1063);
or U1397 (N_1397,In_959,N_1168);
or U1398 (N_1398,N_897,N_950);
nor U1399 (N_1399,In_67,N_731);
and U1400 (N_1400,In_180,N_712);
nor U1401 (N_1401,N_64,N_620);
or U1402 (N_1402,N_464,N_1117);
and U1403 (N_1403,N_990,In_310);
nor U1404 (N_1404,N_901,N_357);
and U1405 (N_1405,N_515,In_1000);
nor U1406 (N_1406,N_1034,N_905);
nand U1407 (N_1407,N_1179,N_1159);
nor U1408 (N_1408,In_348,In_583);
and U1409 (N_1409,In_1070,N_713);
nand U1410 (N_1410,N_680,N_1120);
nor U1411 (N_1411,N_871,N_829);
or U1412 (N_1412,N_471,In_241);
nand U1413 (N_1413,In_595,N_822);
nand U1414 (N_1414,In_116,N_1147);
nand U1415 (N_1415,In_1094,In_380);
or U1416 (N_1416,N_1037,N_366);
or U1417 (N_1417,N_487,In_1192);
nor U1418 (N_1418,N_939,N_686);
or U1419 (N_1419,In_1061,N_963);
nor U1420 (N_1420,N_935,N_1180);
or U1421 (N_1421,N_888,In_1286);
nand U1422 (N_1422,In_785,N_824);
nor U1423 (N_1423,N_1084,N_810);
or U1424 (N_1424,N_555,N_365);
nand U1425 (N_1425,N_1124,N_527);
nand U1426 (N_1426,In_1174,N_1099);
nor U1427 (N_1427,N_1070,N_1026);
or U1428 (N_1428,In_1638,In_249);
or U1429 (N_1429,In_1795,N_868);
or U1430 (N_1430,In_1377,N_1091);
or U1431 (N_1431,In_1382,N_886);
nand U1432 (N_1432,N_292,N_1078);
nor U1433 (N_1433,N_1135,N_1009);
nand U1434 (N_1434,N_8,In_240);
or U1435 (N_1435,N_1056,N_523);
nand U1436 (N_1436,In_1659,N_56);
nor U1437 (N_1437,N_112,N_1050);
nand U1438 (N_1438,N_1128,N_849);
nor U1439 (N_1439,N_854,N_989);
nor U1440 (N_1440,N_830,In_341);
or U1441 (N_1441,N_1097,In_1273);
and U1442 (N_1442,N_1040,N_840);
or U1443 (N_1443,N_1087,N_706);
and U1444 (N_1444,In_1580,N_975);
or U1445 (N_1445,N_614,N_569);
nor U1446 (N_1446,N_1160,N_821);
and U1447 (N_1447,N_1007,In_1615);
nand U1448 (N_1448,N_1093,N_1071);
and U1449 (N_1449,N_1192,In_41);
or U1450 (N_1450,In_1457,N_956);
and U1451 (N_1451,N_635,N_826);
and U1452 (N_1452,In_899,N_117);
nor U1453 (N_1453,In_1063,N_1110);
nor U1454 (N_1454,N_662,N_842);
nand U1455 (N_1455,N_626,N_655);
or U1456 (N_1456,In_793,N_55);
and U1457 (N_1457,N_1133,N_1019);
nand U1458 (N_1458,In_1368,N_1086);
and U1459 (N_1459,N_925,In_686);
and U1460 (N_1460,In_585,In_692);
and U1461 (N_1461,N_1062,N_1113);
nand U1462 (N_1462,N_858,N_895);
xnor U1463 (N_1463,In_765,N_768);
or U1464 (N_1464,In_161,N_1058);
or U1465 (N_1465,N_889,N_806);
and U1466 (N_1466,N_1010,In_1415);
or U1467 (N_1467,In_891,N_131);
or U1468 (N_1468,In_42,In_1576);
nand U1469 (N_1469,In_1901,N_1027);
nand U1470 (N_1470,N_884,N_994);
and U1471 (N_1471,N_834,N_1109);
nor U1472 (N_1472,In_1184,N_1106);
and U1473 (N_1473,N_423,N_1154);
nand U1474 (N_1474,N_750,N_1045);
and U1475 (N_1475,N_820,N_1126);
and U1476 (N_1476,N_831,N_851);
and U1477 (N_1477,In_1621,N_818);
nand U1478 (N_1478,N_814,N_1073);
nand U1479 (N_1479,N_250,In_1525);
nor U1480 (N_1480,In_1275,In_121);
or U1481 (N_1481,In_501,N_911);
nand U1482 (N_1482,N_1096,N_809);
and U1483 (N_1483,N_9,N_813);
nand U1484 (N_1484,N_1001,N_716);
nor U1485 (N_1485,In_467,N_303);
nor U1486 (N_1486,N_1033,N_1018);
and U1487 (N_1487,N_835,N_763);
or U1488 (N_1488,N_672,N_962);
or U1489 (N_1489,N_1108,N_757);
nand U1490 (N_1490,N_852,N_1140);
or U1491 (N_1491,N_966,In_1354);
nor U1492 (N_1492,N_1105,In_1432);
and U1493 (N_1493,N_707,In_1823);
or U1494 (N_1494,N_887,N_1092);
nor U1495 (N_1495,N_1098,N_1047);
or U1496 (N_1496,N_652,In_1178);
and U1497 (N_1497,N_857,In_669);
or U1498 (N_1498,N_805,N_314);
or U1499 (N_1499,N_959,N_891);
nor U1500 (N_1500,N_1130,N_1145);
and U1501 (N_1501,N_987,N_942);
or U1502 (N_1502,N_1072,N_827);
nand U1503 (N_1503,In_1170,In_592);
or U1504 (N_1504,In_679,N_454);
nor U1505 (N_1505,N_1119,N_894);
nor U1506 (N_1506,N_923,N_1178);
nand U1507 (N_1507,N_960,In_1421);
nand U1508 (N_1508,N_566,N_14);
nor U1509 (N_1509,N_332,N_1189);
nand U1510 (N_1510,N_509,In_1888);
nand U1511 (N_1511,N_1049,N_864);
nor U1512 (N_1512,In_126,N_846);
nand U1513 (N_1513,N_1115,N_981);
or U1514 (N_1514,N_877,N_1141);
or U1515 (N_1515,N_976,N_856);
and U1516 (N_1516,In_1216,In_668);
or U1517 (N_1517,In_835,N_288);
nor U1518 (N_1518,In_1682,N_1134);
or U1519 (N_1519,N_921,N_1077);
or U1520 (N_1520,In_1934,N_364);
or U1521 (N_1521,In_1780,N_879);
nor U1522 (N_1522,N_1060,N_934);
nor U1523 (N_1523,N_670,N_1016);
nand U1524 (N_1524,N_524,N_447);
or U1525 (N_1525,N_638,N_1121);
and U1526 (N_1526,N_998,N_836);
or U1527 (N_1527,N_915,N_896);
nor U1528 (N_1528,N_1101,N_179);
and U1529 (N_1529,N_1171,N_841);
nor U1530 (N_1530,N_940,N_899);
nor U1531 (N_1531,In_1131,N_665);
and U1532 (N_1532,In_1282,N_353);
nor U1533 (N_1533,N_700,In_1825);
nor U1534 (N_1534,N_629,N_581);
nor U1535 (N_1535,N_1006,In_1816);
and U1536 (N_1536,N_1095,N_91);
and U1537 (N_1537,In_929,In_1866);
and U1538 (N_1538,In_1589,N_693);
nand U1539 (N_1539,In_1940,N_961);
nor U1540 (N_1540,N_1085,N_979);
and U1541 (N_1541,N_597,N_576);
nand U1542 (N_1542,N_617,N_1149);
and U1543 (N_1543,N_970,N_525);
and U1544 (N_1544,In_411,N_985);
and U1545 (N_1545,In_1095,N_933);
nor U1546 (N_1546,N_883,In_1365);
and U1547 (N_1547,In_1484,In_972);
nand U1548 (N_1548,N_804,N_843);
or U1549 (N_1549,In_797,In_1108);
or U1550 (N_1550,In_1574,N_893);
nand U1551 (N_1551,N_988,N_591);
nor U1552 (N_1552,N_803,N_1195);
and U1553 (N_1553,N_27,In_768);
nand U1554 (N_1554,N_1104,N_311);
nor U1555 (N_1555,In_1588,N_687);
nand U1556 (N_1556,N_986,N_953);
nor U1557 (N_1557,N_1051,In_1418);
nand U1558 (N_1558,N_23,N_1057);
or U1559 (N_1559,N_1136,N_676);
or U1560 (N_1560,N_1188,N_1186);
or U1561 (N_1561,N_1190,N_1155);
nand U1562 (N_1562,In_1187,In_828);
or U1563 (N_1563,N_1052,In_437);
nand U1564 (N_1564,In_537,In_1010);
and U1565 (N_1565,In_1241,N_922);
or U1566 (N_1566,N_982,In_540);
nor U1567 (N_1567,N_227,N_859);
nor U1568 (N_1568,N_1112,N_819);
nand U1569 (N_1569,N_326,N_1090);
and U1570 (N_1570,In_1526,N_784);
and U1571 (N_1571,N_558,In_1918);
or U1572 (N_1572,N_916,N_211);
nor U1573 (N_1573,N_964,N_504);
and U1574 (N_1574,N_946,N_936);
nor U1575 (N_1575,N_151,N_870);
nor U1576 (N_1576,N_325,N_862);
or U1577 (N_1577,N_313,N_678);
xor U1578 (N_1578,In_1604,N_39);
or U1579 (N_1579,N_1122,N_410);
nor U1580 (N_1580,N_991,In_316);
nor U1581 (N_1581,In_1601,N_1157);
and U1582 (N_1582,N_316,N_526);
and U1583 (N_1583,N_1083,N_951);
and U1584 (N_1584,N_890,N_1088);
and U1585 (N_1585,N_882,N_622);
nand U1586 (N_1586,N_958,In_219);
nor U1587 (N_1587,In_1494,In_886);
nand U1588 (N_1588,In_1642,N_801);
nor U1589 (N_1589,In_303,In_1420);
or U1590 (N_1590,In_1798,N_1080);
xnor U1591 (N_1591,In_288,In_1149);
nor U1592 (N_1592,N_1025,N_1116);
nand U1593 (N_1593,N_677,N_800);
nor U1594 (N_1594,N_848,N_1125);
or U1595 (N_1595,N_918,N_562);
nor U1596 (N_1596,In_98,In_775);
nor U1597 (N_1597,N_1004,N_1187);
nand U1598 (N_1598,N_1197,In_702);
and U1599 (N_1599,N_1152,In_1620);
nand U1600 (N_1600,N_1253,N_1312);
nor U1601 (N_1601,N_1328,N_1449);
nand U1602 (N_1602,N_1362,N_1550);
and U1603 (N_1603,N_1396,N_1557);
nand U1604 (N_1604,N_1528,N_1474);
or U1605 (N_1605,N_1233,N_1585);
and U1606 (N_1606,N_1464,N_1336);
nand U1607 (N_1607,N_1489,N_1547);
nor U1608 (N_1608,N_1433,N_1535);
or U1609 (N_1609,N_1333,N_1226);
and U1610 (N_1610,N_1217,N_1581);
nand U1611 (N_1611,N_1439,N_1324);
nor U1612 (N_1612,N_1279,N_1223);
or U1613 (N_1613,N_1388,N_1200);
nand U1614 (N_1614,N_1380,N_1509);
nand U1615 (N_1615,N_1569,N_1366);
or U1616 (N_1616,N_1554,N_1204);
nand U1617 (N_1617,N_1570,N_1292);
or U1618 (N_1618,N_1291,N_1227);
nand U1619 (N_1619,N_1351,N_1371);
and U1620 (N_1620,N_1390,N_1558);
or U1621 (N_1621,N_1468,N_1346);
or U1622 (N_1622,N_1453,N_1205);
or U1623 (N_1623,N_1481,N_1337);
and U1624 (N_1624,N_1465,N_1370);
nand U1625 (N_1625,N_1203,N_1286);
nand U1626 (N_1626,N_1424,N_1395);
or U1627 (N_1627,N_1445,N_1240);
nor U1628 (N_1628,N_1265,N_1207);
nand U1629 (N_1629,N_1456,N_1318);
and U1630 (N_1630,N_1272,N_1443);
nand U1631 (N_1631,N_1350,N_1477);
or U1632 (N_1632,N_1225,N_1364);
nor U1633 (N_1633,N_1495,N_1552);
and U1634 (N_1634,N_1410,N_1532);
nand U1635 (N_1635,N_1431,N_1210);
and U1636 (N_1636,N_1574,N_1549);
nor U1637 (N_1637,N_1471,N_1215);
nor U1638 (N_1638,N_1419,N_1485);
or U1639 (N_1639,N_1442,N_1510);
nand U1640 (N_1640,N_1482,N_1476);
and U1641 (N_1641,N_1266,N_1287);
nand U1642 (N_1642,N_1339,N_1421);
nor U1643 (N_1643,N_1296,N_1344);
or U1644 (N_1644,N_1457,N_1316);
nand U1645 (N_1645,N_1438,N_1459);
nor U1646 (N_1646,N_1248,N_1230);
nor U1647 (N_1647,N_1211,N_1347);
and U1648 (N_1648,N_1486,N_1277);
nand U1649 (N_1649,N_1497,N_1480);
nand U1650 (N_1650,N_1511,N_1377);
nand U1651 (N_1651,N_1586,N_1466);
nand U1652 (N_1652,N_1580,N_1450);
or U1653 (N_1653,N_1407,N_1490);
nor U1654 (N_1654,N_1461,N_1440);
nand U1655 (N_1655,N_1455,N_1268);
nand U1656 (N_1656,N_1437,N_1590);
and U1657 (N_1657,N_1209,N_1392);
and U1658 (N_1658,N_1251,N_1534);
nor U1659 (N_1659,N_1446,N_1417);
or U1660 (N_1660,N_1542,N_1246);
nor U1661 (N_1661,N_1262,N_1483);
and U1662 (N_1662,N_1237,N_1224);
nor U1663 (N_1663,N_1255,N_1214);
and U1664 (N_1664,N_1406,N_1228);
nand U1665 (N_1665,N_1294,N_1589);
nand U1666 (N_1666,N_1303,N_1353);
nor U1667 (N_1667,N_1555,N_1264);
and U1668 (N_1668,N_1413,N_1478);
and U1669 (N_1669,N_1208,N_1301);
or U1670 (N_1670,N_1512,N_1348);
and U1671 (N_1671,N_1447,N_1304);
nand U1672 (N_1672,N_1523,N_1288);
or U1673 (N_1673,N_1571,N_1222);
or U1674 (N_1674,N_1384,N_1520);
and U1675 (N_1675,N_1342,N_1427);
nand U1676 (N_1676,N_1565,N_1435);
nand U1677 (N_1677,N_1331,N_1531);
nor U1678 (N_1678,N_1411,N_1245);
and U1679 (N_1679,N_1373,N_1599);
or U1680 (N_1680,N_1561,N_1420);
or U1681 (N_1681,N_1545,N_1314);
nand U1682 (N_1682,N_1244,N_1235);
or U1683 (N_1683,N_1283,N_1398);
or U1684 (N_1684,N_1400,N_1359);
nor U1685 (N_1685,N_1361,N_1540);
and U1686 (N_1686,N_1521,N_1441);
or U1687 (N_1687,N_1281,N_1238);
nor U1688 (N_1688,N_1463,N_1573);
or U1689 (N_1689,N_1263,N_1280);
nand U1690 (N_1690,N_1556,N_1327);
nand U1691 (N_1691,N_1276,N_1267);
or U1692 (N_1692,N_1213,N_1454);
nor U1693 (N_1693,N_1541,N_1257);
nor U1694 (N_1694,N_1341,N_1340);
or U1695 (N_1695,N_1460,N_1484);
or U1696 (N_1696,N_1504,N_1412);
nor U1697 (N_1697,N_1502,N_1518);
nand U1698 (N_1698,N_1423,N_1329);
nand U1699 (N_1699,N_1335,N_1444);
nand U1700 (N_1700,N_1403,N_1382);
nor U1701 (N_1701,N_1221,N_1472);
nor U1702 (N_1702,N_1343,N_1315);
and U1703 (N_1703,N_1533,N_1234);
or U1704 (N_1704,N_1503,N_1306);
nand U1705 (N_1705,N_1448,N_1367);
and U1706 (N_1706,N_1241,N_1583);
nor U1707 (N_1707,N_1278,N_1313);
and U1708 (N_1708,N_1595,N_1259);
nand U1709 (N_1709,N_1297,N_1357);
and U1710 (N_1710,N_1321,N_1242);
nor U1711 (N_1711,N_1349,N_1404);
and U1712 (N_1712,N_1387,N_1516);
nor U1713 (N_1713,N_1527,N_1260);
or U1714 (N_1714,N_1338,N_1261);
nand U1715 (N_1715,N_1293,N_1475);
or U1716 (N_1716,N_1426,N_1269);
and U1717 (N_1717,N_1354,N_1469);
nor U1718 (N_1718,N_1491,N_1560);
and U1719 (N_1719,N_1375,N_1232);
or U1720 (N_1720,N_1524,N_1372);
nor U1721 (N_1721,N_1575,N_1365);
nand U1722 (N_1722,N_1325,N_1553);
nor U1723 (N_1723,N_1356,N_1492);
and U1724 (N_1724,N_1289,N_1270);
or U1725 (N_1725,N_1374,N_1308);
nand U1726 (N_1726,N_1572,N_1587);
and U1727 (N_1727,N_1479,N_1451);
nand U1728 (N_1728,N_1430,N_1525);
nand U1729 (N_1729,N_1501,N_1218);
and U1730 (N_1730,N_1548,N_1538);
nor U1731 (N_1731,N_1566,N_1529);
and U1732 (N_1732,N_1334,N_1236);
or U1733 (N_1733,N_1298,N_1513);
and U1734 (N_1734,N_1305,N_1559);
nand U1735 (N_1735,N_1567,N_1271);
or U1736 (N_1736,N_1402,N_1522);
nand U1737 (N_1737,N_1389,N_1307);
nor U1738 (N_1738,N_1473,N_1422);
or U1739 (N_1739,N_1526,N_1397);
nor U1740 (N_1740,N_1594,N_1216);
nand U1741 (N_1741,N_1386,N_1201);
or U1742 (N_1742,N_1418,N_1506);
or U1743 (N_1743,N_1425,N_1588);
or U1744 (N_1744,N_1332,N_1409);
nand U1745 (N_1745,N_1416,N_1578);
or U1746 (N_1746,N_1399,N_1243);
nand U1747 (N_1747,N_1393,N_1358);
or U1748 (N_1748,N_1536,N_1285);
and U1749 (N_1749,N_1428,N_1391);
nor U1750 (N_1750,N_1467,N_1546);
nor U1751 (N_1751,N_1385,N_1229);
nand U1752 (N_1752,N_1326,N_1470);
nor U1753 (N_1753,N_1597,N_1514);
nor U1754 (N_1754,N_1505,N_1345);
nand U1755 (N_1755,N_1408,N_1496);
or U1756 (N_1756,N_1352,N_1360);
or U1757 (N_1757,N_1564,N_1519);
and U1758 (N_1758,N_1487,N_1322);
nor U1759 (N_1759,N_1577,N_1551);
nor U1760 (N_1760,N_1537,N_1563);
or U1761 (N_1761,N_1330,N_1539);
or U1762 (N_1762,N_1414,N_1258);
or U1763 (N_1763,N_1282,N_1311);
and U1764 (N_1764,N_1517,N_1206);
and U1765 (N_1765,N_1247,N_1596);
and U1766 (N_1766,N_1317,N_1579);
nand U1767 (N_1767,N_1432,N_1436);
nand U1768 (N_1768,N_1295,N_1507);
xor U1769 (N_1769,N_1381,N_1256);
nand U1770 (N_1770,N_1591,N_1593);
and U1771 (N_1771,N_1320,N_1584);
nor U1772 (N_1772,N_1544,N_1202);
and U1773 (N_1773,N_1378,N_1290);
and U1774 (N_1774,N_1543,N_1394);
nor U1775 (N_1775,N_1250,N_1231);
and U1776 (N_1776,N_1458,N_1220);
or U1777 (N_1777,N_1530,N_1302);
and U1778 (N_1778,N_1415,N_1462);
nor U1779 (N_1779,N_1273,N_1434);
and U1780 (N_1780,N_1309,N_1452);
nor U1781 (N_1781,N_1252,N_1239);
nor U1782 (N_1782,N_1369,N_1568);
and U1783 (N_1783,N_1562,N_1368);
xnor U1784 (N_1784,N_1499,N_1401);
or U1785 (N_1785,N_1508,N_1249);
and U1786 (N_1786,N_1319,N_1488);
nor U1787 (N_1787,N_1254,N_1383);
and U1788 (N_1788,N_1515,N_1598);
nor U1789 (N_1789,N_1494,N_1299);
and U1790 (N_1790,N_1582,N_1493);
nand U1791 (N_1791,N_1363,N_1219);
and U1792 (N_1792,N_1275,N_1592);
or U1793 (N_1793,N_1310,N_1376);
and U1794 (N_1794,N_1300,N_1274);
xor U1795 (N_1795,N_1429,N_1379);
nand U1796 (N_1796,N_1284,N_1576);
nand U1797 (N_1797,N_1355,N_1323);
and U1798 (N_1798,N_1498,N_1405);
or U1799 (N_1799,N_1212,N_1500);
nand U1800 (N_1800,N_1541,N_1376);
or U1801 (N_1801,N_1503,N_1419);
or U1802 (N_1802,N_1493,N_1247);
or U1803 (N_1803,N_1595,N_1318);
nand U1804 (N_1804,N_1329,N_1522);
nor U1805 (N_1805,N_1442,N_1255);
and U1806 (N_1806,N_1235,N_1334);
or U1807 (N_1807,N_1346,N_1275);
nor U1808 (N_1808,N_1231,N_1211);
and U1809 (N_1809,N_1503,N_1591);
nand U1810 (N_1810,N_1574,N_1495);
and U1811 (N_1811,N_1556,N_1473);
nand U1812 (N_1812,N_1418,N_1306);
or U1813 (N_1813,N_1406,N_1201);
or U1814 (N_1814,N_1543,N_1551);
nor U1815 (N_1815,N_1419,N_1268);
nor U1816 (N_1816,N_1271,N_1407);
and U1817 (N_1817,N_1263,N_1407);
and U1818 (N_1818,N_1368,N_1464);
and U1819 (N_1819,N_1490,N_1554);
nor U1820 (N_1820,N_1439,N_1341);
and U1821 (N_1821,N_1308,N_1294);
and U1822 (N_1822,N_1294,N_1256);
nor U1823 (N_1823,N_1298,N_1563);
and U1824 (N_1824,N_1268,N_1279);
nand U1825 (N_1825,N_1540,N_1222);
and U1826 (N_1826,N_1538,N_1508);
and U1827 (N_1827,N_1248,N_1507);
nand U1828 (N_1828,N_1222,N_1594);
and U1829 (N_1829,N_1503,N_1299);
nor U1830 (N_1830,N_1390,N_1490);
and U1831 (N_1831,N_1491,N_1216);
and U1832 (N_1832,N_1498,N_1245);
nand U1833 (N_1833,N_1413,N_1306);
and U1834 (N_1834,N_1479,N_1208);
nand U1835 (N_1835,N_1528,N_1305);
and U1836 (N_1836,N_1438,N_1598);
or U1837 (N_1837,N_1475,N_1531);
nand U1838 (N_1838,N_1432,N_1369);
and U1839 (N_1839,N_1285,N_1560);
or U1840 (N_1840,N_1486,N_1296);
nor U1841 (N_1841,N_1216,N_1355);
and U1842 (N_1842,N_1390,N_1444);
and U1843 (N_1843,N_1584,N_1480);
nor U1844 (N_1844,N_1562,N_1526);
nor U1845 (N_1845,N_1222,N_1498);
nor U1846 (N_1846,N_1481,N_1433);
nand U1847 (N_1847,N_1506,N_1431);
nand U1848 (N_1848,N_1528,N_1459);
and U1849 (N_1849,N_1407,N_1288);
and U1850 (N_1850,N_1410,N_1315);
nor U1851 (N_1851,N_1599,N_1501);
nor U1852 (N_1852,N_1533,N_1212);
xor U1853 (N_1853,N_1214,N_1368);
and U1854 (N_1854,N_1314,N_1587);
nand U1855 (N_1855,N_1326,N_1217);
nand U1856 (N_1856,N_1587,N_1288);
or U1857 (N_1857,N_1486,N_1386);
nand U1858 (N_1858,N_1393,N_1430);
nand U1859 (N_1859,N_1439,N_1426);
and U1860 (N_1860,N_1238,N_1442);
nor U1861 (N_1861,N_1551,N_1538);
and U1862 (N_1862,N_1352,N_1366);
or U1863 (N_1863,N_1489,N_1314);
and U1864 (N_1864,N_1541,N_1252);
nand U1865 (N_1865,N_1583,N_1429);
nand U1866 (N_1866,N_1455,N_1232);
or U1867 (N_1867,N_1475,N_1593);
or U1868 (N_1868,N_1452,N_1474);
nand U1869 (N_1869,N_1553,N_1409);
nor U1870 (N_1870,N_1271,N_1266);
or U1871 (N_1871,N_1421,N_1280);
or U1872 (N_1872,N_1449,N_1386);
and U1873 (N_1873,N_1224,N_1375);
or U1874 (N_1874,N_1499,N_1254);
nand U1875 (N_1875,N_1249,N_1510);
or U1876 (N_1876,N_1326,N_1238);
or U1877 (N_1877,N_1396,N_1376);
and U1878 (N_1878,N_1378,N_1279);
or U1879 (N_1879,N_1568,N_1519);
or U1880 (N_1880,N_1348,N_1541);
nor U1881 (N_1881,N_1287,N_1216);
or U1882 (N_1882,N_1399,N_1431);
and U1883 (N_1883,N_1594,N_1341);
and U1884 (N_1884,N_1517,N_1491);
nand U1885 (N_1885,N_1481,N_1541);
nand U1886 (N_1886,N_1500,N_1275);
or U1887 (N_1887,N_1405,N_1408);
nand U1888 (N_1888,N_1200,N_1466);
and U1889 (N_1889,N_1525,N_1245);
and U1890 (N_1890,N_1260,N_1291);
and U1891 (N_1891,N_1269,N_1309);
nand U1892 (N_1892,N_1396,N_1251);
and U1893 (N_1893,N_1236,N_1309);
nor U1894 (N_1894,N_1221,N_1396);
nor U1895 (N_1895,N_1592,N_1427);
nand U1896 (N_1896,N_1423,N_1410);
and U1897 (N_1897,N_1569,N_1591);
or U1898 (N_1898,N_1429,N_1459);
and U1899 (N_1899,N_1291,N_1353);
or U1900 (N_1900,N_1435,N_1498);
or U1901 (N_1901,N_1289,N_1408);
and U1902 (N_1902,N_1488,N_1442);
nand U1903 (N_1903,N_1404,N_1485);
or U1904 (N_1904,N_1563,N_1246);
or U1905 (N_1905,N_1555,N_1521);
or U1906 (N_1906,N_1338,N_1310);
and U1907 (N_1907,N_1325,N_1552);
nor U1908 (N_1908,N_1455,N_1496);
nor U1909 (N_1909,N_1502,N_1327);
or U1910 (N_1910,N_1377,N_1305);
and U1911 (N_1911,N_1590,N_1535);
nand U1912 (N_1912,N_1369,N_1297);
nor U1913 (N_1913,N_1257,N_1341);
nor U1914 (N_1914,N_1540,N_1300);
or U1915 (N_1915,N_1326,N_1581);
and U1916 (N_1916,N_1294,N_1345);
and U1917 (N_1917,N_1219,N_1507);
or U1918 (N_1918,N_1384,N_1282);
nand U1919 (N_1919,N_1332,N_1436);
or U1920 (N_1920,N_1433,N_1379);
and U1921 (N_1921,N_1305,N_1466);
nor U1922 (N_1922,N_1364,N_1401);
nand U1923 (N_1923,N_1399,N_1565);
nand U1924 (N_1924,N_1366,N_1444);
nand U1925 (N_1925,N_1313,N_1205);
nor U1926 (N_1926,N_1323,N_1212);
nor U1927 (N_1927,N_1476,N_1474);
nand U1928 (N_1928,N_1574,N_1205);
nand U1929 (N_1929,N_1521,N_1334);
or U1930 (N_1930,N_1284,N_1593);
nand U1931 (N_1931,N_1225,N_1205);
and U1932 (N_1932,N_1436,N_1276);
nor U1933 (N_1933,N_1528,N_1258);
and U1934 (N_1934,N_1212,N_1530);
nor U1935 (N_1935,N_1201,N_1539);
nor U1936 (N_1936,N_1591,N_1370);
nor U1937 (N_1937,N_1208,N_1363);
or U1938 (N_1938,N_1512,N_1235);
nor U1939 (N_1939,N_1244,N_1252);
nand U1940 (N_1940,N_1415,N_1208);
and U1941 (N_1941,N_1502,N_1477);
or U1942 (N_1942,N_1309,N_1299);
or U1943 (N_1943,N_1508,N_1539);
or U1944 (N_1944,N_1590,N_1561);
nor U1945 (N_1945,N_1356,N_1564);
and U1946 (N_1946,N_1514,N_1211);
and U1947 (N_1947,N_1309,N_1336);
nor U1948 (N_1948,N_1475,N_1218);
nor U1949 (N_1949,N_1201,N_1554);
nor U1950 (N_1950,N_1336,N_1476);
and U1951 (N_1951,N_1393,N_1571);
nand U1952 (N_1952,N_1332,N_1478);
and U1953 (N_1953,N_1284,N_1224);
and U1954 (N_1954,N_1399,N_1463);
or U1955 (N_1955,N_1299,N_1566);
nand U1956 (N_1956,N_1474,N_1361);
nand U1957 (N_1957,N_1598,N_1335);
and U1958 (N_1958,N_1456,N_1495);
nor U1959 (N_1959,N_1480,N_1245);
and U1960 (N_1960,N_1507,N_1243);
nor U1961 (N_1961,N_1309,N_1463);
nand U1962 (N_1962,N_1482,N_1383);
nor U1963 (N_1963,N_1527,N_1347);
nand U1964 (N_1964,N_1497,N_1265);
or U1965 (N_1965,N_1376,N_1494);
nor U1966 (N_1966,N_1581,N_1342);
xor U1967 (N_1967,N_1445,N_1468);
nand U1968 (N_1968,N_1592,N_1517);
nor U1969 (N_1969,N_1466,N_1318);
nand U1970 (N_1970,N_1476,N_1343);
and U1971 (N_1971,N_1332,N_1230);
and U1972 (N_1972,N_1227,N_1220);
and U1973 (N_1973,N_1598,N_1347);
nor U1974 (N_1974,N_1500,N_1502);
and U1975 (N_1975,N_1338,N_1275);
and U1976 (N_1976,N_1510,N_1416);
and U1977 (N_1977,N_1500,N_1305);
and U1978 (N_1978,N_1542,N_1363);
or U1979 (N_1979,N_1491,N_1382);
and U1980 (N_1980,N_1333,N_1430);
or U1981 (N_1981,N_1353,N_1462);
and U1982 (N_1982,N_1254,N_1341);
nor U1983 (N_1983,N_1560,N_1344);
nand U1984 (N_1984,N_1471,N_1320);
or U1985 (N_1985,N_1214,N_1514);
nand U1986 (N_1986,N_1236,N_1336);
xor U1987 (N_1987,N_1516,N_1273);
nor U1988 (N_1988,N_1207,N_1569);
or U1989 (N_1989,N_1495,N_1306);
nand U1990 (N_1990,N_1526,N_1275);
nand U1991 (N_1991,N_1471,N_1370);
or U1992 (N_1992,N_1578,N_1310);
nand U1993 (N_1993,N_1463,N_1495);
or U1994 (N_1994,N_1235,N_1560);
or U1995 (N_1995,N_1239,N_1412);
and U1996 (N_1996,N_1407,N_1536);
nor U1997 (N_1997,N_1208,N_1388);
or U1998 (N_1998,N_1363,N_1355);
or U1999 (N_1999,N_1480,N_1318);
and U2000 (N_2000,N_1869,N_1894);
and U2001 (N_2001,N_1750,N_1952);
nor U2002 (N_2002,N_1852,N_1886);
and U2003 (N_2003,N_1999,N_1627);
xor U2004 (N_2004,N_1845,N_1936);
or U2005 (N_2005,N_1955,N_1951);
or U2006 (N_2006,N_1910,N_1707);
or U2007 (N_2007,N_1601,N_1621);
nand U2008 (N_2008,N_1946,N_1904);
and U2009 (N_2009,N_1823,N_1629);
or U2010 (N_2010,N_1625,N_1934);
or U2011 (N_2011,N_1930,N_1853);
and U2012 (N_2012,N_1984,N_1828);
or U2013 (N_2013,N_1826,N_1652);
nand U2014 (N_2014,N_1972,N_1892);
or U2015 (N_2015,N_1770,N_1696);
nand U2016 (N_2016,N_1835,N_1643);
nor U2017 (N_2017,N_1772,N_1925);
and U2018 (N_2018,N_1906,N_1868);
nand U2019 (N_2019,N_1626,N_1965);
nor U2020 (N_2020,N_1725,N_1606);
nand U2021 (N_2021,N_1854,N_1807);
and U2022 (N_2022,N_1657,N_1690);
or U2023 (N_2023,N_1858,N_1661);
nand U2024 (N_2024,N_1633,N_1797);
nand U2025 (N_2025,N_1743,N_1648);
nor U2026 (N_2026,N_1677,N_1664);
nor U2027 (N_2027,N_1703,N_1686);
nor U2028 (N_2028,N_1775,N_1866);
nand U2029 (N_2029,N_1982,N_1610);
nor U2030 (N_2030,N_1956,N_1628);
or U2031 (N_2031,N_1996,N_1747);
or U2032 (N_2032,N_1717,N_1815);
nand U2033 (N_2033,N_1758,N_1658);
nor U2034 (N_2034,N_1809,N_1801);
nor U2035 (N_2035,N_1619,N_1979);
nor U2036 (N_2036,N_1649,N_1630);
or U2037 (N_2037,N_1695,N_1613);
and U2038 (N_2038,N_1931,N_1611);
and U2039 (N_2039,N_1709,N_1671);
nor U2040 (N_2040,N_1924,N_1644);
or U2041 (N_2041,N_1986,N_1769);
and U2042 (N_2042,N_1957,N_1918);
or U2043 (N_2043,N_1800,N_1660);
nand U2044 (N_2044,N_1867,N_1898);
nor U2045 (N_2045,N_1961,N_1950);
nor U2046 (N_2046,N_1719,N_1773);
nand U2047 (N_2047,N_1687,N_1749);
nor U2048 (N_2048,N_1865,N_1897);
nand U2049 (N_2049,N_1776,N_1871);
nand U2050 (N_2050,N_1953,N_1857);
and U2051 (N_2051,N_1909,N_1884);
and U2052 (N_2052,N_1939,N_1663);
and U2053 (N_2053,N_1819,N_1942);
or U2054 (N_2054,N_1900,N_1820);
nand U2055 (N_2055,N_1974,N_1822);
and U2056 (N_2056,N_1976,N_1937);
nor U2057 (N_2057,N_1877,N_1981);
and U2058 (N_2058,N_1759,N_1740);
or U2059 (N_2059,N_1736,N_1881);
nand U2060 (N_2060,N_1783,N_1825);
nor U2061 (N_2061,N_1989,N_1899);
or U2062 (N_2062,N_1795,N_1700);
and U2063 (N_2063,N_1812,N_1798);
nand U2064 (N_2064,N_1844,N_1762);
or U2065 (N_2065,N_1802,N_1907);
nor U2066 (N_2066,N_1699,N_1689);
nor U2067 (N_2067,N_1622,N_1817);
and U2068 (N_2068,N_1905,N_1755);
or U2069 (N_2069,N_1679,N_1751);
and U2070 (N_2070,N_1896,N_1855);
nor U2071 (N_2071,N_1670,N_1941);
or U2072 (N_2072,N_1968,N_1742);
nor U2073 (N_2073,N_1814,N_1882);
or U2074 (N_2074,N_1843,N_1718);
nor U2075 (N_2075,N_1832,N_1641);
or U2076 (N_2076,N_1779,N_1875);
or U2077 (N_2077,N_1752,N_1685);
or U2078 (N_2078,N_1929,N_1923);
and U2079 (N_2079,N_1889,N_1806);
nand U2080 (N_2080,N_1603,N_1908);
or U2081 (N_2081,N_1724,N_1993);
nand U2082 (N_2082,N_1780,N_1727);
nor U2083 (N_2083,N_1980,N_1827);
nor U2084 (N_2084,N_1694,N_1919);
and U2085 (N_2085,N_1805,N_1933);
nor U2086 (N_2086,N_1721,N_1616);
or U2087 (N_2087,N_1850,N_1983);
or U2088 (N_2088,N_1997,N_1840);
nand U2089 (N_2089,N_1863,N_1665);
nand U2090 (N_2090,N_1708,N_1682);
or U2091 (N_2091,N_1970,N_1922);
and U2092 (N_2092,N_1887,N_1761);
and U2093 (N_2093,N_1861,N_1739);
nor U2094 (N_2094,N_1796,N_1655);
nand U2095 (N_2095,N_1821,N_1794);
nor U2096 (N_2096,N_1778,N_1920);
and U2097 (N_2097,N_1977,N_1673);
or U2098 (N_2098,N_1711,N_1693);
nor U2099 (N_2099,N_1640,N_1716);
and U2100 (N_2100,N_1880,N_1790);
and U2101 (N_2101,N_1870,N_1838);
nor U2102 (N_2102,N_1831,N_1876);
nor U2103 (N_2103,N_1701,N_1672);
nor U2104 (N_2104,N_1962,N_1959);
and U2105 (N_2105,N_1834,N_1813);
nor U2106 (N_2106,N_1726,N_1833);
nor U2107 (N_2107,N_1960,N_1932);
nand U2108 (N_2108,N_1615,N_1782);
and U2109 (N_2109,N_1729,N_1777);
nor U2110 (N_2110,N_1624,N_1781);
nand U2111 (N_2111,N_1768,N_1738);
and U2112 (N_2112,N_1653,N_1816);
or U2113 (N_2113,N_1666,N_1713);
nor U2114 (N_2114,N_1681,N_1872);
and U2115 (N_2115,N_1901,N_1964);
and U2116 (N_2116,N_1784,N_1792);
or U2117 (N_2117,N_1785,N_1985);
and U2118 (N_2118,N_1893,N_1935);
nor U2119 (N_2119,N_1787,N_1618);
and U2120 (N_2120,N_1754,N_1642);
nor U2121 (N_2121,N_1885,N_1839);
nor U2122 (N_2122,N_1760,N_1915);
and U2123 (N_2123,N_1654,N_1745);
or U2124 (N_2124,N_1966,N_1911);
nand U2125 (N_2125,N_1938,N_1766);
nor U2126 (N_2126,N_1978,N_1879);
or U2127 (N_2127,N_1650,N_1757);
nand U2128 (N_2128,N_1600,N_1829);
nor U2129 (N_2129,N_1969,N_1891);
nor U2130 (N_2130,N_1948,N_1712);
and U2131 (N_2131,N_1926,N_1680);
or U2132 (N_2132,N_1667,N_1612);
nand U2133 (N_2133,N_1856,N_1967);
and U2134 (N_2134,N_1748,N_1646);
nand U2135 (N_2135,N_1958,N_1842);
nand U2136 (N_2136,N_1697,N_1702);
or U2137 (N_2137,N_1676,N_1921);
nand U2138 (N_2138,N_1710,N_1744);
nor U2139 (N_2139,N_1678,N_1620);
nor U2140 (N_2140,N_1927,N_1987);
and U2141 (N_2141,N_1846,N_1604);
or U2142 (N_2142,N_1753,N_1991);
nand U2143 (N_2143,N_1763,N_1940);
and U2144 (N_2144,N_1995,N_1684);
and U2145 (N_2145,N_1674,N_1912);
nor U2146 (N_2146,N_1733,N_1722);
nand U2147 (N_2147,N_1659,N_1614);
nand U2148 (N_2148,N_1998,N_1810);
or U2149 (N_2149,N_1902,N_1990);
nor U2150 (N_2150,N_1849,N_1811);
nor U2151 (N_2151,N_1799,N_1988);
nor U2152 (N_2152,N_1949,N_1714);
nor U2153 (N_2153,N_1698,N_1669);
nor U2154 (N_2154,N_1691,N_1851);
nand U2155 (N_2155,N_1635,N_1994);
or U2156 (N_2156,N_1728,N_1883);
and U2157 (N_2157,N_1947,N_1859);
or U2158 (N_2158,N_1803,N_1715);
or U2159 (N_2159,N_1609,N_1786);
nor U2160 (N_2160,N_1656,N_1765);
nor U2161 (N_2161,N_1645,N_1605);
and U2162 (N_2162,N_1841,N_1632);
and U2163 (N_2163,N_1992,N_1862);
and U2164 (N_2164,N_1873,N_1623);
or U2165 (N_2165,N_1639,N_1975);
nand U2166 (N_2166,N_1737,N_1874);
or U2167 (N_2167,N_1963,N_1848);
nand U2168 (N_2168,N_1973,N_1914);
nand U2169 (N_2169,N_1651,N_1818);
nor U2170 (N_2170,N_1830,N_1608);
nand U2171 (N_2171,N_1636,N_1789);
nand U2172 (N_2172,N_1662,N_1732);
nand U2173 (N_2173,N_1771,N_1735);
and U2174 (N_2174,N_1746,N_1836);
xnor U2175 (N_2175,N_1824,N_1878);
nor U2176 (N_2176,N_1734,N_1890);
or U2177 (N_2177,N_1617,N_1647);
and U2178 (N_2178,N_1631,N_1704);
and U2179 (N_2179,N_1637,N_1788);
nand U2180 (N_2180,N_1607,N_1638);
and U2181 (N_2181,N_1971,N_1723);
nor U2182 (N_2182,N_1943,N_1913);
and U2183 (N_2183,N_1764,N_1804);
and U2184 (N_2184,N_1688,N_1675);
or U2185 (N_2185,N_1916,N_1895);
nand U2186 (N_2186,N_1767,N_1706);
and U2187 (N_2187,N_1720,N_1847);
and U2188 (N_2188,N_1954,N_1668);
and U2189 (N_2189,N_1837,N_1864);
and U2190 (N_2190,N_1741,N_1756);
nand U2191 (N_2191,N_1903,N_1705);
nor U2192 (N_2192,N_1944,N_1692);
or U2193 (N_2193,N_1730,N_1683);
nor U2194 (N_2194,N_1945,N_1791);
and U2195 (N_2195,N_1602,N_1888);
nand U2196 (N_2196,N_1634,N_1774);
or U2197 (N_2197,N_1793,N_1731);
nor U2198 (N_2198,N_1917,N_1860);
nand U2199 (N_2199,N_1928,N_1808);
nand U2200 (N_2200,N_1761,N_1838);
nand U2201 (N_2201,N_1652,N_1600);
or U2202 (N_2202,N_1976,N_1987);
or U2203 (N_2203,N_1840,N_1973);
and U2204 (N_2204,N_1965,N_1673);
or U2205 (N_2205,N_1846,N_1784);
and U2206 (N_2206,N_1951,N_1917);
and U2207 (N_2207,N_1925,N_1659);
or U2208 (N_2208,N_1850,N_1832);
nor U2209 (N_2209,N_1975,N_1659);
and U2210 (N_2210,N_1620,N_1806);
or U2211 (N_2211,N_1707,N_1601);
nor U2212 (N_2212,N_1983,N_1941);
xnor U2213 (N_2213,N_1672,N_1644);
or U2214 (N_2214,N_1624,N_1822);
and U2215 (N_2215,N_1658,N_1791);
xnor U2216 (N_2216,N_1934,N_1854);
or U2217 (N_2217,N_1907,N_1969);
and U2218 (N_2218,N_1960,N_1726);
nand U2219 (N_2219,N_1762,N_1979);
nor U2220 (N_2220,N_1622,N_1963);
nor U2221 (N_2221,N_1884,N_1981);
or U2222 (N_2222,N_1990,N_1852);
nor U2223 (N_2223,N_1674,N_1638);
nor U2224 (N_2224,N_1615,N_1756);
nor U2225 (N_2225,N_1881,N_1691);
nand U2226 (N_2226,N_1890,N_1899);
nor U2227 (N_2227,N_1705,N_1614);
and U2228 (N_2228,N_1923,N_1850);
and U2229 (N_2229,N_1906,N_1675);
nor U2230 (N_2230,N_1667,N_1753);
or U2231 (N_2231,N_1962,N_1740);
and U2232 (N_2232,N_1648,N_1902);
nor U2233 (N_2233,N_1728,N_1956);
nor U2234 (N_2234,N_1946,N_1827);
and U2235 (N_2235,N_1932,N_1979);
nand U2236 (N_2236,N_1746,N_1626);
nand U2237 (N_2237,N_1861,N_1853);
and U2238 (N_2238,N_1795,N_1764);
nor U2239 (N_2239,N_1983,N_1633);
and U2240 (N_2240,N_1774,N_1708);
or U2241 (N_2241,N_1809,N_1707);
and U2242 (N_2242,N_1737,N_1713);
nor U2243 (N_2243,N_1687,N_1667);
nand U2244 (N_2244,N_1831,N_1937);
nand U2245 (N_2245,N_1900,N_1854);
nand U2246 (N_2246,N_1719,N_1943);
nand U2247 (N_2247,N_1808,N_1745);
and U2248 (N_2248,N_1737,N_1832);
xor U2249 (N_2249,N_1873,N_1990);
xor U2250 (N_2250,N_1785,N_1661);
or U2251 (N_2251,N_1737,N_1656);
nand U2252 (N_2252,N_1909,N_1863);
or U2253 (N_2253,N_1744,N_1685);
nand U2254 (N_2254,N_1627,N_1814);
nand U2255 (N_2255,N_1992,N_1919);
and U2256 (N_2256,N_1630,N_1623);
or U2257 (N_2257,N_1859,N_1899);
nor U2258 (N_2258,N_1933,N_1986);
nand U2259 (N_2259,N_1647,N_1815);
or U2260 (N_2260,N_1943,N_1692);
nand U2261 (N_2261,N_1933,N_1608);
nand U2262 (N_2262,N_1980,N_1955);
and U2263 (N_2263,N_1854,N_1811);
and U2264 (N_2264,N_1716,N_1940);
and U2265 (N_2265,N_1611,N_1631);
and U2266 (N_2266,N_1758,N_1779);
or U2267 (N_2267,N_1787,N_1765);
nor U2268 (N_2268,N_1827,N_1729);
and U2269 (N_2269,N_1962,N_1721);
or U2270 (N_2270,N_1782,N_1967);
nor U2271 (N_2271,N_1933,N_1771);
or U2272 (N_2272,N_1971,N_1621);
nand U2273 (N_2273,N_1685,N_1865);
or U2274 (N_2274,N_1611,N_1654);
or U2275 (N_2275,N_1659,N_1847);
and U2276 (N_2276,N_1748,N_1610);
nor U2277 (N_2277,N_1680,N_1646);
and U2278 (N_2278,N_1849,N_1779);
or U2279 (N_2279,N_1670,N_1868);
nand U2280 (N_2280,N_1710,N_1664);
nand U2281 (N_2281,N_1759,N_1905);
or U2282 (N_2282,N_1607,N_1787);
and U2283 (N_2283,N_1757,N_1709);
and U2284 (N_2284,N_1792,N_1626);
and U2285 (N_2285,N_1712,N_1964);
and U2286 (N_2286,N_1679,N_1610);
nor U2287 (N_2287,N_1946,N_1703);
nand U2288 (N_2288,N_1600,N_1801);
xor U2289 (N_2289,N_1994,N_1639);
and U2290 (N_2290,N_1634,N_1838);
or U2291 (N_2291,N_1829,N_1896);
or U2292 (N_2292,N_1862,N_1930);
nor U2293 (N_2293,N_1750,N_1869);
nand U2294 (N_2294,N_1620,N_1936);
and U2295 (N_2295,N_1800,N_1798);
nor U2296 (N_2296,N_1663,N_1664);
or U2297 (N_2297,N_1642,N_1636);
nand U2298 (N_2298,N_1831,N_1852);
nand U2299 (N_2299,N_1904,N_1779);
nor U2300 (N_2300,N_1857,N_1790);
nor U2301 (N_2301,N_1743,N_1871);
nor U2302 (N_2302,N_1602,N_1662);
nand U2303 (N_2303,N_1746,N_1806);
nand U2304 (N_2304,N_1785,N_1698);
nand U2305 (N_2305,N_1954,N_1826);
or U2306 (N_2306,N_1629,N_1609);
nor U2307 (N_2307,N_1758,N_1641);
or U2308 (N_2308,N_1681,N_1956);
nand U2309 (N_2309,N_1711,N_1747);
nand U2310 (N_2310,N_1904,N_1662);
nor U2311 (N_2311,N_1883,N_1738);
and U2312 (N_2312,N_1721,N_1708);
nand U2313 (N_2313,N_1825,N_1638);
or U2314 (N_2314,N_1759,N_1776);
and U2315 (N_2315,N_1987,N_1839);
nand U2316 (N_2316,N_1637,N_1995);
nand U2317 (N_2317,N_1825,N_1974);
nor U2318 (N_2318,N_1962,N_1668);
nor U2319 (N_2319,N_1885,N_1761);
or U2320 (N_2320,N_1682,N_1607);
or U2321 (N_2321,N_1949,N_1882);
or U2322 (N_2322,N_1875,N_1815);
and U2323 (N_2323,N_1698,N_1994);
nor U2324 (N_2324,N_1760,N_1784);
xor U2325 (N_2325,N_1756,N_1910);
or U2326 (N_2326,N_1771,N_1876);
and U2327 (N_2327,N_1888,N_1841);
nor U2328 (N_2328,N_1939,N_1679);
and U2329 (N_2329,N_1781,N_1879);
nand U2330 (N_2330,N_1667,N_1979);
and U2331 (N_2331,N_1814,N_1862);
or U2332 (N_2332,N_1813,N_1600);
nor U2333 (N_2333,N_1718,N_1930);
and U2334 (N_2334,N_1718,N_1918);
nand U2335 (N_2335,N_1768,N_1866);
nand U2336 (N_2336,N_1952,N_1998);
nand U2337 (N_2337,N_1605,N_1930);
nor U2338 (N_2338,N_1710,N_1919);
or U2339 (N_2339,N_1829,N_1768);
and U2340 (N_2340,N_1672,N_1799);
or U2341 (N_2341,N_1848,N_1788);
nand U2342 (N_2342,N_1792,N_1737);
nor U2343 (N_2343,N_1625,N_1829);
nor U2344 (N_2344,N_1904,N_1660);
and U2345 (N_2345,N_1767,N_1968);
or U2346 (N_2346,N_1908,N_1920);
nor U2347 (N_2347,N_1656,N_1790);
nand U2348 (N_2348,N_1672,N_1962);
nor U2349 (N_2349,N_1935,N_1611);
nor U2350 (N_2350,N_1949,N_1919);
and U2351 (N_2351,N_1607,N_1740);
nor U2352 (N_2352,N_1893,N_1991);
nor U2353 (N_2353,N_1642,N_1881);
and U2354 (N_2354,N_1702,N_1924);
nand U2355 (N_2355,N_1975,N_1829);
or U2356 (N_2356,N_1816,N_1904);
nor U2357 (N_2357,N_1913,N_1955);
nand U2358 (N_2358,N_1619,N_1983);
xor U2359 (N_2359,N_1930,N_1696);
or U2360 (N_2360,N_1747,N_1927);
or U2361 (N_2361,N_1673,N_1998);
and U2362 (N_2362,N_1703,N_1854);
nand U2363 (N_2363,N_1803,N_1921);
and U2364 (N_2364,N_1804,N_1896);
nand U2365 (N_2365,N_1682,N_1749);
and U2366 (N_2366,N_1753,N_1648);
and U2367 (N_2367,N_1880,N_1624);
or U2368 (N_2368,N_1782,N_1910);
nand U2369 (N_2369,N_1772,N_1644);
and U2370 (N_2370,N_1860,N_1845);
xnor U2371 (N_2371,N_1955,N_1753);
and U2372 (N_2372,N_1800,N_1650);
nand U2373 (N_2373,N_1767,N_1718);
nand U2374 (N_2374,N_1773,N_1678);
nand U2375 (N_2375,N_1734,N_1670);
or U2376 (N_2376,N_1814,N_1769);
nor U2377 (N_2377,N_1920,N_1907);
and U2378 (N_2378,N_1983,N_1605);
and U2379 (N_2379,N_1610,N_1870);
nand U2380 (N_2380,N_1743,N_1705);
nand U2381 (N_2381,N_1829,N_1834);
nor U2382 (N_2382,N_1955,N_1702);
or U2383 (N_2383,N_1682,N_1611);
nor U2384 (N_2384,N_1681,N_1879);
and U2385 (N_2385,N_1923,N_1975);
and U2386 (N_2386,N_1733,N_1943);
nor U2387 (N_2387,N_1781,N_1972);
and U2388 (N_2388,N_1637,N_1812);
and U2389 (N_2389,N_1767,N_1741);
nor U2390 (N_2390,N_1767,N_1755);
and U2391 (N_2391,N_1608,N_1701);
nand U2392 (N_2392,N_1961,N_1905);
or U2393 (N_2393,N_1735,N_1661);
nand U2394 (N_2394,N_1890,N_1689);
nor U2395 (N_2395,N_1940,N_1989);
nand U2396 (N_2396,N_1986,N_1910);
or U2397 (N_2397,N_1655,N_1946);
nor U2398 (N_2398,N_1625,N_1606);
nand U2399 (N_2399,N_1656,N_1719);
and U2400 (N_2400,N_2080,N_2151);
nand U2401 (N_2401,N_2380,N_2000);
nor U2402 (N_2402,N_2169,N_2199);
or U2403 (N_2403,N_2059,N_2370);
or U2404 (N_2404,N_2094,N_2387);
nor U2405 (N_2405,N_2005,N_2137);
nand U2406 (N_2406,N_2127,N_2092);
nor U2407 (N_2407,N_2099,N_2224);
nor U2408 (N_2408,N_2347,N_2369);
and U2409 (N_2409,N_2046,N_2238);
and U2410 (N_2410,N_2067,N_2084);
nor U2411 (N_2411,N_2147,N_2384);
or U2412 (N_2412,N_2001,N_2177);
or U2413 (N_2413,N_2256,N_2371);
or U2414 (N_2414,N_2276,N_2087);
nand U2415 (N_2415,N_2240,N_2219);
nor U2416 (N_2416,N_2109,N_2189);
nand U2417 (N_2417,N_2161,N_2065);
nor U2418 (N_2418,N_2341,N_2398);
nor U2419 (N_2419,N_2115,N_2023);
nor U2420 (N_2420,N_2133,N_2291);
nand U2421 (N_2421,N_2098,N_2018);
nand U2422 (N_2422,N_2322,N_2011);
or U2423 (N_2423,N_2333,N_2239);
or U2424 (N_2424,N_2212,N_2264);
nand U2425 (N_2425,N_2236,N_2351);
and U2426 (N_2426,N_2363,N_2159);
or U2427 (N_2427,N_2327,N_2213);
or U2428 (N_2428,N_2116,N_2097);
or U2429 (N_2429,N_2376,N_2183);
nand U2430 (N_2430,N_2243,N_2195);
or U2431 (N_2431,N_2292,N_2388);
and U2432 (N_2432,N_2026,N_2385);
and U2433 (N_2433,N_2392,N_2008);
nand U2434 (N_2434,N_2198,N_2299);
nor U2435 (N_2435,N_2383,N_2073);
nand U2436 (N_2436,N_2226,N_2143);
nor U2437 (N_2437,N_2132,N_2180);
or U2438 (N_2438,N_2265,N_2039);
nor U2439 (N_2439,N_2270,N_2220);
nand U2440 (N_2440,N_2128,N_2306);
and U2441 (N_2441,N_2248,N_2129);
and U2442 (N_2442,N_2389,N_2040);
and U2443 (N_2443,N_2048,N_2307);
nor U2444 (N_2444,N_2340,N_2339);
nand U2445 (N_2445,N_2288,N_2163);
and U2446 (N_2446,N_2155,N_2217);
nand U2447 (N_2447,N_2266,N_2300);
nor U2448 (N_2448,N_2148,N_2027);
nor U2449 (N_2449,N_2058,N_2022);
and U2450 (N_2450,N_2375,N_2142);
and U2451 (N_2451,N_2262,N_2395);
or U2452 (N_2452,N_2374,N_2316);
nor U2453 (N_2453,N_2358,N_2253);
or U2454 (N_2454,N_2047,N_2043);
nand U2455 (N_2455,N_2379,N_2372);
and U2456 (N_2456,N_2332,N_2378);
and U2457 (N_2457,N_2344,N_2283);
nand U2458 (N_2458,N_2172,N_2204);
or U2459 (N_2459,N_2321,N_2348);
nor U2460 (N_2460,N_2173,N_2353);
nand U2461 (N_2461,N_2086,N_2202);
or U2462 (N_2462,N_2139,N_2310);
and U2463 (N_2463,N_2287,N_2063);
nor U2464 (N_2464,N_2135,N_2206);
nand U2465 (N_2465,N_2260,N_2165);
or U2466 (N_2466,N_2211,N_2009);
nor U2467 (N_2467,N_2126,N_2136);
nor U2468 (N_2468,N_2263,N_2352);
nor U2469 (N_2469,N_2357,N_2386);
or U2470 (N_2470,N_2313,N_2038);
nor U2471 (N_2471,N_2221,N_2284);
or U2472 (N_2472,N_2308,N_2207);
nor U2473 (N_2473,N_2250,N_2382);
nor U2474 (N_2474,N_2156,N_2293);
and U2475 (N_2475,N_2187,N_2171);
nand U2476 (N_2476,N_2078,N_2294);
or U2477 (N_2477,N_2007,N_2329);
nor U2478 (N_2478,N_2095,N_2324);
nor U2479 (N_2479,N_2366,N_2072);
nand U2480 (N_2480,N_2241,N_2164);
or U2481 (N_2481,N_2326,N_2110);
nand U2482 (N_2482,N_2302,N_2205);
or U2483 (N_2483,N_2054,N_2197);
and U2484 (N_2484,N_2049,N_2235);
nor U2485 (N_2485,N_2315,N_2166);
and U2486 (N_2486,N_2330,N_2051);
nand U2487 (N_2487,N_2175,N_2361);
nor U2488 (N_2488,N_2036,N_2014);
nor U2489 (N_2489,N_2328,N_2013);
nor U2490 (N_2490,N_2319,N_2267);
xor U2491 (N_2491,N_2318,N_2334);
nand U2492 (N_2492,N_2114,N_2274);
nor U2493 (N_2493,N_2160,N_2191);
nand U2494 (N_2494,N_2037,N_2182);
or U2495 (N_2495,N_2365,N_2247);
and U2496 (N_2496,N_2056,N_2230);
nand U2497 (N_2497,N_2185,N_2196);
or U2498 (N_2498,N_2188,N_2157);
nor U2499 (N_2499,N_2050,N_2349);
nor U2500 (N_2500,N_2153,N_2068);
nor U2501 (N_2501,N_2311,N_2024);
or U2502 (N_2502,N_2216,N_2229);
and U2503 (N_2503,N_2006,N_2298);
nand U2504 (N_2504,N_2141,N_2275);
or U2505 (N_2505,N_2179,N_2085);
and U2506 (N_2506,N_2138,N_2301);
nor U2507 (N_2507,N_2228,N_2104);
nand U2508 (N_2508,N_2149,N_2119);
nor U2509 (N_2509,N_2271,N_2140);
nor U2510 (N_2510,N_2071,N_2154);
nand U2511 (N_2511,N_2079,N_2145);
or U2512 (N_2512,N_2096,N_2364);
nor U2513 (N_2513,N_2258,N_2004);
and U2514 (N_2514,N_2304,N_2045);
and U2515 (N_2515,N_2337,N_2064);
and U2516 (N_2516,N_2244,N_2338);
nand U2517 (N_2517,N_2034,N_2131);
nor U2518 (N_2518,N_2391,N_2208);
and U2519 (N_2519,N_2083,N_2261);
nand U2520 (N_2520,N_2190,N_2186);
nor U2521 (N_2521,N_2237,N_2346);
or U2522 (N_2522,N_2373,N_2150);
nand U2523 (N_2523,N_2069,N_2093);
nand U2524 (N_2524,N_2107,N_2393);
and U2525 (N_2525,N_2218,N_2025);
and U2526 (N_2526,N_2033,N_2350);
nor U2527 (N_2527,N_2354,N_2200);
nand U2528 (N_2528,N_2303,N_2254);
nand U2529 (N_2529,N_2360,N_2035);
nand U2530 (N_2530,N_2249,N_2041);
nand U2531 (N_2531,N_2231,N_2223);
or U2532 (N_2532,N_2312,N_2074);
or U2533 (N_2533,N_2090,N_2021);
and U2534 (N_2534,N_2044,N_2323);
nand U2535 (N_2535,N_2146,N_2203);
nor U2536 (N_2536,N_2162,N_2168);
nor U2537 (N_2537,N_2181,N_2210);
nor U2538 (N_2538,N_2245,N_2296);
and U2539 (N_2539,N_2314,N_2060);
nand U2540 (N_2540,N_2289,N_2381);
and U2541 (N_2541,N_2278,N_2215);
nor U2542 (N_2542,N_2081,N_2144);
or U2543 (N_2543,N_2227,N_2345);
or U2544 (N_2544,N_2120,N_2268);
nand U2545 (N_2545,N_2062,N_2320);
or U2546 (N_2546,N_2368,N_2259);
nand U2547 (N_2547,N_2367,N_2246);
nor U2548 (N_2548,N_2222,N_2076);
nor U2549 (N_2549,N_2257,N_2317);
nand U2550 (N_2550,N_2325,N_2053);
or U2551 (N_2551,N_2295,N_2108);
nor U2552 (N_2552,N_2269,N_2124);
or U2553 (N_2553,N_2342,N_2010);
nand U2554 (N_2554,N_2030,N_2070);
and U2555 (N_2555,N_2234,N_2003);
nor U2556 (N_2556,N_2105,N_2075);
or U2557 (N_2557,N_2335,N_2390);
nand U2558 (N_2558,N_2016,N_2103);
or U2559 (N_2559,N_2396,N_2088);
or U2560 (N_2560,N_2193,N_2020);
nor U2561 (N_2561,N_2077,N_2282);
nand U2562 (N_2562,N_2209,N_2019);
nand U2563 (N_2563,N_2130,N_2012);
nor U2564 (N_2564,N_2112,N_2290);
nand U2565 (N_2565,N_2089,N_2362);
nor U2566 (N_2566,N_2279,N_2280);
or U2567 (N_2567,N_2117,N_2285);
and U2568 (N_2568,N_2356,N_2297);
nand U2569 (N_2569,N_2232,N_2082);
nor U2570 (N_2570,N_2201,N_2331);
and U2571 (N_2571,N_2174,N_2152);
nand U2572 (N_2572,N_2042,N_2399);
nor U2573 (N_2573,N_2100,N_2343);
and U2574 (N_2574,N_2336,N_2118);
nand U2575 (N_2575,N_2017,N_2184);
nor U2576 (N_2576,N_2309,N_2394);
nand U2577 (N_2577,N_2091,N_2111);
xnor U2578 (N_2578,N_2106,N_2134);
nand U2579 (N_2579,N_2121,N_2158);
and U2580 (N_2580,N_2233,N_2273);
nand U2581 (N_2581,N_2015,N_2170);
and U2582 (N_2582,N_2255,N_2272);
nor U2583 (N_2583,N_2028,N_2122);
nand U2584 (N_2584,N_2225,N_2355);
nor U2585 (N_2585,N_2101,N_2192);
or U2586 (N_2586,N_2252,N_2242);
nor U2587 (N_2587,N_2066,N_2305);
nor U2588 (N_2588,N_2251,N_2032);
and U2589 (N_2589,N_2281,N_2123);
nor U2590 (N_2590,N_2194,N_2286);
nand U2591 (N_2591,N_2377,N_2277);
and U2592 (N_2592,N_2057,N_2125);
and U2593 (N_2593,N_2031,N_2214);
nand U2594 (N_2594,N_2397,N_2055);
or U2595 (N_2595,N_2061,N_2052);
or U2596 (N_2596,N_2178,N_2102);
nor U2597 (N_2597,N_2176,N_2113);
nor U2598 (N_2598,N_2002,N_2359);
or U2599 (N_2599,N_2167,N_2029);
and U2600 (N_2600,N_2141,N_2372);
or U2601 (N_2601,N_2207,N_2188);
nor U2602 (N_2602,N_2105,N_2092);
or U2603 (N_2603,N_2195,N_2001);
nand U2604 (N_2604,N_2024,N_2219);
and U2605 (N_2605,N_2172,N_2016);
nor U2606 (N_2606,N_2038,N_2047);
nor U2607 (N_2607,N_2351,N_2244);
nand U2608 (N_2608,N_2336,N_2039);
nand U2609 (N_2609,N_2109,N_2001);
nor U2610 (N_2610,N_2304,N_2120);
nor U2611 (N_2611,N_2379,N_2213);
nor U2612 (N_2612,N_2171,N_2337);
nand U2613 (N_2613,N_2212,N_2227);
xnor U2614 (N_2614,N_2056,N_2186);
or U2615 (N_2615,N_2018,N_2000);
nor U2616 (N_2616,N_2119,N_2305);
or U2617 (N_2617,N_2025,N_2038);
nand U2618 (N_2618,N_2266,N_2261);
nand U2619 (N_2619,N_2352,N_2010);
or U2620 (N_2620,N_2188,N_2350);
nor U2621 (N_2621,N_2172,N_2090);
nand U2622 (N_2622,N_2347,N_2291);
nand U2623 (N_2623,N_2262,N_2274);
and U2624 (N_2624,N_2119,N_2045);
nand U2625 (N_2625,N_2163,N_2386);
or U2626 (N_2626,N_2041,N_2363);
nand U2627 (N_2627,N_2130,N_2056);
and U2628 (N_2628,N_2285,N_2058);
nand U2629 (N_2629,N_2379,N_2343);
nand U2630 (N_2630,N_2242,N_2090);
nand U2631 (N_2631,N_2221,N_2279);
and U2632 (N_2632,N_2091,N_2213);
nor U2633 (N_2633,N_2274,N_2220);
or U2634 (N_2634,N_2367,N_2383);
or U2635 (N_2635,N_2021,N_2255);
or U2636 (N_2636,N_2176,N_2321);
and U2637 (N_2637,N_2110,N_2090);
nand U2638 (N_2638,N_2353,N_2070);
nor U2639 (N_2639,N_2146,N_2333);
or U2640 (N_2640,N_2125,N_2344);
and U2641 (N_2641,N_2212,N_2107);
or U2642 (N_2642,N_2205,N_2361);
nand U2643 (N_2643,N_2018,N_2066);
or U2644 (N_2644,N_2046,N_2240);
and U2645 (N_2645,N_2161,N_2114);
or U2646 (N_2646,N_2021,N_2168);
and U2647 (N_2647,N_2136,N_2162);
or U2648 (N_2648,N_2129,N_2326);
or U2649 (N_2649,N_2249,N_2225);
nand U2650 (N_2650,N_2268,N_2344);
nand U2651 (N_2651,N_2349,N_2230);
nand U2652 (N_2652,N_2237,N_2064);
and U2653 (N_2653,N_2289,N_2305);
or U2654 (N_2654,N_2194,N_2115);
or U2655 (N_2655,N_2266,N_2039);
and U2656 (N_2656,N_2339,N_2220);
or U2657 (N_2657,N_2322,N_2066);
or U2658 (N_2658,N_2338,N_2195);
nand U2659 (N_2659,N_2195,N_2222);
nand U2660 (N_2660,N_2199,N_2015);
and U2661 (N_2661,N_2370,N_2023);
and U2662 (N_2662,N_2105,N_2028);
or U2663 (N_2663,N_2013,N_2383);
or U2664 (N_2664,N_2313,N_2040);
nor U2665 (N_2665,N_2399,N_2292);
nor U2666 (N_2666,N_2253,N_2313);
nor U2667 (N_2667,N_2131,N_2180);
nor U2668 (N_2668,N_2044,N_2314);
and U2669 (N_2669,N_2358,N_2332);
nand U2670 (N_2670,N_2395,N_2245);
nand U2671 (N_2671,N_2288,N_2099);
nand U2672 (N_2672,N_2287,N_2097);
and U2673 (N_2673,N_2034,N_2146);
nor U2674 (N_2674,N_2238,N_2387);
or U2675 (N_2675,N_2140,N_2244);
nor U2676 (N_2676,N_2198,N_2056);
nor U2677 (N_2677,N_2160,N_2309);
nand U2678 (N_2678,N_2217,N_2271);
or U2679 (N_2679,N_2211,N_2081);
nand U2680 (N_2680,N_2353,N_2106);
nor U2681 (N_2681,N_2206,N_2297);
or U2682 (N_2682,N_2331,N_2375);
or U2683 (N_2683,N_2153,N_2316);
and U2684 (N_2684,N_2310,N_2365);
or U2685 (N_2685,N_2281,N_2259);
nor U2686 (N_2686,N_2110,N_2015);
or U2687 (N_2687,N_2240,N_2235);
nor U2688 (N_2688,N_2035,N_2130);
nor U2689 (N_2689,N_2199,N_2369);
or U2690 (N_2690,N_2029,N_2082);
xor U2691 (N_2691,N_2120,N_2375);
and U2692 (N_2692,N_2349,N_2326);
nand U2693 (N_2693,N_2229,N_2056);
nor U2694 (N_2694,N_2346,N_2354);
nor U2695 (N_2695,N_2167,N_2186);
nor U2696 (N_2696,N_2030,N_2379);
nand U2697 (N_2697,N_2322,N_2036);
nand U2698 (N_2698,N_2047,N_2104);
or U2699 (N_2699,N_2095,N_2398);
nor U2700 (N_2700,N_2278,N_2287);
and U2701 (N_2701,N_2002,N_2385);
or U2702 (N_2702,N_2289,N_2042);
nand U2703 (N_2703,N_2324,N_2070);
and U2704 (N_2704,N_2009,N_2218);
nand U2705 (N_2705,N_2268,N_2331);
nand U2706 (N_2706,N_2110,N_2344);
nor U2707 (N_2707,N_2286,N_2251);
nand U2708 (N_2708,N_2280,N_2078);
and U2709 (N_2709,N_2236,N_2026);
and U2710 (N_2710,N_2061,N_2323);
nor U2711 (N_2711,N_2186,N_2396);
nand U2712 (N_2712,N_2394,N_2174);
nor U2713 (N_2713,N_2179,N_2217);
xnor U2714 (N_2714,N_2123,N_2370);
nor U2715 (N_2715,N_2285,N_2182);
nand U2716 (N_2716,N_2108,N_2068);
nor U2717 (N_2717,N_2061,N_2260);
and U2718 (N_2718,N_2102,N_2078);
nand U2719 (N_2719,N_2154,N_2159);
nand U2720 (N_2720,N_2392,N_2308);
and U2721 (N_2721,N_2123,N_2171);
or U2722 (N_2722,N_2157,N_2129);
nor U2723 (N_2723,N_2035,N_2075);
nor U2724 (N_2724,N_2216,N_2157);
and U2725 (N_2725,N_2228,N_2185);
nand U2726 (N_2726,N_2052,N_2153);
or U2727 (N_2727,N_2211,N_2267);
and U2728 (N_2728,N_2031,N_2392);
nor U2729 (N_2729,N_2113,N_2239);
and U2730 (N_2730,N_2107,N_2229);
and U2731 (N_2731,N_2036,N_2176);
nor U2732 (N_2732,N_2354,N_2380);
and U2733 (N_2733,N_2314,N_2280);
nand U2734 (N_2734,N_2333,N_2204);
nand U2735 (N_2735,N_2052,N_2225);
nor U2736 (N_2736,N_2047,N_2176);
and U2737 (N_2737,N_2168,N_2311);
or U2738 (N_2738,N_2278,N_2175);
and U2739 (N_2739,N_2224,N_2208);
or U2740 (N_2740,N_2106,N_2129);
and U2741 (N_2741,N_2354,N_2154);
and U2742 (N_2742,N_2172,N_2276);
and U2743 (N_2743,N_2154,N_2138);
and U2744 (N_2744,N_2076,N_2256);
or U2745 (N_2745,N_2309,N_2379);
nand U2746 (N_2746,N_2316,N_2019);
or U2747 (N_2747,N_2311,N_2301);
or U2748 (N_2748,N_2118,N_2134);
nand U2749 (N_2749,N_2157,N_2352);
or U2750 (N_2750,N_2014,N_2271);
and U2751 (N_2751,N_2191,N_2309);
nor U2752 (N_2752,N_2041,N_2129);
or U2753 (N_2753,N_2113,N_2283);
and U2754 (N_2754,N_2141,N_2069);
or U2755 (N_2755,N_2067,N_2344);
and U2756 (N_2756,N_2013,N_2361);
nor U2757 (N_2757,N_2009,N_2294);
nand U2758 (N_2758,N_2039,N_2054);
or U2759 (N_2759,N_2329,N_2260);
or U2760 (N_2760,N_2224,N_2329);
or U2761 (N_2761,N_2214,N_2234);
nand U2762 (N_2762,N_2231,N_2371);
and U2763 (N_2763,N_2025,N_2307);
nor U2764 (N_2764,N_2252,N_2026);
nand U2765 (N_2765,N_2094,N_2239);
nor U2766 (N_2766,N_2187,N_2344);
nand U2767 (N_2767,N_2016,N_2344);
or U2768 (N_2768,N_2291,N_2013);
nand U2769 (N_2769,N_2398,N_2312);
nor U2770 (N_2770,N_2366,N_2028);
or U2771 (N_2771,N_2177,N_2355);
nand U2772 (N_2772,N_2282,N_2352);
or U2773 (N_2773,N_2328,N_2151);
and U2774 (N_2774,N_2359,N_2237);
or U2775 (N_2775,N_2271,N_2155);
or U2776 (N_2776,N_2225,N_2394);
nand U2777 (N_2777,N_2298,N_2002);
and U2778 (N_2778,N_2395,N_2277);
and U2779 (N_2779,N_2186,N_2000);
nand U2780 (N_2780,N_2348,N_2172);
or U2781 (N_2781,N_2049,N_2353);
nand U2782 (N_2782,N_2389,N_2037);
nand U2783 (N_2783,N_2205,N_2068);
nor U2784 (N_2784,N_2183,N_2325);
and U2785 (N_2785,N_2366,N_2011);
or U2786 (N_2786,N_2082,N_2256);
or U2787 (N_2787,N_2035,N_2118);
nand U2788 (N_2788,N_2081,N_2056);
or U2789 (N_2789,N_2027,N_2080);
nand U2790 (N_2790,N_2204,N_2056);
nand U2791 (N_2791,N_2279,N_2259);
and U2792 (N_2792,N_2334,N_2103);
nand U2793 (N_2793,N_2198,N_2385);
or U2794 (N_2794,N_2044,N_2220);
or U2795 (N_2795,N_2221,N_2052);
and U2796 (N_2796,N_2115,N_2330);
and U2797 (N_2797,N_2163,N_2303);
or U2798 (N_2798,N_2212,N_2113);
nor U2799 (N_2799,N_2330,N_2015);
and U2800 (N_2800,N_2766,N_2608);
and U2801 (N_2801,N_2564,N_2617);
nand U2802 (N_2802,N_2727,N_2695);
or U2803 (N_2803,N_2526,N_2578);
and U2804 (N_2804,N_2508,N_2665);
nor U2805 (N_2805,N_2791,N_2437);
and U2806 (N_2806,N_2536,N_2410);
nand U2807 (N_2807,N_2653,N_2655);
nand U2808 (N_2808,N_2794,N_2552);
nor U2809 (N_2809,N_2505,N_2786);
and U2810 (N_2810,N_2560,N_2623);
and U2811 (N_2811,N_2614,N_2668);
or U2812 (N_2812,N_2405,N_2787);
and U2813 (N_2813,N_2458,N_2618);
or U2814 (N_2814,N_2416,N_2544);
or U2815 (N_2815,N_2688,N_2677);
and U2816 (N_2816,N_2561,N_2533);
or U2817 (N_2817,N_2629,N_2640);
or U2818 (N_2818,N_2720,N_2517);
and U2819 (N_2819,N_2563,N_2630);
nand U2820 (N_2820,N_2598,N_2469);
nor U2821 (N_2821,N_2482,N_2797);
and U2822 (N_2822,N_2656,N_2420);
and U2823 (N_2823,N_2584,N_2474);
nand U2824 (N_2824,N_2429,N_2478);
nor U2825 (N_2825,N_2499,N_2481);
and U2826 (N_2826,N_2570,N_2657);
nand U2827 (N_2827,N_2470,N_2734);
nor U2828 (N_2828,N_2631,N_2738);
nand U2829 (N_2829,N_2464,N_2792);
and U2830 (N_2830,N_2520,N_2445);
nand U2831 (N_2831,N_2739,N_2435);
nand U2832 (N_2832,N_2409,N_2406);
nor U2833 (N_2833,N_2597,N_2696);
nand U2834 (N_2834,N_2527,N_2613);
nand U2835 (N_2835,N_2576,N_2730);
nand U2836 (N_2836,N_2615,N_2676);
and U2837 (N_2837,N_2585,N_2486);
and U2838 (N_2838,N_2459,N_2779);
and U2839 (N_2839,N_2782,N_2634);
or U2840 (N_2840,N_2760,N_2412);
or U2841 (N_2841,N_2740,N_2522);
nand U2842 (N_2842,N_2682,N_2546);
and U2843 (N_2843,N_2600,N_2780);
and U2844 (N_2844,N_2492,N_2541);
or U2845 (N_2845,N_2708,N_2693);
and U2846 (N_2846,N_2619,N_2683);
xor U2847 (N_2847,N_2756,N_2471);
and U2848 (N_2848,N_2750,N_2414);
or U2849 (N_2849,N_2594,N_2463);
nand U2850 (N_2850,N_2551,N_2441);
nand U2851 (N_2851,N_2559,N_2711);
or U2852 (N_2852,N_2593,N_2699);
or U2853 (N_2853,N_2515,N_2547);
nor U2854 (N_2854,N_2601,N_2789);
nor U2855 (N_2855,N_2581,N_2663);
nand U2856 (N_2856,N_2778,N_2558);
nand U2857 (N_2857,N_2607,N_2509);
nor U2858 (N_2858,N_2524,N_2698);
or U2859 (N_2859,N_2588,N_2436);
and U2860 (N_2860,N_2624,N_2736);
nor U2861 (N_2861,N_2769,N_2692);
nor U2862 (N_2862,N_2670,N_2709);
nor U2863 (N_2863,N_2504,N_2431);
and U2864 (N_2864,N_2511,N_2702);
and U2865 (N_2865,N_2606,N_2773);
nand U2866 (N_2866,N_2719,N_2785);
and U2867 (N_2867,N_2743,N_2567);
and U2868 (N_2868,N_2427,N_2408);
nor U2869 (N_2869,N_2674,N_2771);
or U2870 (N_2870,N_2438,N_2661);
or U2871 (N_2871,N_2724,N_2513);
nand U2872 (N_2872,N_2506,N_2767);
nand U2873 (N_2873,N_2444,N_2523);
and U2874 (N_2874,N_2641,N_2535);
or U2875 (N_2875,N_2496,N_2799);
or U2876 (N_2876,N_2554,N_2667);
and U2877 (N_2877,N_2647,N_2681);
and U2878 (N_2878,N_2443,N_2484);
nor U2879 (N_2879,N_2611,N_2426);
nand U2880 (N_2880,N_2686,N_2777);
and U2881 (N_2881,N_2604,N_2716);
and U2882 (N_2882,N_2784,N_2555);
or U2883 (N_2883,N_2735,N_2537);
and U2884 (N_2884,N_2400,N_2449);
nor U2885 (N_2885,N_2538,N_2639);
nor U2886 (N_2886,N_2652,N_2574);
nand U2887 (N_2887,N_2746,N_2485);
and U2888 (N_2888,N_2495,N_2691);
or U2889 (N_2889,N_2788,N_2534);
nand U2890 (N_2890,N_2498,N_2425);
nand U2891 (N_2891,N_2660,N_2421);
or U2892 (N_2892,N_2710,N_2599);
or U2893 (N_2893,N_2731,N_2540);
nor U2894 (N_2894,N_2487,N_2562);
and U2895 (N_2895,N_2568,N_2589);
and U2896 (N_2896,N_2772,N_2763);
nor U2897 (N_2897,N_2516,N_2451);
or U2898 (N_2898,N_2573,N_2664);
or U2899 (N_2899,N_2415,N_2501);
nor U2900 (N_2900,N_2654,N_2493);
nand U2901 (N_2901,N_2530,N_2455);
or U2902 (N_2902,N_2553,N_2565);
nand U2903 (N_2903,N_2472,N_2685);
and U2904 (N_2904,N_2662,N_2675);
or U2905 (N_2905,N_2642,N_2602);
nand U2906 (N_2906,N_2793,N_2433);
nor U2907 (N_2907,N_2669,N_2625);
nor U2908 (N_2908,N_2612,N_2759);
nor U2909 (N_2909,N_2467,N_2539);
and U2910 (N_2910,N_2483,N_2590);
and U2911 (N_2911,N_2402,N_2440);
and U2912 (N_2912,N_2783,N_2439);
nor U2913 (N_2913,N_2737,N_2518);
or U2914 (N_2914,N_2419,N_2684);
or U2915 (N_2915,N_2697,N_2770);
and U2916 (N_2916,N_2632,N_2694);
nor U2917 (N_2917,N_2423,N_2745);
and U2918 (N_2918,N_2721,N_2512);
or U2919 (N_2919,N_2411,N_2479);
nor U2920 (N_2920,N_2666,N_2480);
and U2921 (N_2921,N_2579,N_2753);
and U2922 (N_2922,N_2757,N_2502);
or U2923 (N_2923,N_2749,N_2418);
and U2924 (N_2924,N_2548,N_2477);
nand U2925 (N_2925,N_2754,N_2417);
nor U2926 (N_2926,N_2457,N_2532);
nand U2927 (N_2927,N_2627,N_2475);
or U2928 (N_2928,N_2500,N_2672);
and U2929 (N_2929,N_2728,N_2690);
or U2930 (N_2930,N_2447,N_2596);
and U2931 (N_2931,N_2460,N_2529);
and U2932 (N_2932,N_2545,N_2580);
or U2933 (N_2933,N_2622,N_2528);
nand U2934 (N_2934,N_2796,N_2747);
nand U2935 (N_2935,N_2706,N_2489);
or U2936 (N_2936,N_2507,N_2742);
or U2937 (N_2937,N_2543,N_2491);
or U2938 (N_2938,N_2542,N_2610);
or U2939 (N_2939,N_2725,N_2679);
and U2940 (N_2940,N_2466,N_2572);
and U2941 (N_2941,N_2790,N_2550);
and U2942 (N_2942,N_2595,N_2497);
and U2943 (N_2943,N_2718,N_2432);
nand U2944 (N_2944,N_2603,N_2752);
or U2945 (N_2945,N_2671,N_2403);
or U2946 (N_2946,N_2673,N_2450);
nor U2947 (N_2947,N_2658,N_2704);
nand U2948 (N_2948,N_2636,N_2775);
or U2949 (N_2949,N_2776,N_2571);
nor U2950 (N_2950,N_2446,N_2557);
nor U2951 (N_2951,N_2626,N_2490);
or U2952 (N_2952,N_2714,N_2424);
and U2953 (N_2953,N_2659,N_2442);
and U2954 (N_2954,N_2521,N_2687);
nor U2955 (N_2955,N_2705,N_2582);
and U2956 (N_2956,N_2448,N_2758);
or U2957 (N_2957,N_2413,N_2609);
and U2958 (N_2958,N_2605,N_2592);
or U2959 (N_2959,N_2488,N_2726);
nand U2960 (N_2960,N_2722,N_2741);
nor U2961 (N_2961,N_2628,N_2729);
nor U2962 (N_2962,N_2473,N_2700);
nand U2963 (N_2963,N_2650,N_2569);
or U2964 (N_2964,N_2765,N_2407);
nand U2965 (N_2965,N_2525,N_2638);
nor U2966 (N_2966,N_2712,N_2633);
and U2967 (N_2967,N_2514,N_2703);
and U2968 (N_2968,N_2452,N_2510);
nor U2969 (N_2969,N_2651,N_2401);
nor U2970 (N_2970,N_2733,N_2428);
nor U2971 (N_2971,N_2468,N_2707);
or U2972 (N_2972,N_2465,N_2713);
and U2973 (N_2973,N_2494,N_2646);
nor U2974 (N_2974,N_2404,N_2748);
or U2975 (N_2975,N_2701,N_2774);
and U2976 (N_2976,N_2643,N_2453);
nand U2977 (N_2977,N_2556,N_2649);
nor U2978 (N_2978,N_2717,N_2461);
or U2979 (N_2979,N_2587,N_2744);
or U2980 (N_2980,N_2577,N_2616);
nand U2981 (N_2981,N_2755,N_2621);
and U2982 (N_2982,N_2689,N_2456);
and U2983 (N_2983,N_2768,N_2519);
nor U2984 (N_2984,N_2454,N_2644);
and U2985 (N_2985,N_2566,N_2434);
or U2986 (N_2986,N_2620,N_2635);
or U2987 (N_2987,N_2761,N_2781);
nor U2988 (N_2988,N_2680,N_2583);
nand U2989 (N_2989,N_2795,N_2764);
and U2990 (N_2990,N_2637,N_2430);
or U2991 (N_2991,N_2645,N_2751);
or U2992 (N_2992,N_2422,N_2678);
and U2993 (N_2993,N_2531,N_2648);
or U2994 (N_2994,N_2732,N_2549);
and U2995 (N_2995,N_2715,N_2462);
or U2996 (N_2996,N_2723,N_2503);
nor U2997 (N_2997,N_2591,N_2762);
or U2998 (N_2998,N_2575,N_2476);
nand U2999 (N_2999,N_2586,N_2798);
and U3000 (N_3000,N_2728,N_2507);
nand U3001 (N_3001,N_2430,N_2652);
and U3002 (N_3002,N_2416,N_2600);
and U3003 (N_3003,N_2798,N_2670);
nand U3004 (N_3004,N_2751,N_2733);
and U3005 (N_3005,N_2793,N_2483);
and U3006 (N_3006,N_2545,N_2755);
nor U3007 (N_3007,N_2624,N_2555);
or U3008 (N_3008,N_2403,N_2478);
and U3009 (N_3009,N_2571,N_2744);
nor U3010 (N_3010,N_2775,N_2510);
or U3011 (N_3011,N_2767,N_2733);
nand U3012 (N_3012,N_2717,N_2723);
nand U3013 (N_3013,N_2495,N_2731);
or U3014 (N_3014,N_2620,N_2603);
or U3015 (N_3015,N_2539,N_2737);
nand U3016 (N_3016,N_2631,N_2441);
nand U3017 (N_3017,N_2400,N_2560);
nor U3018 (N_3018,N_2545,N_2515);
nand U3019 (N_3019,N_2404,N_2782);
nor U3020 (N_3020,N_2404,N_2420);
nand U3021 (N_3021,N_2685,N_2456);
or U3022 (N_3022,N_2585,N_2607);
nor U3023 (N_3023,N_2688,N_2710);
or U3024 (N_3024,N_2561,N_2492);
nand U3025 (N_3025,N_2638,N_2452);
nor U3026 (N_3026,N_2759,N_2777);
nor U3027 (N_3027,N_2796,N_2604);
or U3028 (N_3028,N_2638,N_2485);
nand U3029 (N_3029,N_2796,N_2618);
nor U3030 (N_3030,N_2597,N_2611);
or U3031 (N_3031,N_2483,N_2653);
nor U3032 (N_3032,N_2686,N_2428);
nand U3033 (N_3033,N_2626,N_2766);
nand U3034 (N_3034,N_2584,N_2670);
and U3035 (N_3035,N_2707,N_2579);
and U3036 (N_3036,N_2581,N_2538);
nor U3037 (N_3037,N_2670,N_2528);
nor U3038 (N_3038,N_2437,N_2688);
or U3039 (N_3039,N_2609,N_2650);
nor U3040 (N_3040,N_2563,N_2421);
nor U3041 (N_3041,N_2605,N_2658);
nand U3042 (N_3042,N_2615,N_2445);
nor U3043 (N_3043,N_2424,N_2584);
and U3044 (N_3044,N_2641,N_2517);
and U3045 (N_3045,N_2417,N_2404);
or U3046 (N_3046,N_2752,N_2690);
nand U3047 (N_3047,N_2689,N_2460);
or U3048 (N_3048,N_2763,N_2792);
and U3049 (N_3049,N_2657,N_2620);
nor U3050 (N_3050,N_2563,N_2530);
nor U3051 (N_3051,N_2645,N_2636);
or U3052 (N_3052,N_2746,N_2635);
or U3053 (N_3053,N_2431,N_2753);
nand U3054 (N_3054,N_2566,N_2791);
and U3055 (N_3055,N_2716,N_2794);
nand U3056 (N_3056,N_2440,N_2518);
and U3057 (N_3057,N_2648,N_2619);
and U3058 (N_3058,N_2425,N_2468);
nor U3059 (N_3059,N_2601,N_2695);
or U3060 (N_3060,N_2617,N_2550);
nand U3061 (N_3061,N_2709,N_2405);
or U3062 (N_3062,N_2653,N_2654);
or U3063 (N_3063,N_2437,N_2641);
nand U3064 (N_3064,N_2521,N_2496);
nand U3065 (N_3065,N_2700,N_2563);
nand U3066 (N_3066,N_2400,N_2761);
nand U3067 (N_3067,N_2445,N_2585);
nor U3068 (N_3068,N_2440,N_2425);
nand U3069 (N_3069,N_2577,N_2540);
and U3070 (N_3070,N_2418,N_2628);
or U3071 (N_3071,N_2646,N_2527);
or U3072 (N_3072,N_2473,N_2589);
and U3073 (N_3073,N_2480,N_2585);
nor U3074 (N_3074,N_2414,N_2428);
or U3075 (N_3075,N_2421,N_2625);
nor U3076 (N_3076,N_2475,N_2401);
or U3077 (N_3077,N_2667,N_2483);
nor U3078 (N_3078,N_2698,N_2563);
and U3079 (N_3079,N_2619,N_2483);
and U3080 (N_3080,N_2525,N_2668);
or U3081 (N_3081,N_2724,N_2512);
or U3082 (N_3082,N_2699,N_2740);
or U3083 (N_3083,N_2623,N_2485);
nand U3084 (N_3084,N_2767,N_2627);
nand U3085 (N_3085,N_2788,N_2618);
xnor U3086 (N_3086,N_2470,N_2703);
nor U3087 (N_3087,N_2661,N_2441);
or U3088 (N_3088,N_2693,N_2703);
nor U3089 (N_3089,N_2529,N_2590);
or U3090 (N_3090,N_2719,N_2451);
or U3091 (N_3091,N_2520,N_2628);
nor U3092 (N_3092,N_2460,N_2411);
or U3093 (N_3093,N_2543,N_2415);
or U3094 (N_3094,N_2680,N_2460);
or U3095 (N_3095,N_2542,N_2593);
or U3096 (N_3096,N_2689,N_2550);
nand U3097 (N_3097,N_2707,N_2767);
nor U3098 (N_3098,N_2674,N_2689);
and U3099 (N_3099,N_2486,N_2452);
nor U3100 (N_3100,N_2428,N_2528);
nand U3101 (N_3101,N_2635,N_2582);
nor U3102 (N_3102,N_2693,N_2614);
nand U3103 (N_3103,N_2635,N_2641);
nand U3104 (N_3104,N_2580,N_2583);
or U3105 (N_3105,N_2629,N_2416);
or U3106 (N_3106,N_2481,N_2596);
nor U3107 (N_3107,N_2508,N_2788);
nand U3108 (N_3108,N_2528,N_2643);
or U3109 (N_3109,N_2411,N_2428);
or U3110 (N_3110,N_2751,N_2449);
or U3111 (N_3111,N_2571,N_2648);
nor U3112 (N_3112,N_2660,N_2718);
nor U3113 (N_3113,N_2668,N_2473);
nand U3114 (N_3114,N_2579,N_2709);
and U3115 (N_3115,N_2610,N_2586);
nand U3116 (N_3116,N_2593,N_2411);
or U3117 (N_3117,N_2796,N_2721);
and U3118 (N_3118,N_2475,N_2792);
nor U3119 (N_3119,N_2686,N_2662);
and U3120 (N_3120,N_2748,N_2470);
or U3121 (N_3121,N_2413,N_2605);
nor U3122 (N_3122,N_2574,N_2579);
and U3123 (N_3123,N_2766,N_2759);
and U3124 (N_3124,N_2799,N_2577);
nor U3125 (N_3125,N_2407,N_2452);
and U3126 (N_3126,N_2640,N_2705);
or U3127 (N_3127,N_2432,N_2419);
nand U3128 (N_3128,N_2608,N_2407);
nor U3129 (N_3129,N_2726,N_2567);
nand U3130 (N_3130,N_2522,N_2694);
nand U3131 (N_3131,N_2690,N_2495);
and U3132 (N_3132,N_2551,N_2764);
or U3133 (N_3133,N_2435,N_2742);
and U3134 (N_3134,N_2637,N_2458);
nand U3135 (N_3135,N_2422,N_2459);
and U3136 (N_3136,N_2611,N_2589);
xor U3137 (N_3137,N_2471,N_2502);
and U3138 (N_3138,N_2601,N_2437);
nor U3139 (N_3139,N_2659,N_2524);
nand U3140 (N_3140,N_2765,N_2505);
nand U3141 (N_3141,N_2619,N_2612);
or U3142 (N_3142,N_2621,N_2557);
nor U3143 (N_3143,N_2781,N_2787);
nor U3144 (N_3144,N_2537,N_2645);
nor U3145 (N_3145,N_2524,N_2759);
and U3146 (N_3146,N_2560,N_2632);
nor U3147 (N_3147,N_2718,N_2521);
nor U3148 (N_3148,N_2656,N_2615);
and U3149 (N_3149,N_2502,N_2408);
nand U3150 (N_3150,N_2530,N_2773);
and U3151 (N_3151,N_2463,N_2743);
nor U3152 (N_3152,N_2627,N_2755);
or U3153 (N_3153,N_2644,N_2767);
nor U3154 (N_3154,N_2521,N_2533);
nand U3155 (N_3155,N_2732,N_2763);
and U3156 (N_3156,N_2772,N_2551);
and U3157 (N_3157,N_2414,N_2713);
nor U3158 (N_3158,N_2603,N_2709);
nor U3159 (N_3159,N_2489,N_2525);
and U3160 (N_3160,N_2513,N_2612);
nor U3161 (N_3161,N_2704,N_2569);
and U3162 (N_3162,N_2584,N_2540);
or U3163 (N_3163,N_2665,N_2767);
xnor U3164 (N_3164,N_2796,N_2749);
nor U3165 (N_3165,N_2536,N_2488);
nor U3166 (N_3166,N_2404,N_2573);
and U3167 (N_3167,N_2590,N_2712);
or U3168 (N_3168,N_2459,N_2606);
nand U3169 (N_3169,N_2444,N_2549);
nand U3170 (N_3170,N_2772,N_2440);
or U3171 (N_3171,N_2505,N_2669);
nand U3172 (N_3172,N_2636,N_2402);
and U3173 (N_3173,N_2508,N_2633);
nand U3174 (N_3174,N_2480,N_2492);
and U3175 (N_3175,N_2476,N_2470);
and U3176 (N_3176,N_2563,N_2708);
nand U3177 (N_3177,N_2570,N_2585);
or U3178 (N_3178,N_2421,N_2476);
nor U3179 (N_3179,N_2556,N_2479);
and U3180 (N_3180,N_2735,N_2669);
nor U3181 (N_3181,N_2589,N_2449);
nor U3182 (N_3182,N_2592,N_2569);
or U3183 (N_3183,N_2668,N_2791);
or U3184 (N_3184,N_2446,N_2434);
nor U3185 (N_3185,N_2716,N_2590);
nor U3186 (N_3186,N_2735,N_2538);
nand U3187 (N_3187,N_2444,N_2659);
nand U3188 (N_3188,N_2575,N_2668);
xor U3189 (N_3189,N_2517,N_2747);
or U3190 (N_3190,N_2417,N_2539);
nor U3191 (N_3191,N_2755,N_2453);
nor U3192 (N_3192,N_2458,N_2692);
and U3193 (N_3193,N_2751,N_2714);
nor U3194 (N_3194,N_2403,N_2791);
nand U3195 (N_3195,N_2559,N_2741);
and U3196 (N_3196,N_2525,N_2660);
or U3197 (N_3197,N_2634,N_2477);
and U3198 (N_3198,N_2785,N_2686);
and U3199 (N_3199,N_2518,N_2774);
and U3200 (N_3200,N_2922,N_3024);
and U3201 (N_3201,N_3167,N_2959);
nor U3202 (N_3202,N_2891,N_2921);
or U3203 (N_3203,N_3067,N_2841);
nor U3204 (N_3204,N_2852,N_2906);
and U3205 (N_3205,N_2816,N_2909);
nand U3206 (N_3206,N_3076,N_3165);
nor U3207 (N_3207,N_2999,N_2970);
and U3208 (N_3208,N_2968,N_2819);
nand U3209 (N_3209,N_3149,N_2877);
nand U3210 (N_3210,N_2808,N_2810);
nor U3211 (N_3211,N_2856,N_3048);
or U3212 (N_3212,N_2935,N_3077);
and U3213 (N_3213,N_2971,N_2826);
nor U3214 (N_3214,N_3125,N_3042);
or U3215 (N_3215,N_2870,N_3029);
or U3216 (N_3216,N_3016,N_2963);
and U3217 (N_3217,N_3050,N_3082);
and U3218 (N_3218,N_3145,N_3113);
and U3219 (N_3219,N_2830,N_2927);
or U3220 (N_3220,N_2855,N_2872);
nor U3221 (N_3221,N_2868,N_2801);
nand U3222 (N_3222,N_3041,N_2951);
and U3223 (N_3223,N_3054,N_2843);
or U3224 (N_3224,N_3101,N_3004);
nand U3225 (N_3225,N_3047,N_2882);
and U3226 (N_3226,N_3034,N_2937);
and U3227 (N_3227,N_2897,N_3063);
nand U3228 (N_3228,N_2978,N_2859);
nand U3229 (N_3229,N_3116,N_2874);
and U3230 (N_3230,N_2892,N_3065);
nand U3231 (N_3231,N_3068,N_3155);
or U3232 (N_3232,N_3123,N_2955);
nor U3233 (N_3233,N_2887,N_2854);
or U3234 (N_3234,N_2840,N_2957);
and U3235 (N_3235,N_2910,N_3127);
nor U3236 (N_3236,N_3179,N_2814);
and U3237 (N_3237,N_3028,N_3006);
or U3238 (N_3238,N_3018,N_3130);
or U3239 (N_3239,N_2938,N_3049);
nand U3240 (N_3240,N_2934,N_2829);
nor U3241 (N_3241,N_2903,N_2871);
or U3242 (N_3242,N_2848,N_3141);
or U3243 (N_3243,N_2881,N_2912);
and U3244 (N_3244,N_3073,N_2976);
nand U3245 (N_3245,N_2905,N_2834);
and U3246 (N_3246,N_3121,N_2981);
or U3247 (N_3247,N_2867,N_3007);
or U3248 (N_3248,N_3015,N_2896);
nand U3249 (N_3249,N_3084,N_3043);
nand U3250 (N_3250,N_3191,N_3119);
nand U3251 (N_3251,N_3071,N_2929);
nand U3252 (N_3252,N_2811,N_3147);
nand U3253 (N_3253,N_3037,N_3008);
nor U3254 (N_3254,N_3107,N_2885);
nand U3255 (N_3255,N_2920,N_2980);
or U3256 (N_3256,N_2888,N_3110);
or U3257 (N_3257,N_3106,N_3170);
or U3258 (N_3258,N_3087,N_2825);
nor U3259 (N_3259,N_2900,N_3097);
nand U3260 (N_3260,N_3036,N_3059);
nor U3261 (N_3261,N_3000,N_3156);
nand U3262 (N_3262,N_3052,N_3033);
or U3263 (N_3263,N_2964,N_3103);
or U3264 (N_3264,N_3099,N_3173);
and U3265 (N_3265,N_3129,N_3005);
nand U3266 (N_3266,N_3138,N_3085);
and U3267 (N_3267,N_3001,N_3003);
or U3268 (N_3268,N_3072,N_3193);
and U3269 (N_3269,N_3075,N_2977);
nor U3270 (N_3270,N_2878,N_3013);
or U3271 (N_3271,N_3090,N_3146);
nor U3272 (N_3272,N_2876,N_2818);
and U3273 (N_3273,N_2925,N_3177);
nor U3274 (N_3274,N_3115,N_3088);
nor U3275 (N_3275,N_3045,N_2879);
nor U3276 (N_3276,N_2932,N_2948);
nand U3277 (N_3277,N_2960,N_2831);
and U3278 (N_3278,N_2974,N_3057);
or U3279 (N_3279,N_2931,N_2817);
and U3280 (N_3280,N_3017,N_3137);
and U3281 (N_3281,N_2918,N_2969);
and U3282 (N_3282,N_3091,N_3180);
and U3283 (N_3283,N_3159,N_2989);
and U3284 (N_3284,N_3089,N_2894);
or U3285 (N_3285,N_2820,N_2943);
or U3286 (N_3286,N_2942,N_3131);
nand U3287 (N_3287,N_3056,N_2994);
nand U3288 (N_3288,N_3198,N_2975);
nor U3289 (N_3289,N_3157,N_3169);
or U3290 (N_3290,N_2839,N_2824);
nor U3291 (N_3291,N_3030,N_3160);
nand U3292 (N_3292,N_3122,N_2907);
nand U3293 (N_3293,N_2886,N_2952);
nor U3294 (N_3294,N_3023,N_3139);
nor U3295 (N_3295,N_3171,N_3164);
and U3296 (N_3296,N_2805,N_2940);
nor U3297 (N_3297,N_3009,N_3181);
or U3298 (N_3298,N_2865,N_2962);
and U3299 (N_3299,N_2853,N_3196);
and U3300 (N_3300,N_3081,N_2812);
nand U3301 (N_3301,N_3002,N_2987);
or U3302 (N_3302,N_3020,N_2847);
nand U3303 (N_3303,N_3078,N_3098);
nand U3304 (N_3304,N_2827,N_3104);
and U3305 (N_3305,N_2983,N_2936);
and U3306 (N_3306,N_2946,N_2973);
or U3307 (N_3307,N_2961,N_3152);
nor U3308 (N_3308,N_3061,N_2908);
nand U3309 (N_3309,N_2883,N_2866);
or U3310 (N_3310,N_3069,N_3158);
or U3311 (N_3311,N_3168,N_2979);
and U3312 (N_3312,N_3166,N_2998);
or U3313 (N_3313,N_3021,N_2835);
or U3314 (N_3314,N_2806,N_3144);
nor U3315 (N_3315,N_3187,N_3150);
or U3316 (N_3316,N_2833,N_2804);
nand U3317 (N_3317,N_3186,N_3175);
and U3318 (N_3318,N_2809,N_2939);
and U3319 (N_3319,N_2923,N_2890);
nor U3320 (N_3320,N_2863,N_3182);
and U3321 (N_3321,N_3128,N_2875);
and U3322 (N_3322,N_2928,N_3022);
xnor U3323 (N_3323,N_2821,N_3195);
or U3324 (N_3324,N_3142,N_3176);
nor U3325 (N_3325,N_3188,N_3161);
nor U3326 (N_3326,N_2884,N_3190);
nor U3327 (N_3327,N_2972,N_2956);
and U3328 (N_3328,N_3051,N_2914);
or U3329 (N_3329,N_3162,N_2924);
or U3330 (N_3330,N_2988,N_2815);
and U3331 (N_3331,N_2954,N_3035);
nor U3332 (N_3332,N_3027,N_3080);
nor U3333 (N_3333,N_3111,N_3058);
nor U3334 (N_3334,N_3011,N_2917);
and U3335 (N_3335,N_3100,N_2945);
and U3336 (N_3336,N_3118,N_2869);
or U3337 (N_3337,N_3070,N_2844);
xor U3338 (N_3338,N_2893,N_2864);
nand U3339 (N_3339,N_2953,N_3132);
and U3340 (N_3340,N_2845,N_3185);
and U3341 (N_3341,N_3092,N_3102);
nor U3342 (N_3342,N_3074,N_3062);
nand U3343 (N_3343,N_2813,N_3189);
nand U3344 (N_3344,N_2933,N_3134);
or U3345 (N_3345,N_3064,N_3153);
and U3346 (N_3346,N_3066,N_2851);
or U3347 (N_3347,N_3079,N_3120);
or U3348 (N_3348,N_3019,N_2992);
or U3349 (N_3349,N_2913,N_2823);
or U3350 (N_3350,N_2889,N_2911);
nor U3351 (N_3351,N_2991,N_3094);
nor U3352 (N_3352,N_2861,N_3192);
nand U3353 (N_3353,N_3014,N_3184);
nand U3354 (N_3354,N_2967,N_3154);
and U3355 (N_3355,N_2995,N_2842);
and U3356 (N_3356,N_3038,N_3040);
nor U3357 (N_3357,N_3135,N_2986);
and U3358 (N_3358,N_2895,N_2857);
and U3359 (N_3359,N_3096,N_2860);
nor U3360 (N_3360,N_3039,N_3174);
or U3361 (N_3361,N_2926,N_3083);
and U3362 (N_3362,N_3172,N_2985);
nand U3363 (N_3363,N_2950,N_3105);
and U3364 (N_3364,N_3151,N_3183);
nor U3365 (N_3365,N_2984,N_3136);
nor U3366 (N_3366,N_2807,N_2916);
or U3367 (N_3367,N_2930,N_2873);
nand U3368 (N_3368,N_3143,N_3108);
or U3369 (N_3369,N_2846,N_3163);
and U3370 (N_3370,N_2915,N_3055);
nor U3371 (N_3371,N_2904,N_3199);
nand U3372 (N_3372,N_2836,N_3046);
and U3373 (N_3373,N_2850,N_3086);
and U3374 (N_3374,N_2996,N_2803);
nand U3375 (N_3375,N_2990,N_3053);
or U3376 (N_3376,N_2901,N_3140);
and U3377 (N_3377,N_3194,N_3124);
or U3378 (N_3378,N_2941,N_2858);
or U3379 (N_3379,N_2849,N_3026);
or U3380 (N_3380,N_3044,N_3025);
xor U3381 (N_3381,N_3117,N_3126);
nor U3382 (N_3382,N_3095,N_2947);
and U3383 (N_3383,N_3178,N_2838);
nand U3384 (N_3384,N_2880,N_2802);
nand U3385 (N_3385,N_2944,N_3109);
or U3386 (N_3386,N_2832,N_2982);
nor U3387 (N_3387,N_2949,N_2898);
or U3388 (N_3388,N_3197,N_2997);
nor U3389 (N_3389,N_2800,N_2837);
or U3390 (N_3390,N_2899,N_2822);
nand U3391 (N_3391,N_2965,N_2862);
or U3392 (N_3392,N_3093,N_3114);
or U3393 (N_3393,N_3112,N_3031);
and U3394 (N_3394,N_2966,N_3060);
or U3395 (N_3395,N_2902,N_3133);
and U3396 (N_3396,N_2993,N_3012);
nand U3397 (N_3397,N_3032,N_3148);
nand U3398 (N_3398,N_2958,N_2919);
and U3399 (N_3399,N_3010,N_2828);
nor U3400 (N_3400,N_3058,N_2948);
nor U3401 (N_3401,N_3120,N_2886);
nand U3402 (N_3402,N_3148,N_3171);
nor U3403 (N_3403,N_3094,N_3176);
nand U3404 (N_3404,N_2975,N_2861);
nor U3405 (N_3405,N_3066,N_3107);
and U3406 (N_3406,N_2825,N_3102);
nor U3407 (N_3407,N_2859,N_3027);
nor U3408 (N_3408,N_2917,N_2831);
and U3409 (N_3409,N_3123,N_3186);
nand U3410 (N_3410,N_3004,N_3099);
or U3411 (N_3411,N_3162,N_2935);
and U3412 (N_3412,N_3067,N_3084);
and U3413 (N_3413,N_3048,N_2827);
nor U3414 (N_3414,N_3156,N_2951);
nor U3415 (N_3415,N_3123,N_3051);
and U3416 (N_3416,N_3075,N_2863);
nand U3417 (N_3417,N_3143,N_3193);
nor U3418 (N_3418,N_2905,N_3026);
nand U3419 (N_3419,N_2960,N_2827);
or U3420 (N_3420,N_2963,N_2843);
nor U3421 (N_3421,N_3121,N_3148);
nand U3422 (N_3422,N_3172,N_2930);
nand U3423 (N_3423,N_3146,N_3133);
nand U3424 (N_3424,N_3139,N_3189);
xnor U3425 (N_3425,N_2844,N_3096);
nor U3426 (N_3426,N_3001,N_2914);
or U3427 (N_3427,N_3168,N_2839);
and U3428 (N_3428,N_3098,N_3120);
nor U3429 (N_3429,N_2896,N_2819);
nor U3430 (N_3430,N_3081,N_3190);
nand U3431 (N_3431,N_2913,N_3095);
nand U3432 (N_3432,N_2848,N_2894);
nand U3433 (N_3433,N_3002,N_3140);
nand U3434 (N_3434,N_3194,N_2974);
nand U3435 (N_3435,N_2886,N_3155);
nor U3436 (N_3436,N_3137,N_2850);
nand U3437 (N_3437,N_3136,N_3193);
nor U3438 (N_3438,N_2899,N_2811);
or U3439 (N_3439,N_2995,N_2849);
nand U3440 (N_3440,N_3090,N_2854);
and U3441 (N_3441,N_3186,N_2978);
nand U3442 (N_3442,N_3172,N_3059);
and U3443 (N_3443,N_3100,N_2915);
and U3444 (N_3444,N_2970,N_3194);
nor U3445 (N_3445,N_2893,N_3023);
nand U3446 (N_3446,N_3189,N_3132);
nand U3447 (N_3447,N_2851,N_3135);
nand U3448 (N_3448,N_2983,N_3130);
nand U3449 (N_3449,N_2889,N_2902);
nor U3450 (N_3450,N_2856,N_2913);
nand U3451 (N_3451,N_2894,N_3186);
nand U3452 (N_3452,N_3045,N_3123);
and U3453 (N_3453,N_3054,N_3031);
nor U3454 (N_3454,N_2976,N_2895);
nand U3455 (N_3455,N_2931,N_2859);
or U3456 (N_3456,N_2837,N_3198);
nor U3457 (N_3457,N_2871,N_2872);
or U3458 (N_3458,N_3184,N_3132);
nor U3459 (N_3459,N_2915,N_3066);
nand U3460 (N_3460,N_3073,N_3020);
nor U3461 (N_3461,N_2875,N_3135);
and U3462 (N_3462,N_3138,N_2863);
nand U3463 (N_3463,N_2808,N_2920);
and U3464 (N_3464,N_2847,N_3083);
and U3465 (N_3465,N_2945,N_2825);
or U3466 (N_3466,N_2874,N_2881);
or U3467 (N_3467,N_3128,N_2849);
and U3468 (N_3468,N_3147,N_2986);
nor U3469 (N_3469,N_2811,N_2955);
or U3470 (N_3470,N_3032,N_2891);
nand U3471 (N_3471,N_2939,N_3014);
nor U3472 (N_3472,N_3080,N_3120);
and U3473 (N_3473,N_2895,N_2856);
and U3474 (N_3474,N_3049,N_3179);
nand U3475 (N_3475,N_2967,N_2969);
or U3476 (N_3476,N_2927,N_2855);
and U3477 (N_3477,N_3151,N_2906);
nand U3478 (N_3478,N_3021,N_2967);
or U3479 (N_3479,N_3031,N_3066);
or U3480 (N_3480,N_2867,N_2985);
nand U3481 (N_3481,N_2963,N_2926);
or U3482 (N_3482,N_2899,N_3069);
nand U3483 (N_3483,N_2973,N_3049);
or U3484 (N_3484,N_3113,N_2818);
or U3485 (N_3485,N_3020,N_3152);
and U3486 (N_3486,N_3079,N_3073);
and U3487 (N_3487,N_2832,N_2991);
nand U3488 (N_3488,N_2814,N_3010);
nand U3489 (N_3489,N_3167,N_3150);
and U3490 (N_3490,N_2875,N_3057);
or U3491 (N_3491,N_3132,N_3091);
or U3492 (N_3492,N_3014,N_3161);
nand U3493 (N_3493,N_3135,N_2804);
nand U3494 (N_3494,N_3162,N_2833);
and U3495 (N_3495,N_2977,N_3152);
and U3496 (N_3496,N_2909,N_3089);
and U3497 (N_3497,N_2991,N_3111);
and U3498 (N_3498,N_3134,N_3063);
nand U3499 (N_3499,N_3000,N_3018);
nor U3500 (N_3500,N_2874,N_2893);
nand U3501 (N_3501,N_3063,N_2933);
nand U3502 (N_3502,N_3117,N_2867);
and U3503 (N_3503,N_2888,N_3121);
nor U3504 (N_3504,N_2947,N_2997);
and U3505 (N_3505,N_3150,N_2839);
nor U3506 (N_3506,N_2866,N_3086);
nor U3507 (N_3507,N_2806,N_2943);
nand U3508 (N_3508,N_3123,N_2926);
or U3509 (N_3509,N_3199,N_3026);
nand U3510 (N_3510,N_3189,N_3097);
and U3511 (N_3511,N_3103,N_3144);
and U3512 (N_3512,N_3071,N_3049);
nand U3513 (N_3513,N_3033,N_2808);
and U3514 (N_3514,N_2919,N_2898);
and U3515 (N_3515,N_2969,N_3198);
nor U3516 (N_3516,N_3137,N_2856);
nor U3517 (N_3517,N_3032,N_2847);
nand U3518 (N_3518,N_2878,N_3155);
and U3519 (N_3519,N_2965,N_2867);
and U3520 (N_3520,N_2810,N_3127);
and U3521 (N_3521,N_2834,N_2972);
nor U3522 (N_3522,N_2869,N_2854);
nand U3523 (N_3523,N_3186,N_2845);
and U3524 (N_3524,N_3131,N_3060);
or U3525 (N_3525,N_2836,N_2955);
nand U3526 (N_3526,N_2914,N_3042);
or U3527 (N_3527,N_2802,N_2901);
and U3528 (N_3528,N_2907,N_2930);
nand U3529 (N_3529,N_3068,N_3167);
nor U3530 (N_3530,N_3196,N_3059);
and U3531 (N_3531,N_2948,N_3032);
and U3532 (N_3532,N_2831,N_2978);
nand U3533 (N_3533,N_3036,N_2840);
and U3534 (N_3534,N_2853,N_2912);
nor U3535 (N_3535,N_3130,N_3039);
or U3536 (N_3536,N_2815,N_3079);
nand U3537 (N_3537,N_3016,N_3089);
nor U3538 (N_3538,N_3087,N_3127);
nor U3539 (N_3539,N_2823,N_3194);
and U3540 (N_3540,N_3025,N_3085);
nand U3541 (N_3541,N_2885,N_3092);
or U3542 (N_3542,N_2811,N_3121);
or U3543 (N_3543,N_3022,N_2882);
and U3544 (N_3544,N_3184,N_3147);
nand U3545 (N_3545,N_3133,N_2976);
or U3546 (N_3546,N_2886,N_2866);
nor U3547 (N_3547,N_3183,N_3024);
and U3548 (N_3548,N_2862,N_3170);
nand U3549 (N_3549,N_3044,N_3196);
nand U3550 (N_3550,N_3035,N_3171);
or U3551 (N_3551,N_2973,N_2846);
nand U3552 (N_3552,N_2877,N_2908);
and U3553 (N_3553,N_3104,N_2845);
nand U3554 (N_3554,N_2882,N_2966);
nor U3555 (N_3555,N_3056,N_2823);
and U3556 (N_3556,N_2879,N_2868);
nand U3557 (N_3557,N_3104,N_3098);
and U3558 (N_3558,N_2896,N_3180);
nor U3559 (N_3559,N_2800,N_3028);
nand U3560 (N_3560,N_2852,N_2959);
nor U3561 (N_3561,N_2904,N_2931);
nand U3562 (N_3562,N_3031,N_3008);
or U3563 (N_3563,N_2965,N_2927);
nand U3564 (N_3564,N_3104,N_2900);
and U3565 (N_3565,N_2946,N_2868);
or U3566 (N_3566,N_2909,N_2903);
nor U3567 (N_3567,N_3043,N_2862);
nand U3568 (N_3568,N_2869,N_2864);
nand U3569 (N_3569,N_2931,N_3021);
and U3570 (N_3570,N_2928,N_2864);
nand U3571 (N_3571,N_2885,N_3026);
xnor U3572 (N_3572,N_3051,N_3184);
nand U3573 (N_3573,N_2977,N_2929);
nor U3574 (N_3574,N_2918,N_2804);
and U3575 (N_3575,N_2926,N_3044);
nand U3576 (N_3576,N_3024,N_3040);
nor U3577 (N_3577,N_2808,N_3057);
or U3578 (N_3578,N_3126,N_3059);
nand U3579 (N_3579,N_2887,N_2857);
and U3580 (N_3580,N_3098,N_2877);
or U3581 (N_3581,N_2997,N_2868);
or U3582 (N_3582,N_2951,N_2830);
nand U3583 (N_3583,N_2845,N_3110);
nor U3584 (N_3584,N_3026,N_3138);
nor U3585 (N_3585,N_2893,N_3038);
and U3586 (N_3586,N_3052,N_2806);
nand U3587 (N_3587,N_2846,N_3125);
nor U3588 (N_3588,N_2929,N_3096);
and U3589 (N_3589,N_2991,N_3119);
nor U3590 (N_3590,N_3139,N_3097);
or U3591 (N_3591,N_2893,N_3094);
nand U3592 (N_3592,N_3009,N_2842);
and U3593 (N_3593,N_2914,N_3146);
nor U3594 (N_3594,N_3152,N_2964);
and U3595 (N_3595,N_3125,N_3020);
nand U3596 (N_3596,N_2803,N_2831);
xnor U3597 (N_3597,N_2854,N_3189);
nor U3598 (N_3598,N_2849,N_3056);
nand U3599 (N_3599,N_2992,N_3044);
or U3600 (N_3600,N_3485,N_3330);
nor U3601 (N_3601,N_3486,N_3325);
nor U3602 (N_3602,N_3461,N_3472);
or U3603 (N_3603,N_3535,N_3430);
and U3604 (N_3604,N_3455,N_3246);
and U3605 (N_3605,N_3326,N_3581);
nor U3606 (N_3606,N_3366,N_3551);
or U3607 (N_3607,N_3312,N_3560);
nand U3608 (N_3608,N_3211,N_3394);
or U3609 (N_3609,N_3360,N_3555);
nand U3610 (N_3610,N_3514,N_3241);
and U3611 (N_3611,N_3423,N_3414);
nand U3612 (N_3612,N_3559,N_3373);
and U3613 (N_3613,N_3565,N_3501);
nor U3614 (N_3614,N_3576,N_3213);
nand U3615 (N_3615,N_3517,N_3382);
and U3616 (N_3616,N_3331,N_3429);
nand U3617 (N_3617,N_3230,N_3309);
or U3618 (N_3618,N_3391,N_3410);
and U3619 (N_3619,N_3425,N_3537);
nor U3620 (N_3620,N_3324,N_3386);
nand U3621 (N_3621,N_3567,N_3436);
nand U3622 (N_3622,N_3541,N_3474);
nor U3623 (N_3623,N_3375,N_3315);
nor U3624 (N_3624,N_3573,N_3469);
and U3625 (N_3625,N_3287,N_3549);
nor U3626 (N_3626,N_3204,N_3243);
or U3627 (N_3627,N_3545,N_3362);
nand U3628 (N_3628,N_3282,N_3553);
nor U3629 (N_3629,N_3234,N_3371);
nand U3630 (N_3630,N_3589,N_3483);
nand U3631 (N_3631,N_3422,N_3277);
nand U3632 (N_3632,N_3363,N_3389);
or U3633 (N_3633,N_3550,N_3240);
nor U3634 (N_3634,N_3507,N_3540);
and U3635 (N_3635,N_3482,N_3340);
nor U3636 (N_3636,N_3520,N_3593);
and U3637 (N_3637,N_3281,N_3433);
nand U3638 (N_3638,N_3367,N_3294);
nor U3639 (N_3639,N_3488,N_3471);
nor U3640 (N_3640,N_3521,N_3466);
nand U3641 (N_3641,N_3300,N_3519);
nor U3642 (N_3642,N_3276,N_3395);
nor U3643 (N_3643,N_3529,N_3225);
or U3644 (N_3644,N_3359,N_3503);
or U3645 (N_3645,N_3558,N_3235);
and U3646 (N_3646,N_3310,N_3296);
and U3647 (N_3647,N_3491,N_3280);
and U3648 (N_3648,N_3318,N_3392);
nor U3649 (N_3649,N_3333,N_3413);
nor U3650 (N_3650,N_3271,N_3267);
nor U3651 (N_3651,N_3354,N_3297);
nor U3652 (N_3652,N_3278,N_3533);
or U3653 (N_3653,N_3512,N_3481);
or U3654 (N_3654,N_3334,N_3390);
nor U3655 (N_3655,N_3442,N_3323);
and U3656 (N_3656,N_3468,N_3252);
and U3657 (N_3657,N_3419,N_3238);
and U3658 (N_3658,N_3592,N_3272);
nand U3659 (N_3659,N_3254,N_3531);
and U3660 (N_3660,N_3229,N_3502);
and U3661 (N_3661,N_3227,N_3465);
or U3662 (N_3662,N_3292,N_3201);
nor U3663 (N_3663,N_3279,N_3351);
or U3664 (N_3664,N_3379,N_3307);
nor U3665 (N_3665,N_3506,N_3579);
and U3666 (N_3666,N_3350,N_3365);
nand U3667 (N_3667,N_3349,N_3441);
nand U3668 (N_3668,N_3329,N_3556);
nor U3669 (N_3669,N_3370,N_3591);
nand U3670 (N_3670,N_3437,N_3219);
or U3671 (N_3671,N_3223,N_3293);
and U3672 (N_3672,N_3364,N_3496);
nand U3673 (N_3673,N_3361,N_3343);
nor U3674 (N_3674,N_3299,N_3542);
nand U3675 (N_3675,N_3402,N_3202);
nand U3676 (N_3676,N_3274,N_3564);
nor U3677 (N_3677,N_3479,N_3554);
and U3678 (N_3678,N_3577,N_3221);
nand U3679 (N_3679,N_3495,N_3536);
and U3680 (N_3680,N_3303,N_3557);
nor U3681 (N_3681,N_3552,N_3291);
or U3682 (N_3682,N_3295,N_3408);
and U3683 (N_3683,N_3518,N_3245);
nor U3684 (N_3684,N_3448,N_3320);
and U3685 (N_3685,N_3269,N_3572);
nor U3686 (N_3686,N_3524,N_3358);
or U3687 (N_3687,N_3393,N_3590);
nor U3688 (N_3688,N_3215,N_3314);
nand U3689 (N_3689,N_3598,N_3490);
or U3690 (N_3690,N_3505,N_3369);
or U3691 (N_3691,N_3487,N_3248);
nor U3692 (N_3692,N_3427,N_3288);
or U3693 (N_3693,N_3377,N_3244);
nor U3694 (N_3694,N_3308,N_3439);
nand U3695 (N_3695,N_3453,N_3412);
nand U3696 (N_3696,N_3415,N_3527);
nand U3697 (N_3697,N_3440,N_3571);
nand U3698 (N_3698,N_3561,N_3345);
and U3699 (N_3699,N_3435,N_3339);
nor U3700 (N_3700,N_3275,N_3304);
or U3701 (N_3701,N_3568,N_3543);
and U3702 (N_3702,N_3477,N_3516);
or U3703 (N_3703,N_3336,N_3301);
nand U3704 (N_3704,N_3580,N_3268);
and U3705 (N_3705,N_3456,N_3473);
nand U3706 (N_3706,N_3587,N_3321);
nor U3707 (N_3707,N_3388,N_3284);
nand U3708 (N_3708,N_3526,N_3378);
and U3709 (N_3709,N_3584,N_3372);
or U3710 (N_3710,N_3508,N_3357);
and U3711 (N_3711,N_3255,N_3528);
nand U3712 (N_3712,N_3210,N_3417);
and U3713 (N_3713,N_3462,N_3327);
nand U3714 (N_3714,N_3588,N_3475);
or U3715 (N_3715,N_3217,N_3356);
nand U3716 (N_3716,N_3311,N_3319);
nand U3717 (N_3717,N_3398,N_3563);
nor U3718 (N_3718,N_3209,N_3266);
nand U3719 (N_3719,N_3237,N_3270);
nand U3720 (N_3720,N_3368,N_3205);
nor U3721 (N_3721,N_3444,N_3352);
and U3722 (N_3722,N_3504,N_3511);
and U3723 (N_3723,N_3214,N_3342);
or U3724 (N_3724,N_3497,N_3332);
nand U3725 (N_3725,N_3463,N_3353);
or U3726 (N_3726,N_3258,N_3431);
nor U3727 (N_3727,N_3374,N_3523);
and U3728 (N_3728,N_3348,N_3585);
nor U3729 (N_3729,N_3597,N_3416);
nor U3730 (N_3730,N_3344,N_3548);
nand U3731 (N_3731,N_3261,N_3257);
or U3732 (N_3732,N_3335,N_3233);
and U3733 (N_3733,N_3489,N_3546);
nor U3734 (N_3734,N_3400,N_3216);
or U3735 (N_3735,N_3260,N_3510);
or U3736 (N_3736,N_3207,N_3454);
nand U3737 (N_3737,N_3222,N_3457);
and U3738 (N_3738,N_3355,N_3224);
nor U3739 (N_3739,N_3409,N_3547);
and U3740 (N_3740,N_3265,N_3251);
and U3741 (N_3741,N_3498,N_3407);
nand U3742 (N_3742,N_3599,N_3494);
and U3743 (N_3743,N_3484,N_3263);
or U3744 (N_3744,N_3583,N_3380);
nand U3745 (N_3745,N_3458,N_3289);
or U3746 (N_3746,N_3247,N_3470);
and U3747 (N_3747,N_3316,N_3399);
nor U3748 (N_3748,N_3420,N_3438);
nand U3749 (N_3749,N_3434,N_3450);
nor U3750 (N_3750,N_3467,N_3544);
nor U3751 (N_3751,N_3259,N_3384);
and U3752 (N_3752,N_3500,N_3566);
nor U3753 (N_3753,N_3200,N_3534);
and U3754 (N_3754,N_3347,N_3586);
nand U3755 (N_3755,N_3232,N_3418);
nor U3756 (N_3756,N_3387,N_3273);
or U3757 (N_3757,N_3525,N_3404);
nand U3758 (N_3758,N_3250,N_3452);
or U3759 (N_3759,N_3403,N_3242);
nand U3760 (N_3760,N_3285,N_3478);
nor U3761 (N_3761,N_3539,N_3231);
nand U3762 (N_3762,N_3509,N_3396);
nor U3763 (N_3763,N_3569,N_3538);
nand U3764 (N_3764,N_3421,N_3451);
and U3765 (N_3765,N_3337,N_3212);
or U3766 (N_3766,N_3596,N_3447);
nand U3767 (N_3767,N_3218,N_3459);
and U3768 (N_3768,N_3515,N_3401);
and U3769 (N_3769,N_3432,N_3341);
or U3770 (N_3770,N_3239,N_3313);
or U3771 (N_3771,N_3253,N_3262);
nand U3772 (N_3772,N_3492,N_3405);
and U3773 (N_3773,N_3226,N_3397);
and U3774 (N_3774,N_3220,N_3290);
nand U3775 (N_3775,N_3522,N_3480);
and U3776 (N_3776,N_3446,N_3499);
nand U3777 (N_3777,N_3228,N_3383);
and U3778 (N_3778,N_3445,N_3283);
or U3779 (N_3779,N_3249,N_3574);
xnor U3780 (N_3780,N_3264,N_3208);
or U3781 (N_3781,N_3428,N_3305);
nand U3782 (N_3782,N_3532,N_3460);
nor U3783 (N_3783,N_3346,N_3582);
and U3784 (N_3784,N_3328,N_3411);
or U3785 (N_3785,N_3530,N_3578);
nand U3786 (N_3786,N_3449,N_3203);
and U3787 (N_3787,N_3575,N_3594);
nand U3788 (N_3788,N_3302,N_3256);
nand U3789 (N_3789,N_3306,N_3424);
nor U3790 (N_3790,N_3562,N_3376);
nor U3791 (N_3791,N_3426,N_3385);
or U3792 (N_3792,N_3298,N_3317);
xnor U3793 (N_3793,N_3322,N_3286);
and U3794 (N_3794,N_3338,N_3406);
nor U3795 (N_3795,N_3476,N_3570);
and U3796 (N_3796,N_3595,N_3513);
nand U3797 (N_3797,N_3206,N_3236);
and U3798 (N_3798,N_3464,N_3381);
xor U3799 (N_3799,N_3493,N_3443);
and U3800 (N_3800,N_3203,N_3363);
nor U3801 (N_3801,N_3277,N_3406);
or U3802 (N_3802,N_3366,N_3202);
nand U3803 (N_3803,N_3273,N_3357);
and U3804 (N_3804,N_3355,N_3451);
or U3805 (N_3805,N_3574,N_3295);
nand U3806 (N_3806,N_3398,N_3516);
nor U3807 (N_3807,N_3419,N_3316);
and U3808 (N_3808,N_3508,N_3479);
nor U3809 (N_3809,N_3410,N_3362);
nand U3810 (N_3810,N_3464,N_3237);
or U3811 (N_3811,N_3488,N_3468);
nand U3812 (N_3812,N_3330,N_3233);
nor U3813 (N_3813,N_3396,N_3279);
nor U3814 (N_3814,N_3412,N_3202);
nand U3815 (N_3815,N_3411,N_3225);
and U3816 (N_3816,N_3310,N_3536);
or U3817 (N_3817,N_3258,N_3556);
nand U3818 (N_3818,N_3506,N_3445);
and U3819 (N_3819,N_3409,N_3270);
nand U3820 (N_3820,N_3359,N_3528);
or U3821 (N_3821,N_3492,N_3530);
and U3822 (N_3822,N_3231,N_3374);
or U3823 (N_3823,N_3388,N_3346);
nand U3824 (N_3824,N_3307,N_3258);
nand U3825 (N_3825,N_3488,N_3315);
or U3826 (N_3826,N_3571,N_3351);
nand U3827 (N_3827,N_3345,N_3479);
or U3828 (N_3828,N_3460,N_3461);
or U3829 (N_3829,N_3510,N_3579);
nor U3830 (N_3830,N_3506,N_3230);
nor U3831 (N_3831,N_3235,N_3516);
and U3832 (N_3832,N_3527,N_3279);
or U3833 (N_3833,N_3214,N_3281);
nand U3834 (N_3834,N_3286,N_3388);
nand U3835 (N_3835,N_3532,N_3539);
and U3836 (N_3836,N_3250,N_3287);
or U3837 (N_3837,N_3217,N_3491);
or U3838 (N_3838,N_3558,N_3256);
and U3839 (N_3839,N_3241,N_3501);
nand U3840 (N_3840,N_3255,N_3312);
nand U3841 (N_3841,N_3284,N_3237);
and U3842 (N_3842,N_3551,N_3560);
nand U3843 (N_3843,N_3561,N_3582);
nor U3844 (N_3844,N_3366,N_3470);
nand U3845 (N_3845,N_3532,N_3440);
and U3846 (N_3846,N_3484,N_3214);
and U3847 (N_3847,N_3436,N_3253);
nor U3848 (N_3848,N_3359,N_3389);
xnor U3849 (N_3849,N_3577,N_3476);
xor U3850 (N_3850,N_3508,N_3322);
and U3851 (N_3851,N_3241,N_3282);
nand U3852 (N_3852,N_3226,N_3503);
or U3853 (N_3853,N_3264,N_3337);
nor U3854 (N_3854,N_3598,N_3316);
or U3855 (N_3855,N_3204,N_3273);
nand U3856 (N_3856,N_3218,N_3317);
nand U3857 (N_3857,N_3414,N_3592);
and U3858 (N_3858,N_3255,N_3595);
nand U3859 (N_3859,N_3522,N_3383);
and U3860 (N_3860,N_3455,N_3485);
nand U3861 (N_3861,N_3388,N_3354);
nand U3862 (N_3862,N_3528,N_3358);
or U3863 (N_3863,N_3453,N_3581);
nor U3864 (N_3864,N_3515,N_3300);
or U3865 (N_3865,N_3428,N_3241);
nor U3866 (N_3866,N_3506,N_3410);
nor U3867 (N_3867,N_3418,N_3456);
or U3868 (N_3868,N_3363,N_3592);
nand U3869 (N_3869,N_3505,N_3332);
or U3870 (N_3870,N_3338,N_3302);
xnor U3871 (N_3871,N_3514,N_3562);
or U3872 (N_3872,N_3345,N_3394);
nand U3873 (N_3873,N_3344,N_3575);
or U3874 (N_3874,N_3356,N_3284);
and U3875 (N_3875,N_3466,N_3569);
or U3876 (N_3876,N_3420,N_3434);
nand U3877 (N_3877,N_3393,N_3226);
nand U3878 (N_3878,N_3576,N_3238);
and U3879 (N_3879,N_3519,N_3523);
nand U3880 (N_3880,N_3267,N_3446);
nand U3881 (N_3881,N_3422,N_3352);
nor U3882 (N_3882,N_3217,N_3429);
and U3883 (N_3883,N_3557,N_3293);
or U3884 (N_3884,N_3351,N_3355);
or U3885 (N_3885,N_3360,N_3267);
nor U3886 (N_3886,N_3277,N_3495);
nand U3887 (N_3887,N_3555,N_3296);
xor U3888 (N_3888,N_3276,N_3477);
or U3889 (N_3889,N_3272,N_3265);
or U3890 (N_3890,N_3342,N_3563);
or U3891 (N_3891,N_3418,N_3235);
or U3892 (N_3892,N_3450,N_3518);
or U3893 (N_3893,N_3341,N_3375);
nor U3894 (N_3894,N_3287,N_3335);
and U3895 (N_3895,N_3461,N_3228);
nand U3896 (N_3896,N_3447,N_3343);
and U3897 (N_3897,N_3518,N_3349);
nor U3898 (N_3898,N_3541,N_3430);
and U3899 (N_3899,N_3269,N_3212);
nor U3900 (N_3900,N_3299,N_3236);
xnor U3901 (N_3901,N_3243,N_3571);
nor U3902 (N_3902,N_3342,N_3294);
nor U3903 (N_3903,N_3393,N_3566);
nor U3904 (N_3904,N_3327,N_3228);
and U3905 (N_3905,N_3283,N_3326);
and U3906 (N_3906,N_3379,N_3373);
nor U3907 (N_3907,N_3400,N_3563);
or U3908 (N_3908,N_3373,N_3272);
nand U3909 (N_3909,N_3292,N_3501);
and U3910 (N_3910,N_3568,N_3525);
nor U3911 (N_3911,N_3540,N_3401);
nor U3912 (N_3912,N_3567,N_3246);
nor U3913 (N_3913,N_3349,N_3323);
nand U3914 (N_3914,N_3542,N_3535);
or U3915 (N_3915,N_3404,N_3424);
and U3916 (N_3916,N_3305,N_3477);
or U3917 (N_3917,N_3349,N_3240);
nor U3918 (N_3918,N_3204,N_3510);
nor U3919 (N_3919,N_3400,N_3346);
or U3920 (N_3920,N_3524,N_3471);
and U3921 (N_3921,N_3421,N_3549);
or U3922 (N_3922,N_3475,N_3464);
or U3923 (N_3923,N_3439,N_3531);
nor U3924 (N_3924,N_3366,N_3259);
and U3925 (N_3925,N_3362,N_3307);
nor U3926 (N_3926,N_3275,N_3205);
and U3927 (N_3927,N_3229,N_3537);
or U3928 (N_3928,N_3259,N_3548);
and U3929 (N_3929,N_3343,N_3490);
xnor U3930 (N_3930,N_3479,N_3551);
and U3931 (N_3931,N_3455,N_3284);
or U3932 (N_3932,N_3416,N_3583);
and U3933 (N_3933,N_3224,N_3373);
or U3934 (N_3934,N_3571,N_3360);
nor U3935 (N_3935,N_3247,N_3553);
nor U3936 (N_3936,N_3284,N_3329);
nand U3937 (N_3937,N_3417,N_3258);
or U3938 (N_3938,N_3582,N_3569);
or U3939 (N_3939,N_3473,N_3528);
nand U3940 (N_3940,N_3242,N_3574);
and U3941 (N_3941,N_3592,N_3554);
or U3942 (N_3942,N_3363,N_3354);
and U3943 (N_3943,N_3523,N_3515);
or U3944 (N_3944,N_3574,N_3320);
nand U3945 (N_3945,N_3565,N_3325);
nor U3946 (N_3946,N_3478,N_3248);
nand U3947 (N_3947,N_3347,N_3214);
and U3948 (N_3948,N_3245,N_3305);
or U3949 (N_3949,N_3506,N_3415);
nor U3950 (N_3950,N_3481,N_3257);
or U3951 (N_3951,N_3514,N_3340);
and U3952 (N_3952,N_3594,N_3261);
nor U3953 (N_3953,N_3562,N_3290);
and U3954 (N_3954,N_3465,N_3200);
nand U3955 (N_3955,N_3332,N_3282);
or U3956 (N_3956,N_3232,N_3386);
or U3957 (N_3957,N_3427,N_3220);
nor U3958 (N_3958,N_3284,N_3381);
or U3959 (N_3959,N_3335,N_3239);
and U3960 (N_3960,N_3246,N_3579);
or U3961 (N_3961,N_3303,N_3295);
nand U3962 (N_3962,N_3307,N_3245);
nor U3963 (N_3963,N_3520,N_3331);
or U3964 (N_3964,N_3563,N_3349);
nor U3965 (N_3965,N_3443,N_3272);
or U3966 (N_3966,N_3484,N_3483);
or U3967 (N_3967,N_3488,N_3484);
nand U3968 (N_3968,N_3344,N_3222);
nor U3969 (N_3969,N_3534,N_3247);
or U3970 (N_3970,N_3489,N_3224);
nor U3971 (N_3971,N_3283,N_3486);
or U3972 (N_3972,N_3533,N_3516);
nand U3973 (N_3973,N_3534,N_3322);
nand U3974 (N_3974,N_3231,N_3215);
and U3975 (N_3975,N_3231,N_3245);
and U3976 (N_3976,N_3288,N_3548);
nor U3977 (N_3977,N_3219,N_3394);
or U3978 (N_3978,N_3401,N_3542);
or U3979 (N_3979,N_3543,N_3467);
nand U3980 (N_3980,N_3443,N_3319);
and U3981 (N_3981,N_3442,N_3475);
nor U3982 (N_3982,N_3567,N_3403);
nand U3983 (N_3983,N_3445,N_3382);
or U3984 (N_3984,N_3251,N_3369);
and U3985 (N_3985,N_3397,N_3526);
or U3986 (N_3986,N_3505,N_3389);
nor U3987 (N_3987,N_3276,N_3417);
and U3988 (N_3988,N_3438,N_3378);
xor U3989 (N_3989,N_3542,N_3352);
nand U3990 (N_3990,N_3371,N_3481);
xnor U3991 (N_3991,N_3362,N_3248);
or U3992 (N_3992,N_3296,N_3301);
nand U3993 (N_3993,N_3543,N_3247);
nand U3994 (N_3994,N_3220,N_3251);
or U3995 (N_3995,N_3536,N_3241);
and U3996 (N_3996,N_3466,N_3587);
nand U3997 (N_3997,N_3554,N_3358);
and U3998 (N_3998,N_3368,N_3396);
nand U3999 (N_3999,N_3410,N_3517);
and U4000 (N_4000,N_3743,N_3927);
and U4001 (N_4001,N_3991,N_3898);
xor U4002 (N_4002,N_3614,N_3651);
nand U4003 (N_4003,N_3807,N_3628);
nor U4004 (N_4004,N_3910,N_3908);
or U4005 (N_4005,N_3709,N_3730);
or U4006 (N_4006,N_3879,N_3600);
nor U4007 (N_4007,N_3876,N_3906);
nor U4008 (N_4008,N_3886,N_3601);
and U4009 (N_4009,N_3641,N_3695);
nand U4010 (N_4010,N_3683,N_3797);
nor U4011 (N_4011,N_3759,N_3720);
nand U4012 (N_4012,N_3928,N_3698);
nand U4013 (N_4013,N_3737,N_3831);
nand U4014 (N_4014,N_3629,N_3657);
nand U4015 (N_4015,N_3659,N_3904);
xor U4016 (N_4016,N_3922,N_3655);
nand U4017 (N_4017,N_3648,N_3633);
nor U4018 (N_4018,N_3757,N_3635);
or U4019 (N_4019,N_3672,N_3630);
and U4020 (N_4020,N_3794,N_3626);
and U4021 (N_4021,N_3692,N_3942);
and U4022 (N_4022,N_3804,N_3950);
or U4023 (N_4023,N_3694,N_3864);
nand U4024 (N_4024,N_3845,N_3682);
nand U4025 (N_4025,N_3763,N_3893);
nor U4026 (N_4026,N_3962,N_3716);
and U4027 (N_4027,N_3812,N_3616);
nand U4028 (N_4028,N_3919,N_3832);
and U4029 (N_4029,N_3921,N_3790);
nand U4030 (N_4030,N_3636,N_3981);
nand U4031 (N_4031,N_3917,N_3912);
and U4032 (N_4032,N_3913,N_3838);
and U4033 (N_4033,N_3795,N_3733);
nand U4034 (N_4034,N_3740,N_3666);
nor U4035 (N_4035,N_3693,N_3789);
or U4036 (N_4036,N_3894,N_3949);
or U4037 (N_4037,N_3829,N_3791);
or U4038 (N_4038,N_3880,N_3788);
nor U4039 (N_4039,N_3994,N_3758);
nand U4040 (N_4040,N_3966,N_3806);
and U4041 (N_4041,N_3847,N_3973);
and U4042 (N_4042,N_3990,N_3982);
and U4043 (N_4043,N_3715,N_3817);
nor U4044 (N_4044,N_3849,N_3874);
xnor U4045 (N_4045,N_3959,N_3933);
nand U4046 (N_4046,N_3739,N_3895);
nor U4047 (N_4047,N_3731,N_3840);
or U4048 (N_4048,N_3735,N_3800);
or U4049 (N_4049,N_3798,N_3852);
or U4050 (N_4050,N_3649,N_3808);
or U4051 (N_4051,N_3993,N_3604);
nand U4052 (N_4052,N_3602,N_3940);
nor U4053 (N_4053,N_3941,N_3680);
and U4054 (N_4054,N_3786,N_3717);
and U4055 (N_4055,N_3667,N_3843);
or U4056 (N_4056,N_3610,N_3955);
nor U4057 (N_4057,N_3828,N_3686);
nor U4058 (N_4058,N_3761,N_3988);
nand U4059 (N_4059,N_3748,N_3664);
nand U4060 (N_4060,N_3859,N_3810);
nor U4061 (N_4061,N_3760,N_3780);
nand U4062 (N_4062,N_3678,N_3677);
and U4063 (N_4063,N_3818,N_3668);
or U4064 (N_4064,N_3764,N_3856);
nor U4065 (N_4065,N_3873,N_3833);
nand U4066 (N_4066,N_3932,N_3699);
or U4067 (N_4067,N_3618,N_3884);
and U4068 (N_4068,N_3696,N_3839);
nand U4069 (N_4069,N_3937,N_3821);
or U4070 (N_4070,N_3768,N_3796);
or U4071 (N_4071,N_3944,N_3957);
or U4072 (N_4072,N_3914,N_3714);
nand U4073 (N_4073,N_3911,N_3787);
or U4074 (N_4074,N_3813,N_3983);
nor U4075 (N_4075,N_3647,N_3650);
nand U4076 (N_4076,N_3861,N_3638);
nand U4077 (N_4077,N_3987,N_3722);
and U4078 (N_4078,N_3738,N_3929);
nand U4079 (N_4079,N_3685,N_3712);
nand U4080 (N_4080,N_3996,N_3784);
nor U4081 (N_4081,N_3968,N_3785);
and U4082 (N_4082,N_3971,N_3984);
or U4083 (N_4083,N_3605,N_3654);
nor U4084 (N_4084,N_3671,N_3896);
nand U4085 (N_4085,N_3972,N_3824);
nor U4086 (N_4086,N_3701,N_3623);
or U4087 (N_4087,N_3844,N_3954);
nand U4088 (N_4088,N_3815,N_3621);
and U4089 (N_4089,N_3872,N_3891);
nand U4090 (N_4090,N_3749,N_3975);
or U4091 (N_4091,N_3920,N_3985);
or U4092 (N_4092,N_3608,N_3978);
nand U4093 (N_4093,N_3943,N_3900);
and U4094 (N_4094,N_3977,N_3903);
and U4095 (N_4095,N_3744,N_3816);
nand U4096 (N_4096,N_3742,N_3639);
and U4097 (N_4097,N_3661,N_3857);
or U4098 (N_4098,N_3835,N_3897);
and U4099 (N_4099,N_3811,N_3774);
or U4100 (N_4100,N_3805,N_3727);
nand U4101 (N_4101,N_3837,N_3842);
or U4102 (N_4102,N_3960,N_3756);
nand U4103 (N_4103,N_3643,N_3770);
nand U4104 (N_4104,N_3995,N_3860);
nand U4105 (N_4105,N_3925,N_3613);
nor U4106 (N_4106,N_3617,N_3889);
nor U4107 (N_4107,N_3778,N_3662);
nand U4108 (N_4108,N_3862,N_3705);
nor U4109 (N_4109,N_3866,N_3867);
and U4110 (N_4110,N_3938,N_3669);
or U4111 (N_4111,N_3826,N_3923);
nand U4112 (N_4112,N_3675,N_3974);
nor U4113 (N_4113,N_3724,N_3750);
or U4114 (N_4114,N_3706,N_3976);
nand U4115 (N_4115,N_3620,N_3939);
or U4116 (N_4116,N_3946,N_3931);
xor U4117 (N_4117,N_3707,N_3718);
nor U4118 (N_4118,N_3644,N_3631);
or U4119 (N_4119,N_3836,N_3710);
and U4120 (N_4120,N_3998,N_3745);
nor U4121 (N_4121,N_3902,N_3767);
xor U4122 (N_4122,N_3684,N_3734);
nand U4123 (N_4123,N_3640,N_3771);
and U4124 (N_4124,N_3704,N_3945);
nor U4125 (N_4125,N_3723,N_3765);
nor U4126 (N_4126,N_3690,N_3827);
nor U4127 (N_4127,N_3646,N_3689);
or U4128 (N_4128,N_3728,N_3766);
or U4129 (N_4129,N_3799,N_3848);
nor U4130 (N_4130,N_3642,N_3711);
and U4131 (N_4131,N_3772,N_3963);
and U4132 (N_4132,N_3951,N_3870);
and U4133 (N_4133,N_3907,N_3953);
or U4134 (N_4134,N_3703,N_3674);
and U4135 (N_4135,N_3634,N_3777);
and U4136 (N_4136,N_3887,N_3607);
nand U4137 (N_4137,N_3665,N_3980);
or U4138 (N_4138,N_3934,N_3736);
and U4139 (N_4139,N_3979,N_3809);
nand U4140 (N_4140,N_3964,N_3755);
and U4141 (N_4141,N_3606,N_3863);
nor U4142 (N_4142,N_3820,N_3881);
or U4143 (N_4143,N_3819,N_3782);
nor U4144 (N_4144,N_3776,N_3885);
or U4145 (N_4145,N_3658,N_3871);
or U4146 (N_4146,N_3846,N_3609);
or U4147 (N_4147,N_3901,N_3909);
nor U4148 (N_4148,N_3924,N_3992);
or U4149 (N_4149,N_3905,N_3823);
and U4150 (N_4150,N_3970,N_3632);
nand U4151 (N_4151,N_3700,N_3930);
or U4152 (N_4152,N_3769,N_3775);
nand U4153 (N_4153,N_3854,N_3673);
or U4154 (N_4154,N_3841,N_3753);
nor U4155 (N_4155,N_3726,N_3691);
nand U4156 (N_4156,N_3754,N_3679);
nor U4157 (N_4157,N_3869,N_3967);
and U4158 (N_4158,N_3624,N_3825);
nor U4159 (N_4159,N_3637,N_3725);
nand U4160 (N_4160,N_3802,N_3746);
nand U4161 (N_4161,N_3989,N_3697);
or U4162 (N_4162,N_3865,N_3947);
and U4163 (N_4163,N_3652,N_3779);
nor U4164 (N_4164,N_3858,N_3935);
and U4165 (N_4165,N_3916,N_3830);
or U4166 (N_4166,N_3969,N_3952);
or U4167 (N_4167,N_3702,N_3783);
nor U4168 (N_4168,N_3850,N_3752);
and U4169 (N_4169,N_3611,N_3965);
or U4170 (N_4170,N_3899,N_3708);
or U4171 (N_4171,N_3732,N_3868);
or U4172 (N_4172,N_3926,N_3801);
and U4173 (N_4173,N_3956,N_3822);
nor U4174 (N_4174,N_3663,N_3721);
nor U4175 (N_4175,N_3877,N_3762);
or U4176 (N_4176,N_3660,N_3803);
and U4177 (N_4177,N_3622,N_3936);
nand U4178 (N_4178,N_3882,N_3681);
or U4179 (N_4179,N_3645,N_3997);
nand U4180 (N_4180,N_3890,N_3948);
or U4181 (N_4181,N_3687,N_3688);
or U4182 (N_4182,N_3892,N_3792);
nand U4183 (N_4183,N_3851,N_3781);
and U4184 (N_4184,N_3670,N_3615);
nor U4185 (N_4185,N_3875,N_3999);
or U4186 (N_4186,N_3773,N_3888);
and U4187 (N_4187,N_3986,N_3878);
or U4188 (N_4188,N_3625,N_3814);
nand U4189 (N_4189,N_3729,N_3612);
nand U4190 (N_4190,N_3751,N_3603);
nand U4191 (N_4191,N_3918,N_3747);
xnor U4192 (N_4192,N_3719,N_3656);
and U4193 (N_4193,N_3958,N_3653);
nand U4194 (N_4194,N_3713,N_3741);
or U4195 (N_4195,N_3627,N_3961);
or U4196 (N_4196,N_3883,N_3676);
or U4197 (N_4197,N_3915,N_3793);
nor U4198 (N_4198,N_3855,N_3619);
nand U4199 (N_4199,N_3834,N_3853);
and U4200 (N_4200,N_3992,N_3974);
nand U4201 (N_4201,N_3941,N_3995);
nor U4202 (N_4202,N_3766,N_3909);
or U4203 (N_4203,N_3763,N_3707);
or U4204 (N_4204,N_3732,N_3979);
nand U4205 (N_4205,N_3714,N_3939);
nand U4206 (N_4206,N_3924,N_3604);
nand U4207 (N_4207,N_3807,N_3794);
or U4208 (N_4208,N_3876,N_3712);
or U4209 (N_4209,N_3992,N_3947);
and U4210 (N_4210,N_3729,N_3689);
or U4211 (N_4211,N_3666,N_3877);
nor U4212 (N_4212,N_3766,N_3641);
xor U4213 (N_4213,N_3916,N_3744);
or U4214 (N_4214,N_3927,N_3679);
and U4215 (N_4215,N_3669,N_3824);
nor U4216 (N_4216,N_3841,N_3961);
nand U4217 (N_4217,N_3666,N_3676);
nand U4218 (N_4218,N_3761,N_3644);
nor U4219 (N_4219,N_3753,N_3631);
and U4220 (N_4220,N_3799,N_3890);
xnor U4221 (N_4221,N_3763,N_3646);
or U4222 (N_4222,N_3804,N_3693);
and U4223 (N_4223,N_3714,N_3696);
and U4224 (N_4224,N_3661,N_3663);
nand U4225 (N_4225,N_3986,N_3670);
nor U4226 (N_4226,N_3885,N_3710);
and U4227 (N_4227,N_3926,N_3614);
or U4228 (N_4228,N_3616,N_3762);
and U4229 (N_4229,N_3923,N_3989);
or U4230 (N_4230,N_3885,N_3896);
and U4231 (N_4231,N_3986,N_3886);
nor U4232 (N_4232,N_3814,N_3970);
and U4233 (N_4233,N_3828,N_3727);
and U4234 (N_4234,N_3776,N_3722);
nor U4235 (N_4235,N_3859,N_3781);
nand U4236 (N_4236,N_3901,N_3978);
and U4237 (N_4237,N_3864,N_3898);
nor U4238 (N_4238,N_3723,N_3621);
or U4239 (N_4239,N_3687,N_3856);
or U4240 (N_4240,N_3948,N_3854);
nand U4241 (N_4241,N_3904,N_3775);
nand U4242 (N_4242,N_3808,N_3813);
or U4243 (N_4243,N_3783,N_3770);
nor U4244 (N_4244,N_3613,N_3780);
nor U4245 (N_4245,N_3857,N_3842);
or U4246 (N_4246,N_3907,N_3761);
nor U4247 (N_4247,N_3753,N_3805);
or U4248 (N_4248,N_3894,N_3919);
nor U4249 (N_4249,N_3844,N_3852);
nand U4250 (N_4250,N_3685,N_3911);
or U4251 (N_4251,N_3981,N_3611);
and U4252 (N_4252,N_3980,N_3876);
nor U4253 (N_4253,N_3757,N_3981);
and U4254 (N_4254,N_3780,N_3833);
and U4255 (N_4255,N_3778,N_3981);
nand U4256 (N_4256,N_3611,N_3953);
nand U4257 (N_4257,N_3656,N_3663);
nor U4258 (N_4258,N_3832,N_3789);
or U4259 (N_4259,N_3917,N_3668);
and U4260 (N_4260,N_3921,N_3712);
and U4261 (N_4261,N_3702,N_3696);
nor U4262 (N_4262,N_3785,N_3762);
nand U4263 (N_4263,N_3612,N_3993);
xor U4264 (N_4264,N_3956,N_3864);
nand U4265 (N_4265,N_3758,N_3923);
nor U4266 (N_4266,N_3651,N_3787);
and U4267 (N_4267,N_3679,N_3745);
and U4268 (N_4268,N_3964,N_3791);
nand U4269 (N_4269,N_3950,N_3964);
or U4270 (N_4270,N_3917,N_3880);
or U4271 (N_4271,N_3646,N_3773);
nand U4272 (N_4272,N_3886,N_3934);
nand U4273 (N_4273,N_3670,N_3913);
and U4274 (N_4274,N_3915,N_3637);
nor U4275 (N_4275,N_3631,N_3880);
and U4276 (N_4276,N_3880,N_3930);
and U4277 (N_4277,N_3626,N_3974);
nor U4278 (N_4278,N_3654,N_3910);
and U4279 (N_4279,N_3675,N_3816);
nor U4280 (N_4280,N_3754,N_3944);
and U4281 (N_4281,N_3848,N_3952);
xnor U4282 (N_4282,N_3904,N_3710);
nor U4283 (N_4283,N_3703,N_3820);
nor U4284 (N_4284,N_3799,N_3990);
xnor U4285 (N_4285,N_3726,N_3617);
nor U4286 (N_4286,N_3820,N_3918);
or U4287 (N_4287,N_3756,N_3993);
and U4288 (N_4288,N_3648,N_3936);
nor U4289 (N_4289,N_3762,N_3900);
and U4290 (N_4290,N_3742,N_3624);
or U4291 (N_4291,N_3708,N_3986);
nor U4292 (N_4292,N_3766,N_3833);
nand U4293 (N_4293,N_3902,N_3715);
nand U4294 (N_4294,N_3880,N_3943);
nor U4295 (N_4295,N_3837,N_3657);
nor U4296 (N_4296,N_3657,N_3850);
and U4297 (N_4297,N_3798,N_3877);
or U4298 (N_4298,N_3916,N_3985);
nand U4299 (N_4299,N_3726,N_3821);
nor U4300 (N_4300,N_3834,N_3899);
nand U4301 (N_4301,N_3716,N_3649);
and U4302 (N_4302,N_3775,N_3964);
nand U4303 (N_4303,N_3723,N_3653);
nor U4304 (N_4304,N_3693,N_3892);
nand U4305 (N_4305,N_3820,N_3834);
and U4306 (N_4306,N_3872,N_3971);
and U4307 (N_4307,N_3741,N_3651);
or U4308 (N_4308,N_3816,N_3655);
nand U4309 (N_4309,N_3778,N_3792);
and U4310 (N_4310,N_3969,N_3946);
nor U4311 (N_4311,N_3881,N_3700);
or U4312 (N_4312,N_3843,N_3996);
nand U4313 (N_4313,N_3737,N_3910);
xor U4314 (N_4314,N_3858,N_3877);
nand U4315 (N_4315,N_3642,N_3759);
nand U4316 (N_4316,N_3863,N_3822);
nand U4317 (N_4317,N_3639,N_3752);
and U4318 (N_4318,N_3815,N_3779);
nand U4319 (N_4319,N_3784,N_3931);
or U4320 (N_4320,N_3927,N_3604);
nor U4321 (N_4321,N_3682,N_3941);
nor U4322 (N_4322,N_3794,N_3810);
or U4323 (N_4323,N_3840,N_3848);
and U4324 (N_4324,N_3951,N_3601);
nor U4325 (N_4325,N_3914,N_3993);
and U4326 (N_4326,N_3910,N_3620);
nand U4327 (N_4327,N_3609,N_3649);
and U4328 (N_4328,N_3753,N_3667);
nor U4329 (N_4329,N_3758,N_3896);
nand U4330 (N_4330,N_3957,N_3738);
and U4331 (N_4331,N_3928,N_3717);
nor U4332 (N_4332,N_3924,N_3975);
nor U4333 (N_4333,N_3615,N_3919);
nand U4334 (N_4334,N_3757,N_3835);
and U4335 (N_4335,N_3807,N_3616);
nand U4336 (N_4336,N_3999,N_3780);
and U4337 (N_4337,N_3728,N_3652);
nand U4338 (N_4338,N_3757,N_3622);
or U4339 (N_4339,N_3946,N_3844);
or U4340 (N_4340,N_3968,N_3954);
or U4341 (N_4341,N_3995,N_3724);
or U4342 (N_4342,N_3841,N_3635);
nand U4343 (N_4343,N_3663,N_3945);
nor U4344 (N_4344,N_3958,N_3859);
nand U4345 (N_4345,N_3906,N_3829);
or U4346 (N_4346,N_3847,N_3683);
nand U4347 (N_4347,N_3825,N_3721);
or U4348 (N_4348,N_3916,N_3971);
nor U4349 (N_4349,N_3922,N_3877);
or U4350 (N_4350,N_3740,N_3712);
nor U4351 (N_4351,N_3663,N_3607);
and U4352 (N_4352,N_3868,N_3666);
or U4353 (N_4353,N_3688,N_3684);
nand U4354 (N_4354,N_3745,N_3862);
nor U4355 (N_4355,N_3842,N_3850);
nand U4356 (N_4356,N_3637,N_3605);
and U4357 (N_4357,N_3867,N_3628);
or U4358 (N_4358,N_3959,N_3619);
and U4359 (N_4359,N_3654,N_3772);
nor U4360 (N_4360,N_3849,N_3602);
or U4361 (N_4361,N_3952,N_3862);
nor U4362 (N_4362,N_3912,N_3779);
nand U4363 (N_4363,N_3942,N_3976);
nor U4364 (N_4364,N_3655,N_3957);
nor U4365 (N_4365,N_3652,N_3970);
nand U4366 (N_4366,N_3754,N_3970);
nand U4367 (N_4367,N_3918,N_3937);
nor U4368 (N_4368,N_3942,N_3985);
and U4369 (N_4369,N_3622,N_3618);
or U4370 (N_4370,N_3607,N_3667);
or U4371 (N_4371,N_3944,N_3767);
xnor U4372 (N_4372,N_3803,N_3701);
or U4373 (N_4373,N_3651,N_3943);
nand U4374 (N_4374,N_3840,N_3601);
nor U4375 (N_4375,N_3624,N_3955);
nor U4376 (N_4376,N_3749,N_3651);
nand U4377 (N_4377,N_3885,N_3853);
or U4378 (N_4378,N_3985,N_3954);
or U4379 (N_4379,N_3722,N_3681);
nor U4380 (N_4380,N_3704,N_3684);
or U4381 (N_4381,N_3682,N_3715);
and U4382 (N_4382,N_3763,N_3692);
nand U4383 (N_4383,N_3665,N_3892);
or U4384 (N_4384,N_3710,N_3671);
or U4385 (N_4385,N_3876,N_3989);
or U4386 (N_4386,N_3841,N_3618);
nand U4387 (N_4387,N_3901,N_3809);
and U4388 (N_4388,N_3617,N_3978);
and U4389 (N_4389,N_3891,N_3726);
or U4390 (N_4390,N_3630,N_3810);
or U4391 (N_4391,N_3978,N_3938);
nor U4392 (N_4392,N_3620,N_3887);
nand U4393 (N_4393,N_3732,N_3643);
nor U4394 (N_4394,N_3911,N_3622);
or U4395 (N_4395,N_3737,N_3866);
nand U4396 (N_4396,N_3657,N_3757);
or U4397 (N_4397,N_3743,N_3705);
and U4398 (N_4398,N_3739,N_3732);
nor U4399 (N_4399,N_3705,N_3920);
nor U4400 (N_4400,N_4117,N_4202);
nor U4401 (N_4401,N_4394,N_4387);
nand U4402 (N_4402,N_4334,N_4335);
or U4403 (N_4403,N_4070,N_4255);
or U4404 (N_4404,N_4185,N_4177);
and U4405 (N_4405,N_4221,N_4010);
or U4406 (N_4406,N_4373,N_4140);
nand U4407 (N_4407,N_4307,N_4105);
or U4408 (N_4408,N_4289,N_4366);
and U4409 (N_4409,N_4098,N_4107);
nor U4410 (N_4410,N_4072,N_4302);
nand U4411 (N_4411,N_4088,N_4019);
or U4412 (N_4412,N_4186,N_4291);
nor U4413 (N_4413,N_4232,N_4397);
or U4414 (N_4414,N_4276,N_4339);
nand U4415 (N_4415,N_4026,N_4131);
and U4416 (N_4416,N_4112,N_4175);
or U4417 (N_4417,N_4049,N_4368);
nand U4418 (N_4418,N_4271,N_4003);
nand U4419 (N_4419,N_4294,N_4396);
nand U4420 (N_4420,N_4187,N_4250);
or U4421 (N_4421,N_4139,N_4369);
nand U4422 (N_4422,N_4133,N_4295);
and U4423 (N_4423,N_4310,N_4017);
nor U4424 (N_4424,N_4337,N_4297);
and U4425 (N_4425,N_4129,N_4227);
nor U4426 (N_4426,N_4304,N_4398);
or U4427 (N_4427,N_4382,N_4204);
or U4428 (N_4428,N_4053,N_4156);
nand U4429 (N_4429,N_4007,N_4096);
or U4430 (N_4430,N_4199,N_4343);
nand U4431 (N_4431,N_4050,N_4099);
nor U4432 (N_4432,N_4321,N_4004);
or U4433 (N_4433,N_4081,N_4196);
and U4434 (N_4434,N_4230,N_4306);
and U4435 (N_4435,N_4275,N_4277);
nor U4436 (N_4436,N_4192,N_4002);
or U4437 (N_4437,N_4205,N_4399);
and U4438 (N_4438,N_4358,N_4086);
nor U4439 (N_4439,N_4251,N_4249);
and U4440 (N_4440,N_4164,N_4032);
and U4441 (N_4441,N_4135,N_4386);
and U4442 (N_4442,N_4217,N_4154);
and U4443 (N_4443,N_4068,N_4045);
or U4444 (N_4444,N_4225,N_4312);
and U4445 (N_4445,N_4371,N_4273);
nor U4446 (N_4446,N_4319,N_4316);
nor U4447 (N_4447,N_4179,N_4143);
nor U4448 (N_4448,N_4285,N_4025);
nor U4449 (N_4449,N_4100,N_4137);
and U4450 (N_4450,N_4111,N_4159);
or U4451 (N_4451,N_4213,N_4238);
and U4452 (N_4452,N_4270,N_4278);
or U4453 (N_4453,N_4233,N_4092);
and U4454 (N_4454,N_4375,N_4360);
or U4455 (N_4455,N_4257,N_4327);
nor U4456 (N_4456,N_4364,N_4228);
nor U4457 (N_4457,N_4259,N_4191);
nand U4458 (N_4458,N_4128,N_4047);
and U4459 (N_4459,N_4207,N_4374);
nand U4460 (N_4460,N_4274,N_4006);
nand U4461 (N_4461,N_4020,N_4384);
or U4462 (N_4462,N_4036,N_4059);
nand U4463 (N_4463,N_4058,N_4342);
nand U4464 (N_4464,N_4283,N_4176);
nor U4465 (N_4465,N_4329,N_4314);
nor U4466 (N_4466,N_4318,N_4293);
nand U4467 (N_4467,N_4263,N_4121);
or U4468 (N_4468,N_4362,N_4180);
and U4469 (N_4469,N_4260,N_4231);
nand U4470 (N_4470,N_4039,N_4146);
and U4471 (N_4471,N_4357,N_4158);
nor U4472 (N_4472,N_4219,N_4269);
and U4473 (N_4473,N_4299,N_4073);
and U4474 (N_4474,N_4016,N_4051);
nor U4475 (N_4475,N_4163,N_4194);
nand U4476 (N_4476,N_4102,N_4011);
and U4477 (N_4477,N_4280,N_4153);
and U4478 (N_4478,N_4282,N_4125);
and U4479 (N_4479,N_4201,N_4168);
nand U4480 (N_4480,N_4268,N_4043);
and U4481 (N_4481,N_4152,N_4388);
nor U4482 (N_4482,N_4054,N_4355);
and U4483 (N_4483,N_4160,N_4008);
nor U4484 (N_4484,N_4169,N_4071);
nor U4485 (N_4485,N_4229,N_4091);
or U4486 (N_4486,N_4211,N_4038);
nand U4487 (N_4487,N_4347,N_4265);
and U4488 (N_4488,N_4042,N_4122);
nand U4489 (N_4489,N_4167,N_4029);
nor U4490 (N_4490,N_4005,N_4301);
and U4491 (N_4491,N_4113,N_4376);
or U4492 (N_4492,N_4134,N_4161);
nor U4493 (N_4493,N_4209,N_4220);
or U4494 (N_4494,N_4303,N_4350);
and U4495 (N_4495,N_4381,N_4315);
or U4496 (N_4496,N_4037,N_4150);
nand U4497 (N_4497,N_4206,N_4379);
and U4498 (N_4498,N_4361,N_4084);
and U4499 (N_4499,N_4279,N_4149);
or U4500 (N_4500,N_4021,N_4332);
nor U4501 (N_4501,N_4145,N_4322);
nor U4502 (N_4502,N_4246,N_4061);
and U4503 (N_4503,N_4261,N_4336);
or U4504 (N_4504,N_4223,N_4027);
nor U4505 (N_4505,N_4023,N_4383);
nor U4506 (N_4506,N_4344,N_4012);
or U4507 (N_4507,N_4138,N_4069);
nand U4508 (N_4508,N_4080,N_4123);
nor U4509 (N_4509,N_4198,N_4242);
nor U4510 (N_4510,N_4200,N_4028);
nor U4511 (N_4511,N_4181,N_4085);
nor U4512 (N_4512,N_4245,N_4262);
and U4513 (N_4513,N_4256,N_4093);
nand U4514 (N_4514,N_4190,N_4320);
or U4515 (N_4515,N_4142,N_4193);
nand U4516 (N_4516,N_4182,N_4252);
and U4517 (N_4517,N_4078,N_4309);
and U4518 (N_4518,N_4218,N_4130);
nor U4519 (N_4519,N_4022,N_4288);
nor U4520 (N_4520,N_4370,N_4147);
nor U4521 (N_4521,N_4377,N_4013);
or U4522 (N_4522,N_4264,N_4014);
nor U4523 (N_4523,N_4074,N_4241);
nand U4524 (N_4524,N_4041,N_4075);
nand U4525 (N_4525,N_4354,N_4046);
nor U4526 (N_4526,N_4248,N_4305);
or U4527 (N_4527,N_4330,N_4141);
nor U4528 (N_4528,N_4065,N_4018);
and U4529 (N_4529,N_4348,N_4067);
nor U4530 (N_4530,N_4101,N_4056);
and U4531 (N_4531,N_4247,N_4083);
or U4532 (N_4532,N_4151,N_4136);
and U4533 (N_4533,N_4254,N_4367);
nor U4534 (N_4534,N_4178,N_4338);
or U4535 (N_4535,N_4090,N_4298);
nand U4536 (N_4536,N_4203,N_4155);
nor U4537 (N_4537,N_4040,N_4237);
or U4538 (N_4538,N_4313,N_4033);
and U4539 (N_4539,N_4290,N_4015);
nand U4540 (N_4540,N_4210,N_4389);
nor U4541 (N_4541,N_4001,N_4226);
nor U4542 (N_4542,N_4195,N_4035);
and U4543 (N_4543,N_4393,N_4057);
nand U4544 (N_4544,N_4236,N_4267);
and U4545 (N_4545,N_4345,N_4224);
or U4546 (N_4546,N_4349,N_4171);
or U4547 (N_4547,N_4300,N_4044);
nand U4548 (N_4548,N_4243,N_4235);
or U4549 (N_4549,N_4391,N_4333);
or U4550 (N_4550,N_4031,N_4120);
nand U4551 (N_4551,N_4184,N_4258);
and U4552 (N_4552,N_4240,N_4030);
or U4553 (N_4553,N_4055,N_4234);
or U4554 (N_4554,N_4127,N_4000);
nand U4555 (N_4555,N_4115,N_4378);
and U4556 (N_4556,N_4183,N_4286);
and U4557 (N_4557,N_4341,N_4064);
and U4558 (N_4558,N_4077,N_4326);
nand U4559 (N_4559,N_4239,N_4188);
nor U4560 (N_4560,N_4272,N_4214);
xnor U4561 (N_4561,N_4317,N_4215);
nand U4562 (N_4562,N_4166,N_4363);
nand U4563 (N_4563,N_4063,N_4076);
nand U4564 (N_4564,N_4116,N_4385);
or U4565 (N_4565,N_4097,N_4108);
or U4566 (N_4566,N_4103,N_4359);
nor U4567 (N_4567,N_4222,N_4189);
and U4568 (N_4568,N_4052,N_4165);
nor U4569 (N_4569,N_4114,N_4060);
nor U4570 (N_4570,N_4340,N_4253);
nor U4571 (N_4571,N_4266,N_4144);
nand U4572 (N_4572,N_4287,N_4380);
or U4573 (N_4573,N_4082,N_4324);
and U4574 (N_4574,N_4048,N_4024);
or U4575 (N_4575,N_4172,N_4079);
nor U4576 (N_4576,N_4392,N_4009);
nor U4577 (N_4577,N_4132,N_4173);
or U4578 (N_4578,N_4104,N_4292);
nor U4579 (N_4579,N_4066,N_4365);
nor U4580 (N_4580,N_4148,N_4351);
or U4581 (N_4581,N_4170,N_4124);
nor U4582 (N_4582,N_4325,N_4331);
nor U4583 (N_4583,N_4281,N_4308);
and U4584 (N_4584,N_4390,N_4162);
nor U4585 (N_4585,N_4106,N_4284);
nor U4586 (N_4586,N_4174,N_4089);
or U4587 (N_4587,N_4296,N_4352);
and U4588 (N_4588,N_4353,N_4356);
nand U4589 (N_4589,N_4244,N_4197);
nand U4590 (N_4590,N_4118,N_4372);
nor U4591 (N_4591,N_4095,N_4216);
and U4592 (N_4592,N_4157,N_4034);
and U4593 (N_4593,N_4212,N_4094);
nor U4594 (N_4594,N_4109,N_4395);
nor U4595 (N_4595,N_4323,N_4311);
nor U4596 (N_4596,N_4087,N_4328);
nand U4597 (N_4597,N_4346,N_4119);
or U4598 (N_4598,N_4110,N_4062);
and U4599 (N_4599,N_4208,N_4126);
and U4600 (N_4600,N_4019,N_4058);
and U4601 (N_4601,N_4110,N_4111);
and U4602 (N_4602,N_4235,N_4282);
nor U4603 (N_4603,N_4318,N_4254);
nor U4604 (N_4604,N_4208,N_4173);
and U4605 (N_4605,N_4332,N_4203);
nor U4606 (N_4606,N_4263,N_4369);
nor U4607 (N_4607,N_4249,N_4398);
nor U4608 (N_4608,N_4119,N_4232);
and U4609 (N_4609,N_4280,N_4030);
nand U4610 (N_4610,N_4018,N_4349);
or U4611 (N_4611,N_4328,N_4279);
nor U4612 (N_4612,N_4203,N_4205);
nor U4613 (N_4613,N_4259,N_4292);
or U4614 (N_4614,N_4173,N_4307);
or U4615 (N_4615,N_4373,N_4054);
or U4616 (N_4616,N_4291,N_4237);
nand U4617 (N_4617,N_4144,N_4332);
nor U4618 (N_4618,N_4020,N_4211);
and U4619 (N_4619,N_4313,N_4354);
nor U4620 (N_4620,N_4281,N_4247);
nor U4621 (N_4621,N_4213,N_4195);
nor U4622 (N_4622,N_4191,N_4001);
or U4623 (N_4623,N_4014,N_4054);
or U4624 (N_4624,N_4110,N_4012);
and U4625 (N_4625,N_4039,N_4387);
nor U4626 (N_4626,N_4177,N_4088);
xnor U4627 (N_4627,N_4344,N_4213);
nor U4628 (N_4628,N_4047,N_4189);
and U4629 (N_4629,N_4121,N_4022);
and U4630 (N_4630,N_4328,N_4152);
and U4631 (N_4631,N_4006,N_4011);
nor U4632 (N_4632,N_4286,N_4384);
nor U4633 (N_4633,N_4272,N_4171);
nor U4634 (N_4634,N_4243,N_4161);
or U4635 (N_4635,N_4288,N_4229);
or U4636 (N_4636,N_4090,N_4331);
or U4637 (N_4637,N_4258,N_4146);
or U4638 (N_4638,N_4308,N_4317);
nor U4639 (N_4639,N_4188,N_4057);
and U4640 (N_4640,N_4243,N_4145);
nand U4641 (N_4641,N_4270,N_4399);
xnor U4642 (N_4642,N_4060,N_4056);
and U4643 (N_4643,N_4003,N_4243);
nand U4644 (N_4644,N_4365,N_4091);
or U4645 (N_4645,N_4361,N_4225);
and U4646 (N_4646,N_4381,N_4050);
and U4647 (N_4647,N_4013,N_4321);
nor U4648 (N_4648,N_4334,N_4223);
nor U4649 (N_4649,N_4027,N_4176);
and U4650 (N_4650,N_4245,N_4017);
nand U4651 (N_4651,N_4085,N_4138);
nor U4652 (N_4652,N_4304,N_4086);
and U4653 (N_4653,N_4211,N_4214);
nor U4654 (N_4654,N_4250,N_4007);
nor U4655 (N_4655,N_4069,N_4055);
nand U4656 (N_4656,N_4142,N_4263);
and U4657 (N_4657,N_4218,N_4251);
nor U4658 (N_4658,N_4136,N_4356);
nand U4659 (N_4659,N_4106,N_4169);
nand U4660 (N_4660,N_4138,N_4309);
nand U4661 (N_4661,N_4037,N_4382);
nor U4662 (N_4662,N_4305,N_4267);
and U4663 (N_4663,N_4372,N_4211);
nand U4664 (N_4664,N_4051,N_4061);
nand U4665 (N_4665,N_4340,N_4114);
nand U4666 (N_4666,N_4396,N_4383);
or U4667 (N_4667,N_4386,N_4205);
nand U4668 (N_4668,N_4180,N_4290);
and U4669 (N_4669,N_4303,N_4354);
nor U4670 (N_4670,N_4135,N_4084);
or U4671 (N_4671,N_4059,N_4159);
or U4672 (N_4672,N_4161,N_4364);
nor U4673 (N_4673,N_4091,N_4307);
and U4674 (N_4674,N_4243,N_4071);
or U4675 (N_4675,N_4151,N_4309);
nand U4676 (N_4676,N_4137,N_4308);
nor U4677 (N_4677,N_4231,N_4014);
and U4678 (N_4678,N_4014,N_4052);
or U4679 (N_4679,N_4360,N_4026);
nor U4680 (N_4680,N_4039,N_4166);
nand U4681 (N_4681,N_4346,N_4071);
or U4682 (N_4682,N_4318,N_4040);
or U4683 (N_4683,N_4321,N_4221);
nand U4684 (N_4684,N_4396,N_4324);
or U4685 (N_4685,N_4269,N_4220);
or U4686 (N_4686,N_4274,N_4034);
and U4687 (N_4687,N_4273,N_4280);
nor U4688 (N_4688,N_4138,N_4227);
and U4689 (N_4689,N_4274,N_4335);
nor U4690 (N_4690,N_4165,N_4099);
nand U4691 (N_4691,N_4235,N_4130);
nor U4692 (N_4692,N_4065,N_4185);
nor U4693 (N_4693,N_4266,N_4314);
or U4694 (N_4694,N_4042,N_4382);
nor U4695 (N_4695,N_4132,N_4232);
nor U4696 (N_4696,N_4182,N_4359);
or U4697 (N_4697,N_4042,N_4017);
and U4698 (N_4698,N_4144,N_4354);
nor U4699 (N_4699,N_4226,N_4158);
or U4700 (N_4700,N_4235,N_4145);
and U4701 (N_4701,N_4064,N_4035);
nand U4702 (N_4702,N_4264,N_4324);
nor U4703 (N_4703,N_4281,N_4219);
nand U4704 (N_4704,N_4015,N_4146);
and U4705 (N_4705,N_4279,N_4092);
and U4706 (N_4706,N_4361,N_4000);
nor U4707 (N_4707,N_4158,N_4214);
or U4708 (N_4708,N_4024,N_4046);
nand U4709 (N_4709,N_4398,N_4092);
or U4710 (N_4710,N_4034,N_4272);
nor U4711 (N_4711,N_4284,N_4386);
or U4712 (N_4712,N_4084,N_4216);
nand U4713 (N_4713,N_4353,N_4260);
nor U4714 (N_4714,N_4320,N_4375);
and U4715 (N_4715,N_4060,N_4140);
or U4716 (N_4716,N_4324,N_4174);
nand U4717 (N_4717,N_4220,N_4057);
nor U4718 (N_4718,N_4055,N_4205);
nor U4719 (N_4719,N_4105,N_4166);
nand U4720 (N_4720,N_4333,N_4233);
or U4721 (N_4721,N_4277,N_4117);
or U4722 (N_4722,N_4096,N_4334);
or U4723 (N_4723,N_4309,N_4147);
or U4724 (N_4724,N_4101,N_4355);
nor U4725 (N_4725,N_4204,N_4008);
nor U4726 (N_4726,N_4235,N_4098);
and U4727 (N_4727,N_4252,N_4207);
nor U4728 (N_4728,N_4241,N_4332);
nand U4729 (N_4729,N_4054,N_4351);
and U4730 (N_4730,N_4019,N_4182);
and U4731 (N_4731,N_4051,N_4106);
or U4732 (N_4732,N_4399,N_4125);
or U4733 (N_4733,N_4087,N_4335);
nand U4734 (N_4734,N_4002,N_4399);
nor U4735 (N_4735,N_4215,N_4377);
nand U4736 (N_4736,N_4370,N_4277);
nand U4737 (N_4737,N_4024,N_4125);
nand U4738 (N_4738,N_4055,N_4019);
and U4739 (N_4739,N_4014,N_4215);
nand U4740 (N_4740,N_4255,N_4188);
and U4741 (N_4741,N_4292,N_4028);
or U4742 (N_4742,N_4116,N_4208);
or U4743 (N_4743,N_4223,N_4052);
or U4744 (N_4744,N_4280,N_4307);
and U4745 (N_4745,N_4215,N_4249);
nor U4746 (N_4746,N_4182,N_4053);
nor U4747 (N_4747,N_4328,N_4052);
or U4748 (N_4748,N_4194,N_4391);
and U4749 (N_4749,N_4045,N_4053);
or U4750 (N_4750,N_4382,N_4224);
or U4751 (N_4751,N_4211,N_4380);
nor U4752 (N_4752,N_4164,N_4076);
or U4753 (N_4753,N_4188,N_4092);
and U4754 (N_4754,N_4117,N_4314);
xor U4755 (N_4755,N_4339,N_4137);
nor U4756 (N_4756,N_4185,N_4348);
nand U4757 (N_4757,N_4361,N_4178);
or U4758 (N_4758,N_4349,N_4012);
and U4759 (N_4759,N_4373,N_4071);
or U4760 (N_4760,N_4349,N_4069);
and U4761 (N_4761,N_4272,N_4225);
nand U4762 (N_4762,N_4236,N_4163);
nor U4763 (N_4763,N_4160,N_4110);
or U4764 (N_4764,N_4323,N_4191);
or U4765 (N_4765,N_4190,N_4075);
and U4766 (N_4766,N_4012,N_4026);
nor U4767 (N_4767,N_4169,N_4398);
nand U4768 (N_4768,N_4061,N_4068);
and U4769 (N_4769,N_4334,N_4137);
nand U4770 (N_4770,N_4077,N_4296);
or U4771 (N_4771,N_4003,N_4176);
or U4772 (N_4772,N_4328,N_4301);
nand U4773 (N_4773,N_4266,N_4267);
and U4774 (N_4774,N_4342,N_4003);
or U4775 (N_4775,N_4282,N_4201);
nand U4776 (N_4776,N_4370,N_4373);
nor U4777 (N_4777,N_4064,N_4102);
or U4778 (N_4778,N_4109,N_4101);
and U4779 (N_4779,N_4048,N_4385);
or U4780 (N_4780,N_4200,N_4109);
nor U4781 (N_4781,N_4300,N_4047);
nand U4782 (N_4782,N_4094,N_4040);
nand U4783 (N_4783,N_4290,N_4005);
or U4784 (N_4784,N_4220,N_4137);
nor U4785 (N_4785,N_4251,N_4312);
nand U4786 (N_4786,N_4172,N_4170);
or U4787 (N_4787,N_4133,N_4080);
xor U4788 (N_4788,N_4391,N_4299);
nor U4789 (N_4789,N_4276,N_4086);
and U4790 (N_4790,N_4316,N_4165);
nand U4791 (N_4791,N_4260,N_4011);
or U4792 (N_4792,N_4358,N_4224);
nor U4793 (N_4793,N_4110,N_4152);
nand U4794 (N_4794,N_4094,N_4308);
nor U4795 (N_4795,N_4100,N_4344);
nor U4796 (N_4796,N_4116,N_4175);
nand U4797 (N_4797,N_4066,N_4340);
nand U4798 (N_4798,N_4055,N_4321);
nand U4799 (N_4799,N_4139,N_4284);
or U4800 (N_4800,N_4514,N_4690);
and U4801 (N_4801,N_4696,N_4588);
or U4802 (N_4802,N_4668,N_4597);
or U4803 (N_4803,N_4438,N_4481);
or U4804 (N_4804,N_4626,N_4407);
or U4805 (N_4805,N_4758,N_4466);
or U4806 (N_4806,N_4491,N_4720);
or U4807 (N_4807,N_4700,N_4463);
nor U4808 (N_4808,N_4787,N_4691);
nand U4809 (N_4809,N_4506,N_4590);
or U4810 (N_4810,N_4759,N_4430);
or U4811 (N_4811,N_4693,N_4670);
nand U4812 (N_4812,N_4410,N_4423);
nor U4813 (N_4813,N_4744,N_4637);
and U4814 (N_4814,N_4684,N_4565);
nand U4815 (N_4815,N_4483,N_4685);
and U4816 (N_4816,N_4456,N_4538);
and U4817 (N_4817,N_4446,N_4639);
nand U4818 (N_4818,N_4716,N_4773);
nor U4819 (N_4819,N_4462,N_4476);
or U4820 (N_4820,N_4553,N_4678);
or U4821 (N_4821,N_4530,N_4757);
and U4822 (N_4822,N_4417,N_4624);
nor U4823 (N_4823,N_4558,N_4609);
nor U4824 (N_4824,N_4405,N_4534);
and U4825 (N_4825,N_4660,N_4733);
and U4826 (N_4826,N_4519,N_4513);
nand U4827 (N_4827,N_4420,N_4702);
nor U4828 (N_4828,N_4649,N_4642);
nor U4829 (N_4829,N_4630,N_4488);
or U4830 (N_4830,N_4546,N_4797);
nor U4831 (N_4831,N_4683,N_4613);
or U4832 (N_4832,N_4485,N_4544);
or U4833 (N_4833,N_4451,N_4748);
and U4834 (N_4834,N_4781,N_4646);
nand U4835 (N_4835,N_4728,N_4421);
nand U4836 (N_4836,N_4676,N_4494);
nor U4837 (N_4837,N_4658,N_4669);
and U4838 (N_4838,N_4708,N_4782);
and U4839 (N_4839,N_4478,N_4612);
nand U4840 (N_4840,N_4729,N_4507);
nor U4841 (N_4841,N_4634,N_4412);
nor U4842 (N_4842,N_4524,N_4661);
and U4843 (N_4843,N_4610,N_4448);
nand U4844 (N_4844,N_4433,N_4577);
and U4845 (N_4845,N_4400,N_4560);
nand U4846 (N_4846,N_4651,N_4486);
and U4847 (N_4847,N_4772,N_4694);
and U4848 (N_4848,N_4500,N_4585);
and U4849 (N_4849,N_4643,N_4575);
nand U4850 (N_4850,N_4746,N_4505);
nor U4851 (N_4851,N_4444,N_4686);
and U4852 (N_4852,N_4606,N_4440);
and U4853 (N_4853,N_4545,N_4449);
xor U4854 (N_4854,N_4452,N_4455);
nand U4855 (N_4855,N_4443,N_4523);
and U4856 (N_4856,N_4766,N_4755);
and U4857 (N_4857,N_4571,N_4719);
nand U4858 (N_4858,N_4460,N_4747);
nor U4859 (N_4859,N_4725,N_4600);
and U4860 (N_4860,N_4415,N_4434);
or U4861 (N_4861,N_4603,N_4601);
nor U4862 (N_4862,N_4619,N_4764);
and U4863 (N_4863,N_4663,N_4633);
and U4864 (N_4864,N_4536,N_4701);
or U4865 (N_4865,N_4672,N_4403);
and U4866 (N_4866,N_4548,N_4628);
and U4867 (N_4867,N_4713,N_4640);
and U4868 (N_4868,N_4586,N_4429);
nand U4869 (N_4869,N_4767,N_4742);
and U4870 (N_4870,N_4699,N_4705);
nand U4871 (N_4871,N_4707,N_4655);
nor U4872 (N_4872,N_4569,N_4441);
nor U4873 (N_4873,N_4795,N_4789);
nand U4874 (N_4874,N_4703,N_4475);
nand U4875 (N_4875,N_4512,N_4510);
nand U4876 (N_4876,N_4539,N_4471);
nand U4877 (N_4877,N_4490,N_4482);
nor U4878 (N_4878,N_4533,N_4776);
and U4879 (N_4879,N_4432,N_4419);
nor U4880 (N_4880,N_4673,N_4737);
and U4881 (N_4881,N_4579,N_4526);
and U4882 (N_4882,N_4679,N_4664);
and U4883 (N_4883,N_4454,N_4652);
or U4884 (N_4884,N_4557,N_4771);
nand U4885 (N_4885,N_4431,N_4469);
nand U4886 (N_4886,N_4723,N_4437);
nand U4887 (N_4887,N_4794,N_4743);
or U4888 (N_4888,N_4516,N_4498);
or U4889 (N_4889,N_4618,N_4559);
nor U4890 (N_4890,N_4641,N_4509);
and U4891 (N_4891,N_4402,N_4572);
nor U4892 (N_4892,N_4735,N_4711);
and U4893 (N_4893,N_4784,N_4654);
and U4894 (N_4894,N_4627,N_4650);
and U4895 (N_4895,N_4712,N_4793);
nor U4896 (N_4896,N_4616,N_4497);
and U4897 (N_4897,N_4467,N_4739);
nand U4898 (N_4898,N_4573,N_4422);
nor U4899 (N_4899,N_4518,N_4662);
and U4900 (N_4900,N_4477,N_4582);
nand U4901 (N_4901,N_4680,N_4542);
nor U4902 (N_4902,N_4620,N_4447);
nor U4903 (N_4903,N_4465,N_4774);
or U4904 (N_4904,N_4608,N_4681);
and U4905 (N_4905,N_4671,N_4593);
nand U4906 (N_4906,N_4749,N_4547);
nor U4907 (N_4907,N_4564,N_4621);
and U4908 (N_4908,N_4413,N_4647);
nand U4909 (N_4909,N_4583,N_4576);
nand U4910 (N_4910,N_4459,N_4788);
nand U4911 (N_4911,N_4710,N_4589);
and U4912 (N_4912,N_4763,N_4596);
or U4913 (N_4913,N_4525,N_4688);
or U4914 (N_4914,N_4734,N_4414);
nand U4915 (N_4915,N_4622,N_4574);
nand U4916 (N_4916,N_4515,N_4783);
or U4917 (N_4917,N_4499,N_4570);
nor U4918 (N_4918,N_4428,N_4566);
or U4919 (N_4919,N_4554,N_4648);
and U4920 (N_4920,N_4473,N_4468);
and U4921 (N_4921,N_4549,N_4552);
nor U4922 (N_4922,N_4792,N_4555);
nor U4923 (N_4923,N_4535,N_4561);
nand U4924 (N_4924,N_4635,N_4568);
or U4925 (N_4925,N_4731,N_4657);
or U4926 (N_4926,N_4595,N_4741);
and U4927 (N_4927,N_4632,N_4502);
and U4928 (N_4928,N_4541,N_4426);
nor U4929 (N_4929,N_4769,N_4745);
or U4930 (N_4930,N_4409,N_4472);
or U4931 (N_4931,N_4425,N_4487);
nand U4932 (N_4932,N_4580,N_4675);
nand U4933 (N_4933,N_4556,N_4581);
or U4934 (N_4934,N_4404,N_4697);
and U4935 (N_4935,N_4495,N_4695);
or U4936 (N_4936,N_4644,N_4464);
nor U4937 (N_4937,N_4717,N_4587);
or U4938 (N_4938,N_4592,N_4638);
or U4939 (N_4939,N_4718,N_4611);
nand U4940 (N_4940,N_4604,N_4562);
and U4941 (N_4941,N_4796,N_4479);
nand U4942 (N_4942,N_4520,N_4416);
nor U4943 (N_4943,N_4435,N_4602);
nand U4944 (N_4944,N_4521,N_4531);
or U4945 (N_4945,N_4424,N_4517);
and U4946 (N_4946,N_4605,N_4754);
or U4947 (N_4947,N_4474,N_4775);
or U4948 (N_4948,N_4779,N_4738);
xnor U4949 (N_4949,N_4724,N_4715);
and U4950 (N_4950,N_4625,N_4778);
and U4951 (N_4951,N_4687,N_4493);
or U4952 (N_4952,N_4427,N_4753);
or U4953 (N_4953,N_4677,N_4791);
and U4954 (N_4954,N_4511,N_4484);
and U4955 (N_4955,N_4631,N_4682);
nor U4956 (N_4956,N_4666,N_4522);
nor U4957 (N_4957,N_4615,N_4629);
and U4958 (N_4958,N_4768,N_4401);
and U4959 (N_4959,N_4667,N_4599);
and U4960 (N_4960,N_4756,N_4503);
and U4961 (N_4961,N_4798,N_4567);
nor U4962 (N_4962,N_4508,N_4765);
nor U4963 (N_4963,N_4411,N_4442);
or U4964 (N_4964,N_4761,N_4461);
nand U4965 (N_4965,N_4740,N_4752);
nand U4966 (N_4966,N_4480,N_4458);
or U4967 (N_4967,N_4607,N_4594);
or U4968 (N_4968,N_4450,N_4732);
and U4969 (N_4969,N_4551,N_4674);
nand U4970 (N_4970,N_4706,N_4408);
nor U4971 (N_4971,N_4750,N_4528);
and U4972 (N_4972,N_4501,N_4799);
nand U4973 (N_4973,N_4645,N_4698);
or U4974 (N_4974,N_4504,N_4418);
nor U4975 (N_4975,N_4656,N_4591);
or U4976 (N_4976,N_4496,N_4760);
nand U4977 (N_4977,N_4730,N_4653);
and U4978 (N_4978,N_4445,N_4785);
nand U4979 (N_4979,N_4540,N_4614);
nand U4980 (N_4980,N_4659,N_4721);
and U4981 (N_4981,N_4762,N_4736);
nor U4982 (N_4982,N_4436,N_4617);
or U4983 (N_4983,N_4489,N_4636);
or U4984 (N_4984,N_4692,N_4537);
or U4985 (N_4985,N_4790,N_4550);
nor U4986 (N_4986,N_4665,N_4470);
or U4987 (N_4987,N_4751,N_4770);
nand U4988 (N_4988,N_4786,N_4689);
nand U4989 (N_4989,N_4543,N_4527);
or U4990 (N_4990,N_4578,N_4722);
nor U4991 (N_4991,N_4714,N_4532);
nor U4992 (N_4992,N_4439,N_4529);
nor U4993 (N_4993,N_4777,N_4780);
and U4994 (N_4994,N_4709,N_4492);
and U4995 (N_4995,N_4457,N_4584);
nand U4996 (N_4996,N_4406,N_4623);
nor U4997 (N_4997,N_4598,N_4453);
nor U4998 (N_4998,N_4563,N_4726);
nor U4999 (N_4999,N_4704,N_4727);
and U5000 (N_5000,N_4793,N_4486);
and U5001 (N_5001,N_4635,N_4669);
nor U5002 (N_5002,N_4462,N_4703);
or U5003 (N_5003,N_4561,N_4513);
nor U5004 (N_5004,N_4474,N_4754);
or U5005 (N_5005,N_4632,N_4513);
xor U5006 (N_5006,N_4779,N_4708);
nand U5007 (N_5007,N_4670,N_4428);
nor U5008 (N_5008,N_4652,N_4458);
or U5009 (N_5009,N_4423,N_4477);
and U5010 (N_5010,N_4517,N_4764);
and U5011 (N_5011,N_4657,N_4582);
or U5012 (N_5012,N_4659,N_4795);
and U5013 (N_5013,N_4598,N_4429);
or U5014 (N_5014,N_4721,N_4677);
or U5015 (N_5015,N_4446,N_4450);
or U5016 (N_5016,N_4770,N_4714);
or U5017 (N_5017,N_4428,N_4793);
nand U5018 (N_5018,N_4622,N_4796);
nor U5019 (N_5019,N_4745,N_4535);
nor U5020 (N_5020,N_4683,N_4662);
or U5021 (N_5021,N_4419,N_4443);
nor U5022 (N_5022,N_4778,N_4451);
nand U5023 (N_5023,N_4477,N_4691);
and U5024 (N_5024,N_4511,N_4714);
nand U5025 (N_5025,N_4588,N_4599);
or U5026 (N_5026,N_4790,N_4727);
nand U5027 (N_5027,N_4712,N_4748);
and U5028 (N_5028,N_4748,N_4622);
and U5029 (N_5029,N_4624,N_4658);
nor U5030 (N_5030,N_4583,N_4561);
or U5031 (N_5031,N_4534,N_4461);
or U5032 (N_5032,N_4456,N_4461);
nand U5033 (N_5033,N_4530,N_4548);
nor U5034 (N_5034,N_4405,N_4481);
and U5035 (N_5035,N_4582,N_4787);
nor U5036 (N_5036,N_4733,N_4601);
nor U5037 (N_5037,N_4639,N_4524);
nand U5038 (N_5038,N_4474,N_4558);
or U5039 (N_5039,N_4721,N_4625);
nor U5040 (N_5040,N_4570,N_4417);
nand U5041 (N_5041,N_4575,N_4635);
nor U5042 (N_5042,N_4563,N_4769);
and U5043 (N_5043,N_4445,N_4620);
and U5044 (N_5044,N_4535,N_4760);
nand U5045 (N_5045,N_4601,N_4673);
and U5046 (N_5046,N_4573,N_4423);
or U5047 (N_5047,N_4407,N_4795);
or U5048 (N_5048,N_4573,N_4697);
nor U5049 (N_5049,N_4681,N_4466);
nand U5050 (N_5050,N_4471,N_4617);
nand U5051 (N_5051,N_4599,N_4567);
nand U5052 (N_5052,N_4759,N_4418);
nor U5053 (N_5053,N_4642,N_4518);
and U5054 (N_5054,N_4532,N_4622);
or U5055 (N_5055,N_4431,N_4606);
or U5056 (N_5056,N_4507,N_4493);
nor U5057 (N_5057,N_4626,N_4492);
or U5058 (N_5058,N_4625,N_4411);
nor U5059 (N_5059,N_4440,N_4762);
and U5060 (N_5060,N_4577,N_4437);
and U5061 (N_5061,N_4614,N_4695);
nor U5062 (N_5062,N_4477,N_4445);
or U5063 (N_5063,N_4792,N_4452);
nand U5064 (N_5064,N_4495,N_4423);
and U5065 (N_5065,N_4672,N_4438);
nor U5066 (N_5066,N_4601,N_4670);
or U5067 (N_5067,N_4531,N_4708);
nand U5068 (N_5068,N_4452,N_4492);
nand U5069 (N_5069,N_4588,N_4793);
and U5070 (N_5070,N_4593,N_4558);
and U5071 (N_5071,N_4551,N_4775);
and U5072 (N_5072,N_4471,N_4489);
and U5073 (N_5073,N_4714,N_4701);
nor U5074 (N_5074,N_4578,N_4759);
and U5075 (N_5075,N_4471,N_4559);
nor U5076 (N_5076,N_4685,N_4776);
nor U5077 (N_5077,N_4626,N_4792);
nor U5078 (N_5078,N_4477,N_4565);
nand U5079 (N_5079,N_4530,N_4612);
nor U5080 (N_5080,N_4546,N_4522);
nor U5081 (N_5081,N_4476,N_4730);
xor U5082 (N_5082,N_4406,N_4566);
or U5083 (N_5083,N_4484,N_4617);
nor U5084 (N_5084,N_4620,N_4429);
nand U5085 (N_5085,N_4521,N_4557);
nor U5086 (N_5086,N_4765,N_4556);
and U5087 (N_5087,N_4550,N_4597);
nand U5088 (N_5088,N_4413,N_4575);
nor U5089 (N_5089,N_4797,N_4634);
nand U5090 (N_5090,N_4459,N_4500);
nand U5091 (N_5091,N_4619,N_4624);
and U5092 (N_5092,N_4586,N_4496);
nand U5093 (N_5093,N_4706,N_4580);
nand U5094 (N_5094,N_4746,N_4734);
or U5095 (N_5095,N_4573,N_4464);
nor U5096 (N_5096,N_4492,N_4412);
or U5097 (N_5097,N_4578,N_4691);
and U5098 (N_5098,N_4585,N_4579);
nand U5099 (N_5099,N_4740,N_4520);
and U5100 (N_5100,N_4511,N_4573);
and U5101 (N_5101,N_4797,N_4407);
nor U5102 (N_5102,N_4747,N_4404);
nor U5103 (N_5103,N_4728,N_4494);
nand U5104 (N_5104,N_4643,N_4459);
or U5105 (N_5105,N_4612,N_4558);
nand U5106 (N_5106,N_4461,N_4462);
nand U5107 (N_5107,N_4743,N_4568);
and U5108 (N_5108,N_4519,N_4488);
nand U5109 (N_5109,N_4535,N_4528);
and U5110 (N_5110,N_4657,N_4687);
nor U5111 (N_5111,N_4442,N_4645);
nand U5112 (N_5112,N_4777,N_4647);
or U5113 (N_5113,N_4749,N_4426);
nor U5114 (N_5114,N_4680,N_4580);
nand U5115 (N_5115,N_4553,N_4488);
nor U5116 (N_5116,N_4521,N_4593);
and U5117 (N_5117,N_4665,N_4638);
nor U5118 (N_5118,N_4461,N_4515);
or U5119 (N_5119,N_4761,N_4425);
or U5120 (N_5120,N_4547,N_4773);
nor U5121 (N_5121,N_4548,N_4721);
nor U5122 (N_5122,N_4754,N_4413);
nor U5123 (N_5123,N_4619,N_4777);
nor U5124 (N_5124,N_4526,N_4723);
or U5125 (N_5125,N_4524,N_4505);
or U5126 (N_5126,N_4782,N_4487);
or U5127 (N_5127,N_4594,N_4445);
or U5128 (N_5128,N_4441,N_4423);
and U5129 (N_5129,N_4720,N_4702);
or U5130 (N_5130,N_4509,N_4495);
and U5131 (N_5131,N_4581,N_4569);
and U5132 (N_5132,N_4644,N_4563);
and U5133 (N_5133,N_4441,N_4655);
or U5134 (N_5134,N_4704,N_4423);
or U5135 (N_5135,N_4459,N_4542);
nor U5136 (N_5136,N_4730,N_4798);
nor U5137 (N_5137,N_4512,N_4725);
and U5138 (N_5138,N_4589,N_4688);
nand U5139 (N_5139,N_4491,N_4639);
or U5140 (N_5140,N_4401,N_4426);
nor U5141 (N_5141,N_4702,N_4647);
and U5142 (N_5142,N_4695,N_4512);
nor U5143 (N_5143,N_4711,N_4486);
or U5144 (N_5144,N_4749,N_4628);
or U5145 (N_5145,N_4588,N_4688);
nand U5146 (N_5146,N_4745,N_4674);
and U5147 (N_5147,N_4592,N_4780);
nor U5148 (N_5148,N_4473,N_4593);
or U5149 (N_5149,N_4507,N_4564);
nor U5150 (N_5150,N_4458,N_4749);
nand U5151 (N_5151,N_4428,N_4402);
and U5152 (N_5152,N_4729,N_4505);
or U5153 (N_5153,N_4497,N_4619);
nor U5154 (N_5154,N_4484,N_4608);
or U5155 (N_5155,N_4690,N_4762);
and U5156 (N_5156,N_4616,N_4663);
nand U5157 (N_5157,N_4443,N_4668);
and U5158 (N_5158,N_4500,N_4416);
and U5159 (N_5159,N_4794,N_4726);
xor U5160 (N_5160,N_4530,N_4771);
or U5161 (N_5161,N_4486,N_4739);
or U5162 (N_5162,N_4481,N_4560);
nand U5163 (N_5163,N_4631,N_4402);
and U5164 (N_5164,N_4682,N_4514);
nand U5165 (N_5165,N_4497,N_4600);
and U5166 (N_5166,N_4675,N_4568);
and U5167 (N_5167,N_4681,N_4667);
or U5168 (N_5168,N_4671,N_4669);
or U5169 (N_5169,N_4416,N_4664);
nor U5170 (N_5170,N_4449,N_4418);
nor U5171 (N_5171,N_4732,N_4628);
or U5172 (N_5172,N_4419,N_4771);
nor U5173 (N_5173,N_4458,N_4451);
and U5174 (N_5174,N_4545,N_4623);
nand U5175 (N_5175,N_4561,N_4727);
xnor U5176 (N_5176,N_4428,N_4724);
and U5177 (N_5177,N_4592,N_4761);
nand U5178 (N_5178,N_4629,N_4545);
or U5179 (N_5179,N_4547,N_4595);
and U5180 (N_5180,N_4797,N_4425);
and U5181 (N_5181,N_4498,N_4708);
and U5182 (N_5182,N_4614,N_4628);
or U5183 (N_5183,N_4615,N_4465);
or U5184 (N_5184,N_4443,N_4440);
nor U5185 (N_5185,N_4723,N_4598);
or U5186 (N_5186,N_4592,N_4583);
and U5187 (N_5187,N_4648,N_4411);
nand U5188 (N_5188,N_4450,N_4684);
and U5189 (N_5189,N_4490,N_4715);
or U5190 (N_5190,N_4441,N_4749);
and U5191 (N_5191,N_4544,N_4717);
nand U5192 (N_5192,N_4740,N_4518);
nor U5193 (N_5193,N_4661,N_4686);
nand U5194 (N_5194,N_4665,N_4754);
nand U5195 (N_5195,N_4740,N_4407);
nand U5196 (N_5196,N_4496,N_4714);
nor U5197 (N_5197,N_4511,N_4663);
and U5198 (N_5198,N_4460,N_4570);
and U5199 (N_5199,N_4457,N_4530);
nor U5200 (N_5200,N_4898,N_4916);
and U5201 (N_5201,N_4997,N_4897);
nand U5202 (N_5202,N_5050,N_5015);
and U5203 (N_5203,N_4991,N_5170);
or U5204 (N_5204,N_4944,N_4955);
nand U5205 (N_5205,N_5160,N_4988);
nand U5206 (N_5206,N_5081,N_5136);
or U5207 (N_5207,N_5158,N_4970);
nor U5208 (N_5208,N_4879,N_5053);
nor U5209 (N_5209,N_4844,N_4823);
or U5210 (N_5210,N_5022,N_4873);
nor U5211 (N_5211,N_4836,N_4815);
nand U5212 (N_5212,N_4971,N_4866);
nor U5213 (N_5213,N_5094,N_4811);
or U5214 (N_5214,N_4943,N_5182);
and U5215 (N_5215,N_4804,N_5043);
and U5216 (N_5216,N_5028,N_5061);
and U5217 (N_5217,N_4978,N_5163);
nor U5218 (N_5218,N_5169,N_4874);
or U5219 (N_5219,N_4965,N_5176);
nand U5220 (N_5220,N_5185,N_5102);
nand U5221 (N_5221,N_4888,N_4882);
and U5222 (N_5222,N_4968,N_4973);
and U5223 (N_5223,N_4856,N_5197);
nor U5224 (N_5224,N_5054,N_4993);
nor U5225 (N_5225,N_5069,N_5035);
nand U5226 (N_5226,N_5171,N_4829);
and U5227 (N_5227,N_5067,N_4816);
nor U5228 (N_5228,N_4999,N_4869);
nand U5229 (N_5229,N_5079,N_4826);
and U5230 (N_5230,N_4863,N_4837);
and U5231 (N_5231,N_4875,N_5036);
nand U5232 (N_5232,N_4867,N_4979);
and U5233 (N_5233,N_4919,N_4987);
nand U5234 (N_5234,N_4995,N_4957);
and U5235 (N_5235,N_5082,N_4903);
nand U5236 (N_5236,N_4982,N_4905);
or U5237 (N_5237,N_5075,N_4959);
nand U5238 (N_5238,N_5190,N_4914);
nand U5239 (N_5239,N_5140,N_5117);
nor U5240 (N_5240,N_5047,N_4901);
and U5241 (N_5241,N_4977,N_4877);
nor U5242 (N_5242,N_5121,N_5162);
nand U5243 (N_5243,N_4893,N_4820);
nand U5244 (N_5244,N_4807,N_5196);
nand U5245 (N_5245,N_5107,N_4937);
or U5246 (N_5246,N_4813,N_5045);
and U5247 (N_5247,N_5099,N_5145);
nor U5248 (N_5248,N_4899,N_4885);
nand U5249 (N_5249,N_4953,N_4950);
nor U5250 (N_5250,N_4803,N_4932);
and U5251 (N_5251,N_5151,N_5023);
or U5252 (N_5252,N_4825,N_5006);
nor U5253 (N_5253,N_4906,N_4894);
or U5254 (N_5254,N_4946,N_4969);
and U5255 (N_5255,N_5156,N_5146);
or U5256 (N_5256,N_5115,N_5177);
nor U5257 (N_5257,N_5126,N_4831);
nand U5258 (N_5258,N_5192,N_5180);
nor U5259 (N_5259,N_4835,N_4850);
and U5260 (N_5260,N_4994,N_5071);
and U5261 (N_5261,N_5051,N_5063);
nor U5262 (N_5262,N_5175,N_5065);
or U5263 (N_5263,N_5038,N_5168);
or U5264 (N_5264,N_4832,N_5000);
nand U5265 (N_5265,N_5132,N_5157);
nor U5266 (N_5266,N_4886,N_5076);
or U5267 (N_5267,N_5110,N_5090);
nand U5268 (N_5268,N_5116,N_4819);
nor U5269 (N_5269,N_4839,N_5141);
nand U5270 (N_5270,N_5129,N_4954);
nand U5271 (N_5271,N_5007,N_4830);
and U5272 (N_5272,N_4814,N_4920);
and U5273 (N_5273,N_4864,N_4849);
or U5274 (N_5274,N_4872,N_5031);
or U5275 (N_5275,N_5037,N_5167);
and U5276 (N_5276,N_4917,N_5093);
or U5277 (N_5277,N_5096,N_4868);
nand U5278 (N_5278,N_4834,N_5166);
nand U5279 (N_5279,N_4876,N_4865);
nand U5280 (N_5280,N_4890,N_5186);
nor U5281 (N_5281,N_4860,N_4808);
nand U5282 (N_5282,N_5021,N_5144);
and U5283 (N_5283,N_5080,N_4871);
nand U5284 (N_5284,N_4900,N_4847);
or U5285 (N_5285,N_4922,N_4948);
nand U5286 (N_5286,N_5155,N_5147);
nor U5287 (N_5287,N_5143,N_5084);
or U5288 (N_5288,N_5120,N_4881);
xor U5289 (N_5289,N_4908,N_4904);
nor U5290 (N_5290,N_4818,N_4800);
or U5291 (N_5291,N_4909,N_5009);
and U5292 (N_5292,N_4845,N_4984);
nand U5293 (N_5293,N_4891,N_5173);
nand U5294 (N_5294,N_4851,N_5193);
nor U5295 (N_5295,N_4801,N_5026);
nand U5296 (N_5296,N_4930,N_5113);
or U5297 (N_5297,N_5077,N_4921);
and U5298 (N_5298,N_4805,N_4840);
or U5299 (N_5299,N_5034,N_4859);
or U5300 (N_5300,N_4989,N_5033);
nor U5301 (N_5301,N_5001,N_5060);
nand U5302 (N_5302,N_4974,N_4887);
nand U5303 (N_5303,N_4967,N_5064);
nand U5304 (N_5304,N_5072,N_4963);
and U5305 (N_5305,N_4843,N_4951);
or U5306 (N_5306,N_5152,N_5052);
nor U5307 (N_5307,N_5040,N_5103);
and U5308 (N_5308,N_4940,N_4927);
nor U5309 (N_5309,N_4822,N_4956);
or U5310 (N_5310,N_5044,N_4812);
or U5311 (N_5311,N_4929,N_5085);
or U5312 (N_5312,N_4964,N_5105);
and U5313 (N_5313,N_5165,N_5059);
nand U5314 (N_5314,N_4941,N_5008);
nor U5315 (N_5315,N_4936,N_5057);
nand U5316 (N_5316,N_5199,N_5097);
and U5317 (N_5317,N_5139,N_4966);
nand U5318 (N_5318,N_4870,N_5055);
nand U5319 (N_5319,N_5024,N_5003);
nor U5320 (N_5320,N_4842,N_4896);
nor U5321 (N_5321,N_5066,N_4880);
and U5322 (N_5322,N_5112,N_4923);
nand U5323 (N_5323,N_4809,N_4821);
nand U5324 (N_5324,N_5154,N_4857);
nand U5325 (N_5325,N_5106,N_4972);
xnor U5326 (N_5326,N_4910,N_5164);
nor U5327 (N_5327,N_4878,N_5127);
nor U5328 (N_5328,N_4961,N_5013);
and U5329 (N_5329,N_5184,N_5130);
nor U5330 (N_5330,N_5118,N_4895);
nand U5331 (N_5331,N_5138,N_5017);
nor U5332 (N_5332,N_5042,N_5133);
nor U5333 (N_5333,N_5068,N_4817);
nor U5334 (N_5334,N_5111,N_5091);
or U5335 (N_5335,N_4931,N_5131);
nor U5336 (N_5336,N_5029,N_5083);
and U5337 (N_5337,N_4949,N_4996);
or U5338 (N_5338,N_4985,N_5124);
and U5339 (N_5339,N_5187,N_4855);
and U5340 (N_5340,N_5191,N_4976);
or U5341 (N_5341,N_5010,N_4848);
nor U5342 (N_5342,N_4861,N_5020);
and U5343 (N_5343,N_4924,N_4810);
nor U5344 (N_5344,N_5161,N_4913);
nor U5345 (N_5345,N_5195,N_5062);
and U5346 (N_5346,N_4939,N_4938);
nand U5347 (N_5347,N_4992,N_5027);
or U5348 (N_5348,N_5188,N_4841);
or U5349 (N_5349,N_4962,N_5086);
and U5350 (N_5350,N_5014,N_5189);
and U5351 (N_5351,N_4942,N_5032);
nor U5352 (N_5352,N_5012,N_5074);
nor U5353 (N_5353,N_5088,N_4926);
or U5354 (N_5354,N_5135,N_5178);
or U5355 (N_5355,N_4852,N_4915);
or U5356 (N_5356,N_4986,N_5016);
nor U5357 (N_5357,N_5058,N_4892);
or U5358 (N_5358,N_5181,N_4907);
and U5359 (N_5359,N_4958,N_5049);
nor U5360 (N_5360,N_5114,N_5056);
nand U5361 (N_5361,N_5122,N_5070);
nand U5362 (N_5362,N_5041,N_5179);
and U5363 (N_5363,N_4854,N_5198);
or U5364 (N_5364,N_5101,N_5039);
or U5365 (N_5365,N_5078,N_4824);
nand U5366 (N_5366,N_4918,N_5087);
and U5367 (N_5367,N_4806,N_5046);
or U5368 (N_5368,N_5011,N_4975);
nor U5369 (N_5369,N_4858,N_5092);
or U5370 (N_5370,N_5183,N_5128);
or U5371 (N_5371,N_4853,N_5108);
and U5372 (N_5372,N_4838,N_5150);
nor U5373 (N_5373,N_4980,N_4990);
nor U5374 (N_5374,N_5089,N_5153);
or U5375 (N_5375,N_4884,N_4934);
or U5376 (N_5376,N_5172,N_5104);
and U5377 (N_5377,N_4935,N_5119);
and U5378 (N_5378,N_5174,N_4952);
nor U5379 (N_5379,N_4827,N_5149);
or U5380 (N_5380,N_5098,N_4902);
or U5381 (N_5381,N_5048,N_5137);
or U5382 (N_5382,N_5019,N_4889);
and U5383 (N_5383,N_4802,N_5005);
or U5384 (N_5384,N_4912,N_5148);
nor U5385 (N_5385,N_5004,N_4933);
nor U5386 (N_5386,N_5030,N_4883);
nand U5387 (N_5387,N_5142,N_4862);
or U5388 (N_5388,N_5002,N_5194);
and U5389 (N_5389,N_4828,N_4960);
or U5390 (N_5390,N_4911,N_5134);
nand U5391 (N_5391,N_4928,N_4983);
nor U5392 (N_5392,N_4925,N_4945);
nand U5393 (N_5393,N_5018,N_5100);
nor U5394 (N_5394,N_5109,N_4846);
nand U5395 (N_5395,N_4998,N_5123);
nand U5396 (N_5396,N_5025,N_5073);
or U5397 (N_5397,N_5095,N_4833);
nor U5398 (N_5398,N_4981,N_4947);
and U5399 (N_5399,N_5125,N_5159);
nor U5400 (N_5400,N_4847,N_5154);
nand U5401 (N_5401,N_5175,N_5057);
or U5402 (N_5402,N_4832,N_4938);
and U5403 (N_5403,N_5159,N_5149);
nor U5404 (N_5404,N_5134,N_5057);
xnor U5405 (N_5405,N_4828,N_4888);
nand U5406 (N_5406,N_5180,N_5030);
nor U5407 (N_5407,N_4967,N_5076);
or U5408 (N_5408,N_4919,N_4857);
nand U5409 (N_5409,N_4946,N_4875);
xnor U5410 (N_5410,N_5045,N_4947);
nor U5411 (N_5411,N_4911,N_4839);
nor U5412 (N_5412,N_5078,N_5096);
nor U5413 (N_5413,N_4996,N_5198);
or U5414 (N_5414,N_5138,N_5061);
or U5415 (N_5415,N_5117,N_5000);
nor U5416 (N_5416,N_5104,N_5129);
or U5417 (N_5417,N_5093,N_5137);
nor U5418 (N_5418,N_4921,N_4867);
nor U5419 (N_5419,N_5097,N_4828);
and U5420 (N_5420,N_5033,N_4822);
nor U5421 (N_5421,N_5004,N_4805);
nor U5422 (N_5422,N_5111,N_4874);
or U5423 (N_5423,N_4904,N_4815);
or U5424 (N_5424,N_5197,N_5023);
nor U5425 (N_5425,N_5085,N_5046);
or U5426 (N_5426,N_4833,N_5150);
and U5427 (N_5427,N_5011,N_5012);
nand U5428 (N_5428,N_5100,N_5176);
or U5429 (N_5429,N_5134,N_5060);
nand U5430 (N_5430,N_4986,N_4953);
and U5431 (N_5431,N_4853,N_5044);
or U5432 (N_5432,N_5094,N_5120);
and U5433 (N_5433,N_5122,N_4911);
nor U5434 (N_5434,N_5154,N_5001);
nor U5435 (N_5435,N_4965,N_4911);
and U5436 (N_5436,N_5032,N_4825);
and U5437 (N_5437,N_4832,N_4807);
nor U5438 (N_5438,N_4914,N_4995);
and U5439 (N_5439,N_5123,N_4847);
or U5440 (N_5440,N_4873,N_4932);
nor U5441 (N_5441,N_4818,N_4991);
nor U5442 (N_5442,N_5047,N_5079);
and U5443 (N_5443,N_4891,N_5062);
nor U5444 (N_5444,N_4840,N_5022);
nor U5445 (N_5445,N_4904,N_5030);
xnor U5446 (N_5446,N_4934,N_5031);
nand U5447 (N_5447,N_5005,N_5126);
or U5448 (N_5448,N_5088,N_5083);
nand U5449 (N_5449,N_4984,N_5087);
and U5450 (N_5450,N_4906,N_5171);
or U5451 (N_5451,N_5051,N_5148);
nor U5452 (N_5452,N_5162,N_5032);
nor U5453 (N_5453,N_5085,N_5148);
and U5454 (N_5454,N_5139,N_4906);
nand U5455 (N_5455,N_5121,N_5083);
nor U5456 (N_5456,N_4916,N_4819);
xnor U5457 (N_5457,N_4921,N_4856);
or U5458 (N_5458,N_5012,N_4860);
nand U5459 (N_5459,N_5100,N_5029);
or U5460 (N_5460,N_5113,N_5199);
nor U5461 (N_5461,N_5164,N_5036);
nor U5462 (N_5462,N_4964,N_5096);
and U5463 (N_5463,N_4970,N_4949);
nand U5464 (N_5464,N_4902,N_4884);
nor U5465 (N_5465,N_4913,N_5040);
or U5466 (N_5466,N_4977,N_5196);
nor U5467 (N_5467,N_4892,N_5094);
nand U5468 (N_5468,N_4950,N_5194);
and U5469 (N_5469,N_5037,N_4824);
and U5470 (N_5470,N_5094,N_5119);
and U5471 (N_5471,N_5060,N_5077);
or U5472 (N_5472,N_5171,N_5152);
nand U5473 (N_5473,N_5004,N_4842);
or U5474 (N_5474,N_4934,N_4894);
and U5475 (N_5475,N_5193,N_5095);
or U5476 (N_5476,N_4951,N_4898);
nor U5477 (N_5477,N_5017,N_5021);
or U5478 (N_5478,N_4930,N_4974);
nor U5479 (N_5479,N_5109,N_5099);
and U5480 (N_5480,N_5092,N_4851);
or U5481 (N_5481,N_4931,N_4806);
and U5482 (N_5482,N_4920,N_5105);
and U5483 (N_5483,N_5028,N_4859);
nor U5484 (N_5484,N_5066,N_5149);
and U5485 (N_5485,N_4967,N_5126);
nand U5486 (N_5486,N_4820,N_4941);
nand U5487 (N_5487,N_5132,N_5078);
nand U5488 (N_5488,N_4969,N_5144);
or U5489 (N_5489,N_4970,N_4906);
or U5490 (N_5490,N_5191,N_5044);
and U5491 (N_5491,N_5184,N_5028);
nand U5492 (N_5492,N_5008,N_5169);
and U5493 (N_5493,N_4941,N_4952);
nor U5494 (N_5494,N_5138,N_4814);
and U5495 (N_5495,N_4821,N_4832);
or U5496 (N_5496,N_4992,N_4875);
nand U5497 (N_5497,N_5035,N_4929);
nand U5498 (N_5498,N_5014,N_4869);
nor U5499 (N_5499,N_5162,N_4873);
or U5500 (N_5500,N_5057,N_5093);
nand U5501 (N_5501,N_5087,N_5049);
nand U5502 (N_5502,N_4899,N_5199);
and U5503 (N_5503,N_5106,N_5152);
nand U5504 (N_5504,N_4800,N_4817);
or U5505 (N_5505,N_4938,N_4906);
nand U5506 (N_5506,N_5195,N_5087);
and U5507 (N_5507,N_5113,N_5030);
or U5508 (N_5508,N_5047,N_5198);
and U5509 (N_5509,N_4920,N_4892);
nand U5510 (N_5510,N_5064,N_4881);
and U5511 (N_5511,N_5064,N_4988);
and U5512 (N_5512,N_5161,N_5149);
or U5513 (N_5513,N_5102,N_5019);
nor U5514 (N_5514,N_4922,N_5062);
and U5515 (N_5515,N_5068,N_5050);
nand U5516 (N_5516,N_4841,N_5050);
nor U5517 (N_5517,N_4916,N_4841);
nor U5518 (N_5518,N_4880,N_4922);
and U5519 (N_5519,N_4852,N_4969);
nor U5520 (N_5520,N_5153,N_4922);
or U5521 (N_5521,N_4984,N_4885);
and U5522 (N_5522,N_5031,N_4820);
nand U5523 (N_5523,N_4904,N_5077);
or U5524 (N_5524,N_4878,N_4929);
nor U5525 (N_5525,N_4927,N_5048);
nor U5526 (N_5526,N_5089,N_4970);
nor U5527 (N_5527,N_4819,N_5112);
nor U5528 (N_5528,N_5129,N_5037);
and U5529 (N_5529,N_4900,N_5023);
or U5530 (N_5530,N_4818,N_5036);
nor U5531 (N_5531,N_4888,N_5047);
or U5532 (N_5532,N_5191,N_5045);
and U5533 (N_5533,N_4815,N_4898);
or U5534 (N_5534,N_5160,N_4940);
or U5535 (N_5535,N_5057,N_4924);
nand U5536 (N_5536,N_4834,N_4999);
and U5537 (N_5537,N_5043,N_5097);
and U5538 (N_5538,N_4828,N_5091);
or U5539 (N_5539,N_5168,N_5147);
nand U5540 (N_5540,N_5197,N_4820);
and U5541 (N_5541,N_5043,N_4890);
and U5542 (N_5542,N_4993,N_5027);
nand U5543 (N_5543,N_4990,N_4817);
or U5544 (N_5544,N_5161,N_4831);
nand U5545 (N_5545,N_5125,N_5131);
nor U5546 (N_5546,N_4941,N_5171);
or U5547 (N_5547,N_5068,N_4935);
and U5548 (N_5548,N_4819,N_4885);
or U5549 (N_5549,N_5071,N_4981);
and U5550 (N_5550,N_5196,N_5063);
nand U5551 (N_5551,N_4888,N_4863);
nor U5552 (N_5552,N_4999,N_5169);
or U5553 (N_5553,N_5025,N_4982);
or U5554 (N_5554,N_4896,N_5055);
and U5555 (N_5555,N_4821,N_5039);
nand U5556 (N_5556,N_5078,N_5051);
and U5557 (N_5557,N_4886,N_5018);
nand U5558 (N_5558,N_5163,N_5126);
nand U5559 (N_5559,N_5082,N_5015);
nand U5560 (N_5560,N_5043,N_5109);
nor U5561 (N_5561,N_5166,N_5113);
nand U5562 (N_5562,N_5024,N_4828);
or U5563 (N_5563,N_4989,N_4903);
or U5564 (N_5564,N_4961,N_4910);
nor U5565 (N_5565,N_4826,N_4854);
nor U5566 (N_5566,N_5035,N_5056);
nor U5567 (N_5567,N_4898,N_4803);
nand U5568 (N_5568,N_4849,N_4891);
and U5569 (N_5569,N_4889,N_5080);
and U5570 (N_5570,N_5015,N_4823);
and U5571 (N_5571,N_5165,N_5083);
nor U5572 (N_5572,N_5050,N_4875);
or U5573 (N_5573,N_5102,N_4933);
nor U5574 (N_5574,N_5159,N_4933);
and U5575 (N_5575,N_4816,N_4842);
or U5576 (N_5576,N_5038,N_5147);
nor U5577 (N_5577,N_4964,N_4872);
nor U5578 (N_5578,N_5147,N_5000);
nand U5579 (N_5579,N_5072,N_4922);
nor U5580 (N_5580,N_5110,N_5174);
or U5581 (N_5581,N_5108,N_5051);
or U5582 (N_5582,N_4998,N_5085);
and U5583 (N_5583,N_4976,N_5080);
nand U5584 (N_5584,N_4996,N_5117);
or U5585 (N_5585,N_4855,N_4982);
nand U5586 (N_5586,N_5117,N_5142);
nor U5587 (N_5587,N_5162,N_5073);
and U5588 (N_5588,N_5064,N_5096);
nand U5589 (N_5589,N_4835,N_5042);
nor U5590 (N_5590,N_4817,N_4948);
nand U5591 (N_5591,N_5189,N_4833);
nand U5592 (N_5592,N_4921,N_5071);
or U5593 (N_5593,N_5179,N_4867);
and U5594 (N_5594,N_4965,N_4889);
nor U5595 (N_5595,N_5193,N_5133);
nand U5596 (N_5596,N_5192,N_5141);
nor U5597 (N_5597,N_4967,N_5089);
and U5598 (N_5598,N_5015,N_5094);
nor U5599 (N_5599,N_4873,N_5038);
or U5600 (N_5600,N_5267,N_5405);
or U5601 (N_5601,N_5575,N_5293);
nand U5602 (N_5602,N_5412,N_5542);
or U5603 (N_5603,N_5493,N_5561);
or U5604 (N_5604,N_5282,N_5509);
nand U5605 (N_5605,N_5582,N_5315);
or U5606 (N_5606,N_5284,N_5215);
nand U5607 (N_5607,N_5480,N_5216);
and U5608 (N_5608,N_5342,N_5511);
or U5609 (N_5609,N_5323,N_5523);
nor U5610 (N_5610,N_5201,N_5428);
nand U5611 (N_5611,N_5253,N_5246);
nand U5612 (N_5612,N_5371,N_5564);
or U5613 (N_5613,N_5461,N_5551);
nor U5614 (N_5614,N_5592,N_5465);
or U5615 (N_5615,N_5485,N_5273);
or U5616 (N_5616,N_5257,N_5500);
and U5617 (N_5617,N_5319,N_5567);
nor U5618 (N_5618,N_5346,N_5470);
nor U5619 (N_5619,N_5502,N_5382);
nand U5620 (N_5620,N_5334,N_5489);
nor U5621 (N_5621,N_5361,N_5539);
and U5622 (N_5622,N_5492,N_5488);
or U5623 (N_5623,N_5331,N_5579);
nand U5624 (N_5624,N_5270,N_5358);
or U5625 (N_5625,N_5439,N_5325);
or U5626 (N_5626,N_5530,N_5240);
and U5627 (N_5627,N_5395,N_5288);
or U5628 (N_5628,N_5340,N_5208);
nor U5629 (N_5629,N_5341,N_5256);
or U5630 (N_5630,N_5343,N_5455);
nor U5631 (N_5631,N_5406,N_5312);
or U5632 (N_5632,N_5454,N_5360);
and U5633 (N_5633,N_5233,N_5307);
or U5634 (N_5634,N_5247,N_5200);
or U5635 (N_5635,N_5392,N_5271);
or U5636 (N_5636,N_5469,N_5234);
or U5637 (N_5637,N_5593,N_5232);
nor U5638 (N_5638,N_5269,N_5448);
and U5639 (N_5639,N_5495,N_5329);
and U5640 (N_5640,N_5432,N_5259);
and U5641 (N_5641,N_5436,N_5518);
or U5642 (N_5642,N_5421,N_5403);
or U5643 (N_5643,N_5338,N_5496);
or U5644 (N_5644,N_5396,N_5276);
and U5645 (N_5645,N_5344,N_5423);
and U5646 (N_5646,N_5444,N_5241);
or U5647 (N_5647,N_5598,N_5353);
or U5648 (N_5648,N_5373,N_5433);
nand U5649 (N_5649,N_5224,N_5352);
and U5650 (N_5650,N_5497,N_5554);
nor U5651 (N_5651,N_5532,N_5377);
and U5652 (N_5652,N_5220,N_5417);
and U5653 (N_5653,N_5393,N_5278);
or U5654 (N_5654,N_5449,N_5498);
or U5655 (N_5655,N_5437,N_5547);
nor U5656 (N_5656,N_5491,N_5481);
nand U5657 (N_5657,N_5265,N_5588);
or U5658 (N_5658,N_5571,N_5223);
nor U5659 (N_5659,N_5387,N_5538);
and U5660 (N_5660,N_5418,N_5431);
and U5661 (N_5661,N_5205,N_5471);
nand U5662 (N_5662,N_5553,N_5583);
nand U5663 (N_5663,N_5524,N_5504);
or U5664 (N_5664,N_5472,N_5484);
nor U5665 (N_5665,N_5379,N_5348);
nor U5666 (N_5666,N_5306,N_5308);
nor U5667 (N_5667,N_5225,N_5209);
and U5668 (N_5668,N_5441,N_5467);
nand U5669 (N_5669,N_5254,N_5398);
nor U5670 (N_5670,N_5295,N_5384);
or U5671 (N_5671,N_5355,N_5536);
and U5672 (N_5672,N_5228,N_5580);
and U5673 (N_5673,N_5457,N_5578);
nand U5674 (N_5674,N_5451,N_5559);
and U5675 (N_5675,N_5272,N_5243);
or U5676 (N_5676,N_5490,N_5522);
nor U5677 (N_5677,N_5560,N_5237);
and U5678 (N_5678,N_5236,N_5450);
nor U5679 (N_5679,N_5242,N_5221);
nand U5680 (N_5680,N_5408,N_5506);
nand U5681 (N_5681,N_5277,N_5499);
and U5682 (N_5682,N_5266,N_5462);
nor U5683 (N_5683,N_5268,N_5519);
and U5684 (N_5684,N_5318,N_5501);
or U5685 (N_5685,N_5263,N_5245);
nand U5686 (N_5686,N_5517,N_5581);
nor U5687 (N_5687,N_5548,N_5314);
nor U5688 (N_5688,N_5456,N_5570);
or U5689 (N_5689,N_5594,N_5591);
nand U5690 (N_5690,N_5364,N_5248);
or U5691 (N_5691,N_5414,N_5305);
nand U5692 (N_5692,N_5573,N_5375);
nand U5693 (N_5693,N_5213,N_5328);
nand U5694 (N_5694,N_5238,N_5541);
and U5695 (N_5695,N_5376,N_5332);
and U5696 (N_5696,N_5239,N_5244);
or U5697 (N_5697,N_5370,N_5291);
nor U5698 (N_5698,N_5320,N_5516);
and U5699 (N_5699,N_5285,N_5218);
and U5700 (N_5700,N_5584,N_5557);
and U5701 (N_5701,N_5300,N_5311);
nor U5702 (N_5702,N_5357,N_5280);
nand U5703 (N_5703,N_5464,N_5363);
or U5704 (N_5704,N_5563,N_5350);
or U5705 (N_5705,N_5204,N_5415);
or U5706 (N_5706,N_5585,N_5458);
nor U5707 (N_5707,N_5321,N_5262);
or U5708 (N_5708,N_5521,N_5531);
nand U5709 (N_5709,N_5427,N_5482);
nand U5710 (N_5710,N_5258,N_5550);
or U5711 (N_5711,N_5302,N_5424);
nand U5712 (N_5712,N_5381,N_5235);
nand U5713 (N_5713,N_5211,N_5558);
or U5714 (N_5714,N_5203,N_5586);
nor U5715 (N_5715,N_5438,N_5394);
nor U5716 (N_5716,N_5401,N_5407);
or U5717 (N_5717,N_5478,N_5569);
nor U5718 (N_5718,N_5525,N_5316);
and U5719 (N_5719,N_5362,N_5335);
or U5720 (N_5720,N_5459,N_5386);
and U5721 (N_5721,N_5359,N_5446);
nand U5722 (N_5722,N_5324,N_5250);
or U5723 (N_5723,N_5351,N_5426);
or U5724 (N_5724,N_5230,N_5599);
and U5725 (N_5725,N_5231,N_5336);
nor U5726 (N_5726,N_5366,N_5565);
and U5727 (N_5727,N_5445,N_5577);
nor U5728 (N_5728,N_5333,N_5313);
or U5729 (N_5729,N_5413,N_5283);
or U5730 (N_5730,N_5543,N_5447);
nand U5731 (N_5731,N_5349,N_5466);
or U5732 (N_5732,N_5510,N_5549);
nor U5733 (N_5733,N_5255,N_5390);
nand U5734 (N_5734,N_5369,N_5347);
nor U5735 (N_5735,N_5251,N_5528);
or U5736 (N_5736,N_5527,N_5222);
nand U5737 (N_5737,N_5327,N_5298);
nor U5738 (N_5738,N_5430,N_5494);
nand U5739 (N_5739,N_5322,N_5317);
nand U5740 (N_5740,N_5529,N_5420);
nand U5741 (N_5741,N_5526,N_5287);
and U5742 (N_5742,N_5388,N_5562);
and U5743 (N_5743,N_5574,N_5545);
nand U5744 (N_5744,N_5309,N_5546);
and U5745 (N_5745,N_5597,N_5540);
nor U5746 (N_5746,N_5217,N_5207);
and U5747 (N_5747,N_5249,N_5576);
or U5748 (N_5748,N_5210,N_5389);
and U5749 (N_5749,N_5261,N_5568);
nor U5750 (N_5750,N_5368,N_5544);
or U5751 (N_5751,N_5483,N_5294);
or U5752 (N_5752,N_5212,N_5587);
nor U5753 (N_5753,N_5345,N_5595);
nor U5754 (N_5754,N_5290,N_5537);
and U5755 (N_5755,N_5589,N_5229);
nor U5756 (N_5756,N_5372,N_5555);
or U5757 (N_5757,N_5463,N_5385);
nand U5758 (N_5758,N_5508,N_5292);
or U5759 (N_5759,N_5503,N_5274);
nand U5760 (N_5760,N_5411,N_5400);
and U5761 (N_5761,N_5505,N_5468);
and U5762 (N_5762,N_5297,N_5513);
and U5763 (N_5763,N_5378,N_5416);
or U5764 (N_5764,N_5202,N_5304);
nor U5765 (N_5765,N_5303,N_5520);
nor U5766 (N_5766,N_5442,N_5219);
and U5767 (N_5767,N_5419,N_5275);
or U5768 (N_5768,N_5227,N_5440);
and U5769 (N_5769,N_5367,N_5339);
and U5770 (N_5770,N_5264,N_5402);
nor U5771 (N_5771,N_5397,N_5410);
or U5772 (N_5772,N_5487,N_5281);
nor U5773 (N_5773,N_5535,N_5404);
or U5774 (N_5774,N_5429,N_5473);
xnor U5775 (N_5775,N_5391,N_5301);
nor U5776 (N_5776,N_5475,N_5572);
and U5777 (N_5777,N_5443,N_5310);
or U5778 (N_5778,N_5534,N_5434);
and U5779 (N_5779,N_5453,N_5289);
nor U5780 (N_5780,N_5337,N_5356);
nand U5781 (N_5781,N_5326,N_5460);
and U5782 (N_5782,N_5214,N_5512);
or U5783 (N_5783,N_5596,N_5330);
and U5784 (N_5784,N_5514,N_5590);
nor U5785 (N_5785,N_5452,N_5299);
or U5786 (N_5786,N_5279,N_5383);
or U5787 (N_5787,N_5479,N_5533);
or U5788 (N_5788,N_5425,N_5476);
nor U5789 (N_5789,N_5422,N_5552);
or U5790 (N_5790,N_5566,N_5354);
nand U5791 (N_5791,N_5286,N_5206);
or U5792 (N_5792,N_5260,N_5399);
nand U5793 (N_5793,N_5477,N_5409);
and U5794 (N_5794,N_5515,N_5486);
nor U5795 (N_5795,N_5374,N_5226);
nor U5796 (N_5796,N_5435,N_5296);
nor U5797 (N_5797,N_5474,N_5365);
and U5798 (N_5798,N_5507,N_5252);
nor U5799 (N_5799,N_5556,N_5380);
and U5800 (N_5800,N_5471,N_5567);
or U5801 (N_5801,N_5580,N_5265);
nor U5802 (N_5802,N_5351,N_5215);
or U5803 (N_5803,N_5512,N_5438);
nand U5804 (N_5804,N_5335,N_5519);
nand U5805 (N_5805,N_5241,N_5358);
and U5806 (N_5806,N_5421,N_5587);
or U5807 (N_5807,N_5317,N_5507);
nor U5808 (N_5808,N_5326,N_5264);
nor U5809 (N_5809,N_5205,N_5290);
and U5810 (N_5810,N_5454,N_5478);
or U5811 (N_5811,N_5272,N_5578);
and U5812 (N_5812,N_5430,N_5380);
nand U5813 (N_5813,N_5265,N_5271);
or U5814 (N_5814,N_5432,N_5542);
nand U5815 (N_5815,N_5313,N_5370);
nand U5816 (N_5816,N_5408,N_5248);
nor U5817 (N_5817,N_5495,N_5292);
nor U5818 (N_5818,N_5372,N_5595);
and U5819 (N_5819,N_5363,N_5515);
and U5820 (N_5820,N_5528,N_5208);
or U5821 (N_5821,N_5385,N_5258);
or U5822 (N_5822,N_5521,N_5339);
or U5823 (N_5823,N_5418,N_5348);
nor U5824 (N_5824,N_5589,N_5351);
nand U5825 (N_5825,N_5271,N_5461);
and U5826 (N_5826,N_5534,N_5395);
nand U5827 (N_5827,N_5354,N_5552);
nand U5828 (N_5828,N_5420,N_5225);
nand U5829 (N_5829,N_5452,N_5335);
and U5830 (N_5830,N_5278,N_5334);
nand U5831 (N_5831,N_5518,N_5303);
or U5832 (N_5832,N_5399,N_5381);
nor U5833 (N_5833,N_5407,N_5389);
or U5834 (N_5834,N_5488,N_5566);
and U5835 (N_5835,N_5335,N_5507);
and U5836 (N_5836,N_5543,N_5295);
nor U5837 (N_5837,N_5379,N_5558);
nand U5838 (N_5838,N_5249,N_5339);
nand U5839 (N_5839,N_5502,N_5460);
and U5840 (N_5840,N_5515,N_5572);
nand U5841 (N_5841,N_5224,N_5533);
or U5842 (N_5842,N_5544,N_5212);
nor U5843 (N_5843,N_5306,N_5572);
nor U5844 (N_5844,N_5519,N_5353);
nand U5845 (N_5845,N_5332,N_5404);
nand U5846 (N_5846,N_5341,N_5597);
nor U5847 (N_5847,N_5556,N_5450);
or U5848 (N_5848,N_5282,N_5344);
nor U5849 (N_5849,N_5340,N_5315);
or U5850 (N_5850,N_5469,N_5504);
nand U5851 (N_5851,N_5418,N_5500);
nor U5852 (N_5852,N_5370,N_5535);
nor U5853 (N_5853,N_5503,N_5359);
or U5854 (N_5854,N_5305,N_5533);
nor U5855 (N_5855,N_5491,N_5418);
or U5856 (N_5856,N_5466,N_5373);
nand U5857 (N_5857,N_5271,N_5558);
and U5858 (N_5858,N_5412,N_5414);
nor U5859 (N_5859,N_5466,N_5306);
nor U5860 (N_5860,N_5252,N_5473);
nand U5861 (N_5861,N_5340,N_5579);
nor U5862 (N_5862,N_5528,N_5265);
and U5863 (N_5863,N_5360,N_5228);
nor U5864 (N_5864,N_5475,N_5225);
or U5865 (N_5865,N_5364,N_5237);
and U5866 (N_5866,N_5206,N_5542);
nor U5867 (N_5867,N_5490,N_5400);
nor U5868 (N_5868,N_5218,N_5357);
or U5869 (N_5869,N_5574,N_5233);
nor U5870 (N_5870,N_5388,N_5401);
and U5871 (N_5871,N_5200,N_5569);
and U5872 (N_5872,N_5470,N_5390);
and U5873 (N_5873,N_5347,N_5335);
or U5874 (N_5874,N_5297,N_5546);
or U5875 (N_5875,N_5348,N_5259);
nor U5876 (N_5876,N_5280,N_5202);
nor U5877 (N_5877,N_5526,N_5470);
and U5878 (N_5878,N_5524,N_5459);
nand U5879 (N_5879,N_5487,N_5406);
or U5880 (N_5880,N_5480,N_5565);
nand U5881 (N_5881,N_5234,N_5244);
and U5882 (N_5882,N_5496,N_5363);
and U5883 (N_5883,N_5474,N_5443);
or U5884 (N_5884,N_5538,N_5367);
or U5885 (N_5885,N_5523,N_5320);
nand U5886 (N_5886,N_5327,N_5324);
nor U5887 (N_5887,N_5373,N_5267);
and U5888 (N_5888,N_5304,N_5221);
nor U5889 (N_5889,N_5291,N_5282);
nor U5890 (N_5890,N_5468,N_5375);
nand U5891 (N_5891,N_5348,N_5385);
nand U5892 (N_5892,N_5253,N_5385);
xnor U5893 (N_5893,N_5204,N_5324);
or U5894 (N_5894,N_5491,N_5490);
and U5895 (N_5895,N_5449,N_5551);
nand U5896 (N_5896,N_5271,N_5418);
nor U5897 (N_5897,N_5362,N_5269);
nand U5898 (N_5898,N_5266,N_5530);
xnor U5899 (N_5899,N_5221,N_5297);
and U5900 (N_5900,N_5489,N_5270);
nand U5901 (N_5901,N_5554,N_5283);
or U5902 (N_5902,N_5353,N_5537);
or U5903 (N_5903,N_5469,N_5431);
or U5904 (N_5904,N_5257,N_5585);
or U5905 (N_5905,N_5207,N_5558);
nand U5906 (N_5906,N_5304,N_5516);
or U5907 (N_5907,N_5398,N_5539);
nor U5908 (N_5908,N_5485,N_5260);
or U5909 (N_5909,N_5504,N_5270);
or U5910 (N_5910,N_5343,N_5344);
nor U5911 (N_5911,N_5516,N_5241);
nand U5912 (N_5912,N_5545,N_5287);
and U5913 (N_5913,N_5404,N_5223);
or U5914 (N_5914,N_5245,N_5541);
and U5915 (N_5915,N_5576,N_5492);
or U5916 (N_5916,N_5382,N_5460);
or U5917 (N_5917,N_5237,N_5216);
and U5918 (N_5918,N_5496,N_5536);
or U5919 (N_5919,N_5307,N_5354);
or U5920 (N_5920,N_5261,N_5492);
and U5921 (N_5921,N_5525,N_5479);
or U5922 (N_5922,N_5478,N_5272);
nand U5923 (N_5923,N_5273,N_5368);
and U5924 (N_5924,N_5489,N_5223);
nand U5925 (N_5925,N_5374,N_5497);
and U5926 (N_5926,N_5294,N_5471);
or U5927 (N_5927,N_5221,N_5400);
nor U5928 (N_5928,N_5333,N_5431);
nand U5929 (N_5929,N_5261,N_5249);
nand U5930 (N_5930,N_5240,N_5447);
and U5931 (N_5931,N_5401,N_5545);
or U5932 (N_5932,N_5556,N_5586);
and U5933 (N_5933,N_5231,N_5568);
nor U5934 (N_5934,N_5374,N_5359);
or U5935 (N_5935,N_5398,N_5212);
nand U5936 (N_5936,N_5538,N_5274);
or U5937 (N_5937,N_5329,N_5426);
nor U5938 (N_5938,N_5569,N_5587);
and U5939 (N_5939,N_5420,N_5344);
nand U5940 (N_5940,N_5264,N_5356);
nand U5941 (N_5941,N_5423,N_5337);
or U5942 (N_5942,N_5593,N_5390);
or U5943 (N_5943,N_5583,N_5438);
nand U5944 (N_5944,N_5272,N_5475);
nand U5945 (N_5945,N_5430,N_5598);
nor U5946 (N_5946,N_5227,N_5490);
or U5947 (N_5947,N_5299,N_5414);
nand U5948 (N_5948,N_5368,N_5337);
or U5949 (N_5949,N_5358,N_5554);
and U5950 (N_5950,N_5533,N_5341);
nand U5951 (N_5951,N_5598,N_5236);
nand U5952 (N_5952,N_5493,N_5575);
nand U5953 (N_5953,N_5458,N_5420);
and U5954 (N_5954,N_5206,N_5298);
nor U5955 (N_5955,N_5338,N_5237);
and U5956 (N_5956,N_5267,N_5202);
nand U5957 (N_5957,N_5340,N_5227);
nor U5958 (N_5958,N_5397,N_5475);
and U5959 (N_5959,N_5307,N_5382);
nor U5960 (N_5960,N_5462,N_5500);
and U5961 (N_5961,N_5283,N_5367);
nor U5962 (N_5962,N_5431,N_5474);
or U5963 (N_5963,N_5341,N_5570);
or U5964 (N_5964,N_5279,N_5369);
nor U5965 (N_5965,N_5495,N_5248);
nand U5966 (N_5966,N_5349,N_5221);
nand U5967 (N_5967,N_5398,N_5451);
and U5968 (N_5968,N_5498,N_5422);
and U5969 (N_5969,N_5568,N_5385);
or U5970 (N_5970,N_5381,N_5392);
nor U5971 (N_5971,N_5539,N_5341);
and U5972 (N_5972,N_5557,N_5524);
or U5973 (N_5973,N_5579,N_5444);
nor U5974 (N_5974,N_5233,N_5526);
or U5975 (N_5975,N_5362,N_5401);
nor U5976 (N_5976,N_5249,N_5343);
and U5977 (N_5977,N_5362,N_5575);
and U5978 (N_5978,N_5320,N_5309);
or U5979 (N_5979,N_5575,N_5596);
nor U5980 (N_5980,N_5294,N_5445);
nand U5981 (N_5981,N_5543,N_5330);
and U5982 (N_5982,N_5501,N_5478);
and U5983 (N_5983,N_5441,N_5368);
or U5984 (N_5984,N_5326,N_5500);
nor U5985 (N_5985,N_5349,N_5275);
nand U5986 (N_5986,N_5541,N_5408);
or U5987 (N_5987,N_5321,N_5388);
or U5988 (N_5988,N_5508,N_5368);
and U5989 (N_5989,N_5340,N_5408);
nand U5990 (N_5990,N_5494,N_5597);
nor U5991 (N_5991,N_5527,N_5215);
nand U5992 (N_5992,N_5490,N_5308);
or U5993 (N_5993,N_5311,N_5565);
nor U5994 (N_5994,N_5320,N_5314);
nor U5995 (N_5995,N_5554,N_5383);
or U5996 (N_5996,N_5448,N_5455);
and U5997 (N_5997,N_5480,N_5430);
nor U5998 (N_5998,N_5221,N_5544);
nand U5999 (N_5999,N_5382,N_5278);
nor U6000 (N_6000,N_5842,N_5927);
nor U6001 (N_6001,N_5967,N_5951);
and U6002 (N_6002,N_5863,N_5788);
nor U6003 (N_6003,N_5745,N_5876);
nand U6004 (N_6004,N_5739,N_5642);
nor U6005 (N_6005,N_5614,N_5632);
or U6006 (N_6006,N_5705,N_5771);
nor U6007 (N_6007,N_5701,N_5791);
nor U6008 (N_6008,N_5982,N_5829);
and U6009 (N_6009,N_5796,N_5601);
and U6010 (N_6010,N_5895,N_5986);
nor U6011 (N_6011,N_5925,N_5960);
nand U6012 (N_6012,N_5975,N_5819);
or U6013 (N_6013,N_5749,N_5779);
nand U6014 (N_6014,N_5893,N_5622);
or U6015 (N_6015,N_5710,N_5688);
or U6016 (N_6016,N_5767,N_5897);
nand U6017 (N_6017,N_5994,N_5912);
nand U6018 (N_6018,N_5811,N_5720);
and U6019 (N_6019,N_5914,N_5718);
or U6020 (N_6020,N_5877,N_5890);
nor U6021 (N_6021,N_5887,N_5643);
nor U6022 (N_6022,N_5706,N_5784);
and U6023 (N_6023,N_5916,N_5915);
or U6024 (N_6024,N_5891,N_5750);
nor U6025 (N_6025,N_5618,N_5786);
or U6026 (N_6026,N_5963,N_5898);
nor U6027 (N_6027,N_5689,N_5792);
or U6028 (N_6028,N_5899,N_5972);
and U6029 (N_6029,N_5755,N_5873);
and U6030 (N_6030,N_5879,N_5735);
and U6031 (N_6031,N_5996,N_5861);
nor U6032 (N_6032,N_5690,N_5657);
or U6033 (N_6033,N_5823,N_5947);
nand U6034 (N_6034,N_5764,N_5874);
nor U6035 (N_6035,N_5797,N_5609);
nand U6036 (N_6036,N_5827,N_5653);
and U6037 (N_6037,N_5644,N_5987);
nand U6038 (N_6038,N_5738,N_5699);
and U6039 (N_6039,N_5984,N_5837);
nor U6040 (N_6040,N_5623,N_5712);
nor U6041 (N_6041,N_5911,N_5978);
and U6042 (N_6042,N_5841,N_5668);
nor U6043 (N_6043,N_5757,N_5789);
or U6044 (N_6044,N_5940,N_5765);
or U6045 (N_6045,N_5851,N_5880);
or U6046 (N_6046,N_5626,N_5651);
and U6047 (N_6047,N_5684,N_5807);
nor U6048 (N_6048,N_5773,N_5950);
and U6049 (N_6049,N_5840,N_5806);
nor U6050 (N_6050,N_5658,N_5781);
nor U6051 (N_6051,N_5969,N_5956);
or U6052 (N_6052,N_5646,N_5721);
or U6053 (N_6053,N_5606,N_5761);
nand U6054 (N_6054,N_5838,N_5681);
nor U6055 (N_6055,N_5962,N_5707);
nand U6056 (N_6056,N_5865,N_5857);
nand U6057 (N_6057,N_5785,N_5920);
and U6058 (N_6058,N_5741,N_5907);
nor U6059 (N_6059,N_5848,N_5926);
or U6060 (N_6060,N_5736,N_5787);
nor U6061 (N_6061,N_5669,N_5654);
nor U6062 (N_6062,N_5812,N_5624);
or U6063 (N_6063,N_5871,N_5989);
or U6064 (N_6064,N_5939,N_5852);
nand U6065 (N_6065,N_5621,N_5656);
nand U6066 (N_6066,N_5748,N_5620);
nand U6067 (N_6067,N_5683,N_5952);
nand U6068 (N_6068,N_5930,N_5869);
or U6069 (N_6069,N_5918,N_5696);
or U6070 (N_6070,N_5846,N_5760);
nand U6071 (N_6071,N_5961,N_5948);
and U6072 (N_6072,N_5875,N_5988);
and U6073 (N_6073,N_5909,N_5850);
or U6074 (N_6074,N_5886,N_5715);
and U6075 (N_6075,N_5900,N_5803);
nand U6076 (N_6076,N_5866,N_5665);
nor U6077 (N_6077,N_5983,N_5763);
or U6078 (N_6078,N_5816,N_5636);
or U6079 (N_6079,N_5999,N_5768);
and U6080 (N_6080,N_5923,N_5769);
nand U6081 (N_6081,N_5700,N_5673);
and U6082 (N_6082,N_5815,N_5800);
and U6083 (N_6083,N_5667,N_5862);
nor U6084 (N_6084,N_5743,N_5966);
or U6085 (N_6085,N_5727,N_5648);
or U6086 (N_6086,N_5835,N_5611);
or U6087 (N_6087,N_5889,N_5725);
or U6088 (N_6088,N_5698,N_5619);
nand U6089 (N_6089,N_5839,N_5600);
or U6090 (N_6090,N_5946,N_5671);
nand U6091 (N_6091,N_5603,N_5659);
nor U6092 (N_6092,N_5808,N_5938);
nor U6093 (N_6093,N_5702,N_5997);
nor U6094 (N_6094,N_5830,N_5828);
and U6095 (N_6095,N_5678,N_5780);
or U6096 (N_6096,N_5809,N_5954);
nand U6097 (N_6097,N_5981,N_5904);
or U6098 (N_6098,N_5697,N_5752);
nand U6099 (N_6099,N_5663,N_5709);
and U6100 (N_6100,N_5722,N_5958);
nand U6101 (N_6101,N_5854,N_5868);
and U6102 (N_6102,N_5836,N_5881);
nand U6103 (N_6103,N_5790,N_5717);
or U6104 (N_6104,N_5856,N_5953);
nor U6105 (N_6105,N_5729,N_5637);
nor U6106 (N_6106,N_5731,N_5759);
nor U6107 (N_6107,N_5936,N_5719);
nor U6108 (N_6108,N_5730,N_5617);
nand U6109 (N_6109,N_5998,N_5903);
or U6110 (N_6110,N_5630,N_5793);
and U6111 (N_6111,N_5977,N_5777);
and U6112 (N_6112,N_5813,N_5616);
nor U6113 (N_6113,N_5728,N_5804);
nand U6114 (N_6114,N_5782,N_5716);
or U6115 (N_6115,N_5666,N_5703);
or U6116 (N_6116,N_5686,N_5919);
or U6117 (N_6117,N_5825,N_5691);
nor U6118 (N_6118,N_5670,N_5753);
nor U6119 (N_6119,N_5645,N_5882);
nor U6120 (N_6120,N_5802,N_5694);
and U6121 (N_6121,N_5737,N_5704);
nand U6122 (N_6122,N_5894,N_5766);
or U6123 (N_6123,N_5860,N_5732);
and U6124 (N_6124,N_5713,N_5992);
nor U6125 (N_6125,N_5831,N_5993);
nand U6126 (N_6126,N_5849,N_5746);
or U6127 (N_6127,N_5845,N_5896);
xnor U6128 (N_6128,N_5995,N_5762);
nor U6129 (N_6129,N_5754,N_5964);
or U6130 (N_6130,N_5607,N_5902);
or U6131 (N_6131,N_5968,N_5708);
and U6132 (N_6132,N_5693,N_5633);
nor U6133 (N_6133,N_5625,N_5641);
nand U6134 (N_6134,N_5959,N_5794);
and U6135 (N_6135,N_5744,N_5685);
nand U6136 (N_6136,N_5833,N_5774);
nand U6137 (N_6137,N_5908,N_5870);
or U6138 (N_6138,N_5884,N_5859);
and U6139 (N_6139,N_5605,N_5855);
nand U6140 (N_6140,N_5628,N_5921);
nor U6141 (N_6141,N_5602,N_5991);
nor U6142 (N_6142,N_5844,N_5979);
nor U6143 (N_6143,N_5935,N_5740);
and U6144 (N_6144,N_5758,N_5649);
nor U6145 (N_6145,N_5858,N_5652);
and U6146 (N_6146,N_5615,N_5957);
or U6147 (N_6147,N_5672,N_5949);
or U6148 (N_6148,N_5726,N_5677);
nor U6149 (N_6149,N_5980,N_5783);
nand U6150 (N_6150,N_5817,N_5734);
nand U6151 (N_6151,N_5610,N_5799);
nor U6152 (N_6152,N_5878,N_5775);
and U6153 (N_6153,N_5627,N_5679);
nor U6154 (N_6154,N_5928,N_5826);
nand U6155 (N_6155,N_5795,N_5660);
nand U6156 (N_6156,N_5824,N_5772);
nor U6157 (N_6157,N_5818,N_5711);
nand U6158 (N_6158,N_5676,N_5942);
or U6159 (N_6159,N_5932,N_5937);
and U6160 (N_6160,N_5650,N_5687);
nor U6161 (N_6161,N_5798,N_5943);
nor U6162 (N_6162,N_5820,N_5747);
nand U6163 (N_6163,N_5631,N_5872);
xor U6164 (N_6164,N_5821,N_5613);
nor U6165 (N_6165,N_5634,N_5955);
or U6166 (N_6166,N_5974,N_5941);
and U6167 (N_6167,N_5913,N_5742);
or U6168 (N_6168,N_5985,N_5864);
and U6169 (N_6169,N_5629,N_5822);
or U6170 (N_6170,N_5810,N_5682);
nor U6171 (N_6171,N_5971,N_5695);
and U6172 (N_6172,N_5885,N_5664);
nand U6173 (N_6173,N_5834,N_5608);
nand U6174 (N_6174,N_5976,N_5883);
nand U6175 (N_6175,N_5814,N_5910);
or U6176 (N_6176,N_5639,N_5724);
nand U6177 (N_6177,N_5612,N_5692);
nor U6178 (N_6178,N_5733,N_5680);
nor U6179 (N_6179,N_5906,N_5945);
nor U6180 (N_6180,N_5970,N_5905);
nand U6181 (N_6181,N_5723,N_5674);
nor U6182 (N_6182,N_5662,N_5832);
or U6183 (N_6183,N_5924,N_5714);
nand U6184 (N_6184,N_5929,N_5604);
or U6185 (N_6185,N_5933,N_5901);
nor U6186 (N_6186,N_5675,N_5944);
nor U6187 (N_6187,N_5655,N_5847);
nand U6188 (N_6188,N_5778,N_5934);
and U6189 (N_6189,N_5922,N_5867);
nand U6190 (N_6190,N_5647,N_5776);
and U6191 (N_6191,N_5770,N_5640);
and U6192 (N_6192,N_5853,N_5917);
nor U6193 (N_6193,N_5888,N_5801);
nand U6194 (N_6194,N_5990,N_5635);
and U6195 (N_6195,N_5965,N_5892);
and U6196 (N_6196,N_5751,N_5931);
or U6197 (N_6197,N_5843,N_5805);
and U6198 (N_6198,N_5638,N_5973);
and U6199 (N_6199,N_5756,N_5661);
and U6200 (N_6200,N_5703,N_5966);
nor U6201 (N_6201,N_5787,N_5777);
nand U6202 (N_6202,N_5899,N_5703);
and U6203 (N_6203,N_5630,N_5752);
and U6204 (N_6204,N_5931,N_5927);
or U6205 (N_6205,N_5702,N_5913);
nand U6206 (N_6206,N_5872,N_5912);
or U6207 (N_6207,N_5925,N_5726);
nor U6208 (N_6208,N_5653,N_5823);
nand U6209 (N_6209,N_5992,N_5873);
and U6210 (N_6210,N_5798,N_5753);
nor U6211 (N_6211,N_5998,N_5694);
and U6212 (N_6212,N_5959,N_5762);
nand U6213 (N_6213,N_5815,N_5727);
nor U6214 (N_6214,N_5784,N_5630);
or U6215 (N_6215,N_5943,N_5725);
nor U6216 (N_6216,N_5727,N_5728);
nand U6217 (N_6217,N_5758,N_5966);
nand U6218 (N_6218,N_5801,N_5723);
and U6219 (N_6219,N_5600,N_5924);
and U6220 (N_6220,N_5847,N_5890);
or U6221 (N_6221,N_5747,N_5738);
xnor U6222 (N_6222,N_5881,N_5740);
nand U6223 (N_6223,N_5750,N_5980);
nor U6224 (N_6224,N_5741,N_5913);
and U6225 (N_6225,N_5988,N_5907);
nand U6226 (N_6226,N_5943,N_5767);
or U6227 (N_6227,N_5657,N_5668);
nand U6228 (N_6228,N_5831,N_5693);
and U6229 (N_6229,N_5768,N_5741);
nand U6230 (N_6230,N_5741,N_5643);
nor U6231 (N_6231,N_5889,N_5799);
or U6232 (N_6232,N_5757,N_5672);
nor U6233 (N_6233,N_5791,N_5975);
nor U6234 (N_6234,N_5899,N_5969);
nand U6235 (N_6235,N_5872,N_5981);
or U6236 (N_6236,N_5804,N_5605);
and U6237 (N_6237,N_5835,N_5829);
nor U6238 (N_6238,N_5949,N_5774);
or U6239 (N_6239,N_5842,N_5978);
nor U6240 (N_6240,N_5843,N_5970);
nand U6241 (N_6241,N_5891,N_5884);
nor U6242 (N_6242,N_5978,N_5776);
and U6243 (N_6243,N_5818,N_5781);
and U6244 (N_6244,N_5658,N_5855);
nor U6245 (N_6245,N_5929,N_5830);
nor U6246 (N_6246,N_5825,N_5689);
and U6247 (N_6247,N_5620,N_5737);
or U6248 (N_6248,N_5982,N_5977);
nand U6249 (N_6249,N_5951,N_5680);
nor U6250 (N_6250,N_5696,N_5961);
nand U6251 (N_6251,N_5827,N_5689);
and U6252 (N_6252,N_5804,N_5754);
nand U6253 (N_6253,N_5646,N_5691);
or U6254 (N_6254,N_5756,N_5867);
nand U6255 (N_6255,N_5977,N_5761);
or U6256 (N_6256,N_5870,N_5739);
or U6257 (N_6257,N_5932,N_5613);
and U6258 (N_6258,N_5889,N_5711);
and U6259 (N_6259,N_5662,N_5804);
nand U6260 (N_6260,N_5908,N_5953);
nand U6261 (N_6261,N_5697,N_5658);
nand U6262 (N_6262,N_5691,N_5729);
or U6263 (N_6263,N_5834,N_5894);
nor U6264 (N_6264,N_5668,N_5695);
and U6265 (N_6265,N_5818,N_5640);
nor U6266 (N_6266,N_5898,N_5816);
or U6267 (N_6267,N_5867,N_5757);
and U6268 (N_6268,N_5850,N_5890);
and U6269 (N_6269,N_5973,N_5710);
nor U6270 (N_6270,N_5916,N_5715);
and U6271 (N_6271,N_5748,N_5993);
or U6272 (N_6272,N_5993,N_5729);
nor U6273 (N_6273,N_5824,N_5760);
or U6274 (N_6274,N_5666,N_5796);
nor U6275 (N_6275,N_5754,N_5778);
or U6276 (N_6276,N_5931,N_5824);
nand U6277 (N_6277,N_5621,N_5883);
nor U6278 (N_6278,N_5752,N_5852);
nand U6279 (N_6279,N_5701,N_5980);
nand U6280 (N_6280,N_5991,N_5664);
or U6281 (N_6281,N_5758,N_5937);
nand U6282 (N_6282,N_5701,N_5901);
or U6283 (N_6283,N_5702,N_5862);
or U6284 (N_6284,N_5896,N_5747);
and U6285 (N_6285,N_5733,N_5667);
and U6286 (N_6286,N_5936,N_5785);
nor U6287 (N_6287,N_5916,N_5997);
nand U6288 (N_6288,N_5605,N_5777);
and U6289 (N_6289,N_5967,N_5707);
nor U6290 (N_6290,N_5950,N_5976);
nand U6291 (N_6291,N_5954,N_5774);
or U6292 (N_6292,N_5620,N_5912);
nor U6293 (N_6293,N_5949,N_5686);
nor U6294 (N_6294,N_5758,N_5651);
or U6295 (N_6295,N_5620,N_5811);
or U6296 (N_6296,N_5772,N_5723);
nand U6297 (N_6297,N_5904,N_5746);
and U6298 (N_6298,N_5646,N_5823);
nor U6299 (N_6299,N_5954,N_5746);
nor U6300 (N_6300,N_5781,N_5626);
nand U6301 (N_6301,N_5668,N_5855);
and U6302 (N_6302,N_5654,N_5734);
or U6303 (N_6303,N_5981,N_5610);
or U6304 (N_6304,N_5772,N_5685);
and U6305 (N_6305,N_5609,N_5883);
and U6306 (N_6306,N_5985,N_5614);
nor U6307 (N_6307,N_5976,N_5764);
or U6308 (N_6308,N_5732,N_5959);
or U6309 (N_6309,N_5833,N_5791);
nor U6310 (N_6310,N_5944,N_5914);
and U6311 (N_6311,N_5618,N_5721);
nor U6312 (N_6312,N_5776,N_5927);
nand U6313 (N_6313,N_5903,N_5676);
and U6314 (N_6314,N_5789,N_5839);
or U6315 (N_6315,N_5957,N_5925);
or U6316 (N_6316,N_5895,N_5605);
or U6317 (N_6317,N_5673,N_5971);
or U6318 (N_6318,N_5698,N_5925);
or U6319 (N_6319,N_5942,N_5808);
or U6320 (N_6320,N_5999,N_5879);
nor U6321 (N_6321,N_5680,N_5873);
and U6322 (N_6322,N_5805,N_5672);
or U6323 (N_6323,N_5774,N_5827);
and U6324 (N_6324,N_5810,N_5878);
xnor U6325 (N_6325,N_5726,N_5762);
nand U6326 (N_6326,N_5704,N_5903);
or U6327 (N_6327,N_5941,N_5802);
or U6328 (N_6328,N_5883,N_5950);
nor U6329 (N_6329,N_5685,N_5897);
and U6330 (N_6330,N_5984,N_5757);
or U6331 (N_6331,N_5711,N_5972);
and U6332 (N_6332,N_5601,N_5635);
nor U6333 (N_6333,N_5745,N_5782);
and U6334 (N_6334,N_5860,N_5776);
or U6335 (N_6335,N_5985,N_5650);
and U6336 (N_6336,N_5681,N_5678);
nor U6337 (N_6337,N_5601,N_5931);
nand U6338 (N_6338,N_5891,N_5617);
or U6339 (N_6339,N_5966,N_5950);
or U6340 (N_6340,N_5958,N_5629);
nand U6341 (N_6341,N_5652,N_5622);
nor U6342 (N_6342,N_5645,N_5651);
nand U6343 (N_6343,N_5713,N_5791);
nor U6344 (N_6344,N_5978,N_5762);
nand U6345 (N_6345,N_5868,N_5990);
nand U6346 (N_6346,N_5818,N_5759);
and U6347 (N_6347,N_5775,N_5958);
and U6348 (N_6348,N_5802,N_5811);
or U6349 (N_6349,N_5921,N_5817);
nor U6350 (N_6350,N_5730,N_5761);
or U6351 (N_6351,N_5634,N_5652);
nand U6352 (N_6352,N_5691,N_5951);
or U6353 (N_6353,N_5911,N_5616);
nand U6354 (N_6354,N_5884,N_5792);
or U6355 (N_6355,N_5741,N_5775);
or U6356 (N_6356,N_5982,N_5706);
nor U6357 (N_6357,N_5817,N_5972);
nor U6358 (N_6358,N_5873,N_5615);
and U6359 (N_6359,N_5951,N_5794);
or U6360 (N_6360,N_5618,N_5604);
and U6361 (N_6361,N_5889,N_5837);
or U6362 (N_6362,N_5798,N_5748);
and U6363 (N_6363,N_5950,N_5756);
or U6364 (N_6364,N_5995,N_5968);
nand U6365 (N_6365,N_5710,N_5677);
nand U6366 (N_6366,N_5997,N_5811);
xor U6367 (N_6367,N_5752,N_5631);
and U6368 (N_6368,N_5976,N_5933);
or U6369 (N_6369,N_5829,N_5637);
or U6370 (N_6370,N_5882,N_5971);
or U6371 (N_6371,N_5628,N_5753);
nor U6372 (N_6372,N_5814,N_5663);
nand U6373 (N_6373,N_5875,N_5968);
nor U6374 (N_6374,N_5926,N_5750);
and U6375 (N_6375,N_5730,N_5940);
or U6376 (N_6376,N_5932,N_5984);
or U6377 (N_6377,N_5684,N_5898);
nand U6378 (N_6378,N_5958,N_5605);
or U6379 (N_6379,N_5853,N_5940);
nand U6380 (N_6380,N_5977,N_5633);
nand U6381 (N_6381,N_5731,N_5872);
or U6382 (N_6382,N_5719,N_5737);
nand U6383 (N_6383,N_5712,N_5602);
or U6384 (N_6384,N_5959,N_5755);
nand U6385 (N_6385,N_5871,N_5865);
nor U6386 (N_6386,N_5821,N_5987);
nand U6387 (N_6387,N_5753,N_5727);
or U6388 (N_6388,N_5790,N_5744);
and U6389 (N_6389,N_5906,N_5893);
and U6390 (N_6390,N_5859,N_5827);
nand U6391 (N_6391,N_5796,N_5677);
nor U6392 (N_6392,N_5600,N_5751);
nand U6393 (N_6393,N_5789,N_5847);
and U6394 (N_6394,N_5838,N_5916);
nor U6395 (N_6395,N_5738,N_5686);
nand U6396 (N_6396,N_5809,N_5798);
nor U6397 (N_6397,N_5991,N_5881);
nand U6398 (N_6398,N_5628,N_5636);
and U6399 (N_6399,N_5901,N_5616);
nand U6400 (N_6400,N_6097,N_6101);
nor U6401 (N_6401,N_6047,N_6172);
or U6402 (N_6402,N_6324,N_6376);
nor U6403 (N_6403,N_6132,N_6086);
nor U6404 (N_6404,N_6362,N_6010);
nor U6405 (N_6405,N_6291,N_6051);
or U6406 (N_6406,N_6219,N_6107);
nand U6407 (N_6407,N_6346,N_6260);
nor U6408 (N_6408,N_6121,N_6142);
and U6409 (N_6409,N_6261,N_6072);
or U6410 (N_6410,N_6082,N_6158);
xnor U6411 (N_6411,N_6169,N_6211);
nand U6412 (N_6412,N_6202,N_6012);
and U6413 (N_6413,N_6256,N_6125);
and U6414 (N_6414,N_6283,N_6371);
nand U6415 (N_6415,N_6109,N_6159);
and U6416 (N_6416,N_6166,N_6286);
and U6417 (N_6417,N_6262,N_6021);
nor U6418 (N_6418,N_6041,N_6223);
or U6419 (N_6419,N_6066,N_6395);
nor U6420 (N_6420,N_6263,N_6322);
nor U6421 (N_6421,N_6009,N_6329);
and U6422 (N_6422,N_6335,N_6191);
or U6423 (N_6423,N_6083,N_6186);
and U6424 (N_6424,N_6251,N_6259);
nand U6425 (N_6425,N_6278,N_6111);
nand U6426 (N_6426,N_6077,N_6019);
or U6427 (N_6427,N_6363,N_6124);
and U6428 (N_6428,N_6060,N_6252);
nand U6429 (N_6429,N_6373,N_6198);
nand U6430 (N_6430,N_6178,N_6182);
or U6431 (N_6431,N_6184,N_6225);
nor U6432 (N_6432,N_6217,N_6315);
nor U6433 (N_6433,N_6087,N_6255);
or U6434 (N_6434,N_6033,N_6175);
nand U6435 (N_6435,N_6037,N_6200);
or U6436 (N_6436,N_6079,N_6243);
nand U6437 (N_6437,N_6341,N_6030);
or U6438 (N_6438,N_6215,N_6145);
and U6439 (N_6439,N_6342,N_6026);
nand U6440 (N_6440,N_6314,N_6359);
and U6441 (N_6441,N_6059,N_6129);
and U6442 (N_6442,N_6284,N_6053);
nor U6443 (N_6443,N_6323,N_6011);
nor U6444 (N_6444,N_6375,N_6289);
nand U6445 (N_6445,N_6133,N_6234);
nand U6446 (N_6446,N_6282,N_6366);
nor U6447 (N_6447,N_6193,N_6056);
and U6448 (N_6448,N_6380,N_6139);
nand U6449 (N_6449,N_6365,N_6049);
or U6450 (N_6450,N_6239,N_6295);
or U6451 (N_6451,N_6005,N_6013);
nand U6452 (N_6452,N_6331,N_6271);
or U6453 (N_6453,N_6247,N_6391);
nand U6454 (N_6454,N_6212,N_6078);
or U6455 (N_6455,N_6112,N_6382);
and U6456 (N_6456,N_6280,N_6088);
nand U6457 (N_6457,N_6258,N_6165);
nor U6458 (N_6458,N_6339,N_6214);
or U6459 (N_6459,N_6361,N_6020);
and U6460 (N_6460,N_6250,N_6140);
and U6461 (N_6461,N_6038,N_6045);
or U6462 (N_6462,N_6245,N_6277);
and U6463 (N_6463,N_6167,N_6096);
and U6464 (N_6464,N_6170,N_6242);
and U6465 (N_6465,N_6399,N_6270);
nand U6466 (N_6466,N_6292,N_6398);
nand U6467 (N_6467,N_6321,N_6151);
nand U6468 (N_6468,N_6057,N_6143);
or U6469 (N_6469,N_6226,N_6073);
and U6470 (N_6470,N_6328,N_6094);
and U6471 (N_6471,N_6296,N_6352);
nor U6472 (N_6472,N_6288,N_6055);
nand U6473 (N_6473,N_6067,N_6332);
and U6474 (N_6474,N_6188,N_6034);
nand U6475 (N_6475,N_6189,N_6171);
nand U6476 (N_6476,N_6377,N_6353);
nand U6477 (N_6477,N_6046,N_6205);
or U6478 (N_6478,N_6192,N_6108);
nand U6479 (N_6479,N_6075,N_6357);
nand U6480 (N_6480,N_6319,N_6199);
and U6481 (N_6481,N_6048,N_6181);
nor U6482 (N_6482,N_6179,N_6320);
or U6483 (N_6483,N_6150,N_6340);
or U6484 (N_6484,N_6122,N_6378);
nor U6485 (N_6485,N_6275,N_6136);
and U6486 (N_6486,N_6274,N_6204);
and U6487 (N_6487,N_6209,N_6264);
or U6488 (N_6488,N_6155,N_6338);
nor U6489 (N_6489,N_6031,N_6257);
or U6490 (N_6490,N_6210,N_6311);
and U6491 (N_6491,N_6302,N_6134);
nor U6492 (N_6492,N_6146,N_6253);
or U6493 (N_6493,N_6232,N_6036);
or U6494 (N_6494,N_6091,N_6392);
nand U6495 (N_6495,N_6074,N_6195);
nor U6496 (N_6496,N_6333,N_6208);
xnor U6497 (N_6497,N_6309,N_6039);
or U6498 (N_6498,N_6160,N_6387);
or U6499 (N_6499,N_6114,N_6183);
and U6500 (N_6500,N_6196,N_6233);
or U6501 (N_6501,N_6203,N_6100);
nor U6502 (N_6502,N_6393,N_6099);
and U6503 (N_6503,N_6093,N_6326);
nor U6504 (N_6504,N_6040,N_6222);
or U6505 (N_6505,N_6297,N_6218);
and U6506 (N_6506,N_6081,N_6236);
nand U6507 (N_6507,N_6207,N_6374);
or U6508 (N_6508,N_6098,N_6002);
nor U6509 (N_6509,N_6349,N_6069);
nor U6510 (N_6510,N_6241,N_6367);
nand U6511 (N_6511,N_6293,N_6187);
nand U6512 (N_6512,N_6384,N_6113);
nor U6513 (N_6513,N_6254,N_6272);
or U6514 (N_6514,N_6344,N_6154);
nor U6515 (N_6515,N_6213,N_6070);
or U6516 (N_6516,N_6206,N_6080);
and U6517 (N_6517,N_6042,N_6246);
or U6518 (N_6518,N_6281,N_6156);
nand U6519 (N_6519,N_6138,N_6318);
and U6520 (N_6520,N_6240,N_6058);
nand U6521 (N_6521,N_6001,N_6249);
nor U6522 (N_6522,N_6054,N_6347);
or U6523 (N_6523,N_6294,N_6032);
or U6524 (N_6524,N_6383,N_6244);
nor U6525 (N_6525,N_6161,N_6117);
or U6526 (N_6526,N_6174,N_6024);
nor U6527 (N_6527,N_6168,N_6052);
nor U6528 (N_6528,N_6220,N_6381);
nor U6529 (N_6529,N_6364,N_6325);
nor U6530 (N_6530,N_6316,N_6290);
nor U6531 (N_6531,N_6265,N_6299);
nand U6532 (N_6532,N_6164,N_6103);
nor U6533 (N_6533,N_6229,N_6317);
nor U6534 (N_6534,N_6016,N_6076);
nor U6535 (N_6535,N_6388,N_6372);
nand U6536 (N_6536,N_6095,N_6354);
xnor U6537 (N_6537,N_6235,N_6023);
and U6538 (N_6538,N_6084,N_6137);
and U6539 (N_6539,N_6303,N_6287);
nor U6540 (N_6540,N_6268,N_6000);
or U6541 (N_6541,N_6089,N_6221);
nand U6542 (N_6542,N_6301,N_6141);
or U6543 (N_6543,N_6014,N_6368);
or U6544 (N_6544,N_6279,N_6304);
and U6545 (N_6545,N_6063,N_6153);
or U6546 (N_6546,N_6120,N_6201);
and U6547 (N_6547,N_6131,N_6334);
nor U6548 (N_6548,N_6064,N_6285);
nor U6549 (N_6549,N_6061,N_6119);
and U6550 (N_6550,N_6248,N_6118);
nor U6551 (N_6551,N_6231,N_6018);
or U6552 (N_6552,N_6152,N_6337);
and U6553 (N_6553,N_6298,N_6327);
nand U6554 (N_6554,N_6173,N_6050);
and U6555 (N_6555,N_6345,N_6148);
and U6556 (N_6556,N_6035,N_6043);
nor U6557 (N_6557,N_6115,N_6090);
nand U6558 (N_6558,N_6369,N_6228);
and U6559 (N_6559,N_6276,N_6025);
nand U6560 (N_6560,N_6007,N_6238);
and U6561 (N_6561,N_6062,N_6343);
or U6562 (N_6562,N_6227,N_6300);
nor U6563 (N_6563,N_6336,N_6135);
nand U6564 (N_6564,N_6180,N_6102);
nor U6565 (N_6565,N_6389,N_6348);
and U6566 (N_6566,N_6351,N_6029);
nor U6567 (N_6567,N_6106,N_6104);
and U6568 (N_6568,N_6386,N_6397);
or U6569 (N_6569,N_6273,N_6163);
and U6570 (N_6570,N_6379,N_6355);
nand U6571 (N_6571,N_6123,N_6190);
nand U6572 (N_6572,N_6267,N_6350);
nand U6573 (N_6573,N_6216,N_6224);
nor U6574 (N_6574,N_6157,N_6330);
or U6575 (N_6575,N_6004,N_6008);
and U6576 (N_6576,N_6307,N_6015);
nor U6577 (N_6577,N_6360,N_6394);
and U6578 (N_6578,N_6312,N_6194);
nor U6579 (N_6579,N_6105,N_6313);
nor U6580 (N_6580,N_6127,N_6065);
nand U6581 (N_6581,N_6110,N_6128);
and U6582 (N_6582,N_6068,N_6147);
or U6583 (N_6583,N_6162,N_6266);
and U6584 (N_6584,N_6085,N_6305);
or U6585 (N_6585,N_6022,N_6176);
or U6586 (N_6586,N_6385,N_6028);
nor U6587 (N_6587,N_6126,N_6370);
nor U6588 (N_6588,N_6144,N_6177);
nand U6589 (N_6589,N_6396,N_6358);
and U6590 (N_6590,N_6197,N_6237);
or U6591 (N_6591,N_6306,N_6017);
and U6592 (N_6592,N_6310,N_6390);
nor U6593 (N_6593,N_6185,N_6130);
nand U6594 (N_6594,N_6116,N_6356);
or U6595 (N_6595,N_6269,N_6044);
nand U6596 (N_6596,N_6092,N_6003);
nor U6597 (N_6597,N_6230,N_6006);
nand U6598 (N_6598,N_6071,N_6308);
and U6599 (N_6599,N_6149,N_6027);
and U6600 (N_6600,N_6228,N_6101);
and U6601 (N_6601,N_6095,N_6021);
or U6602 (N_6602,N_6274,N_6171);
or U6603 (N_6603,N_6360,N_6315);
or U6604 (N_6604,N_6359,N_6195);
nor U6605 (N_6605,N_6131,N_6399);
nor U6606 (N_6606,N_6182,N_6391);
nor U6607 (N_6607,N_6186,N_6357);
nand U6608 (N_6608,N_6096,N_6393);
nor U6609 (N_6609,N_6107,N_6233);
or U6610 (N_6610,N_6374,N_6163);
or U6611 (N_6611,N_6065,N_6228);
and U6612 (N_6612,N_6069,N_6382);
and U6613 (N_6613,N_6226,N_6172);
or U6614 (N_6614,N_6184,N_6271);
and U6615 (N_6615,N_6376,N_6295);
nand U6616 (N_6616,N_6087,N_6175);
nor U6617 (N_6617,N_6035,N_6031);
nor U6618 (N_6618,N_6250,N_6312);
or U6619 (N_6619,N_6277,N_6138);
nand U6620 (N_6620,N_6338,N_6181);
nor U6621 (N_6621,N_6188,N_6305);
and U6622 (N_6622,N_6260,N_6140);
or U6623 (N_6623,N_6389,N_6104);
nand U6624 (N_6624,N_6392,N_6064);
nand U6625 (N_6625,N_6098,N_6304);
nor U6626 (N_6626,N_6288,N_6278);
or U6627 (N_6627,N_6244,N_6229);
nor U6628 (N_6628,N_6368,N_6297);
nor U6629 (N_6629,N_6088,N_6229);
nand U6630 (N_6630,N_6231,N_6317);
nor U6631 (N_6631,N_6048,N_6164);
nor U6632 (N_6632,N_6044,N_6226);
or U6633 (N_6633,N_6385,N_6146);
nor U6634 (N_6634,N_6046,N_6219);
and U6635 (N_6635,N_6229,N_6093);
nand U6636 (N_6636,N_6188,N_6263);
nand U6637 (N_6637,N_6169,N_6146);
nand U6638 (N_6638,N_6056,N_6236);
nand U6639 (N_6639,N_6311,N_6294);
nor U6640 (N_6640,N_6153,N_6136);
nor U6641 (N_6641,N_6090,N_6086);
nand U6642 (N_6642,N_6297,N_6223);
nor U6643 (N_6643,N_6317,N_6375);
and U6644 (N_6644,N_6069,N_6301);
and U6645 (N_6645,N_6346,N_6261);
nand U6646 (N_6646,N_6003,N_6032);
nor U6647 (N_6647,N_6291,N_6079);
and U6648 (N_6648,N_6043,N_6221);
and U6649 (N_6649,N_6080,N_6286);
and U6650 (N_6650,N_6056,N_6391);
nor U6651 (N_6651,N_6343,N_6100);
and U6652 (N_6652,N_6150,N_6053);
and U6653 (N_6653,N_6031,N_6186);
and U6654 (N_6654,N_6358,N_6383);
nand U6655 (N_6655,N_6100,N_6303);
or U6656 (N_6656,N_6054,N_6025);
nor U6657 (N_6657,N_6024,N_6183);
or U6658 (N_6658,N_6124,N_6095);
nand U6659 (N_6659,N_6313,N_6348);
or U6660 (N_6660,N_6001,N_6266);
nand U6661 (N_6661,N_6276,N_6130);
nand U6662 (N_6662,N_6343,N_6211);
xor U6663 (N_6663,N_6361,N_6011);
or U6664 (N_6664,N_6300,N_6242);
and U6665 (N_6665,N_6265,N_6209);
nand U6666 (N_6666,N_6391,N_6140);
or U6667 (N_6667,N_6198,N_6168);
or U6668 (N_6668,N_6383,N_6156);
or U6669 (N_6669,N_6313,N_6133);
nand U6670 (N_6670,N_6105,N_6233);
nor U6671 (N_6671,N_6119,N_6147);
and U6672 (N_6672,N_6200,N_6270);
nand U6673 (N_6673,N_6315,N_6118);
and U6674 (N_6674,N_6074,N_6221);
or U6675 (N_6675,N_6173,N_6074);
or U6676 (N_6676,N_6029,N_6390);
nor U6677 (N_6677,N_6281,N_6170);
nand U6678 (N_6678,N_6395,N_6155);
or U6679 (N_6679,N_6324,N_6218);
and U6680 (N_6680,N_6011,N_6082);
nand U6681 (N_6681,N_6316,N_6001);
and U6682 (N_6682,N_6164,N_6168);
nor U6683 (N_6683,N_6302,N_6129);
nor U6684 (N_6684,N_6017,N_6042);
xor U6685 (N_6685,N_6347,N_6278);
xor U6686 (N_6686,N_6130,N_6215);
or U6687 (N_6687,N_6301,N_6390);
nor U6688 (N_6688,N_6358,N_6110);
or U6689 (N_6689,N_6291,N_6085);
nor U6690 (N_6690,N_6221,N_6384);
nand U6691 (N_6691,N_6186,N_6173);
nand U6692 (N_6692,N_6240,N_6122);
nor U6693 (N_6693,N_6141,N_6364);
xor U6694 (N_6694,N_6326,N_6216);
nand U6695 (N_6695,N_6182,N_6378);
nor U6696 (N_6696,N_6119,N_6378);
nand U6697 (N_6697,N_6224,N_6191);
or U6698 (N_6698,N_6114,N_6118);
or U6699 (N_6699,N_6058,N_6312);
nand U6700 (N_6700,N_6290,N_6341);
or U6701 (N_6701,N_6272,N_6316);
and U6702 (N_6702,N_6391,N_6226);
or U6703 (N_6703,N_6039,N_6065);
or U6704 (N_6704,N_6370,N_6215);
nand U6705 (N_6705,N_6132,N_6358);
nand U6706 (N_6706,N_6148,N_6203);
nand U6707 (N_6707,N_6212,N_6386);
and U6708 (N_6708,N_6216,N_6375);
or U6709 (N_6709,N_6252,N_6283);
nor U6710 (N_6710,N_6157,N_6207);
and U6711 (N_6711,N_6027,N_6070);
nand U6712 (N_6712,N_6389,N_6394);
nor U6713 (N_6713,N_6396,N_6111);
or U6714 (N_6714,N_6203,N_6126);
nand U6715 (N_6715,N_6145,N_6176);
and U6716 (N_6716,N_6137,N_6160);
or U6717 (N_6717,N_6382,N_6261);
or U6718 (N_6718,N_6077,N_6291);
nor U6719 (N_6719,N_6364,N_6300);
nand U6720 (N_6720,N_6256,N_6220);
or U6721 (N_6721,N_6160,N_6366);
and U6722 (N_6722,N_6225,N_6117);
nand U6723 (N_6723,N_6049,N_6315);
nand U6724 (N_6724,N_6084,N_6024);
or U6725 (N_6725,N_6200,N_6147);
or U6726 (N_6726,N_6227,N_6344);
nand U6727 (N_6727,N_6138,N_6072);
or U6728 (N_6728,N_6367,N_6206);
nor U6729 (N_6729,N_6215,N_6055);
nor U6730 (N_6730,N_6298,N_6025);
and U6731 (N_6731,N_6110,N_6152);
and U6732 (N_6732,N_6362,N_6371);
and U6733 (N_6733,N_6107,N_6118);
nor U6734 (N_6734,N_6260,N_6350);
or U6735 (N_6735,N_6378,N_6031);
and U6736 (N_6736,N_6018,N_6264);
and U6737 (N_6737,N_6275,N_6043);
or U6738 (N_6738,N_6181,N_6176);
nor U6739 (N_6739,N_6336,N_6394);
nor U6740 (N_6740,N_6319,N_6147);
nor U6741 (N_6741,N_6116,N_6285);
nor U6742 (N_6742,N_6037,N_6169);
nor U6743 (N_6743,N_6121,N_6127);
nand U6744 (N_6744,N_6198,N_6181);
or U6745 (N_6745,N_6342,N_6332);
nand U6746 (N_6746,N_6024,N_6132);
nor U6747 (N_6747,N_6308,N_6122);
or U6748 (N_6748,N_6391,N_6305);
or U6749 (N_6749,N_6277,N_6151);
nor U6750 (N_6750,N_6020,N_6129);
and U6751 (N_6751,N_6163,N_6317);
nor U6752 (N_6752,N_6338,N_6130);
and U6753 (N_6753,N_6293,N_6221);
or U6754 (N_6754,N_6174,N_6288);
and U6755 (N_6755,N_6205,N_6043);
or U6756 (N_6756,N_6341,N_6228);
nor U6757 (N_6757,N_6064,N_6319);
nand U6758 (N_6758,N_6109,N_6029);
or U6759 (N_6759,N_6081,N_6098);
nor U6760 (N_6760,N_6190,N_6288);
and U6761 (N_6761,N_6377,N_6258);
or U6762 (N_6762,N_6208,N_6307);
nor U6763 (N_6763,N_6227,N_6011);
and U6764 (N_6764,N_6320,N_6233);
or U6765 (N_6765,N_6019,N_6244);
nand U6766 (N_6766,N_6009,N_6268);
or U6767 (N_6767,N_6261,N_6390);
or U6768 (N_6768,N_6032,N_6028);
or U6769 (N_6769,N_6110,N_6223);
nand U6770 (N_6770,N_6159,N_6379);
and U6771 (N_6771,N_6169,N_6369);
nor U6772 (N_6772,N_6339,N_6397);
or U6773 (N_6773,N_6152,N_6165);
nor U6774 (N_6774,N_6138,N_6187);
or U6775 (N_6775,N_6161,N_6374);
nor U6776 (N_6776,N_6299,N_6053);
or U6777 (N_6777,N_6112,N_6372);
nor U6778 (N_6778,N_6247,N_6340);
nand U6779 (N_6779,N_6084,N_6085);
nor U6780 (N_6780,N_6102,N_6090);
and U6781 (N_6781,N_6352,N_6272);
nand U6782 (N_6782,N_6282,N_6353);
or U6783 (N_6783,N_6086,N_6040);
or U6784 (N_6784,N_6362,N_6105);
and U6785 (N_6785,N_6101,N_6325);
nor U6786 (N_6786,N_6089,N_6021);
xor U6787 (N_6787,N_6013,N_6022);
nor U6788 (N_6788,N_6127,N_6119);
or U6789 (N_6789,N_6390,N_6362);
nor U6790 (N_6790,N_6311,N_6022);
and U6791 (N_6791,N_6120,N_6147);
nor U6792 (N_6792,N_6171,N_6163);
or U6793 (N_6793,N_6190,N_6211);
and U6794 (N_6794,N_6384,N_6238);
and U6795 (N_6795,N_6255,N_6108);
and U6796 (N_6796,N_6040,N_6078);
nor U6797 (N_6797,N_6166,N_6079);
or U6798 (N_6798,N_6229,N_6295);
and U6799 (N_6799,N_6233,N_6198);
and U6800 (N_6800,N_6698,N_6631);
and U6801 (N_6801,N_6718,N_6666);
nor U6802 (N_6802,N_6525,N_6764);
nor U6803 (N_6803,N_6412,N_6438);
nand U6804 (N_6804,N_6475,N_6783);
and U6805 (N_6805,N_6639,N_6683);
or U6806 (N_6806,N_6780,N_6401);
and U6807 (N_6807,N_6769,N_6744);
or U6808 (N_6808,N_6479,N_6507);
or U6809 (N_6809,N_6502,N_6561);
and U6810 (N_6810,N_6721,N_6456);
or U6811 (N_6811,N_6523,N_6573);
or U6812 (N_6812,N_6633,N_6776);
or U6813 (N_6813,N_6680,N_6459);
and U6814 (N_6814,N_6681,N_6733);
or U6815 (N_6815,N_6710,N_6537);
or U6816 (N_6816,N_6553,N_6434);
nand U6817 (N_6817,N_6725,N_6752);
and U6818 (N_6818,N_6559,N_6761);
and U6819 (N_6819,N_6758,N_6403);
or U6820 (N_6820,N_6748,N_6707);
or U6821 (N_6821,N_6447,N_6518);
or U6822 (N_6822,N_6599,N_6751);
nand U6823 (N_6823,N_6597,N_6706);
or U6824 (N_6824,N_6612,N_6477);
nand U6825 (N_6825,N_6539,N_6750);
nand U6826 (N_6826,N_6689,N_6517);
nor U6827 (N_6827,N_6515,N_6510);
and U6828 (N_6828,N_6608,N_6560);
and U6829 (N_6829,N_6749,N_6448);
and U6830 (N_6830,N_6745,N_6732);
nor U6831 (N_6831,N_6742,N_6670);
or U6832 (N_6832,N_6641,N_6770);
and U6833 (N_6833,N_6419,N_6674);
nor U6834 (N_6834,N_6413,N_6684);
and U6835 (N_6835,N_6593,N_6509);
and U6836 (N_6836,N_6657,N_6577);
nor U6837 (N_6837,N_6486,N_6695);
nand U6838 (N_6838,N_6451,N_6627);
and U6839 (N_6839,N_6554,N_6431);
and U6840 (N_6840,N_6501,N_6402);
nor U6841 (N_6841,N_6566,N_6784);
nor U6842 (N_6842,N_6587,N_6708);
and U6843 (N_6843,N_6555,N_6636);
xor U6844 (N_6844,N_6632,N_6478);
nand U6845 (N_6845,N_6755,N_6454);
nand U6846 (N_6846,N_6427,N_6669);
and U6847 (N_6847,N_6583,N_6663);
nand U6848 (N_6848,N_6647,N_6425);
and U6849 (N_6849,N_6580,N_6405);
nor U6850 (N_6850,N_6458,N_6495);
nand U6851 (N_6851,N_6659,N_6508);
or U6852 (N_6852,N_6439,N_6487);
nand U6853 (N_6853,N_6450,N_6716);
and U6854 (N_6854,N_6430,N_6704);
xor U6855 (N_6855,N_6414,N_6685);
nand U6856 (N_6856,N_6420,N_6463);
or U6857 (N_6857,N_6584,N_6714);
nor U6858 (N_6858,N_6675,N_6775);
nand U6859 (N_6859,N_6408,N_6490);
nor U6860 (N_6860,N_6505,N_6773);
and U6861 (N_6861,N_6452,N_6529);
nand U6862 (N_6862,N_6422,N_6796);
nor U6863 (N_6863,N_6467,N_6491);
or U6864 (N_6864,N_6480,N_6544);
nand U6865 (N_6865,N_6794,N_6562);
or U6866 (N_6866,N_6741,N_6492);
and U6867 (N_6867,N_6446,N_6441);
xor U6868 (N_6868,N_6581,N_6740);
nor U6869 (N_6869,N_6609,N_6570);
nor U6870 (N_6870,N_6410,N_6563);
or U6871 (N_6871,N_6760,N_6528);
and U6872 (N_6872,N_6791,N_6432);
or U6873 (N_6873,N_6453,N_6585);
nor U6874 (N_6874,N_6664,N_6460);
and U6875 (N_6875,N_6542,N_6603);
nor U6876 (N_6876,N_6653,N_6620);
or U6877 (N_6877,N_6787,N_6437);
or U6878 (N_6878,N_6634,N_6404);
and U6879 (N_6879,N_6702,N_6496);
nor U6880 (N_6880,N_6682,N_6737);
or U6881 (N_6881,N_6457,N_6499);
nor U6882 (N_6882,N_6615,N_6556);
and U6883 (N_6883,N_6646,N_6435);
and U6884 (N_6884,N_6652,N_6471);
nand U6885 (N_6885,N_6739,N_6619);
nand U6886 (N_6886,N_6688,N_6734);
nor U6887 (N_6887,N_6527,N_6648);
and U6888 (N_6888,N_6598,N_6595);
and U6889 (N_6889,N_6763,N_6483);
nand U6890 (N_6890,N_6484,N_6416);
or U6891 (N_6891,N_6444,N_6645);
nand U6892 (N_6892,N_6582,N_6579);
nor U6893 (N_6893,N_6602,N_6470);
nand U6894 (N_6894,N_6743,N_6601);
and U6895 (N_6895,N_6443,N_6638);
or U6896 (N_6896,N_6735,N_6482);
or U6897 (N_6897,N_6694,N_6747);
nor U6898 (N_6898,N_6738,N_6798);
or U6899 (N_6899,N_6606,N_6488);
and U6900 (N_6900,N_6626,N_6726);
or U6901 (N_6901,N_6692,N_6771);
nor U6902 (N_6902,N_6790,N_6709);
or U6903 (N_6903,N_6711,N_6665);
or U6904 (N_6904,N_6530,N_6691);
and U6905 (N_6905,N_6567,N_6618);
and U6906 (N_6906,N_6616,N_6712);
or U6907 (N_6907,N_6569,N_6531);
and U6908 (N_6908,N_6594,N_6536);
nor U6909 (N_6909,N_6696,N_6604);
nor U6910 (N_6910,N_6736,N_6406);
or U6911 (N_6911,N_6719,N_6503);
nand U6912 (N_6912,N_6651,N_6588);
and U6913 (N_6913,N_6565,N_6779);
nor U6914 (N_6914,N_6644,N_6468);
nand U6915 (N_6915,N_6538,N_6524);
xor U6916 (N_6916,N_6642,N_6715);
nor U6917 (N_6917,N_6596,N_6591);
and U6918 (N_6918,N_6455,N_6564);
nand U6919 (N_6919,N_6407,N_6720);
nor U6920 (N_6920,N_6759,N_6624);
nor U6921 (N_6921,N_6557,N_6500);
nor U6922 (N_6922,N_6762,N_6799);
and U6923 (N_6923,N_6436,N_6723);
or U6924 (N_6924,N_6550,N_6672);
nand U6925 (N_6925,N_6793,N_6476);
or U6926 (N_6926,N_6429,N_6534);
and U6927 (N_6927,N_6440,N_6650);
nor U6928 (N_6928,N_6772,N_6679);
nor U6929 (N_6929,N_6717,N_6660);
nor U6930 (N_6930,N_6673,N_6705);
or U6931 (N_6931,N_6797,N_6415);
and U6932 (N_6932,N_6513,N_6605);
nand U6933 (N_6933,N_6781,N_6466);
and U6934 (N_6934,N_6535,N_6722);
or U6935 (N_6935,N_6774,N_6592);
nor U6936 (N_6936,N_6661,N_6678);
nor U6937 (N_6937,N_6782,N_6445);
nand U6938 (N_6938,N_6754,N_6610);
nand U6939 (N_6939,N_6789,N_6469);
and U6940 (N_6940,N_6767,N_6586);
nor U6941 (N_6941,N_6549,N_6558);
or U6942 (N_6942,N_6611,N_6568);
nor U6943 (N_6943,N_6727,N_6600);
or U6944 (N_6944,N_6623,N_6643);
and U6945 (N_6945,N_6428,N_6654);
nor U6946 (N_6946,N_6551,N_6526);
nor U6947 (N_6947,N_6697,N_6788);
nand U6948 (N_6948,N_6617,N_6520);
nand U6949 (N_6949,N_6677,N_6589);
and U6950 (N_6950,N_6543,N_6786);
or U6951 (N_6951,N_6686,N_6671);
and U6952 (N_6952,N_6699,N_6655);
nor U6953 (N_6953,N_6700,N_6637);
nand U6954 (N_6954,N_6522,N_6630);
nand U6955 (N_6955,N_6497,N_6622);
nand U6956 (N_6956,N_6607,N_6629);
and U6957 (N_6957,N_6656,N_6703);
nand U6958 (N_6958,N_6713,N_6576);
nand U6959 (N_6959,N_6621,N_6512);
nand U6960 (N_6960,N_6730,N_6668);
nor U6961 (N_6961,N_6521,N_6548);
nor U6962 (N_6962,N_6461,N_6417);
or U6963 (N_6963,N_6777,N_6792);
and U6964 (N_6964,N_6540,N_6728);
and U6965 (N_6965,N_6546,N_6552);
or U6966 (N_6966,N_6640,N_6731);
or U6967 (N_6967,N_6424,N_6693);
nand U6968 (N_6968,N_6474,N_6473);
or U6969 (N_6969,N_6768,N_6409);
nand U6970 (N_6970,N_6423,N_6613);
or U6971 (N_6971,N_6433,N_6545);
nor U6972 (N_6972,N_6571,N_6785);
or U6973 (N_6973,N_6493,N_6514);
or U6974 (N_6974,N_6578,N_6778);
or U6975 (N_6975,N_6472,N_6511);
nand U6976 (N_6976,N_6662,N_6442);
xor U6977 (N_6977,N_6421,N_6449);
nand U6978 (N_6978,N_6485,N_6462);
nand U6979 (N_6979,N_6614,N_6547);
nor U6980 (N_6980,N_6690,N_6519);
or U6981 (N_6981,N_6516,N_6757);
nor U6982 (N_6982,N_6687,N_6498);
nor U6983 (N_6983,N_6746,N_6481);
nor U6984 (N_6984,N_6572,N_6494);
xnor U6985 (N_6985,N_6756,N_6575);
nor U6986 (N_6986,N_6753,N_6724);
nand U6987 (N_6987,N_6766,N_6489);
and U6988 (N_6988,N_6729,N_6628);
or U6989 (N_6989,N_6504,N_6701);
nand U6990 (N_6990,N_6667,N_6649);
nor U6991 (N_6991,N_6765,N_6533);
and U6992 (N_6992,N_6506,N_6464);
or U6993 (N_6993,N_6795,N_6465);
or U6994 (N_6994,N_6426,N_6635);
xnor U6995 (N_6995,N_6625,N_6541);
and U6996 (N_6996,N_6590,N_6532);
nand U6997 (N_6997,N_6411,N_6574);
nor U6998 (N_6998,N_6658,N_6676);
and U6999 (N_6999,N_6400,N_6418);
and U7000 (N_7000,N_6578,N_6646);
and U7001 (N_7001,N_6722,N_6578);
nand U7002 (N_7002,N_6482,N_6741);
and U7003 (N_7003,N_6580,N_6402);
nor U7004 (N_7004,N_6401,N_6660);
nand U7005 (N_7005,N_6732,N_6636);
or U7006 (N_7006,N_6746,N_6742);
nor U7007 (N_7007,N_6472,N_6464);
and U7008 (N_7008,N_6696,N_6520);
nor U7009 (N_7009,N_6668,N_6700);
nand U7010 (N_7010,N_6563,N_6795);
nor U7011 (N_7011,N_6566,N_6450);
and U7012 (N_7012,N_6550,N_6754);
nand U7013 (N_7013,N_6703,N_6608);
or U7014 (N_7014,N_6746,N_6503);
nor U7015 (N_7015,N_6434,N_6523);
and U7016 (N_7016,N_6446,N_6522);
nand U7017 (N_7017,N_6779,N_6590);
or U7018 (N_7018,N_6476,N_6537);
and U7019 (N_7019,N_6476,N_6659);
nand U7020 (N_7020,N_6662,N_6535);
nor U7021 (N_7021,N_6763,N_6641);
and U7022 (N_7022,N_6714,N_6753);
and U7023 (N_7023,N_6639,N_6600);
nand U7024 (N_7024,N_6692,N_6719);
nor U7025 (N_7025,N_6752,N_6772);
nand U7026 (N_7026,N_6607,N_6504);
or U7027 (N_7027,N_6559,N_6494);
nor U7028 (N_7028,N_6790,N_6792);
or U7029 (N_7029,N_6742,N_6445);
and U7030 (N_7030,N_6782,N_6435);
or U7031 (N_7031,N_6564,N_6438);
or U7032 (N_7032,N_6542,N_6611);
nand U7033 (N_7033,N_6592,N_6744);
or U7034 (N_7034,N_6741,N_6758);
and U7035 (N_7035,N_6743,N_6438);
and U7036 (N_7036,N_6687,N_6545);
and U7037 (N_7037,N_6491,N_6677);
nor U7038 (N_7038,N_6592,N_6716);
nand U7039 (N_7039,N_6784,N_6432);
and U7040 (N_7040,N_6577,N_6417);
nor U7041 (N_7041,N_6711,N_6600);
or U7042 (N_7042,N_6727,N_6724);
or U7043 (N_7043,N_6522,N_6636);
nor U7044 (N_7044,N_6791,N_6704);
or U7045 (N_7045,N_6547,N_6439);
nand U7046 (N_7046,N_6729,N_6619);
nor U7047 (N_7047,N_6493,N_6474);
and U7048 (N_7048,N_6736,N_6421);
nor U7049 (N_7049,N_6759,N_6549);
nor U7050 (N_7050,N_6467,N_6592);
nand U7051 (N_7051,N_6678,N_6447);
nor U7052 (N_7052,N_6593,N_6403);
and U7053 (N_7053,N_6628,N_6738);
and U7054 (N_7054,N_6447,N_6636);
or U7055 (N_7055,N_6647,N_6748);
or U7056 (N_7056,N_6572,N_6639);
nand U7057 (N_7057,N_6616,N_6494);
nor U7058 (N_7058,N_6662,N_6780);
nor U7059 (N_7059,N_6462,N_6420);
nand U7060 (N_7060,N_6590,N_6475);
nand U7061 (N_7061,N_6557,N_6570);
and U7062 (N_7062,N_6718,N_6567);
and U7063 (N_7063,N_6696,N_6722);
nor U7064 (N_7064,N_6458,N_6476);
nor U7065 (N_7065,N_6462,N_6413);
and U7066 (N_7066,N_6622,N_6432);
and U7067 (N_7067,N_6712,N_6686);
and U7068 (N_7068,N_6771,N_6680);
and U7069 (N_7069,N_6722,N_6600);
nand U7070 (N_7070,N_6776,N_6473);
and U7071 (N_7071,N_6428,N_6569);
or U7072 (N_7072,N_6432,N_6437);
and U7073 (N_7073,N_6470,N_6485);
and U7074 (N_7074,N_6459,N_6435);
nand U7075 (N_7075,N_6472,N_6601);
nor U7076 (N_7076,N_6614,N_6747);
nand U7077 (N_7077,N_6497,N_6571);
nand U7078 (N_7078,N_6757,N_6751);
and U7079 (N_7079,N_6740,N_6626);
nor U7080 (N_7080,N_6551,N_6700);
nor U7081 (N_7081,N_6665,N_6408);
or U7082 (N_7082,N_6439,N_6621);
or U7083 (N_7083,N_6727,N_6634);
and U7084 (N_7084,N_6484,N_6494);
nand U7085 (N_7085,N_6745,N_6799);
nand U7086 (N_7086,N_6626,N_6468);
or U7087 (N_7087,N_6641,N_6444);
and U7088 (N_7088,N_6726,N_6472);
or U7089 (N_7089,N_6442,N_6752);
and U7090 (N_7090,N_6602,N_6778);
or U7091 (N_7091,N_6699,N_6563);
or U7092 (N_7092,N_6631,N_6682);
nand U7093 (N_7093,N_6551,N_6426);
and U7094 (N_7094,N_6656,N_6706);
nor U7095 (N_7095,N_6440,N_6620);
and U7096 (N_7096,N_6431,N_6636);
nor U7097 (N_7097,N_6504,N_6749);
nand U7098 (N_7098,N_6586,N_6463);
nor U7099 (N_7099,N_6542,N_6532);
nand U7100 (N_7100,N_6640,N_6553);
and U7101 (N_7101,N_6631,N_6577);
nand U7102 (N_7102,N_6599,N_6720);
nor U7103 (N_7103,N_6611,N_6779);
and U7104 (N_7104,N_6427,N_6461);
or U7105 (N_7105,N_6403,N_6662);
and U7106 (N_7106,N_6673,N_6560);
nor U7107 (N_7107,N_6758,N_6564);
nor U7108 (N_7108,N_6761,N_6445);
and U7109 (N_7109,N_6773,N_6487);
and U7110 (N_7110,N_6463,N_6649);
or U7111 (N_7111,N_6521,N_6584);
or U7112 (N_7112,N_6727,N_6766);
nand U7113 (N_7113,N_6579,N_6702);
and U7114 (N_7114,N_6691,N_6413);
nor U7115 (N_7115,N_6788,N_6670);
or U7116 (N_7116,N_6440,N_6715);
nor U7117 (N_7117,N_6704,N_6642);
and U7118 (N_7118,N_6650,N_6682);
nand U7119 (N_7119,N_6471,N_6636);
or U7120 (N_7120,N_6715,N_6552);
nor U7121 (N_7121,N_6480,N_6501);
nand U7122 (N_7122,N_6646,N_6758);
or U7123 (N_7123,N_6471,N_6702);
nor U7124 (N_7124,N_6527,N_6524);
or U7125 (N_7125,N_6549,N_6734);
and U7126 (N_7126,N_6458,N_6739);
and U7127 (N_7127,N_6696,N_6709);
or U7128 (N_7128,N_6453,N_6793);
or U7129 (N_7129,N_6718,N_6521);
and U7130 (N_7130,N_6434,N_6492);
and U7131 (N_7131,N_6434,N_6676);
nand U7132 (N_7132,N_6476,N_6682);
or U7133 (N_7133,N_6784,N_6495);
nand U7134 (N_7134,N_6722,N_6440);
and U7135 (N_7135,N_6622,N_6741);
or U7136 (N_7136,N_6504,N_6470);
nand U7137 (N_7137,N_6705,N_6494);
and U7138 (N_7138,N_6421,N_6472);
nand U7139 (N_7139,N_6624,N_6728);
nor U7140 (N_7140,N_6572,N_6433);
nor U7141 (N_7141,N_6650,N_6683);
and U7142 (N_7142,N_6552,N_6442);
nor U7143 (N_7143,N_6646,N_6418);
or U7144 (N_7144,N_6728,N_6436);
and U7145 (N_7145,N_6435,N_6794);
and U7146 (N_7146,N_6443,N_6732);
and U7147 (N_7147,N_6532,N_6628);
nand U7148 (N_7148,N_6487,N_6542);
nand U7149 (N_7149,N_6490,N_6469);
or U7150 (N_7150,N_6799,N_6727);
xor U7151 (N_7151,N_6678,N_6627);
nand U7152 (N_7152,N_6635,N_6524);
or U7153 (N_7153,N_6483,N_6798);
or U7154 (N_7154,N_6593,N_6793);
or U7155 (N_7155,N_6592,N_6410);
or U7156 (N_7156,N_6598,N_6404);
nand U7157 (N_7157,N_6779,N_6661);
nand U7158 (N_7158,N_6785,N_6549);
or U7159 (N_7159,N_6442,N_6663);
or U7160 (N_7160,N_6658,N_6730);
nor U7161 (N_7161,N_6745,N_6548);
and U7162 (N_7162,N_6696,N_6418);
nor U7163 (N_7163,N_6511,N_6707);
nor U7164 (N_7164,N_6476,N_6630);
nand U7165 (N_7165,N_6580,N_6496);
or U7166 (N_7166,N_6472,N_6466);
nand U7167 (N_7167,N_6479,N_6630);
nand U7168 (N_7168,N_6629,N_6712);
and U7169 (N_7169,N_6500,N_6779);
nand U7170 (N_7170,N_6658,N_6546);
and U7171 (N_7171,N_6518,N_6410);
or U7172 (N_7172,N_6527,N_6544);
nor U7173 (N_7173,N_6476,N_6430);
or U7174 (N_7174,N_6431,N_6637);
and U7175 (N_7175,N_6569,N_6461);
nor U7176 (N_7176,N_6783,N_6411);
nand U7177 (N_7177,N_6560,N_6452);
nand U7178 (N_7178,N_6658,N_6595);
or U7179 (N_7179,N_6711,N_6717);
and U7180 (N_7180,N_6492,N_6705);
and U7181 (N_7181,N_6523,N_6522);
nand U7182 (N_7182,N_6543,N_6478);
nor U7183 (N_7183,N_6532,N_6427);
and U7184 (N_7184,N_6593,N_6665);
or U7185 (N_7185,N_6735,N_6715);
nand U7186 (N_7186,N_6773,N_6593);
or U7187 (N_7187,N_6598,N_6650);
or U7188 (N_7188,N_6718,N_6765);
nand U7189 (N_7189,N_6437,N_6697);
nor U7190 (N_7190,N_6653,N_6547);
nand U7191 (N_7191,N_6471,N_6496);
nor U7192 (N_7192,N_6671,N_6593);
nor U7193 (N_7193,N_6756,N_6447);
and U7194 (N_7194,N_6468,N_6441);
nand U7195 (N_7195,N_6759,N_6681);
or U7196 (N_7196,N_6708,N_6451);
nand U7197 (N_7197,N_6682,N_6558);
or U7198 (N_7198,N_6496,N_6586);
or U7199 (N_7199,N_6491,N_6653);
or U7200 (N_7200,N_7107,N_7130);
and U7201 (N_7201,N_7142,N_7102);
and U7202 (N_7202,N_7149,N_6960);
nand U7203 (N_7203,N_6836,N_7194);
and U7204 (N_7204,N_7168,N_7068);
nor U7205 (N_7205,N_7025,N_7159);
nand U7206 (N_7206,N_6878,N_7059);
or U7207 (N_7207,N_6942,N_7166);
or U7208 (N_7208,N_7177,N_7139);
or U7209 (N_7209,N_7040,N_7011);
nand U7210 (N_7210,N_6818,N_6990);
nand U7211 (N_7211,N_7188,N_7113);
nor U7212 (N_7212,N_6957,N_6964);
and U7213 (N_7213,N_7002,N_7086);
nor U7214 (N_7214,N_7078,N_7193);
or U7215 (N_7215,N_7164,N_6808);
nand U7216 (N_7216,N_6930,N_6926);
and U7217 (N_7217,N_6999,N_6854);
nor U7218 (N_7218,N_6851,N_7010);
or U7219 (N_7219,N_6920,N_6868);
and U7220 (N_7220,N_7091,N_6865);
or U7221 (N_7221,N_6945,N_6955);
nor U7222 (N_7222,N_6988,N_7112);
and U7223 (N_7223,N_7156,N_7187);
or U7224 (N_7224,N_6992,N_6911);
nor U7225 (N_7225,N_6966,N_7079);
nor U7226 (N_7226,N_7101,N_7183);
or U7227 (N_7227,N_6863,N_6895);
nand U7228 (N_7228,N_7090,N_6912);
nand U7229 (N_7229,N_7172,N_6946);
or U7230 (N_7230,N_6838,N_7105);
and U7231 (N_7231,N_7152,N_6901);
nor U7232 (N_7232,N_7128,N_6963);
nand U7233 (N_7233,N_6903,N_6896);
nor U7234 (N_7234,N_7144,N_7004);
and U7235 (N_7235,N_6846,N_7046);
or U7236 (N_7236,N_7057,N_6932);
or U7237 (N_7237,N_6847,N_6884);
or U7238 (N_7238,N_6931,N_6914);
or U7239 (N_7239,N_7012,N_7154);
nor U7240 (N_7240,N_7135,N_6991);
nor U7241 (N_7241,N_6864,N_6977);
or U7242 (N_7242,N_6962,N_6909);
nand U7243 (N_7243,N_6858,N_7153);
and U7244 (N_7244,N_7071,N_6954);
or U7245 (N_7245,N_6804,N_7191);
or U7246 (N_7246,N_6828,N_6853);
nand U7247 (N_7247,N_6859,N_6915);
and U7248 (N_7248,N_6841,N_6885);
nor U7249 (N_7249,N_7176,N_6829);
and U7250 (N_7250,N_6902,N_7151);
or U7251 (N_7251,N_7036,N_7083);
nor U7252 (N_7252,N_6965,N_7018);
nand U7253 (N_7253,N_6972,N_7089);
and U7254 (N_7254,N_6917,N_6876);
or U7255 (N_7255,N_7048,N_6817);
nor U7256 (N_7256,N_6813,N_6950);
nand U7257 (N_7257,N_6934,N_6807);
nand U7258 (N_7258,N_7100,N_7127);
nor U7259 (N_7259,N_7087,N_7140);
or U7260 (N_7260,N_7131,N_7062);
nand U7261 (N_7261,N_6969,N_7126);
and U7262 (N_7262,N_6898,N_7008);
nand U7263 (N_7263,N_6834,N_6855);
nor U7264 (N_7264,N_7192,N_6810);
xor U7265 (N_7265,N_7095,N_7138);
and U7266 (N_7266,N_7019,N_7015);
and U7267 (N_7267,N_6971,N_7041);
xor U7268 (N_7268,N_7064,N_7109);
nor U7269 (N_7269,N_6979,N_6883);
or U7270 (N_7270,N_6982,N_6887);
nand U7271 (N_7271,N_6975,N_7161);
or U7272 (N_7272,N_7052,N_7022);
nor U7273 (N_7273,N_6837,N_6984);
or U7274 (N_7274,N_6918,N_6871);
nor U7275 (N_7275,N_6852,N_6822);
and U7276 (N_7276,N_7050,N_7180);
and U7277 (N_7277,N_6956,N_7070);
or U7278 (N_7278,N_7063,N_6893);
nor U7279 (N_7279,N_7077,N_7115);
nor U7280 (N_7280,N_7021,N_6815);
or U7281 (N_7281,N_6987,N_7124);
nor U7282 (N_7282,N_7125,N_6881);
or U7283 (N_7283,N_7199,N_6941);
nor U7284 (N_7284,N_7088,N_6897);
nand U7285 (N_7285,N_7158,N_7104);
nand U7286 (N_7286,N_6831,N_6940);
and U7287 (N_7287,N_7185,N_7175);
nand U7288 (N_7288,N_7076,N_6843);
or U7289 (N_7289,N_7157,N_6973);
nor U7290 (N_7290,N_6899,N_7000);
and U7291 (N_7291,N_6959,N_6900);
or U7292 (N_7292,N_6850,N_7134);
nor U7293 (N_7293,N_6840,N_6907);
or U7294 (N_7294,N_6839,N_7034);
nand U7295 (N_7295,N_6805,N_6921);
nor U7296 (N_7296,N_6905,N_7181);
xor U7297 (N_7297,N_6886,N_6939);
nor U7298 (N_7298,N_7098,N_7190);
and U7299 (N_7299,N_6821,N_6882);
nand U7300 (N_7300,N_7038,N_6970);
nand U7301 (N_7301,N_7005,N_6806);
or U7302 (N_7302,N_6812,N_7061);
nand U7303 (N_7303,N_6860,N_6943);
or U7304 (N_7304,N_7007,N_7137);
nor U7305 (N_7305,N_6922,N_6936);
nor U7306 (N_7306,N_7020,N_7055);
and U7307 (N_7307,N_6980,N_6978);
nor U7308 (N_7308,N_6873,N_7032);
or U7309 (N_7309,N_7106,N_7111);
and U7310 (N_7310,N_6874,N_7058);
nor U7311 (N_7311,N_6869,N_7043);
nor U7312 (N_7312,N_7155,N_7047);
xor U7313 (N_7313,N_6923,N_7119);
nand U7314 (N_7314,N_6870,N_7184);
nor U7315 (N_7315,N_6924,N_6862);
nand U7316 (N_7316,N_6995,N_7027);
and U7317 (N_7317,N_7121,N_7170);
and U7318 (N_7318,N_6832,N_6944);
or U7319 (N_7319,N_7035,N_7001);
or U7320 (N_7320,N_6996,N_7029);
and U7321 (N_7321,N_6927,N_7195);
nand U7322 (N_7322,N_7174,N_6997);
and U7323 (N_7323,N_7081,N_7065);
and U7324 (N_7324,N_7129,N_6830);
nand U7325 (N_7325,N_7147,N_6989);
nand U7326 (N_7326,N_7120,N_7053);
or U7327 (N_7327,N_7013,N_7044);
nand U7328 (N_7328,N_6949,N_7026);
nand U7329 (N_7329,N_6937,N_6872);
or U7330 (N_7330,N_6824,N_7073);
or U7331 (N_7331,N_6833,N_7072);
nor U7332 (N_7332,N_7096,N_6994);
nand U7333 (N_7333,N_6952,N_6848);
nand U7334 (N_7334,N_6906,N_7179);
nor U7335 (N_7335,N_7189,N_7094);
or U7336 (N_7336,N_6951,N_7082);
or U7337 (N_7337,N_7118,N_7162);
or U7338 (N_7338,N_7009,N_7103);
and U7339 (N_7339,N_7031,N_6875);
nand U7340 (N_7340,N_6826,N_6801);
and U7341 (N_7341,N_7030,N_6820);
and U7342 (N_7342,N_7092,N_6935);
nand U7343 (N_7343,N_6857,N_6919);
and U7344 (N_7344,N_7148,N_6967);
or U7345 (N_7345,N_7173,N_7037);
or U7346 (N_7346,N_6835,N_7171);
nor U7347 (N_7347,N_6986,N_6861);
or U7348 (N_7348,N_7028,N_6845);
nand U7349 (N_7349,N_7033,N_7136);
nor U7350 (N_7350,N_6948,N_7051);
nor U7351 (N_7351,N_7097,N_7075);
and U7352 (N_7352,N_7150,N_7146);
nor U7353 (N_7353,N_6856,N_7017);
nor U7354 (N_7354,N_7039,N_7123);
nand U7355 (N_7355,N_7169,N_7060);
nand U7356 (N_7356,N_7196,N_6889);
or U7357 (N_7357,N_6892,N_7074);
nor U7358 (N_7358,N_6803,N_7045);
nand U7359 (N_7359,N_6849,N_7014);
nand U7360 (N_7360,N_6933,N_6916);
and U7361 (N_7361,N_7067,N_7122);
nor U7362 (N_7362,N_6844,N_6974);
or U7363 (N_7363,N_7197,N_7049);
nand U7364 (N_7364,N_7056,N_6802);
and U7365 (N_7365,N_6866,N_7163);
nand U7366 (N_7366,N_7042,N_7080);
nand U7367 (N_7367,N_6814,N_6968);
nor U7368 (N_7368,N_7023,N_6880);
and U7369 (N_7369,N_7084,N_7132);
and U7370 (N_7370,N_7003,N_6925);
nor U7371 (N_7371,N_7069,N_7198);
or U7372 (N_7372,N_6928,N_7099);
nor U7373 (N_7373,N_6825,N_6993);
and U7374 (N_7374,N_6947,N_7117);
nor U7375 (N_7375,N_6800,N_6811);
and U7376 (N_7376,N_7178,N_7016);
or U7377 (N_7377,N_6867,N_6985);
or U7378 (N_7378,N_6842,N_7141);
or U7379 (N_7379,N_6809,N_6961);
nand U7380 (N_7380,N_7054,N_6910);
and U7381 (N_7381,N_6894,N_7133);
nand U7382 (N_7382,N_6890,N_6976);
and U7383 (N_7383,N_7093,N_6953);
or U7384 (N_7384,N_7165,N_7145);
nor U7385 (N_7385,N_7116,N_6913);
or U7386 (N_7386,N_7110,N_7066);
nand U7387 (N_7387,N_6998,N_7160);
and U7388 (N_7388,N_6958,N_6877);
nor U7389 (N_7389,N_6904,N_7024);
or U7390 (N_7390,N_6888,N_6823);
and U7391 (N_7391,N_6879,N_7182);
nand U7392 (N_7392,N_6983,N_6938);
nand U7393 (N_7393,N_7114,N_7108);
and U7394 (N_7394,N_7143,N_7167);
or U7395 (N_7395,N_6908,N_6891);
nor U7396 (N_7396,N_7085,N_6819);
or U7397 (N_7397,N_6816,N_6929);
or U7398 (N_7398,N_7006,N_6981);
and U7399 (N_7399,N_6827,N_7186);
nand U7400 (N_7400,N_7176,N_6838);
xor U7401 (N_7401,N_7107,N_7014);
and U7402 (N_7402,N_7129,N_6928);
or U7403 (N_7403,N_6874,N_7050);
nand U7404 (N_7404,N_6831,N_6933);
and U7405 (N_7405,N_7167,N_6891);
and U7406 (N_7406,N_6916,N_7044);
nand U7407 (N_7407,N_6847,N_7002);
or U7408 (N_7408,N_7013,N_7012);
nor U7409 (N_7409,N_6979,N_6937);
or U7410 (N_7410,N_6936,N_6811);
or U7411 (N_7411,N_6958,N_6860);
xnor U7412 (N_7412,N_6984,N_7135);
xor U7413 (N_7413,N_7086,N_6979);
nor U7414 (N_7414,N_6846,N_6863);
nand U7415 (N_7415,N_6821,N_6918);
xor U7416 (N_7416,N_6975,N_7198);
nand U7417 (N_7417,N_7137,N_6971);
and U7418 (N_7418,N_7094,N_6817);
and U7419 (N_7419,N_7091,N_6858);
nand U7420 (N_7420,N_7138,N_6977);
or U7421 (N_7421,N_7070,N_7170);
or U7422 (N_7422,N_6905,N_6868);
or U7423 (N_7423,N_7017,N_7048);
or U7424 (N_7424,N_7131,N_6951);
and U7425 (N_7425,N_6924,N_7002);
nor U7426 (N_7426,N_7022,N_6843);
and U7427 (N_7427,N_6927,N_6832);
nand U7428 (N_7428,N_6815,N_6894);
nand U7429 (N_7429,N_6905,N_7192);
nand U7430 (N_7430,N_6921,N_7126);
or U7431 (N_7431,N_6977,N_7129);
nor U7432 (N_7432,N_7199,N_7006);
nor U7433 (N_7433,N_6983,N_7076);
or U7434 (N_7434,N_7044,N_7014);
nor U7435 (N_7435,N_7088,N_6862);
and U7436 (N_7436,N_6836,N_7177);
or U7437 (N_7437,N_7157,N_6808);
nand U7438 (N_7438,N_7067,N_6899);
nor U7439 (N_7439,N_7170,N_6902);
and U7440 (N_7440,N_6820,N_7133);
nand U7441 (N_7441,N_6917,N_6862);
nand U7442 (N_7442,N_6806,N_7089);
and U7443 (N_7443,N_6960,N_7011);
nand U7444 (N_7444,N_7160,N_6885);
nor U7445 (N_7445,N_6833,N_6916);
nand U7446 (N_7446,N_6832,N_7119);
and U7447 (N_7447,N_7004,N_6820);
or U7448 (N_7448,N_6972,N_6877);
and U7449 (N_7449,N_6913,N_7020);
and U7450 (N_7450,N_7064,N_6950);
nand U7451 (N_7451,N_6863,N_6812);
nand U7452 (N_7452,N_6937,N_6814);
nand U7453 (N_7453,N_6864,N_7013);
nand U7454 (N_7454,N_7140,N_6954);
xor U7455 (N_7455,N_6864,N_6943);
nor U7456 (N_7456,N_6821,N_7106);
nand U7457 (N_7457,N_7177,N_7130);
or U7458 (N_7458,N_7097,N_7008);
and U7459 (N_7459,N_7098,N_6976);
or U7460 (N_7460,N_6801,N_6847);
nor U7461 (N_7461,N_6986,N_7141);
and U7462 (N_7462,N_7148,N_7137);
nand U7463 (N_7463,N_7135,N_6935);
or U7464 (N_7464,N_6807,N_7039);
nor U7465 (N_7465,N_7008,N_6850);
nand U7466 (N_7466,N_7157,N_6814);
nand U7467 (N_7467,N_7111,N_7010);
nor U7468 (N_7468,N_7110,N_7126);
nor U7469 (N_7469,N_7177,N_7182);
nor U7470 (N_7470,N_7153,N_6918);
or U7471 (N_7471,N_7056,N_6934);
nor U7472 (N_7472,N_6984,N_6970);
or U7473 (N_7473,N_6942,N_6854);
nor U7474 (N_7474,N_6892,N_7144);
and U7475 (N_7475,N_7168,N_6874);
nor U7476 (N_7476,N_7076,N_6824);
nand U7477 (N_7477,N_7171,N_7174);
nor U7478 (N_7478,N_7169,N_7139);
or U7479 (N_7479,N_7186,N_7017);
nor U7480 (N_7480,N_6905,N_7144);
and U7481 (N_7481,N_6924,N_7145);
nand U7482 (N_7482,N_6853,N_6927);
and U7483 (N_7483,N_7005,N_6882);
nand U7484 (N_7484,N_7054,N_7001);
and U7485 (N_7485,N_6837,N_6891);
nand U7486 (N_7486,N_7146,N_6987);
or U7487 (N_7487,N_7079,N_6974);
nor U7488 (N_7488,N_7194,N_7148);
nand U7489 (N_7489,N_7180,N_6911);
or U7490 (N_7490,N_7103,N_6844);
or U7491 (N_7491,N_6849,N_7090);
nand U7492 (N_7492,N_7136,N_6874);
and U7493 (N_7493,N_6880,N_6813);
or U7494 (N_7494,N_7162,N_6938);
or U7495 (N_7495,N_7117,N_7034);
or U7496 (N_7496,N_6843,N_7006);
and U7497 (N_7497,N_7100,N_7020);
and U7498 (N_7498,N_7001,N_6933);
or U7499 (N_7499,N_7188,N_7121);
or U7500 (N_7500,N_6914,N_6996);
nor U7501 (N_7501,N_6900,N_6836);
nand U7502 (N_7502,N_6894,N_6848);
nor U7503 (N_7503,N_6913,N_6874);
nand U7504 (N_7504,N_6908,N_7150);
nor U7505 (N_7505,N_7058,N_7179);
or U7506 (N_7506,N_6913,N_6802);
and U7507 (N_7507,N_6855,N_7192);
or U7508 (N_7508,N_6913,N_6976);
and U7509 (N_7509,N_7012,N_6940);
and U7510 (N_7510,N_7090,N_6835);
and U7511 (N_7511,N_6811,N_6864);
nand U7512 (N_7512,N_6945,N_7086);
or U7513 (N_7513,N_7012,N_6943);
nor U7514 (N_7514,N_6838,N_7050);
nor U7515 (N_7515,N_6898,N_6863);
and U7516 (N_7516,N_6904,N_7163);
nand U7517 (N_7517,N_7037,N_7078);
and U7518 (N_7518,N_7130,N_6927);
or U7519 (N_7519,N_6960,N_7109);
nor U7520 (N_7520,N_6837,N_7123);
and U7521 (N_7521,N_6939,N_7045);
nor U7522 (N_7522,N_6949,N_7093);
nand U7523 (N_7523,N_6805,N_6863);
nor U7524 (N_7524,N_6868,N_6831);
nor U7525 (N_7525,N_6959,N_6889);
or U7526 (N_7526,N_6864,N_6801);
and U7527 (N_7527,N_6954,N_7034);
and U7528 (N_7528,N_7130,N_6894);
or U7529 (N_7529,N_7155,N_6835);
nand U7530 (N_7530,N_7146,N_7065);
and U7531 (N_7531,N_6931,N_6980);
nor U7532 (N_7532,N_7088,N_6908);
nor U7533 (N_7533,N_6993,N_6890);
and U7534 (N_7534,N_7063,N_7062);
and U7535 (N_7535,N_6819,N_6922);
nand U7536 (N_7536,N_7194,N_6958);
and U7537 (N_7537,N_6900,N_7029);
and U7538 (N_7538,N_7097,N_7041);
and U7539 (N_7539,N_7008,N_7069);
nand U7540 (N_7540,N_7062,N_6950);
nor U7541 (N_7541,N_6858,N_7097);
nor U7542 (N_7542,N_7070,N_6969);
xor U7543 (N_7543,N_6978,N_6919);
nand U7544 (N_7544,N_6908,N_7032);
nand U7545 (N_7545,N_7152,N_6807);
nor U7546 (N_7546,N_6978,N_6972);
nand U7547 (N_7547,N_6811,N_6976);
and U7548 (N_7548,N_7104,N_6990);
nand U7549 (N_7549,N_7080,N_6856);
nand U7550 (N_7550,N_6857,N_7069);
and U7551 (N_7551,N_7073,N_7001);
nand U7552 (N_7552,N_7170,N_6802);
nor U7553 (N_7553,N_6905,N_7104);
and U7554 (N_7554,N_6928,N_7183);
nor U7555 (N_7555,N_6899,N_6820);
nor U7556 (N_7556,N_6856,N_6914);
and U7557 (N_7557,N_6964,N_6952);
nand U7558 (N_7558,N_6975,N_6957);
nand U7559 (N_7559,N_7165,N_6918);
or U7560 (N_7560,N_6804,N_7066);
nor U7561 (N_7561,N_6918,N_7053);
xnor U7562 (N_7562,N_7050,N_6963);
nor U7563 (N_7563,N_7045,N_6935);
or U7564 (N_7564,N_6940,N_6885);
and U7565 (N_7565,N_7159,N_6804);
nand U7566 (N_7566,N_7012,N_6878);
nand U7567 (N_7567,N_7138,N_7114);
or U7568 (N_7568,N_6996,N_7185);
nand U7569 (N_7569,N_6869,N_6837);
or U7570 (N_7570,N_6918,N_7125);
nand U7571 (N_7571,N_7152,N_6984);
and U7572 (N_7572,N_6835,N_7055);
and U7573 (N_7573,N_7124,N_7005);
and U7574 (N_7574,N_6839,N_6895);
and U7575 (N_7575,N_7099,N_7096);
and U7576 (N_7576,N_7078,N_7176);
and U7577 (N_7577,N_6885,N_6913);
and U7578 (N_7578,N_6860,N_6836);
and U7579 (N_7579,N_6800,N_6924);
nor U7580 (N_7580,N_6917,N_7097);
nand U7581 (N_7581,N_6888,N_7153);
and U7582 (N_7582,N_7114,N_7056);
or U7583 (N_7583,N_7081,N_7019);
and U7584 (N_7584,N_7134,N_6926);
nor U7585 (N_7585,N_7015,N_7001);
or U7586 (N_7586,N_6960,N_6912);
nand U7587 (N_7587,N_7117,N_6904);
nor U7588 (N_7588,N_6994,N_7167);
nor U7589 (N_7589,N_7143,N_7046);
nand U7590 (N_7590,N_7006,N_6966);
nor U7591 (N_7591,N_6909,N_7054);
nand U7592 (N_7592,N_6844,N_7086);
nand U7593 (N_7593,N_7189,N_7025);
and U7594 (N_7594,N_7143,N_7080);
nand U7595 (N_7595,N_6807,N_6845);
and U7596 (N_7596,N_7050,N_7097);
nor U7597 (N_7597,N_7182,N_6894);
nor U7598 (N_7598,N_7173,N_7000);
nand U7599 (N_7599,N_6828,N_6872);
nor U7600 (N_7600,N_7419,N_7331);
or U7601 (N_7601,N_7411,N_7350);
nor U7602 (N_7602,N_7562,N_7508);
and U7603 (N_7603,N_7263,N_7208);
and U7604 (N_7604,N_7438,N_7403);
nor U7605 (N_7605,N_7566,N_7270);
nor U7606 (N_7606,N_7353,N_7576);
nand U7607 (N_7607,N_7445,N_7288);
and U7608 (N_7608,N_7559,N_7256);
nand U7609 (N_7609,N_7429,N_7289);
nor U7610 (N_7610,N_7332,N_7565);
nor U7611 (N_7611,N_7236,N_7540);
and U7612 (N_7612,N_7390,N_7202);
nand U7613 (N_7613,N_7221,N_7587);
nand U7614 (N_7614,N_7447,N_7328);
nand U7615 (N_7615,N_7364,N_7584);
nor U7616 (N_7616,N_7423,N_7317);
nor U7617 (N_7617,N_7502,N_7303);
nand U7618 (N_7618,N_7501,N_7491);
and U7619 (N_7619,N_7254,N_7389);
and U7620 (N_7620,N_7302,N_7301);
and U7621 (N_7621,N_7467,N_7518);
nor U7622 (N_7622,N_7228,N_7441);
or U7623 (N_7623,N_7510,N_7235);
and U7624 (N_7624,N_7568,N_7500);
nor U7625 (N_7625,N_7229,N_7227);
and U7626 (N_7626,N_7570,N_7539);
nand U7627 (N_7627,N_7422,N_7201);
or U7628 (N_7628,N_7347,N_7535);
and U7629 (N_7629,N_7489,N_7431);
and U7630 (N_7630,N_7581,N_7203);
nand U7631 (N_7631,N_7346,N_7395);
and U7632 (N_7632,N_7291,N_7385);
or U7633 (N_7633,N_7307,N_7554);
and U7634 (N_7634,N_7567,N_7529);
and U7635 (N_7635,N_7585,N_7264);
and U7636 (N_7636,N_7433,N_7564);
nand U7637 (N_7637,N_7583,N_7267);
or U7638 (N_7638,N_7448,N_7382);
nor U7639 (N_7639,N_7355,N_7246);
nor U7640 (N_7640,N_7375,N_7416);
or U7641 (N_7641,N_7504,N_7394);
nor U7642 (N_7642,N_7315,N_7408);
nand U7643 (N_7643,N_7524,N_7522);
nor U7644 (N_7644,N_7440,N_7473);
nand U7645 (N_7645,N_7420,N_7401);
or U7646 (N_7646,N_7404,N_7297);
nor U7647 (N_7647,N_7439,N_7250);
and U7648 (N_7648,N_7470,N_7362);
nand U7649 (N_7649,N_7245,N_7294);
or U7650 (N_7650,N_7369,N_7262);
or U7651 (N_7651,N_7455,N_7471);
nand U7652 (N_7652,N_7387,N_7333);
nand U7653 (N_7653,N_7209,N_7573);
nand U7654 (N_7654,N_7240,N_7225);
and U7655 (N_7655,N_7530,N_7571);
nor U7656 (N_7656,N_7378,N_7357);
or U7657 (N_7657,N_7280,N_7271);
nand U7658 (N_7658,N_7223,N_7268);
and U7659 (N_7659,N_7278,N_7233);
nor U7660 (N_7660,N_7205,N_7552);
or U7661 (N_7661,N_7457,N_7374);
or U7662 (N_7662,N_7586,N_7244);
nand U7663 (N_7663,N_7406,N_7373);
nor U7664 (N_7664,N_7360,N_7476);
nand U7665 (N_7665,N_7396,N_7546);
and U7666 (N_7666,N_7442,N_7452);
and U7667 (N_7667,N_7300,N_7204);
and U7668 (N_7668,N_7596,N_7239);
and U7669 (N_7669,N_7407,N_7511);
or U7670 (N_7670,N_7388,N_7451);
or U7671 (N_7671,N_7252,N_7575);
or U7672 (N_7672,N_7437,N_7480);
nor U7673 (N_7673,N_7287,N_7474);
or U7674 (N_7674,N_7578,N_7509);
and U7675 (N_7675,N_7277,N_7290);
and U7676 (N_7676,N_7323,N_7220);
and U7677 (N_7677,N_7496,N_7541);
nor U7678 (N_7678,N_7409,N_7495);
and U7679 (N_7679,N_7354,N_7479);
nand U7680 (N_7680,N_7545,N_7515);
nor U7681 (N_7681,N_7349,N_7417);
or U7682 (N_7682,N_7595,N_7593);
or U7683 (N_7683,N_7563,N_7306);
nand U7684 (N_7684,N_7241,N_7557);
nor U7685 (N_7685,N_7370,N_7391);
and U7686 (N_7686,N_7402,N_7215);
nand U7687 (N_7687,N_7547,N_7230);
nand U7688 (N_7688,N_7218,N_7327);
nand U7689 (N_7689,N_7342,N_7363);
or U7690 (N_7690,N_7550,N_7248);
or U7691 (N_7691,N_7274,N_7324);
or U7692 (N_7692,N_7326,N_7210);
nand U7693 (N_7693,N_7365,N_7341);
and U7694 (N_7694,N_7525,N_7200);
nand U7695 (N_7695,N_7213,N_7386);
and U7696 (N_7696,N_7499,N_7591);
nand U7697 (N_7697,N_7466,N_7296);
nor U7698 (N_7698,N_7206,N_7392);
or U7699 (N_7699,N_7358,N_7492);
nor U7700 (N_7700,N_7582,N_7275);
or U7701 (N_7701,N_7519,N_7597);
nand U7702 (N_7702,N_7222,N_7465);
or U7703 (N_7703,N_7232,N_7536);
nor U7704 (N_7704,N_7361,N_7265);
or U7705 (N_7705,N_7310,N_7325);
or U7706 (N_7706,N_7531,N_7444);
or U7707 (N_7707,N_7574,N_7432);
and U7708 (N_7708,N_7381,N_7322);
nand U7709 (N_7709,N_7488,N_7556);
or U7710 (N_7710,N_7285,N_7376);
nand U7711 (N_7711,N_7456,N_7526);
nor U7712 (N_7712,N_7311,N_7397);
or U7713 (N_7713,N_7249,N_7588);
nor U7714 (N_7714,N_7283,N_7458);
and U7715 (N_7715,N_7366,N_7478);
and U7716 (N_7716,N_7295,N_7413);
nor U7717 (N_7717,N_7352,N_7405);
or U7718 (N_7718,N_7255,N_7421);
nand U7719 (N_7719,N_7207,N_7534);
or U7720 (N_7720,N_7313,N_7312);
nor U7721 (N_7721,N_7334,N_7462);
or U7722 (N_7722,N_7292,N_7279);
or U7723 (N_7723,N_7314,N_7453);
or U7724 (N_7724,N_7548,N_7538);
and U7725 (N_7725,N_7266,N_7475);
and U7726 (N_7726,N_7211,N_7594);
nor U7727 (N_7727,N_7592,N_7212);
nand U7728 (N_7728,N_7286,N_7468);
and U7729 (N_7729,N_7503,N_7482);
nand U7730 (N_7730,N_7304,N_7494);
nor U7731 (N_7731,N_7426,N_7486);
nor U7732 (N_7732,N_7549,N_7464);
or U7733 (N_7733,N_7259,N_7589);
or U7734 (N_7734,N_7537,N_7398);
and U7735 (N_7735,N_7418,N_7553);
and U7736 (N_7736,N_7414,N_7393);
and U7737 (N_7737,N_7425,N_7598);
and U7738 (N_7738,N_7521,N_7226);
and U7739 (N_7739,N_7412,N_7400);
and U7740 (N_7740,N_7590,N_7399);
nand U7741 (N_7741,N_7558,N_7371);
nand U7742 (N_7742,N_7384,N_7430);
or U7743 (N_7743,N_7542,N_7377);
nand U7744 (N_7744,N_7513,N_7336);
nand U7745 (N_7745,N_7348,N_7356);
nor U7746 (N_7746,N_7528,N_7351);
nand U7747 (N_7747,N_7368,N_7450);
and U7748 (N_7748,N_7216,N_7320);
and U7749 (N_7749,N_7238,N_7309);
or U7750 (N_7750,N_7293,N_7298);
or U7751 (N_7751,N_7551,N_7497);
nor U7752 (N_7752,N_7446,N_7517);
nor U7753 (N_7753,N_7579,N_7247);
nand U7754 (N_7754,N_7380,N_7485);
nor U7755 (N_7755,N_7454,N_7459);
nand U7756 (N_7756,N_7506,N_7477);
nand U7757 (N_7757,N_7507,N_7316);
nand U7758 (N_7758,N_7415,N_7514);
or U7759 (N_7759,N_7276,N_7428);
nor U7760 (N_7760,N_7577,N_7214);
or U7761 (N_7761,N_7367,N_7481);
and U7762 (N_7762,N_7435,N_7580);
nor U7763 (N_7763,N_7234,N_7305);
and U7764 (N_7764,N_7318,N_7273);
or U7765 (N_7765,N_7449,N_7231);
nor U7766 (N_7766,N_7560,N_7572);
nand U7767 (N_7767,N_7261,N_7484);
and U7768 (N_7768,N_7527,N_7308);
nand U7769 (N_7769,N_7561,N_7461);
or U7770 (N_7770,N_7490,N_7512);
or U7771 (N_7771,N_7463,N_7344);
and U7772 (N_7772,N_7434,N_7487);
and U7773 (N_7773,N_7257,N_7284);
or U7774 (N_7774,N_7253,N_7219);
or U7775 (N_7775,N_7330,N_7321);
nand U7776 (N_7776,N_7282,N_7343);
and U7777 (N_7777,N_7505,N_7543);
nor U7778 (N_7778,N_7469,N_7443);
and U7779 (N_7779,N_7243,N_7383);
or U7780 (N_7780,N_7345,N_7340);
and U7781 (N_7781,N_7272,N_7460);
nor U7782 (N_7782,N_7258,N_7217);
and U7783 (N_7783,N_7555,N_7427);
nand U7784 (N_7784,N_7319,N_7224);
nand U7785 (N_7785,N_7493,N_7242);
or U7786 (N_7786,N_7237,N_7338);
or U7787 (N_7787,N_7329,N_7483);
or U7788 (N_7788,N_7569,N_7532);
or U7789 (N_7789,N_7372,N_7523);
nor U7790 (N_7790,N_7516,N_7337);
and U7791 (N_7791,N_7520,N_7260);
nand U7792 (N_7792,N_7424,N_7379);
nand U7793 (N_7793,N_7335,N_7339);
nand U7794 (N_7794,N_7436,N_7359);
and U7795 (N_7795,N_7533,N_7498);
and U7796 (N_7796,N_7472,N_7281);
and U7797 (N_7797,N_7299,N_7251);
nand U7798 (N_7798,N_7410,N_7599);
and U7799 (N_7799,N_7544,N_7269);
or U7800 (N_7800,N_7513,N_7542);
or U7801 (N_7801,N_7494,N_7586);
nor U7802 (N_7802,N_7277,N_7242);
and U7803 (N_7803,N_7210,N_7241);
nor U7804 (N_7804,N_7428,N_7304);
or U7805 (N_7805,N_7358,N_7474);
nor U7806 (N_7806,N_7322,N_7215);
nand U7807 (N_7807,N_7254,N_7266);
nor U7808 (N_7808,N_7535,N_7240);
nor U7809 (N_7809,N_7572,N_7372);
nor U7810 (N_7810,N_7253,N_7307);
nor U7811 (N_7811,N_7369,N_7537);
nor U7812 (N_7812,N_7452,N_7470);
or U7813 (N_7813,N_7488,N_7422);
or U7814 (N_7814,N_7232,N_7560);
nor U7815 (N_7815,N_7559,N_7276);
nand U7816 (N_7816,N_7231,N_7228);
nand U7817 (N_7817,N_7294,N_7285);
nor U7818 (N_7818,N_7207,N_7486);
nor U7819 (N_7819,N_7530,N_7412);
nor U7820 (N_7820,N_7320,N_7572);
or U7821 (N_7821,N_7483,N_7538);
or U7822 (N_7822,N_7271,N_7410);
nand U7823 (N_7823,N_7217,N_7453);
and U7824 (N_7824,N_7401,N_7332);
nand U7825 (N_7825,N_7411,N_7546);
and U7826 (N_7826,N_7564,N_7332);
nand U7827 (N_7827,N_7348,N_7246);
and U7828 (N_7828,N_7405,N_7418);
nor U7829 (N_7829,N_7267,N_7352);
and U7830 (N_7830,N_7519,N_7323);
nor U7831 (N_7831,N_7236,N_7561);
and U7832 (N_7832,N_7235,N_7582);
or U7833 (N_7833,N_7528,N_7593);
nor U7834 (N_7834,N_7504,N_7467);
nand U7835 (N_7835,N_7464,N_7216);
or U7836 (N_7836,N_7298,N_7212);
nand U7837 (N_7837,N_7331,N_7581);
and U7838 (N_7838,N_7230,N_7228);
or U7839 (N_7839,N_7353,N_7224);
and U7840 (N_7840,N_7524,N_7560);
nand U7841 (N_7841,N_7437,N_7435);
or U7842 (N_7842,N_7244,N_7465);
or U7843 (N_7843,N_7404,N_7571);
nor U7844 (N_7844,N_7533,N_7532);
nand U7845 (N_7845,N_7509,N_7280);
or U7846 (N_7846,N_7385,N_7532);
nand U7847 (N_7847,N_7431,N_7425);
nand U7848 (N_7848,N_7577,N_7490);
or U7849 (N_7849,N_7412,N_7480);
and U7850 (N_7850,N_7282,N_7459);
or U7851 (N_7851,N_7353,N_7434);
nor U7852 (N_7852,N_7472,N_7371);
nand U7853 (N_7853,N_7218,N_7467);
or U7854 (N_7854,N_7536,N_7244);
nand U7855 (N_7855,N_7594,N_7337);
nor U7856 (N_7856,N_7411,N_7306);
and U7857 (N_7857,N_7551,N_7493);
nand U7858 (N_7858,N_7218,N_7256);
and U7859 (N_7859,N_7542,N_7281);
and U7860 (N_7860,N_7229,N_7595);
nand U7861 (N_7861,N_7530,N_7346);
or U7862 (N_7862,N_7503,N_7350);
nand U7863 (N_7863,N_7593,N_7442);
nor U7864 (N_7864,N_7546,N_7514);
nor U7865 (N_7865,N_7376,N_7565);
nor U7866 (N_7866,N_7462,N_7401);
nand U7867 (N_7867,N_7375,N_7246);
or U7868 (N_7868,N_7210,N_7282);
and U7869 (N_7869,N_7423,N_7237);
or U7870 (N_7870,N_7342,N_7402);
nor U7871 (N_7871,N_7307,N_7581);
or U7872 (N_7872,N_7399,N_7221);
or U7873 (N_7873,N_7477,N_7219);
nand U7874 (N_7874,N_7253,N_7519);
nand U7875 (N_7875,N_7549,N_7523);
and U7876 (N_7876,N_7480,N_7221);
and U7877 (N_7877,N_7296,N_7257);
and U7878 (N_7878,N_7456,N_7341);
nand U7879 (N_7879,N_7452,N_7255);
nor U7880 (N_7880,N_7477,N_7355);
nor U7881 (N_7881,N_7205,N_7219);
or U7882 (N_7882,N_7545,N_7220);
nor U7883 (N_7883,N_7449,N_7216);
nor U7884 (N_7884,N_7394,N_7570);
nor U7885 (N_7885,N_7532,N_7425);
or U7886 (N_7886,N_7234,N_7512);
nand U7887 (N_7887,N_7582,N_7229);
nor U7888 (N_7888,N_7220,N_7286);
nor U7889 (N_7889,N_7445,N_7483);
nand U7890 (N_7890,N_7330,N_7217);
nor U7891 (N_7891,N_7431,N_7339);
nand U7892 (N_7892,N_7384,N_7582);
and U7893 (N_7893,N_7380,N_7469);
and U7894 (N_7894,N_7379,N_7429);
and U7895 (N_7895,N_7288,N_7369);
nand U7896 (N_7896,N_7528,N_7589);
or U7897 (N_7897,N_7474,N_7249);
nand U7898 (N_7898,N_7513,N_7439);
or U7899 (N_7899,N_7256,N_7262);
and U7900 (N_7900,N_7380,N_7409);
and U7901 (N_7901,N_7501,N_7226);
nor U7902 (N_7902,N_7376,N_7576);
nor U7903 (N_7903,N_7339,N_7241);
nand U7904 (N_7904,N_7339,N_7451);
or U7905 (N_7905,N_7368,N_7292);
nand U7906 (N_7906,N_7257,N_7573);
or U7907 (N_7907,N_7518,N_7421);
nor U7908 (N_7908,N_7348,N_7595);
or U7909 (N_7909,N_7262,N_7248);
nand U7910 (N_7910,N_7474,N_7536);
and U7911 (N_7911,N_7445,N_7434);
or U7912 (N_7912,N_7324,N_7471);
nand U7913 (N_7913,N_7291,N_7567);
and U7914 (N_7914,N_7253,N_7487);
and U7915 (N_7915,N_7352,N_7266);
or U7916 (N_7916,N_7207,N_7219);
nand U7917 (N_7917,N_7432,N_7414);
or U7918 (N_7918,N_7448,N_7519);
nand U7919 (N_7919,N_7398,N_7494);
nor U7920 (N_7920,N_7281,N_7509);
nor U7921 (N_7921,N_7398,N_7578);
and U7922 (N_7922,N_7512,N_7404);
nor U7923 (N_7923,N_7572,N_7422);
nand U7924 (N_7924,N_7298,N_7486);
nor U7925 (N_7925,N_7564,N_7343);
or U7926 (N_7926,N_7586,N_7247);
or U7927 (N_7927,N_7379,N_7203);
or U7928 (N_7928,N_7326,N_7357);
xor U7929 (N_7929,N_7254,N_7355);
and U7930 (N_7930,N_7552,N_7510);
nand U7931 (N_7931,N_7435,N_7318);
or U7932 (N_7932,N_7563,N_7426);
nand U7933 (N_7933,N_7560,N_7266);
or U7934 (N_7934,N_7317,N_7375);
nand U7935 (N_7935,N_7379,N_7286);
and U7936 (N_7936,N_7481,N_7493);
and U7937 (N_7937,N_7512,N_7555);
nand U7938 (N_7938,N_7502,N_7553);
or U7939 (N_7939,N_7334,N_7449);
nor U7940 (N_7940,N_7445,N_7262);
or U7941 (N_7941,N_7371,N_7551);
nand U7942 (N_7942,N_7521,N_7263);
nand U7943 (N_7943,N_7508,N_7396);
and U7944 (N_7944,N_7440,N_7284);
xor U7945 (N_7945,N_7214,N_7509);
or U7946 (N_7946,N_7213,N_7295);
nand U7947 (N_7947,N_7491,N_7473);
nor U7948 (N_7948,N_7400,N_7212);
or U7949 (N_7949,N_7535,N_7490);
nor U7950 (N_7950,N_7546,N_7452);
and U7951 (N_7951,N_7405,N_7401);
nand U7952 (N_7952,N_7499,N_7434);
or U7953 (N_7953,N_7235,N_7229);
nor U7954 (N_7954,N_7224,N_7368);
or U7955 (N_7955,N_7254,N_7486);
nor U7956 (N_7956,N_7569,N_7323);
nand U7957 (N_7957,N_7505,N_7382);
nand U7958 (N_7958,N_7470,N_7279);
or U7959 (N_7959,N_7472,N_7246);
and U7960 (N_7960,N_7557,N_7215);
nand U7961 (N_7961,N_7533,N_7244);
nand U7962 (N_7962,N_7434,N_7519);
or U7963 (N_7963,N_7388,N_7314);
and U7964 (N_7964,N_7377,N_7464);
and U7965 (N_7965,N_7212,N_7425);
or U7966 (N_7966,N_7287,N_7408);
nor U7967 (N_7967,N_7532,N_7244);
nand U7968 (N_7968,N_7509,N_7299);
and U7969 (N_7969,N_7224,N_7424);
and U7970 (N_7970,N_7505,N_7287);
or U7971 (N_7971,N_7411,N_7447);
nor U7972 (N_7972,N_7494,N_7238);
or U7973 (N_7973,N_7338,N_7450);
and U7974 (N_7974,N_7512,N_7380);
nor U7975 (N_7975,N_7382,N_7327);
nand U7976 (N_7976,N_7596,N_7420);
nor U7977 (N_7977,N_7212,N_7524);
or U7978 (N_7978,N_7276,N_7521);
and U7979 (N_7979,N_7260,N_7592);
or U7980 (N_7980,N_7423,N_7477);
nand U7981 (N_7981,N_7400,N_7479);
or U7982 (N_7982,N_7465,N_7218);
and U7983 (N_7983,N_7523,N_7457);
nor U7984 (N_7984,N_7448,N_7566);
or U7985 (N_7985,N_7378,N_7313);
or U7986 (N_7986,N_7245,N_7569);
nand U7987 (N_7987,N_7410,N_7588);
and U7988 (N_7988,N_7428,N_7448);
nor U7989 (N_7989,N_7431,N_7565);
nand U7990 (N_7990,N_7235,N_7416);
and U7991 (N_7991,N_7586,N_7356);
nand U7992 (N_7992,N_7459,N_7313);
xor U7993 (N_7993,N_7358,N_7250);
nand U7994 (N_7994,N_7499,N_7253);
nor U7995 (N_7995,N_7269,N_7531);
or U7996 (N_7996,N_7215,N_7471);
nor U7997 (N_7997,N_7388,N_7581);
nor U7998 (N_7998,N_7577,N_7516);
and U7999 (N_7999,N_7399,N_7294);
nand U8000 (N_8000,N_7942,N_7772);
and U8001 (N_8001,N_7924,N_7793);
or U8002 (N_8002,N_7652,N_7969);
or U8003 (N_8003,N_7918,N_7648);
nand U8004 (N_8004,N_7619,N_7862);
and U8005 (N_8005,N_7878,N_7814);
and U8006 (N_8006,N_7792,N_7769);
xor U8007 (N_8007,N_7638,N_7857);
nand U8008 (N_8008,N_7828,N_7940);
nand U8009 (N_8009,N_7995,N_7982);
or U8010 (N_8010,N_7600,N_7958);
and U8011 (N_8011,N_7836,N_7926);
or U8012 (N_8012,N_7865,N_7839);
nand U8013 (N_8013,N_7740,N_7938);
nor U8014 (N_8014,N_7985,N_7650);
nor U8015 (N_8015,N_7907,N_7894);
and U8016 (N_8016,N_7722,N_7917);
and U8017 (N_8017,N_7800,N_7873);
and U8018 (N_8018,N_7645,N_7935);
nand U8019 (N_8019,N_7758,N_7630);
xnor U8020 (N_8020,N_7668,N_7887);
or U8021 (N_8021,N_7923,N_7734);
nand U8022 (N_8022,N_7892,N_7877);
or U8023 (N_8023,N_7978,N_7714);
nor U8024 (N_8024,N_7971,N_7750);
nand U8025 (N_8025,N_7846,N_7962);
and U8026 (N_8026,N_7756,N_7884);
or U8027 (N_8027,N_7929,N_7941);
nand U8028 (N_8028,N_7915,N_7670);
or U8029 (N_8029,N_7869,N_7897);
and U8030 (N_8030,N_7854,N_7972);
xnor U8031 (N_8031,N_7933,N_7678);
nor U8032 (N_8032,N_7711,N_7739);
nand U8033 (N_8033,N_7890,N_7781);
and U8034 (N_8034,N_7888,N_7639);
nor U8035 (N_8035,N_7623,N_7899);
xnor U8036 (N_8036,N_7851,N_7720);
and U8037 (N_8037,N_7980,N_7767);
nor U8038 (N_8038,N_7687,N_7715);
nor U8039 (N_8039,N_7761,N_7868);
and U8040 (N_8040,N_7747,N_7984);
nor U8041 (N_8041,N_7805,N_7817);
nand U8042 (N_8042,N_7610,N_7647);
and U8043 (N_8043,N_7803,N_7948);
or U8044 (N_8044,N_7694,N_7603);
nand U8045 (N_8045,N_7932,N_7867);
nor U8046 (N_8046,N_7795,N_7755);
and U8047 (N_8047,N_7601,N_7724);
nand U8048 (N_8048,N_7957,N_7961);
and U8049 (N_8049,N_7659,N_7880);
and U8050 (N_8050,N_7680,N_7927);
and U8051 (N_8051,N_7859,N_7777);
or U8052 (N_8052,N_7665,N_7766);
or U8053 (N_8053,N_7901,N_7611);
or U8054 (N_8054,N_7733,N_7841);
or U8055 (N_8055,N_7872,N_7970);
and U8056 (N_8056,N_7742,N_7672);
and U8057 (N_8057,N_7626,N_7625);
nor U8058 (N_8058,N_7629,N_7912);
and U8059 (N_8059,N_7864,N_7685);
and U8060 (N_8060,N_7621,N_7796);
nor U8061 (N_8061,N_7847,N_7667);
and U8062 (N_8062,N_7661,N_7662);
nor U8063 (N_8063,N_7820,N_7891);
or U8064 (N_8064,N_7736,N_7956);
nor U8065 (N_8065,N_7908,N_7807);
and U8066 (N_8066,N_7968,N_7690);
or U8067 (N_8067,N_7752,N_7748);
and U8068 (N_8068,N_7641,N_7987);
or U8069 (N_8069,N_7951,N_7993);
or U8070 (N_8070,N_7698,N_7785);
nor U8071 (N_8071,N_7997,N_7673);
nor U8072 (N_8072,N_7804,N_7778);
or U8073 (N_8073,N_7963,N_7966);
nor U8074 (N_8074,N_7773,N_7605);
nand U8075 (N_8075,N_7677,N_7770);
nor U8076 (N_8076,N_7823,N_7949);
nor U8077 (N_8077,N_7906,N_7879);
nand U8078 (N_8078,N_7719,N_7848);
nor U8079 (N_8079,N_7954,N_7620);
nand U8080 (N_8080,N_7794,N_7693);
nor U8081 (N_8081,N_7689,N_7920);
nand U8082 (N_8082,N_7635,N_7824);
or U8083 (N_8083,N_7764,N_7644);
nor U8084 (N_8084,N_7708,N_7754);
or U8085 (N_8085,N_7835,N_7905);
and U8086 (N_8086,N_7822,N_7808);
and U8087 (N_8087,N_7717,N_7910);
or U8088 (N_8088,N_7759,N_7886);
and U8089 (N_8089,N_7612,N_7992);
nand U8090 (N_8090,N_7973,N_7922);
nand U8091 (N_8091,N_7660,N_7852);
nor U8092 (N_8092,N_7840,N_7947);
or U8093 (N_8093,N_7723,N_7919);
nand U8094 (N_8094,N_7831,N_7893);
or U8095 (N_8095,N_7815,N_7700);
nand U8096 (N_8096,N_7735,N_7729);
nand U8097 (N_8097,N_7850,N_7682);
and U8098 (N_8098,N_7704,N_7943);
nor U8099 (N_8099,N_7651,N_7990);
and U8100 (N_8100,N_7712,N_7885);
nor U8101 (N_8101,N_7640,N_7676);
nor U8102 (N_8102,N_7701,N_7959);
or U8103 (N_8103,N_7911,N_7743);
nand U8104 (N_8104,N_7686,N_7881);
and U8105 (N_8105,N_7654,N_7692);
nor U8106 (N_8106,N_7696,N_7697);
nor U8107 (N_8107,N_7809,N_7679);
nor U8108 (N_8108,N_7979,N_7856);
or U8109 (N_8109,N_7633,N_7751);
nand U8110 (N_8110,N_7928,N_7707);
or U8111 (N_8111,N_7806,N_7898);
nor U8112 (N_8112,N_7783,N_7937);
or U8113 (N_8113,N_7730,N_7861);
nor U8114 (N_8114,N_7691,N_7606);
nand U8115 (N_8115,N_7613,N_7904);
nor U8116 (N_8116,N_7797,N_7858);
nand U8117 (N_8117,N_7607,N_7774);
and U8118 (N_8118,N_7802,N_7882);
and U8119 (N_8119,N_7812,N_7965);
and U8120 (N_8120,N_7991,N_7934);
nor U8121 (N_8121,N_7632,N_7616);
or U8122 (N_8122,N_7779,N_7731);
nand U8123 (N_8123,N_7983,N_7709);
nand U8124 (N_8124,N_7986,N_7614);
or U8125 (N_8125,N_7728,N_7666);
nor U8126 (N_8126,N_7914,N_7870);
and U8127 (N_8127,N_7830,N_7790);
nor U8128 (N_8128,N_7875,N_7843);
nand U8129 (N_8129,N_7964,N_7902);
and U8130 (N_8130,N_7953,N_7945);
nor U8131 (N_8131,N_7624,N_7604);
and U8132 (N_8132,N_7950,N_7627);
and U8133 (N_8133,N_7936,N_7727);
and U8134 (N_8134,N_7646,N_7798);
and U8135 (N_8135,N_7998,N_7816);
nor U8136 (N_8136,N_7713,N_7845);
or U8137 (N_8137,N_7977,N_7810);
nand U8138 (N_8138,N_7702,N_7976);
nor U8139 (N_8139,N_7669,N_7746);
or U8140 (N_8140,N_7771,N_7732);
nor U8141 (N_8141,N_7921,N_7671);
nand U8142 (N_8142,N_7784,N_7716);
or U8143 (N_8143,N_7726,N_7819);
nor U8144 (N_8144,N_7721,N_7749);
nor U8145 (N_8145,N_7674,N_7705);
nand U8146 (N_8146,N_7788,N_7622);
and U8147 (N_8147,N_7744,N_7786);
nand U8148 (N_8148,N_7725,N_7653);
and U8149 (N_8149,N_7903,N_7710);
and U8150 (N_8150,N_7813,N_7683);
nand U8151 (N_8151,N_7706,N_7900);
or U8152 (N_8152,N_7913,N_7849);
nand U8153 (N_8153,N_7826,N_7791);
and U8154 (N_8154,N_7829,N_7999);
and U8155 (N_8155,N_7655,N_7981);
nand U8156 (N_8156,N_7842,N_7946);
or U8157 (N_8157,N_7642,N_7617);
nand U8158 (N_8158,N_7762,N_7989);
nand U8159 (N_8159,N_7838,N_7699);
nand U8160 (N_8160,N_7818,N_7637);
nor U8161 (N_8161,N_7628,N_7787);
or U8162 (N_8162,N_7618,N_7703);
and U8163 (N_8163,N_7960,N_7782);
nor U8164 (N_8164,N_7695,N_7874);
nor U8165 (N_8165,N_7834,N_7657);
nor U8166 (N_8166,N_7684,N_7883);
and U8167 (N_8167,N_7801,N_7895);
nor U8168 (N_8168,N_7643,N_7658);
and U8169 (N_8169,N_7925,N_7768);
and U8170 (N_8170,N_7896,N_7688);
or U8171 (N_8171,N_7825,N_7663);
and U8172 (N_8172,N_7837,N_7827);
nor U8173 (N_8173,N_7745,N_7944);
nor U8174 (N_8174,N_7780,N_7939);
or U8175 (N_8175,N_7876,N_7681);
nand U8176 (N_8176,N_7675,N_7602);
nor U8177 (N_8177,N_7649,N_7634);
or U8178 (N_8178,N_7737,N_7909);
and U8179 (N_8179,N_7889,N_7863);
or U8180 (N_8180,N_7775,N_7916);
nand U8181 (N_8181,N_7952,N_7763);
nor U8182 (N_8182,N_7988,N_7636);
and U8183 (N_8183,N_7832,N_7615);
or U8184 (N_8184,N_7994,N_7664);
or U8185 (N_8185,N_7871,N_7789);
and U8186 (N_8186,N_7753,N_7738);
nand U8187 (N_8187,N_7844,N_7931);
nor U8188 (N_8188,N_7760,N_7974);
xnor U8189 (N_8189,N_7955,N_7855);
nor U8190 (N_8190,N_7608,N_7967);
nor U8191 (N_8191,N_7799,N_7860);
and U8192 (N_8192,N_7776,N_7821);
or U8193 (N_8193,N_7930,N_7609);
nand U8194 (N_8194,N_7765,N_7996);
and U8195 (N_8195,N_7741,N_7866);
or U8196 (N_8196,N_7811,N_7975);
nor U8197 (N_8197,N_7833,N_7631);
and U8198 (N_8198,N_7853,N_7656);
nand U8199 (N_8199,N_7718,N_7757);
xnor U8200 (N_8200,N_7917,N_7841);
nand U8201 (N_8201,N_7722,N_7873);
or U8202 (N_8202,N_7823,N_7623);
nor U8203 (N_8203,N_7697,N_7609);
nand U8204 (N_8204,N_7769,N_7963);
or U8205 (N_8205,N_7723,N_7939);
nand U8206 (N_8206,N_7945,N_7935);
and U8207 (N_8207,N_7695,N_7806);
nor U8208 (N_8208,N_7759,N_7985);
nor U8209 (N_8209,N_7664,N_7908);
nor U8210 (N_8210,N_7892,N_7899);
or U8211 (N_8211,N_7631,N_7856);
nor U8212 (N_8212,N_7768,N_7712);
xor U8213 (N_8213,N_7635,N_7779);
and U8214 (N_8214,N_7705,N_7820);
nor U8215 (N_8215,N_7743,N_7757);
nand U8216 (N_8216,N_7823,N_7844);
and U8217 (N_8217,N_7908,N_7896);
or U8218 (N_8218,N_7844,N_7752);
and U8219 (N_8219,N_7658,N_7909);
nand U8220 (N_8220,N_7771,N_7765);
nand U8221 (N_8221,N_7929,N_7810);
nand U8222 (N_8222,N_7897,N_7991);
nor U8223 (N_8223,N_7951,N_7658);
nand U8224 (N_8224,N_7678,N_7885);
nand U8225 (N_8225,N_7740,N_7607);
nor U8226 (N_8226,N_7749,N_7750);
nor U8227 (N_8227,N_7893,N_7686);
or U8228 (N_8228,N_7791,N_7780);
or U8229 (N_8229,N_7924,N_7746);
or U8230 (N_8230,N_7885,N_7924);
or U8231 (N_8231,N_7845,N_7933);
and U8232 (N_8232,N_7610,N_7854);
or U8233 (N_8233,N_7640,N_7620);
nor U8234 (N_8234,N_7686,N_7774);
or U8235 (N_8235,N_7809,N_7990);
or U8236 (N_8236,N_7693,N_7741);
nor U8237 (N_8237,N_7958,N_7836);
or U8238 (N_8238,N_7768,N_7780);
and U8239 (N_8239,N_7837,N_7653);
or U8240 (N_8240,N_7650,N_7870);
and U8241 (N_8241,N_7920,N_7656);
nand U8242 (N_8242,N_7861,N_7789);
nor U8243 (N_8243,N_7978,N_7873);
or U8244 (N_8244,N_7817,N_7983);
or U8245 (N_8245,N_7882,N_7737);
nand U8246 (N_8246,N_7654,N_7770);
or U8247 (N_8247,N_7718,N_7950);
nand U8248 (N_8248,N_7801,N_7614);
nor U8249 (N_8249,N_7995,N_7833);
nor U8250 (N_8250,N_7929,N_7898);
or U8251 (N_8251,N_7779,N_7959);
or U8252 (N_8252,N_7855,N_7777);
or U8253 (N_8253,N_7669,N_7684);
or U8254 (N_8254,N_7841,N_7762);
nand U8255 (N_8255,N_7774,N_7756);
or U8256 (N_8256,N_7767,N_7806);
or U8257 (N_8257,N_7605,N_7951);
or U8258 (N_8258,N_7681,N_7854);
nor U8259 (N_8259,N_7629,N_7764);
and U8260 (N_8260,N_7882,N_7726);
nand U8261 (N_8261,N_7662,N_7714);
nand U8262 (N_8262,N_7785,N_7960);
and U8263 (N_8263,N_7994,N_7903);
and U8264 (N_8264,N_7972,N_7744);
and U8265 (N_8265,N_7716,N_7749);
and U8266 (N_8266,N_7764,N_7610);
or U8267 (N_8267,N_7789,N_7900);
nand U8268 (N_8268,N_7779,N_7611);
nand U8269 (N_8269,N_7996,N_7958);
and U8270 (N_8270,N_7997,N_7765);
nand U8271 (N_8271,N_7886,N_7747);
and U8272 (N_8272,N_7752,N_7728);
and U8273 (N_8273,N_7601,N_7751);
xor U8274 (N_8274,N_7600,N_7626);
nand U8275 (N_8275,N_7757,N_7963);
or U8276 (N_8276,N_7792,N_7923);
nand U8277 (N_8277,N_7735,N_7919);
or U8278 (N_8278,N_7689,N_7959);
and U8279 (N_8279,N_7854,N_7625);
and U8280 (N_8280,N_7824,N_7886);
nand U8281 (N_8281,N_7760,N_7755);
nand U8282 (N_8282,N_7807,N_7950);
or U8283 (N_8283,N_7729,N_7647);
nand U8284 (N_8284,N_7935,N_7927);
or U8285 (N_8285,N_7919,N_7626);
and U8286 (N_8286,N_7926,N_7979);
or U8287 (N_8287,N_7661,N_7803);
nand U8288 (N_8288,N_7871,N_7681);
nand U8289 (N_8289,N_7864,N_7876);
or U8290 (N_8290,N_7841,N_7709);
or U8291 (N_8291,N_7769,N_7658);
and U8292 (N_8292,N_7919,N_7797);
and U8293 (N_8293,N_7756,N_7725);
and U8294 (N_8294,N_7839,N_7837);
or U8295 (N_8295,N_7733,N_7850);
or U8296 (N_8296,N_7814,N_7831);
or U8297 (N_8297,N_7673,N_7897);
and U8298 (N_8298,N_7716,N_7842);
or U8299 (N_8299,N_7835,N_7956);
nand U8300 (N_8300,N_7602,N_7742);
and U8301 (N_8301,N_7725,N_7673);
and U8302 (N_8302,N_7859,N_7991);
nor U8303 (N_8303,N_7761,N_7824);
and U8304 (N_8304,N_7805,N_7624);
nor U8305 (N_8305,N_7967,N_7797);
or U8306 (N_8306,N_7639,N_7902);
nor U8307 (N_8307,N_7800,N_7941);
or U8308 (N_8308,N_7990,N_7943);
and U8309 (N_8309,N_7702,N_7838);
or U8310 (N_8310,N_7715,N_7617);
nand U8311 (N_8311,N_7617,N_7624);
or U8312 (N_8312,N_7782,N_7912);
and U8313 (N_8313,N_7806,N_7981);
nand U8314 (N_8314,N_7932,N_7995);
or U8315 (N_8315,N_7727,N_7846);
nor U8316 (N_8316,N_7668,N_7883);
nand U8317 (N_8317,N_7613,N_7722);
and U8318 (N_8318,N_7766,N_7816);
and U8319 (N_8319,N_7951,N_7833);
nand U8320 (N_8320,N_7935,N_7982);
or U8321 (N_8321,N_7849,N_7977);
nor U8322 (N_8322,N_7790,N_7977);
nor U8323 (N_8323,N_7634,N_7763);
or U8324 (N_8324,N_7828,N_7869);
or U8325 (N_8325,N_7885,N_7769);
or U8326 (N_8326,N_7821,N_7751);
and U8327 (N_8327,N_7793,N_7690);
nor U8328 (N_8328,N_7680,N_7876);
nor U8329 (N_8329,N_7892,N_7849);
nor U8330 (N_8330,N_7696,N_7755);
or U8331 (N_8331,N_7911,N_7744);
or U8332 (N_8332,N_7983,N_7703);
nor U8333 (N_8333,N_7891,N_7964);
nor U8334 (N_8334,N_7664,N_7682);
nand U8335 (N_8335,N_7921,N_7885);
and U8336 (N_8336,N_7890,N_7846);
and U8337 (N_8337,N_7638,N_7701);
nor U8338 (N_8338,N_7909,N_7786);
and U8339 (N_8339,N_7894,N_7606);
and U8340 (N_8340,N_7817,N_7653);
or U8341 (N_8341,N_7830,N_7829);
or U8342 (N_8342,N_7877,N_7856);
nor U8343 (N_8343,N_7850,N_7693);
nand U8344 (N_8344,N_7661,N_7676);
nor U8345 (N_8345,N_7764,N_7943);
or U8346 (N_8346,N_7614,N_7639);
nor U8347 (N_8347,N_7609,N_7894);
nor U8348 (N_8348,N_7982,N_7887);
or U8349 (N_8349,N_7858,N_7644);
nor U8350 (N_8350,N_7790,N_7744);
or U8351 (N_8351,N_7958,N_7737);
nor U8352 (N_8352,N_7610,N_7972);
and U8353 (N_8353,N_7956,N_7696);
or U8354 (N_8354,N_7735,N_7770);
nor U8355 (N_8355,N_7994,N_7862);
or U8356 (N_8356,N_7659,N_7639);
nor U8357 (N_8357,N_7931,N_7690);
nand U8358 (N_8358,N_7854,N_7804);
nand U8359 (N_8359,N_7778,N_7617);
or U8360 (N_8360,N_7918,N_7896);
nand U8361 (N_8361,N_7905,N_7607);
xor U8362 (N_8362,N_7858,N_7813);
or U8363 (N_8363,N_7937,N_7667);
nand U8364 (N_8364,N_7839,N_7938);
and U8365 (N_8365,N_7940,N_7993);
nor U8366 (N_8366,N_7990,N_7650);
and U8367 (N_8367,N_7763,N_7971);
nand U8368 (N_8368,N_7700,N_7629);
nand U8369 (N_8369,N_7931,N_7781);
and U8370 (N_8370,N_7600,N_7965);
and U8371 (N_8371,N_7767,N_7835);
nor U8372 (N_8372,N_7627,N_7687);
or U8373 (N_8373,N_7661,N_7653);
and U8374 (N_8374,N_7803,N_7879);
and U8375 (N_8375,N_7961,N_7922);
or U8376 (N_8376,N_7657,N_7909);
or U8377 (N_8377,N_7849,N_7639);
and U8378 (N_8378,N_7737,N_7769);
nor U8379 (N_8379,N_7688,N_7835);
or U8380 (N_8380,N_7673,N_7612);
nand U8381 (N_8381,N_7764,N_7690);
and U8382 (N_8382,N_7910,N_7831);
and U8383 (N_8383,N_7696,N_7726);
or U8384 (N_8384,N_7987,N_7638);
or U8385 (N_8385,N_7625,N_7883);
or U8386 (N_8386,N_7688,N_7912);
nor U8387 (N_8387,N_7950,N_7749);
or U8388 (N_8388,N_7693,N_7993);
nor U8389 (N_8389,N_7653,N_7818);
or U8390 (N_8390,N_7986,N_7789);
nand U8391 (N_8391,N_7857,N_7826);
nand U8392 (N_8392,N_7763,N_7658);
and U8393 (N_8393,N_7893,N_7623);
nand U8394 (N_8394,N_7687,N_7607);
or U8395 (N_8395,N_7652,N_7607);
nand U8396 (N_8396,N_7786,N_7673);
nor U8397 (N_8397,N_7680,N_7783);
nor U8398 (N_8398,N_7685,N_7954);
or U8399 (N_8399,N_7616,N_7896);
xor U8400 (N_8400,N_8321,N_8078);
nor U8401 (N_8401,N_8201,N_8179);
and U8402 (N_8402,N_8003,N_8237);
and U8403 (N_8403,N_8039,N_8159);
and U8404 (N_8404,N_8164,N_8045);
nand U8405 (N_8405,N_8210,N_8280);
nor U8406 (N_8406,N_8154,N_8376);
nor U8407 (N_8407,N_8354,N_8263);
and U8408 (N_8408,N_8370,N_8057);
or U8409 (N_8409,N_8310,N_8181);
and U8410 (N_8410,N_8291,N_8099);
nor U8411 (N_8411,N_8026,N_8233);
nand U8412 (N_8412,N_8002,N_8234);
and U8413 (N_8413,N_8082,N_8115);
nor U8414 (N_8414,N_8117,N_8343);
nand U8415 (N_8415,N_8085,N_8202);
or U8416 (N_8416,N_8007,N_8023);
nand U8417 (N_8417,N_8194,N_8292);
nor U8418 (N_8418,N_8329,N_8006);
and U8419 (N_8419,N_8130,N_8256);
or U8420 (N_8420,N_8389,N_8177);
or U8421 (N_8421,N_8037,N_8012);
or U8422 (N_8422,N_8157,N_8107);
nand U8423 (N_8423,N_8076,N_8294);
or U8424 (N_8424,N_8249,N_8196);
nand U8425 (N_8425,N_8273,N_8010);
and U8426 (N_8426,N_8379,N_8308);
nand U8427 (N_8427,N_8024,N_8261);
nand U8428 (N_8428,N_8183,N_8298);
and U8429 (N_8429,N_8255,N_8001);
and U8430 (N_8430,N_8300,N_8351);
and U8431 (N_8431,N_8288,N_8088);
nand U8432 (N_8432,N_8284,N_8034);
or U8433 (N_8433,N_8043,N_8283);
nor U8434 (N_8434,N_8165,N_8189);
and U8435 (N_8435,N_8213,N_8250);
or U8436 (N_8436,N_8173,N_8035);
nor U8437 (N_8437,N_8286,N_8374);
nand U8438 (N_8438,N_8050,N_8339);
and U8439 (N_8439,N_8268,N_8209);
nor U8440 (N_8440,N_8277,N_8315);
nand U8441 (N_8441,N_8146,N_8048);
and U8442 (N_8442,N_8191,N_8136);
nor U8443 (N_8443,N_8295,N_8122);
or U8444 (N_8444,N_8242,N_8391);
nand U8445 (N_8445,N_8325,N_8208);
or U8446 (N_8446,N_8028,N_8015);
and U8447 (N_8447,N_8276,N_8285);
nor U8448 (N_8448,N_8333,N_8172);
nor U8449 (N_8449,N_8124,N_8114);
nand U8450 (N_8450,N_8128,N_8005);
nand U8451 (N_8451,N_8320,N_8075);
and U8452 (N_8452,N_8086,N_8131);
nor U8453 (N_8453,N_8153,N_8394);
and U8454 (N_8454,N_8123,N_8017);
nor U8455 (N_8455,N_8305,N_8171);
nand U8456 (N_8456,N_8218,N_8365);
or U8457 (N_8457,N_8254,N_8104);
nand U8458 (N_8458,N_8323,N_8383);
or U8459 (N_8459,N_8169,N_8135);
or U8460 (N_8460,N_8054,N_8205);
xor U8461 (N_8461,N_8342,N_8200);
nand U8462 (N_8462,N_8299,N_8101);
nand U8463 (N_8463,N_8113,N_8143);
and U8464 (N_8464,N_8190,N_8373);
and U8465 (N_8465,N_8390,N_8160);
nand U8466 (N_8466,N_8060,N_8144);
and U8467 (N_8467,N_8064,N_8396);
nand U8468 (N_8468,N_8059,N_8000);
nand U8469 (N_8469,N_8009,N_8049);
or U8470 (N_8470,N_8334,N_8161);
nand U8471 (N_8471,N_8386,N_8223);
nand U8472 (N_8472,N_8366,N_8367);
or U8473 (N_8473,N_8182,N_8167);
nand U8474 (N_8474,N_8170,N_8248);
nand U8475 (N_8475,N_8092,N_8041);
and U8476 (N_8476,N_8369,N_8047);
nor U8477 (N_8477,N_8175,N_8044);
and U8478 (N_8478,N_8225,N_8281);
or U8479 (N_8479,N_8080,N_8303);
or U8480 (N_8480,N_8253,N_8073);
nor U8481 (N_8481,N_8304,N_8319);
and U8482 (N_8482,N_8258,N_8068);
or U8483 (N_8483,N_8055,N_8166);
nand U8484 (N_8484,N_8061,N_8004);
and U8485 (N_8485,N_8081,N_8235);
nand U8486 (N_8486,N_8014,N_8228);
or U8487 (N_8487,N_8387,N_8309);
or U8488 (N_8488,N_8178,N_8158);
or U8489 (N_8489,N_8397,N_8262);
nor U8490 (N_8490,N_8239,N_8251);
nor U8491 (N_8491,N_8382,N_8030);
and U8492 (N_8492,N_8069,N_8100);
nor U8493 (N_8493,N_8332,N_8274);
or U8494 (N_8494,N_8188,N_8021);
nor U8495 (N_8495,N_8247,N_8380);
nor U8496 (N_8496,N_8241,N_8138);
nor U8497 (N_8497,N_8053,N_8216);
or U8498 (N_8498,N_8150,N_8119);
or U8499 (N_8499,N_8363,N_8331);
or U8500 (N_8500,N_8011,N_8349);
nand U8501 (N_8501,N_8312,N_8013);
nor U8502 (N_8502,N_8084,N_8290);
nand U8503 (N_8503,N_8065,N_8140);
nor U8504 (N_8504,N_8199,N_8067);
nor U8505 (N_8505,N_8240,N_8317);
nand U8506 (N_8506,N_8350,N_8032);
nand U8507 (N_8507,N_8186,N_8212);
nand U8508 (N_8508,N_8215,N_8324);
nand U8509 (N_8509,N_8192,N_8203);
nor U8510 (N_8510,N_8125,N_8353);
and U8511 (N_8511,N_8279,N_8344);
nand U8512 (N_8512,N_8307,N_8244);
or U8513 (N_8513,N_8066,N_8377);
and U8514 (N_8514,N_8381,N_8058);
nor U8515 (N_8515,N_8220,N_8145);
nand U8516 (N_8516,N_8393,N_8340);
or U8517 (N_8517,N_8091,N_8127);
or U8518 (N_8518,N_8302,N_8133);
nand U8519 (N_8519,N_8222,N_8266);
and U8520 (N_8520,N_8278,N_8384);
nor U8521 (N_8521,N_8371,N_8226);
nand U8522 (N_8522,N_8301,N_8399);
or U8523 (N_8523,N_8090,N_8282);
and U8524 (N_8524,N_8163,N_8306);
and U8525 (N_8525,N_8198,N_8327);
nand U8526 (N_8526,N_8033,N_8108);
and U8527 (N_8527,N_8142,N_8094);
and U8528 (N_8528,N_8347,N_8093);
nor U8529 (N_8529,N_8042,N_8341);
nand U8530 (N_8530,N_8388,N_8176);
nand U8531 (N_8531,N_8185,N_8238);
and U8532 (N_8532,N_8105,N_8008);
nand U8533 (N_8533,N_8195,N_8120);
and U8534 (N_8534,N_8134,N_8027);
or U8535 (N_8535,N_8221,N_8072);
nand U8536 (N_8536,N_8378,N_8155);
or U8537 (N_8537,N_8022,N_8345);
nand U8538 (N_8538,N_8264,N_8265);
or U8539 (N_8539,N_8296,N_8230);
nand U8540 (N_8540,N_8020,N_8311);
nand U8541 (N_8541,N_8246,N_8174);
nand U8542 (N_8542,N_8346,N_8031);
nor U8543 (N_8543,N_8063,N_8089);
nor U8544 (N_8544,N_8180,N_8335);
and U8545 (N_8545,N_8079,N_8252);
nor U8546 (N_8546,N_8214,N_8372);
xor U8547 (N_8547,N_8187,N_8260);
and U8548 (N_8548,N_8168,N_8025);
and U8549 (N_8549,N_8217,N_8207);
nor U8550 (N_8550,N_8074,N_8149);
nand U8551 (N_8551,N_8368,N_8197);
nand U8552 (N_8552,N_8110,N_8129);
nand U8553 (N_8553,N_8243,N_8356);
and U8554 (N_8554,N_8137,N_8359);
and U8555 (N_8555,N_8109,N_8018);
nand U8556 (N_8556,N_8052,N_8193);
xor U8557 (N_8557,N_8102,N_8257);
nor U8558 (N_8558,N_8126,N_8267);
xnor U8559 (N_8559,N_8231,N_8147);
and U8560 (N_8560,N_8152,N_8271);
xor U8561 (N_8561,N_8019,N_8337);
and U8562 (N_8562,N_8322,N_8070);
nand U8563 (N_8563,N_8375,N_8211);
and U8564 (N_8564,N_8358,N_8316);
nand U8565 (N_8565,N_8336,N_8098);
and U8566 (N_8566,N_8330,N_8361);
nand U8567 (N_8567,N_8224,N_8040);
nor U8568 (N_8568,N_8132,N_8206);
and U8569 (N_8569,N_8272,N_8116);
or U8570 (N_8570,N_8095,N_8156);
or U8571 (N_8571,N_8227,N_8289);
nand U8572 (N_8572,N_8111,N_8259);
and U8573 (N_8573,N_8364,N_8385);
and U8574 (N_8574,N_8270,N_8297);
nand U8575 (N_8575,N_8229,N_8348);
and U8576 (N_8576,N_8232,N_8083);
xor U8577 (N_8577,N_8318,N_8293);
and U8578 (N_8578,N_8121,N_8269);
nand U8579 (N_8579,N_8275,N_8355);
and U8580 (N_8580,N_8357,N_8219);
and U8581 (N_8581,N_8314,N_8071);
nand U8582 (N_8582,N_8112,N_8326);
nand U8583 (N_8583,N_8392,N_8245);
and U8584 (N_8584,N_8148,N_8360);
and U8585 (N_8585,N_8139,N_8362);
nor U8586 (N_8586,N_8016,N_8106);
nor U8587 (N_8587,N_8151,N_8204);
nand U8588 (N_8588,N_8352,N_8395);
or U8589 (N_8589,N_8313,N_8051);
xor U8590 (N_8590,N_8077,N_8062);
and U8591 (N_8591,N_8103,N_8056);
or U8592 (N_8592,N_8087,N_8184);
nor U8593 (N_8593,N_8328,N_8398);
and U8594 (N_8594,N_8141,N_8118);
or U8595 (N_8595,N_8046,N_8096);
and U8596 (N_8596,N_8236,N_8097);
nand U8597 (N_8597,N_8338,N_8162);
nand U8598 (N_8598,N_8036,N_8287);
or U8599 (N_8599,N_8029,N_8038);
nor U8600 (N_8600,N_8189,N_8079);
or U8601 (N_8601,N_8109,N_8186);
nand U8602 (N_8602,N_8045,N_8060);
nor U8603 (N_8603,N_8191,N_8020);
nor U8604 (N_8604,N_8213,N_8091);
nor U8605 (N_8605,N_8186,N_8112);
or U8606 (N_8606,N_8338,N_8230);
or U8607 (N_8607,N_8029,N_8233);
and U8608 (N_8608,N_8007,N_8334);
nor U8609 (N_8609,N_8142,N_8234);
or U8610 (N_8610,N_8079,N_8341);
and U8611 (N_8611,N_8286,N_8145);
xnor U8612 (N_8612,N_8044,N_8303);
nand U8613 (N_8613,N_8212,N_8262);
nor U8614 (N_8614,N_8118,N_8074);
or U8615 (N_8615,N_8284,N_8197);
or U8616 (N_8616,N_8323,N_8224);
and U8617 (N_8617,N_8108,N_8066);
nand U8618 (N_8618,N_8306,N_8288);
nand U8619 (N_8619,N_8303,N_8143);
and U8620 (N_8620,N_8238,N_8209);
nor U8621 (N_8621,N_8072,N_8231);
or U8622 (N_8622,N_8089,N_8160);
nand U8623 (N_8623,N_8048,N_8333);
nand U8624 (N_8624,N_8355,N_8040);
nor U8625 (N_8625,N_8191,N_8342);
nor U8626 (N_8626,N_8228,N_8393);
nand U8627 (N_8627,N_8195,N_8011);
or U8628 (N_8628,N_8290,N_8139);
nor U8629 (N_8629,N_8119,N_8017);
or U8630 (N_8630,N_8106,N_8038);
and U8631 (N_8631,N_8232,N_8329);
and U8632 (N_8632,N_8182,N_8337);
and U8633 (N_8633,N_8052,N_8014);
or U8634 (N_8634,N_8104,N_8151);
nand U8635 (N_8635,N_8295,N_8188);
or U8636 (N_8636,N_8132,N_8228);
and U8637 (N_8637,N_8168,N_8073);
nor U8638 (N_8638,N_8289,N_8336);
and U8639 (N_8639,N_8350,N_8105);
xnor U8640 (N_8640,N_8298,N_8042);
nand U8641 (N_8641,N_8357,N_8248);
nor U8642 (N_8642,N_8145,N_8043);
nor U8643 (N_8643,N_8353,N_8086);
nand U8644 (N_8644,N_8292,N_8033);
or U8645 (N_8645,N_8193,N_8323);
nand U8646 (N_8646,N_8042,N_8080);
or U8647 (N_8647,N_8318,N_8272);
or U8648 (N_8648,N_8353,N_8197);
or U8649 (N_8649,N_8061,N_8266);
and U8650 (N_8650,N_8143,N_8377);
nor U8651 (N_8651,N_8329,N_8376);
nand U8652 (N_8652,N_8122,N_8246);
nand U8653 (N_8653,N_8131,N_8351);
and U8654 (N_8654,N_8305,N_8343);
or U8655 (N_8655,N_8272,N_8242);
and U8656 (N_8656,N_8133,N_8181);
nor U8657 (N_8657,N_8237,N_8397);
or U8658 (N_8658,N_8208,N_8049);
or U8659 (N_8659,N_8123,N_8103);
or U8660 (N_8660,N_8030,N_8199);
nand U8661 (N_8661,N_8125,N_8323);
and U8662 (N_8662,N_8277,N_8254);
nand U8663 (N_8663,N_8006,N_8154);
nand U8664 (N_8664,N_8134,N_8254);
nand U8665 (N_8665,N_8097,N_8081);
or U8666 (N_8666,N_8178,N_8029);
nor U8667 (N_8667,N_8163,N_8012);
nor U8668 (N_8668,N_8262,N_8394);
nand U8669 (N_8669,N_8217,N_8277);
or U8670 (N_8670,N_8348,N_8240);
nand U8671 (N_8671,N_8114,N_8281);
nor U8672 (N_8672,N_8134,N_8308);
nor U8673 (N_8673,N_8231,N_8159);
nor U8674 (N_8674,N_8223,N_8366);
nor U8675 (N_8675,N_8307,N_8350);
nand U8676 (N_8676,N_8390,N_8317);
nand U8677 (N_8677,N_8135,N_8108);
or U8678 (N_8678,N_8143,N_8263);
and U8679 (N_8679,N_8204,N_8011);
nand U8680 (N_8680,N_8321,N_8212);
and U8681 (N_8681,N_8219,N_8090);
and U8682 (N_8682,N_8098,N_8335);
or U8683 (N_8683,N_8188,N_8041);
nor U8684 (N_8684,N_8271,N_8227);
nor U8685 (N_8685,N_8330,N_8114);
and U8686 (N_8686,N_8388,N_8151);
and U8687 (N_8687,N_8303,N_8114);
nand U8688 (N_8688,N_8311,N_8016);
and U8689 (N_8689,N_8157,N_8224);
or U8690 (N_8690,N_8275,N_8185);
or U8691 (N_8691,N_8121,N_8350);
nand U8692 (N_8692,N_8083,N_8175);
nand U8693 (N_8693,N_8164,N_8356);
nor U8694 (N_8694,N_8242,N_8204);
or U8695 (N_8695,N_8256,N_8057);
or U8696 (N_8696,N_8342,N_8316);
or U8697 (N_8697,N_8065,N_8394);
nor U8698 (N_8698,N_8164,N_8332);
or U8699 (N_8699,N_8181,N_8204);
nand U8700 (N_8700,N_8121,N_8048);
or U8701 (N_8701,N_8334,N_8133);
or U8702 (N_8702,N_8066,N_8146);
and U8703 (N_8703,N_8346,N_8185);
nor U8704 (N_8704,N_8246,N_8057);
and U8705 (N_8705,N_8324,N_8336);
xnor U8706 (N_8706,N_8264,N_8308);
nor U8707 (N_8707,N_8013,N_8391);
or U8708 (N_8708,N_8168,N_8153);
and U8709 (N_8709,N_8271,N_8023);
and U8710 (N_8710,N_8190,N_8125);
nand U8711 (N_8711,N_8270,N_8378);
nand U8712 (N_8712,N_8389,N_8235);
nor U8713 (N_8713,N_8022,N_8329);
and U8714 (N_8714,N_8331,N_8220);
nor U8715 (N_8715,N_8230,N_8126);
and U8716 (N_8716,N_8086,N_8144);
or U8717 (N_8717,N_8127,N_8238);
nand U8718 (N_8718,N_8208,N_8334);
nor U8719 (N_8719,N_8032,N_8330);
nand U8720 (N_8720,N_8147,N_8168);
nor U8721 (N_8721,N_8206,N_8275);
nand U8722 (N_8722,N_8114,N_8046);
or U8723 (N_8723,N_8277,N_8088);
nand U8724 (N_8724,N_8078,N_8059);
or U8725 (N_8725,N_8109,N_8004);
nand U8726 (N_8726,N_8359,N_8095);
nand U8727 (N_8727,N_8093,N_8078);
and U8728 (N_8728,N_8293,N_8350);
or U8729 (N_8729,N_8307,N_8030);
or U8730 (N_8730,N_8389,N_8212);
nand U8731 (N_8731,N_8341,N_8197);
and U8732 (N_8732,N_8392,N_8184);
nand U8733 (N_8733,N_8174,N_8375);
or U8734 (N_8734,N_8167,N_8145);
nor U8735 (N_8735,N_8123,N_8171);
and U8736 (N_8736,N_8210,N_8236);
nor U8737 (N_8737,N_8281,N_8387);
or U8738 (N_8738,N_8264,N_8152);
and U8739 (N_8739,N_8176,N_8315);
nand U8740 (N_8740,N_8331,N_8172);
or U8741 (N_8741,N_8348,N_8074);
nand U8742 (N_8742,N_8206,N_8078);
nor U8743 (N_8743,N_8046,N_8369);
or U8744 (N_8744,N_8123,N_8168);
or U8745 (N_8745,N_8332,N_8243);
nand U8746 (N_8746,N_8164,N_8302);
and U8747 (N_8747,N_8377,N_8241);
nand U8748 (N_8748,N_8189,N_8124);
and U8749 (N_8749,N_8236,N_8039);
xnor U8750 (N_8750,N_8012,N_8225);
and U8751 (N_8751,N_8204,N_8340);
or U8752 (N_8752,N_8020,N_8263);
nand U8753 (N_8753,N_8123,N_8142);
or U8754 (N_8754,N_8042,N_8115);
nor U8755 (N_8755,N_8048,N_8369);
nor U8756 (N_8756,N_8117,N_8394);
nor U8757 (N_8757,N_8122,N_8294);
nor U8758 (N_8758,N_8266,N_8123);
and U8759 (N_8759,N_8346,N_8322);
nand U8760 (N_8760,N_8025,N_8124);
nand U8761 (N_8761,N_8200,N_8011);
nor U8762 (N_8762,N_8013,N_8080);
nor U8763 (N_8763,N_8224,N_8024);
or U8764 (N_8764,N_8282,N_8177);
and U8765 (N_8765,N_8265,N_8225);
nor U8766 (N_8766,N_8291,N_8109);
and U8767 (N_8767,N_8374,N_8316);
and U8768 (N_8768,N_8128,N_8348);
or U8769 (N_8769,N_8190,N_8225);
nor U8770 (N_8770,N_8135,N_8274);
or U8771 (N_8771,N_8147,N_8379);
or U8772 (N_8772,N_8133,N_8271);
nand U8773 (N_8773,N_8177,N_8089);
nand U8774 (N_8774,N_8063,N_8261);
nand U8775 (N_8775,N_8369,N_8291);
nand U8776 (N_8776,N_8191,N_8269);
and U8777 (N_8777,N_8131,N_8270);
and U8778 (N_8778,N_8380,N_8034);
nand U8779 (N_8779,N_8009,N_8167);
and U8780 (N_8780,N_8150,N_8014);
and U8781 (N_8781,N_8271,N_8278);
xor U8782 (N_8782,N_8218,N_8190);
nor U8783 (N_8783,N_8281,N_8319);
and U8784 (N_8784,N_8017,N_8280);
nor U8785 (N_8785,N_8144,N_8365);
and U8786 (N_8786,N_8154,N_8105);
and U8787 (N_8787,N_8218,N_8051);
nand U8788 (N_8788,N_8209,N_8101);
or U8789 (N_8789,N_8011,N_8199);
or U8790 (N_8790,N_8075,N_8140);
or U8791 (N_8791,N_8088,N_8231);
or U8792 (N_8792,N_8343,N_8135);
nor U8793 (N_8793,N_8090,N_8133);
and U8794 (N_8794,N_8099,N_8262);
nor U8795 (N_8795,N_8189,N_8275);
or U8796 (N_8796,N_8291,N_8365);
nand U8797 (N_8797,N_8308,N_8091);
nand U8798 (N_8798,N_8210,N_8361);
or U8799 (N_8799,N_8258,N_8313);
nor U8800 (N_8800,N_8748,N_8709);
or U8801 (N_8801,N_8542,N_8445);
and U8802 (N_8802,N_8655,N_8713);
and U8803 (N_8803,N_8467,N_8762);
or U8804 (N_8804,N_8423,N_8565);
and U8805 (N_8805,N_8403,N_8418);
or U8806 (N_8806,N_8737,N_8407);
nor U8807 (N_8807,N_8450,N_8618);
nor U8808 (N_8808,N_8797,N_8624);
nand U8809 (N_8809,N_8634,N_8643);
nor U8810 (N_8810,N_8796,N_8436);
nor U8811 (N_8811,N_8465,N_8558);
or U8812 (N_8812,N_8688,N_8476);
or U8813 (N_8813,N_8587,N_8752);
and U8814 (N_8814,N_8656,N_8678);
nand U8815 (N_8815,N_8612,N_8607);
or U8816 (N_8816,N_8440,N_8720);
nor U8817 (N_8817,N_8771,N_8480);
and U8818 (N_8818,N_8710,N_8726);
nand U8819 (N_8819,N_8590,N_8416);
nor U8820 (N_8820,N_8576,N_8522);
and U8821 (N_8821,N_8511,N_8616);
or U8822 (N_8822,N_8553,N_8591);
and U8823 (N_8823,N_8657,N_8615);
or U8824 (N_8824,N_8438,N_8794);
nor U8825 (N_8825,N_8516,N_8547);
and U8826 (N_8826,N_8722,N_8583);
and U8827 (N_8827,N_8550,N_8686);
nand U8828 (N_8828,N_8602,N_8673);
nand U8829 (N_8829,N_8441,N_8484);
or U8830 (N_8830,N_8543,N_8617);
nor U8831 (N_8831,N_8654,N_8652);
nor U8832 (N_8832,N_8408,N_8533);
nor U8833 (N_8833,N_8404,N_8665);
nand U8834 (N_8834,N_8676,N_8473);
nor U8835 (N_8835,N_8498,N_8585);
nor U8836 (N_8836,N_8700,N_8798);
and U8837 (N_8837,N_8462,N_8777);
or U8838 (N_8838,N_8515,N_8589);
and U8839 (N_8839,N_8548,N_8672);
and U8840 (N_8840,N_8733,N_8660);
and U8841 (N_8841,N_8429,N_8491);
and U8842 (N_8842,N_8468,N_8725);
or U8843 (N_8843,N_8717,N_8756);
and U8844 (N_8844,N_8471,N_8708);
or U8845 (N_8845,N_8577,N_8651);
nand U8846 (N_8846,N_8417,N_8513);
nor U8847 (N_8847,N_8744,N_8446);
nand U8848 (N_8848,N_8639,N_8755);
nand U8849 (N_8849,N_8563,N_8691);
and U8850 (N_8850,N_8714,N_8782);
nor U8851 (N_8851,N_8723,N_8781);
or U8852 (N_8852,N_8568,N_8409);
and U8853 (N_8853,N_8443,N_8658);
or U8854 (N_8854,N_8734,N_8598);
nand U8855 (N_8855,N_8431,N_8411);
or U8856 (N_8856,N_8420,N_8694);
nand U8857 (N_8857,N_8736,N_8560);
and U8858 (N_8858,N_8791,N_8746);
and U8859 (N_8859,N_8638,N_8758);
nand U8860 (N_8860,N_8627,N_8519);
or U8861 (N_8861,N_8728,N_8432);
and U8862 (N_8862,N_8456,N_8427);
and U8863 (N_8863,N_8489,N_8721);
and U8864 (N_8864,N_8626,N_8479);
nor U8865 (N_8865,N_8493,N_8697);
nor U8866 (N_8866,N_8631,N_8650);
and U8867 (N_8867,N_8772,N_8597);
nand U8868 (N_8868,N_8584,N_8502);
nor U8869 (N_8869,N_8580,N_8716);
and U8870 (N_8870,N_8641,N_8774);
nor U8871 (N_8871,N_8754,N_8463);
nor U8872 (N_8872,N_8768,N_8689);
or U8873 (N_8873,N_8646,N_8606);
nand U8874 (N_8874,N_8569,N_8570);
and U8875 (N_8875,N_8653,N_8464);
nand U8876 (N_8876,N_8659,N_8595);
nor U8877 (N_8877,N_8472,N_8444);
and U8878 (N_8878,N_8727,N_8452);
nor U8879 (N_8879,N_8559,N_8766);
and U8880 (N_8880,N_8698,N_8434);
or U8881 (N_8881,N_8719,N_8675);
and U8882 (N_8882,N_8501,N_8644);
and U8883 (N_8883,N_8786,N_8776);
nor U8884 (N_8884,N_8545,N_8740);
nor U8885 (N_8885,N_8753,N_8635);
nand U8886 (N_8886,N_8622,N_8611);
nor U8887 (N_8887,N_8566,N_8537);
nor U8888 (N_8888,N_8579,N_8425);
nor U8889 (N_8889,N_8799,N_8745);
nor U8890 (N_8890,N_8681,N_8410);
nor U8891 (N_8891,N_8601,N_8625);
or U8892 (N_8892,N_8790,N_8668);
and U8893 (N_8893,N_8594,N_8731);
nor U8894 (N_8894,N_8402,N_8704);
or U8895 (N_8895,N_8421,N_8680);
nand U8896 (N_8896,N_8603,N_8507);
and U8897 (N_8897,N_8629,N_8414);
or U8898 (N_8898,N_8690,N_8715);
and U8899 (N_8899,N_8663,N_8599);
nand U8900 (N_8900,N_8750,N_8509);
nor U8901 (N_8901,N_8706,N_8481);
or U8902 (N_8902,N_8767,N_8729);
nand U8903 (N_8903,N_8453,N_8751);
nor U8904 (N_8904,N_8564,N_8460);
and U8905 (N_8905,N_8496,N_8632);
nor U8906 (N_8906,N_8492,N_8528);
nand U8907 (N_8907,N_8705,N_8536);
and U8908 (N_8908,N_8439,N_8670);
nand U8909 (N_8909,N_8621,N_8422);
or U8910 (N_8910,N_8490,N_8712);
nand U8911 (N_8911,N_8741,N_8400);
and U8912 (N_8912,N_8764,N_8412);
and U8913 (N_8913,N_8649,N_8765);
or U8914 (N_8914,N_8524,N_8692);
nor U8915 (N_8915,N_8699,N_8572);
or U8916 (N_8916,N_8784,N_8451);
nor U8917 (N_8917,N_8711,N_8529);
nor U8918 (N_8918,N_8592,N_8544);
nor U8919 (N_8919,N_8466,N_8459);
or U8920 (N_8920,N_8695,N_8671);
nand U8921 (N_8921,N_8783,N_8415);
nand U8922 (N_8922,N_8426,N_8555);
and U8923 (N_8923,N_8578,N_8795);
nand U8924 (N_8924,N_8534,N_8787);
nor U8925 (N_8925,N_8619,N_8478);
nand U8926 (N_8926,N_8494,N_8623);
nor U8927 (N_8927,N_8541,N_8428);
nor U8928 (N_8928,N_8549,N_8401);
or U8929 (N_8929,N_8682,N_8495);
nand U8930 (N_8930,N_8530,N_8769);
nand U8931 (N_8931,N_8455,N_8551);
nor U8932 (N_8932,N_8540,N_8556);
or U8933 (N_8933,N_8525,N_8730);
nand U8934 (N_8934,N_8770,N_8454);
nor U8935 (N_8935,N_8596,N_8527);
or U8936 (N_8936,N_8669,N_8789);
nor U8937 (N_8937,N_8779,N_8664);
or U8938 (N_8938,N_8510,N_8531);
nand U8939 (N_8939,N_8469,N_8437);
nor U8940 (N_8940,N_8505,N_8503);
nor U8941 (N_8941,N_8461,N_8546);
or U8942 (N_8942,N_8637,N_8512);
or U8943 (N_8943,N_8645,N_8487);
or U8944 (N_8944,N_8647,N_8683);
and U8945 (N_8945,N_8486,N_8482);
nor U8946 (N_8946,N_8539,N_8488);
nor U8947 (N_8947,N_8620,N_8588);
and U8948 (N_8948,N_8778,N_8447);
or U8949 (N_8949,N_8574,N_8636);
xnor U8950 (N_8950,N_8506,N_8448);
nor U8951 (N_8951,N_8442,N_8604);
and U8952 (N_8952,N_8773,N_8593);
or U8953 (N_8953,N_8483,N_8609);
nor U8954 (N_8954,N_8633,N_8757);
and U8955 (N_8955,N_8517,N_8685);
nand U8956 (N_8956,N_8424,N_8605);
nand U8957 (N_8957,N_8608,N_8666);
nor U8958 (N_8958,N_8735,N_8780);
or U8959 (N_8959,N_8687,N_8732);
nor U8960 (N_8960,N_8693,N_8648);
or U8961 (N_8961,N_8497,N_8743);
nand U8962 (N_8962,N_8433,N_8475);
nand U8963 (N_8963,N_8586,N_8413);
nor U8964 (N_8964,N_8739,N_8661);
nor U8965 (N_8965,N_8535,N_8667);
nor U8966 (N_8966,N_8600,N_8514);
nand U8967 (N_8967,N_8457,N_8523);
and U8968 (N_8968,N_8788,N_8696);
nand U8969 (N_8969,N_8747,N_8526);
nor U8970 (N_8970,N_8724,N_8742);
or U8971 (N_8971,N_8775,N_8642);
nand U8972 (N_8972,N_8573,N_8581);
or U8973 (N_8973,N_8701,N_8749);
nor U8974 (N_8974,N_8405,N_8485);
nor U8975 (N_8975,N_8759,N_8521);
nor U8976 (N_8976,N_8458,N_8562);
and U8977 (N_8977,N_8640,N_8435);
and U8978 (N_8978,N_8449,N_8793);
nor U8979 (N_8979,N_8504,N_8738);
and U8980 (N_8980,N_8785,N_8718);
or U8981 (N_8981,N_8499,N_8792);
and U8982 (N_8982,N_8520,N_8474);
or U8983 (N_8983,N_8500,N_8703);
nand U8984 (N_8984,N_8430,N_8707);
or U8985 (N_8985,N_8684,N_8508);
or U8986 (N_8986,N_8406,N_8532);
nand U8987 (N_8987,N_8610,N_8614);
and U8988 (N_8988,N_8470,N_8477);
or U8989 (N_8989,N_8582,N_8763);
nor U8990 (N_8990,N_8538,N_8419);
nor U8991 (N_8991,N_8702,N_8571);
or U8992 (N_8992,N_8677,N_8557);
nand U8993 (N_8993,N_8567,N_8575);
or U8994 (N_8994,N_8561,N_8662);
nand U8995 (N_8995,N_8679,N_8613);
nand U8996 (N_8996,N_8630,N_8518);
or U8997 (N_8997,N_8760,N_8761);
nand U8998 (N_8998,N_8552,N_8554);
and U8999 (N_8999,N_8628,N_8674);
nand U9000 (N_9000,N_8798,N_8539);
and U9001 (N_9001,N_8665,N_8558);
or U9002 (N_9002,N_8488,N_8670);
nor U9003 (N_9003,N_8573,N_8790);
nand U9004 (N_9004,N_8411,N_8427);
xor U9005 (N_9005,N_8416,N_8473);
nand U9006 (N_9006,N_8758,N_8410);
and U9007 (N_9007,N_8409,N_8532);
and U9008 (N_9008,N_8432,N_8701);
and U9009 (N_9009,N_8423,N_8443);
nor U9010 (N_9010,N_8659,N_8550);
nand U9011 (N_9011,N_8486,N_8736);
nor U9012 (N_9012,N_8417,N_8620);
or U9013 (N_9013,N_8776,N_8553);
and U9014 (N_9014,N_8687,N_8778);
nor U9015 (N_9015,N_8586,N_8508);
or U9016 (N_9016,N_8770,N_8518);
or U9017 (N_9017,N_8637,N_8542);
nor U9018 (N_9018,N_8713,N_8618);
nand U9019 (N_9019,N_8586,N_8616);
nand U9020 (N_9020,N_8430,N_8718);
nor U9021 (N_9021,N_8602,N_8537);
nand U9022 (N_9022,N_8799,N_8519);
nand U9023 (N_9023,N_8485,N_8636);
nor U9024 (N_9024,N_8681,N_8545);
and U9025 (N_9025,N_8408,N_8440);
nor U9026 (N_9026,N_8512,N_8721);
nor U9027 (N_9027,N_8658,N_8400);
nand U9028 (N_9028,N_8544,N_8629);
or U9029 (N_9029,N_8624,N_8603);
or U9030 (N_9030,N_8553,N_8667);
nor U9031 (N_9031,N_8618,N_8562);
nand U9032 (N_9032,N_8427,N_8505);
nor U9033 (N_9033,N_8583,N_8523);
nor U9034 (N_9034,N_8502,N_8408);
nand U9035 (N_9035,N_8747,N_8642);
or U9036 (N_9036,N_8472,N_8425);
nor U9037 (N_9037,N_8472,N_8750);
nand U9038 (N_9038,N_8783,N_8768);
or U9039 (N_9039,N_8726,N_8518);
nor U9040 (N_9040,N_8656,N_8602);
or U9041 (N_9041,N_8608,N_8565);
nand U9042 (N_9042,N_8777,N_8554);
or U9043 (N_9043,N_8784,N_8577);
nand U9044 (N_9044,N_8549,N_8768);
and U9045 (N_9045,N_8733,N_8719);
nor U9046 (N_9046,N_8485,N_8513);
or U9047 (N_9047,N_8713,N_8615);
and U9048 (N_9048,N_8514,N_8433);
nor U9049 (N_9049,N_8747,N_8719);
or U9050 (N_9050,N_8646,N_8755);
or U9051 (N_9051,N_8763,N_8456);
or U9052 (N_9052,N_8401,N_8718);
nand U9053 (N_9053,N_8676,N_8591);
nor U9054 (N_9054,N_8412,N_8704);
and U9055 (N_9055,N_8445,N_8708);
and U9056 (N_9056,N_8758,N_8708);
and U9057 (N_9057,N_8736,N_8651);
or U9058 (N_9058,N_8424,N_8408);
nor U9059 (N_9059,N_8564,N_8578);
nor U9060 (N_9060,N_8410,N_8457);
and U9061 (N_9061,N_8734,N_8600);
nand U9062 (N_9062,N_8480,N_8665);
nand U9063 (N_9063,N_8404,N_8754);
nor U9064 (N_9064,N_8528,N_8695);
nand U9065 (N_9065,N_8559,N_8429);
or U9066 (N_9066,N_8771,N_8454);
nor U9067 (N_9067,N_8775,N_8522);
and U9068 (N_9068,N_8732,N_8674);
or U9069 (N_9069,N_8786,N_8539);
or U9070 (N_9070,N_8766,N_8661);
nor U9071 (N_9071,N_8442,N_8668);
nor U9072 (N_9072,N_8437,N_8704);
nor U9073 (N_9073,N_8605,N_8619);
nor U9074 (N_9074,N_8495,N_8580);
or U9075 (N_9075,N_8509,N_8542);
nor U9076 (N_9076,N_8725,N_8538);
nand U9077 (N_9077,N_8668,N_8558);
and U9078 (N_9078,N_8615,N_8534);
and U9079 (N_9079,N_8517,N_8512);
and U9080 (N_9080,N_8594,N_8649);
and U9081 (N_9081,N_8454,N_8596);
nand U9082 (N_9082,N_8756,N_8603);
and U9083 (N_9083,N_8789,N_8420);
or U9084 (N_9084,N_8642,N_8486);
nor U9085 (N_9085,N_8761,N_8436);
nor U9086 (N_9086,N_8606,N_8777);
or U9087 (N_9087,N_8671,N_8722);
nor U9088 (N_9088,N_8591,N_8590);
or U9089 (N_9089,N_8551,N_8711);
and U9090 (N_9090,N_8756,N_8426);
nor U9091 (N_9091,N_8559,N_8623);
nor U9092 (N_9092,N_8476,N_8653);
and U9093 (N_9093,N_8492,N_8742);
nor U9094 (N_9094,N_8535,N_8462);
or U9095 (N_9095,N_8648,N_8796);
and U9096 (N_9096,N_8554,N_8402);
nand U9097 (N_9097,N_8415,N_8603);
nor U9098 (N_9098,N_8702,N_8796);
and U9099 (N_9099,N_8570,N_8727);
or U9100 (N_9100,N_8611,N_8770);
nand U9101 (N_9101,N_8664,N_8489);
or U9102 (N_9102,N_8530,N_8607);
nor U9103 (N_9103,N_8610,N_8743);
or U9104 (N_9104,N_8408,N_8751);
nor U9105 (N_9105,N_8774,N_8435);
nand U9106 (N_9106,N_8435,N_8460);
nand U9107 (N_9107,N_8553,N_8567);
nor U9108 (N_9108,N_8423,N_8764);
or U9109 (N_9109,N_8764,N_8441);
nand U9110 (N_9110,N_8539,N_8462);
nor U9111 (N_9111,N_8779,N_8616);
nor U9112 (N_9112,N_8568,N_8521);
and U9113 (N_9113,N_8700,N_8463);
or U9114 (N_9114,N_8492,N_8734);
nor U9115 (N_9115,N_8523,N_8469);
nor U9116 (N_9116,N_8416,N_8463);
and U9117 (N_9117,N_8618,N_8532);
nor U9118 (N_9118,N_8659,N_8481);
nand U9119 (N_9119,N_8460,N_8737);
and U9120 (N_9120,N_8608,N_8563);
or U9121 (N_9121,N_8511,N_8765);
or U9122 (N_9122,N_8580,N_8529);
nand U9123 (N_9123,N_8498,N_8529);
or U9124 (N_9124,N_8598,N_8561);
nand U9125 (N_9125,N_8412,N_8494);
and U9126 (N_9126,N_8715,N_8653);
nand U9127 (N_9127,N_8417,N_8580);
nor U9128 (N_9128,N_8606,N_8578);
and U9129 (N_9129,N_8470,N_8453);
nand U9130 (N_9130,N_8711,N_8602);
and U9131 (N_9131,N_8440,N_8772);
nand U9132 (N_9132,N_8457,N_8595);
or U9133 (N_9133,N_8548,N_8793);
nor U9134 (N_9134,N_8724,N_8473);
nor U9135 (N_9135,N_8492,N_8513);
nor U9136 (N_9136,N_8651,N_8743);
nor U9137 (N_9137,N_8592,N_8453);
or U9138 (N_9138,N_8462,N_8733);
nor U9139 (N_9139,N_8640,N_8497);
nand U9140 (N_9140,N_8728,N_8630);
nand U9141 (N_9141,N_8754,N_8539);
nand U9142 (N_9142,N_8430,N_8421);
and U9143 (N_9143,N_8792,N_8428);
and U9144 (N_9144,N_8696,N_8652);
nor U9145 (N_9145,N_8560,N_8772);
nand U9146 (N_9146,N_8575,N_8475);
nor U9147 (N_9147,N_8663,N_8724);
and U9148 (N_9148,N_8718,N_8406);
nand U9149 (N_9149,N_8595,N_8684);
nand U9150 (N_9150,N_8732,N_8635);
nand U9151 (N_9151,N_8729,N_8531);
nor U9152 (N_9152,N_8546,N_8690);
nor U9153 (N_9153,N_8462,N_8405);
nand U9154 (N_9154,N_8629,N_8762);
or U9155 (N_9155,N_8459,N_8510);
nor U9156 (N_9156,N_8536,N_8467);
nor U9157 (N_9157,N_8741,N_8405);
or U9158 (N_9158,N_8773,N_8638);
and U9159 (N_9159,N_8710,N_8670);
nor U9160 (N_9160,N_8528,N_8459);
or U9161 (N_9161,N_8774,N_8520);
or U9162 (N_9162,N_8433,N_8686);
and U9163 (N_9163,N_8408,N_8543);
nand U9164 (N_9164,N_8642,N_8669);
nand U9165 (N_9165,N_8690,N_8786);
nor U9166 (N_9166,N_8558,N_8654);
nand U9167 (N_9167,N_8774,N_8775);
nand U9168 (N_9168,N_8418,N_8657);
nand U9169 (N_9169,N_8690,N_8512);
or U9170 (N_9170,N_8602,N_8592);
or U9171 (N_9171,N_8561,N_8433);
and U9172 (N_9172,N_8775,N_8692);
or U9173 (N_9173,N_8588,N_8407);
or U9174 (N_9174,N_8571,N_8490);
nand U9175 (N_9175,N_8412,N_8492);
or U9176 (N_9176,N_8550,N_8579);
and U9177 (N_9177,N_8684,N_8487);
and U9178 (N_9178,N_8498,N_8503);
nand U9179 (N_9179,N_8575,N_8597);
nor U9180 (N_9180,N_8408,N_8584);
nand U9181 (N_9181,N_8660,N_8681);
nand U9182 (N_9182,N_8552,N_8421);
and U9183 (N_9183,N_8739,N_8534);
or U9184 (N_9184,N_8734,N_8414);
nand U9185 (N_9185,N_8480,N_8789);
nand U9186 (N_9186,N_8593,N_8797);
and U9187 (N_9187,N_8596,N_8483);
nand U9188 (N_9188,N_8443,N_8503);
and U9189 (N_9189,N_8552,N_8485);
or U9190 (N_9190,N_8680,N_8755);
or U9191 (N_9191,N_8620,N_8673);
or U9192 (N_9192,N_8699,N_8681);
nand U9193 (N_9193,N_8711,N_8631);
or U9194 (N_9194,N_8427,N_8533);
nand U9195 (N_9195,N_8644,N_8586);
nor U9196 (N_9196,N_8519,N_8409);
or U9197 (N_9197,N_8595,N_8458);
and U9198 (N_9198,N_8610,N_8455);
or U9199 (N_9199,N_8406,N_8432);
nand U9200 (N_9200,N_9003,N_8929);
and U9201 (N_9201,N_9101,N_8836);
or U9202 (N_9202,N_9141,N_8897);
nand U9203 (N_9203,N_9179,N_9162);
and U9204 (N_9204,N_8862,N_8900);
or U9205 (N_9205,N_8916,N_8899);
nand U9206 (N_9206,N_9180,N_8935);
or U9207 (N_9207,N_8936,N_8927);
nand U9208 (N_9208,N_8866,N_8944);
or U9209 (N_9209,N_8963,N_8951);
nor U9210 (N_9210,N_9111,N_9077);
and U9211 (N_9211,N_9036,N_8908);
nor U9212 (N_9212,N_8975,N_8956);
or U9213 (N_9213,N_9194,N_8955);
nor U9214 (N_9214,N_9035,N_9044);
nor U9215 (N_9215,N_8925,N_8923);
nand U9216 (N_9216,N_8864,N_9055);
and U9217 (N_9217,N_8873,N_9132);
or U9218 (N_9218,N_9178,N_8877);
and U9219 (N_9219,N_8855,N_8930);
and U9220 (N_9220,N_9063,N_9183);
or U9221 (N_9221,N_9142,N_8835);
and U9222 (N_9222,N_8945,N_8902);
nand U9223 (N_9223,N_8978,N_9193);
or U9224 (N_9224,N_9197,N_8952);
and U9225 (N_9225,N_8840,N_9145);
or U9226 (N_9226,N_8903,N_8852);
or U9227 (N_9227,N_9074,N_9081);
and U9228 (N_9228,N_9150,N_9015);
and U9229 (N_9229,N_8977,N_9115);
and U9230 (N_9230,N_9023,N_8878);
nand U9231 (N_9231,N_8827,N_9076);
nand U9232 (N_9232,N_8904,N_8882);
nor U9233 (N_9233,N_8806,N_8898);
nand U9234 (N_9234,N_9087,N_9041);
nand U9235 (N_9235,N_9149,N_8831);
or U9236 (N_9236,N_9169,N_9059);
or U9237 (N_9237,N_9028,N_8808);
and U9238 (N_9238,N_9102,N_8843);
nor U9239 (N_9239,N_8921,N_8879);
nand U9240 (N_9240,N_9113,N_9026);
nand U9241 (N_9241,N_8822,N_9070);
and U9242 (N_9242,N_8815,N_8931);
and U9243 (N_9243,N_8809,N_8830);
nand U9244 (N_9244,N_9112,N_8894);
and U9245 (N_9245,N_9109,N_9153);
or U9246 (N_9246,N_8807,N_8847);
nor U9247 (N_9247,N_9008,N_8957);
nor U9248 (N_9248,N_8803,N_8987);
xnor U9249 (N_9249,N_8950,N_8967);
nor U9250 (N_9250,N_8909,N_9122);
and U9251 (N_9251,N_9029,N_9147);
nor U9252 (N_9252,N_9098,N_9006);
nand U9253 (N_9253,N_8871,N_8823);
or U9254 (N_9254,N_8805,N_9065);
nor U9255 (N_9255,N_9110,N_8856);
nand U9256 (N_9256,N_9182,N_8971);
nand U9257 (N_9257,N_9130,N_9095);
nor U9258 (N_9258,N_8932,N_8942);
and U9259 (N_9259,N_9128,N_9199);
and U9260 (N_9260,N_8886,N_9089);
or U9261 (N_9261,N_9016,N_9037);
or U9262 (N_9262,N_8915,N_9158);
nor U9263 (N_9263,N_9117,N_9108);
and U9264 (N_9264,N_9120,N_9084);
nor U9265 (N_9265,N_8889,N_8844);
nand U9266 (N_9266,N_8985,N_8853);
nor U9267 (N_9267,N_8954,N_8905);
nand U9268 (N_9268,N_9103,N_9165);
and U9269 (N_9269,N_8842,N_8992);
xor U9270 (N_9270,N_9176,N_8892);
and U9271 (N_9271,N_9184,N_9067);
and U9272 (N_9272,N_8914,N_8891);
or U9273 (N_9273,N_9043,N_8863);
nor U9274 (N_9274,N_8854,N_9133);
or U9275 (N_9275,N_9146,N_8920);
nand U9276 (N_9276,N_8825,N_8820);
nand U9277 (N_9277,N_8861,N_8926);
or U9278 (N_9278,N_8874,N_8858);
and U9279 (N_9279,N_9156,N_8826);
xnor U9280 (N_9280,N_8867,N_8872);
nor U9281 (N_9281,N_8964,N_9118);
nand U9282 (N_9282,N_9097,N_9060);
nor U9283 (N_9283,N_9093,N_8965);
nor U9284 (N_9284,N_9160,N_9068);
and U9285 (N_9285,N_8962,N_9107);
or U9286 (N_9286,N_9017,N_8993);
and U9287 (N_9287,N_8875,N_9022);
nand U9288 (N_9288,N_9009,N_9058);
and U9289 (N_9289,N_9002,N_9123);
nor U9290 (N_9290,N_9078,N_8982);
or U9291 (N_9291,N_9012,N_8959);
or U9292 (N_9292,N_9061,N_9054);
and U9293 (N_9293,N_9088,N_8913);
and U9294 (N_9294,N_8890,N_8845);
nand U9295 (N_9295,N_8851,N_8841);
nand U9296 (N_9296,N_8974,N_9053);
nand U9297 (N_9297,N_9192,N_9137);
or U9298 (N_9298,N_8990,N_8961);
and U9299 (N_9299,N_9000,N_9094);
and U9300 (N_9300,N_9086,N_9186);
nand U9301 (N_9301,N_9187,N_9191);
or U9302 (N_9302,N_9148,N_9119);
nand U9303 (N_9303,N_9040,N_9140);
nand U9304 (N_9304,N_8819,N_8860);
or U9305 (N_9305,N_9196,N_9091);
or U9306 (N_9306,N_9030,N_8810);
and U9307 (N_9307,N_9048,N_8981);
and U9308 (N_9308,N_9066,N_8996);
and U9309 (N_9309,N_9106,N_8876);
nor U9310 (N_9310,N_8850,N_8994);
nand U9311 (N_9311,N_8804,N_9027);
nand U9312 (N_9312,N_9001,N_9100);
nor U9313 (N_9313,N_9129,N_9104);
xor U9314 (N_9314,N_8800,N_9127);
or U9315 (N_9315,N_9011,N_9047);
nand U9316 (N_9316,N_9151,N_8917);
nand U9317 (N_9317,N_9092,N_9173);
nor U9318 (N_9318,N_8829,N_9139);
nand U9319 (N_9319,N_8918,N_9004);
nand U9320 (N_9320,N_8979,N_9114);
nor U9321 (N_9321,N_8973,N_8969);
xor U9322 (N_9322,N_9134,N_8999);
or U9323 (N_9323,N_8924,N_9057);
nor U9324 (N_9324,N_9175,N_9062);
and U9325 (N_9325,N_9025,N_8988);
and U9326 (N_9326,N_9039,N_9190);
nor U9327 (N_9327,N_8888,N_9021);
nor U9328 (N_9328,N_8901,N_8937);
or U9329 (N_9329,N_9161,N_9116);
or U9330 (N_9330,N_9085,N_8958);
and U9331 (N_9331,N_9013,N_8801);
nor U9332 (N_9332,N_8859,N_9075);
nand U9333 (N_9333,N_9083,N_9072);
nand U9334 (N_9334,N_8911,N_8910);
or U9335 (N_9335,N_8848,N_9135);
xor U9336 (N_9336,N_8837,N_8939);
or U9337 (N_9337,N_9033,N_9071);
nand U9338 (N_9338,N_9005,N_9090);
or U9339 (N_9339,N_9105,N_8972);
nand U9340 (N_9340,N_8966,N_8849);
and U9341 (N_9341,N_9031,N_8885);
and U9342 (N_9342,N_9155,N_9045);
nand U9343 (N_9343,N_9166,N_8970);
nand U9344 (N_9344,N_9121,N_8869);
or U9345 (N_9345,N_8865,N_9007);
nand U9346 (N_9346,N_9082,N_8976);
or U9347 (N_9347,N_8839,N_9159);
nand U9348 (N_9348,N_8833,N_8943);
nor U9349 (N_9349,N_9144,N_8834);
nor U9350 (N_9350,N_8940,N_8989);
or U9351 (N_9351,N_8887,N_9188);
and U9352 (N_9352,N_9024,N_8948);
nor U9353 (N_9353,N_8821,N_9154);
or U9354 (N_9354,N_9010,N_9046);
or U9355 (N_9355,N_9080,N_9157);
nor U9356 (N_9356,N_8953,N_8802);
nand U9357 (N_9357,N_9174,N_8912);
and U9358 (N_9358,N_9185,N_9143);
and U9359 (N_9359,N_8941,N_9018);
nand U9360 (N_9360,N_9051,N_8893);
nor U9361 (N_9361,N_9164,N_9052);
and U9362 (N_9362,N_9014,N_9126);
or U9363 (N_9363,N_8998,N_8813);
nand U9364 (N_9364,N_8846,N_8857);
and U9365 (N_9365,N_8907,N_8934);
or U9366 (N_9366,N_9034,N_9177);
or U9367 (N_9367,N_9172,N_8980);
nor U9368 (N_9368,N_9138,N_8983);
and U9369 (N_9369,N_9019,N_8997);
and U9370 (N_9370,N_8919,N_9069);
xnor U9371 (N_9371,N_9198,N_8814);
nand U9372 (N_9372,N_8938,N_8895);
nand U9373 (N_9373,N_9099,N_9170);
or U9374 (N_9374,N_8933,N_9064);
nor U9375 (N_9375,N_8880,N_9020);
nand U9376 (N_9376,N_8968,N_8817);
nor U9377 (N_9377,N_8896,N_8984);
or U9378 (N_9378,N_9189,N_8960);
nand U9379 (N_9379,N_9152,N_8922);
or U9380 (N_9380,N_8832,N_9163);
and U9381 (N_9381,N_8828,N_9042);
nor U9382 (N_9382,N_8991,N_9136);
or U9383 (N_9383,N_9195,N_8868);
nand U9384 (N_9384,N_9073,N_8838);
nand U9385 (N_9385,N_9049,N_8906);
nand U9386 (N_9386,N_8881,N_9181);
and U9387 (N_9387,N_9125,N_8812);
or U9388 (N_9388,N_8883,N_9096);
nand U9389 (N_9389,N_8928,N_8870);
nor U9390 (N_9390,N_9131,N_8811);
and U9391 (N_9391,N_9056,N_9171);
nand U9392 (N_9392,N_8824,N_8884);
or U9393 (N_9393,N_8816,N_8947);
and U9394 (N_9394,N_9032,N_9050);
nand U9395 (N_9395,N_9124,N_8995);
or U9396 (N_9396,N_8818,N_9168);
and U9397 (N_9397,N_8946,N_8949);
nand U9398 (N_9398,N_8986,N_9167);
and U9399 (N_9399,N_9038,N_9079);
and U9400 (N_9400,N_9190,N_8878);
or U9401 (N_9401,N_8891,N_8812);
nor U9402 (N_9402,N_9064,N_9082);
or U9403 (N_9403,N_9114,N_8926);
nand U9404 (N_9404,N_8860,N_9167);
nand U9405 (N_9405,N_9177,N_8878);
or U9406 (N_9406,N_9106,N_9167);
nand U9407 (N_9407,N_8950,N_8911);
and U9408 (N_9408,N_9178,N_8804);
nand U9409 (N_9409,N_8957,N_8866);
nor U9410 (N_9410,N_9027,N_8882);
or U9411 (N_9411,N_9171,N_8883);
nand U9412 (N_9412,N_8812,N_9106);
nor U9413 (N_9413,N_8898,N_9125);
nor U9414 (N_9414,N_9061,N_9164);
nand U9415 (N_9415,N_8819,N_8813);
nor U9416 (N_9416,N_8916,N_9193);
or U9417 (N_9417,N_9104,N_9000);
or U9418 (N_9418,N_8878,N_8856);
nor U9419 (N_9419,N_9093,N_8867);
or U9420 (N_9420,N_9059,N_9110);
or U9421 (N_9421,N_9100,N_8850);
and U9422 (N_9422,N_8900,N_8846);
nor U9423 (N_9423,N_8877,N_9039);
nand U9424 (N_9424,N_8824,N_9022);
nand U9425 (N_9425,N_9030,N_9053);
and U9426 (N_9426,N_9076,N_8944);
nand U9427 (N_9427,N_9081,N_8885);
nand U9428 (N_9428,N_9169,N_8952);
or U9429 (N_9429,N_9109,N_9041);
nand U9430 (N_9430,N_8809,N_9041);
or U9431 (N_9431,N_9008,N_9103);
nand U9432 (N_9432,N_8839,N_8880);
and U9433 (N_9433,N_9086,N_9029);
or U9434 (N_9434,N_9126,N_9194);
and U9435 (N_9435,N_9075,N_9144);
or U9436 (N_9436,N_9018,N_8818);
or U9437 (N_9437,N_8835,N_9021);
and U9438 (N_9438,N_9021,N_8852);
and U9439 (N_9439,N_9139,N_9180);
nand U9440 (N_9440,N_8949,N_8814);
nor U9441 (N_9441,N_8811,N_8862);
and U9442 (N_9442,N_9038,N_8849);
nor U9443 (N_9443,N_9163,N_8871);
nand U9444 (N_9444,N_9115,N_8914);
and U9445 (N_9445,N_9174,N_8961);
and U9446 (N_9446,N_8868,N_8946);
nand U9447 (N_9447,N_8947,N_8924);
or U9448 (N_9448,N_8995,N_9119);
nand U9449 (N_9449,N_8867,N_8909);
nor U9450 (N_9450,N_9038,N_9136);
nand U9451 (N_9451,N_9182,N_8951);
or U9452 (N_9452,N_8832,N_9125);
nor U9453 (N_9453,N_9075,N_9198);
nor U9454 (N_9454,N_9159,N_8817);
and U9455 (N_9455,N_9027,N_8868);
or U9456 (N_9456,N_8944,N_9077);
nand U9457 (N_9457,N_8853,N_8877);
nor U9458 (N_9458,N_9042,N_9141);
nor U9459 (N_9459,N_8996,N_9010);
nand U9460 (N_9460,N_8863,N_9026);
or U9461 (N_9461,N_9175,N_9079);
or U9462 (N_9462,N_9091,N_8848);
nor U9463 (N_9463,N_8924,N_8919);
nand U9464 (N_9464,N_9091,N_8896);
nor U9465 (N_9465,N_8834,N_9071);
and U9466 (N_9466,N_9014,N_9016);
nand U9467 (N_9467,N_8823,N_9175);
nor U9468 (N_9468,N_9064,N_8911);
nand U9469 (N_9469,N_9044,N_8867);
and U9470 (N_9470,N_9001,N_8833);
nor U9471 (N_9471,N_9033,N_8882);
nand U9472 (N_9472,N_9097,N_8837);
and U9473 (N_9473,N_9103,N_8829);
and U9474 (N_9474,N_9072,N_9091);
nor U9475 (N_9475,N_9040,N_8914);
nand U9476 (N_9476,N_8967,N_9027);
and U9477 (N_9477,N_9135,N_9157);
nor U9478 (N_9478,N_8934,N_9199);
or U9479 (N_9479,N_8962,N_9128);
and U9480 (N_9480,N_8804,N_8867);
or U9481 (N_9481,N_8916,N_8860);
nand U9482 (N_9482,N_8949,N_9079);
nor U9483 (N_9483,N_9029,N_9089);
and U9484 (N_9484,N_9007,N_8986);
and U9485 (N_9485,N_9016,N_8845);
or U9486 (N_9486,N_9022,N_9010);
nand U9487 (N_9487,N_9171,N_8936);
nor U9488 (N_9488,N_8829,N_9075);
nor U9489 (N_9489,N_9002,N_8949);
nand U9490 (N_9490,N_9105,N_9045);
or U9491 (N_9491,N_9098,N_9152);
and U9492 (N_9492,N_8928,N_8903);
or U9493 (N_9493,N_9134,N_8958);
and U9494 (N_9494,N_8864,N_9098);
nand U9495 (N_9495,N_8804,N_9022);
and U9496 (N_9496,N_8864,N_8850);
nand U9497 (N_9497,N_8929,N_8836);
nor U9498 (N_9498,N_9025,N_8928);
nand U9499 (N_9499,N_9050,N_8889);
nor U9500 (N_9500,N_9023,N_8845);
or U9501 (N_9501,N_9131,N_8996);
or U9502 (N_9502,N_8965,N_9024);
nand U9503 (N_9503,N_8888,N_8832);
and U9504 (N_9504,N_8877,N_9073);
nor U9505 (N_9505,N_9132,N_9107);
and U9506 (N_9506,N_9144,N_9108);
nor U9507 (N_9507,N_9011,N_8952);
and U9508 (N_9508,N_8945,N_8887);
or U9509 (N_9509,N_8971,N_9021);
nand U9510 (N_9510,N_8978,N_9145);
nand U9511 (N_9511,N_9130,N_8868);
and U9512 (N_9512,N_9193,N_8866);
and U9513 (N_9513,N_9006,N_9177);
and U9514 (N_9514,N_8830,N_9170);
nor U9515 (N_9515,N_8878,N_8945);
and U9516 (N_9516,N_8856,N_8885);
and U9517 (N_9517,N_8896,N_8999);
nor U9518 (N_9518,N_9192,N_8949);
and U9519 (N_9519,N_9154,N_8830);
or U9520 (N_9520,N_8942,N_8955);
xnor U9521 (N_9521,N_9049,N_8915);
nand U9522 (N_9522,N_9060,N_9115);
nand U9523 (N_9523,N_9175,N_8898);
nor U9524 (N_9524,N_9109,N_8812);
and U9525 (N_9525,N_8813,N_9166);
and U9526 (N_9526,N_9170,N_8987);
nand U9527 (N_9527,N_8973,N_9111);
nor U9528 (N_9528,N_9141,N_8814);
or U9529 (N_9529,N_9029,N_8832);
nor U9530 (N_9530,N_8901,N_8941);
nor U9531 (N_9531,N_8818,N_8977);
nand U9532 (N_9532,N_8929,N_9073);
nor U9533 (N_9533,N_8951,N_8815);
and U9534 (N_9534,N_9099,N_9064);
nor U9535 (N_9535,N_8907,N_8975);
or U9536 (N_9536,N_9059,N_8888);
and U9537 (N_9537,N_9128,N_9042);
nand U9538 (N_9538,N_8930,N_9098);
or U9539 (N_9539,N_9096,N_9127);
and U9540 (N_9540,N_9032,N_9097);
nand U9541 (N_9541,N_8880,N_9006);
and U9542 (N_9542,N_8928,N_9108);
or U9543 (N_9543,N_9018,N_8802);
nand U9544 (N_9544,N_9198,N_8900);
and U9545 (N_9545,N_8893,N_9112);
nor U9546 (N_9546,N_8842,N_9016);
nor U9547 (N_9547,N_9023,N_8877);
nor U9548 (N_9548,N_8851,N_9143);
and U9549 (N_9549,N_9148,N_9103);
or U9550 (N_9550,N_8986,N_8956);
xor U9551 (N_9551,N_9071,N_9075);
and U9552 (N_9552,N_8884,N_9106);
and U9553 (N_9553,N_9085,N_8844);
and U9554 (N_9554,N_9109,N_8995);
nor U9555 (N_9555,N_9156,N_9044);
or U9556 (N_9556,N_8869,N_9044);
nor U9557 (N_9557,N_9162,N_8965);
nor U9558 (N_9558,N_8996,N_9182);
and U9559 (N_9559,N_8879,N_9066);
xor U9560 (N_9560,N_9140,N_8866);
nor U9561 (N_9561,N_9133,N_8891);
and U9562 (N_9562,N_9026,N_9197);
nand U9563 (N_9563,N_8882,N_8990);
or U9564 (N_9564,N_8975,N_9159);
nand U9565 (N_9565,N_9148,N_9009);
nand U9566 (N_9566,N_9186,N_8919);
nand U9567 (N_9567,N_9168,N_8988);
nor U9568 (N_9568,N_9185,N_9060);
or U9569 (N_9569,N_8907,N_9024);
nor U9570 (N_9570,N_8911,N_9120);
or U9571 (N_9571,N_9196,N_9148);
and U9572 (N_9572,N_9004,N_8801);
nor U9573 (N_9573,N_8956,N_9134);
or U9574 (N_9574,N_9161,N_9003);
nand U9575 (N_9575,N_8804,N_8936);
and U9576 (N_9576,N_8955,N_8876);
nand U9577 (N_9577,N_8950,N_9184);
nor U9578 (N_9578,N_9061,N_9127);
and U9579 (N_9579,N_8917,N_9091);
nand U9580 (N_9580,N_9003,N_8851);
nor U9581 (N_9581,N_9040,N_9063);
or U9582 (N_9582,N_9027,N_9182);
nor U9583 (N_9583,N_8853,N_9078);
and U9584 (N_9584,N_8810,N_9149);
nand U9585 (N_9585,N_9183,N_8980);
and U9586 (N_9586,N_8870,N_9032);
and U9587 (N_9587,N_8916,N_9088);
nor U9588 (N_9588,N_9106,N_9022);
or U9589 (N_9589,N_8949,N_9038);
or U9590 (N_9590,N_9103,N_9044);
and U9591 (N_9591,N_8856,N_9086);
or U9592 (N_9592,N_8844,N_9084);
and U9593 (N_9593,N_8854,N_9182);
nor U9594 (N_9594,N_9007,N_9182);
and U9595 (N_9595,N_8866,N_9076);
nand U9596 (N_9596,N_8877,N_8892);
or U9597 (N_9597,N_8901,N_9152);
nor U9598 (N_9598,N_9173,N_9011);
nand U9599 (N_9599,N_8964,N_9126);
or U9600 (N_9600,N_9446,N_9426);
or U9601 (N_9601,N_9314,N_9254);
and U9602 (N_9602,N_9396,N_9533);
or U9603 (N_9603,N_9264,N_9500);
nand U9604 (N_9604,N_9481,N_9403);
or U9605 (N_9605,N_9432,N_9453);
or U9606 (N_9606,N_9351,N_9469);
or U9607 (N_9607,N_9245,N_9413);
nand U9608 (N_9608,N_9544,N_9408);
nor U9609 (N_9609,N_9480,N_9369);
and U9610 (N_9610,N_9231,N_9423);
nand U9611 (N_9611,N_9447,N_9411);
nor U9612 (N_9612,N_9315,N_9506);
nand U9613 (N_9613,N_9491,N_9294);
or U9614 (N_9614,N_9508,N_9206);
and U9615 (N_9615,N_9329,N_9594);
or U9616 (N_9616,N_9399,N_9363);
nand U9617 (N_9617,N_9402,N_9542);
nand U9618 (N_9618,N_9452,N_9581);
or U9619 (N_9619,N_9551,N_9285);
or U9620 (N_9620,N_9289,N_9582);
and U9621 (N_9621,N_9256,N_9203);
nand U9622 (N_9622,N_9407,N_9400);
and U9623 (N_9623,N_9472,N_9483);
nand U9624 (N_9624,N_9205,N_9416);
nor U9625 (N_9625,N_9317,N_9441);
nand U9626 (N_9626,N_9507,N_9489);
or U9627 (N_9627,N_9252,N_9553);
nor U9628 (N_9628,N_9589,N_9577);
or U9629 (N_9629,N_9377,N_9342);
or U9630 (N_9630,N_9211,N_9295);
and U9631 (N_9631,N_9232,N_9296);
or U9632 (N_9632,N_9283,N_9328);
and U9633 (N_9633,N_9558,N_9379);
and U9634 (N_9634,N_9515,N_9404);
nand U9635 (N_9635,N_9521,N_9485);
or U9636 (N_9636,N_9534,N_9345);
nand U9637 (N_9637,N_9478,N_9234);
and U9638 (N_9638,N_9561,N_9456);
nor U9639 (N_9639,N_9536,N_9299);
nand U9640 (N_9640,N_9312,N_9214);
nand U9641 (N_9641,N_9380,N_9444);
nand U9642 (N_9642,N_9414,N_9578);
nand U9643 (N_9643,N_9307,N_9219);
nor U9644 (N_9644,N_9431,N_9383);
nand U9645 (N_9645,N_9512,N_9367);
or U9646 (N_9646,N_9261,N_9430);
or U9647 (N_9647,N_9488,N_9236);
nand U9648 (N_9648,N_9286,N_9373);
or U9649 (N_9649,N_9549,N_9409);
nor U9650 (N_9650,N_9398,N_9424);
and U9651 (N_9651,N_9226,N_9439);
nor U9652 (N_9652,N_9209,N_9579);
nand U9653 (N_9653,N_9279,N_9591);
nor U9654 (N_9654,N_9248,N_9401);
and U9655 (N_9655,N_9548,N_9576);
xor U9656 (N_9656,N_9498,N_9352);
nand U9657 (N_9657,N_9525,N_9545);
nand U9658 (N_9658,N_9273,N_9266);
or U9659 (N_9659,N_9280,N_9514);
and U9660 (N_9660,N_9204,N_9599);
and U9661 (N_9661,N_9490,N_9249);
and U9662 (N_9662,N_9465,N_9572);
or U9663 (N_9663,N_9215,N_9223);
and U9664 (N_9664,N_9596,N_9366);
nor U9665 (N_9665,N_9332,N_9437);
or U9666 (N_9666,N_9590,N_9271);
and U9667 (N_9667,N_9301,N_9371);
and U9668 (N_9668,N_9201,N_9421);
xor U9669 (N_9669,N_9537,N_9356);
or U9670 (N_9670,N_9334,N_9584);
or U9671 (N_9671,N_9550,N_9365);
nand U9672 (N_9672,N_9524,N_9208);
or U9673 (N_9673,N_9540,N_9461);
or U9674 (N_9674,N_9547,N_9517);
nor U9675 (N_9675,N_9422,N_9381);
nand U9676 (N_9676,N_9598,N_9333);
and U9677 (N_9677,N_9360,N_9346);
nor U9678 (N_9678,N_9392,N_9355);
and U9679 (N_9679,N_9238,N_9412);
nand U9680 (N_9680,N_9291,N_9348);
nand U9681 (N_9681,N_9418,N_9393);
nand U9682 (N_9682,N_9313,N_9493);
nor U9683 (N_9683,N_9270,N_9224);
and U9684 (N_9684,N_9405,N_9257);
nor U9685 (N_9685,N_9523,N_9428);
or U9686 (N_9686,N_9565,N_9511);
nand U9687 (N_9687,N_9425,N_9323);
and U9688 (N_9688,N_9237,N_9258);
nor U9689 (N_9689,N_9319,N_9557);
or U9690 (N_9690,N_9504,N_9267);
or U9691 (N_9691,N_9388,N_9357);
or U9692 (N_9692,N_9494,N_9477);
xnor U9693 (N_9693,N_9281,N_9353);
nand U9694 (N_9694,N_9415,N_9499);
nand U9695 (N_9695,N_9250,N_9420);
nand U9696 (N_9696,N_9336,N_9435);
and U9697 (N_9697,N_9560,N_9530);
or U9698 (N_9698,N_9220,N_9592);
and U9699 (N_9699,N_9227,N_9510);
or U9700 (N_9700,N_9397,N_9559);
or U9701 (N_9701,N_9454,N_9362);
nand U9702 (N_9702,N_9538,N_9391);
nor U9703 (N_9703,N_9484,N_9298);
and U9704 (N_9704,N_9513,N_9337);
nand U9705 (N_9705,N_9569,N_9546);
or U9706 (N_9706,N_9574,N_9450);
or U9707 (N_9707,N_9496,N_9320);
and U9708 (N_9708,N_9364,N_9374);
nor U9709 (N_9709,N_9288,N_9567);
nand U9710 (N_9710,N_9275,N_9570);
nand U9711 (N_9711,N_9247,N_9361);
nand U9712 (N_9712,N_9233,N_9274);
and U9713 (N_9713,N_9330,N_9466);
nand U9714 (N_9714,N_9390,N_9468);
or U9715 (N_9715,N_9573,N_9503);
nand U9716 (N_9716,N_9442,N_9293);
nand U9717 (N_9717,N_9242,N_9476);
nor U9718 (N_9718,N_9229,N_9529);
nor U9719 (N_9719,N_9427,N_9554);
and U9720 (N_9720,N_9230,N_9213);
nand U9721 (N_9721,N_9518,N_9309);
or U9722 (N_9722,N_9308,N_9327);
and U9723 (N_9723,N_9376,N_9335);
or U9724 (N_9724,N_9482,N_9520);
or U9725 (N_9725,N_9338,N_9262);
and U9726 (N_9726,N_9445,N_9585);
and U9727 (N_9727,N_9277,N_9359);
nand U9728 (N_9728,N_9474,N_9304);
and U9729 (N_9729,N_9593,N_9265);
xnor U9730 (N_9730,N_9539,N_9516);
nand U9731 (N_9731,N_9222,N_9470);
nand U9732 (N_9732,N_9487,N_9386);
or U9733 (N_9733,N_9349,N_9458);
nor U9734 (N_9734,N_9475,N_9527);
nand U9735 (N_9735,N_9406,N_9419);
nor U9736 (N_9736,N_9325,N_9410);
and U9737 (N_9737,N_9519,N_9322);
or U9738 (N_9738,N_9316,N_9350);
nand U9739 (N_9739,N_9347,N_9340);
or U9740 (N_9740,N_9240,N_9448);
or U9741 (N_9741,N_9455,N_9278);
xnor U9742 (N_9742,N_9387,N_9532);
nor U9743 (N_9743,N_9246,N_9394);
or U9744 (N_9744,N_9341,N_9210);
nand U9745 (N_9745,N_9339,N_9241);
and U9746 (N_9746,N_9300,N_9378);
or U9747 (N_9747,N_9251,N_9492);
nor U9748 (N_9748,N_9225,N_9479);
or U9749 (N_9749,N_9228,N_9526);
and U9750 (N_9750,N_9505,N_9311);
nor U9751 (N_9751,N_9429,N_9384);
and U9752 (N_9752,N_9575,N_9436);
and U9753 (N_9753,N_9284,N_9568);
nor U9754 (N_9754,N_9276,N_9541);
nor U9755 (N_9755,N_9358,N_9297);
and U9756 (N_9756,N_9268,N_9372);
and U9757 (N_9757,N_9566,N_9321);
nor U9758 (N_9758,N_9287,N_9221);
nand U9759 (N_9759,N_9306,N_9259);
nor U9760 (N_9760,N_9449,N_9556);
and U9761 (N_9761,N_9260,N_9462);
nor U9762 (N_9762,N_9310,N_9202);
nor U9763 (N_9763,N_9459,N_9235);
nand U9764 (N_9764,N_9486,N_9451);
nor U9765 (N_9765,N_9443,N_9272);
nand U9766 (N_9766,N_9555,N_9562);
nor U9767 (N_9767,N_9344,N_9433);
nor U9768 (N_9768,N_9588,N_9324);
or U9769 (N_9769,N_9263,N_9467);
nand U9770 (N_9770,N_9583,N_9326);
nand U9771 (N_9771,N_9244,N_9382);
nor U9772 (N_9772,N_9586,N_9501);
and U9773 (N_9773,N_9563,N_9571);
nand U9774 (N_9774,N_9552,N_9255);
nor U9775 (N_9775,N_9463,N_9522);
and U9776 (N_9776,N_9587,N_9389);
nor U9777 (N_9777,N_9354,N_9217);
nand U9778 (N_9778,N_9303,N_9595);
or U9779 (N_9779,N_9302,N_9495);
or U9780 (N_9780,N_9218,N_9375);
nor U9781 (N_9781,N_9343,N_9543);
nor U9782 (N_9782,N_9434,N_9216);
or U9783 (N_9783,N_9531,N_9253);
and U9784 (N_9784,N_9580,N_9207);
nand U9785 (N_9785,N_9385,N_9471);
nor U9786 (N_9786,N_9597,N_9212);
or U9787 (N_9787,N_9368,N_9464);
and U9788 (N_9788,N_9282,N_9239);
nand U9789 (N_9789,N_9395,N_9269);
or U9790 (N_9790,N_9292,N_9535);
nand U9791 (N_9791,N_9243,N_9564);
or U9792 (N_9792,N_9318,N_9457);
or U9793 (N_9793,N_9460,N_9200);
or U9794 (N_9794,N_9440,N_9370);
nor U9795 (N_9795,N_9509,N_9290);
and U9796 (N_9796,N_9473,N_9438);
or U9797 (N_9797,N_9497,N_9502);
and U9798 (N_9798,N_9528,N_9331);
nor U9799 (N_9799,N_9305,N_9417);
nand U9800 (N_9800,N_9372,N_9218);
nor U9801 (N_9801,N_9296,N_9441);
or U9802 (N_9802,N_9403,N_9557);
nor U9803 (N_9803,N_9584,N_9393);
nand U9804 (N_9804,N_9525,N_9520);
nor U9805 (N_9805,N_9516,N_9594);
or U9806 (N_9806,N_9245,N_9335);
and U9807 (N_9807,N_9313,N_9430);
nor U9808 (N_9808,N_9237,N_9248);
and U9809 (N_9809,N_9521,N_9404);
or U9810 (N_9810,N_9583,N_9229);
nand U9811 (N_9811,N_9445,N_9448);
or U9812 (N_9812,N_9329,N_9457);
or U9813 (N_9813,N_9591,N_9289);
and U9814 (N_9814,N_9530,N_9390);
and U9815 (N_9815,N_9355,N_9317);
or U9816 (N_9816,N_9406,N_9353);
or U9817 (N_9817,N_9454,N_9449);
nand U9818 (N_9818,N_9358,N_9235);
or U9819 (N_9819,N_9580,N_9524);
and U9820 (N_9820,N_9238,N_9203);
nand U9821 (N_9821,N_9430,N_9409);
nand U9822 (N_9822,N_9244,N_9432);
nor U9823 (N_9823,N_9467,N_9337);
nor U9824 (N_9824,N_9335,N_9569);
nor U9825 (N_9825,N_9514,N_9583);
or U9826 (N_9826,N_9525,N_9547);
and U9827 (N_9827,N_9245,N_9536);
and U9828 (N_9828,N_9534,N_9331);
and U9829 (N_9829,N_9532,N_9295);
nor U9830 (N_9830,N_9516,N_9277);
nand U9831 (N_9831,N_9319,N_9515);
and U9832 (N_9832,N_9509,N_9446);
nand U9833 (N_9833,N_9568,N_9337);
nand U9834 (N_9834,N_9258,N_9228);
or U9835 (N_9835,N_9321,N_9390);
and U9836 (N_9836,N_9499,N_9246);
or U9837 (N_9837,N_9543,N_9442);
or U9838 (N_9838,N_9566,N_9269);
or U9839 (N_9839,N_9200,N_9516);
or U9840 (N_9840,N_9365,N_9338);
nor U9841 (N_9841,N_9216,N_9396);
and U9842 (N_9842,N_9597,N_9577);
nand U9843 (N_9843,N_9411,N_9262);
and U9844 (N_9844,N_9216,N_9416);
or U9845 (N_9845,N_9333,N_9484);
nand U9846 (N_9846,N_9405,N_9547);
nand U9847 (N_9847,N_9547,N_9266);
nor U9848 (N_9848,N_9258,N_9269);
nand U9849 (N_9849,N_9339,N_9383);
nor U9850 (N_9850,N_9344,N_9384);
or U9851 (N_9851,N_9599,N_9314);
or U9852 (N_9852,N_9569,N_9536);
and U9853 (N_9853,N_9204,N_9314);
nor U9854 (N_9854,N_9599,N_9372);
nor U9855 (N_9855,N_9383,N_9422);
and U9856 (N_9856,N_9282,N_9478);
nor U9857 (N_9857,N_9563,N_9351);
or U9858 (N_9858,N_9431,N_9305);
or U9859 (N_9859,N_9530,N_9311);
or U9860 (N_9860,N_9545,N_9491);
nor U9861 (N_9861,N_9477,N_9218);
nand U9862 (N_9862,N_9502,N_9553);
nor U9863 (N_9863,N_9335,N_9476);
nand U9864 (N_9864,N_9589,N_9455);
or U9865 (N_9865,N_9367,N_9318);
or U9866 (N_9866,N_9359,N_9347);
nand U9867 (N_9867,N_9249,N_9598);
or U9868 (N_9868,N_9524,N_9430);
nor U9869 (N_9869,N_9569,N_9329);
nand U9870 (N_9870,N_9310,N_9245);
nor U9871 (N_9871,N_9212,N_9353);
and U9872 (N_9872,N_9291,N_9507);
nor U9873 (N_9873,N_9536,N_9580);
or U9874 (N_9874,N_9252,N_9340);
or U9875 (N_9875,N_9252,N_9271);
and U9876 (N_9876,N_9486,N_9568);
or U9877 (N_9877,N_9566,N_9418);
and U9878 (N_9878,N_9498,N_9231);
nor U9879 (N_9879,N_9567,N_9448);
nor U9880 (N_9880,N_9429,N_9587);
nor U9881 (N_9881,N_9223,N_9561);
nor U9882 (N_9882,N_9308,N_9247);
nand U9883 (N_9883,N_9366,N_9257);
nor U9884 (N_9884,N_9595,N_9252);
nand U9885 (N_9885,N_9327,N_9455);
and U9886 (N_9886,N_9313,N_9377);
or U9887 (N_9887,N_9587,N_9483);
or U9888 (N_9888,N_9222,N_9418);
xor U9889 (N_9889,N_9480,N_9539);
or U9890 (N_9890,N_9595,N_9578);
and U9891 (N_9891,N_9530,N_9445);
or U9892 (N_9892,N_9359,N_9596);
nand U9893 (N_9893,N_9456,N_9560);
nor U9894 (N_9894,N_9359,N_9574);
and U9895 (N_9895,N_9263,N_9552);
nand U9896 (N_9896,N_9286,N_9337);
and U9897 (N_9897,N_9544,N_9491);
or U9898 (N_9898,N_9560,N_9282);
nand U9899 (N_9899,N_9352,N_9437);
or U9900 (N_9900,N_9544,N_9371);
or U9901 (N_9901,N_9333,N_9282);
or U9902 (N_9902,N_9594,N_9308);
or U9903 (N_9903,N_9396,N_9217);
and U9904 (N_9904,N_9372,N_9306);
nand U9905 (N_9905,N_9422,N_9432);
or U9906 (N_9906,N_9555,N_9328);
and U9907 (N_9907,N_9449,N_9246);
nand U9908 (N_9908,N_9349,N_9277);
nor U9909 (N_9909,N_9472,N_9547);
nor U9910 (N_9910,N_9387,N_9319);
and U9911 (N_9911,N_9313,N_9340);
nor U9912 (N_9912,N_9540,N_9310);
nor U9913 (N_9913,N_9410,N_9405);
nor U9914 (N_9914,N_9461,N_9586);
or U9915 (N_9915,N_9478,N_9470);
or U9916 (N_9916,N_9385,N_9556);
or U9917 (N_9917,N_9559,N_9264);
nand U9918 (N_9918,N_9246,N_9517);
nor U9919 (N_9919,N_9311,N_9271);
xor U9920 (N_9920,N_9345,N_9536);
or U9921 (N_9921,N_9270,N_9452);
and U9922 (N_9922,N_9476,N_9252);
nor U9923 (N_9923,N_9267,N_9241);
nor U9924 (N_9924,N_9405,N_9479);
or U9925 (N_9925,N_9385,N_9340);
nor U9926 (N_9926,N_9589,N_9466);
and U9927 (N_9927,N_9335,N_9222);
nand U9928 (N_9928,N_9490,N_9407);
or U9929 (N_9929,N_9537,N_9388);
nor U9930 (N_9930,N_9374,N_9386);
nand U9931 (N_9931,N_9496,N_9484);
or U9932 (N_9932,N_9375,N_9409);
or U9933 (N_9933,N_9367,N_9453);
and U9934 (N_9934,N_9288,N_9552);
nand U9935 (N_9935,N_9292,N_9520);
or U9936 (N_9936,N_9355,N_9420);
nand U9937 (N_9937,N_9506,N_9460);
nor U9938 (N_9938,N_9224,N_9307);
nor U9939 (N_9939,N_9304,N_9404);
or U9940 (N_9940,N_9457,N_9442);
or U9941 (N_9941,N_9509,N_9334);
and U9942 (N_9942,N_9243,N_9477);
or U9943 (N_9943,N_9263,N_9498);
nand U9944 (N_9944,N_9232,N_9461);
and U9945 (N_9945,N_9366,N_9537);
nand U9946 (N_9946,N_9329,N_9460);
and U9947 (N_9947,N_9287,N_9515);
or U9948 (N_9948,N_9579,N_9522);
xnor U9949 (N_9949,N_9449,N_9233);
nand U9950 (N_9950,N_9435,N_9566);
nor U9951 (N_9951,N_9200,N_9390);
or U9952 (N_9952,N_9598,N_9330);
and U9953 (N_9953,N_9208,N_9437);
or U9954 (N_9954,N_9542,N_9331);
nand U9955 (N_9955,N_9393,N_9262);
and U9956 (N_9956,N_9240,N_9338);
and U9957 (N_9957,N_9430,N_9541);
or U9958 (N_9958,N_9257,N_9468);
and U9959 (N_9959,N_9587,N_9294);
or U9960 (N_9960,N_9218,N_9343);
and U9961 (N_9961,N_9481,N_9375);
or U9962 (N_9962,N_9405,N_9219);
or U9963 (N_9963,N_9492,N_9263);
and U9964 (N_9964,N_9502,N_9257);
or U9965 (N_9965,N_9401,N_9543);
nor U9966 (N_9966,N_9234,N_9328);
nand U9967 (N_9967,N_9558,N_9425);
nor U9968 (N_9968,N_9574,N_9559);
nor U9969 (N_9969,N_9476,N_9504);
or U9970 (N_9970,N_9408,N_9493);
or U9971 (N_9971,N_9207,N_9442);
nand U9972 (N_9972,N_9244,N_9402);
nor U9973 (N_9973,N_9510,N_9562);
nor U9974 (N_9974,N_9292,N_9478);
nand U9975 (N_9975,N_9453,N_9211);
or U9976 (N_9976,N_9427,N_9215);
and U9977 (N_9977,N_9519,N_9241);
nor U9978 (N_9978,N_9301,N_9310);
or U9979 (N_9979,N_9505,N_9426);
and U9980 (N_9980,N_9442,N_9284);
nand U9981 (N_9981,N_9542,N_9442);
and U9982 (N_9982,N_9558,N_9578);
and U9983 (N_9983,N_9458,N_9412);
or U9984 (N_9984,N_9254,N_9214);
and U9985 (N_9985,N_9384,N_9557);
and U9986 (N_9986,N_9444,N_9324);
nand U9987 (N_9987,N_9410,N_9426);
nand U9988 (N_9988,N_9348,N_9240);
or U9989 (N_9989,N_9225,N_9376);
nor U9990 (N_9990,N_9249,N_9473);
nor U9991 (N_9991,N_9527,N_9242);
or U9992 (N_9992,N_9292,N_9388);
or U9993 (N_9993,N_9574,N_9473);
nor U9994 (N_9994,N_9398,N_9242);
and U9995 (N_9995,N_9525,N_9536);
or U9996 (N_9996,N_9354,N_9410);
nor U9997 (N_9997,N_9585,N_9284);
nor U9998 (N_9998,N_9236,N_9260);
or U9999 (N_9999,N_9404,N_9472);
nand U10000 (N_10000,N_9640,N_9768);
or U10001 (N_10001,N_9760,N_9748);
nand U10002 (N_10002,N_9743,N_9823);
nor U10003 (N_10003,N_9704,N_9687);
or U10004 (N_10004,N_9999,N_9624);
nor U10005 (N_10005,N_9930,N_9634);
or U10006 (N_10006,N_9706,N_9708);
or U10007 (N_10007,N_9792,N_9869);
nor U10008 (N_10008,N_9881,N_9899);
nor U10009 (N_10009,N_9826,N_9841);
and U10010 (N_10010,N_9829,N_9783);
and U10011 (N_10011,N_9987,N_9809);
nand U10012 (N_10012,N_9867,N_9749);
nor U10013 (N_10013,N_9682,N_9985);
nor U10014 (N_10014,N_9971,N_9794);
nand U10015 (N_10015,N_9834,N_9775);
and U10016 (N_10016,N_9996,N_9782);
nand U10017 (N_10017,N_9671,N_9645);
nand U10018 (N_10018,N_9931,N_9790);
or U10019 (N_10019,N_9769,N_9911);
nand U10020 (N_10020,N_9620,N_9946);
nor U10021 (N_10021,N_9913,N_9993);
or U10022 (N_10022,N_9844,N_9685);
and U10023 (N_10023,N_9968,N_9954);
and U10024 (N_10024,N_9811,N_9723);
nor U10025 (N_10025,N_9615,N_9952);
nor U10026 (N_10026,N_9644,N_9716);
and U10027 (N_10027,N_9733,N_9779);
nand U10028 (N_10028,N_9902,N_9746);
nand U10029 (N_10029,N_9653,N_9870);
or U10030 (N_10030,N_9879,N_9874);
nand U10031 (N_10031,N_9833,N_9859);
nor U10032 (N_10032,N_9614,N_9732);
nor U10033 (N_10033,N_9764,N_9835);
nand U10034 (N_10034,N_9681,N_9696);
nand U10035 (N_10035,N_9961,N_9621);
and U10036 (N_10036,N_9938,N_9808);
nor U10037 (N_10037,N_9991,N_9994);
and U10038 (N_10038,N_9857,N_9817);
and U10039 (N_10039,N_9969,N_9892);
nand U10040 (N_10040,N_9837,N_9876);
nand U10041 (N_10041,N_9639,N_9630);
nand U10042 (N_10042,N_9818,N_9658);
or U10043 (N_10043,N_9676,N_9607);
and U10044 (N_10044,N_9661,N_9830);
or U10045 (N_10045,N_9836,N_9997);
nand U10046 (N_10046,N_9988,N_9699);
or U10047 (N_10047,N_9788,N_9616);
or U10048 (N_10048,N_9942,N_9861);
or U10049 (N_10049,N_9939,N_9686);
and U10050 (N_10050,N_9774,N_9962);
or U10051 (N_10051,N_9669,N_9904);
nand U10052 (N_10052,N_9619,N_9893);
nand U10053 (N_10053,N_9872,N_9629);
nand U10054 (N_10054,N_9737,N_9878);
and U10055 (N_10055,N_9989,N_9649);
xnor U10056 (N_10056,N_9903,N_9995);
and U10057 (N_10057,N_9941,N_9928);
and U10058 (N_10058,N_9744,N_9868);
and U10059 (N_10059,N_9807,N_9670);
nand U10060 (N_10060,N_9672,N_9784);
nand U10061 (N_10061,N_9875,N_9683);
and U10062 (N_10062,N_9666,N_9828);
nand U10063 (N_10063,N_9650,N_9710);
nor U10064 (N_10064,N_9777,N_9771);
nand U10065 (N_10065,N_9780,N_9745);
and U10066 (N_10066,N_9973,N_9984);
or U10067 (N_10067,N_9883,N_9695);
nor U10068 (N_10068,N_9812,N_9885);
nor U10069 (N_10069,N_9786,N_9714);
nand U10070 (N_10070,N_9887,N_9998);
or U10071 (N_10071,N_9729,N_9724);
or U10072 (N_10072,N_9715,N_9785);
nor U10073 (N_10073,N_9776,N_9720);
and U10074 (N_10074,N_9947,N_9707);
or U10075 (N_10075,N_9647,N_9851);
nand U10076 (N_10076,N_9900,N_9896);
nand U10077 (N_10077,N_9909,N_9965);
and U10078 (N_10078,N_9719,N_9978);
nor U10079 (N_10079,N_9972,N_9943);
nand U10080 (N_10080,N_9901,N_9726);
or U10081 (N_10081,N_9605,N_9635);
nor U10082 (N_10082,N_9956,N_9798);
and U10083 (N_10083,N_9692,N_9960);
nand U10084 (N_10084,N_9934,N_9778);
and U10085 (N_10085,N_9608,N_9622);
and U10086 (N_10086,N_9871,N_9664);
nor U10087 (N_10087,N_9628,N_9923);
or U10088 (N_10088,N_9802,N_9637);
nor U10089 (N_10089,N_9839,N_9703);
and U10090 (N_10090,N_9898,N_9945);
or U10091 (N_10091,N_9684,N_9843);
nor U10092 (N_10092,N_9757,N_9814);
nor U10093 (N_10093,N_9625,N_9915);
nor U10094 (N_10094,N_9604,N_9747);
or U10095 (N_10095,N_9983,N_9709);
and U10096 (N_10096,N_9611,N_9966);
nor U10097 (N_10097,N_9753,N_9977);
and U10098 (N_10098,N_9789,N_9717);
nor U10099 (N_10099,N_9854,N_9980);
and U10100 (N_10100,N_9602,N_9662);
nor U10101 (N_10101,N_9958,N_9705);
nand U10102 (N_10102,N_9617,N_9722);
or U10103 (N_10103,N_9765,N_9797);
nand U10104 (N_10104,N_9950,N_9725);
and U10105 (N_10105,N_9643,N_9754);
or U10106 (N_10106,N_9654,N_9813);
and U10107 (N_10107,N_9642,N_9603);
or U10108 (N_10108,N_9949,N_9912);
and U10109 (N_10109,N_9741,N_9601);
or U10110 (N_10110,N_9986,N_9927);
and U10111 (N_10111,N_9819,N_9713);
and U10112 (N_10112,N_9990,N_9890);
or U10113 (N_10113,N_9825,N_9940);
and U10114 (N_10114,N_9652,N_9667);
nor U10115 (N_10115,N_9690,N_9679);
nor U10116 (N_10116,N_9755,N_9711);
or U10117 (N_10117,N_9860,N_9751);
nor U10118 (N_10118,N_9728,N_9864);
and U10119 (N_10119,N_9816,N_9845);
and U10120 (N_10120,N_9739,N_9668);
and U10121 (N_10121,N_9659,N_9894);
nor U10122 (N_10122,N_9763,N_9791);
or U10123 (N_10123,N_9736,N_9865);
nor U10124 (N_10124,N_9674,N_9948);
nor U10125 (N_10125,N_9822,N_9907);
xnor U10126 (N_10126,N_9925,N_9863);
or U10127 (N_10127,N_9922,N_9734);
xor U10128 (N_10128,N_9804,N_9889);
nand U10129 (N_10129,N_9663,N_9651);
nand U10130 (N_10130,N_9810,N_9656);
nor U10131 (N_10131,N_9606,N_9842);
and U10132 (N_10132,N_9623,N_9675);
nor U10133 (N_10133,N_9935,N_9908);
nand U10134 (N_10134,N_9873,N_9727);
nor U10135 (N_10135,N_9853,N_9756);
nor U10136 (N_10136,N_9895,N_9959);
nor U10137 (N_10137,N_9916,N_9924);
nand U10138 (N_10138,N_9975,N_9944);
nor U10139 (N_10139,N_9806,N_9955);
or U10140 (N_10140,N_9759,N_9600);
nand U10141 (N_10141,N_9858,N_9648);
nand U10142 (N_10142,N_9799,N_9933);
nor U10143 (N_10143,N_9920,N_9852);
and U10144 (N_10144,N_9884,N_9932);
nand U10145 (N_10145,N_9742,N_9824);
nor U10146 (N_10146,N_9700,N_9701);
nor U10147 (N_10147,N_9951,N_9731);
and U10148 (N_10148,N_9698,N_9917);
and U10149 (N_10149,N_9641,N_9805);
nor U10150 (N_10150,N_9773,N_9891);
or U10151 (N_10151,N_9735,N_9803);
nand U10152 (N_10152,N_9957,N_9626);
nand U10153 (N_10153,N_9758,N_9800);
nor U10154 (N_10154,N_9979,N_9680);
nand U10155 (N_10155,N_9982,N_9787);
or U10156 (N_10156,N_9847,N_9914);
or U10157 (N_10157,N_9638,N_9612);
nand U10158 (N_10158,N_9762,N_9655);
nand U10159 (N_10159,N_9689,N_9849);
or U10160 (N_10160,N_9693,N_9730);
nand U10161 (N_10161,N_9929,N_9831);
nor U10162 (N_10162,N_9918,N_9636);
or U10163 (N_10163,N_9761,N_9926);
nand U10164 (N_10164,N_9795,N_9974);
nand U10165 (N_10165,N_9721,N_9866);
or U10166 (N_10166,N_9963,N_9678);
nor U10167 (N_10167,N_9801,N_9752);
or U10168 (N_10168,N_9850,N_9815);
or U10169 (N_10169,N_9772,N_9953);
nor U10170 (N_10170,N_9738,N_9781);
nand U10171 (N_10171,N_9855,N_9691);
or U10172 (N_10172,N_9796,N_9688);
or U10173 (N_10173,N_9886,N_9906);
or U10174 (N_10174,N_9609,N_9610);
or U10175 (N_10175,N_9882,N_9846);
nand U10176 (N_10176,N_9770,N_9910);
nand U10177 (N_10177,N_9665,N_9793);
or U10178 (N_10178,N_9712,N_9967);
nor U10179 (N_10179,N_9992,N_9627);
or U10180 (N_10180,N_9937,N_9702);
and U10181 (N_10181,N_9856,N_9970);
nor U10182 (N_10182,N_9677,N_9827);
nand U10183 (N_10183,N_9832,N_9880);
or U10184 (N_10184,N_9718,N_9660);
nor U10185 (N_10185,N_9631,N_9697);
nand U10186 (N_10186,N_9613,N_9840);
nor U10187 (N_10187,N_9976,N_9673);
nor U10188 (N_10188,N_9877,N_9633);
and U10189 (N_10189,N_9862,N_9767);
or U10190 (N_10190,N_9820,N_9632);
nor U10191 (N_10191,N_9750,N_9618);
nor U10192 (N_10192,N_9740,N_9921);
nor U10193 (N_10193,N_9905,N_9888);
nor U10194 (N_10194,N_9838,N_9766);
nand U10195 (N_10195,N_9897,N_9919);
nor U10196 (N_10196,N_9848,N_9981);
and U10197 (N_10197,N_9821,N_9964);
or U10198 (N_10198,N_9936,N_9657);
nor U10199 (N_10199,N_9646,N_9694);
nand U10200 (N_10200,N_9876,N_9657);
nand U10201 (N_10201,N_9967,N_9851);
or U10202 (N_10202,N_9727,N_9996);
nand U10203 (N_10203,N_9741,N_9914);
and U10204 (N_10204,N_9791,N_9866);
and U10205 (N_10205,N_9891,N_9663);
nand U10206 (N_10206,N_9717,N_9604);
nand U10207 (N_10207,N_9773,N_9721);
nor U10208 (N_10208,N_9897,N_9914);
nor U10209 (N_10209,N_9933,N_9898);
and U10210 (N_10210,N_9727,N_9675);
nor U10211 (N_10211,N_9807,N_9614);
and U10212 (N_10212,N_9947,N_9729);
nand U10213 (N_10213,N_9677,N_9729);
nand U10214 (N_10214,N_9668,N_9949);
nand U10215 (N_10215,N_9650,N_9707);
nor U10216 (N_10216,N_9912,N_9967);
nand U10217 (N_10217,N_9949,N_9850);
nand U10218 (N_10218,N_9935,N_9642);
or U10219 (N_10219,N_9629,N_9897);
and U10220 (N_10220,N_9889,N_9771);
nand U10221 (N_10221,N_9982,N_9627);
and U10222 (N_10222,N_9954,N_9874);
nor U10223 (N_10223,N_9651,N_9791);
nor U10224 (N_10224,N_9684,N_9982);
or U10225 (N_10225,N_9731,N_9619);
nand U10226 (N_10226,N_9668,N_9944);
or U10227 (N_10227,N_9645,N_9985);
nand U10228 (N_10228,N_9853,N_9719);
nand U10229 (N_10229,N_9830,N_9969);
and U10230 (N_10230,N_9706,N_9723);
nor U10231 (N_10231,N_9690,N_9646);
nand U10232 (N_10232,N_9881,N_9785);
nand U10233 (N_10233,N_9858,N_9708);
nand U10234 (N_10234,N_9971,N_9874);
or U10235 (N_10235,N_9771,N_9696);
and U10236 (N_10236,N_9696,N_9639);
nor U10237 (N_10237,N_9836,N_9751);
and U10238 (N_10238,N_9672,N_9737);
and U10239 (N_10239,N_9972,N_9773);
nor U10240 (N_10240,N_9909,N_9960);
and U10241 (N_10241,N_9858,N_9707);
or U10242 (N_10242,N_9634,N_9905);
and U10243 (N_10243,N_9777,N_9635);
nand U10244 (N_10244,N_9643,N_9991);
nor U10245 (N_10245,N_9806,N_9819);
nor U10246 (N_10246,N_9958,N_9766);
nand U10247 (N_10247,N_9728,N_9759);
or U10248 (N_10248,N_9811,N_9952);
or U10249 (N_10249,N_9888,N_9894);
nor U10250 (N_10250,N_9902,N_9959);
nand U10251 (N_10251,N_9913,N_9635);
nor U10252 (N_10252,N_9801,N_9846);
or U10253 (N_10253,N_9776,N_9711);
or U10254 (N_10254,N_9658,N_9961);
and U10255 (N_10255,N_9686,N_9835);
or U10256 (N_10256,N_9893,N_9948);
and U10257 (N_10257,N_9778,N_9650);
nor U10258 (N_10258,N_9992,N_9781);
nor U10259 (N_10259,N_9653,N_9855);
nor U10260 (N_10260,N_9878,N_9839);
and U10261 (N_10261,N_9654,N_9606);
or U10262 (N_10262,N_9716,N_9722);
nand U10263 (N_10263,N_9914,N_9687);
and U10264 (N_10264,N_9677,N_9755);
and U10265 (N_10265,N_9682,N_9876);
nor U10266 (N_10266,N_9950,N_9749);
and U10267 (N_10267,N_9920,N_9977);
and U10268 (N_10268,N_9859,N_9972);
nand U10269 (N_10269,N_9845,N_9907);
or U10270 (N_10270,N_9913,N_9971);
nor U10271 (N_10271,N_9869,N_9773);
or U10272 (N_10272,N_9680,N_9998);
and U10273 (N_10273,N_9766,N_9933);
nor U10274 (N_10274,N_9632,N_9678);
nor U10275 (N_10275,N_9899,N_9890);
nand U10276 (N_10276,N_9841,N_9767);
or U10277 (N_10277,N_9756,N_9901);
and U10278 (N_10278,N_9732,N_9616);
nor U10279 (N_10279,N_9765,N_9708);
or U10280 (N_10280,N_9685,N_9999);
nand U10281 (N_10281,N_9767,N_9875);
or U10282 (N_10282,N_9731,N_9659);
nor U10283 (N_10283,N_9624,N_9874);
nand U10284 (N_10284,N_9829,N_9650);
or U10285 (N_10285,N_9755,N_9870);
nand U10286 (N_10286,N_9657,N_9933);
nor U10287 (N_10287,N_9658,N_9788);
nand U10288 (N_10288,N_9724,N_9668);
and U10289 (N_10289,N_9793,N_9965);
and U10290 (N_10290,N_9827,N_9950);
and U10291 (N_10291,N_9642,N_9946);
nand U10292 (N_10292,N_9701,N_9862);
nor U10293 (N_10293,N_9665,N_9695);
nand U10294 (N_10294,N_9862,N_9997);
or U10295 (N_10295,N_9807,N_9620);
nand U10296 (N_10296,N_9926,N_9830);
and U10297 (N_10297,N_9875,N_9782);
or U10298 (N_10298,N_9819,N_9638);
nor U10299 (N_10299,N_9689,N_9631);
and U10300 (N_10300,N_9804,N_9872);
or U10301 (N_10301,N_9613,N_9758);
nor U10302 (N_10302,N_9914,N_9600);
and U10303 (N_10303,N_9619,N_9871);
nand U10304 (N_10304,N_9632,N_9951);
nor U10305 (N_10305,N_9988,N_9774);
and U10306 (N_10306,N_9689,N_9894);
or U10307 (N_10307,N_9618,N_9702);
nor U10308 (N_10308,N_9604,N_9864);
nand U10309 (N_10309,N_9744,N_9901);
nor U10310 (N_10310,N_9718,N_9832);
nor U10311 (N_10311,N_9612,N_9708);
nor U10312 (N_10312,N_9940,N_9768);
and U10313 (N_10313,N_9962,N_9956);
nand U10314 (N_10314,N_9784,N_9961);
nor U10315 (N_10315,N_9672,N_9988);
nand U10316 (N_10316,N_9808,N_9663);
or U10317 (N_10317,N_9646,N_9634);
nor U10318 (N_10318,N_9685,N_9851);
and U10319 (N_10319,N_9853,N_9628);
or U10320 (N_10320,N_9690,N_9942);
or U10321 (N_10321,N_9728,N_9779);
and U10322 (N_10322,N_9933,N_9891);
nor U10323 (N_10323,N_9837,N_9742);
or U10324 (N_10324,N_9904,N_9994);
or U10325 (N_10325,N_9915,N_9870);
or U10326 (N_10326,N_9816,N_9805);
nand U10327 (N_10327,N_9832,N_9630);
and U10328 (N_10328,N_9861,N_9753);
nor U10329 (N_10329,N_9919,N_9898);
nor U10330 (N_10330,N_9967,N_9987);
and U10331 (N_10331,N_9816,N_9621);
or U10332 (N_10332,N_9691,N_9735);
or U10333 (N_10333,N_9954,N_9642);
nand U10334 (N_10334,N_9906,N_9654);
nand U10335 (N_10335,N_9656,N_9669);
nor U10336 (N_10336,N_9793,N_9963);
nor U10337 (N_10337,N_9940,N_9689);
and U10338 (N_10338,N_9611,N_9985);
and U10339 (N_10339,N_9621,N_9664);
nor U10340 (N_10340,N_9826,N_9929);
and U10341 (N_10341,N_9936,N_9931);
or U10342 (N_10342,N_9822,N_9751);
and U10343 (N_10343,N_9866,N_9994);
nand U10344 (N_10344,N_9781,N_9884);
nor U10345 (N_10345,N_9881,N_9601);
and U10346 (N_10346,N_9719,N_9644);
nand U10347 (N_10347,N_9836,N_9999);
nand U10348 (N_10348,N_9889,N_9984);
and U10349 (N_10349,N_9672,N_9664);
nor U10350 (N_10350,N_9690,N_9923);
or U10351 (N_10351,N_9917,N_9984);
or U10352 (N_10352,N_9739,N_9787);
nor U10353 (N_10353,N_9731,N_9738);
nand U10354 (N_10354,N_9602,N_9854);
or U10355 (N_10355,N_9726,N_9779);
nand U10356 (N_10356,N_9792,N_9881);
nand U10357 (N_10357,N_9822,N_9672);
nor U10358 (N_10358,N_9961,N_9947);
or U10359 (N_10359,N_9908,N_9817);
nor U10360 (N_10360,N_9750,N_9763);
or U10361 (N_10361,N_9716,N_9946);
and U10362 (N_10362,N_9778,N_9654);
and U10363 (N_10363,N_9844,N_9692);
and U10364 (N_10364,N_9791,N_9863);
nor U10365 (N_10365,N_9776,N_9691);
or U10366 (N_10366,N_9736,N_9879);
nor U10367 (N_10367,N_9659,N_9767);
nor U10368 (N_10368,N_9800,N_9609);
nand U10369 (N_10369,N_9906,N_9863);
nor U10370 (N_10370,N_9815,N_9729);
nor U10371 (N_10371,N_9920,N_9742);
or U10372 (N_10372,N_9985,N_9751);
nor U10373 (N_10373,N_9636,N_9816);
nor U10374 (N_10374,N_9953,N_9716);
nor U10375 (N_10375,N_9694,N_9861);
nand U10376 (N_10376,N_9680,N_9619);
and U10377 (N_10377,N_9788,N_9776);
or U10378 (N_10378,N_9760,N_9608);
or U10379 (N_10379,N_9849,N_9817);
nand U10380 (N_10380,N_9756,N_9790);
or U10381 (N_10381,N_9911,N_9803);
and U10382 (N_10382,N_9679,N_9641);
or U10383 (N_10383,N_9686,N_9614);
or U10384 (N_10384,N_9728,N_9952);
and U10385 (N_10385,N_9754,N_9934);
nor U10386 (N_10386,N_9910,N_9661);
and U10387 (N_10387,N_9714,N_9970);
or U10388 (N_10388,N_9623,N_9938);
nor U10389 (N_10389,N_9770,N_9890);
nand U10390 (N_10390,N_9927,N_9750);
or U10391 (N_10391,N_9759,N_9989);
or U10392 (N_10392,N_9887,N_9711);
and U10393 (N_10393,N_9978,N_9844);
nor U10394 (N_10394,N_9638,N_9962);
nand U10395 (N_10395,N_9621,N_9622);
and U10396 (N_10396,N_9859,N_9877);
nor U10397 (N_10397,N_9812,N_9660);
nand U10398 (N_10398,N_9775,N_9875);
nor U10399 (N_10399,N_9971,N_9837);
and U10400 (N_10400,N_10336,N_10309);
nand U10401 (N_10401,N_10060,N_10086);
nor U10402 (N_10402,N_10390,N_10220);
nor U10403 (N_10403,N_10372,N_10117);
and U10404 (N_10404,N_10205,N_10001);
or U10405 (N_10405,N_10111,N_10080);
nor U10406 (N_10406,N_10025,N_10053);
or U10407 (N_10407,N_10352,N_10260);
and U10408 (N_10408,N_10023,N_10049);
nor U10409 (N_10409,N_10156,N_10145);
nand U10410 (N_10410,N_10254,N_10138);
nor U10411 (N_10411,N_10213,N_10276);
nor U10412 (N_10412,N_10379,N_10386);
nor U10413 (N_10413,N_10020,N_10356);
or U10414 (N_10414,N_10241,N_10291);
nand U10415 (N_10415,N_10341,N_10246);
nor U10416 (N_10416,N_10087,N_10264);
and U10417 (N_10417,N_10282,N_10362);
and U10418 (N_10418,N_10107,N_10056);
nand U10419 (N_10419,N_10158,N_10378);
or U10420 (N_10420,N_10209,N_10244);
xor U10421 (N_10421,N_10189,N_10028);
xor U10422 (N_10422,N_10012,N_10344);
nand U10423 (N_10423,N_10286,N_10251);
nand U10424 (N_10424,N_10228,N_10345);
or U10425 (N_10425,N_10069,N_10383);
nor U10426 (N_10426,N_10338,N_10215);
and U10427 (N_10427,N_10162,N_10150);
or U10428 (N_10428,N_10201,N_10234);
nand U10429 (N_10429,N_10112,N_10275);
nand U10430 (N_10430,N_10248,N_10253);
nand U10431 (N_10431,N_10230,N_10108);
nand U10432 (N_10432,N_10240,N_10174);
and U10433 (N_10433,N_10302,N_10231);
nor U10434 (N_10434,N_10222,N_10333);
nor U10435 (N_10435,N_10081,N_10224);
and U10436 (N_10436,N_10292,N_10301);
or U10437 (N_10437,N_10211,N_10051);
nor U10438 (N_10438,N_10153,N_10398);
nor U10439 (N_10439,N_10126,N_10316);
nor U10440 (N_10440,N_10365,N_10116);
and U10441 (N_10441,N_10115,N_10035);
and U10442 (N_10442,N_10274,N_10340);
and U10443 (N_10443,N_10270,N_10018);
or U10444 (N_10444,N_10159,N_10212);
and U10445 (N_10445,N_10332,N_10010);
and U10446 (N_10446,N_10393,N_10245);
nand U10447 (N_10447,N_10307,N_10299);
xor U10448 (N_10448,N_10261,N_10180);
or U10449 (N_10449,N_10290,N_10247);
and U10450 (N_10450,N_10311,N_10088);
nand U10451 (N_10451,N_10142,N_10078);
nand U10452 (N_10452,N_10041,N_10042);
and U10453 (N_10453,N_10155,N_10385);
nand U10454 (N_10454,N_10024,N_10195);
or U10455 (N_10455,N_10318,N_10040);
nor U10456 (N_10456,N_10085,N_10170);
or U10457 (N_10457,N_10062,N_10368);
nand U10458 (N_10458,N_10308,N_10337);
nand U10459 (N_10459,N_10288,N_10119);
and U10460 (N_10460,N_10033,N_10273);
nand U10461 (N_10461,N_10163,N_10037);
and U10462 (N_10462,N_10278,N_10054);
and U10463 (N_10463,N_10330,N_10339);
or U10464 (N_10464,N_10166,N_10026);
nor U10465 (N_10465,N_10237,N_10191);
nor U10466 (N_10466,N_10347,N_10187);
or U10467 (N_10467,N_10359,N_10343);
nor U10468 (N_10468,N_10384,N_10052);
nand U10469 (N_10469,N_10169,N_10165);
or U10470 (N_10470,N_10090,N_10095);
nor U10471 (N_10471,N_10321,N_10197);
nand U10472 (N_10472,N_10249,N_10227);
and U10473 (N_10473,N_10216,N_10271);
nand U10474 (N_10474,N_10185,N_10003);
and U10475 (N_10475,N_10016,N_10118);
or U10476 (N_10476,N_10008,N_10262);
or U10477 (N_10477,N_10196,N_10179);
nor U10478 (N_10478,N_10329,N_10004);
nand U10479 (N_10479,N_10233,N_10141);
nor U10480 (N_10480,N_10289,N_10312);
nor U10481 (N_10481,N_10357,N_10171);
and U10482 (N_10482,N_10218,N_10198);
and U10483 (N_10483,N_10125,N_10203);
nand U10484 (N_10484,N_10055,N_10015);
or U10485 (N_10485,N_10031,N_10143);
and U10486 (N_10486,N_10148,N_10265);
nor U10487 (N_10487,N_10272,N_10206);
or U10488 (N_10488,N_10223,N_10050);
or U10489 (N_10489,N_10334,N_10214);
and U10490 (N_10490,N_10190,N_10252);
and U10491 (N_10491,N_10006,N_10225);
nand U10492 (N_10492,N_10181,N_10394);
nand U10493 (N_10493,N_10124,N_10146);
nand U10494 (N_10494,N_10120,N_10135);
or U10495 (N_10495,N_10101,N_10217);
nor U10496 (N_10496,N_10131,N_10239);
nor U10497 (N_10497,N_10065,N_10317);
nor U10498 (N_10498,N_10114,N_10202);
nor U10499 (N_10499,N_10236,N_10154);
nor U10500 (N_10500,N_10096,N_10326);
nor U10501 (N_10501,N_10331,N_10349);
or U10502 (N_10502,N_10300,N_10375);
nor U10503 (N_10503,N_10192,N_10039);
nand U10504 (N_10504,N_10259,N_10380);
nor U10505 (N_10505,N_10057,N_10168);
nand U10506 (N_10506,N_10335,N_10034);
nand U10507 (N_10507,N_10173,N_10296);
and U10508 (N_10508,N_10036,N_10200);
nand U10509 (N_10509,N_10066,N_10005);
nor U10510 (N_10510,N_10281,N_10367);
nor U10511 (N_10511,N_10027,N_10161);
or U10512 (N_10512,N_10167,N_10235);
nor U10513 (N_10513,N_10268,N_10194);
nand U10514 (N_10514,N_10269,N_10139);
and U10515 (N_10515,N_10106,N_10075);
nor U10516 (N_10516,N_10103,N_10044);
nand U10517 (N_10517,N_10284,N_10280);
and U10518 (N_10518,N_10364,N_10129);
nor U10519 (N_10519,N_10019,N_10152);
nor U10520 (N_10520,N_10000,N_10243);
nor U10521 (N_10521,N_10105,N_10250);
nor U10522 (N_10522,N_10188,N_10097);
or U10523 (N_10523,N_10058,N_10029);
nor U10524 (N_10524,N_10032,N_10193);
xnor U10525 (N_10525,N_10184,N_10315);
and U10526 (N_10526,N_10009,N_10151);
and U10527 (N_10527,N_10313,N_10391);
and U10528 (N_10528,N_10371,N_10207);
or U10529 (N_10529,N_10350,N_10346);
or U10530 (N_10530,N_10387,N_10396);
or U10531 (N_10531,N_10017,N_10038);
or U10532 (N_10532,N_10083,N_10160);
and U10533 (N_10533,N_10370,N_10325);
xnor U10534 (N_10534,N_10132,N_10133);
and U10535 (N_10535,N_10182,N_10073);
and U10536 (N_10536,N_10011,N_10342);
nor U10537 (N_10537,N_10082,N_10395);
or U10538 (N_10538,N_10305,N_10063);
nand U10539 (N_10539,N_10149,N_10045);
and U10540 (N_10540,N_10186,N_10100);
nor U10541 (N_10541,N_10226,N_10279);
or U10542 (N_10542,N_10283,N_10221);
nand U10543 (N_10543,N_10388,N_10068);
or U10544 (N_10544,N_10084,N_10210);
nor U10545 (N_10545,N_10079,N_10091);
or U10546 (N_10546,N_10102,N_10092);
and U10547 (N_10547,N_10071,N_10059);
or U10548 (N_10548,N_10122,N_10285);
or U10549 (N_10549,N_10157,N_10295);
or U10550 (N_10550,N_10013,N_10258);
nor U10551 (N_10551,N_10098,N_10319);
nor U10552 (N_10552,N_10067,N_10121);
nor U10553 (N_10553,N_10070,N_10110);
nand U10554 (N_10554,N_10074,N_10002);
and U10555 (N_10555,N_10293,N_10361);
and U10556 (N_10556,N_10164,N_10094);
nor U10557 (N_10557,N_10113,N_10183);
and U10558 (N_10558,N_10376,N_10229);
nor U10559 (N_10559,N_10320,N_10354);
nor U10560 (N_10560,N_10363,N_10366);
nand U10561 (N_10561,N_10392,N_10199);
nor U10562 (N_10562,N_10021,N_10324);
nand U10563 (N_10563,N_10369,N_10351);
nand U10564 (N_10564,N_10381,N_10397);
nand U10565 (N_10565,N_10373,N_10263);
nand U10566 (N_10566,N_10130,N_10328);
nor U10567 (N_10567,N_10064,N_10014);
nand U10568 (N_10568,N_10007,N_10172);
nand U10569 (N_10569,N_10238,N_10104);
or U10570 (N_10570,N_10348,N_10177);
nand U10571 (N_10571,N_10399,N_10310);
nor U10572 (N_10572,N_10136,N_10140);
nor U10573 (N_10573,N_10046,N_10304);
and U10574 (N_10574,N_10144,N_10266);
nor U10575 (N_10575,N_10353,N_10048);
and U10576 (N_10576,N_10178,N_10093);
or U10577 (N_10577,N_10355,N_10256);
and U10578 (N_10578,N_10072,N_10323);
and U10579 (N_10579,N_10358,N_10123);
and U10580 (N_10580,N_10389,N_10327);
and U10581 (N_10581,N_10298,N_10137);
nand U10582 (N_10582,N_10099,N_10208);
nor U10583 (N_10583,N_10109,N_10176);
or U10584 (N_10584,N_10077,N_10297);
and U10585 (N_10585,N_10204,N_10374);
nand U10586 (N_10586,N_10242,N_10232);
nand U10587 (N_10587,N_10267,N_10294);
nor U10588 (N_10588,N_10022,N_10047);
nor U10589 (N_10589,N_10030,N_10382);
or U10590 (N_10590,N_10175,N_10089);
or U10591 (N_10591,N_10043,N_10287);
nor U10592 (N_10592,N_10303,N_10255);
and U10593 (N_10593,N_10377,N_10219);
and U10594 (N_10594,N_10314,N_10306);
or U10595 (N_10595,N_10322,N_10147);
and U10596 (N_10596,N_10257,N_10061);
nor U10597 (N_10597,N_10127,N_10277);
nand U10598 (N_10598,N_10128,N_10134);
nand U10599 (N_10599,N_10076,N_10360);
or U10600 (N_10600,N_10212,N_10070);
or U10601 (N_10601,N_10385,N_10054);
or U10602 (N_10602,N_10075,N_10170);
nand U10603 (N_10603,N_10283,N_10248);
nand U10604 (N_10604,N_10190,N_10315);
and U10605 (N_10605,N_10260,N_10259);
nor U10606 (N_10606,N_10226,N_10388);
nand U10607 (N_10607,N_10138,N_10372);
nor U10608 (N_10608,N_10230,N_10189);
and U10609 (N_10609,N_10304,N_10254);
nor U10610 (N_10610,N_10359,N_10260);
nor U10611 (N_10611,N_10323,N_10024);
or U10612 (N_10612,N_10316,N_10092);
and U10613 (N_10613,N_10375,N_10234);
or U10614 (N_10614,N_10387,N_10233);
and U10615 (N_10615,N_10229,N_10394);
nand U10616 (N_10616,N_10352,N_10100);
or U10617 (N_10617,N_10125,N_10181);
and U10618 (N_10618,N_10341,N_10396);
nor U10619 (N_10619,N_10333,N_10000);
and U10620 (N_10620,N_10210,N_10079);
nor U10621 (N_10621,N_10138,N_10299);
or U10622 (N_10622,N_10010,N_10311);
nor U10623 (N_10623,N_10026,N_10058);
nor U10624 (N_10624,N_10161,N_10121);
and U10625 (N_10625,N_10098,N_10208);
nor U10626 (N_10626,N_10206,N_10229);
or U10627 (N_10627,N_10368,N_10111);
and U10628 (N_10628,N_10141,N_10241);
and U10629 (N_10629,N_10141,N_10394);
and U10630 (N_10630,N_10039,N_10243);
and U10631 (N_10631,N_10043,N_10120);
nor U10632 (N_10632,N_10324,N_10284);
nand U10633 (N_10633,N_10255,N_10225);
nand U10634 (N_10634,N_10282,N_10306);
and U10635 (N_10635,N_10353,N_10123);
nor U10636 (N_10636,N_10188,N_10320);
nor U10637 (N_10637,N_10109,N_10220);
nor U10638 (N_10638,N_10065,N_10123);
nor U10639 (N_10639,N_10142,N_10081);
nand U10640 (N_10640,N_10118,N_10063);
nand U10641 (N_10641,N_10255,N_10133);
nor U10642 (N_10642,N_10072,N_10107);
or U10643 (N_10643,N_10369,N_10004);
or U10644 (N_10644,N_10162,N_10234);
nand U10645 (N_10645,N_10385,N_10250);
and U10646 (N_10646,N_10360,N_10335);
nand U10647 (N_10647,N_10031,N_10032);
nor U10648 (N_10648,N_10382,N_10027);
and U10649 (N_10649,N_10187,N_10314);
and U10650 (N_10650,N_10369,N_10266);
nor U10651 (N_10651,N_10064,N_10046);
nor U10652 (N_10652,N_10025,N_10139);
and U10653 (N_10653,N_10177,N_10246);
or U10654 (N_10654,N_10379,N_10307);
nor U10655 (N_10655,N_10302,N_10002);
and U10656 (N_10656,N_10344,N_10339);
nand U10657 (N_10657,N_10149,N_10125);
and U10658 (N_10658,N_10014,N_10042);
and U10659 (N_10659,N_10109,N_10282);
or U10660 (N_10660,N_10134,N_10227);
and U10661 (N_10661,N_10266,N_10119);
nand U10662 (N_10662,N_10034,N_10063);
nand U10663 (N_10663,N_10099,N_10293);
or U10664 (N_10664,N_10156,N_10002);
nor U10665 (N_10665,N_10141,N_10161);
or U10666 (N_10666,N_10134,N_10120);
nor U10667 (N_10667,N_10246,N_10247);
nor U10668 (N_10668,N_10273,N_10262);
or U10669 (N_10669,N_10042,N_10377);
or U10670 (N_10670,N_10171,N_10212);
nand U10671 (N_10671,N_10032,N_10138);
nor U10672 (N_10672,N_10342,N_10068);
or U10673 (N_10673,N_10174,N_10200);
and U10674 (N_10674,N_10391,N_10140);
nand U10675 (N_10675,N_10338,N_10161);
and U10676 (N_10676,N_10126,N_10066);
nand U10677 (N_10677,N_10333,N_10367);
nor U10678 (N_10678,N_10292,N_10053);
nand U10679 (N_10679,N_10223,N_10390);
or U10680 (N_10680,N_10076,N_10157);
nor U10681 (N_10681,N_10154,N_10345);
nor U10682 (N_10682,N_10376,N_10173);
or U10683 (N_10683,N_10022,N_10186);
or U10684 (N_10684,N_10262,N_10333);
nand U10685 (N_10685,N_10019,N_10099);
nand U10686 (N_10686,N_10242,N_10099);
and U10687 (N_10687,N_10350,N_10302);
nand U10688 (N_10688,N_10067,N_10101);
nor U10689 (N_10689,N_10084,N_10151);
and U10690 (N_10690,N_10388,N_10096);
and U10691 (N_10691,N_10325,N_10213);
or U10692 (N_10692,N_10254,N_10153);
or U10693 (N_10693,N_10220,N_10383);
nor U10694 (N_10694,N_10392,N_10202);
or U10695 (N_10695,N_10201,N_10296);
or U10696 (N_10696,N_10259,N_10245);
nand U10697 (N_10697,N_10372,N_10016);
nor U10698 (N_10698,N_10370,N_10364);
or U10699 (N_10699,N_10188,N_10008);
or U10700 (N_10700,N_10150,N_10052);
nor U10701 (N_10701,N_10261,N_10196);
nor U10702 (N_10702,N_10347,N_10124);
and U10703 (N_10703,N_10275,N_10198);
and U10704 (N_10704,N_10367,N_10186);
nor U10705 (N_10705,N_10269,N_10147);
or U10706 (N_10706,N_10365,N_10183);
nand U10707 (N_10707,N_10187,N_10258);
or U10708 (N_10708,N_10036,N_10163);
and U10709 (N_10709,N_10385,N_10345);
nor U10710 (N_10710,N_10324,N_10062);
and U10711 (N_10711,N_10362,N_10349);
nor U10712 (N_10712,N_10299,N_10376);
nand U10713 (N_10713,N_10267,N_10182);
nor U10714 (N_10714,N_10243,N_10099);
nand U10715 (N_10715,N_10187,N_10230);
and U10716 (N_10716,N_10303,N_10328);
or U10717 (N_10717,N_10139,N_10003);
and U10718 (N_10718,N_10144,N_10259);
nor U10719 (N_10719,N_10155,N_10004);
or U10720 (N_10720,N_10135,N_10026);
and U10721 (N_10721,N_10102,N_10236);
or U10722 (N_10722,N_10305,N_10317);
nor U10723 (N_10723,N_10171,N_10069);
nor U10724 (N_10724,N_10026,N_10124);
or U10725 (N_10725,N_10048,N_10099);
nand U10726 (N_10726,N_10384,N_10289);
and U10727 (N_10727,N_10003,N_10078);
nand U10728 (N_10728,N_10318,N_10029);
nor U10729 (N_10729,N_10274,N_10334);
or U10730 (N_10730,N_10335,N_10200);
nand U10731 (N_10731,N_10372,N_10201);
or U10732 (N_10732,N_10069,N_10300);
nor U10733 (N_10733,N_10075,N_10058);
nand U10734 (N_10734,N_10318,N_10007);
nand U10735 (N_10735,N_10319,N_10161);
and U10736 (N_10736,N_10305,N_10087);
and U10737 (N_10737,N_10342,N_10105);
nand U10738 (N_10738,N_10317,N_10184);
nand U10739 (N_10739,N_10257,N_10197);
or U10740 (N_10740,N_10208,N_10371);
and U10741 (N_10741,N_10038,N_10149);
and U10742 (N_10742,N_10088,N_10243);
nor U10743 (N_10743,N_10276,N_10322);
and U10744 (N_10744,N_10298,N_10358);
nor U10745 (N_10745,N_10016,N_10164);
nor U10746 (N_10746,N_10103,N_10071);
and U10747 (N_10747,N_10346,N_10193);
nor U10748 (N_10748,N_10273,N_10388);
and U10749 (N_10749,N_10311,N_10314);
or U10750 (N_10750,N_10294,N_10078);
nand U10751 (N_10751,N_10149,N_10048);
or U10752 (N_10752,N_10122,N_10182);
and U10753 (N_10753,N_10392,N_10382);
and U10754 (N_10754,N_10077,N_10054);
nand U10755 (N_10755,N_10078,N_10358);
nand U10756 (N_10756,N_10075,N_10266);
and U10757 (N_10757,N_10126,N_10381);
nand U10758 (N_10758,N_10329,N_10330);
nor U10759 (N_10759,N_10040,N_10185);
nand U10760 (N_10760,N_10071,N_10108);
or U10761 (N_10761,N_10360,N_10213);
or U10762 (N_10762,N_10108,N_10103);
or U10763 (N_10763,N_10320,N_10146);
or U10764 (N_10764,N_10290,N_10099);
or U10765 (N_10765,N_10010,N_10002);
nor U10766 (N_10766,N_10149,N_10243);
and U10767 (N_10767,N_10177,N_10065);
or U10768 (N_10768,N_10179,N_10272);
and U10769 (N_10769,N_10109,N_10329);
nand U10770 (N_10770,N_10304,N_10028);
or U10771 (N_10771,N_10273,N_10139);
nand U10772 (N_10772,N_10054,N_10068);
nor U10773 (N_10773,N_10151,N_10361);
and U10774 (N_10774,N_10225,N_10098);
nor U10775 (N_10775,N_10243,N_10142);
nand U10776 (N_10776,N_10322,N_10028);
nand U10777 (N_10777,N_10323,N_10398);
and U10778 (N_10778,N_10112,N_10079);
nand U10779 (N_10779,N_10373,N_10247);
or U10780 (N_10780,N_10359,N_10079);
nand U10781 (N_10781,N_10053,N_10367);
nor U10782 (N_10782,N_10317,N_10376);
and U10783 (N_10783,N_10073,N_10151);
and U10784 (N_10784,N_10339,N_10056);
or U10785 (N_10785,N_10137,N_10016);
or U10786 (N_10786,N_10147,N_10390);
and U10787 (N_10787,N_10365,N_10386);
nor U10788 (N_10788,N_10232,N_10112);
or U10789 (N_10789,N_10037,N_10273);
nand U10790 (N_10790,N_10204,N_10259);
and U10791 (N_10791,N_10121,N_10192);
nand U10792 (N_10792,N_10184,N_10253);
nand U10793 (N_10793,N_10183,N_10004);
nand U10794 (N_10794,N_10320,N_10298);
nand U10795 (N_10795,N_10384,N_10261);
nor U10796 (N_10796,N_10225,N_10019);
and U10797 (N_10797,N_10228,N_10292);
or U10798 (N_10798,N_10166,N_10146);
nor U10799 (N_10799,N_10286,N_10191);
and U10800 (N_10800,N_10560,N_10701);
or U10801 (N_10801,N_10605,N_10575);
nor U10802 (N_10802,N_10625,N_10699);
nor U10803 (N_10803,N_10726,N_10542);
nor U10804 (N_10804,N_10450,N_10505);
and U10805 (N_10805,N_10449,N_10617);
nor U10806 (N_10806,N_10659,N_10741);
and U10807 (N_10807,N_10703,N_10720);
or U10808 (N_10808,N_10700,N_10459);
and U10809 (N_10809,N_10656,N_10432);
and U10810 (N_10810,N_10643,N_10756);
and U10811 (N_10811,N_10568,N_10710);
and U10812 (N_10812,N_10424,N_10429);
and U10813 (N_10813,N_10418,N_10722);
xnor U10814 (N_10814,N_10408,N_10472);
and U10815 (N_10815,N_10727,N_10520);
nor U10816 (N_10816,N_10503,N_10463);
nand U10817 (N_10817,N_10614,N_10721);
nand U10818 (N_10818,N_10532,N_10436);
or U10819 (N_10819,N_10653,N_10538);
and U10820 (N_10820,N_10517,N_10431);
nand U10821 (N_10821,N_10404,N_10446);
nand U10822 (N_10822,N_10524,N_10594);
or U10823 (N_10823,N_10546,N_10790);
and U10824 (N_10824,N_10685,N_10563);
or U10825 (N_10825,N_10640,N_10655);
or U10826 (N_10826,N_10521,N_10670);
nor U10827 (N_10827,N_10508,N_10416);
nand U10828 (N_10828,N_10519,N_10476);
nor U10829 (N_10829,N_10777,N_10554);
and U10830 (N_10830,N_10526,N_10717);
or U10831 (N_10831,N_10552,N_10651);
or U10832 (N_10832,N_10786,N_10737);
and U10833 (N_10833,N_10799,N_10510);
and U10834 (N_10834,N_10781,N_10636);
or U10835 (N_10835,N_10584,N_10414);
and U10836 (N_10836,N_10448,N_10602);
or U10837 (N_10837,N_10691,N_10473);
or U10838 (N_10838,N_10761,N_10627);
nor U10839 (N_10839,N_10465,N_10797);
or U10840 (N_10840,N_10783,N_10582);
or U10841 (N_10841,N_10724,N_10599);
nand U10842 (N_10842,N_10425,N_10740);
nand U10843 (N_10843,N_10671,N_10588);
nor U10844 (N_10844,N_10528,N_10662);
nor U10845 (N_10845,N_10693,N_10591);
or U10846 (N_10846,N_10491,N_10742);
or U10847 (N_10847,N_10674,N_10587);
and U10848 (N_10848,N_10657,N_10489);
nand U10849 (N_10849,N_10712,N_10497);
nor U10850 (N_10850,N_10539,N_10445);
nor U10851 (N_10851,N_10628,N_10547);
or U10852 (N_10852,N_10695,N_10441);
or U10853 (N_10853,N_10597,N_10401);
or U10854 (N_10854,N_10557,N_10725);
nand U10855 (N_10855,N_10745,N_10707);
nor U10856 (N_10856,N_10577,N_10458);
nand U10857 (N_10857,N_10647,N_10555);
nor U10858 (N_10858,N_10788,N_10637);
or U10859 (N_10859,N_10744,N_10677);
nor U10860 (N_10860,N_10567,N_10456);
nand U10861 (N_10861,N_10439,N_10772);
nor U10862 (N_10862,N_10496,N_10665);
nand U10863 (N_10863,N_10791,N_10775);
nand U10864 (N_10864,N_10768,N_10592);
or U10865 (N_10865,N_10603,N_10421);
nand U10866 (N_10866,N_10733,N_10709);
or U10867 (N_10867,N_10753,N_10534);
nor U10868 (N_10868,N_10752,N_10624);
nand U10869 (N_10869,N_10646,N_10470);
and U10870 (N_10870,N_10481,N_10440);
nand U10871 (N_10871,N_10748,N_10593);
and U10872 (N_10872,N_10638,N_10686);
and U10873 (N_10873,N_10420,N_10410);
nand U10874 (N_10874,N_10518,N_10796);
and U10875 (N_10875,N_10711,N_10457);
nand U10876 (N_10876,N_10688,N_10664);
nand U10877 (N_10877,N_10596,N_10762);
nand U10878 (N_10878,N_10409,N_10434);
nand U10879 (N_10879,N_10447,N_10760);
nor U10880 (N_10880,N_10641,N_10773);
or U10881 (N_10881,N_10732,N_10715);
or U10882 (N_10882,N_10723,N_10407);
nor U10883 (N_10883,N_10702,N_10649);
nor U10884 (N_10884,N_10494,N_10525);
and U10885 (N_10885,N_10586,N_10570);
nor U10886 (N_10886,N_10573,N_10704);
nor U10887 (N_10887,N_10765,N_10739);
or U10888 (N_10888,N_10566,N_10415);
nand U10889 (N_10889,N_10750,N_10442);
or U10890 (N_10890,N_10572,N_10585);
and U10891 (N_10891,N_10530,N_10606);
and U10892 (N_10892,N_10474,N_10716);
or U10893 (N_10893,N_10589,N_10776);
or U10894 (N_10894,N_10697,N_10569);
or U10895 (N_10895,N_10611,N_10734);
and U10896 (N_10896,N_10738,N_10438);
or U10897 (N_10897,N_10444,N_10405);
nand U10898 (N_10898,N_10559,N_10679);
or U10899 (N_10899,N_10486,N_10485);
or U10900 (N_10900,N_10619,N_10435);
or U10901 (N_10901,N_10549,N_10654);
nand U10902 (N_10902,N_10523,N_10574);
and U10903 (N_10903,N_10652,N_10464);
and U10904 (N_10904,N_10479,N_10692);
nor U10905 (N_10905,N_10488,N_10499);
nor U10906 (N_10906,N_10427,N_10437);
or U10907 (N_10907,N_10419,N_10764);
and U10908 (N_10908,N_10504,N_10561);
or U10909 (N_10909,N_10749,N_10675);
or U10910 (N_10910,N_10512,N_10634);
nand U10911 (N_10911,N_10422,N_10668);
nand U10912 (N_10912,N_10607,N_10751);
or U10913 (N_10913,N_10779,N_10430);
nand U10914 (N_10914,N_10527,N_10551);
nand U10915 (N_10915,N_10579,N_10713);
or U10916 (N_10916,N_10537,N_10471);
and U10917 (N_10917,N_10669,N_10622);
and U10918 (N_10918,N_10729,N_10792);
nand U10919 (N_10919,N_10580,N_10564);
nand U10920 (N_10920,N_10730,N_10660);
nand U10921 (N_10921,N_10482,N_10412);
xnor U10922 (N_10922,N_10536,N_10601);
and U10923 (N_10923,N_10644,N_10746);
nor U10924 (N_10924,N_10774,N_10453);
or U10925 (N_10925,N_10452,N_10475);
nand U10926 (N_10926,N_10633,N_10565);
nor U10927 (N_10927,N_10492,N_10500);
nand U10928 (N_10928,N_10658,N_10728);
nor U10929 (N_10929,N_10502,N_10680);
and U10930 (N_10930,N_10506,N_10516);
nor U10931 (N_10931,N_10477,N_10501);
or U10932 (N_10932,N_10763,N_10608);
nor U10933 (N_10933,N_10618,N_10469);
and U10934 (N_10934,N_10583,N_10681);
and U10935 (N_10935,N_10642,N_10787);
and U10936 (N_10936,N_10443,N_10609);
and U10937 (N_10937,N_10639,N_10755);
and U10938 (N_10938,N_10400,N_10632);
nor U10939 (N_10939,N_10694,N_10648);
and U10940 (N_10940,N_10548,N_10667);
nand U10941 (N_10941,N_10795,N_10461);
nor U10942 (N_10942,N_10417,N_10630);
nand U10943 (N_10943,N_10758,N_10770);
nor U10944 (N_10944,N_10507,N_10454);
nor U10945 (N_10945,N_10682,N_10478);
and U10946 (N_10946,N_10426,N_10413);
and U10947 (N_10947,N_10615,N_10498);
nor U10948 (N_10948,N_10631,N_10511);
nand U10949 (N_10949,N_10698,N_10673);
nand U10950 (N_10950,N_10696,N_10541);
and U10951 (N_10951,N_10754,N_10544);
nor U10952 (N_10952,N_10621,N_10714);
and U10953 (N_10953,N_10483,N_10793);
nand U10954 (N_10954,N_10533,N_10610);
or U10955 (N_10955,N_10411,N_10433);
or U10956 (N_10956,N_10490,N_10645);
nand U10957 (N_10957,N_10543,N_10403);
or U10958 (N_10958,N_10626,N_10798);
or U10959 (N_10959,N_10529,N_10576);
nor U10960 (N_10960,N_10757,N_10487);
or U10961 (N_10961,N_10612,N_10629);
nand U10962 (N_10962,N_10689,N_10620);
nor U10963 (N_10963,N_10598,N_10778);
nand U10964 (N_10964,N_10406,N_10635);
and U10965 (N_10965,N_10545,N_10785);
and U10966 (N_10966,N_10731,N_10767);
or U10967 (N_10967,N_10402,N_10661);
nor U10968 (N_10968,N_10706,N_10515);
or U10969 (N_10969,N_10581,N_10613);
and U10970 (N_10970,N_10460,N_10759);
and U10971 (N_10971,N_10535,N_10604);
and U10972 (N_10972,N_10719,N_10540);
or U10973 (N_10973,N_10467,N_10623);
nand U10974 (N_10974,N_10766,N_10743);
or U10975 (N_10975,N_10769,N_10571);
and U10976 (N_10976,N_10553,N_10708);
and U10977 (N_10977,N_10531,N_10690);
and U10978 (N_10978,N_10794,N_10784);
nor U10979 (N_10979,N_10663,N_10678);
nand U10980 (N_10980,N_10484,N_10466);
or U10981 (N_10981,N_10514,N_10578);
or U10982 (N_10982,N_10480,N_10771);
nor U10983 (N_10983,N_10495,N_10513);
nand U10984 (N_10984,N_10687,N_10600);
nand U10985 (N_10985,N_10683,N_10595);
and U10986 (N_10986,N_10705,N_10493);
nor U10987 (N_10987,N_10509,N_10558);
or U10988 (N_10988,N_10616,N_10650);
xor U10989 (N_10989,N_10736,N_10782);
and U10990 (N_10990,N_10562,N_10590);
or U10991 (N_10991,N_10735,N_10718);
nor U10992 (N_10992,N_10789,N_10780);
and U10993 (N_10993,N_10522,N_10676);
or U10994 (N_10994,N_10423,N_10462);
nand U10995 (N_10995,N_10747,N_10550);
nand U10996 (N_10996,N_10556,N_10684);
nor U10997 (N_10997,N_10468,N_10666);
and U10998 (N_10998,N_10451,N_10455);
and U10999 (N_10999,N_10428,N_10672);
nand U11000 (N_11000,N_10792,N_10513);
or U11001 (N_11001,N_10691,N_10463);
and U11002 (N_11002,N_10693,N_10744);
nor U11003 (N_11003,N_10794,N_10544);
nand U11004 (N_11004,N_10436,N_10597);
or U11005 (N_11005,N_10751,N_10418);
or U11006 (N_11006,N_10767,N_10419);
or U11007 (N_11007,N_10477,N_10412);
nor U11008 (N_11008,N_10669,N_10687);
nor U11009 (N_11009,N_10597,N_10509);
or U11010 (N_11010,N_10643,N_10677);
nor U11011 (N_11011,N_10513,N_10425);
nor U11012 (N_11012,N_10536,N_10570);
nor U11013 (N_11013,N_10525,N_10745);
nor U11014 (N_11014,N_10445,N_10718);
nor U11015 (N_11015,N_10689,N_10597);
and U11016 (N_11016,N_10565,N_10674);
or U11017 (N_11017,N_10771,N_10572);
or U11018 (N_11018,N_10783,N_10790);
nor U11019 (N_11019,N_10752,N_10413);
or U11020 (N_11020,N_10603,N_10679);
and U11021 (N_11021,N_10762,N_10788);
nor U11022 (N_11022,N_10675,N_10728);
and U11023 (N_11023,N_10647,N_10764);
and U11024 (N_11024,N_10512,N_10687);
and U11025 (N_11025,N_10487,N_10566);
and U11026 (N_11026,N_10403,N_10710);
and U11027 (N_11027,N_10441,N_10422);
nand U11028 (N_11028,N_10612,N_10560);
nand U11029 (N_11029,N_10756,N_10633);
nor U11030 (N_11030,N_10491,N_10635);
nand U11031 (N_11031,N_10738,N_10471);
and U11032 (N_11032,N_10736,N_10457);
or U11033 (N_11033,N_10661,N_10571);
and U11034 (N_11034,N_10508,N_10794);
nor U11035 (N_11035,N_10580,N_10640);
or U11036 (N_11036,N_10788,N_10594);
nand U11037 (N_11037,N_10564,N_10542);
or U11038 (N_11038,N_10486,N_10456);
or U11039 (N_11039,N_10402,N_10670);
nor U11040 (N_11040,N_10565,N_10455);
nand U11041 (N_11041,N_10629,N_10651);
and U11042 (N_11042,N_10601,N_10512);
nand U11043 (N_11043,N_10784,N_10652);
nor U11044 (N_11044,N_10598,N_10482);
and U11045 (N_11045,N_10439,N_10534);
and U11046 (N_11046,N_10683,N_10597);
or U11047 (N_11047,N_10611,N_10621);
nor U11048 (N_11048,N_10613,N_10526);
nand U11049 (N_11049,N_10604,N_10495);
nor U11050 (N_11050,N_10575,N_10790);
xor U11051 (N_11051,N_10732,N_10499);
nand U11052 (N_11052,N_10617,N_10572);
and U11053 (N_11053,N_10505,N_10409);
nor U11054 (N_11054,N_10647,N_10626);
nand U11055 (N_11055,N_10405,N_10740);
nor U11056 (N_11056,N_10685,N_10687);
nor U11057 (N_11057,N_10554,N_10446);
nor U11058 (N_11058,N_10649,N_10716);
nand U11059 (N_11059,N_10459,N_10737);
nor U11060 (N_11060,N_10486,N_10632);
or U11061 (N_11061,N_10439,N_10481);
nand U11062 (N_11062,N_10404,N_10753);
or U11063 (N_11063,N_10743,N_10780);
nor U11064 (N_11064,N_10412,N_10521);
or U11065 (N_11065,N_10721,N_10485);
or U11066 (N_11066,N_10798,N_10691);
or U11067 (N_11067,N_10592,N_10622);
or U11068 (N_11068,N_10679,N_10784);
and U11069 (N_11069,N_10609,N_10581);
and U11070 (N_11070,N_10773,N_10785);
nand U11071 (N_11071,N_10410,N_10520);
or U11072 (N_11072,N_10694,N_10742);
nand U11073 (N_11073,N_10707,N_10771);
and U11074 (N_11074,N_10780,N_10475);
nand U11075 (N_11075,N_10789,N_10717);
and U11076 (N_11076,N_10766,N_10564);
and U11077 (N_11077,N_10594,N_10719);
and U11078 (N_11078,N_10604,N_10481);
and U11079 (N_11079,N_10495,N_10584);
and U11080 (N_11080,N_10652,N_10580);
or U11081 (N_11081,N_10663,N_10662);
nand U11082 (N_11082,N_10503,N_10548);
nand U11083 (N_11083,N_10561,N_10573);
nand U11084 (N_11084,N_10795,N_10735);
and U11085 (N_11085,N_10649,N_10570);
nor U11086 (N_11086,N_10589,N_10544);
nand U11087 (N_11087,N_10704,N_10543);
and U11088 (N_11088,N_10798,N_10675);
nor U11089 (N_11089,N_10725,N_10681);
or U11090 (N_11090,N_10673,N_10652);
nand U11091 (N_11091,N_10593,N_10709);
nand U11092 (N_11092,N_10596,N_10589);
and U11093 (N_11093,N_10409,N_10678);
nor U11094 (N_11094,N_10615,N_10603);
nand U11095 (N_11095,N_10507,N_10408);
or U11096 (N_11096,N_10727,N_10756);
nand U11097 (N_11097,N_10477,N_10614);
nor U11098 (N_11098,N_10530,N_10509);
nand U11099 (N_11099,N_10763,N_10425);
nor U11100 (N_11100,N_10785,N_10442);
xor U11101 (N_11101,N_10732,N_10656);
nor U11102 (N_11102,N_10551,N_10627);
or U11103 (N_11103,N_10719,N_10406);
nor U11104 (N_11104,N_10634,N_10541);
and U11105 (N_11105,N_10649,N_10492);
nand U11106 (N_11106,N_10521,N_10692);
and U11107 (N_11107,N_10747,N_10585);
and U11108 (N_11108,N_10488,N_10454);
nor U11109 (N_11109,N_10675,N_10460);
nor U11110 (N_11110,N_10646,N_10607);
nor U11111 (N_11111,N_10458,N_10791);
nand U11112 (N_11112,N_10687,N_10583);
nor U11113 (N_11113,N_10713,N_10530);
nand U11114 (N_11114,N_10509,N_10617);
nand U11115 (N_11115,N_10759,N_10646);
nor U11116 (N_11116,N_10527,N_10609);
nor U11117 (N_11117,N_10683,N_10556);
and U11118 (N_11118,N_10478,N_10552);
and U11119 (N_11119,N_10712,N_10693);
or U11120 (N_11120,N_10470,N_10623);
nor U11121 (N_11121,N_10417,N_10401);
or U11122 (N_11122,N_10613,N_10792);
nor U11123 (N_11123,N_10659,N_10405);
and U11124 (N_11124,N_10624,N_10508);
or U11125 (N_11125,N_10721,N_10585);
nor U11126 (N_11126,N_10491,N_10597);
nand U11127 (N_11127,N_10697,N_10455);
or U11128 (N_11128,N_10620,N_10736);
or U11129 (N_11129,N_10531,N_10725);
or U11130 (N_11130,N_10400,N_10438);
or U11131 (N_11131,N_10428,N_10779);
nand U11132 (N_11132,N_10605,N_10783);
and U11133 (N_11133,N_10795,N_10669);
and U11134 (N_11134,N_10792,N_10571);
nand U11135 (N_11135,N_10517,N_10565);
or U11136 (N_11136,N_10716,N_10664);
and U11137 (N_11137,N_10668,N_10552);
nand U11138 (N_11138,N_10498,N_10738);
nand U11139 (N_11139,N_10730,N_10519);
nand U11140 (N_11140,N_10644,N_10769);
and U11141 (N_11141,N_10432,N_10754);
nor U11142 (N_11142,N_10490,N_10571);
nand U11143 (N_11143,N_10483,N_10593);
and U11144 (N_11144,N_10524,N_10629);
nand U11145 (N_11145,N_10791,N_10513);
or U11146 (N_11146,N_10533,N_10460);
nor U11147 (N_11147,N_10714,N_10577);
or U11148 (N_11148,N_10483,N_10648);
or U11149 (N_11149,N_10406,N_10535);
nand U11150 (N_11150,N_10559,N_10521);
and U11151 (N_11151,N_10640,N_10507);
nand U11152 (N_11152,N_10553,N_10630);
nand U11153 (N_11153,N_10665,N_10444);
and U11154 (N_11154,N_10507,N_10757);
nand U11155 (N_11155,N_10750,N_10792);
nand U11156 (N_11156,N_10589,N_10513);
or U11157 (N_11157,N_10568,N_10750);
or U11158 (N_11158,N_10493,N_10522);
or U11159 (N_11159,N_10486,N_10453);
and U11160 (N_11160,N_10523,N_10705);
nor U11161 (N_11161,N_10417,N_10406);
nor U11162 (N_11162,N_10671,N_10778);
or U11163 (N_11163,N_10682,N_10751);
nor U11164 (N_11164,N_10510,N_10407);
and U11165 (N_11165,N_10516,N_10709);
and U11166 (N_11166,N_10662,N_10616);
nor U11167 (N_11167,N_10608,N_10755);
nor U11168 (N_11168,N_10614,N_10788);
and U11169 (N_11169,N_10776,N_10428);
or U11170 (N_11170,N_10704,N_10760);
nor U11171 (N_11171,N_10647,N_10769);
nor U11172 (N_11172,N_10491,N_10415);
and U11173 (N_11173,N_10717,N_10758);
and U11174 (N_11174,N_10747,N_10533);
nor U11175 (N_11175,N_10435,N_10418);
or U11176 (N_11176,N_10729,N_10609);
nor U11177 (N_11177,N_10762,N_10611);
and U11178 (N_11178,N_10580,N_10627);
or U11179 (N_11179,N_10565,N_10671);
or U11180 (N_11180,N_10658,N_10491);
nor U11181 (N_11181,N_10430,N_10530);
nand U11182 (N_11182,N_10465,N_10515);
and U11183 (N_11183,N_10737,N_10777);
nor U11184 (N_11184,N_10658,N_10750);
or U11185 (N_11185,N_10756,N_10597);
or U11186 (N_11186,N_10469,N_10475);
and U11187 (N_11187,N_10747,N_10642);
nor U11188 (N_11188,N_10517,N_10758);
nand U11189 (N_11189,N_10531,N_10765);
nor U11190 (N_11190,N_10438,N_10409);
and U11191 (N_11191,N_10413,N_10525);
or U11192 (N_11192,N_10671,N_10529);
or U11193 (N_11193,N_10529,N_10721);
or U11194 (N_11194,N_10587,N_10485);
and U11195 (N_11195,N_10714,N_10522);
xor U11196 (N_11196,N_10564,N_10779);
nand U11197 (N_11197,N_10635,N_10693);
nor U11198 (N_11198,N_10657,N_10585);
or U11199 (N_11199,N_10535,N_10766);
nand U11200 (N_11200,N_11095,N_11087);
and U11201 (N_11201,N_11141,N_10858);
and U11202 (N_11202,N_10932,N_10879);
nand U11203 (N_11203,N_10815,N_10871);
nor U11204 (N_11204,N_10803,N_10863);
or U11205 (N_11205,N_10820,N_10845);
and U11206 (N_11206,N_11011,N_11037);
and U11207 (N_11207,N_10853,N_10850);
and U11208 (N_11208,N_11038,N_11181);
and U11209 (N_11209,N_11100,N_11086);
nand U11210 (N_11210,N_10951,N_10891);
nor U11211 (N_11211,N_10811,N_10905);
xor U11212 (N_11212,N_11122,N_11066);
nor U11213 (N_11213,N_11159,N_10913);
nor U11214 (N_11214,N_10971,N_11179);
nor U11215 (N_11215,N_11025,N_11083);
nand U11216 (N_11216,N_11151,N_11171);
nor U11217 (N_11217,N_11187,N_11174);
nor U11218 (N_11218,N_11175,N_11137);
nand U11219 (N_11219,N_11144,N_11048);
and U11220 (N_11220,N_10800,N_10958);
and U11221 (N_11221,N_10847,N_10983);
and U11222 (N_11222,N_10824,N_10935);
and U11223 (N_11223,N_10816,N_10894);
nor U11224 (N_11224,N_11135,N_11126);
nor U11225 (N_11225,N_11125,N_10985);
nor U11226 (N_11226,N_10939,N_11019);
or U11227 (N_11227,N_11013,N_10862);
nand U11228 (N_11228,N_11153,N_11184);
nor U11229 (N_11229,N_10989,N_11186);
nor U11230 (N_11230,N_11057,N_10825);
nor U11231 (N_11231,N_11041,N_10952);
nand U11232 (N_11232,N_10868,N_11018);
nor U11233 (N_11233,N_11056,N_11076);
nor U11234 (N_11234,N_10967,N_11118);
nand U11235 (N_11235,N_11177,N_11132);
nor U11236 (N_11236,N_10940,N_11069);
or U11237 (N_11237,N_11136,N_10882);
and U11238 (N_11238,N_11047,N_11110);
or U11239 (N_11239,N_11005,N_10835);
and U11240 (N_11240,N_11101,N_10990);
nor U11241 (N_11241,N_10867,N_11052);
and U11242 (N_11242,N_10901,N_11124);
nand U11243 (N_11243,N_11073,N_11189);
or U11244 (N_11244,N_10978,N_11060);
or U11245 (N_11245,N_10878,N_10836);
and U11246 (N_11246,N_11152,N_10949);
nand U11247 (N_11247,N_10801,N_10916);
nand U11248 (N_11248,N_11198,N_10922);
nor U11249 (N_11249,N_10831,N_10995);
and U11250 (N_11250,N_11072,N_10827);
and U11251 (N_11251,N_10906,N_11096);
or U11252 (N_11252,N_10822,N_11067);
and U11253 (N_11253,N_11007,N_10838);
nand U11254 (N_11254,N_10819,N_10991);
nand U11255 (N_11255,N_11170,N_11142);
nand U11256 (N_11256,N_10931,N_10870);
nand U11257 (N_11257,N_10981,N_10866);
and U11258 (N_11258,N_10807,N_11167);
and U11259 (N_11259,N_11113,N_10988);
nor U11260 (N_11260,N_11032,N_10875);
or U11261 (N_11261,N_11042,N_11003);
and U11262 (N_11262,N_10980,N_11117);
or U11263 (N_11263,N_11040,N_11197);
and U11264 (N_11264,N_10970,N_11090);
and U11265 (N_11265,N_10826,N_10959);
nor U11266 (N_11266,N_10823,N_11046);
nand U11267 (N_11267,N_11140,N_10883);
nand U11268 (N_11268,N_10938,N_11094);
or U11269 (N_11269,N_10928,N_11089);
xor U11270 (N_11270,N_11129,N_10885);
and U11271 (N_11271,N_11084,N_10987);
and U11272 (N_11272,N_10911,N_10984);
and U11273 (N_11273,N_10856,N_10921);
and U11274 (N_11274,N_11078,N_11004);
or U11275 (N_11275,N_11149,N_10806);
or U11276 (N_11276,N_11017,N_11128);
and U11277 (N_11277,N_10936,N_11121);
nand U11278 (N_11278,N_11099,N_11102);
nor U11279 (N_11279,N_11188,N_10979);
nor U11280 (N_11280,N_11006,N_10977);
nand U11281 (N_11281,N_10814,N_11199);
and U11282 (N_11282,N_11164,N_10805);
or U11283 (N_11283,N_10884,N_11105);
nor U11284 (N_11284,N_10966,N_11120);
nand U11285 (N_11285,N_10963,N_10934);
xor U11286 (N_11286,N_11027,N_11012);
or U11287 (N_11287,N_10930,N_11115);
and U11288 (N_11288,N_10975,N_10834);
and U11289 (N_11289,N_10802,N_10889);
nor U11290 (N_11290,N_10896,N_10973);
nand U11291 (N_11291,N_11092,N_11157);
nand U11292 (N_11292,N_10840,N_10837);
xor U11293 (N_11293,N_11138,N_11190);
nand U11294 (N_11294,N_10897,N_11178);
nand U11295 (N_11295,N_10874,N_11192);
or U11296 (N_11296,N_11074,N_10898);
nor U11297 (N_11297,N_10809,N_11160);
nor U11298 (N_11298,N_10869,N_10843);
nor U11299 (N_11299,N_11111,N_10960);
nor U11300 (N_11300,N_10888,N_10914);
or U11301 (N_11301,N_10957,N_11143);
nor U11302 (N_11302,N_10842,N_10945);
nor U11303 (N_11303,N_11080,N_10818);
nand U11304 (N_11304,N_11131,N_11191);
nor U11305 (N_11305,N_11127,N_10964);
or U11306 (N_11306,N_11169,N_11195);
and U11307 (N_11307,N_10998,N_10904);
nand U11308 (N_11308,N_10865,N_11193);
nor U11309 (N_11309,N_11182,N_10854);
nand U11310 (N_11310,N_10848,N_10893);
nand U11311 (N_11311,N_10941,N_10821);
nor U11312 (N_11312,N_11055,N_10999);
and U11313 (N_11313,N_10919,N_11033);
and U11314 (N_11314,N_11114,N_11075);
nand U11315 (N_11315,N_10876,N_11058);
nand U11316 (N_11316,N_11062,N_10812);
and U11317 (N_11317,N_11053,N_11172);
nand U11318 (N_11318,N_11010,N_10920);
or U11319 (N_11319,N_10918,N_10857);
nand U11320 (N_11320,N_11176,N_10860);
nand U11321 (N_11321,N_10852,N_11036);
or U11322 (N_11322,N_11168,N_11098);
nand U11323 (N_11323,N_11020,N_11045);
and U11324 (N_11324,N_10942,N_10909);
nor U11325 (N_11325,N_11022,N_11147);
and U11326 (N_11326,N_11002,N_10910);
xor U11327 (N_11327,N_10986,N_10993);
or U11328 (N_11328,N_10947,N_11001);
or U11329 (N_11329,N_10907,N_11021);
nor U11330 (N_11330,N_10946,N_11146);
nand U11331 (N_11331,N_11034,N_10996);
and U11332 (N_11332,N_11061,N_10968);
nand U11333 (N_11333,N_10828,N_11014);
or U11334 (N_11334,N_11082,N_10926);
nor U11335 (N_11335,N_10899,N_11063);
nand U11336 (N_11336,N_10861,N_10873);
and U11337 (N_11337,N_11134,N_11043);
nor U11338 (N_11338,N_10830,N_11166);
nor U11339 (N_11339,N_10912,N_11039);
nor U11340 (N_11340,N_11081,N_11161);
or U11341 (N_11341,N_11156,N_11049);
nand U11342 (N_11342,N_11194,N_10813);
and U11343 (N_11343,N_11123,N_10890);
nor U11344 (N_11344,N_10937,N_10915);
and U11345 (N_11345,N_11008,N_11029);
or U11346 (N_11346,N_10961,N_10955);
or U11347 (N_11347,N_11088,N_11119);
and U11348 (N_11348,N_11028,N_10864);
nor U11349 (N_11349,N_11106,N_10841);
or U11350 (N_11350,N_11024,N_11109);
and U11351 (N_11351,N_11030,N_10908);
nor U11352 (N_11352,N_10927,N_10948);
and U11353 (N_11353,N_11079,N_11183);
nand U11354 (N_11354,N_10829,N_11091);
nor U11355 (N_11355,N_11085,N_11093);
nand U11356 (N_11356,N_11015,N_11180);
and U11357 (N_11357,N_10851,N_10954);
nor U11358 (N_11358,N_10900,N_10872);
and U11359 (N_11359,N_11158,N_11097);
or U11360 (N_11360,N_10839,N_10804);
and U11361 (N_11361,N_11044,N_11130);
or U11362 (N_11362,N_11154,N_11108);
and U11363 (N_11363,N_11009,N_10956);
and U11364 (N_11364,N_10892,N_10992);
and U11365 (N_11365,N_11116,N_10969);
nor U11366 (N_11366,N_11054,N_10923);
nor U11367 (N_11367,N_11150,N_10953);
nand U11368 (N_11368,N_10881,N_11148);
nand U11369 (N_11369,N_11077,N_11103);
nor U11370 (N_11370,N_10844,N_11196);
or U11371 (N_11371,N_10887,N_10924);
or U11372 (N_11372,N_11104,N_10925);
nand U11373 (N_11373,N_10808,N_11065);
nor U11374 (N_11374,N_10903,N_11026);
and U11375 (N_11375,N_10976,N_11000);
nand U11376 (N_11376,N_10972,N_11023);
nor U11377 (N_11377,N_11162,N_10929);
nor U11378 (N_11378,N_10943,N_10994);
nand U11379 (N_11379,N_11155,N_11050);
xnor U11380 (N_11380,N_10933,N_11165);
or U11381 (N_11381,N_11173,N_10832);
nand U11382 (N_11382,N_10895,N_11107);
xor U11383 (N_11383,N_11016,N_10997);
and U11384 (N_11384,N_10817,N_11071);
or U11385 (N_11385,N_11051,N_10944);
or U11386 (N_11386,N_10880,N_10962);
or U11387 (N_11387,N_11070,N_10902);
and U11388 (N_11388,N_10974,N_10950);
or U11389 (N_11389,N_10859,N_10849);
nor U11390 (N_11390,N_11059,N_10846);
nand U11391 (N_11391,N_10982,N_11139);
nand U11392 (N_11392,N_11035,N_10965);
nor U11393 (N_11393,N_11185,N_10877);
or U11394 (N_11394,N_10833,N_11145);
or U11395 (N_11395,N_10855,N_11163);
or U11396 (N_11396,N_11031,N_10886);
or U11397 (N_11397,N_10917,N_10810);
nor U11398 (N_11398,N_11112,N_11068);
nand U11399 (N_11399,N_11064,N_11133);
or U11400 (N_11400,N_10832,N_10900);
nand U11401 (N_11401,N_11062,N_10905);
and U11402 (N_11402,N_10994,N_10828);
xnor U11403 (N_11403,N_11089,N_10898);
nor U11404 (N_11404,N_10827,N_10891);
or U11405 (N_11405,N_10901,N_10896);
nand U11406 (N_11406,N_10996,N_11147);
nand U11407 (N_11407,N_11139,N_10828);
and U11408 (N_11408,N_11018,N_11114);
or U11409 (N_11409,N_10895,N_11088);
and U11410 (N_11410,N_11145,N_11108);
or U11411 (N_11411,N_10931,N_10972);
and U11412 (N_11412,N_10975,N_11055);
or U11413 (N_11413,N_10898,N_11024);
nand U11414 (N_11414,N_11109,N_10845);
or U11415 (N_11415,N_10894,N_11109);
and U11416 (N_11416,N_10872,N_10914);
and U11417 (N_11417,N_11164,N_10984);
and U11418 (N_11418,N_11012,N_11110);
nor U11419 (N_11419,N_10980,N_10918);
or U11420 (N_11420,N_11122,N_11156);
or U11421 (N_11421,N_10807,N_11188);
nor U11422 (N_11422,N_10909,N_10887);
nand U11423 (N_11423,N_10961,N_11137);
nand U11424 (N_11424,N_11098,N_11190);
and U11425 (N_11425,N_11063,N_10998);
and U11426 (N_11426,N_11056,N_10915);
or U11427 (N_11427,N_10932,N_11100);
or U11428 (N_11428,N_11004,N_10863);
nand U11429 (N_11429,N_10832,N_11185);
nor U11430 (N_11430,N_10817,N_10864);
and U11431 (N_11431,N_10828,N_11072);
or U11432 (N_11432,N_11053,N_10993);
nand U11433 (N_11433,N_11198,N_11125);
nand U11434 (N_11434,N_10905,N_11134);
or U11435 (N_11435,N_11112,N_10825);
or U11436 (N_11436,N_11103,N_11005);
nand U11437 (N_11437,N_11016,N_10929);
nand U11438 (N_11438,N_10833,N_10890);
xor U11439 (N_11439,N_10827,N_10973);
nor U11440 (N_11440,N_10866,N_10843);
nand U11441 (N_11441,N_10928,N_11129);
nor U11442 (N_11442,N_11039,N_10997);
or U11443 (N_11443,N_10870,N_11080);
and U11444 (N_11444,N_10917,N_10842);
nand U11445 (N_11445,N_11180,N_10958);
or U11446 (N_11446,N_11114,N_10997);
nor U11447 (N_11447,N_10970,N_10877);
nor U11448 (N_11448,N_11026,N_11048);
or U11449 (N_11449,N_10976,N_11006);
nor U11450 (N_11450,N_10866,N_11189);
and U11451 (N_11451,N_11184,N_11156);
nand U11452 (N_11452,N_10802,N_11183);
and U11453 (N_11453,N_11029,N_10880);
and U11454 (N_11454,N_10967,N_10877);
or U11455 (N_11455,N_11005,N_10801);
and U11456 (N_11456,N_10805,N_11138);
and U11457 (N_11457,N_11052,N_11102);
nor U11458 (N_11458,N_11095,N_10899);
nor U11459 (N_11459,N_10849,N_10936);
or U11460 (N_11460,N_11088,N_11021);
and U11461 (N_11461,N_11160,N_10841);
or U11462 (N_11462,N_11015,N_10933);
nor U11463 (N_11463,N_10995,N_10992);
and U11464 (N_11464,N_10965,N_11145);
nor U11465 (N_11465,N_11096,N_10953);
nor U11466 (N_11466,N_11036,N_11166);
nor U11467 (N_11467,N_10905,N_11138);
or U11468 (N_11468,N_11097,N_10898);
or U11469 (N_11469,N_11050,N_11186);
nor U11470 (N_11470,N_11039,N_10865);
and U11471 (N_11471,N_10816,N_10991);
nor U11472 (N_11472,N_11051,N_10806);
nand U11473 (N_11473,N_10885,N_10858);
nand U11474 (N_11474,N_10895,N_11100);
or U11475 (N_11475,N_10849,N_11015);
or U11476 (N_11476,N_10935,N_11002);
xnor U11477 (N_11477,N_10907,N_10911);
nor U11478 (N_11478,N_11164,N_10830);
and U11479 (N_11479,N_11073,N_10863);
nand U11480 (N_11480,N_10952,N_10870);
or U11481 (N_11481,N_11016,N_11123);
nor U11482 (N_11482,N_11081,N_11101);
and U11483 (N_11483,N_10925,N_11137);
nor U11484 (N_11484,N_10922,N_11058);
and U11485 (N_11485,N_10962,N_11024);
nand U11486 (N_11486,N_10933,N_11160);
or U11487 (N_11487,N_11101,N_10949);
and U11488 (N_11488,N_11065,N_11096);
nand U11489 (N_11489,N_10840,N_11164);
nand U11490 (N_11490,N_10978,N_11043);
and U11491 (N_11491,N_11096,N_10876);
nand U11492 (N_11492,N_10872,N_11122);
nor U11493 (N_11493,N_10983,N_11008);
and U11494 (N_11494,N_11084,N_11129);
or U11495 (N_11495,N_11132,N_10948);
nand U11496 (N_11496,N_10927,N_11015);
nor U11497 (N_11497,N_11091,N_10918);
or U11498 (N_11498,N_11152,N_11195);
nand U11499 (N_11499,N_11156,N_10962);
or U11500 (N_11500,N_10820,N_10971);
nand U11501 (N_11501,N_11028,N_10834);
nand U11502 (N_11502,N_10869,N_10927);
or U11503 (N_11503,N_10938,N_10965);
nand U11504 (N_11504,N_11077,N_10965);
or U11505 (N_11505,N_11064,N_11046);
and U11506 (N_11506,N_11172,N_10940);
or U11507 (N_11507,N_11174,N_11076);
or U11508 (N_11508,N_11166,N_10829);
nand U11509 (N_11509,N_11160,N_11070);
nand U11510 (N_11510,N_11001,N_11175);
or U11511 (N_11511,N_11001,N_10803);
nor U11512 (N_11512,N_11148,N_10923);
and U11513 (N_11513,N_10906,N_11058);
nand U11514 (N_11514,N_10874,N_10982);
nor U11515 (N_11515,N_11021,N_11033);
nor U11516 (N_11516,N_10893,N_10960);
and U11517 (N_11517,N_10802,N_11156);
and U11518 (N_11518,N_11023,N_11199);
and U11519 (N_11519,N_11038,N_11117);
and U11520 (N_11520,N_11151,N_11081);
and U11521 (N_11521,N_11136,N_10963);
nand U11522 (N_11522,N_11118,N_10897);
nand U11523 (N_11523,N_11167,N_11142);
or U11524 (N_11524,N_10869,N_10900);
and U11525 (N_11525,N_10927,N_11132);
or U11526 (N_11526,N_10824,N_10846);
nand U11527 (N_11527,N_11050,N_11018);
nand U11528 (N_11528,N_11003,N_10852);
nor U11529 (N_11529,N_10977,N_10886);
nor U11530 (N_11530,N_11099,N_11114);
nor U11531 (N_11531,N_11015,N_11082);
and U11532 (N_11532,N_11110,N_11099);
or U11533 (N_11533,N_11084,N_11050);
and U11534 (N_11534,N_11039,N_11054);
nor U11535 (N_11535,N_11151,N_11146);
nand U11536 (N_11536,N_10889,N_11123);
nor U11537 (N_11537,N_10929,N_11185);
nor U11538 (N_11538,N_11098,N_11071);
nor U11539 (N_11539,N_10850,N_11173);
or U11540 (N_11540,N_10920,N_10956);
and U11541 (N_11541,N_10908,N_10986);
or U11542 (N_11542,N_11005,N_11167);
nor U11543 (N_11543,N_11187,N_10945);
nand U11544 (N_11544,N_11074,N_11182);
nand U11545 (N_11545,N_10891,N_11091);
or U11546 (N_11546,N_11120,N_11055);
nand U11547 (N_11547,N_10992,N_11040);
or U11548 (N_11548,N_10976,N_10876);
nor U11549 (N_11549,N_10862,N_10974);
or U11550 (N_11550,N_11052,N_11001);
xor U11551 (N_11551,N_11082,N_10824);
nor U11552 (N_11552,N_11102,N_10886);
nor U11553 (N_11553,N_11013,N_10984);
nor U11554 (N_11554,N_10936,N_10829);
or U11555 (N_11555,N_11175,N_11017);
and U11556 (N_11556,N_11023,N_10872);
nor U11557 (N_11557,N_11192,N_10931);
and U11558 (N_11558,N_11003,N_11199);
nor U11559 (N_11559,N_10954,N_11071);
nand U11560 (N_11560,N_10990,N_10802);
nand U11561 (N_11561,N_10804,N_10945);
nand U11562 (N_11562,N_10943,N_11067);
and U11563 (N_11563,N_10835,N_11151);
and U11564 (N_11564,N_10898,N_10865);
nand U11565 (N_11565,N_10861,N_11109);
and U11566 (N_11566,N_11186,N_10982);
and U11567 (N_11567,N_10966,N_10921);
nand U11568 (N_11568,N_11102,N_11008);
nand U11569 (N_11569,N_11008,N_11192);
or U11570 (N_11570,N_10859,N_10897);
and U11571 (N_11571,N_10987,N_10841);
nor U11572 (N_11572,N_11093,N_10852);
and U11573 (N_11573,N_10953,N_10982);
nor U11574 (N_11574,N_11053,N_10997);
nand U11575 (N_11575,N_11100,N_11141);
or U11576 (N_11576,N_10982,N_11088);
or U11577 (N_11577,N_10812,N_10891);
and U11578 (N_11578,N_11125,N_11070);
nand U11579 (N_11579,N_10925,N_11102);
nor U11580 (N_11580,N_11189,N_10925);
and U11581 (N_11581,N_10831,N_11180);
or U11582 (N_11582,N_11121,N_10906);
or U11583 (N_11583,N_11109,N_10929);
xnor U11584 (N_11584,N_10947,N_10987);
nor U11585 (N_11585,N_10920,N_11152);
nor U11586 (N_11586,N_10852,N_10904);
nor U11587 (N_11587,N_11090,N_10950);
and U11588 (N_11588,N_11092,N_11171);
or U11589 (N_11589,N_10958,N_10967);
or U11590 (N_11590,N_11175,N_11144);
and U11591 (N_11591,N_10977,N_11023);
nor U11592 (N_11592,N_10977,N_10852);
or U11593 (N_11593,N_10927,N_10943);
nand U11594 (N_11594,N_11141,N_11093);
nor U11595 (N_11595,N_11080,N_10874);
nor U11596 (N_11596,N_11111,N_11019);
nand U11597 (N_11597,N_10858,N_11192);
nand U11598 (N_11598,N_10852,N_10877);
or U11599 (N_11599,N_10962,N_11105);
and U11600 (N_11600,N_11355,N_11330);
or U11601 (N_11601,N_11254,N_11221);
and U11602 (N_11602,N_11400,N_11259);
nor U11603 (N_11603,N_11404,N_11308);
or U11604 (N_11604,N_11206,N_11244);
and U11605 (N_11605,N_11504,N_11530);
or U11606 (N_11606,N_11305,N_11352);
nand U11607 (N_11607,N_11487,N_11285);
or U11608 (N_11608,N_11324,N_11433);
nor U11609 (N_11609,N_11593,N_11312);
and U11610 (N_11610,N_11439,N_11597);
or U11611 (N_11611,N_11226,N_11223);
nand U11612 (N_11612,N_11260,N_11576);
and U11613 (N_11613,N_11202,N_11574);
or U11614 (N_11614,N_11451,N_11389);
and U11615 (N_11615,N_11559,N_11539);
nor U11616 (N_11616,N_11271,N_11314);
and U11617 (N_11617,N_11429,N_11533);
or U11618 (N_11618,N_11449,N_11387);
nand U11619 (N_11619,N_11476,N_11291);
nand U11620 (N_11620,N_11544,N_11479);
nor U11621 (N_11621,N_11458,N_11380);
nor U11622 (N_11622,N_11201,N_11397);
nor U11623 (N_11623,N_11456,N_11251);
or U11624 (N_11624,N_11266,N_11339);
nand U11625 (N_11625,N_11300,N_11406);
and U11626 (N_11626,N_11495,N_11463);
nand U11627 (N_11627,N_11445,N_11467);
nand U11628 (N_11628,N_11407,N_11493);
nor U11629 (N_11629,N_11513,N_11343);
or U11630 (N_11630,N_11516,N_11503);
or U11631 (N_11631,N_11542,N_11419);
nor U11632 (N_11632,N_11425,N_11359);
nor U11633 (N_11633,N_11470,N_11519);
and U11634 (N_11634,N_11273,N_11410);
and U11635 (N_11635,N_11486,N_11340);
nand U11636 (N_11636,N_11210,N_11537);
or U11637 (N_11637,N_11284,N_11394);
nor U11638 (N_11638,N_11520,N_11306);
and U11639 (N_11639,N_11379,N_11596);
nand U11640 (N_11640,N_11497,N_11220);
nand U11641 (N_11641,N_11346,N_11408);
and U11642 (N_11642,N_11437,N_11211);
nor U11643 (N_11643,N_11462,N_11442);
or U11644 (N_11644,N_11573,N_11491);
nor U11645 (N_11645,N_11317,N_11413);
and U11646 (N_11646,N_11207,N_11534);
nor U11647 (N_11647,N_11233,N_11238);
or U11648 (N_11648,N_11370,N_11447);
nor U11649 (N_11649,N_11547,N_11357);
and U11650 (N_11650,N_11468,N_11351);
nand U11651 (N_11651,N_11332,N_11358);
nor U11652 (N_11652,N_11292,N_11554);
nor U11653 (N_11653,N_11327,N_11241);
nand U11654 (N_11654,N_11441,N_11325);
nand U11655 (N_11655,N_11381,N_11489);
nand U11656 (N_11656,N_11274,N_11235);
and U11657 (N_11657,N_11249,N_11423);
nand U11658 (N_11658,N_11286,N_11364);
nand U11659 (N_11659,N_11320,N_11420);
nand U11660 (N_11660,N_11309,N_11382);
and U11661 (N_11661,N_11572,N_11371);
and U11662 (N_11662,N_11552,N_11250);
or U11663 (N_11663,N_11555,N_11374);
nor U11664 (N_11664,N_11322,N_11548);
or U11665 (N_11665,N_11248,N_11512);
nand U11666 (N_11666,N_11477,N_11511);
and U11667 (N_11667,N_11452,N_11577);
nand U11668 (N_11668,N_11589,N_11427);
and U11669 (N_11669,N_11390,N_11569);
nand U11670 (N_11670,N_11252,N_11281);
nor U11671 (N_11671,N_11313,N_11277);
nor U11672 (N_11672,N_11328,N_11229);
nand U11673 (N_11673,N_11236,N_11564);
or U11674 (N_11674,N_11438,N_11599);
and U11675 (N_11675,N_11298,N_11480);
nor U11676 (N_11676,N_11311,N_11431);
nor U11677 (N_11677,N_11591,N_11461);
and U11678 (N_11678,N_11301,N_11414);
nor U11679 (N_11679,N_11475,N_11335);
nor U11680 (N_11680,N_11218,N_11347);
and U11681 (N_11681,N_11490,N_11570);
or U11682 (N_11682,N_11526,N_11436);
nor U11683 (N_11683,N_11543,N_11538);
nand U11684 (N_11684,N_11556,N_11455);
nor U11685 (N_11685,N_11209,N_11278);
and U11686 (N_11686,N_11588,N_11293);
and U11687 (N_11687,N_11230,N_11416);
nor U11688 (N_11688,N_11453,N_11345);
and U11689 (N_11689,N_11510,N_11567);
or U11690 (N_11690,N_11213,N_11337);
or U11691 (N_11691,N_11578,N_11483);
and U11692 (N_11692,N_11246,N_11203);
nor U11693 (N_11693,N_11227,N_11532);
nor U11694 (N_11694,N_11466,N_11415);
nand U11695 (N_11695,N_11469,N_11217);
and U11696 (N_11696,N_11336,N_11396);
nand U11697 (N_11697,N_11372,N_11446);
and U11698 (N_11698,N_11256,N_11296);
or U11699 (N_11699,N_11257,N_11258);
or U11700 (N_11700,N_11460,N_11360);
and U11701 (N_11701,N_11212,N_11540);
and U11702 (N_11702,N_11454,N_11498);
nor U11703 (N_11703,N_11316,N_11272);
and U11704 (N_11704,N_11386,N_11571);
and U11705 (N_11705,N_11354,N_11523);
nor U11706 (N_11706,N_11377,N_11344);
and U11707 (N_11707,N_11443,N_11541);
or U11708 (N_11708,N_11261,N_11373);
nand U11709 (N_11709,N_11485,N_11517);
nand U11710 (N_11710,N_11240,N_11398);
and U11711 (N_11711,N_11402,N_11412);
nand U11712 (N_11712,N_11598,N_11264);
nor U11713 (N_11713,N_11582,N_11518);
nor U11714 (N_11714,N_11204,N_11562);
nor U11715 (N_11715,N_11494,N_11424);
or U11716 (N_11716,N_11581,N_11349);
nor U11717 (N_11717,N_11592,N_11522);
or U11718 (N_11718,N_11385,N_11208);
nor U11719 (N_11719,N_11514,N_11275);
nor U11720 (N_11720,N_11393,N_11265);
nand U11721 (N_11721,N_11321,N_11580);
nand U11722 (N_11722,N_11383,N_11568);
or U11723 (N_11723,N_11488,N_11342);
or U11724 (N_11724,N_11392,N_11341);
or U11725 (N_11725,N_11585,N_11289);
and U11726 (N_11726,N_11500,N_11245);
and U11727 (N_11727,N_11575,N_11550);
or U11728 (N_11728,N_11524,N_11214);
nor U11729 (N_11729,N_11565,N_11269);
nand U11730 (N_11730,N_11561,N_11528);
or U11731 (N_11731,N_11361,N_11409);
nor U11732 (N_11732,N_11362,N_11465);
and U11733 (N_11733,N_11478,N_11403);
nor U11734 (N_11734,N_11366,N_11496);
and U11735 (N_11735,N_11302,N_11243);
nand U11736 (N_11736,N_11563,N_11560);
nand U11737 (N_11737,N_11376,N_11283);
or U11738 (N_11738,N_11237,N_11363);
or U11739 (N_11739,N_11215,N_11492);
and U11740 (N_11740,N_11267,N_11405);
and U11741 (N_11741,N_11457,N_11595);
and U11742 (N_11742,N_11551,N_11297);
nor U11743 (N_11743,N_11558,N_11557);
nor U11744 (N_11744,N_11444,N_11428);
or U11745 (N_11745,N_11587,N_11529);
and U11746 (N_11746,N_11432,N_11474);
nor U11747 (N_11747,N_11594,N_11280);
nand U11748 (N_11748,N_11234,N_11326);
nor U11749 (N_11749,N_11307,N_11279);
or U11750 (N_11750,N_11464,N_11287);
nor U11751 (N_11751,N_11531,N_11482);
or U11752 (N_11752,N_11319,N_11232);
nand U11753 (N_11753,N_11507,N_11276);
nand U11754 (N_11754,N_11239,N_11501);
and U11755 (N_11755,N_11348,N_11586);
or U11756 (N_11756,N_11481,N_11282);
or U11757 (N_11757,N_11448,N_11242);
nor U11758 (N_11758,N_11549,N_11472);
or U11759 (N_11759,N_11294,N_11459);
or U11760 (N_11760,N_11471,N_11536);
or U11761 (N_11761,N_11418,N_11499);
nand U11762 (N_11762,N_11417,N_11579);
or U11763 (N_11763,N_11521,N_11205);
and U11764 (N_11764,N_11401,N_11365);
and U11765 (N_11765,N_11224,N_11566);
or U11766 (N_11766,N_11535,N_11253);
nor U11767 (N_11767,N_11270,N_11262);
or U11768 (N_11768,N_11334,N_11315);
nor U11769 (N_11769,N_11421,N_11440);
or U11770 (N_11770,N_11545,N_11411);
nand U11771 (N_11771,N_11590,N_11525);
and U11772 (N_11772,N_11329,N_11502);
and U11773 (N_11773,N_11515,N_11268);
and U11774 (N_11774,N_11434,N_11304);
nor U11775 (N_11775,N_11583,N_11263);
or U11776 (N_11776,N_11200,N_11338);
and U11777 (N_11777,N_11225,N_11584);
or U11778 (N_11778,N_11399,N_11303);
nand U11779 (N_11779,N_11367,N_11353);
and U11780 (N_11780,N_11333,N_11422);
nand U11781 (N_11781,N_11231,N_11255);
and U11782 (N_11782,N_11378,N_11553);
nor U11783 (N_11783,N_11484,N_11222);
nand U11784 (N_11784,N_11391,N_11384);
nand U11785 (N_11785,N_11527,N_11310);
nand U11786 (N_11786,N_11450,N_11288);
nand U11787 (N_11787,N_11368,N_11473);
nor U11788 (N_11788,N_11216,N_11430);
nor U11789 (N_11789,N_11509,N_11247);
nand U11790 (N_11790,N_11395,N_11318);
nor U11791 (N_11791,N_11388,N_11219);
nand U11792 (N_11792,N_11331,N_11323);
and U11793 (N_11793,N_11435,N_11228);
nand U11794 (N_11794,N_11505,N_11506);
nand U11795 (N_11795,N_11426,N_11356);
nand U11796 (N_11796,N_11350,N_11295);
nand U11797 (N_11797,N_11290,N_11546);
or U11798 (N_11798,N_11375,N_11299);
and U11799 (N_11799,N_11508,N_11369);
and U11800 (N_11800,N_11463,N_11485);
and U11801 (N_11801,N_11218,N_11329);
nand U11802 (N_11802,N_11491,N_11206);
nand U11803 (N_11803,N_11318,N_11593);
nand U11804 (N_11804,N_11589,N_11416);
nor U11805 (N_11805,N_11475,N_11571);
or U11806 (N_11806,N_11275,N_11281);
nand U11807 (N_11807,N_11367,N_11246);
and U11808 (N_11808,N_11268,N_11585);
or U11809 (N_11809,N_11445,N_11200);
or U11810 (N_11810,N_11540,N_11219);
nand U11811 (N_11811,N_11293,N_11425);
and U11812 (N_11812,N_11456,N_11596);
and U11813 (N_11813,N_11248,N_11234);
and U11814 (N_11814,N_11418,N_11336);
and U11815 (N_11815,N_11581,N_11433);
and U11816 (N_11816,N_11326,N_11549);
and U11817 (N_11817,N_11519,N_11238);
and U11818 (N_11818,N_11244,N_11417);
nor U11819 (N_11819,N_11338,N_11519);
or U11820 (N_11820,N_11386,N_11596);
nor U11821 (N_11821,N_11501,N_11536);
nand U11822 (N_11822,N_11371,N_11462);
and U11823 (N_11823,N_11429,N_11263);
nor U11824 (N_11824,N_11243,N_11477);
nor U11825 (N_11825,N_11260,N_11259);
or U11826 (N_11826,N_11232,N_11567);
nor U11827 (N_11827,N_11317,N_11468);
or U11828 (N_11828,N_11265,N_11242);
and U11829 (N_11829,N_11376,N_11540);
and U11830 (N_11830,N_11247,N_11592);
and U11831 (N_11831,N_11316,N_11402);
nand U11832 (N_11832,N_11299,N_11520);
and U11833 (N_11833,N_11241,N_11518);
nor U11834 (N_11834,N_11446,N_11598);
nand U11835 (N_11835,N_11583,N_11355);
nor U11836 (N_11836,N_11372,N_11328);
or U11837 (N_11837,N_11360,N_11274);
nand U11838 (N_11838,N_11326,N_11518);
and U11839 (N_11839,N_11385,N_11302);
or U11840 (N_11840,N_11253,N_11460);
nor U11841 (N_11841,N_11579,N_11524);
nand U11842 (N_11842,N_11511,N_11261);
and U11843 (N_11843,N_11539,N_11598);
nand U11844 (N_11844,N_11400,N_11485);
and U11845 (N_11845,N_11452,N_11405);
and U11846 (N_11846,N_11274,N_11498);
nand U11847 (N_11847,N_11322,N_11293);
nand U11848 (N_11848,N_11578,N_11260);
nor U11849 (N_11849,N_11396,N_11397);
and U11850 (N_11850,N_11314,N_11325);
nand U11851 (N_11851,N_11420,N_11298);
and U11852 (N_11852,N_11299,N_11537);
nor U11853 (N_11853,N_11230,N_11466);
nor U11854 (N_11854,N_11268,N_11540);
nor U11855 (N_11855,N_11512,N_11241);
nand U11856 (N_11856,N_11318,N_11416);
or U11857 (N_11857,N_11292,N_11523);
and U11858 (N_11858,N_11521,N_11223);
or U11859 (N_11859,N_11484,N_11405);
or U11860 (N_11860,N_11514,N_11525);
and U11861 (N_11861,N_11274,N_11512);
nor U11862 (N_11862,N_11525,N_11478);
nor U11863 (N_11863,N_11202,N_11391);
nand U11864 (N_11864,N_11527,N_11463);
nor U11865 (N_11865,N_11296,N_11376);
nand U11866 (N_11866,N_11578,N_11347);
and U11867 (N_11867,N_11512,N_11358);
nor U11868 (N_11868,N_11297,N_11522);
and U11869 (N_11869,N_11280,N_11515);
nand U11870 (N_11870,N_11309,N_11384);
nand U11871 (N_11871,N_11498,N_11577);
nand U11872 (N_11872,N_11378,N_11498);
and U11873 (N_11873,N_11477,N_11312);
or U11874 (N_11874,N_11367,N_11384);
nor U11875 (N_11875,N_11239,N_11435);
and U11876 (N_11876,N_11259,N_11312);
and U11877 (N_11877,N_11307,N_11266);
and U11878 (N_11878,N_11590,N_11319);
nand U11879 (N_11879,N_11267,N_11414);
or U11880 (N_11880,N_11302,N_11472);
and U11881 (N_11881,N_11250,N_11353);
and U11882 (N_11882,N_11573,N_11402);
xor U11883 (N_11883,N_11327,N_11433);
or U11884 (N_11884,N_11260,N_11313);
nor U11885 (N_11885,N_11519,N_11594);
nand U11886 (N_11886,N_11498,N_11420);
nor U11887 (N_11887,N_11301,N_11352);
or U11888 (N_11888,N_11284,N_11545);
or U11889 (N_11889,N_11555,N_11248);
and U11890 (N_11890,N_11393,N_11336);
or U11891 (N_11891,N_11487,N_11357);
xnor U11892 (N_11892,N_11478,N_11256);
or U11893 (N_11893,N_11508,N_11211);
nand U11894 (N_11894,N_11240,N_11237);
nand U11895 (N_11895,N_11329,N_11248);
and U11896 (N_11896,N_11269,N_11446);
or U11897 (N_11897,N_11471,N_11408);
nor U11898 (N_11898,N_11382,N_11221);
and U11899 (N_11899,N_11535,N_11344);
nand U11900 (N_11900,N_11438,N_11351);
nor U11901 (N_11901,N_11512,N_11458);
or U11902 (N_11902,N_11470,N_11548);
nor U11903 (N_11903,N_11409,N_11349);
nor U11904 (N_11904,N_11209,N_11459);
nand U11905 (N_11905,N_11541,N_11317);
and U11906 (N_11906,N_11298,N_11337);
and U11907 (N_11907,N_11371,N_11350);
and U11908 (N_11908,N_11214,N_11576);
and U11909 (N_11909,N_11268,N_11349);
and U11910 (N_11910,N_11386,N_11458);
and U11911 (N_11911,N_11227,N_11447);
and U11912 (N_11912,N_11361,N_11358);
nand U11913 (N_11913,N_11327,N_11436);
nor U11914 (N_11914,N_11393,N_11489);
or U11915 (N_11915,N_11444,N_11249);
or U11916 (N_11916,N_11329,N_11569);
or U11917 (N_11917,N_11391,N_11345);
nor U11918 (N_11918,N_11427,N_11291);
or U11919 (N_11919,N_11567,N_11425);
and U11920 (N_11920,N_11471,N_11553);
nand U11921 (N_11921,N_11297,N_11435);
nor U11922 (N_11922,N_11216,N_11245);
nor U11923 (N_11923,N_11423,N_11298);
nor U11924 (N_11924,N_11477,N_11425);
or U11925 (N_11925,N_11240,N_11517);
and U11926 (N_11926,N_11399,N_11489);
and U11927 (N_11927,N_11574,N_11566);
nor U11928 (N_11928,N_11251,N_11537);
nand U11929 (N_11929,N_11443,N_11500);
nor U11930 (N_11930,N_11487,N_11272);
or U11931 (N_11931,N_11532,N_11427);
or U11932 (N_11932,N_11313,N_11228);
nand U11933 (N_11933,N_11468,N_11405);
and U11934 (N_11934,N_11268,N_11373);
nand U11935 (N_11935,N_11204,N_11229);
or U11936 (N_11936,N_11562,N_11578);
and U11937 (N_11937,N_11253,N_11292);
and U11938 (N_11938,N_11465,N_11205);
and U11939 (N_11939,N_11514,N_11437);
and U11940 (N_11940,N_11203,N_11457);
and U11941 (N_11941,N_11356,N_11339);
and U11942 (N_11942,N_11353,N_11237);
nor U11943 (N_11943,N_11286,N_11341);
or U11944 (N_11944,N_11471,N_11545);
and U11945 (N_11945,N_11580,N_11245);
nand U11946 (N_11946,N_11507,N_11231);
nor U11947 (N_11947,N_11482,N_11492);
nand U11948 (N_11948,N_11527,N_11490);
or U11949 (N_11949,N_11202,N_11463);
nor U11950 (N_11950,N_11229,N_11435);
or U11951 (N_11951,N_11200,N_11258);
and U11952 (N_11952,N_11425,N_11275);
and U11953 (N_11953,N_11318,N_11409);
or U11954 (N_11954,N_11249,N_11386);
or U11955 (N_11955,N_11387,N_11496);
and U11956 (N_11956,N_11508,N_11382);
nand U11957 (N_11957,N_11479,N_11459);
nand U11958 (N_11958,N_11336,N_11205);
nor U11959 (N_11959,N_11502,N_11256);
nor U11960 (N_11960,N_11534,N_11579);
nand U11961 (N_11961,N_11541,N_11323);
nor U11962 (N_11962,N_11293,N_11301);
nor U11963 (N_11963,N_11513,N_11288);
nor U11964 (N_11964,N_11388,N_11426);
or U11965 (N_11965,N_11310,N_11206);
and U11966 (N_11966,N_11504,N_11277);
nor U11967 (N_11967,N_11319,N_11583);
or U11968 (N_11968,N_11518,N_11426);
nor U11969 (N_11969,N_11258,N_11533);
and U11970 (N_11970,N_11554,N_11467);
and U11971 (N_11971,N_11302,N_11394);
and U11972 (N_11972,N_11486,N_11264);
nor U11973 (N_11973,N_11219,N_11599);
or U11974 (N_11974,N_11239,N_11461);
and U11975 (N_11975,N_11258,N_11284);
nor U11976 (N_11976,N_11444,N_11204);
nand U11977 (N_11977,N_11234,N_11453);
and U11978 (N_11978,N_11365,N_11546);
nor U11979 (N_11979,N_11558,N_11360);
nand U11980 (N_11980,N_11478,N_11221);
nand U11981 (N_11981,N_11531,N_11357);
and U11982 (N_11982,N_11333,N_11258);
nor U11983 (N_11983,N_11272,N_11491);
nand U11984 (N_11984,N_11561,N_11200);
or U11985 (N_11985,N_11415,N_11536);
and U11986 (N_11986,N_11522,N_11566);
or U11987 (N_11987,N_11307,N_11504);
and U11988 (N_11988,N_11298,N_11500);
nand U11989 (N_11989,N_11355,N_11353);
nand U11990 (N_11990,N_11261,N_11538);
or U11991 (N_11991,N_11280,N_11432);
and U11992 (N_11992,N_11280,N_11531);
or U11993 (N_11993,N_11569,N_11513);
or U11994 (N_11994,N_11301,N_11341);
nor U11995 (N_11995,N_11530,N_11219);
nor U11996 (N_11996,N_11388,N_11586);
nand U11997 (N_11997,N_11223,N_11487);
or U11998 (N_11998,N_11200,N_11439);
and U11999 (N_11999,N_11442,N_11494);
nor U12000 (N_12000,N_11909,N_11795);
or U12001 (N_12001,N_11894,N_11675);
or U12002 (N_12002,N_11661,N_11948);
nand U12003 (N_12003,N_11729,N_11707);
and U12004 (N_12004,N_11664,N_11834);
nand U12005 (N_12005,N_11907,N_11670);
nor U12006 (N_12006,N_11825,N_11954);
nand U12007 (N_12007,N_11897,N_11783);
nor U12008 (N_12008,N_11898,N_11865);
nand U12009 (N_12009,N_11977,N_11970);
nand U12010 (N_12010,N_11677,N_11787);
or U12011 (N_12011,N_11963,N_11690);
nand U12012 (N_12012,N_11790,N_11821);
nand U12013 (N_12013,N_11855,N_11934);
and U12014 (N_12014,N_11960,N_11867);
nand U12015 (N_12015,N_11702,N_11671);
and U12016 (N_12016,N_11940,N_11654);
and U12017 (N_12017,N_11765,N_11618);
and U12018 (N_12018,N_11725,N_11775);
or U12019 (N_12019,N_11818,N_11959);
nand U12020 (N_12020,N_11822,N_11622);
and U12021 (N_12021,N_11974,N_11657);
and U12022 (N_12022,N_11848,N_11924);
nand U12023 (N_12023,N_11711,N_11908);
or U12024 (N_12024,N_11992,N_11709);
or U12025 (N_12025,N_11852,N_11944);
and U12026 (N_12026,N_11806,N_11923);
or U12027 (N_12027,N_11910,N_11653);
nand U12028 (N_12028,N_11650,N_11824);
nor U12029 (N_12029,N_11995,N_11800);
nor U12030 (N_12030,N_11916,N_11745);
nand U12031 (N_12031,N_11856,N_11627);
and U12032 (N_12032,N_11912,N_11638);
and U12033 (N_12033,N_11836,N_11918);
nand U12034 (N_12034,N_11686,N_11639);
nand U12035 (N_12035,N_11864,N_11844);
nand U12036 (N_12036,N_11901,N_11764);
and U12037 (N_12037,N_11863,N_11648);
nor U12038 (N_12038,N_11724,N_11895);
or U12039 (N_12039,N_11920,N_11956);
nand U12040 (N_12040,N_11667,N_11733);
and U12041 (N_12041,N_11946,N_11643);
nand U12042 (N_12042,N_11830,N_11760);
or U12043 (N_12043,N_11708,N_11616);
or U12044 (N_12044,N_11750,N_11752);
nor U12045 (N_12045,N_11665,N_11973);
nor U12046 (N_12046,N_11820,N_11996);
or U12047 (N_12047,N_11826,N_11829);
and U12048 (N_12048,N_11942,N_11780);
nor U12049 (N_12049,N_11735,N_11939);
nor U12050 (N_12050,N_11936,N_11805);
nor U12051 (N_12051,N_11781,N_11635);
or U12052 (N_12052,N_11849,N_11982);
nor U12053 (N_12053,N_11857,N_11719);
nand U12054 (N_12054,N_11911,N_11990);
nor U12055 (N_12055,N_11727,N_11640);
and U12056 (N_12056,N_11641,N_11985);
nor U12057 (N_12057,N_11740,N_11603);
nand U12058 (N_12058,N_11943,N_11935);
and U12059 (N_12059,N_11986,N_11619);
nand U12060 (N_12060,N_11813,N_11791);
nand U12061 (N_12061,N_11634,N_11703);
nand U12062 (N_12062,N_11613,N_11947);
or U12063 (N_12063,N_11839,N_11718);
nand U12064 (N_12064,N_11621,N_11828);
nor U12065 (N_12065,N_11662,N_11833);
or U12066 (N_12066,N_11882,N_11652);
or U12067 (N_12067,N_11880,N_11681);
nand U12068 (N_12068,N_11971,N_11757);
and U12069 (N_12069,N_11815,N_11647);
or U12070 (N_12070,N_11927,N_11604);
or U12071 (N_12071,N_11792,N_11701);
or U12072 (N_12072,N_11810,N_11845);
nand U12073 (N_12073,N_11688,N_11890);
nand U12074 (N_12074,N_11770,N_11949);
or U12075 (N_12075,N_11788,N_11929);
and U12076 (N_12076,N_11628,N_11888);
nand U12077 (N_12077,N_11793,N_11987);
and U12078 (N_12078,N_11967,N_11840);
nand U12079 (N_12079,N_11704,N_11732);
or U12080 (N_12080,N_11605,N_11997);
nor U12081 (N_12081,N_11969,N_11789);
nand U12082 (N_12082,N_11877,N_11832);
nand U12083 (N_12083,N_11607,N_11769);
nor U12084 (N_12084,N_11905,N_11953);
nor U12085 (N_12085,N_11951,N_11819);
nand U12086 (N_12086,N_11958,N_11984);
nand U12087 (N_12087,N_11955,N_11767);
nand U12088 (N_12088,N_11649,N_11608);
nor U12089 (N_12089,N_11682,N_11779);
nand U12090 (N_12090,N_11957,N_11730);
or U12091 (N_12091,N_11873,N_11816);
nand U12092 (N_12092,N_11917,N_11919);
or U12093 (N_12093,N_11660,N_11705);
nor U12094 (N_12094,N_11642,N_11874);
and U12095 (N_12095,N_11876,N_11913);
and U12096 (N_12096,N_11978,N_11689);
nor U12097 (N_12097,N_11807,N_11797);
or U12098 (N_12098,N_11712,N_11858);
or U12099 (N_12099,N_11799,N_11734);
and U12100 (N_12100,N_11698,N_11674);
or U12101 (N_12101,N_11950,N_11902);
nand U12102 (N_12102,N_11827,N_11624);
nand U12103 (N_12103,N_11759,N_11843);
or U12104 (N_12104,N_11979,N_11636);
nand U12105 (N_12105,N_11786,N_11866);
and U12106 (N_12106,N_11926,N_11646);
nand U12107 (N_12107,N_11776,N_11742);
nor U12108 (N_12108,N_11714,N_11685);
nand U12109 (N_12109,N_11663,N_11758);
and U12110 (N_12110,N_11617,N_11630);
and U12111 (N_12111,N_11921,N_11717);
and U12112 (N_12112,N_11612,N_11842);
and U12113 (N_12113,N_11861,N_11893);
nand U12114 (N_12114,N_11726,N_11754);
nor U12115 (N_12115,N_11976,N_11771);
nor U12116 (N_12116,N_11886,N_11846);
or U12117 (N_12117,N_11904,N_11763);
nor U12118 (N_12118,N_11903,N_11747);
nor U12119 (N_12119,N_11965,N_11676);
or U12120 (N_12120,N_11772,N_11737);
nor U12121 (N_12121,N_11838,N_11964);
and U12122 (N_12122,N_11611,N_11785);
nor U12123 (N_12123,N_11610,N_11900);
nor U12124 (N_12124,N_11673,N_11989);
or U12125 (N_12125,N_11837,N_11802);
xor U12126 (N_12126,N_11645,N_11906);
nand U12127 (N_12127,N_11801,N_11966);
and U12128 (N_12128,N_11716,N_11869);
nor U12129 (N_12129,N_11669,N_11835);
or U12130 (N_12130,N_11988,N_11739);
and U12131 (N_12131,N_11961,N_11656);
or U12132 (N_12132,N_11931,N_11854);
nand U12133 (N_12133,N_11975,N_11887);
or U12134 (N_12134,N_11879,N_11631);
nor U12135 (N_12135,N_11922,N_11778);
and U12136 (N_12136,N_11694,N_11614);
or U12137 (N_12137,N_11892,N_11762);
nand U12138 (N_12138,N_11672,N_11875);
nor U12139 (N_12139,N_11626,N_11766);
nand U12140 (N_12140,N_11796,N_11687);
or U12141 (N_12141,N_11755,N_11868);
nand U12142 (N_12142,N_11655,N_11808);
nand U12143 (N_12143,N_11889,N_11881);
and U12144 (N_12144,N_11683,N_11883);
and U12145 (N_12145,N_11720,N_11722);
or U12146 (N_12146,N_11993,N_11850);
nand U12147 (N_12147,N_11713,N_11695);
or U12148 (N_12148,N_11710,N_11700);
and U12149 (N_12149,N_11847,N_11633);
nand U12150 (N_12150,N_11817,N_11715);
nor U12151 (N_12151,N_11684,N_11862);
or U12152 (N_12152,N_11600,N_11666);
and U12153 (N_12153,N_11831,N_11999);
nor U12154 (N_12154,N_11915,N_11798);
or U12155 (N_12155,N_11878,N_11678);
nor U12156 (N_12156,N_11812,N_11644);
nand U12157 (N_12157,N_11823,N_11841);
or U12158 (N_12158,N_11738,N_11991);
xnor U12159 (N_12159,N_11659,N_11615);
or U12160 (N_12160,N_11896,N_11851);
nand U12161 (N_12161,N_11870,N_11761);
and U12162 (N_12162,N_11743,N_11744);
and U12163 (N_12163,N_11928,N_11637);
or U12164 (N_12164,N_11891,N_11692);
and U12165 (N_12165,N_11809,N_11602);
and U12166 (N_12166,N_11803,N_11629);
and U12167 (N_12167,N_11968,N_11691);
and U12168 (N_12168,N_11623,N_11699);
and U12169 (N_12169,N_11625,N_11937);
or U12170 (N_12170,N_11751,N_11723);
nor U12171 (N_12171,N_11784,N_11768);
and U12172 (N_12172,N_11774,N_11632);
and U12173 (N_12173,N_11693,N_11620);
or U12174 (N_12174,N_11804,N_11914);
nor U12175 (N_12175,N_11668,N_11860);
and U12176 (N_12176,N_11601,N_11930);
nand U12177 (N_12177,N_11938,N_11983);
nand U12178 (N_12178,N_11952,N_11756);
or U12179 (N_12179,N_11859,N_11728);
nand U12180 (N_12180,N_11932,N_11885);
nand U12181 (N_12181,N_11980,N_11736);
and U12182 (N_12182,N_11962,N_11933);
nor U12183 (N_12183,N_11696,N_11899);
or U12184 (N_12184,N_11871,N_11794);
and U12185 (N_12185,N_11782,N_11680);
xnor U12186 (N_12186,N_11753,N_11777);
and U12187 (N_12187,N_11814,N_11741);
and U12188 (N_12188,N_11941,N_11697);
and U12189 (N_12189,N_11998,N_11811);
or U12190 (N_12190,N_11706,N_11721);
nand U12191 (N_12191,N_11972,N_11679);
or U12192 (N_12192,N_11884,N_11853);
and U12193 (N_12193,N_11731,N_11749);
nor U12194 (N_12194,N_11981,N_11945);
nor U12195 (N_12195,N_11773,N_11606);
nor U12196 (N_12196,N_11651,N_11746);
nand U12197 (N_12197,N_11748,N_11925);
nand U12198 (N_12198,N_11609,N_11872);
nor U12199 (N_12199,N_11658,N_11994);
and U12200 (N_12200,N_11706,N_11838);
nand U12201 (N_12201,N_11909,N_11650);
nand U12202 (N_12202,N_11873,N_11740);
nand U12203 (N_12203,N_11600,N_11731);
nand U12204 (N_12204,N_11629,N_11672);
nor U12205 (N_12205,N_11711,N_11702);
nor U12206 (N_12206,N_11827,N_11851);
nand U12207 (N_12207,N_11982,N_11990);
and U12208 (N_12208,N_11797,N_11831);
nor U12209 (N_12209,N_11793,N_11606);
nor U12210 (N_12210,N_11791,N_11832);
nand U12211 (N_12211,N_11924,N_11738);
and U12212 (N_12212,N_11667,N_11916);
or U12213 (N_12213,N_11900,N_11779);
nor U12214 (N_12214,N_11974,N_11724);
and U12215 (N_12215,N_11924,N_11767);
and U12216 (N_12216,N_11624,N_11636);
or U12217 (N_12217,N_11728,N_11976);
nor U12218 (N_12218,N_11793,N_11648);
and U12219 (N_12219,N_11908,N_11825);
nor U12220 (N_12220,N_11959,N_11948);
and U12221 (N_12221,N_11902,N_11917);
and U12222 (N_12222,N_11719,N_11706);
nor U12223 (N_12223,N_11832,N_11689);
nand U12224 (N_12224,N_11831,N_11615);
or U12225 (N_12225,N_11786,N_11988);
and U12226 (N_12226,N_11757,N_11968);
or U12227 (N_12227,N_11662,N_11829);
nor U12228 (N_12228,N_11891,N_11958);
or U12229 (N_12229,N_11698,N_11726);
or U12230 (N_12230,N_11727,N_11662);
and U12231 (N_12231,N_11945,N_11765);
and U12232 (N_12232,N_11967,N_11703);
nand U12233 (N_12233,N_11687,N_11754);
nand U12234 (N_12234,N_11817,N_11658);
and U12235 (N_12235,N_11645,N_11828);
nor U12236 (N_12236,N_11875,N_11709);
and U12237 (N_12237,N_11814,N_11908);
nor U12238 (N_12238,N_11675,N_11965);
nor U12239 (N_12239,N_11976,N_11930);
nand U12240 (N_12240,N_11864,N_11693);
nand U12241 (N_12241,N_11845,N_11694);
and U12242 (N_12242,N_11756,N_11844);
xor U12243 (N_12243,N_11917,N_11800);
nor U12244 (N_12244,N_11838,N_11746);
nand U12245 (N_12245,N_11689,N_11890);
nand U12246 (N_12246,N_11683,N_11759);
nand U12247 (N_12247,N_11691,N_11742);
or U12248 (N_12248,N_11952,N_11605);
nand U12249 (N_12249,N_11892,N_11850);
nand U12250 (N_12250,N_11829,N_11943);
and U12251 (N_12251,N_11882,N_11952);
and U12252 (N_12252,N_11991,N_11903);
or U12253 (N_12253,N_11631,N_11689);
nor U12254 (N_12254,N_11738,N_11863);
or U12255 (N_12255,N_11906,N_11776);
and U12256 (N_12256,N_11996,N_11889);
nand U12257 (N_12257,N_11931,N_11707);
nor U12258 (N_12258,N_11617,N_11661);
nor U12259 (N_12259,N_11618,N_11606);
or U12260 (N_12260,N_11681,N_11840);
nor U12261 (N_12261,N_11775,N_11691);
nor U12262 (N_12262,N_11857,N_11607);
or U12263 (N_12263,N_11903,N_11992);
or U12264 (N_12264,N_11626,N_11952);
nor U12265 (N_12265,N_11793,N_11985);
nand U12266 (N_12266,N_11700,N_11946);
nor U12267 (N_12267,N_11678,N_11926);
nor U12268 (N_12268,N_11660,N_11631);
or U12269 (N_12269,N_11807,N_11645);
or U12270 (N_12270,N_11940,N_11718);
or U12271 (N_12271,N_11759,N_11741);
and U12272 (N_12272,N_11866,N_11808);
nor U12273 (N_12273,N_11892,N_11921);
nor U12274 (N_12274,N_11964,N_11914);
nand U12275 (N_12275,N_11837,N_11967);
and U12276 (N_12276,N_11753,N_11949);
nand U12277 (N_12277,N_11610,N_11884);
nand U12278 (N_12278,N_11744,N_11617);
nand U12279 (N_12279,N_11724,N_11721);
and U12280 (N_12280,N_11878,N_11754);
nor U12281 (N_12281,N_11723,N_11918);
nand U12282 (N_12282,N_11978,N_11881);
or U12283 (N_12283,N_11970,N_11824);
or U12284 (N_12284,N_11759,N_11795);
nor U12285 (N_12285,N_11884,N_11956);
or U12286 (N_12286,N_11831,N_11697);
or U12287 (N_12287,N_11617,N_11729);
nand U12288 (N_12288,N_11838,N_11942);
or U12289 (N_12289,N_11743,N_11992);
nand U12290 (N_12290,N_11794,N_11683);
and U12291 (N_12291,N_11764,N_11685);
nand U12292 (N_12292,N_11719,N_11702);
or U12293 (N_12293,N_11672,N_11745);
nand U12294 (N_12294,N_11794,N_11868);
nand U12295 (N_12295,N_11779,N_11766);
nor U12296 (N_12296,N_11894,N_11757);
nand U12297 (N_12297,N_11838,N_11604);
or U12298 (N_12298,N_11953,N_11821);
nor U12299 (N_12299,N_11948,N_11736);
nand U12300 (N_12300,N_11926,N_11897);
or U12301 (N_12301,N_11889,N_11948);
nand U12302 (N_12302,N_11762,N_11642);
nor U12303 (N_12303,N_11799,N_11702);
or U12304 (N_12304,N_11763,N_11949);
and U12305 (N_12305,N_11682,N_11896);
and U12306 (N_12306,N_11733,N_11937);
nand U12307 (N_12307,N_11653,N_11993);
or U12308 (N_12308,N_11686,N_11633);
or U12309 (N_12309,N_11932,N_11956);
nand U12310 (N_12310,N_11658,N_11735);
or U12311 (N_12311,N_11629,N_11948);
nor U12312 (N_12312,N_11698,N_11936);
nor U12313 (N_12313,N_11966,N_11609);
or U12314 (N_12314,N_11722,N_11725);
and U12315 (N_12315,N_11852,N_11922);
nor U12316 (N_12316,N_11764,N_11748);
nor U12317 (N_12317,N_11852,N_11865);
or U12318 (N_12318,N_11964,N_11814);
or U12319 (N_12319,N_11698,N_11873);
nor U12320 (N_12320,N_11793,N_11803);
nand U12321 (N_12321,N_11862,N_11819);
nor U12322 (N_12322,N_11916,N_11840);
or U12323 (N_12323,N_11964,N_11982);
and U12324 (N_12324,N_11811,N_11711);
and U12325 (N_12325,N_11622,N_11629);
nor U12326 (N_12326,N_11846,N_11949);
or U12327 (N_12327,N_11752,N_11888);
nand U12328 (N_12328,N_11711,N_11603);
or U12329 (N_12329,N_11826,N_11815);
nand U12330 (N_12330,N_11882,N_11610);
or U12331 (N_12331,N_11800,N_11869);
and U12332 (N_12332,N_11848,N_11986);
nor U12333 (N_12333,N_11723,N_11672);
or U12334 (N_12334,N_11822,N_11836);
and U12335 (N_12335,N_11958,N_11971);
and U12336 (N_12336,N_11692,N_11762);
and U12337 (N_12337,N_11819,N_11973);
and U12338 (N_12338,N_11753,N_11676);
nor U12339 (N_12339,N_11637,N_11815);
nor U12340 (N_12340,N_11673,N_11777);
and U12341 (N_12341,N_11791,N_11851);
nor U12342 (N_12342,N_11666,N_11622);
nor U12343 (N_12343,N_11928,N_11817);
nor U12344 (N_12344,N_11903,N_11610);
nand U12345 (N_12345,N_11631,N_11909);
or U12346 (N_12346,N_11664,N_11898);
or U12347 (N_12347,N_11651,N_11774);
and U12348 (N_12348,N_11928,N_11654);
nor U12349 (N_12349,N_11928,N_11896);
nand U12350 (N_12350,N_11934,N_11657);
nor U12351 (N_12351,N_11947,N_11622);
nand U12352 (N_12352,N_11636,N_11631);
or U12353 (N_12353,N_11897,N_11672);
nor U12354 (N_12354,N_11821,N_11841);
or U12355 (N_12355,N_11711,N_11830);
or U12356 (N_12356,N_11894,N_11878);
nand U12357 (N_12357,N_11827,N_11747);
nor U12358 (N_12358,N_11775,N_11992);
nor U12359 (N_12359,N_11928,N_11756);
and U12360 (N_12360,N_11739,N_11878);
and U12361 (N_12361,N_11862,N_11795);
nor U12362 (N_12362,N_11760,N_11927);
nand U12363 (N_12363,N_11673,N_11836);
or U12364 (N_12364,N_11954,N_11749);
nor U12365 (N_12365,N_11876,N_11658);
nor U12366 (N_12366,N_11612,N_11680);
nand U12367 (N_12367,N_11917,N_11877);
nor U12368 (N_12368,N_11950,N_11990);
nor U12369 (N_12369,N_11950,N_11614);
nor U12370 (N_12370,N_11670,N_11823);
or U12371 (N_12371,N_11887,N_11835);
and U12372 (N_12372,N_11701,N_11724);
nand U12373 (N_12373,N_11859,N_11665);
and U12374 (N_12374,N_11699,N_11698);
and U12375 (N_12375,N_11636,N_11889);
or U12376 (N_12376,N_11757,N_11629);
nor U12377 (N_12377,N_11694,N_11635);
and U12378 (N_12378,N_11685,N_11695);
and U12379 (N_12379,N_11787,N_11844);
nand U12380 (N_12380,N_11676,N_11907);
nand U12381 (N_12381,N_11724,N_11718);
and U12382 (N_12382,N_11810,N_11646);
or U12383 (N_12383,N_11730,N_11744);
nand U12384 (N_12384,N_11822,N_11745);
xor U12385 (N_12385,N_11790,N_11690);
or U12386 (N_12386,N_11914,N_11685);
or U12387 (N_12387,N_11939,N_11989);
and U12388 (N_12388,N_11955,N_11918);
nand U12389 (N_12389,N_11767,N_11729);
nand U12390 (N_12390,N_11818,N_11700);
or U12391 (N_12391,N_11606,N_11835);
nand U12392 (N_12392,N_11837,N_11840);
and U12393 (N_12393,N_11601,N_11671);
and U12394 (N_12394,N_11861,N_11786);
and U12395 (N_12395,N_11702,N_11865);
nand U12396 (N_12396,N_11752,N_11880);
or U12397 (N_12397,N_11995,N_11610);
nand U12398 (N_12398,N_11769,N_11656);
or U12399 (N_12399,N_11914,N_11987);
nor U12400 (N_12400,N_12101,N_12105);
nand U12401 (N_12401,N_12096,N_12288);
and U12402 (N_12402,N_12262,N_12392);
and U12403 (N_12403,N_12373,N_12064);
or U12404 (N_12404,N_12110,N_12348);
nand U12405 (N_12405,N_12084,N_12363);
and U12406 (N_12406,N_12019,N_12005);
nand U12407 (N_12407,N_12237,N_12258);
nor U12408 (N_12408,N_12073,N_12075);
nand U12409 (N_12409,N_12024,N_12012);
nand U12410 (N_12410,N_12203,N_12260);
and U12411 (N_12411,N_12275,N_12234);
or U12412 (N_12412,N_12303,N_12290);
or U12413 (N_12413,N_12062,N_12010);
or U12414 (N_12414,N_12380,N_12383);
or U12415 (N_12415,N_12013,N_12050);
and U12416 (N_12416,N_12365,N_12281);
and U12417 (N_12417,N_12001,N_12305);
or U12418 (N_12418,N_12367,N_12386);
nand U12419 (N_12419,N_12280,N_12081);
nor U12420 (N_12420,N_12014,N_12117);
nand U12421 (N_12421,N_12332,N_12335);
nand U12422 (N_12422,N_12023,N_12201);
nor U12423 (N_12423,N_12277,N_12146);
nand U12424 (N_12424,N_12176,N_12236);
nor U12425 (N_12425,N_12265,N_12178);
or U12426 (N_12426,N_12187,N_12035);
and U12427 (N_12427,N_12209,N_12042);
nand U12428 (N_12428,N_12033,N_12169);
xnor U12429 (N_12429,N_12197,N_12229);
and U12430 (N_12430,N_12111,N_12056);
or U12431 (N_12431,N_12204,N_12104);
nor U12432 (N_12432,N_12051,N_12192);
nor U12433 (N_12433,N_12099,N_12045);
and U12434 (N_12434,N_12221,N_12261);
nor U12435 (N_12435,N_12137,N_12108);
or U12436 (N_12436,N_12271,N_12317);
nand U12437 (N_12437,N_12185,N_12061);
nand U12438 (N_12438,N_12227,N_12021);
xnor U12439 (N_12439,N_12202,N_12313);
nand U12440 (N_12440,N_12315,N_12299);
or U12441 (N_12441,N_12166,N_12055);
nor U12442 (N_12442,N_12341,N_12145);
nand U12443 (N_12443,N_12196,N_12331);
nor U12444 (N_12444,N_12232,N_12256);
or U12445 (N_12445,N_12195,N_12011);
or U12446 (N_12446,N_12279,N_12393);
or U12447 (N_12447,N_12330,N_12162);
nor U12448 (N_12448,N_12250,N_12246);
and U12449 (N_12449,N_12004,N_12038);
nand U12450 (N_12450,N_12396,N_12048);
nand U12451 (N_12451,N_12297,N_12339);
nand U12452 (N_12452,N_12328,N_12337);
nor U12453 (N_12453,N_12200,N_12346);
nor U12454 (N_12454,N_12352,N_12316);
and U12455 (N_12455,N_12116,N_12296);
and U12456 (N_12456,N_12274,N_12268);
or U12457 (N_12457,N_12027,N_12144);
and U12458 (N_12458,N_12127,N_12054);
or U12459 (N_12459,N_12183,N_12003);
or U12460 (N_12460,N_12319,N_12378);
nand U12461 (N_12461,N_12385,N_12077);
and U12462 (N_12462,N_12189,N_12345);
and U12463 (N_12463,N_12002,N_12164);
or U12464 (N_12464,N_12376,N_12006);
nand U12465 (N_12465,N_12366,N_12304);
or U12466 (N_12466,N_12351,N_12031);
nand U12467 (N_12467,N_12368,N_12138);
or U12468 (N_12468,N_12121,N_12302);
nand U12469 (N_12469,N_12134,N_12143);
nor U12470 (N_12470,N_12177,N_12308);
and U12471 (N_12471,N_12210,N_12287);
or U12472 (N_12472,N_12220,N_12282);
or U12473 (N_12473,N_12211,N_12206);
or U12474 (N_12474,N_12284,N_12344);
xor U12475 (N_12475,N_12253,N_12102);
nand U12476 (N_12476,N_12283,N_12039);
or U12477 (N_12477,N_12349,N_12312);
or U12478 (N_12478,N_12047,N_12087);
or U12479 (N_12479,N_12159,N_12394);
nor U12480 (N_12480,N_12184,N_12285);
nor U12481 (N_12481,N_12235,N_12037);
nor U12482 (N_12482,N_12133,N_12388);
nor U12483 (N_12483,N_12090,N_12094);
nand U12484 (N_12484,N_12015,N_12292);
nor U12485 (N_12485,N_12359,N_12286);
and U12486 (N_12486,N_12217,N_12357);
and U12487 (N_12487,N_12018,N_12314);
or U12488 (N_12488,N_12088,N_12186);
or U12489 (N_12489,N_12079,N_12245);
or U12490 (N_12490,N_12172,N_12242);
or U12491 (N_12491,N_12072,N_12318);
nand U12492 (N_12492,N_12028,N_12109);
and U12493 (N_12493,N_12240,N_12374);
and U12494 (N_12494,N_12198,N_12160);
and U12495 (N_12495,N_12149,N_12148);
nor U12496 (N_12496,N_12151,N_12100);
and U12497 (N_12497,N_12324,N_12125);
nor U12498 (N_12498,N_12059,N_12255);
nand U12499 (N_12499,N_12362,N_12112);
and U12500 (N_12500,N_12294,N_12307);
nand U12501 (N_12501,N_12158,N_12239);
nor U12502 (N_12502,N_12171,N_12043);
nor U12503 (N_12503,N_12301,N_12263);
or U12504 (N_12504,N_12129,N_12371);
nor U12505 (N_12505,N_12377,N_12289);
nand U12506 (N_12506,N_12068,N_12040);
or U12507 (N_12507,N_12174,N_12278);
or U12508 (N_12508,N_12218,N_12132);
and U12509 (N_12509,N_12030,N_12325);
and U12510 (N_12510,N_12016,N_12122);
nand U12511 (N_12511,N_12334,N_12182);
or U12512 (N_12512,N_12120,N_12071);
and U12513 (N_12513,N_12060,N_12194);
and U12514 (N_12514,N_12092,N_12049);
and U12515 (N_12515,N_12347,N_12340);
and U12516 (N_12516,N_12252,N_12141);
nor U12517 (N_12517,N_12381,N_12170);
nor U12518 (N_12518,N_12078,N_12089);
and U12519 (N_12519,N_12276,N_12191);
or U12520 (N_12520,N_12085,N_12139);
and U12521 (N_12521,N_12364,N_12032);
or U12522 (N_12522,N_12025,N_12193);
nand U12523 (N_12523,N_12074,N_12390);
nand U12524 (N_12524,N_12399,N_12008);
nand U12525 (N_12525,N_12052,N_12226);
or U12526 (N_12526,N_12215,N_12336);
nor U12527 (N_12527,N_12382,N_12058);
nor U12528 (N_12528,N_12029,N_12343);
and U12529 (N_12529,N_12241,N_12310);
and U12530 (N_12530,N_12333,N_12167);
xnor U12531 (N_12531,N_12208,N_12179);
xor U12532 (N_12532,N_12213,N_12248);
or U12533 (N_12533,N_12273,N_12257);
nand U12534 (N_12534,N_12173,N_12267);
nor U12535 (N_12535,N_12130,N_12152);
nand U12536 (N_12536,N_12247,N_12065);
and U12537 (N_12537,N_12266,N_12395);
nand U12538 (N_12538,N_12327,N_12119);
nor U12539 (N_12539,N_12326,N_12026);
or U12540 (N_12540,N_12036,N_12175);
or U12541 (N_12541,N_12113,N_12387);
nor U12542 (N_12542,N_12207,N_12020);
and U12543 (N_12543,N_12041,N_12205);
nand U12544 (N_12544,N_12291,N_12095);
or U12545 (N_12545,N_12007,N_12228);
and U12546 (N_12546,N_12165,N_12069);
or U12547 (N_12547,N_12034,N_12153);
and U12548 (N_12548,N_12358,N_12369);
nor U12549 (N_12549,N_12398,N_12123);
and U12550 (N_12550,N_12293,N_12259);
and U12551 (N_12551,N_12321,N_12103);
and U12552 (N_12552,N_12370,N_12251);
nor U12553 (N_12553,N_12353,N_12212);
and U12554 (N_12554,N_12180,N_12124);
and U12555 (N_12555,N_12233,N_12156);
xnor U12556 (N_12556,N_12391,N_12136);
nor U12557 (N_12557,N_12131,N_12126);
or U12558 (N_12558,N_12067,N_12379);
nor U12559 (N_12559,N_12243,N_12107);
and U12560 (N_12560,N_12300,N_12115);
nand U12561 (N_12561,N_12161,N_12350);
and U12562 (N_12562,N_12157,N_12118);
and U12563 (N_12563,N_12354,N_12091);
or U12564 (N_12564,N_12222,N_12188);
nand U12565 (N_12565,N_12181,N_12356);
or U12566 (N_12566,N_12295,N_12066);
or U12567 (N_12567,N_12298,N_12070);
or U12568 (N_12568,N_12140,N_12106);
nand U12569 (N_12569,N_12306,N_12168);
nor U12570 (N_12570,N_12231,N_12322);
nand U12571 (N_12571,N_12372,N_12214);
and U12572 (N_12572,N_12223,N_12224);
nand U12573 (N_12573,N_12311,N_12083);
and U12574 (N_12574,N_12086,N_12128);
nand U12575 (N_12575,N_12046,N_12269);
and U12576 (N_12576,N_12142,N_12190);
and U12577 (N_12577,N_12375,N_12320);
nor U12578 (N_12578,N_12397,N_12163);
nor U12579 (N_12579,N_12355,N_12135);
and U12580 (N_12580,N_12053,N_12230);
nand U12581 (N_12581,N_12154,N_12097);
and U12582 (N_12582,N_12323,N_12244);
nor U12583 (N_12583,N_12238,N_12254);
nor U12584 (N_12584,N_12249,N_12093);
nand U12585 (N_12585,N_12360,N_12309);
or U12586 (N_12586,N_12225,N_12000);
and U12587 (N_12587,N_12022,N_12342);
nand U12588 (N_12588,N_12384,N_12270);
nor U12589 (N_12589,N_12009,N_12082);
nor U12590 (N_12590,N_12216,N_12338);
or U12591 (N_12591,N_12155,N_12063);
and U12592 (N_12592,N_12098,N_12199);
nor U12593 (N_12593,N_12017,N_12219);
and U12594 (N_12594,N_12389,N_12329);
xnor U12595 (N_12595,N_12264,N_12150);
and U12596 (N_12596,N_12076,N_12044);
or U12597 (N_12597,N_12114,N_12080);
nor U12598 (N_12598,N_12147,N_12272);
or U12599 (N_12599,N_12361,N_12057);
nor U12600 (N_12600,N_12154,N_12286);
nand U12601 (N_12601,N_12025,N_12393);
or U12602 (N_12602,N_12109,N_12329);
or U12603 (N_12603,N_12343,N_12099);
nand U12604 (N_12604,N_12282,N_12067);
and U12605 (N_12605,N_12218,N_12305);
or U12606 (N_12606,N_12294,N_12170);
or U12607 (N_12607,N_12200,N_12293);
or U12608 (N_12608,N_12068,N_12151);
nor U12609 (N_12609,N_12182,N_12133);
nor U12610 (N_12610,N_12320,N_12219);
nand U12611 (N_12611,N_12087,N_12071);
and U12612 (N_12612,N_12226,N_12170);
nand U12613 (N_12613,N_12185,N_12046);
nor U12614 (N_12614,N_12179,N_12167);
and U12615 (N_12615,N_12107,N_12195);
nor U12616 (N_12616,N_12331,N_12116);
or U12617 (N_12617,N_12394,N_12069);
and U12618 (N_12618,N_12370,N_12387);
or U12619 (N_12619,N_12248,N_12355);
nor U12620 (N_12620,N_12216,N_12227);
nand U12621 (N_12621,N_12305,N_12288);
nor U12622 (N_12622,N_12052,N_12223);
or U12623 (N_12623,N_12024,N_12308);
and U12624 (N_12624,N_12338,N_12326);
nor U12625 (N_12625,N_12271,N_12121);
nor U12626 (N_12626,N_12021,N_12009);
nand U12627 (N_12627,N_12077,N_12051);
or U12628 (N_12628,N_12070,N_12140);
and U12629 (N_12629,N_12167,N_12141);
or U12630 (N_12630,N_12089,N_12364);
or U12631 (N_12631,N_12351,N_12098);
nor U12632 (N_12632,N_12146,N_12123);
or U12633 (N_12633,N_12286,N_12269);
nand U12634 (N_12634,N_12169,N_12006);
nand U12635 (N_12635,N_12360,N_12042);
or U12636 (N_12636,N_12182,N_12205);
nor U12637 (N_12637,N_12144,N_12048);
nand U12638 (N_12638,N_12325,N_12066);
or U12639 (N_12639,N_12258,N_12295);
nor U12640 (N_12640,N_12226,N_12253);
nor U12641 (N_12641,N_12397,N_12185);
and U12642 (N_12642,N_12084,N_12184);
and U12643 (N_12643,N_12173,N_12194);
or U12644 (N_12644,N_12299,N_12147);
and U12645 (N_12645,N_12235,N_12271);
nor U12646 (N_12646,N_12171,N_12190);
nand U12647 (N_12647,N_12008,N_12039);
and U12648 (N_12648,N_12188,N_12046);
or U12649 (N_12649,N_12123,N_12084);
nor U12650 (N_12650,N_12094,N_12379);
nor U12651 (N_12651,N_12178,N_12252);
nor U12652 (N_12652,N_12093,N_12060);
nor U12653 (N_12653,N_12180,N_12278);
or U12654 (N_12654,N_12195,N_12059);
nand U12655 (N_12655,N_12263,N_12207);
or U12656 (N_12656,N_12282,N_12223);
and U12657 (N_12657,N_12338,N_12129);
nor U12658 (N_12658,N_12086,N_12243);
and U12659 (N_12659,N_12033,N_12168);
and U12660 (N_12660,N_12395,N_12396);
or U12661 (N_12661,N_12267,N_12230);
and U12662 (N_12662,N_12019,N_12124);
and U12663 (N_12663,N_12049,N_12207);
or U12664 (N_12664,N_12101,N_12344);
nor U12665 (N_12665,N_12002,N_12273);
nand U12666 (N_12666,N_12257,N_12356);
nand U12667 (N_12667,N_12102,N_12278);
nor U12668 (N_12668,N_12372,N_12307);
nand U12669 (N_12669,N_12215,N_12268);
or U12670 (N_12670,N_12215,N_12131);
and U12671 (N_12671,N_12207,N_12234);
or U12672 (N_12672,N_12172,N_12194);
and U12673 (N_12673,N_12379,N_12152);
or U12674 (N_12674,N_12105,N_12188);
and U12675 (N_12675,N_12207,N_12317);
nand U12676 (N_12676,N_12385,N_12287);
and U12677 (N_12677,N_12274,N_12202);
nand U12678 (N_12678,N_12121,N_12197);
nor U12679 (N_12679,N_12278,N_12285);
nand U12680 (N_12680,N_12166,N_12301);
or U12681 (N_12681,N_12179,N_12291);
nor U12682 (N_12682,N_12319,N_12277);
and U12683 (N_12683,N_12338,N_12078);
nor U12684 (N_12684,N_12068,N_12094);
nor U12685 (N_12685,N_12313,N_12110);
and U12686 (N_12686,N_12061,N_12037);
or U12687 (N_12687,N_12040,N_12324);
nor U12688 (N_12688,N_12195,N_12085);
nor U12689 (N_12689,N_12318,N_12220);
nand U12690 (N_12690,N_12389,N_12050);
or U12691 (N_12691,N_12081,N_12075);
nor U12692 (N_12692,N_12028,N_12114);
or U12693 (N_12693,N_12074,N_12052);
xnor U12694 (N_12694,N_12365,N_12258);
and U12695 (N_12695,N_12275,N_12348);
nor U12696 (N_12696,N_12024,N_12382);
nor U12697 (N_12697,N_12353,N_12092);
nor U12698 (N_12698,N_12014,N_12009);
nand U12699 (N_12699,N_12343,N_12329);
nor U12700 (N_12700,N_12149,N_12229);
nand U12701 (N_12701,N_12002,N_12009);
nand U12702 (N_12702,N_12020,N_12235);
nand U12703 (N_12703,N_12345,N_12332);
nor U12704 (N_12704,N_12290,N_12016);
nor U12705 (N_12705,N_12079,N_12168);
and U12706 (N_12706,N_12041,N_12105);
or U12707 (N_12707,N_12063,N_12079);
and U12708 (N_12708,N_12169,N_12170);
nand U12709 (N_12709,N_12127,N_12040);
nor U12710 (N_12710,N_12270,N_12226);
or U12711 (N_12711,N_12148,N_12122);
nand U12712 (N_12712,N_12301,N_12081);
nor U12713 (N_12713,N_12239,N_12284);
nand U12714 (N_12714,N_12152,N_12192);
or U12715 (N_12715,N_12380,N_12248);
nand U12716 (N_12716,N_12266,N_12247);
nand U12717 (N_12717,N_12118,N_12095);
and U12718 (N_12718,N_12273,N_12114);
or U12719 (N_12719,N_12226,N_12163);
and U12720 (N_12720,N_12184,N_12351);
and U12721 (N_12721,N_12313,N_12174);
nor U12722 (N_12722,N_12069,N_12107);
nand U12723 (N_12723,N_12295,N_12054);
nand U12724 (N_12724,N_12359,N_12077);
or U12725 (N_12725,N_12361,N_12119);
nor U12726 (N_12726,N_12046,N_12094);
nor U12727 (N_12727,N_12353,N_12360);
and U12728 (N_12728,N_12016,N_12114);
and U12729 (N_12729,N_12199,N_12372);
nor U12730 (N_12730,N_12140,N_12329);
nor U12731 (N_12731,N_12196,N_12163);
nand U12732 (N_12732,N_12386,N_12102);
and U12733 (N_12733,N_12027,N_12173);
and U12734 (N_12734,N_12176,N_12367);
and U12735 (N_12735,N_12101,N_12200);
nor U12736 (N_12736,N_12271,N_12139);
nand U12737 (N_12737,N_12030,N_12065);
nor U12738 (N_12738,N_12002,N_12292);
nand U12739 (N_12739,N_12330,N_12267);
nor U12740 (N_12740,N_12157,N_12201);
nor U12741 (N_12741,N_12227,N_12093);
or U12742 (N_12742,N_12262,N_12342);
or U12743 (N_12743,N_12050,N_12087);
nand U12744 (N_12744,N_12313,N_12042);
nor U12745 (N_12745,N_12387,N_12058);
nor U12746 (N_12746,N_12370,N_12388);
and U12747 (N_12747,N_12069,N_12339);
and U12748 (N_12748,N_12178,N_12047);
or U12749 (N_12749,N_12097,N_12245);
and U12750 (N_12750,N_12315,N_12320);
or U12751 (N_12751,N_12298,N_12370);
or U12752 (N_12752,N_12250,N_12370);
or U12753 (N_12753,N_12284,N_12272);
xor U12754 (N_12754,N_12113,N_12085);
nor U12755 (N_12755,N_12291,N_12101);
nor U12756 (N_12756,N_12148,N_12125);
nand U12757 (N_12757,N_12265,N_12135);
nor U12758 (N_12758,N_12334,N_12080);
nor U12759 (N_12759,N_12122,N_12010);
or U12760 (N_12760,N_12014,N_12317);
or U12761 (N_12761,N_12128,N_12277);
nand U12762 (N_12762,N_12090,N_12380);
and U12763 (N_12763,N_12142,N_12311);
nand U12764 (N_12764,N_12265,N_12266);
nor U12765 (N_12765,N_12113,N_12287);
or U12766 (N_12766,N_12201,N_12141);
nor U12767 (N_12767,N_12104,N_12162);
or U12768 (N_12768,N_12226,N_12312);
nor U12769 (N_12769,N_12346,N_12168);
or U12770 (N_12770,N_12183,N_12006);
and U12771 (N_12771,N_12195,N_12361);
or U12772 (N_12772,N_12337,N_12263);
and U12773 (N_12773,N_12342,N_12055);
and U12774 (N_12774,N_12235,N_12273);
or U12775 (N_12775,N_12194,N_12377);
and U12776 (N_12776,N_12360,N_12284);
and U12777 (N_12777,N_12146,N_12360);
nand U12778 (N_12778,N_12227,N_12277);
nor U12779 (N_12779,N_12265,N_12234);
nand U12780 (N_12780,N_12046,N_12189);
nand U12781 (N_12781,N_12255,N_12230);
or U12782 (N_12782,N_12041,N_12310);
nor U12783 (N_12783,N_12381,N_12330);
nand U12784 (N_12784,N_12257,N_12005);
or U12785 (N_12785,N_12022,N_12118);
nor U12786 (N_12786,N_12103,N_12004);
nor U12787 (N_12787,N_12163,N_12023);
or U12788 (N_12788,N_12250,N_12259);
or U12789 (N_12789,N_12265,N_12173);
and U12790 (N_12790,N_12080,N_12199);
nor U12791 (N_12791,N_12236,N_12382);
and U12792 (N_12792,N_12258,N_12214);
nor U12793 (N_12793,N_12084,N_12294);
nor U12794 (N_12794,N_12297,N_12225);
and U12795 (N_12795,N_12030,N_12173);
nor U12796 (N_12796,N_12160,N_12371);
nand U12797 (N_12797,N_12071,N_12190);
nand U12798 (N_12798,N_12350,N_12059);
or U12799 (N_12799,N_12139,N_12388);
or U12800 (N_12800,N_12724,N_12727);
and U12801 (N_12801,N_12471,N_12771);
xnor U12802 (N_12802,N_12472,N_12411);
and U12803 (N_12803,N_12638,N_12692);
nand U12804 (N_12804,N_12442,N_12599);
or U12805 (N_12805,N_12513,N_12779);
and U12806 (N_12806,N_12538,N_12548);
and U12807 (N_12807,N_12636,N_12447);
nor U12808 (N_12808,N_12796,N_12459);
or U12809 (N_12809,N_12432,N_12506);
nand U12810 (N_12810,N_12569,N_12429);
nor U12811 (N_12811,N_12512,N_12700);
and U12812 (N_12812,N_12463,N_12424);
or U12813 (N_12813,N_12642,N_12468);
nand U12814 (N_12814,N_12798,N_12628);
nand U12815 (N_12815,N_12577,N_12756);
and U12816 (N_12816,N_12522,N_12631);
and U12817 (N_12817,N_12458,N_12606);
or U12818 (N_12818,N_12768,N_12466);
nand U12819 (N_12819,N_12658,N_12763);
or U12820 (N_12820,N_12684,N_12477);
nand U12821 (N_12821,N_12561,N_12706);
or U12822 (N_12822,N_12567,N_12774);
and U12823 (N_12823,N_12738,N_12669);
or U12824 (N_12824,N_12467,N_12528);
nand U12825 (N_12825,N_12640,N_12721);
nand U12826 (N_12826,N_12593,N_12720);
or U12827 (N_12827,N_12537,N_12409);
or U12828 (N_12828,N_12649,N_12535);
nand U12829 (N_12829,N_12427,N_12621);
nand U12830 (N_12830,N_12685,N_12697);
nor U12831 (N_12831,N_12540,N_12408);
nand U12832 (N_12832,N_12634,N_12438);
and U12833 (N_12833,N_12602,N_12465);
nor U12834 (N_12834,N_12435,N_12541);
or U12835 (N_12835,N_12770,N_12558);
xor U12836 (N_12836,N_12683,N_12710);
nand U12837 (N_12837,N_12562,N_12469);
nand U12838 (N_12838,N_12603,N_12713);
or U12839 (N_12839,N_12436,N_12783);
or U12840 (N_12840,N_12641,N_12709);
nand U12841 (N_12841,N_12671,N_12677);
nor U12842 (N_12842,N_12550,N_12417);
or U12843 (N_12843,N_12475,N_12648);
or U12844 (N_12844,N_12610,N_12782);
and U12845 (N_12845,N_12691,N_12462);
nor U12846 (N_12846,N_12674,N_12682);
and U12847 (N_12847,N_12410,N_12554);
or U12848 (N_12848,N_12696,N_12553);
nor U12849 (N_12849,N_12443,N_12711);
nor U12850 (N_12850,N_12460,N_12736);
and U12851 (N_12851,N_12620,N_12423);
or U12852 (N_12852,N_12643,N_12769);
or U12853 (N_12853,N_12699,N_12483);
xnor U12854 (N_12854,N_12737,N_12413);
nor U12855 (N_12855,N_12662,N_12492);
nand U12856 (N_12856,N_12747,N_12547);
or U12857 (N_12857,N_12406,N_12639);
and U12858 (N_12858,N_12725,N_12729);
and U12859 (N_12859,N_12637,N_12786);
xor U12860 (N_12860,N_12480,N_12624);
or U12861 (N_12861,N_12470,N_12474);
nor U12862 (N_12862,N_12543,N_12510);
nor U12863 (N_12863,N_12440,N_12404);
and U12864 (N_12864,N_12627,N_12579);
nor U12865 (N_12865,N_12430,N_12485);
nor U12866 (N_12866,N_12461,N_12446);
or U12867 (N_12867,N_12735,N_12743);
and U12868 (N_12868,N_12767,N_12644);
nand U12869 (N_12869,N_12758,N_12766);
or U12870 (N_12870,N_12751,N_12712);
xor U12871 (N_12871,N_12657,N_12740);
or U12872 (N_12872,N_12418,N_12500);
nand U12873 (N_12873,N_12437,N_12784);
or U12874 (N_12874,N_12525,N_12434);
nor U12875 (N_12875,N_12672,N_12645);
or U12876 (N_12876,N_12650,N_12493);
or U12877 (N_12877,N_12777,N_12601);
nor U12878 (N_12878,N_12633,N_12714);
nand U12879 (N_12879,N_12557,N_12791);
and U12880 (N_12880,N_12464,N_12514);
and U12881 (N_12881,N_12688,N_12733);
nor U12882 (N_12882,N_12455,N_12625);
and U12883 (N_12883,N_12750,N_12450);
nor U12884 (N_12884,N_12589,N_12584);
nor U12885 (N_12885,N_12635,N_12539);
nor U12886 (N_12886,N_12509,N_12545);
and U12887 (N_12887,N_12481,N_12582);
nor U12888 (N_12888,N_12753,N_12761);
and U12889 (N_12889,N_12520,N_12705);
and U12890 (N_12890,N_12665,N_12694);
nand U12891 (N_12891,N_12646,N_12679);
or U12892 (N_12892,N_12615,N_12670);
nand U12893 (N_12893,N_12667,N_12619);
and U12894 (N_12894,N_12583,N_12564);
or U12895 (N_12895,N_12505,N_12702);
or U12896 (N_12896,N_12746,N_12789);
or U12897 (N_12897,N_12530,N_12673);
and U12898 (N_12898,N_12715,N_12489);
and U12899 (N_12899,N_12487,N_12590);
nor U12900 (N_12900,N_12653,N_12403);
nand U12901 (N_12901,N_12734,N_12703);
nor U12902 (N_12902,N_12686,N_12723);
and U12903 (N_12903,N_12654,N_12778);
nor U12904 (N_12904,N_12580,N_12776);
nand U12905 (N_12905,N_12659,N_12533);
or U12906 (N_12906,N_12581,N_12596);
and U12907 (N_12907,N_12799,N_12515);
nand U12908 (N_12908,N_12412,N_12503);
or U12909 (N_12909,N_12402,N_12604);
nand U12910 (N_12910,N_12431,N_12749);
or U12911 (N_12911,N_12400,N_12707);
nor U12912 (N_12912,N_12575,N_12422);
nand U12913 (N_12913,N_12594,N_12491);
and U12914 (N_12914,N_12676,N_12698);
or U12915 (N_12915,N_12521,N_12598);
nand U12916 (N_12916,N_12524,N_12797);
or U12917 (N_12917,N_12526,N_12419);
xor U12918 (N_12918,N_12785,N_12661);
nand U12919 (N_12919,N_12586,N_12597);
or U12920 (N_12920,N_12551,N_12792);
nand U12921 (N_12921,N_12563,N_12453);
nand U12922 (N_12922,N_12511,N_12498);
and U12923 (N_12923,N_12484,N_12608);
nor U12924 (N_12924,N_12660,N_12508);
and U12925 (N_12925,N_12687,N_12701);
nor U12926 (N_12926,N_12433,N_12616);
or U12927 (N_12927,N_12428,N_12739);
nand U12928 (N_12928,N_12574,N_12780);
and U12929 (N_12929,N_12401,N_12719);
nand U12930 (N_12930,N_12742,N_12717);
nor U12931 (N_12931,N_12523,N_12656);
nor U12932 (N_12932,N_12448,N_12445);
and U12933 (N_12933,N_12632,N_12416);
and U12934 (N_12934,N_12741,N_12516);
nand U12935 (N_12935,N_12678,N_12745);
nor U12936 (N_12936,N_12405,N_12629);
or U12937 (N_12937,N_12675,N_12668);
nand U12938 (N_12938,N_12421,N_12693);
nand U12939 (N_12939,N_12591,N_12587);
or U12940 (N_12940,N_12726,N_12479);
and U12941 (N_12941,N_12759,N_12454);
or U12942 (N_12942,N_12571,N_12732);
or U12943 (N_12943,N_12555,N_12663);
or U12944 (N_12944,N_12499,N_12614);
or U12945 (N_12945,N_12690,N_12755);
and U12946 (N_12946,N_12731,N_12552);
nand U12947 (N_12947,N_12490,N_12630);
and U12948 (N_12948,N_12572,N_12718);
or U12949 (N_12949,N_12415,N_12452);
and U12950 (N_12950,N_12542,N_12708);
nor U12951 (N_12951,N_12529,N_12494);
nor U12952 (N_12952,N_12781,N_12559);
nand U12953 (N_12953,N_12793,N_12560);
nand U12954 (N_12954,N_12772,N_12451);
and U12955 (N_12955,N_12612,N_12478);
or U12956 (N_12956,N_12689,N_12518);
or U12957 (N_12957,N_12764,N_12600);
and U12958 (N_12958,N_12534,N_12794);
nand U12959 (N_12959,N_12795,N_12546);
nor U12960 (N_12960,N_12651,N_12549);
and U12961 (N_12961,N_12502,N_12544);
nor U12962 (N_12962,N_12444,N_12488);
nand U12963 (N_12963,N_12655,N_12473);
nand U12964 (N_12964,N_12609,N_12449);
nor U12965 (N_12965,N_12425,N_12496);
nor U12966 (N_12966,N_12595,N_12556);
or U12967 (N_12967,N_12607,N_12617);
and U12968 (N_12968,N_12457,N_12748);
nand U12969 (N_12969,N_12578,N_12762);
nand U12970 (N_12970,N_12565,N_12476);
and U12971 (N_12971,N_12618,N_12744);
nor U12972 (N_12972,N_12652,N_12765);
or U12973 (N_12973,N_12622,N_12592);
nor U12974 (N_12974,N_12695,N_12507);
or U12975 (N_12975,N_12588,N_12722);
or U12976 (N_12976,N_12716,N_12788);
nor U12977 (N_12977,N_12754,N_12420);
nand U12978 (N_12978,N_12626,N_12773);
nor U12979 (N_12979,N_12536,N_12482);
nor U12980 (N_12980,N_12752,N_12730);
nand U12981 (N_12981,N_12757,N_12568);
nor U12982 (N_12982,N_12611,N_12497);
nor U12983 (N_12983,N_12407,N_12486);
or U12984 (N_12984,N_12576,N_12704);
nand U12985 (N_12985,N_12728,N_12531);
nor U12986 (N_12986,N_12664,N_12790);
nand U12987 (N_12987,N_12517,N_12441);
and U12988 (N_12988,N_12647,N_12519);
nand U12989 (N_12989,N_12681,N_12570);
and U12990 (N_12990,N_12426,N_12456);
nor U12991 (N_12991,N_12527,N_12573);
or U12992 (N_12992,N_12605,N_12680);
or U12993 (N_12993,N_12566,N_12495);
nand U12994 (N_12994,N_12504,N_12501);
nand U12995 (N_12995,N_12532,N_12775);
nand U12996 (N_12996,N_12666,N_12623);
and U12997 (N_12997,N_12613,N_12760);
and U12998 (N_12998,N_12414,N_12439);
or U12999 (N_12999,N_12787,N_12585);
and U13000 (N_13000,N_12635,N_12771);
or U13001 (N_13001,N_12509,N_12550);
nor U13002 (N_13002,N_12575,N_12782);
and U13003 (N_13003,N_12639,N_12408);
and U13004 (N_13004,N_12532,N_12586);
nand U13005 (N_13005,N_12581,N_12671);
or U13006 (N_13006,N_12788,N_12499);
or U13007 (N_13007,N_12437,N_12601);
or U13008 (N_13008,N_12510,N_12430);
and U13009 (N_13009,N_12463,N_12504);
nor U13010 (N_13010,N_12706,N_12588);
nor U13011 (N_13011,N_12587,N_12623);
or U13012 (N_13012,N_12501,N_12416);
nand U13013 (N_13013,N_12429,N_12441);
and U13014 (N_13014,N_12702,N_12474);
or U13015 (N_13015,N_12674,N_12459);
and U13016 (N_13016,N_12446,N_12567);
nand U13017 (N_13017,N_12697,N_12492);
nand U13018 (N_13018,N_12555,N_12698);
or U13019 (N_13019,N_12440,N_12524);
or U13020 (N_13020,N_12759,N_12575);
or U13021 (N_13021,N_12443,N_12446);
or U13022 (N_13022,N_12482,N_12627);
and U13023 (N_13023,N_12465,N_12768);
and U13024 (N_13024,N_12458,N_12574);
and U13025 (N_13025,N_12589,N_12577);
and U13026 (N_13026,N_12753,N_12525);
nand U13027 (N_13027,N_12472,N_12602);
nand U13028 (N_13028,N_12769,N_12678);
nand U13029 (N_13029,N_12402,N_12758);
and U13030 (N_13030,N_12618,N_12790);
or U13031 (N_13031,N_12792,N_12709);
nand U13032 (N_13032,N_12627,N_12785);
nand U13033 (N_13033,N_12618,N_12619);
nor U13034 (N_13034,N_12554,N_12682);
and U13035 (N_13035,N_12718,N_12793);
nor U13036 (N_13036,N_12757,N_12552);
or U13037 (N_13037,N_12545,N_12489);
nor U13038 (N_13038,N_12649,N_12606);
and U13039 (N_13039,N_12655,N_12589);
or U13040 (N_13040,N_12457,N_12573);
nor U13041 (N_13041,N_12449,N_12657);
nand U13042 (N_13042,N_12403,N_12568);
or U13043 (N_13043,N_12764,N_12449);
and U13044 (N_13044,N_12684,N_12611);
nand U13045 (N_13045,N_12453,N_12489);
or U13046 (N_13046,N_12791,N_12441);
nand U13047 (N_13047,N_12603,N_12683);
and U13048 (N_13048,N_12655,N_12424);
nand U13049 (N_13049,N_12682,N_12751);
nand U13050 (N_13050,N_12524,N_12645);
nor U13051 (N_13051,N_12576,N_12669);
nor U13052 (N_13052,N_12661,N_12663);
nand U13053 (N_13053,N_12434,N_12660);
or U13054 (N_13054,N_12756,N_12786);
or U13055 (N_13055,N_12778,N_12662);
or U13056 (N_13056,N_12732,N_12712);
nand U13057 (N_13057,N_12578,N_12638);
nor U13058 (N_13058,N_12633,N_12469);
or U13059 (N_13059,N_12609,N_12430);
nand U13060 (N_13060,N_12602,N_12542);
and U13061 (N_13061,N_12781,N_12494);
or U13062 (N_13062,N_12655,N_12416);
or U13063 (N_13063,N_12470,N_12417);
and U13064 (N_13064,N_12464,N_12707);
nand U13065 (N_13065,N_12643,N_12458);
nor U13066 (N_13066,N_12768,N_12595);
or U13067 (N_13067,N_12562,N_12692);
xnor U13068 (N_13068,N_12669,N_12425);
nand U13069 (N_13069,N_12510,N_12434);
and U13070 (N_13070,N_12419,N_12700);
nand U13071 (N_13071,N_12643,N_12793);
nand U13072 (N_13072,N_12617,N_12722);
and U13073 (N_13073,N_12739,N_12485);
nand U13074 (N_13074,N_12552,N_12742);
and U13075 (N_13075,N_12705,N_12416);
nand U13076 (N_13076,N_12766,N_12421);
or U13077 (N_13077,N_12407,N_12401);
and U13078 (N_13078,N_12691,N_12741);
or U13079 (N_13079,N_12492,N_12693);
nor U13080 (N_13080,N_12535,N_12722);
and U13081 (N_13081,N_12749,N_12455);
nor U13082 (N_13082,N_12795,N_12516);
and U13083 (N_13083,N_12740,N_12713);
nor U13084 (N_13084,N_12447,N_12797);
or U13085 (N_13085,N_12429,N_12606);
nand U13086 (N_13086,N_12598,N_12483);
nor U13087 (N_13087,N_12475,N_12506);
nor U13088 (N_13088,N_12526,N_12551);
and U13089 (N_13089,N_12660,N_12799);
or U13090 (N_13090,N_12544,N_12693);
or U13091 (N_13091,N_12445,N_12746);
nor U13092 (N_13092,N_12671,N_12633);
or U13093 (N_13093,N_12714,N_12557);
or U13094 (N_13094,N_12706,N_12401);
nor U13095 (N_13095,N_12774,N_12421);
nor U13096 (N_13096,N_12591,N_12738);
nand U13097 (N_13097,N_12556,N_12671);
nand U13098 (N_13098,N_12664,N_12464);
nor U13099 (N_13099,N_12506,N_12676);
and U13100 (N_13100,N_12657,N_12517);
and U13101 (N_13101,N_12442,N_12754);
and U13102 (N_13102,N_12762,N_12442);
xnor U13103 (N_13103,N_12545,N_12543);
and U13104 (N_13104,N_12718,N_12627);
nor U13105 (N_13105,N_12426,N_12792);
nor U13106 (N_13106,N_12620,N_12751);
nor U13107 (N_13107,N_12794,N_12704);
and U13108 (N_13108,N_12416,N_12672);
nand U13109 (N_13109,N_12727,N_12467);
nand U13110 (N_13110,N_12438,N_12580);
nor U13111 (N_13111,N_12715,N_12526);
nor U13112 (N_13112,N_12649,N_12793);
nor U13113 (N_13113,N_12431,N_12476);
or U13114 (N_13114,N_12412,N_12434);
and U13115 (N_13115,N_12584,N_12570);
nand U13116 (N_13116,N_12771,N_12568);
nand U13117 (N_13117,N_12609,N_12583);
xor U13118 (N_13118,N_12418,N_12540);
nor U13119 (N_13119,N_12777,N_12700);
nand U13120 (N_13120,N_12758,N_12697);
nor U13121 (N_13121,N_12559,N_12425);
and U13122 (N_13122,N_12709,N_12666);
nand U13123 (N_13123,N_12549,N_12467);
nand U13124 (N_13124,N_12645,N_12781);
nor U13125 (N_13125,N_12682,N_12695);
and U13126 (N_13126,N_12596,N_12482);
nor U13127 (N_13127,N_12737,N_12414);
or U13128 (N_13128,N_12481,N_12457);
nand U13129 (N_13129,N_12426,N_12728);
and U13130 (N_13130,N_12460,N_12529);
or U13131 (N_13131,N_12759,N_12484);
or U13132 (N_13132,N_12490,N_12475);
and U13133 (N_13133,N_12713,N_12411);
and U13134 (N_13134,N_12441,N_12794);
nor U13135 (N_13135,N_12700,N_12724);
nand U13136 (N_13136,N_12629,N_12684);
or U13137 (N_13137,N_12688,N_12676);
or U13138 (N_13138,N_12439,N_12628);
or U13139 (N_13139,N_12692,N_12781);
or U13140 (N_13140,N_12507,N_12443);
or U13141 (N_13141,N_12609,N_12766);
or U13142 (N_13142,N_12426,N_12580);
nand U13143 (N_13143,N_12743,N_12401);
or U13144 (N_13144,N_12656,N_12608);
nor U13145 (N_13145,N_12563,N_12709);
nor U13146 (N_13146,N_12798,N_12505);
or U13147 (N_13147,N_12416,N_12733);
and U13148 (N_13148,N_12756,N_12775);
nand U13149 (N_13149,N_12680,N_12786);
nor U13150 (N_13150,N_12578,N_12484);
nand U13151 (N_13151,N_12484,N_12453);
nor U13152 (N_13152,N_12606,N_12783);
or U13153 (N_13153,N_12754,N_12668);
nor U13154 (N_13154,N_12712,N_12671);
nor U13155 (N_13155,N_12502,N_12442);
xor U13156 (N_13156,N_12427,N_12436);
nand U13157 (N_13157,N_12589,N_12654);
or U13158 (N_13158,N_12457,N_12561);
and U13159 (N_13159,N_12452,N_12488);
or U13160 (N_13160,N_12476,N_12557);
and U13161 (N_13161,N_12603,N_12531);
xnor U13162 (N_13162,N_12518,N_12515);
nand U13163 (N_13163,N_12466,N_12758);
nor U13164 (N_13164,N_12682,N_12434);
nand U13165 (N_13165,N_12443,N_12478);
and U13166 (N_13166,N_12646,N_12500);
or U13167 (N_13167,N_12754,N_12740);
and U13168 (N_13168,N_12472,N_12475);
nor U13169 (N_13169,N_12417,N_12787);
nor U13170 (N_13170,N_12719,N_12726);
and U13171 (N_13171,N_12585,N_12404);
nor U13172 (N_13172,N_12676,N_12456);
or U13173 (N_13173,N_12794,N_12647);
nand U13174 (N_13174,N_12654,N_12498);
and U13175 (N_13175,N_12720,N_12521);
nand U13176 (N_13176,N_12485,N_12489);
nand U13177 (N_13177,N_12653,N_12609);
or U13178 (N_13178,N_12765,N_12405);
or U13179 (N_13179,N_12692,N_12598);
nor U13180 (N_13180,N_12525,N_12742);
nor U13181 (N_13181,N_12478,N_12403);
or U13182 (N_13182,N_12736,N_12632);
nand U13183 (N_13183,N_12464,N_12564);
nor U13184 (N_13184,N_12608,N_12436);
nand U13185 (N_13185,N_12529,N_12469);
nor U13186 (N_13186,N_12692,N_12430);
and U13187 (N_13187,N_12773,N_12669);
and U13188 (N_13188,N_12670,N_12543);
or U13189 (N_13189,N_12759,N_12571);
and U13190 (N_13190,N_12468,N_12607);
and U13191 (N_13191,N_12781,N_12554);
and U13192 (N_13192,N_12546,N_12700);
or U13193 (N_13193,N_12436,N_12472);
nor U13194 (N_13194,N_12653,N_12749);
and U13195 (N_13195,N_12419,N_12782);
or U13196 (N_13196,N_12538,N_12506);
nand U13197 (N_13197,N_12693,N_12572);
nor U13198 (N_13198,N_12461,N_12701);
nor U13199 (N_13199,N_12609,N_12768);
or U13200 (N_13200,N_12802,N_13168);
nor U13201 (N_13201,N_12833,N_13140);
and U13202 (N_13202,N_13154,N_12904);
and U13203 (N_13203,N_13107,N_13192);
nor U13204 (N_13204,N_13133,N_12821);
or U13205 (N_13205,N_13127,N_13189);
nor U13206 (N_13206,N_12935,N_13056);
nor U13207 (N_13207,N_13052,N_13025);
nor U13208 (N_13208,N_12927,N_12863);
nor U13209 (N_13209,N_13009,N_13100);
nand U13210 (N_13210,N_12999,N_13180);
nor U13211 (N_13211,N_12916,N_12881);
and U13212 (N_13212,N_13182,N_12900);
or U13213 (N_13213,N_12800,N_12929);
or U13214 (N_13214,N_12956,N_12901);
and U13215 (N_13215,N_13124,N_13044);
or U13216 (N_13216,N_12869,N_13010);
and U13217 (N_13217,N_13195,N_13038);
or U13218 (N_13218,N_13125,N_12948);
nor U13219 (N_13219,N_13197,N_13057);
or U13220 (N_13220,N_13033,N_12827);
nor U13221 (N_13221,N_13071,N_13128);
and U13222 (N_13222,N_12878,N_13155);
and U13223 (N_13223,N_12842,N_12921);
or U13224 (N_13224,N_12848,N_12942);
nor U13225 (N_13225,N_13121,N_12940);
or U13226 (N_13226,N_12811,N_12857);
nor U13227 (N_13227,N_12889,N_12925);
and U13228 (N_13228,N_13097,N_12977);
nor U13229 (N_13229,N_12974,N_13015);
nand U13230 (N_13230,N_13074,N_13007);
nand U13231 (N_13231,N_12941,N_12832);
xor U13232 (N_13232,N_13162,N_12895);
nor U13233 (N_13233,N_13031,N_12840);
and U13234 (N_13234,N_13043,N_13148);
or U13235 (N_13235,N_13013,N_12815);
or U13236 (N_13236,N_12947,N_13153);
nand U13237 (N_13237,N_12897,N_12960);
nor U13238 (N_13238,N_13032,N_13085);
and U13239 (N_13239,N_13048,N_13086);
xnor U13240 (N_13240,N_13185,N_13190);
nand U13241 (N_13241,N_13080,N_12908);
and U13242 (N_13242,N_13144,N_12907);
nand U13243 (N_13243,N_12971,N_13171);
and U13244 (N_13244,N_12975,N_13002);
nand U13245 (N_13245,N_12831,N_12870);
nand U13246 (N_13246,N_12843,N_13012);
xnor U13247 (N_13247,N_12893,N_12970);
nand U13248 (N_13248,N_12953,N_13167);
and U13249 (N_13249,N_12814,N_13053);
or U13250 (N_13250,N_13003,N_13017);
nand U13251 (N_13251,N_13020,N_12823);
nor U13252 (N_13252,N_12852,N_12818);
or U13253 (N_13253,N_12939,N_12891);
and U13254 (N_13254,N_12973,N_12911);
nor U13255 (N_13255,N_12986,N_13082);
or U13256 (N_13256,N_12862,N_13123);
nor U13257 (N_13257,N_13076,N_12820);
and U13258 (N_13258,N_12898,N_12928);
nand U13259 (N_13259,N_13161,N_13118);
nor U13260 (N_13260,N_13041,N_13170);
nand U13261 (N_13261,N_13094,N_12903);
or U13262 (N_13262,N_12995,N_13034);
and U13263 (N_13263,N_12855,N_13198);
or U13264 (N_13264,N_13199,N_13112);
nor U13265 (N_13265,N_12932,N_13036);
or U13266 (N_13266,N_13131,N_12980);
or U13267 (N_13267,N_12896,N_12899);
xnor U13268 (N_13268,N_13169,N_13194);
or U13269 (N_13269,N_12844,N_13023);
and U13270 (N_13270,N_13087,N_13152);
nor U13271 (N_13271,N_13050,N_12981);
nor U13272 (N_13272,N_13058,N_12946);
nand U13273 (N_13273,N_13178,N_13011);
or U13274 (N_13274,N_12882,N_13062);
nor U13275 (N_13275,N_13102,N_12860);
nor U13276 (N_13276,N_12867,N_13037);
and U13277 (N_13277,N_13114,N_12957);
nand U13278 (N_13278,N_13141,N_12849);
and U13279 (N_13279,N_12915,N_12991);
nor U13280 (N_13280,N_13084,N_13186);
nand U13281 (N_13281,N_13088,N_12978);
or U13282 (N_13282,N_13181,N_12819);
and U13283 (N_13283,N_12805,N_12822);
or U13284 (N_13284,N_13019,N_12873);
or U13285 (N_13285,N_13177,N_12879);
nor U13286 (N_13286,N_12997,N_13092);
nor U13287 (N_13287,N_13039,N_13024);
nand U13288 (N_13288,N_12983,N_13159);
nor U13289 (N_13289,N_12825,N_12871);
and U13290 (N_13290,N_12979,N_12910);
nand U13291 (N_13291,N_12830,N_12838);
or U13292 (N_13292,N_13175,N_13143);
nand U13293 (N_13293,N_12924,N_13077);
nor U13294 (N_13294,N_12945,N_12874);
nor U13295 (N_13295,N_13089,N_13098);
or U13296 (N_13296,N_13078,N_13113);
xnor U13297 (N_13297,N_13183,N_12807);
nor U13298 (N_13298,N_12865,N_12905);
and U13299 (N_13299,N_13116,N_13008);
nand U13300 (N_13300,N_12868,N_12919);
or U13301 (N_13301,N_12998,N_13069);
nand U13302 (N_13302,N_13018,N_13166);
nor U13303 (N_13303,N_13163,N_13022);
nor U13304 (N_13304,N_12834,N_12959);
xor U13305 (N_13305,N_12824,N_12906);
nor U13306 (N_13306,N_12949,N_12875);
nor U13307 (N_13307,N_13035,N_13176);
nor U13308 (N_13308,N_13054,N_12965);
and U13309 (N_13309,N_13051,N_12828);
and U13310 (N_13310,N_12885,N_12955);
nor U13311 (N_13311,N_12990,N_13106);
or U13312 (N_13312,N_12938,N_13014);
nand U13313 (N_13313,N_13122,N_12839);
and U13314 (N_13314,N_12841,N_13105);
or U13315 (N_13315,N_12853,N_12813);
nor U13316 (N_13316,N_12950,N_12877);
nand U13317 (N_13317,N_13158,N_12951);
or U13318 (N_13318,N_13173,N_13063);
or U13319 (N_13319,N_12926,N_13095);
and U13320 (N_13320,N_12985,N_12968);
and U13321 (N_13321,N_12887,N_12866);
nor U13322 (N_13322,N_12854,N_13179);
and U13323 (N_13323,N_12846,N_13142);
nand U13324 (N_13324,N_12861,N_13047);
nor U13325 (N_13325,N_12984,N_12884);
nand U13326 (N_13326,N_13081,N_13064);
nand U13327 (N_13327,N_12803,N_12993);
nand U13328 (N_13328,N_12851,N_12936);
nand U13329 (N_13329,N_13042,N_12850);
nand U13330 (N_13330,N_12847,N_13110);
or U13331 (N_13331,N_12826,N_13067);
nor U13332 (N_13332,N_12994,N_13165);
and U13333 (N_13333,N_13060,N_12835);
nand U13334 (N_13334,N_12902,N_12934);
or U13335 (N_13335,N_13109,N_13126);
nand U13336 (N_13336,N_13061,N_13196);
nand U13337 (N_13337,N_12914,N_13030);
nor U13338 (N_13338,N_13117,N_12883);
nor U13339 (N_13339,N_13066,N_12817);
and U13340 (N_13340,N_13172,N_12961);
and U13341 (N_13341,N_13111,N_13193);
and U13342 (N_13342,N_12812,N_13104);
or U13343 (N_13343,N_13065,N_13145);
xor U13344 (N_13344,N_12920,N_12806);
or U13345 (N_13345,N_13059,N_13187);
nor U13346 (N_13346,N_13029,N_12845);
nand U13347 (N_13347,N_12969,N_13164);
nor U13348 (N_13348,N_13160,N_12886);
or U13349 (N_13349,N_13108,N_12837);
or U13350 (N_13350,N_12989,N_12864);
nand U13351 (N_13351,N_12808,N_12810);
or U13352 (N_13352,N_12872,N_12963);
or U13353 (N_13353,N_13103,N_12966);
nand U13354 (N_13354,N_12913,N_13115);
or U13355 (N_13355,N_12931,N_12836);
nor U13356 (N_13356,N_13184,N_13157);
and U13357 (N_13357,N_13135,N_12892);
or U13358 (N_13358,N_12890,N_13045);
nor U13359 (N_13359,N_13072,N_13132);
nor U13360 (N_13360,N_12972,N_13049);
or U13361 (N_13361,N_12912,N_13134);
and U13362 (N_13362,N_13146,N_13138);
or U13363 (N_13363,N_13136,N_12888);
or U13364 (N_13364,N_12856,N_12976);
nor U13365 (N_13365,N_12982,N_12952);
and U13366 (N_13366,N_12958,N_13055);
nor U13367 (N_13367,N_13101,N_13090);
nand U13368 (N_13368,N_13005,N_12816);
or U13369 (N_13369,N_12922,N_12964);
nand U13370 (N_13370,N_12933,N_13149);
nor U13371 (N_13371,N_13119,N_12992);
nor U13372 (N_13372,N_13174,N_13073);
nor U13373 (N_13373,N_13001,N_12809);
or U13374 (N_13374,N_13046,N_13150);
and U13375 (N_13375,N_12962,N_12801);
nand U13376 (N_13376,N_12967,N_12917);
or U13377 (N_13377,N_13120,N_12923);
nand U13378 (N_13378,N_12858,N_13188);
or U13379 (N_13379,N_13156,N_13000);
nand U13380 (N_13380,N_13093,N_13083);
nor U13381 (N_13381,N_12937,N_13099);
nand U13382 (N_13382,N_13070,N_13191);
and U13383 (N_13383,N_13068,N_13040);
nor U13384 (N_13384,N_12987,N_12943);
or U13385 (N_13385,N_13139,N_12880);
nand U13386 (N_13386,N_13006,N_12918);
nand U13387 (N_13387,N_13075,N_12829);
nand U13388 (N_13388,N_12876,N_13026);
nor U13389 (N_13389,N_12894,N_12954);
and U13390 (N_13390,N_12996,N_13079);
nand U13391 (N_13391,N_13129,N_12859);
or U13392 (N_13392,N_13137,N_13130);
nand U13393 (N_13393,N_13147,N_13027);
or U13394 (N_13394,N_12804,N_12909);
nand U13395 (N_13395,N_13021,N_13016);
nand U13396 (N_13396,N_13028,N_13091);
and U13397 (N_13397,N_12930,N_13151);
nor U13398 (N_13398,N_12944,N_13096);
or U13399 (N_13399,N_12988,N_13004);
nand U13400 (N_13400,N_12874,N_13121);
or U13401 (N_13401,N_12908,N_13032);
nand U13402 (N_13402,N_12904,N_13046);
or U13403 (N_13403,N_13025,N_13180);
and U13404 (N_13404,N_13024,N_13052);
nand U13405 (N_13405,N_13064,N_12884);
nor U13406 (N_13406,N_13080,N_12954);
nor U13407 (N_13407,N_12808,N_12957);
xor U13408 (N_13408,N_13152,N_12835);
nand U13409 (N_13409,N_12843,N_12961);
and U13410 (N_13410,N_13170,N_13087);
nand U13411 (N_13411,N_13187,N_13077);
or U13412 (N_13412,N_13192,N_12991);
xnor U13413 (N_13413,N_12815,N_13185);
and U13414 (N_13414,N_13047,N_12837);
or U13415 (N_13415,N_13154,N_13082);
nand U13416 (N_13416,N_12950,N_12990);
and U13417 (N_13417,N_13040,N_13148);
and U13418 (N_13418,N_12909,N_13040);
and U13419 (N_13419,N_12979,N_13094);
nor U13420 (N_13420,N_13012,N_12954);
nor U13421 (N_13421,N_12976,N_13017);
nand U13422 (N_13422,N_12921,N_12928);
nor U13423 (N_13423,N_12862,N_12963);
and U13424 (N_13424,N_13135,N_12864);
or U13425 (N_13425,N_12871,N_13015);
or U13426 (N_13426,N_12972,N_13126);
nand U13427 (N_13427,N_13038,N_13199);
and U13428 (N_13428,N_12902,N_12963);
and U13429 (N_13429,N_13190,N_13116);
or U13430 (N_13430,N_12891,N_12802);
and U13431 (N_13431,N_13127,N_12975);
nor U13432 (N_13432,N_12865,N_12806);
nor U13433 (N_13433,N_12864,N_12972);
nor U13434 (N_13434,N_12913,N_13014);
nor U13435 (N_13435,N_12803,N_12900);
nor U13436 (N_13436,N_13118,N_13188);
and U13437 (N_13437,N_12910,N_13115);
and U13438 (N_13438,N_13060,N_12940);
nand U13439 (N_13439,N_12947,N_13068);
nand U13440 (N_13440,N_13015,N_12880);
or U13441 (N_13441,N_13191,N_12923);
or U13442 (N_13442,N_12827,N_12825);
nand U13443 (N_13443,N_12970,N_13102);
or U13444 (N_13444,N_13040,N_12898);
and U13445 (N_13445,N_12870,N_13194);
and U13446 (N_13446,N_12900,N_13130);
and U13447 (N_13447,N_12872,N_13066);
nor U13448 (N_13448,N_13010,N_13071);
nor U13449 (N_13449,N_12930,N_13046);
nor U13450 (N_13450,N_13142,N_13156);
nor U13451 (N_13451,N_12927,N_13085);
nand U13452 (N_13452,N_13070,N_13031);
nand U13453 (N_13453,N_12888,N_12930);
nor U13454 (N_13454,N_12803,N_13005);
nor U13455 (N_13455,N_12893,N_12827);
and U13456 (N_13456,N_12872,N_12976);
or U13457 (N_13457,N_12864,N_13173);
or U13458 (N_13458,N_12849,N_13135);
nand U13459 (N_13459,N_13014,N_13069);
or U13460 (N_13460,N_12950,N_12862);
nor U13461 (N_13461,N_12878,N_13058);
and U13462 (N_13462,N_13077,N_13032);
and U13463 (N_13463,N_13002,N_12992);
and U13464 (N_13464,N_13053,N_12864);
or U13465 (N_13465,N_13018,N_13071);
nand U13466 (N_13466,N_12971,N_12970);
nand U13467 (N_13467,N_12836,N_12972);
or U13468 (N_13468,N_12919,N_13112);
nand U13469 (N_13469,N_13089,N_13159);
or U13470 (N_13470,N_13197,N_12885);
or U13471 (N_13471,N_13069,N_12932);
nor U13472 (N_13472,N_13138,N_13041);
nor U13473 (N_13473,N_13111,N_12898);
and U13474 (N_13474,N_12894,N_13120);
or U13475 (N_13475,N_12997,N_12845);
nor U13476 (N_13476,N_12893,N_13126);
nor U13477 (N_13477,N_12875,N_13055);
nand U13478 (N_13478,N_13155,N_13122);
or U13479 (N_13479,N_12883,N_12929);
or U13480 (N_13480,N_12982,N_12919);
and U13481 (N_13481,N_12953,N_12856);
or U13482 (N_13482,N_12853,N_12857);
and U13483 (N_13483,N_12993,N_12986);
or U13484 (N_13484,N_12917,N_13077);
nor U13485 (N_13485,N_12823,N_12882);
nor U13486 (N_13486,N_13159,N_13061);
nor U13487 (N_13487,N_13180,N_12938);
or U13488 (N_13488,N_12926,N_12915);
nor U13489 (N_13489,N_13112,N_13145);
or U13490 (N_13490,N_12851,N_12862);
nand U13491 (N_13491,N_12903,N_12851);
nor U13492 (N_13492,N_12933,N_13164);
nor U13493 (N_13493,N_13073,N_13057);
nand U13494 (N_13494,N_13057,N_12937);
and U13495 (N_13495,N_13087,N_12850);
or U13496 (N_13496,N_12874,N_12855);
and U13497 (N_13497,N_13092,N_13136);
nand U13498 (N_13498,N_12864,N_13037);
and U13499 (N_13499,N_12926,N_13022);
nand U13500 (N_13500,N_13120,N_13013);
or U13501 (N_13501,N_12804,N_13027);
nor U13502 (N_13502,N_13148,N_13112);
nand U13503 (N_13503,N_12859,N_13190);
or U13504 (N_13504,N_13042,N_12928);
nand U13505 (N_13505,N_13070,N_13039);
nand U13506 (N_13506,N_13091,N_12843);
nor U13507 (N_13507,N_12855,N_13108);
nor U13508 (N_13508,N_13111,N_12815);
or U13509 (N_13509,N_13145,N_13000);
and U13510 (N_13510,N_13057,N_13056);
and U13511 (N_13511,N_12920,N_12808);
nand U13512 (N_13512,N_12912,N_12824);
and U13513 (N_13513,N_13172,N_13014);
and U13514 (N_13514,N_13000,N_13082);
and U13515 (N_13515,N_13152,N_12931);
and U13516 (N_13516,N_12918,N_13168);
nand U13517 (N_13517,N_13181,N_13058);
or U13518 (N_13518,N_12898,N_12839);
nand U13519 (N_13519,N_13114,N_12808);
and U13520 (N_13520,N_12807,N_12932);
or U13521 (N_13521,N_13140,N_13115);
and U13522 (N_13522,N_12989,N_12825);
nor U13523 (N_13523,N_12927,N_13045);
or U13524 (N_13524,N_13037,N_13121);
nor U13525 (N_13525,N_12872,N_12953);
nand U13526 (N_13526,N_13003,N_12997);
nand U13527 (N_13527,N_12865,N_13115);
nand U13528 (N_13528,N_12957,N_12996);
or U13529 (N_13529,N_12855,N_13082);
and U13530 (N_13530,N_12935,N_12847);
nor U13531 (N_13531,N_12821,N_13147);
nand U13532 (N_13532,N_12957,N_12864);
nor U13533 (N_13533,N_13060,N_12974);
nor U13534 (N_13534,N_13070,N_12965);
nand U13535 (N_13535,N_12998,N_12941);
and U13536 (N_13536,N_13102,N_13139);
or U13537 (N_13537,N_13072,N_12862);
or U13538 (N_13538,N_12820,N_13152);
and U13539 (N_13539,N_13143,N_12875);
nor U13540 (N_13540,N_13112,N_12811);
nor U13541 (N_13541,N_12931,N_13173);
nand U13542 (N_13542,N_13031,N_12854);
nand U13543 (N_13543,N_13082,N_12866);
and U13544 (N_13544,N_12852,N_12812);
or U13545 (N_13545,N_12989,N_13016);
nand U13546 (N_13546,N_13033,N_13104);
nor U13547 (N_13547,N_12818,N_13075);
nand U13548 (N_13548,N_12860,N_12963);
or U13549 (N_13549,N_12824,N_12966);
or U13550 (N_13550,N_13118,N_12971);
and U13551 (N_13551,N_12950,N_12860);
and U13552 (N_13552,N_12871,N_12926);
or U13553 (N_13553,N_12880,N_13180);
nand U13554 (N_13554,N_12933,N_13025);
and U13555 (N_13555,N_13061,N_13150);
nand U13556 (N_13556,N_13126,N_13000);
or U13557 (N_13557,N_12842,N_12932);
nor U13558 (N_13558,N_13066,N_13027);
or U13559 (N_13559,N_12891,N_13020);
nand U13560 (N_13560,N_13056,N_12852);
and U13561 (N_13561,N_12870,N_12825);
and U13562 (N_13562,N_12925,N_12917);
nor U13563 (N_13563,N_12974,N_12806);
and U13564 (N_13564,N_12986,N_13136);
or U13565 (N_13565,N_13185,N_13112);
and U13566 (N_13566,N_13193,N_12971);
and U13567 (N_13567,N_12953,N_13194);
or U13568 (N_13568,N_12882,N_12982);
or U13569 (N_13569,N_13155,N_12873);
nor U13570 (N_13570,N_13006,N_12855);
nand U13571 (N_13571,N_12898,N_12860);
or U13572 (N_13572,N_13168,N_13052);
or U13573 (N_13573,N_13140,N_12825);
nor U13574 (N_13574,N_13024,N_13174);
nand U13575 (N_13575,N_13134,N_13189);
or U13576 (N_13576,N_13012,N_12823);
and U13577 (N_13577,N_13190,N_12817);
or U13578 (N_13578,N_12876,N_12836);
nor U13579 (N_13579,N_12885,N_12932);
or U13580 (N_13580,N_12979,N_13109);
and U13581 (N_13581,N_12981,N_13101);
nand U13582 (N_13582,N_12999,N_12907);
and U13583 (N_13583,N_12910,N_12954);
nand U13584 (N_13584,N_12815,N_13125);
nor U13585 (N_13585,N_13021,N_12914);
nor U13586 (N_13586,N_13143,N_12843);
or U13587 (N_13587,N_13158,N_12947);
nor U13588 (N_13588,N_12803,N_12984);
or U13589 (N_13589,N_13119,N_13166);
nor U13590 (N_13590,N_12896,N_13177);
nor U13591 (N_13591,N_13107,N_13188);
and U13592 (N_13592,N_13191,N_13198);
nand U13593 (N_13593,N_13054,N_13061);
nand U13594 (N_13594,N_13044,N_13059);
nor U13595 (N_13595,N_12925,N_12866);
and U13596 (N_13596,N_12989,N_12898);
or U13597 (N_13597,N_12900,N_12980);
nor U13598 (N_13598,N_13083,N_12805);
and U13599 (N_13599,N_13116,N_13004);
or U13600 (N_13600,N_13303,N_13483);
and U13601 (N_13601,N_13586,N_13371);
and U13602 (N_13602,N_13284,N_13367);
or U13603 (N_13603,N_13564,N_13584);
and U13604 (N_13604,N_13309,N_13451);
nand U13605 (N_13605,N_13414,N_13551);
or U13606 (N_13606,N_13337,N_13506);
xor U13607 (N_13607,N_13445,N_13476);
or U13608 (N_13608,N_13539,N_13228);
or U13609 (N_13609,N_13434,N_13323);
or U13610 (N_13610,N_13307,N_13226);
nand U13611 (N_13611,N_13599,N_13413);
nor U13612 (N_13612,N_13428,N_13381);
or U13613 (N_13613,N_13544,N_13457);
nor U13614 (N_13614,N_13396,N_13566);
nand U13615 (N_13615,N_13289,N_13547);
nand U13616 (N_13616,N_13569,N_13562);
and U13617 (N_13617,N_13221,N_13262);
and U13618 (N_13618,N_13285,N_13433);
nor U13619 (N_13619,N_13248,N_13220);
or U13620 (N_13620,N_13342,N_13589);
and U13621 (N_13621,N_13347,N_13438);
nand U13622 (N_13622,N_13505,N_13204);
or U13623 (N_13623,N_13352,N_13200);
nand U13624 (N_13624,N_13391,N_13207);
and U13625 (N_13625,N_13444,N_13540);
nand U13626 (N_13626,N_13295,N_13417);
nand U13627 (N_13627,N_13530,N_13594);
and U13628 (N_13628,N_13430,N_13479);
nand U13629 (N_13629,N_13465,N_13420);
and U13630 (N_13630,N_13443,N_13240);
nor U13631 (N_13631,N_13321,N_13355);
or U13632 (N_13632,N_13514,N_13350);
nor U13633 (N_13633,N_13526,N_13593);
nor U13634 (N_13634,N_13480,N_13233);
nand U13635 (N_13635,N_13344,N_13597);
and U13636 (N_13636,N_13518,N_13249);
nand U13637 (N_13637,N_13432,N_13494);
and U13638 (N_13638,N_13570,N_13275);
and U13639 (N_13639,N_13582,N_13472);
or U13640 (N_13640,N_13409,N_13332);
nor U13641 (N_13641,N_13283,N_13203);
nand U13642 (N_13642,N_13251,N_13500);
nor U13643 (N_13643,N_13508,N_13255);
nand U13644 (N_13644,N_13531,N_13360);
nor U13645 (N_13645,N_13477,N_13528);
or U13646 (N_13646,N_13296,N_13496);
nor U13647 (N_13647,N_13473,N_13462);
or U13648 (N_13648,N_13598,N_13209);
or U13649 (N_13649,N_13202,N_13426);
or U13650 (N_13650,N_13304,N_13591);
nor U13651 (N_13651,N_13592,N_13449);
and U13652 (N_13652,N_13229,N_13583);
nand U13653 (N_13653,N_13448,N_13557);
and U13654 (N_13654,N_13581,N_13537);
and U13655 (N_13655,N_13561,N_13542);
or U13656 (N_13656,N_13231,N_13520);
nor U13657 (N_13657,N_13471,N_13287);
nand U13658 (N_13658,N_13401,N_13468);
nand U13659 (N_13659,N_13305,N_13382);
nand U13660 (N_13660,N_13574,N_13234);
and U13661 (N_13661,N_13595,N_13392);
nand U13662 (N_13662,N_13554,N_13334);
and U13663 (N_13663,N_13458,N_13293);
and U13664 (N_13664,N_13230,N_13560);
nand U13665 (N_13665,N_13298,N_13292);
nand U13666 (N_13666,N_13374,N_13340);
and U13667 (N_13667,N_13276,N_13559);
or U13668 (N_13668,N_13386,N_13365);
nand U13669 (N_13669,N_13288,N_13308);
or U13670 (N_13670,N_13380,N_13330);
nand U13671 (N_13671,N_13400,N_13453);
and U13672 (N_13672,N_13407,N_13241);
nor U13673 (N_13673,N_13403,N_13336);
and U13674 (N_13674,N_13349,N_13546);
nor U13675 (N_13675,N_13238,N_13545);
and U13676 (N_13676,N_13268,N_13259);
or U13677 (N_13677,N_13378,N_13455);
and U13678 (N_13678,N_13524,N_13447);
and U13679 (N_13679,N_13243,N_13213);
and U13680 (N_13680,N_13406,N_13441);
or U13681 (N_13681,N_13568,N_13523);
or U13682 (N_13682,N_13246,N_13541);
nor U13683 (N_13683,N_13356,N_13343);
or U13684 (N_13684,N_13266,N_13532);
or U13685 (N_13685,N_13370,N_13394);
and U13686 (N_13686,N_13281,N_13326);
nand U13687 (N_13687,N_13489,N_13511);
nor U13688 (N_13688,N_13237,N_13482);
nor U13689 (N_13689,N_13300,N_13442);
nand U13690 (N_13690,N_13206,N_13533);
or U13691 (N_13691,N_13317,N_13521);
and U13692 (N_13692,N_13390,N_13236);
nand U13693 (N_13693,N_13527,N_13258);
xor U13694 (N_13694,N_13214,N_13478);
or U13695 (N_13695,N_13205,N_13429);
or U13696 (N_13696,N_13492,N_13577);
nor U13697 (N_13697,N_13516,N_13253);
and U13698 (N_13698,N_13215,N_13579);
nor U13699 (N_13699,N_13211,N_13421);
and U13700 (N_13700,N_13398,N_13498);
nand U13701 (N_13701,N_13459,N_13565);
nand U13702 (N_13702,N_13439,N_13486);
nand U13703 (N_13703,N_13265,N_13452);
or U13704 (N_13704,N_13331,N_13484);
nor U13705 (N_13705,N_13339,N_13558);
or U13706 (N_13706,N_13286,N_13387);
nand U13707 (N_13707,N_13510,N_13252);
nor U13708 (N_13708,N_13219,N_13495);
or U13709 (N_13709,N_13280,N_13201);
nand U13710 (N_13710,N_13454,N_13299);
and U13711 (N_13711,N_13263,N_13502);
nand U13712 (N_13712,N_13416,N_13515);
nand U13713 (N_13713,N_13311,N_13385);
or U13714 (N_13714,N_13315,N_13488);
nor U13715 (N_13715,N_13273,N_13411);
nand U13716 (N_13716,N_13210,N_13440);
and U13717 (N_13717,N_13456,N_13556);
and U13718 (N_13718,N_13519,N_13306);
nor U13719 (N_13719,N_13366,N_13436);
nand U13720 (N_13720,N_13377,N_13320);
nor U13721 (N_13721,N_13277,N_13522);
nor U13722 (N_13722,N_13427,N_13422);
nor U13723 (N_13723,N_13571,N_13379);
or U13724 (N_13724,N_13278,N_13501);
or U13725 (N_13725,N_13250,N_13338);
and U13726 (N_13726,N_13232,N_13239);
and U13727 (N_13727,N_13503,N_13242);
or U13728 (N_13728,N_13590,N_13368);
nand U13729 (N_13729,N_13481,N_13318);
or U13730 (N_13730,N_13322,N_13329);
nor U13731 (N_13731,N_13576,N_13376);
nor U13732 (N_13732,N_13563,N_13314);
or U13733 (N_13733,N_13549,N_13359);
or U13734 (N_13734,N_13464,N_13254);
nor U13735 (N_13735,N_13269,N_13389);
nor U13736 (N_13736,N_13575,N_13474);
nand U13737 (N_13737,N_13497,N_13467);
nor U13738 (N_13738,N_13354,N_13548);
nor U13739 (N_13739,N_13247,N_13450);
nor U13740 (N_13740,N_13372,N_13543);
nor U13741 (N_13741,N_13279,N_13310);
nand U13742 (N_13742,N_13297,N_13225);
or U13743 (N_13743,N_13395,N_13271);
and U13744 (N_13744,N_13325,N_13404);
and U13745 (N_13745,N_13256,N_13312);
and U13746 (N_13746,N_13388,N_13425);
nor U13747 (N_13747,N_13316,N_13357);
nor U13748 (N_13748,N_13529,N_13573);
nand U13749 (N_13749,N_13493,N_13302);
nor U13750 (N_13750,N_13399,N_13517);
and U13751 (N_13751,N_13588,N_13383);
nand U13752 (N_13752,N_13460,N_13536);
and U13753 (N_13753,N_13274,N_13550);
nor U13754 (N_13754,N_13294,N_13423);
and U13755 (N_13755,N_13208,N_13218);
or U13756 (N_13756,N_13487,N_13509);
and U13757 (N_13757,N_13319,N_13410);
or U13758 (N_13758,N_13345,N_13408);
and U13759 (N_13759,N_13555,N_13353);
nand U13760 (N_13760,N_13424,N_13437);
nor U13761 (N_13761,N_13301,N_13333);
nand U13762 (N_13762,N_13270,N_13596);
nor U13763 (N_13763,N_13470,N_13553);
and U13764 (N_13764,N_13405,N_13235);
xnor U13765 (N_13765,N_13290,N_13538);
nand U13766 (N_13766,N_13418,N_13327);
and U13767 (N_13767,N_13580,N_13341);
nor U13768 (N_13768,N_13475,N_13217);
and U13769 (N_13769,N_13504,N_13485);
nor U13770 (N_13770,N_13324,N_13313);
nand U13771 (N_13771,N_13375,N_13412);
nand U13772 (N_13772,N_13261,N_13535);
and U13773 (N_13773,N_13351,N_13373);
nand U13774 (N_13774,N_13578,N_13490);
nand U13775 (N_13775,N_13402,N_13272);
nand U13776 (N_13776,N_13431,N_13267);
nor U13777 (N_13777,N_13348,N_13397);
or U13778 (N_13778,N_13585,N_13525);
and U13779 (N_13779,N_13461,N_13364);
nand U13780 (N_13780,N_13507,N_13245);
nor U13781 (N_13781,N_13534,N_13572);
or U13782 (N_13782,N_13335,N_13328);
nand U13783 (N_13783,N_13216,N_13363);
and U13784 (N_13784,N_13346,N_13257);
and U13785 (N_13785,N_13361,N_13415);
or U13786 (N_13786,N_13291,N_13587);
and U13787 (N_13787,N_13362,N_13469);
and U13788 (N_13788,N_13393,N_13227);
or U13789 (N_13789,N_13463,N_13260);
or U13790 (N_13790,N_13491,N_13212);
nor U13791 (N_13791,N_13223,N_13419);
and U13792 (N_13792,N_13466,N_13567);
nand U13793 (N_13793,N_13512,N_13446);
or U13794 (N_13794,N_13264,N_13369);
or U13795 (N_13795,N_13499,N_13244);
and U13796 (N_13796,N_13222,N_13384);
or U13797 (N_13797,N_13435,N_13513);
or U13798 (N_13798,N_13552,N_13282);
nand U13799 (N_13799,N_13224,N_13358);
or U13800 (N_13800,N_13450,N_13272);
and U13801 (N_13801,N_13445,N_13271);
and U13802 (N_13802,N_13433,N_13453);
nor U13803 (N_13803,N_13582,N_13316);
nand U13804 (N_13804,N_13310,N_13325);
nor U13805 (N_13805,N_13359,N_13277);
or U13806 (N_13806,N_13270,N_13244);
or U13807 (N_13807,N_13522,N_13307);
nand U13808 (N_13808,N_13492,N_13352);
or U13809 (N_13809,N_13431,N_13221);
or U13810 (N_13810,N_13434,N_13300);
and U13811 (N_13811,N_13357,N_13570);
nor U13812 (N_13812,N_13562,N_13383);
or U13813 (N_13813,N_13479,N_13523);
nor U13814 (N_13814,N_13372,N_13567);
and U13815 (N_13815,N_13505,N_13579);
nor U13816 (N_13816,N_13495,N_13331);
nand U13817 (N_13817,N_13492,N_13382);
and U13818 (N_13818,N_13575,N_13424);
nand U13819 (N_13819,N_13370,N_13443);
or U13820 (N_13820,N_13204,N_13217);
nor U13821 (N_13821,N_13419,N_13217);
and U13822 (N_13822,N_13500,N_13448);
and U13823 (N_13823,N_13308,N_13234);
and U13824 (N_13824,N_13398,N_13216);
xnor U13825 (N_13825,N_13489,N_13277);
nor U13826 (N_13826,N_13438,N_13295);
and U13827 (N_13827,N_13217,N_13384);
nand U13828 (N_13828,N_13273,N_13287);
and U13829 (N_13829,N_13515,N_13553);
or U13830 (N_13830,N_13371,N_13200);
or U13831 (N_13831,N_13304,N_13336);
and U13832 (N_13832,N_13244,N_13474);
and U13833 (N_13833,N_13592,N_13575);
nor U13834 (N_13834,N_13404,N_13326);
or U13835 (N_13835,N_13320,N_13267);
nor U13836 (N_13836,N_13323,N_13213);
nand U13837 (N_13837,N_13448,N_13560);
nand U13838 (N_13838,N_13330,N_13493);
nand U13839 (N_13839,N_13426,N_13312);
nor U13840 (N_13840,N_13313,N_13591);
or U13841 (N_13841,N_13413,N_13255);
nand U13842 (N_13842,N_13323,N_13302);
or U13843 (N_13843,N_13585,N_13245);
nor U13844 (N_13844,N_13447,N_13530);
and U13845 (N_13845,N_13281,N_13478);
nand U13846 (N_13846,N_13251,N_13491);
nand U13847 (N_13847,N_13388,N_13572);
nand U13848 (N_13848,N_13215,N_13329);
nor U13849 (N_13849,N_13417,N_13274);
nand U13850 (N_13850,N_13249,N_13396);
nand U13851 (N_13851,N_13374,N_13328);
or U13852 (N_13852,N_13435,N_13250);
and U13853 (N_13853,N_13505,N_13434);
nand U13854 (N_13854,N_13518,N_13423);
nand U13855 (N_13855,N_13581,N_13208);
nand U13856 (N_13856,N_13346,N_13415);
nor U13857 (N_13857,N_13389,N_13350);
nand U13858 (N_13858,N_13409,N_13521);
or U13859 (N_13859,N_13484,N_13207);
or U13860 (N_13860,N_13376,N_13537);
or U13861 (N_13861,N_13562,N_13519);
or U13862 (N_13862,N_13542,N_13206);
nand U13863 (N_13863,N_13374,N_13591);
nand U13864 (N_13864,N_13328,N_13515);
nor U13865 (N_13865,N_13470,N_13531);
nor U13866 (N_13866,N_13364,N_13424);
nor U13867 (N_13867,N_13556,N_13316);
or U13868 (N_13868,N_13297,N_13426);
and U13869 (N_13869,N_13319,N_13315);
nand U13870 (N_13870,N_13465,N_13375);
nor U13871 (N_13871,N_13557,N_13356);
nand U13872 (N_13872,N_13305,N_13394);
and U13873 (N_13873,N_13201,N_13296);
nor U13874 (N_13874,N_13396,N_13454);
nand U13875 (N_13875,N_13439,N_13582);
nor U13876 (N_13876,N_13509,N_13417);
and U13877 (N_13877,N_13488,N_13245);
or U13878 (N_13878,N_13369,N_13301);
nand U13879 (N_13879,N_13311,N_13438);
and U13880 (N_13880,N_13310,N_13566);
nor U13881 (N_13881,N_13444,N_13452);
nor U13882 (N_13882,N_13536,N_13511);
and U13883 (N_13883,N_13460,N_13324);
nor U13884 (N_13884,N_13207,N_13252);
nand U13885 (N_13885,N_13342,N_13521);
and U13886 (N_13886,N_13360,N_13596);
or U13887 (N_13887,N_13409,N_13353);
nor U13888 (N_13888,N_13598,N_13272);
and U13889 (N_13889,N_13446,N_13450);
or U13890 (N_13890,N_13302,N_13318);
or U13891 (N_13891,N_13258,N_13296);
or U13892 (N_13892,N_13348,N_13491);
nor U13893 (N_13893,N_13547,N_13539);
nor U13894 (N_13894,N_13487,N_13303);
and U13895 (N_13895,N_13285,N_13490);
nor U13896 (N_13896,N_13506,N_13283);
nor U13897 (N_13897,N_13330,N_13458);
nor U13898 (N_13898,N_13314,N_13420);
nand U13899 (N_13899,N_13428,N_13296);
or U13900 (N_13900,N_13450,N_13492);
nand U13901 (N_13901,N_13565,N_13448);
and U13902 (N_13902,N_13485,N_13399);
or U13903 (N_13903,N_13580,N_13465);
nor U13904 (N_13904,N_13484,N_13295);
and U13905 (N_13905,N_13590,N_13572);
nand U13906 (N_13906,N_13550,N_13302);
or U13907 (N_13907,N_13509,N_13395);
or U13908 (N_13908,N_13252,N_13592);
nand U13909 (N_13909,N_13291,N_13403);
nand U13910 (N_13910,N_13474,N_13583);
nand U13911 (N_13911,N_13463,N_13591);
nor U13912 (N_13912,N_13324,N_13283);
nor U13913 (N_13913,N_13329,N_13262);
nand U13914 (N_13914,N_13397,N_13376);
nor U13915 (N_13915,N_13275,N_13374);
or U13916 (N_13916,N_13593,N_13278);
nand U13917 (N_13917,N_13335,N_13200);
nor U13918 (N_13918,N_13205,N_13318);
and U13919 (N_13919,N_13343,N_13391);
nor U13920 (N_13920,N_13388,N_13550);
or U13921 (N_13921,N_13298,N_13200);
nand U13922 (N_13922,N_13553,N_13471);
and U13923 (N_13923,N_13450,N_13383);
nor U13924 (N_13924,N_13285,N_13477);
or U13925 (N_13925,N_13307,N_13476);
and U13926 (N_13926,N_13589,N_13430);
nor U13927 (N_13927,N_13371,N_13273);
nor U13928 (N_13928,N_13497,N_13548);
or U13929 (N_13929,N_13594,N_13269);
nand U13930 (N_13930,N_13304,N_13438);
nand U13931 (N_13931,N_13399,N_13477);
or U13932 (N_13932,N_13217,N_13452);
nand U13933 (N_13933,N_13263,N_13374);
and U13934 (N_13934,N_13289,N_13561);
nand U13935 (N_13935,N_13232,N_13212);
nor U13936 (N_13936,N_13336,N_13227);
or U13937 (N_13937,N_13401,N_13558);
or U13938 (N_13938,N_13208,N_13565);
nor U13939 (N_13939,N_13477,N_13372);
and U13940 (N_13940,N_13528,N_13380);
or U13941 (N_13941,N_13352,N_13528);
nand U13942 (N_13942,N_13466,N_13518);
or U13943 (N_13943,N_13549,N_13576);
and U13944 (N_13944,N_13416,N_13596);
nand U13945 (N_13945,N_13335,N_13558);
nand U13946 (N_13946,N_13306,N_13415);
nand U13947 (N_13947,N_13305,N_13461);
and U13948 (N_13948,N_13529,N_13592);
or U13949 (N_13949,N_13370,N_13467);
nand U13950 (N_13950,N_13421,N_13273);
and U13951 (N_13951,N_13497,N_13314);
nand U13952 (N_13952,N_13253,N_13223);
nor U13953 (N_13953,N_13514,N_13562);
and U13954 (N_13954,N_13571,N_13400);
or U13955 (N_13955,N_13232,N_13236);
and U13956 (N_13956,N_13470,N_13494);
and U13957 (N_13957,N_13384,N_13363);
nand U13958 (N_13958,N_13391,N_13321);
nor U13959 (N_13959,N_13386,N_13401);
nand U13960 (N_13960,N_13387,N_13270);
nand U13961 (N_13961,N_13237,N_13563);
and U13962 (N_13962,N_13518,N_13384);
or U13963 (N_13963,N_13447,N_13533);
and U13964 (N_13964,N_13236,N_13330);
nor U13965 (N_13965,N_13452,N_13398);
and U13966 (N_13966,N_13235,N_13545);
nand U13967 (N_13967,N_13430,N_13284);
nand U13968 (N_13968,N_13375,N_13431);
nand U13969 (N_13969,N_13359,N_13367);
or U13970 (N_13970,N_13236,N_13551);
nand U13971 (N_13971,N_13305,N_13584);
or U13972 (N_13972,N_13479,N_13335);
nor U13973 (N_13973,N_13202,N_13384);
nor U13974 (N_13974,N_13313,N_13416);
nor U13975 (N_13975,N_13268,N_13452);
and U13976 (N_13976,N_13450,N_13580);
nor U13977 (N_13977,N_13265,N_13555);
nand U13978 (N_13978,N_13596,N_13586);
nand U13979 (N_13979,N_13587,N_13271);
nand U13980 (N_13980,N_13532,N_13290);
nor U13981 (N_13981,N_13506,N_13550);
nor U13982 (N_13982,N_13460,N_13296);
or U13983 (N_13983,N_13403,N_13476);
and U13984 (N_13984,N_13580,N_13265);
nor U13985 (N_13985,N_13571,N_13567);
or U13986 (N_13986,N_13406,N_13463);
xnor U13987 (N_13987,N_13379,N_13474);
nand U13988 (N_13988,N_13486,N_13476);
and U13989 (N_13989,N_13236,N_13428);
nor U13990 (N_13990,N_13480,N_13372);
nand U13991 (N_13991,N_13211,N_13497);
or U13992 (N_13992,N_13442,N_13359);
nor U13993 (N_13993,N_13367,N_13507);
and U13994 (N_13994,N_13298,N_13278);
or U13995 (N_13995,N_13213,N_13568);
and U13996 (N_13996,N_13449,N_13360);
nor U13997 (N_13997,N_13326,N_13519);
nor U13998 (N_13998,N_13239,N_13593);
or U13999 (N_13999,N_13276,N_13446);
nor U14000 (N_14000,N_13643,N_13631);
nand U14001 (N_14001,N_13966,N_13805);
nor U14002 (N_14002,N_13611,N_13777);
and U14003 (N_14003,N_13645,N_13670);
or U14004 (N_14004,N_13740,N_13957);
nand U14005 (N_14005,N_13801,N_13739);
nand U14006 (N_14006,N_13871,N_13616);
nor U14007 (N_14007,N_13936,N_13843);
or U14008 (N_14008,N_13730,N_13771);
or U14009 (N_14009,N_13747,N_13889);
xnor U14010 (N_14010,N_13917,N_13899);
and U14011 (N_14011,N_13911,N_13931);
nand U14012 (N_14012,N_13683,N_13703);
nand U14013 (N_14013,N_13835,N_13902);
nand U14014 (N_14014,N_13685,N_13792);
and U14015 (N_14015,N_13733,N_13692);
or U14016 (N_14016,N_13811,N_13967);
and U14017 (N_14017,N_13992,N_13769);
or U14018 (N_14018,N_13656,N_13767);
nor U14019 (N_14019,N_13676,N_13925);
nand U14020 (N_14020,N_13999,N_13738);
nor U14021 (N_14021,N_13726,N_13824);
nand U14022 (N_14022,N_13695,N_13655);
nand U14023 (N_14023,N_13648,N_13834);
nand U14024 (N_14024,N_13632,N_13618);
nand U14025 (N_14025,N_13723,N_13875);
nor U14026 (N_14026,N_13704,N_13634);
nor U14027 (N_14027,N_13937,N_13849);
and U14028 (N_14028,N_13839,N_13660);
and U14029 (N_14029,N_13946,N_13831);
and U14030 (N_14030,N_13793,N_13714);
or U14031 (N_14031,N_13995,N_13786);
nor U14032 (N_14032,N_13880,N_13705);
or U14033 (N_14033,N_13844,N_13797);
or U14034 (N_14034,N_13859,N_13753);
nor U14035 (N_14035,N_13898,N_13668);
nand U14036 (N_14036,N_13894,N_13809);
or U14037 (N_14037,N_13850,N_13601);
or U14038 (N_14038,N_13744,N_13633);
nand U14039 (N_14039,N_13900,N_13972);
and U14040 (N_14040,N_13680,N_13641);
and U14041 (N_14041,N_13851,N_13847);
or U14042 (N_14042,N_13840,N_13830);
and U14043 (N_14043,N_13855,N_13816);
and U14044 (N_14044,N_13798,N_13841);
and U14045 (N_14045,N_13788,N_13861);
and U14046 (N_14046,N_13803,N_13615);
and U14047 (N_14047,N_13672,N_13884);
or U14048 (N_14048,N_13944,N_13838);
nor U14049 (N_14049,N_13605,N_13940);
nand U14050 (N_14050,N_13784,N_13970);
nand U14051 (N_14051,N_13993,N_13761);
nand U14052 (N_14052,N_13954,N_13895);
nand U14053 (N_14053,N_13709,N_13909);
or U14054 (N_14054,N_13780,N_13918);
nand U14055 (N_14055,N_13958,N_13657);
or U14056 (N_14056,N_13883,N_13653);
nand U14057 (N_14057,N_13845,N_13650);
and U14058 (N_14058,N_13912,N_13825);
nand U14059 (N_14059,N_13983,N_13949);
nor U14060 (N_14060,N_13699,N_13906);
and U14061 (N_14061,N_13916,N_13901);
nand U14062 (N_14062,N_13987,N_13613);
or U14063 (N_14063,N_13752,N_13913);
or U14064 (N_14064,N_13642,N_13904);
nand U14065 (N_14065,N_13727,N_13969);
and U14066 (N_14066,N_13819,N_13971);
nand U14067 (N_14067,N_13757,N_13735);
nand U14068 (N_14068,N_13823,N_13896);
nand U14069 (N_14069,N_13742,N_13951);
nor U14070 (N_14070,N_13688,N_13998);
nor U14071 (N_14071,N_13905,N_13796);
and U14072 (N_14072,N_13930,N_13827);
nor U14073 (N_14073,N_13789,N_13927);
and U14074 (N_14074,N_13887,N_13921);
nor U14075 (N_14075,N_13626,N_13684);
nor U14076 (N_14076,N_13713,N_13669);
and U14077 (N_14077,N_13867,N_13890);
nor U14078 (N_14078,N_13678,N_13873);
nand U14079 (N_14079,N_13860,N_13857);
nor U14080 (N_14080,N_13609,N_13746);
nand U14081 (N_14081,N_13817,N_13624);
nand U14082 (N_14082,N_13700,N_13636);
and U14083 (N_14083,N_13920,N_13745);
nand U14084 (N_14084,N_13782,N_13960);
nor U14085 (N_14085,N_13988,N_13625);
nand U14086 (N_14086,N_13863,N_13986);
or U14087 (N_14087,N_13687,N_13852);
or U14088 (N_14088,N_13622,N_13929);
or U14089 (N_14089,N_13897,N_13996);
and U14090 (N_14090,N_13846,N_13608);
or U14091 (N_14091,N_13759,N_13985);
or U14092 (N_14092,N_13702,N_13720);
nor U14093 (N_14093,N_13962,N_13778);
and U14094 (N_14094,N_13952,N_13749);
nand U14095 (N_14095,N_13681,N_13978);
nand U14096 (N_14096,N_13935,N_13724);
or U14097 (N_14097,N_13603,N_13812);
nand U14098 (N_14098,N_13964,N_13828);
nand U14099 (N_14099,N_13984,N_13800);
nor U14100 (N_14100,N_13785,N_13600);
and U14101 (N_14101,N_13674,N_13804);
nand U14102 (N_14102,N_13950,N_13829);
nor U14103 (N_14103,N_13820,N_13891);
xnor U14104 (N_14104,N_13821,N_13639);
nand U14105 (N_14105,N_13725,N_13955);
nor U14106 (N_14106,N_13664,N_13832);
or U14107 (N_14107,N_13651,N_13776);
or U14108 (N_14108,N_13652,N_13886);
nand U14109 (N_14109,N_13647,N_13719);
or U14110 (N_14110,N_13848,N_13864);
and U14111 (N_14111,N_13619,N_13662);
or U14112 (N_14112,N_13976,N_13926);
nor U14113 (N_14113,N_13961,N_13721);
or U14114 (N_14114,N_13799,N_13659);
or U14115 (N_14115,N_13773,N_13748);
and U14116 (N_14116,N_13826,N_13696);
nor U14117 (N_14117,N_13856,N_13602);
nand U14118 (N_14118,N_13706,N_13649);
nand U14119 (N_14119,N_13693,N_13661);
nor U14120 (N_14120,N_13965,N_13722);
or U14121 (N_14121,N_13667,N_13712);
nor U14122 (N_14122,N_13663,N_13837);
nand U14123 (N_14123,N_13677,N_13945);
nand U14124 (N_14124,N_13754,N_13914);
or U14125 (N_14125,N_13710,N_13932);
and U14126 (N_14126,N_13948,N_13666);
nor U14127 (N_14127,N_13617,N_13635);
nor U14128 (N_14128,N_13818,N_13628);
or U14129 (N_14129,N_13963,N_13637);
and U14130 (N_14130,N_13795,N_13853);
nor U14131 (N_14131,N_13729,N_13878);
or U14132 (N_14132,N_13689,N_13833);
nor U14133 (N_14133,N_13755,N_13708);
nand U14134 (N_14134,N_13968,N_13815);
nor U14135 (N_14135,N_13989,N_13694);
nor U14136 (N_14136,N_13981,N_13743);
or U14137 (N_14137,N_13974,N_13881);
nor U14138 (N_14138,N_13934,N_13893);
and U14139 (N_14139,N_13686,N_13922);
and U14140 (N_14140,N_13953,N_13865);
and U14141 (N_14141,N_13903,N_13770);
or U14142 (N_14142,N_13716,N_13715);
or U14143 (N_14143,N_13774,N_13604);
and U14144 (N_14144,N_13933,N_13858);
or U14145 (N_14145,N_13790,N_13763);
and U14146 (N_14146,N_13679,N_13766);
or U14147 (N_14147,N_13781,N_13607);
and U14148 (N_14148,N_13783,N_13938);
nor U14149 (N_14149,N_13764,N_13736);
nand U14150 (N_14150,N_13959,N_13814);
or U14151 (N_14151,N_13640,N_13658);
nor U14152 (N_14152,N_13813,N_13928);
or U14153 (N_14153,N_13673,N_13697);
nand U14154 (N_14154,N_13870,N_13731);
and U14155 (N_14155,N_13924,N_13734);
or U14156 (N_14156,N_13977,N_13760);
nand U14157 (N_14157,N_13810,N_13997);
nor U14158 (N_14158,N_13779,N_13939);
nor U14159 (N_14159,N_13876,N_13758);
nand U14160 (N_14160,N_13888,N_13943);
or U14161 (N_14161,N_13947,N_13629);
nand U14162 (N_14162,N_13610,N_13623);
and U14163 (N_14163,N_13872,N_13718);
nor U14164 (N_14164,N_13606,N_13630);
or U14165 (N_14165,N_13942,N_13806);
and U14166 (N_14166,N_13750,N_13711);
and U14167 (N_14167,N_13941,N_13682);
nor U14168 (N_14168,N_13802,N_13980);
nor U14169 (N_14169,N_13866,N_13741);
or U14170 (N_14170,N_13638,N_13762);
nor U14171 (N_14171,N_13885,N_13791);
and U14172 (N_14172,N_13807,N_13671);
or U14173 (N_14173,N_13775,N_13701);
nor U14174 (N_14174,N_13908,N_13654);
nor U14175 (N_14175,N_13874,N_13994);
nand U14176 (N_14176,N_13836,N_13627);
and U14177 (N_14177,N_13691,N_13665);
or U14178 (N_14178,N_13862,N_13620);
and U14179 (N_14179,N_13772,N_13717);
or U14180 (N_14180,N_13910,N_13892);
nor U14181 (N_14181,N_13614,N_13868);
nor U14182 (N_14182,N_13822,N_13675);
or U14183 (N_14183,N_13756,N_13973);
and U14184 (N_14184,N_13765,N_13923);
or U14185 (N_14185,N_13991,N_13907);
or U14186 (N_14186,N_13915,N_13982);
nor U14187 (N_14187,N_13794,N_13737);
nand U14188 (N_14188,N_13707,N_13751);
or U14189 (N_14189,N_13787,N_13869);
nand U14190 (N_14190,N_13732,N_13990);
nor U14191 (N_14191,N_13854,N_13975);
or U14192 (N_14192,N_13879,N_13808);
and U14193 (N_14193,N_13877,N_13842);
nor U14194 (N_14194,N_13612,N_13768);
and U14195 (N_14195,N_13698,N_13646);
or U14196 (N_14196,N_13882,N_13956);
or U14197 (N_14197,N_13728,N_13690);
or U14198 (N_14198,N_13919,N_13644);
and U14199 (N_14199,N_13979,N_13621);
or U14200 (N_14200,N_13766,N_13616);
or U14201 (N_14201,N_13974,N_13877);
xnor U14202 (N_14202,N_13826,N_13879);
and U14203 (N_14203,N_13976,N_13686);
and U14204 (N_14204,N_13659,N_13682);
and U14205 (N_14205,N_13616,N_13944);
and U14206 (N_14206,N_13624,N_13884);
nor U14207 (N_14207,N_13827,N_13730);
nand U14208 (N_14208,N_13737,N_13810);
nand U14209 (N_14209,N_13657,N_13734);
nor U14210 (N_14210,N_13882,N_13691);
or U14211 (N_14211,N_13820,N_13842);
nor U14212 (N_14212,N_13956,N_13659);
nor U14213 (N_14213,N_13761,N_13738);
nor U14214 (N_14214,N_13933,N_13725);
xor U14215 (N_14215,N_13706,N_13780);
nor U14216 (N_14216,N_13872,N_13719);
nand U14217 (N_14217,N_13701,N_13746);
nor U14218 (N_14218,N_13901,N_13927);
nand U14219 (N_14219,N_13670,N_13879);
and U14220 (N_14220,N_13958,N_13736);
or U14221 (N_14221,N_13701,N_13781);
and U14222 (N_14222,N_13642,N_13835);
nor U14223 (N_14223,N_13760,N_13998);
or U14224 (N_14224,N_13778,N_13805);
nor U14225 (N_14225,N_13618,N_13893);
nand U14226 (N_14226,N_13882,N_13904);
nand U14227 (N_14227,N_13906,N_13611);
nor U14228 (N_14228,N_13952,N_13785);
nor U14229 (N_14229,N_13630,N_13692);
nand U14230 (N_14230,N_13645,N_13965);
or U14231 (N_14231,N_13889,N_13773);
or U14232 (N_14232,N_13811,N_13946);
nand U14233 (N_14233,N_13953,N_13601);
or U14234 (N_14234,N_13897,N_13637);
or U14235 (N_14235,N_13901,N_13799);
nor U14236 (N_14236,N_13987,N_13656);
xnor U14237 (N_14237,N_13835,N_13761);
nand U14238 (N_14238,N_13780,N_13866);
nand U14239 (N_14239,N_13930,N_13934);
and U14240 (N_14240,N_13624,N_13770);
or U14241 (N_14241,N_13855,N_13651);
nor U14242 (N_14242,N_13712,N_13833);
nand U14243 (N_14243,N_13811,N_13876);
or U14244 (N_14244,N_13831,N_13659);
nand U14245 (N_14245,N_13661,N_13678);
nor U14246 (N_14246,N_13869,N_13725);
and U14247 (N_14247,N_13991,N_13757);
or U14248 (N_14248,N_13634,N_13652);
nand U14249 (N_14249,N_13947,N_13608);
and U14250 (N_14250,N_13710,N_13897);
nand U14251 (N_14251,N_13633,N_13785);
nand U14252 (N_14252,N_13659,N_13668);
nand U14253 (N_14253,N_13751,N_13692);
and U14254 (N_14254,N_13657,N_13676);
and U14255 (N_14255,N_13642,N_13920);
and U14256 (N_14256,N_13802,N_13855);
nor U14257 (N_14257,N_13670,N_13849);
and U14258 (N_14258,N_13671,N_13955);
nand U14259 (N_14259,N_13814,N_13850);
nand U14260 (N_14260,N_13757,N_13954);
nor U14261 (N_14261,N_13790,N_13833);
nor U14262 (N_14262,N_13910,N_13972);
nand U14263 (N_14263,N_13896,N_13830);
nand U14264 (N_14264,N_13949,N_13740);
xor U14265 (N_14265,N_13902,N_13855);
or U14266 (N_14266,N_13924,N_13631);
nand U14267 (N_14267,N_13974,N_13958);
nand U14268 (N_14268,N_13869,N_13777);
and U14269 (N_14269,N_13617,N_13784);
and U14270 (N_14270,N_13612,N_13688);
nor U14271 (N_14271,N_13777,N_13975);
nand U14272 (N_14272,N_13627,N_13647);
nand U14273 (N_14273,N_13687,N_13667);
nor U14274 (N_14274,N_13728,N_13619);
nand U14275 (N_14275,N_13944,N_13621);
nor U14276 (N_14276,N_13743,N_13856);
nand U14277 (N_14277,N_13978,N_13925);
nand U14278 (N_14278,N_13760,N_13861);
nor U14279 (N_14279,N_13987,N_13971);
and U14280 (N_14280,N_13976,N_13787);
nor U14281 (N_14281,N_13623,N_13642);
nand U14282 (N_14282,N_13810,N_13697);
xor U14283 (N_14283,N_13777,N_13972);
nand U14284 (N_14284,N_13848,N_13922);
or U14285 (N_14285,N_13777,N_13985);
or U14286 (N_14286,N_13915,N_13953);
and U14287 (N_14287,N_13844,N_13846);
or U14288 (N_14288,N_13771,N_13742);
nor U14289 (N_14289,N_13998,N_13924);
or U14290 (N_14290,N_13820,N_13847);
nor U14291 (N_14291,N_13954,N_13824);
or U14292 (N_14292,N_13995,N_13627);
or U14293 (N_14293,N_13810,N_13688);
nand U14294 (N_14294,N_13907,N_13915);
or U14295 (N_14295,N_13849,N_13666);
or U14296 (N_14296,N_13863,N_13825);
nor U14297 (N_14297,N_13938,N_13932);
nor U14298 (N_14298,N_13993,N_13870);
nand U14299 (N_14299,N_13657,N_13710);
and U14300 (N_14300,N_13699,N_13998);
nor U14301 (N_14301,N_13938,N_13770);
or U14302 (N_14302,N_13706,N_13776);
nand U14303 (N_14303,N_13620,N_13984);
nand U14304 (N_14304,N_13612,N_13982);
nand U14305 (N_14305,N_13720,N_13766);
and U14306 (N_14306,N_13816,N_13868);
or U14307 (N_14307,N_13738,N_13863);
and U14308 (N_14308,N_13895,N_13769);
or U14309 (N_14309,N_13731,N_13847);
or U14310 (N_14310,N_13920,N_13609);
nand U14311 (N_14311,N_13639,N_13832);
nand U14312 (N_14312,N_13929,N_13698);
nor U14313 (N_14313,N_13823,N_13793);
and U14314 (N_14314,N_13736,N_13711);
or U14315 (N_14315,N_13751,N_13720);
nor U14316 (N_14316,N_13989,N_13997);
nand U14317 (N_14317,N_13909,N_13668);
or U14318 (N_14318,N_13681,N_13893);
nor U14319 (N_14319,N_13884,N_13853);
and U14320 (N_14320,N_13799,N_13847);
nand U14321 (N_14321,N_13660,N_13755);
and U14322 (N_14322,N_13892,N_13737);
nor U14323 (N_14323,N_13742,N_13840);
or U14324 (N_14324,N_13932,N_13796);
or U14325 (N_14325,N_13811,N_13740);
or U14326 (N_14326,N_13928,N_13951);
nand U14327 (N_14327,N_13960,N_13815);
nor U14328 (N_14328,N_13603,N_13665);
or U14329 (N_14329,N_13600,N_13633);
nand U14330 (N_14330,N_13957,N_13937);
nand U14331 (N_14331,N_13737,N_13727);
or U14332 (N_14332,N_13885,N_13631);
nor U14333 (N_14333,N_13757,N_13825);
and U14334 (N_14334,N_13793,N_13741);
nand U14335 (N_14335,N_13747,N_13855);
nor U14336 (N_14336,N_13940,N_13704);
nor U14337 (N_14337,N_13897,N_13924);
nand U14338 (N_14338,N_13822,N_13859);
nand U14339 (N_14339,N_13603,N_13821);
or U14340 (N_14340,N_13913,N_13903);
nand U14341 (N_14341,N_13876,N_13879);
nor U14342 (N_14342,N_13669,N_13797);
and U14343 (N_14343,N_13873,N_13893);
and U14344 (N_14344,N_13610,N_13684);
or U14345 (N_14345,N_13896,N_13861);
nor U14346 (N_14346,N_13725,N_13718);
nor U14347 (N_14347,N_13721,N_13849);
or U14348 (N_14348,N_13972,N_13729);
nand U14349 (N_14349,N_13670,N_13903);
and U14350 (N_14350,N_13849,N_13829);
nor U14351 (N_14351,N_13747,N_13832);
and U14352 (N_14352,N_13943,N_13939);
nand U14353 (N_14353,N_13966,N_13942);
nor U14354 (N_14354,N_13906,N_13620);
and U14355 (N_14355,N_13630,N_13837);
nand U14356 (N_14356,N_13854,N_13851);
nand U14357 (N_14357,N_13959,N_13620);
or U14358 (N_14358,N_13619,N_13819);
nand U14359 (N_14359,N_13805,N_13887);
xnor U14360 (N_14360,N_13865,N_13746);
nor U14361 (N_14361,N_13972,N_13934);
xor U14362 (N_14362,N_13847,N_13879);
nand U14363 (N_14363,N_13786,N_13905);
nand U14364 (N_14364,N_13907,N_13811);
nand U14365 (N_14365,N_13934,N_13980);
or U14366 (N_14366,N_13676,N_13844);
nor U14367 (N_14367,N_13759,N_13803);
or U14368 (N_14368,N_13614,N_13816);
and U14369 (N_14369,N_13983,N_13761);
or U14370 (N_14370,N_13615,N_13824);
nand U14371 (N_14371,N_13897,N_13739);
and U14372 (N_14372,N_13825,N_13747);
and U14373 (N_14373,N_13602,N_13653);
and U14374 (N_14374,N_13828,N_13796);
nor U14375 (N_14375,N_13751,N_13908);
or U14376 (N_14376,N_13724,N_13766);
nand U14377 (N_14377,N_13981,N_13971);
nor U14378 (N_14378,N_13912,N_13963);
nor U14379 (N_14379,N_13618,N_13984);
nand U14380 (N_14380,N_13778,N_13730);
or U14381 (N_14381,N_13926,N_13961);
or U14382 (N_14382,N_13645,N_13732);
nor U14383 (N_14383,N_13699,N_13817);
or U14384 (N_14384,N_13831,N_13988);
and U14385 (N_14385,N_13746,N_13674);
or U14386 (N_14386,N_13931,N_13949);
nor U14387 (N_14387,N_13707,N_13852);
nor U14388 (N_14388,N_13637,N_13870);
nor U14389 (N_14389,N_13682,N_13650);
and U14390 (N_14390,N_13683,N_13727);
or U14391 (N_14391,N_13993,N_13752);
and U14392 (N_14392,N_13647,N_13865);
nor U14393 (N_14393,N_13884,N_13694);
xnor U14394 (N_14394,N_13854,N_13849);
and U14395 (N_14395,N_13651,N_13960);
or U14396 (N_14396,N_13655,N_13621);
and U14397 (N_14397,N_13892,N_13829);
or U14398 (N_14398,N_13779,N_13933);
or U14399 (N_14399,N_13861,N_13827);
and U14400 (N_14400,N_14154,N_14391);
or U14401 (N_14401,N_14146,N_14346);
or U14402 (N_14402,N_14311,N_14290);
or U14403 (N_14403,N_14174,N_14240);
or U14404 (N_14404,N_14087,N_14375);
and U14405 (N_14405,N_14245,N_14171);
nand U14406 (N_14406,N_14166,N_14210);
and U14407 (N_14407,N_14119,N_14093);
or U14408 (N_14408,N_14058,N_14274);
and U14409 (N_14409,N_14017,N_14080);
and U14410 (N_14410,N_14392,N_14239);
and U14411 (N_14411,N_14161,N_14047);
nor U14412 (N_14412,N_14264,N_14013);
and U14413 (N_14413,N_14106,N_14066);
or U14414 (N_14414,N_14319,N_14000);
and U14415 (N_14415,N_14082,N_14107);
nor U14416 (N_14416,N_14307,N_14374);
or U14417 (N_14417,N_14026,N_14004);
and U14418 (N_14418,N_14155,N_14356);
nor U14419 (N_14419,N_14257,N_14123);
nand U14420 (N_14420,N_14387,N_14362);
nor U14421 (N_14421,N_14364,N_14286);
or U14422 (N_14422,N_14011,N_14014);
or U14423 (N_14423,N_14215,N_14353);
or U14424 (N_14424,N_14042,N_14332);
nand U14425 (N_14425,N_14037,N_14149);
or U14426 (N_14426,N_14313,N_14314);
or U14427 (N_14427,N_14061,N_14041);
nor U14428 (N_14428,N_14358,N_14233);
nand U14429 (N_14429,N_14386,N_14191);
or U14430 (N_14430,N_14381,N_14323);
or U14431 (N_14431,N_14320,N_14009);
and U14432 (N_14432,N_14018,N_14217);
and U14433 (N_14433,N_14095,N_14071);
and U14434 (N_14434,N_14310,N_14388);
nor U14435 (N_14435,N_14044,N_14079);
nor U14436 (N_14436,N_14331,N_14135);
or U14437 (N_14437,N_14315,N_14393);
and U14438 (N_14438,N_14198,N_14345);
nand U14439 (N_14439,N_14192,N_14275);
and U14440 (N_14440,N_14163,N_14228);
nor U14441 (N_14441,N_14103,N_14196);
or U14442 (N_14442,N_14350,N_14060);
nand U14443 (N_14443,N_14394,N_14202);
or U14444 (N_14444,N_14164,N_14033);
nand U14445 (N_14445,N_14298,N_14039);
nand U14446 (N_14446,N_14136,N_14302);
or U14447 (N_14447,N_14281,N_14074);
or U14448 (N_14448,N_14208,N_14390);
nand U14449 (N_14449,N_14351,N_14325);
and U14450 (N_14450,N_14005,N_14175);
nor U14451 (N_14451,N_14069,N_14101);
and U14452 (N_14452,N_14089,N_14102);
nor U14453 (N_14453,N_14088,N_14295);
nand U14454 (N_14454,N_14382,N_14186);
or U14455 (N_14455,N_14024,N_14395);
or U14456 (N_14456,N_14316,N_14040);
and U14457 (N_14457,N_14100,N_14188);
and U14458 (N_14458,N_14104,N_14105);
and U14459 (N_14459,N_14068,N_14056);
or U14460 (N_14460,N_14299,N_14214);
nand U14461 (N_14461,N_14229,N_14195);
nand U14462 (N_14462,N_14283,N_14049);
nand U14463 (N_14463,N_14126,N_14322);
and U14464 (N_14464,N_14021,N_14031);
or U14465 (N_14465,N_14296,N_14083);
nand U14466 (N_14466,N_14055,N_14389);
and U14467 (N_14467,N_14212,N_14054);
xor U14468 (N_14468,N_14289,N_14029);
nand U14469 (N_14469,N_14181,N_14179);
nand U14470 (N_14470,N_14177,N_14365);
nor U14471 (N_14471,N_14063,N_14216);
nor U14472 (N_14472,N_14222,N_14372);
nand U14473 (N_14473,N_14232,N_14246);
or U14474 (N_14474,N_14151,N_14006);
nor U14475 (N_14475,N_14116,N_14184);
or U14476 (N_14476,N_14197,N_14248);
nor U14477 (N_14477,N_14090,N_14007);
and U14478 (N_14478,N_14237,N_14273);
or U14479 (N_14479,N_14276,N_14303);
nor U14480 (N_14480,N_14140,N_14287);
nor U14481 (N_14481,N_14318,N_14204);
nor U14482 (N_14482,N_14213,N_14280);
nor U14483 (N_14483,N_14050,N_14189);
nand U14484 (N_14484,N_14262,N_14277);
nor U14485 (N_14485,N_14341,N_14397);
or U14486 (N_14486,N_14003,N_14027);
and U14487 (N_14487,N_14187,N_14019);
nor U14488 (N_14488,N_14131,N_14371);
or U14489 (N_14489,N_14025,N_14373);
and U14490 (N_14490,N_14355,N_14279);
or U14491 (N_14491,N_14053,N_14225);
nand U14492 (N_14492,N_14002,N_14183);
or U14493 (N_14493,N_14010,N_14162);
and U14494 (N_14494,N_14076,N_14038);
nand U14495 (N_14495,N_14152,N_14122);
nand U14496 (N_14496,N_14261,N_14172);
nand U14497 (N_14497,N_14270,N_14130);
or U14498 (N_14498,N_14156,N_14115);
or U14499 (N_14499,N_14267,N_14340);
and U14500 (N_14500,N_14297,N_14221);
nand U14501 (N_14501,N_14160,N_14158);
or U14502 (N_14502,N_14059,N_14159);
and U14503 (N_14503,N_14361,N_14255);
or U14504 (N_14504,N_14075,N_14077);
nor U14505 (N_14505,N_14343,N_14078);
and U14506 (N_14506,N_14167,N_14224);
nor U14507 (N_14507,N_14098,N_14070);
nand U14508 (N_14508,N_14134,N_14338);
or U14509 (N_14509,N_14265,N_14327);
and U14510 (N_14510,N_14032,N_14384);
nand U14511 (N_14511,N_14243,N_14133);
and U14512 (N_14512,N_14023,N_14293);
or U14513 (N_14513,N_14052,N_14157);
nor U14514 (N_14514,N_14139,N_14112);
nand U14515 (N_14515,N_14263,N_14118);
or U14516 (N_14516,N_14370,N_14254);
or U14517 (N_14517,N_14241,N_14178);
nand U14518 (N_14518,N_14148,N_14360);
and U14519 (N_14519,N_14120,N_14234);
or U14520 (N_14520,N_14301,N_14312);
or U14521 (N_14521,N_14352,N_14142);
nor U14522 (N_14522,N_14128,N_14269);
nand U14523 (N_14523,N_14342,N_14097);
nor U14524 (N_14524,N_14376,N_14073);
nand U14525 (N_14525,N_14236,N_14380);
and U14526 (N_14526,N_14379,N_14207);
nand U14527 (N_14527,N_14008,N_14141);
nor U14528 (N_14528,N_14253,N_14121);
nand U14529 (N_14529,N_14377,N_14266);
nor U14530 (N_14530,N_14190,N_14094);
nor U14531 (N_14531,N_14045,N_14194);
or U14532 (N_14532,N_14304,N_14065);
and U14533 (N_14533,N_14334,N_14231);
or U14534 (N_14534,N_14125,N_14200);
and U14535 (N_14535,N_14220,N_14369);
or U14536 (N_14536,N_14317,N_14012);
or U14537 (N_14537,N_14051,N_14099);
and U14538 (N_14538,N_14378,N_14034);
nor U14539 (N_14539,N_14367,N_14291);
nor U14540 (N_14540,N_14258,N_14235);
nor U14541 (N_14541,N_14227,N_14336);
or U14542 (N_14542,N_14064,N_14242);
and U14543 (N_14543,N_14249,N_14288);
nor U14544 (N_14544,N_14043,N_14169);
or U14545 (N_14545,N_14294,N_14137);
nand U14546 (N_14546,N_14305,N_14324);
or U14547 (N_14547,N_14252,N_14330);
nand U14548 (N_14548,N_14218,N_14205);
and U14549 (N_14549,N_14359,N_14337);
nand U14550 (N_14550,N_14272,N_14201);
or U14551 (N_14551,N_14015,N_14357);
or U14552 (N_14552,N_14284,N_14339);
nand U14553 (N_14553,N_14247,N_14129);
xnor U14554 (N_14554,N_14030,N_14399);
nand U14555 (N_14555,N_14092,N_14072);
nand U14556 (N_14556,N_14168,N_14259);
nand U14557 (N_14557,N_14117,N_14292);
or U14558 (N_14558,N_14203,N_14383);
or U14559 (N_14559,N_14036,N_14271);
nor U14560 (N_14560,N_14348,N_14385);
and U14561 (N_14561,N_14326,N_14109);
or U14562 (N_14562,N_14182,N_14321);
nor U14563 (N_14563,N_14022,N_14165);
and U14564 (N_14564,N_14368,N_14084);
or U14565 (N_14565,N_14085,N_14398);
and U14566 (N_14566,N_14354,N_14028);
or U14567 (N_14567,N_14329,N_14211);
nor U14568 (N_14568,N_14108,N_14113);
and U14569 (N_14569,N_14244,N_14285);
and U14570 (N_14570,N_14153,N_14268);
and U14571 (N_14571,N_14138,N_14173);
and U14572 (N_14572,N_14335,N_14086);
nor U14573 (N_14573,N_14176,N_14127);
or U14574 (N_14574,N_14219,N_14349);
nand U14575 (N_14575,N_14111,N_14250);
or U14576 (N_14576,N_14150,N_14209);
or U14577 (N_14577,N_14396,N_14282);
nand U14578 (N_14578,N_14230,N_14020);
or U14579 (N_14579,N_14260,N_14180);
nand U14580 (N_14580,N_14147,N_14016);
and U14581 (N_14581,N_14223,N_14057);
or U14582 (N_14582,N_14143,N_14226);
nor U14583 (N_14583,N_14001,N_14035);
nand U14584 (N_14584,N_14096,N_14251);
nor U14585 (N_14585,N_14132,N_14193);
nand U14586 (N_14586,N_14110,N_14300);
and U14587 (N_14587,N_14046,N_14067);
nor U14588 (N_14588,N_14145,N_14363);
and U14589 (N_14589,N_14124,N_14048);
or U14590 (N_14590,N_14333,N_14344);
nand U14591 (N_14591,N_14185,N_14309);
and U14592 (N_14592,N_14366,N_14278);
nor U14593 (N_14593,N_14062,N_14170);
and U14594 (N_14594,N_14256,N_14206);
nor U14595 (N_14595,N_14347,N_14081);
nor U14596 (N_14596,N_14199,N_14328);
nor U14597 (N_14597,N_14114,N_14238);
nand U14598 (N_14598,N_14144,N_14306);
nor U14599 (N_14599,N_14091,N_14308);
nand U14600 (N_14600,N_14124,N_14147);
nor U14601 (N_14601,N_14300,N_14214);
nor U14602 (N_14602,N_14275,N_14207);
or U14603 (N_14603,N_14284,N_14312);
nand U14604 (N_14604,N_14332,N_14312);
or U14605 (N_14605,N_14262,N_14128);
nand U14606 (N_14606,N_14275,N_14120);
and U14607 (N_14607,N_14369,N_14123);
and U14608 (N_14608,N_14153,N_14200);
and U14609 (N_14609,N_14383,N_14195);
nor U14610 (N_14610,N_14195,N_14063);
or U14611 (N_14611,N_14300,N_14210);
nand U14612 (N_14612,N_14089,N_14148);
or U14613 (N_14613,N_14379,N_14022);
nand U14614 (N_14614,N_14040,N_14329);
or U14615 (N_14615,N_14320,N_14308);
or U14616 (N_14616,N_14039,N_14068);
and U14617 (N_14617,N_14053,N_14061);
nand U14618 (N_14618,N_14308,N_14143);
and U14619 (N_14619,N_14157,N_14213);
or U14620 (N_14620,N_14154,N_14181);
nand U14621 (N_14621,N_14076,N_14391);
and U14622 (N_14622,N_14019,N_14110);
or U14623 (N_14623,N_14169,N_14175);
nor U14624 (N_14624,N_14263,N_14115);
and U14625 (N_14625,N_14040,N_14240);
nand U14626 (N_14626,N_14115,N_14352);
or U14627 (N_14627,N_14138,N_14041);
or U14628 (N_14628,N_14198,N_14365);
or U14629 (N_14629,N_14060,N_14079);
and U14630 (N_14630,N_14043,N_14305);
and U14631 (N_14631,N_14270,N_14235);
and U14632 (N_14632,N_14101,N_14117);
or U14633 (N_14633,N_14252,N_14340);
and U14634 (N_14634,N_14354,N_14157);
nor U14635 (N_14635,N_14220,N_14136);
and U14636 (N_14636,N_14123,N_14111);
xnor U14637 (N_14637,N_14169,N_14218);
and U14638 (N_14638,N_14214,N_14363);
or U14639 (N_14639,N_14183,N_14063);
nand U14640 (N_14640,N_14154,N_14341);
nand U14641 (N_14641,N_14394,N_14215);
or U14642 (N_14642,N_14133,N_14227);
and U14643 (N_14643,N_14275,N_14239);
nand U14644 (N_14644,N_14055,N_14078);
or U14645 (N_14645,N_14369,N_14170);
nor U14646 (N_14646,N_14094,N_14033);
nand U14647 (N_14647,N_14147,N_14371);
and U14648 (N_14648,N_14074,N_14067);
nor U14649 (N_14649,N_14275,N_14008);
and U14650 (N_14650,N_14286,N_14395);
and U14651 (N_14651,N_14390,N_14233);
or U14652 (N_14652,N_14341,N_14076);
or U14653 (N_14653,N_14316,N_14063);
nand U14654 (N_14654,N_14000,N_14303);
and U14655 (N_14655,N_14345,N_14172);
and U14656 (N_14656,N_14188,N_14159);
or U14657 (N_14657,N_14121,N_14206);
or U14658 (N_14658,N_14178,N_14048);
and U14659 (N_14659,N_14099,N_14056);
or U14660 (N_14660,N_14096,N_14150);
nand U14661 (N_14661,N_14167,N_14225);
and U14662 (N_14662,N_14184,N_14026);
nand U14663 (N_14663,N_14312,N_14242);
nor U14664 (N_14664,N_14122,N_14370);
or U14665 (N_14665,N_14158,N_14032);
nand U14666 (N_14666,N_14154,N_14158);
nor U14667 (N_14667,N_14144,N_14346);
nand U14668 (N_14668,N_14270,N_14125);
nand U14669 (N_14669,N_14291,N_14035);
and U14670 (N_14670,N_14279,N_14117);
nor U14671 (N_14671,N_14393,N_14225);
nand U14672 (N_14672,N_14012,N_14292);
or U14673 (N_14673,N_14228,N_14115);
nor U14674 (N_14674,N_14369,N_14146);
or U14675 (N_14675,N_14055,N_14163);
nor U14676 (N_14676,N_14095,N_14185);
and U14677 (N_14677,N_14136,N_14131);
nand U14678 (N_14678,N_14016,N_14309);
or U14679 (N_14679,N_14044,N_14048);
and U14680 (N_14680,N_14319,N_14390);
and U14681 (N_14681,N_14068,N_14262);
or U14682 (N_14682,N_14026,N_14074);
nor U14683 (N_14683,N_14056,N_14242);
nor U14684 (N_14684,N_14360,N_14341);
and U14685 (N_14685,N_14397,N_14320);
or U14686 (N_14686,N_14383,N_14284);
or U14687 (N_14687,N_14115,N_14099);
and U14688 (N_14688,N_14106,N_14368);
nand U14689 (N_14689,N_14367,N_14047);
nor U14690 (N_14690,N_14101,N_14240);
and U14691 (N_14691,N_14388,N_14108);
or U14692 (N_14692,N_14217,N_14152);
nor U14693 (N_14693,N_14294,N_14389);
or U14694 (N_14694,N_14272,N_14000);
or U14695 (N_14695,N_14238,N_14010);
nor U14696 (N_14696,N_14382,N_14335);
and U14697 (N_14697,N_14113,N_14227);
and U14698 (N_14698,N_14092,N_14194);
nand U14699 (N_14699,N_14239,N_14290);
nor U14700 (N_14700,N_14212,N_14142);
or U14701 (N_14701,N_14081,N_14284);
or U14702 (N_14702,N_14125,N_14123);
nor U14703 (N_14703,N_14256,N_14325);
or U14704 (N_14704,N_14376,N_14220);
xnor U14705 (N_14705,N_14366,N_14190);
nand U14706 (N_14706,N_14194,N_14181);
nand U14707 (N_14707,N_14374,N_14294);
nor U14708 (N_14708,N_14107,N_14047);
or U14709 (N_14709,N_14300,N_14087);
nor U14710 (N_14710,N_14048,N_14095);
or U14711 (N_14711,N_14009,N_14072);
nand U14712 (N_14712,N_14282,N_14382);
nand U14713 (N_14713,N_14339,N_14116);
or U14714 (N_14714,N_14076,N_14161);
or U14715 (N_14715,N_14295,N_14004);
nor U14716 (N_14716,N_14268,N_14277);
nor U14717 (N_14717,N_14042,N_14099);
and U14718 (N_14718,N_14093,N_14153);
nor U14719 (N_14719,N_14146,N_14389);
nor U14720 (N_14720,N_14138,N_14099);
nand U14721 (N_14721,N_14357,N_14398);
and U14722 (N_14722,N_14033,N_14293);
xnor U14723 (N_14723,N_14313,N_14078);
or U14724 (N_14724,N_14070,N_14075);
nor U14725 (N_14725,N_14132,N_14094);
nor U14726 (N_14726,N_14150,N_14352);
or U14727 (N_14727,N_14004,N_14041);
nand U14728 (N_14728,N_14324,N_14126);
or U14729 (N_14729,N_14345,N_14382);
or U14730 (N_14730,N_14298,N_14287);
nor U14731 (N_14731,N_14148,N_14190);
nand U14732 (N_14732,N_14231,N_14365);
and U14733 (N_14733,N_14190,N_14167);
nor U14734 (N_14734,N_14366,N_14353);
or U14735 (N_14735,N_14051,N_14215);
and U14736 (N_14736,N_14076,N_14031);
or U14737 (N_14737,N_14364,N_14021);
nand U14738 (N_14738,N_14353,N_14314);
or U14739 (N_14739,N_14260,N_14005);
or U14740 (N_14740,N_14383,N_14236);
nor U14741 (N_14741,N_14361,N_14219);
nor U14742 (N_14742,N_14278,N_14049);
nand U14743 (N_14743,N_14225,N_14130);
nor U14744 (N_14744,N_14376,N_14224);
nand U14745 (N_14745,N_14186,N_14227);
nor U14746 (N_14746,N_14292,N_14176);
and U14747 (N_14747,N_14131,N_14149);
and U14748 (N_14748,N_14055,N_14300);
and U14749 (N_14749,N_14252,N_14229);
nand U14750 (N_14750,N_14230,N_14052);
nand U14751 (N_14751,N_14058,N_14008);
and U14752 (N_14752,N_14293,N_14325);
nor U14753 (N_14753,N_14067,N_14092);
nor U14754 (N_14754,N_14341,N_14149);
and U14755 (N_14755,N_14115,N_14054);
nor U14756 (N_14756,N_14112,N_14178);
and U14757 (N_14757,N_14318,N_14052);
xor U14758 (N_14758,N_14271,N_14286);
nor U14759 (N_14759,N_14329,N_14212);
nand U14760 (N_14760,N_14254,N_14208);
and U14761 (N_14761,N_14187,N_14374);
or U14762 (N_14762,N_14335,N_14176);
nor U14763 (N_14763,N_14186,N_14061);
and U14764 (N_14764,N_14106,N_14212);
nor U14765 (N_14765,N_14192,N_14232);
and U14766 (N_14766,N_14255,N_14138);
nand U14767 (N_14767,N_14039,N_14087);
or U14768 (N_14768,N_14347,N_14094);
nand U14769 (N_14769,N_14180,N_14385);
and U14770 (N_14770,N_14382,N_14249);
nand U14771 (N_14771,N_14206,N_14039);
nand U14772 (N_14772,N_14033,N_14038);
nand U14773 (N_14773,N_14202,N_14241);
or U14774 (N_14774,N_14382,N_14213);
nand U14775 (N_14775,N_14322,N_14174);
or U14776 (N_14776,N_14165,N_14003);
and U14777 (N_14777,N_14038,N_14182);
nor U14778 (N_14778,N_14104,N_14066);
nand U14779 (N_14779,N_14187,N_14185);
or U14780 (N_14780,N_14200,N_14245);
and U14781 (N_14781,N_14270,N_14338);
nand U14782 (N_14782,N_14148,N_14124);
or U14783 (N_14783,N_14035,N_14378);
or U14784 (N_14784,N_14173,N_14186);
or U14785 (N_14785,N_14286,N_14134);
or U14786 (N_14786,N_14200,N_14372);
or U14787 (N_14787,N_14210,N_14121);
or U14788 (N_14788,N_14336,N_14077);
and U14789 (N_14789,N_14377,N_14378);
or U14790 (N_14790,N_14257,N_14027);
nor U14791 (N_14791,N_14166,N_14379);
and U14792 (N_14792,N_14314,N_14345);
or U14793 (N_14793,N_14276,N_14048);
nand U14794 (N_14794,N_14179,N_14390);
or U14795 (N_14795,N_14240,N_14287);
nand U14796 (N_14796,N_14279,N_14320);
xnor U14797 (N_14797,N_14295,N_14040);
nand U14798 (N_14798,N_14396,N_14073);
nor U14799 (N_14799,N_14029,N_14151);
or U14800 (N_14800,N_14493,N_14476);
nand U14801 (N_14801,N_14485,N_14488);
nand U14802 (N_14802,N_14451,N_14696);
nor U14803 (N_14803,N_14791,N_14763);
or U14804 (N_14804,N_14608,N_14446);
and U14805 (N_14805,N_14531,N_14680);
nand U14806 (N_14806,N_14430,N_14676);
or U14807 (N_14807,N_14606,N_14486);
nor U14808 (N_14808,N_14668,N_14675);
nor U14809 (N_14809,N_14428,N_14739);
or U14810 (N_14810,N_14586,N_14778);
nor U14811 (N_14811,N_14655,N_14695);
nand U14812 (N_14812,N_14556,N_14706);
nand U14813 (N_14813,N_14440,N_14536);
or U14814 (N_14814,N_14458,N_14713);
nor U14815 (N_14815,N_14429,N_14513);
and U14816 (N_14816,N_14540,N_14403);
nand U14817 (N_14817,N_14424,N_14756);
and U14818 (N_14818,N_14598,N_14745);
or U14819 (N_14819,N_14770,N_14640);
nor U14820 (N_14820,N_14677,N_14688);
and U14821 (N_14821,N_14617,N_14738);
nand U14822 (N_14822,N_14457,N_14796);
nand U14823 (N_14823,N_14495,N_14682);
nand U14824 (N_14824,N_14666,N_14492);
or U14825 (N_14825,N_14530,N_14632);
or U14826 (N_14826,N_14413,N_14714);
nand U14827 (N_14827,N_14523,N_14537);
and U14828 (N_14828,N_14623,N_14498);
nand U14829 (N_14829,N_14538,N_14618);
nor U14830 (N_14830,N_14605,N_14471);
or U14831 (N_14831,N_14400,N_14685);
nor U14832 (N_14832,N_14636,N_14544);
nand U14833 (N_14833,N_14559,N_14445);
nor U14834 (N_14834,N_14644,N_14542);
nand U14835 (N_14835,N_14747,N_14438);
xnor U14836 (N_14836,N_14522,N_14748);
and U14837 (N_14837,N_14405,N_14555);
nor U14838 (N_14838,N_14726,N_14669);
nor U14839 (N_14839,N_14639,N_14592);
or U14840 (N_14840,N_14734,N_14594);
or U14841 (N_14841,N_14414,N_14715);
nand U14842 (N_14842,N_14506,N_14466);
and U14843 (N_14843,N_14736,N_14401);
nand U14844 (N_14844,N_14439,N_14661);
and U14845 (N_14845,N_14443,N_14690);
and U14846 (N_14846,N_14474,N_14742);
and U14847 (N_14847,N_14683,N_14731);
nor U14848 (N_14848,N_14590,N_14789);
nand U14849 (N_14849,N_14664,N_14601);
nand U14850 (N_14850,N_14635,N_14681);
nand U14851 (N_14851,N_14417,N_14477);
or U14852 (N_14852,N_14535,N_14779);
nand U14853 (N_14853,N_14546,N_14660);
nor U14854 (N_14854,N_14648,N_14687);
and U14855 (N_14855,N_14580,N_14702);
nor U14856 (N_14856,N_14479,N_14788);
nand U14857 (N_14857,N_14557,N_14735);
nand U14858 (N_14858,N_14615,N_14565);
nand U14859 (N_14859,N_14525,N_14611);
or U14860 (N_14860,N_14693,N_14689);
and U14861 (N_14861,N_14776,N_14434);
and U14862 (N_14862,N_14646,N_14772);
and U14863 (N_14863,N_14613,N_14780);
or U14864 (N_14864,N_14614,N_14470);
nand U14865 (N_14865,N_14781,N_14785);
nor U14866 (N_14866,N_14421,N_14643);
and U14867 (N_14867,N_14743,N_14444);
nand U14868 (N_14868,N_14452,N_14799);
nor U14869 (N_14869,N_14566,N_14719);
or U14870 (N_14870,N_14751,N_14459);
nand U14871 (N_14871,N_14449,N_14497);
nand U14872 (N_14872,N_14589,N_14765);
nor U14873 (N_14873,N_14588,N_14600);
or U14874 (N_14874,N_14496,N_14527);
and U14875 (N_14875,N_14626,N_14610);
and U14876 (N_14876,N_14411,N_14408);
nand U14877 (N_14877,N_14460,N_14732);
nor U14878 (N_14878,N_14532,N_14426);
nand U14879 (N_14879,N_14754,N_14563);
nand U14880 (N_14880,N_14774,N_14507);
nand U14881 (N_14881,N_14679,N_14575);
and U14882 (N_14882,N_14698,N_14511);
and U14883 (N_14883,N_14427,N_14553);
and U14884 (N_14884,N_14447,N_14435);
and U14885 (N_14885,N_14595,N_14518);
and U14886 (N_14886,N_14528,N_14755);
nor U14887 (N_14887,N_14673,N_14609);
nor U14888 (N_14888,N_14746,N_14656);
and U14889 (N_14889,N_14490,N_14415);
and U14890 (N_14890,N_14771,N_14792);
nand U14891 (N_14891,N_14436,N_14469);
and U14892 (N_14892,N_14450,N_14412);
nand U14893 (N_14893,N_14596,N_14637);
or U14894 (N_14894,N_14455,N_14517);
or U14895 (N_14895,N_14684,N_14521);
nand U14896 (N_14896,N_14552,N_14561);
or U14897 (N_14897,N_14797,N_14597);
nor U14898 (N_14898,N_14541,N_14549);
nand U14899 (N_14899,N_14501,N_14749);
nand U14900 (N_14900,N_14509,N_14691);
nor U14901 (N_14901,N_14694,N_14423);
nand U14902 (N_14902,N_14526,N_14651);
nand U14903 (N_14903,N_14489,N_14621);
nand U14904 (N_14904,N_14456,N_14578);
and U14905 (N_14905,N_14573,N_14599);
and U14906 (N_14906,N_14545,N_14551);
nor U14907 (N_14907,N_14583,N_14422);
nand U14908 (N_14908,N_14692,N_14409);
or U14909 (N_14909,N_14529,N_14464);
and U14910 (N_14910,N_14753,N_14487);
nor U14911 (N_14911,N_14752,N_14767);
nand U14912 (N_14912,N_14775,N_14560);
and U14913 (N_14913,N_14725,N_14524);
and U14914 (N_14914,N_14473,N_14442);
or U14915 (N_14915,N_14625,N_14783);
or U14916 (N_14916,N_14717,N_14795);
or U14917 (N_14917,N_14463,N_14678);
or U14918 (N_14918,N_14494,N_14520);
and U14919 (N_14919,N_14558,N_14467);
nor U14920 (N_14920,N_14758,N_14570);
nand U14921 (N_14921,N_14616,N_14480);
nor U14922 (N_14922,N_14441,N_14432);
nand U14923 (N_14923,N_14708,N_14741);
nand U14924 (N_14924,N_14483,N_14645);
nand U14925 (N_14925,N_14419,N_14711);
and U14926 (N_14926,N_14550,N_14571);
or U14927 (N_14927,N_14649,N_14554);
or U14928 (N_14928,N_14504,N_14612);
or U14929 (N_14929,N_14505,N_14630);
and U14930 (N_14930,N_14663,N_14420);
nand U14931 (N_14931,N_14707,N_14410);
and U14932 (N_14932,N_14431,N_14515);
nor U14933 (N_14933,N_14574,N_14568);
nor U14934 (N_14934,N_14777,N_14634);
nor U14935 (N_14935,N_14622,N_14737);
xor U14936 (N_14936,N_14603,N_14500);
nand U14937 (N_14937,N_14567,N_14629);
nor U14938 (N_14938,N_14654,N_14465);
nor U14939 (N_14939,N_14516,N_14760);
and U14940 (N_14940,N_14533,N_14723);
and U14941 (N_14941,N_14740,N_14703);
nor U14942 (N_14942,N_14793,N_14562);
and U14943 (N_14943,N_14667,N_14712);
nor U14944 (N_14944,N_14461,N_14786);
nor U14945 (N_14945,N_14733,N_14619);
and U14946 (N_14946,N_14468,N_14766);
nand U14947 (N_14947,N_14425,N_14761);
nor U14948 (N_14948,N_14718,N_14462);
and U14949 (N_14949,N_14716,N_14728);
or U14950 (N_14950,N_14478,N_14404);
or U14951 (N_14951,N_14638,N_14534);
nand U14952 (N_14952,N_14699,N_14674);
or U14953 (N_14953,N_14790,N_14794);
nor U14954 (N_14954,N_14482,N_14407);
or U14955 (N_14955,N_14631,N_14647);
and U14956 (N_14956,N_14710,N_14577);
and U14957 (N_14957,N_14762,N_14508);
nor U14958 (N_14958,N_14579,N_14769);
nor U14959 (N_14959,N_14418,N_14481);
and U14960 (N_14960,N_14670,N_14484);
nand U14961 (N_14961,N_14593,N_14620);
nand U14962 (N_14962,N_14642,N_14650);
nand U14963 (N_14963,N_14773,N_14705);
and U14964 (N_14964,N_14709,N_14416);
or U14965 (N_14965,N_14433,N_14581);
and U14966 (N_14966,N_14624,N_14502);
or U14967 (N_14967,N_14744,N_14548);
nand U14968 (N_14968,N_14491,N_14759);
and U14969 (N_14969,N_14700,N_14787);
nand U14970 (N_14970,N_14628,N_14768);
nor U14971 (N_14971,N_14627,N_14569);
or U14972 (N_14972,N_14453,N_14582);
nand U14973 (N_14973,N_14727,N_14475);
and U14974 (N_14974,N_14437,N_14704);
or U14975 (N_14975,N_14662,N_14730);
nand U14976 (N_14976,N_14503,N_14701);
or U14977 (N_14977,N_14454,N_14672);
nor U14978 (N_14978,N_14607,N_14543);
or U14979 (N_14979,N_14697,N_14499);
and U14980 (N_14980,N_14729,N_14572);
nor U14981 (N_14981,N_14750,N_14539);
and U14982 (N_14982,N_14721,N_14764);
nand U14983 (N_14983,N_14585,N_14653);
nand U14984 (N_14984,N_14402,N_14576);
and U14985 (N_14985,N_14798,N_14720);
and U14986 (N_14986,N_14406,N_14724);
nand U14987 (N_14987,N_14686,N_14652);
nor U14988 (N_14988,N_14510,N_14448);
and U14989 (N_14989,N_14472,N_14591);
nand U14990 (N_14990,N_14519,N_14514);
and U14991 (N_14991,N_14659,N_14658);
and U14992 (N_14992,N_14757,N_14584);
and U14993 (N_14993,N_14784,N_14512);
nor U14994 (N_14994,N_14665,N_14657);
nor U14995 (N_14995,N_14604,N_14641);
nor U14996 (N_14996,N_14547,N_14602);
and U14997 (N_14997,N_14564,N_14782);
and U14998 (N_14998,N_14722,N_14633);
nor U14999 (N_14999,N_14587,N_14671);
and U15000 (N_15000,N_14440,N_14786);
xnor U15001 (N_15001,N_14745,N_14522);
or U15002 (N_15002,N_14617,N_14489);
or U15003 (N_15003,N_14404,N_14454);
or U15004 (N_15004,N_14554,N_14571);
nor U15005 (N_15005,N_14457,N_14703);
nand U15006 (N_15006,N_14424,N_14582);
nor U15007 (N_15007,N_14630,N_14689);
or U15008 (N_15008,N_14685,N_14608);
or U15009 (N_15009,N_14451,N_14523);
nand U15010 (N_15010,N_14495,N_14633);
or U15011 (N_15011,N_14686,N_14514);
nand U15012 (N_15012,N_14425,N_14418);
nor U15013 (N_15013,N_14753,N_14455);
or U15014 (N_15014,N_14650,N_14745);
and U15015 (N_15015,N_14704,N_14438);
and U15016 (N_15016,N_14795,N_14460);
or U15017 (N_15017,N_14451,N_14699);
nor U15018 (N_15018,N_14436,N_14617);
or U15019 (N_15019,N_14707,N_14709);
xor U15020 (N_15020,N_14539,N_14599);
nand U15021 (N_15021,N_14500,N_14514);
nand U15022 (N_15022,N_14486,N_14615);
nand U15023 (N_15023,N_14419,N_14652);
nor U15024 (N_15024,N_14719,N_14524);
nand U15025 (N_15025,N_14667,N_14697);
and U15026 (N_15026,N_14481,N_14475);
nor U15027 (N_15027,N_14570,N_14703);
or U15028 (N_15028,N_14707,N_14660);
nand U15029 (N_15029,N_14720,N_14658);
or U15030 (N_15030,N_14688,N_14639);
nand U15031 (N_15031,N_14402,N_14536);
nand U15032 (N_15032,N_14701,N_14741);
and U15033 (N_15033,N_14408,N_14515);
nor U15034 (N_15034,N_14781,N_14639);
and U15035 (N_15035,N_14410,N_14546);
nand U15036 (N_15036,N_14506,N_14669);
nand U15037 (N_15037,N_14415,N_14613);
or U15038 (N_15038,N_14426,N_14469);
and U15039 (N_15039,N_14635,N_14658);
nor U15040 (N_15040,N_14695,N_14753);
or U15041 (N_15041,N_14551,N_14452);
and U15042 (N_15042,N_14453,N_14539);
nor U15043 (N_15043,N_14599,N_14767);
nor U15044 (N_15044,N_14625,N_14701);
or U15045 (N_15045,N_14598,N_14516);
and U15046 (N_15046,N_14775,N_14670);
or U15047 (N_15047,N_14770,N_14747);
nor U15048 (N_15048,N_14592,N_14734);
or U15049 (N_15049,N_14486,N_14559);
nand U15050 (N_15050,N_14400,N_14609);
nand U15051 (N_15051,N_14502,N_14769);
or U15052 (N_15052,N_14425,N_14615);
or U15053 (N_15053,N_14708,N_14798);
nand U15054 (N_15054,N_14741,N_14753);
or U15055 (N_15055,N_14786,N_14435);
nand U15056 (N_15056,N_14795,N_14405);
or U15057 (N_15057,N_14429,N_14404);
and U15058 (N_15058,N_14720,N_14750);
or U15059 (N_15059,N_14556,N_14694);
and U15060 (N_15060,N_14731,N_14689);
and U15061 (N_15061,N_14733,N_14533);
nor U15062 (N_15062,N_14538,N_14707);
or U15063 (N_15063,N_14416,N_14459);
or U15064 (N_15064,N_14662,N_14731);
and U15065 (N_15065,N_14716,N_14422);
or U15066 (N_15066,N_14509,N_14702);
nand U15067 (N_15067,N_14539,N_14682);
nor U15068 (N_15068,N_14771,N_14454);
nand U15069 (N_15069,N_14420,N_14488);
nand U15070 (N_15070,N_14509,N_14563);
nand U15071 (N_15071,N_14526,N_14718);
nand U15072 (N_15072,N_14648,N_14651);
and U15073 (N_15073,N_14618,N_14565);
nand U15074 (N_15074,N_14791,N_14579);
and U15075 (N_15075,N_14671,N_14462);
and U15076 (N_15076,N_14589,N_14532);
nor U15077 (N_15077,N_14727,N_14524);
and U15078 (N_15078,N_14508,N_14406);
nand U15079 (N_15079,N_14773,N_14730);
nor U15080 (N_15080,N_14610,N_14718);
nor U15081 (N_15081,N_14498,N_14799);
nor U15082 (N_15082,N_14696,N_14756);
nor U15083 (N_15083,N_14554,N_14494);
and U15084 (N_15084,N_14547,N_14701);
and U15085 (N_15085,N_14455,N_14764);
or U15086 (N_15086,N_14485,N_14607);
and U15087 (N_15087,N_14599,N_14422);
or U15088 (N_15088,N_14601,N_14752);
nand U15089 (N_15089,N_14444,N_14799);
and U15090 (N_15090,N_14513,N_14545);
nand U15091 (N_15091,N_14637,N_14714);
or U15092 (N_15092,N_14464,N_14691);
nand U15093 (N_15093,N_14539,N_14581);
nand U15094 (N_15094,N_14608,N_14554);
nand U15095 (N_15095,N_14752,N_14475);
and U15096 (N_15096,N_14508,N_14594);
or U15097 (N_15097,N_14786,N_14423);
nand U15098 (N_15098,N_14441,N_14474);
or U15099 (N_15099,N_14702,N_14575);
nor U15100 (N_15100,N_14597,N_14456);
and U15101 (N_15101,N_14698,N_14631);
or U15102 (N_15102,N_14788,N_14413);
nor U15103 (N_15103,N_14455,N_14794);
or U15104 (N_15104,N_14523,N_14684);
nand U15105 (N_15105,N_14632,N_14481);
and U15106 (N_15106,N_14636,N_14796);
and U15107 (N_15107,N_14426,N_14787);
and U15108 (N_15108,N_14509,N_14709);
nor U15109 (N_15109,N_14680,N_14731);
and U15110 (N_15110,N_14767,N_14474);
and U15111 (N_15111,N_14789,N_14495);
nand U15112 (N_15112,N_14610,N_14745);
nor U15113 (N_15113,N_14482,N_14516);
nor U15114 (N_15114,N_14780,N_14528);
nor U15115 (N_15115,N_14506,N_14653);
or U15116 (N_15116,N_14768,N_14734);
nor U15117 (N_15117,N_14731,N_14745);
or U15118 (N_15118,N_14739,N_14513);
or U15119 (N_15119,N_14653,N_14420);
nand U15120 (N_15120,N_14621,N_14665);
nand U15121 (N_15121,N_14748,N_14452);
nand U15122 (N_15122,N_14560,N_14401);
nand U15123 (N_15123,N_14631,N_14518);
and U15124 (N_15124,N_14777,N_14675);
and U15125 (N_15125,N_14510,N_14734);
nor U15126 (N_15126,N_14490,N_14432);
nand U15127 (N_15127,N_14693,N_14512);
nor U15128 (N_15128,N_14440,N_14407);
nor U15129 (N_15129,N_14448,N_14484);
nor U15130 (N_15130,N_14479,N_14405);
or U15131 (N_15131,N_14613,N_14453);
and U15132 (N_15132,N_14592,N_14423);
and U15133 (N_15133,N_14511,N_14691);
and U15134 (N_15134,N_14409,N_14421);
nor U15135 (N_15135,N_14772,N_14556);
or U15136 (N_15136,N_14643,N_14761);
nand U15137 (N_15137,N_14668,N_14501);
or U15138 (N_15138,N_14779,N_14700);
nor U15139 (N_15139,N_14560,N_14748);
or U15140 (N_15140,N_14749,N_14518);
or U15141 (N_15141,N_14614,N_14762);
nor U15142 (N_15142,N_14759,N_14786);
nand U15143 (N_15143,N_14567,N_14660);
nor U15144 (N_15144,N_14560,N_14679);
or U15145 (N_15145,N_14672,N_14497);
nand U15146 (N_15146,N_14799,N_14759);
nor U15147 (N_15147,N_14732,N_14404);
and U15148 (N_15148,N_14783,N_14614);
or U15149 (N_15149,N_14477,N_14743);
or U15150 (N_15150,N_14472,N_14651);
nor U15151 (N_15151,N_14536,N_14541);
and U15152 (N_15152,N_14530,N_14795);
or U15153 (N_15153,N_14730,N_14731);
nor U15154 (N_15154,N_14493,N_14531);
nand U15155 (N_15155,N_14447,N_14742);
nor U15156 (N_15156,N_14418,N_14656);
and U15157 (N_15157,N_14754,N_14444);
nor U15158 (N_15158,N_14770,N_14425);
and U15159 (N_15159,N_14575,N_14777);
nand U15160 (N_15160,N_14649,N_14787);
and U15161 (N_15161,N_14425,N_14667);
and U15162 (N_15162,N_14695,N_14551);
nor U15163 (N_15163,N_14712,N_14512);
and U15164 (N_15164,N_14674,N_14665);
or U15165 (N_15165,N_14490,N_14568);
or U15166 (N_15166,N_14769,N_14655);
nor U15167 (N_15167,N_14719,N_14643);
nor U15168 (N_15168,N_14596,N_14554);
and U15169 (N_15169,N_14617,N_14673);
nand U15170 (N_15170,N_14406,N_14530);
and U15171 (N_15171,N_14521,N_14630);
or U15172 (N_15172,N_14688,N_14708);
and U15173 (N_15173,N_14722,N_14610);
or U15174 (N_15174,N_14491,N_14768);
or U15175 (N_15175,N_14675,N_14406);
or U15176 (N_15176,N_14614,N_14495);
nor U15177 (N_15177,N_14642,N_14703);
and U15178 (N_15178,N_14666,N_14735);
and U15179 (N_15179,N_14754,N_14695);
nor U15180 (N_15180,N_14735,N_14746);
nand U15181 (N_15181,N_14706,N_14502);
nor U15182 (N_15182,N_14444,N_14565);
nand U15183 (N_15183,N_14693,N_14416);
or U15184 (N_15184,N_14463,N_14715);
and U15185 (N_15185,N_14672,N_14583);
or U15186 (N_15186,N_14752,N_14764);
nand U15187 (N_15187,N_14511,N_14553);
nand U15188 (N_15188,N_14690,N_14543);
and U15189 (N_15189,N_14739,N_14436);
and U15190 (N_15190,N_14631,N_14510);
nor U15191 (N_15191,N_14792,N_14646);
nand U15192 (N_15192,N_14499,N_14418);
nor U15193 (N_15193,N_14764,N_14715);
or U15194 (N_15194,N_14571,N_14406);
nand U15195 (N_15195,N_14670,N_14413);
nand U15196 (N_15196,N_14417,N_14653);
nor U15197 (N_15197,N_14628,N_14461);
or U15198 (N_15198,N_14600,N_14425);
nor U15199 (N_15199,N_14746,N_14467);
or U15200 (N_15200,N_15160,N_14994);
and U15201 (N_15201,N_14999,N_15033);
and U15202 (N_15202,N_14825,N_14801);
or U15203 (N_15203,N_15132,N_14865);
nand U15204 (N_15204,N_14817,N_15001);
nor U15205 (N_15205,N_14880,N_14902);
and U15206 (N_15206,N_14976,N_15028);
and U15207 (N_15207,N_14898,N_14997);
nor U15208 (N_15208,N_14978,N_14953);
nor U15209 (N_15209,N_15081,N_15049);
or U15210 (N_15210,N_14831,N_15117);
or U15211 (N_15211,N_15147,N_14908);
and U15212 (N_15212,N_15040,N_14963);
nand U15213 (N_15213,N_14847,N_15064);
nand U15214 (N_15214,N_14893,N_14934);
nor U15215 (N_15215,N_15076,N_15013);
and U15216 (N_15216,N_15120,N_15005);
or U15217 (N_15217,N_14995,N_14967);
nor U15218 (N_15218,N_14919,N_15089);
nand U15219 (N_15219,N_15181,N_14837);
nand U15220 (N_15220,N_15090,N_14887);
nand U15221 (N_15221,N_15138,N_14805);
nand U15222 (N_15222,N_14958,N_15145);
nand U15223 (N_15223,N_15131,N_14855);
or U15224 (N_15224,N_15115,N_14952);
and U15225 (N_15225,N_15103,N_15079);
and U15226 (N_15226,N_15135,N_15058);
nor U15227 (N_15227,N_14867,N_15182);
nor U15228 (N_15228,N_15169,N_15193);
nand U15229 (N_15229,N_14907,N_14929);
nand U15230 (N_15230,N_15163,N_14948);
or U15231 (N_15231,N_14913,N_14957);
nor U15232 (N_15232,N_14906,N_15039);
and U15233 (N_15233,N_15096,N_14981);
and U15234 (N_15234,N_15124,N_15179);
nand U15235 (N_15235,N_15188,N_15004);
or U15236 (N_15236,N_14979,N_15198);
nor U15237 (N_15237,N_15123,N_15034);
nor U15238 (N_15238,N_15091,N_15199);
and U15239 (N_15239,N_15152,N_14941);
and U15240 (N_15240,N_14858,N_15080);
or U15241 (N_15241,N_14848,N_14917);
nand U15242 (N_15242,N_15111,N_14925);
nand U15243 (N_15243,N_15038,N_14947);
nor U15244 (N_15244,N_15171,N_15055);
nand U15245 (N_15245,N_15108,N_14922);
nand U15246 (N_15246,N_14846,N_14830);
nand U15247 (N_15247,N_14881,N_15186);
nand U15248 (N_15248,N_15042,N_14871);
nor U15249 (N_15249,N_15074,N_15037);
nand U15250 (N_15250,N_15069,N_14804);
nor U15251 (N_15251,N_14809,N_14959);
nand U15252 (N_15252,N_15178,N_14828);
nand U15253 (N_15253,N_15194,N_15121);
nor U15254 (N_15254,N_14950,N_14905);
and U15255 (N_15255,N_14819,N_14818);
or U15256 (N_15256,N_14816,N_14935);
or U15257 (N_15257,N_14824,N_15011);
or U15258 (N_15258,N_14849,N_14859);
nor U15259 (N_15259,N_15094,N_15156);
or U15260 (N_15260,N_14872,N_14891);
nor U15261 (N_15261,N_15030,N_14875);
nand U15262 (N_15262,N_14843,N_14895);
nand U15263 (N_15263,N_14983,N_15019);
nand U15264 (N_15264,N_14856,N_15035);
and U15265 (N_15265,N_14903,N_15085);
and U15266 (N_15266,N_15029,N_15027);
nor U15267 (N_15267,N_14829,N_14901);
and U15268 (N_15268,N_15050,N_15082);
or U15269 (N_15269,N_15032,N_15105);
nor U15270 (N_15270,N_14966,N_14894);
or U15271 (N_15271,N_15003,N_14923);
nand U15272 (N_15272,N_14892,N_14803);
or U15273 (N_15273,N_15073,N_15095);
or U15274 (N_15274,N_15083,N_15067);
or U15275 (N_15275,N_15128,N_14940);
nand U15276 (N_15276,N_14810,N_14869);
nor U15277 (N_15277,N_14927,N_14971);
nor U15278 (N_15278,N_15077,N_14883);
or U15279 (N_15279,N_14945,N_15142);
nand U15280 (N_15280,N_14954,N_15144);
nand U15281 (N_15281,N_14860,N_15093);
nand U15282 (N_15282,N_14811,N_15164);
nand U15283 (N_15283,N_15018,N_15059);
or U15284 (N_15284,N_15114,N_14899);
or U15285 (N_15285,N_14862,N_14868);
nor U15286 (N_15286,N_14841,N_15167);
nor U15287 (N_15287,N_15098,N_14975);
and U15288 (N_15288,N_15158,N_14969);
and U15289 (N_15289,N_15045,N_14909);
or U15290 (N_15290,N_15066,N_15071);
or U15291 (N_15291,N_14938,N_14851);
or U15292 (N_15292,N_15173,N_14806);
or U15293 (N_15293,N_14854,N_14939);
nand U15294 (N_15294,N_14836,N_15023);
nand U15295 (N_15295,N_15172,N_15112);
nor U15296 (N_15296,N_15161,N_15187);
nand U15297 (N_15297,N_15149,N_14873);
nor U15298 (N_15298,N_15166,N_14916);
and U15299 (N_15299,N_14800,N_15168);
or U15300 (N_15300,N_15014,N_14943);
and U15301 (N_15301,N_15084,N_15010);
or U15302 (N_15302,N_14914,N_14815);
and U15303 (N_15303,N_15025,N_15107);
or U15304 (N_15304,N_14968,N_14885);
or U15305 (N_15305,N_14937,N_15113);
and U15306 (N_15306,N_15063,N_15155);
nand U15307 (N_15307,N_15002,N_15015);
nor U15308 (N_15308,N_14986,N_15136);
or U15309 (N_15309,N_14821,N_15134);
nand U15310 (N_15310,N_15106,N_14827);
nand U15311 (N_15311,N_15065,N_14834);
and U15312 (N_15312,N_14990,N_15092);
or U15313 (N_15313,N_14850,N_15052);
and U15314 (N_15314,N_14965,N_14951);
nor U15315 (N_15315,N_15129,N_15060);
nand U15316 (N_15316,N_15070,N_14845);
nand U15317 (N_15317,N_14946,N_15053);
nor U15318 (N_15318,N_15101,N_14822);
and U15319 (N_15319,N_14989,N_15174);
and U15320 (N_15320,N_14991,N_14863);
or U15321 (N_15321,N_15150,N_15009);
nor U15322 (N_15322,N_15031,N_15189);
xnor U15323 (N_15323,N_15051,N_14980);
or U15324 (N_15324,N_15097,N_15017);
or U15325 (N_15325,N_14993,N_15046);
nor U15326 (N_15326,N_14839,N_14844);
and U15327 (N_15327,N_15012,N_14866);
nor U15328 (N_15328,N_15056,N_14814);
and U15329 (N_15329,N_14942,N_14985);
or U15330 (N_15330,N_15165,N_15176);
and U15331 (N_15331,N_15127,N_15139);
nor U15332 (N_15332,N_15153,N_14802);
nand U15333 (N_15333,N_14870,N_14933);
and U15334 (N_15334,N_15148,N_15104);
nor U15335 (N_15335,N_15102,N_15020);
or U15336 (N_15336,N_14920,N_15026);
nor U15337 (N_15337,N_14921,N_14955);
nand U15338 (N_15338,N_15143,N_15125);
nand U15339 (N_15339,N_14974,N_15109);
nor U15340 (N_15340,N_15022,N_14911);
nor U15341 (N_15341,N_14879,N_15184);
and U15342 (N_15342,N_14926,N_15054);
and U15343 (N_15343,N_15110,N_14984);
or U15344 (N_15344,N_14910,N_14964);
or U15345 (N_15345,N_14884,N_15008);
or U15346 (N_15346,N_14900,N_14998);
or U15347 (N_15347,N_14813,N_14832);
nor U15348 (N_15348,N_15062,N_14931);
nand U15349 (N_15349,N_14853,N_14877);
nor U15350 (N_15350,N_14992,N_15047);
or U15351 (N_15351,N_14912,N_14932);
or U15352 (N_15352,N_14886,N_14944);
or U15353 (N_15353,N_14888,N_15075);
nand U15354 (N_15354,N_14972,N_15151);
nor U15355 (N_15355,N_14808,N_15183);
and U15356 (N_15356,N_15000,N_14823);
nor U15357 (N_15357,N_14874,N_15043);
nand U15358 (N_15358,N_14962,N_15175);
nand U15359 (N_15359,N_14960,N_15068);
nand U15360 (N_15360,N_15170,N_15087);
nand U15361 (N_15361,N_14961,N_15141);
nor U15362 (N_15362,N_15021,N_15196);
nand U15363 (N_15363,N_15086,N_15041);
nand U15364 (N_15364,N_14864,N_15061);
nor U15365 (N_15365,N_15190,N_15185);
and U15366 (N_15366,N_14982,N_14896);
and U15367 (N_15367,N_15007,N_14807);
and U15368 (N_15368,N_15197,N_15100);
nor U15369 (N_15369,N_14861,N_15146);
nor U15370 (N_15370,N_15126,N_14820);
nor U15371 (N_15371,N_15195,N_15044);
nor U15372 (N_15372,N_14897,N_14988);
or U15373 (N_15373,N_15057,N_14956);
nand U15374 (N_15374,N_15130,N_15036);
or U15375 (N_15375,N_14977,N_14915);
nor U15376 (N_15376,N_15088,N_14812);
or U15377 (N_15377,N_14949,N_15157);
nor U15378 (N_15378,N_15180,N_14842);
nand U15379 (N_15379,N_14882,N_14852);
or U15380 (N_15380,N_14890,N_14838);
nor U15381 (N_15381,N_15048,N_14930);
nor U15382 (N_15382,N_15116,N_14973);
nand U15383 (N_15383,N_15006,N_15192);
nor U15384 (N_15384,N_15137,N_14996);
or U15385 (N_15385,N_15118,N_14857);
or U15386 (N_15386,N_15072,N_14889);
nand U15387 (N_15387,N_14928,N_15162);
or U15388 (N_15388,N_15024,N_15177);
nor U15389 (N_15389,N_14876,N_14918);
and U15390 (N_15390,N_15099,N_14936);
and U15391 (N_15391,N_15016,N_15122);
nor U15392 (N_15392,N_14970,N_14878);
nor U15393 (N_15393,N_14826,N_14840);
nor U15394 (N_15394,N_15119,N_14987);
nor U15395 (N_15395,N_15078,N_15140);
nor U15396 (N_15396,N_15191,N_14904);
nor U15397 (N_15397,N_15133,N_15154);
xnor U15398 (N_15398,N_14924,N_14835);
nor U15399 (N_15399,N_14833,N_15159);
or U15400 (N_15400,N_15101,N_15161);
or U15401 (N_15401,N_14890,N_15196);
and U15402 (N_15402,N_14939,N_14917);
or U15403 (N_15403,N_15126,N_14981);
nor U15404 (N_15404,N_14972,N_14815);
nand U15405 (N_15405,N_14870,N_14978);
nand U15406 (N_15406,N_15058,N_15014);
nand U15407 (N_15407,N_15199,N_15194);
xnor U15408 (N_15408,N_14872,N_14822);
and U15409 (N_15409,N_14924,N_14945);
or U15410 (N_15410,N_15185,N_15187);
nor U15411 (N_15411,N_15165,N_15087);
and U15412 (N_15412,N_14953,N_15096);
nor U15413 (N_15413,N_14899,N_15033);
and U15414 (N_15414,N_14895,N_15074);
nand U15415 (N_15415,N_14900,N_15156);
or U15416 (N_15416,N_15184,N_15047);
or U15417 (N_15417,N_14826,N_15070);
or U15418 (N_15418,N_14866,N_15124);
or U15419 (N_15419,N_15054,N_15126);
or U15420 (N_15420,N_15117,N_14938);
or U15421 (N_15421,N_15028,N_14982);
nor U15422 (N_15422,N_14887,N_14908);
and U15423 (N_15423,N_15005,N_14802);
nand U15424 (N_15424,N_14910,N_15037);
and U15425 (N_15425,N_14927,N_14877);
nor U15426 (N_15426,N_14829,N_14967);
nor U15427 (N_15427,N_14947,N_14818);
and U15428 (N_15428,N_14975,N_14919);
nor U15429 (N_15429,N_15028,N_15065);
nand U15430 (N_15430,N_14915,N_15052);
and U15431 (N_15431,N_14810,N_14955);
nor U15432 (N_15432,N_14861,N_15061);
nor U15433 (N_15433,N_15017,N_15199);
nor U15434 (N_15434,N_14909,N_14800);
or U15435 (N_15435,N_15143,N_14907);
and U15436 (N_15436,N_14854,N_14923);
and U15437 (N_15437,N_14914,N_14922);
nand U15438 (N_15438,N_15067,N_14879);
or U15439 (N_15439,N_15167,N_15042);
nor U15440 (N_15440,N_14951,N_15142);
nor U15441 (N_15441,N_14844,N_14989);
or U15442 (N_15442,N_15048,N_14939);
or U15443 (N_15443,N_15109,N_15055);
and U15444 (N_15444,N_15023,N_14937);
nor U15445 (N_15445,N_14933,N_14895);
nand U15446 (N_15446,N_14971,N_15093);
and U15447 (N_15447,N_15106,N_15011);
and U15448 (N_15448,N_15151,N_14926);
and U15449 (N_15449,N_14994,N_14959);
nor U15450 (N_15450,N_14872,N_14859);
nand U15451 (N_15451,N_14961,N_15101);
nand U15452 (N_15452,N_14992,N_15141);
nor U15453 (N_15453,N_15180,N_14931);
or U15454 (N_15454,N_15116,N_15115);
nor U15455 (N_15455,N_15159,N_14902);
nor U15456 (N_15456,N_14948,N_14971);
nand U15457 (N_15457,N_14815,N_14968);
nand U15458 (N_15458,N_14978,N_14908);
and U15459 (N_15459,N_15033,N_14863);
nor U15460 (N_15460,N_14823,N_14924);
nand U15461 (N_15461,N_14978,N_15115);
and U15462 (N_15462,N_15115,N_14858);
nand U15463 (N_15463,N_14821,N_15004);
and U15464 (N_15464,N_15055,N_15070);
nand U15465 (N_15465,N_14881,N_14909);
nand U15466 (N_15466,N_14835,N_14906);
nand U15467 (N_15467,N_15189,N_14877);
nand U15468 (N_15468,N_14901,N_15005);
nand U15469 (N_15469,N_15089,N_15095);
or U15470 (N_15470,N_15189,N_14870);
nor U15471 (N_15471,N_14910,N_15186);
or U15472 (N_15472,N_15120,N_14810);
and U15473 (N_15473,N_14966,N_15091);
or U15474 (N_15474,N_14978,N_14945);
nor U15475 (N_15475,N_15068,N_15115);
or U15476 (N_15476,N_15027,N_15110);
and U15477 (N_15477,N_14932,N_15178);
nor U15478 (N_15478,N_14849,N_15198);
and U15479 (N_15479,N_15027,N_15122);
or U15480 (N_15480,N_15012,N_15119);
nand U15481 (N_15481,N_15063,N_14980);
and U15482 (N_15482,N_14945,N_15161);
xnor U15483 (N_15483,N_15156,N_15112);
nand U15484 (N_15484,N_15166,N_14878);
or U15485 (N_15485,N_15098,N_15000);
nand U15486 (N_15486,N_15187,N_14833);
nor U15487 (N_15487,N_15101,N_15187);
or U15488 (N_15488,N_14966,N_15105);
or U15489 (N_15489,N_15079,N_14883);
or U15490 (N_15490,N_14835,N_15004);
or U15491 (N_15491,N_15096,N_15057);
or U15492 (N_15492,N_15109,N_14973);
nand U15493 (N_15493,N_15187,N_15031);
or U15494 (N_15494,N_15019,N_14825);
or U15495 (N_15495,N_15155,N_15048);
or U15496 (N_15496,N_14891,N_15041);
nor U15497 (N_15497,N_14999,N_14836);
or U15498 (N_15498,N_15004,N_15050);
nand U15499 (N_15499,N_14879,N_15131);
and U15500 (N_15500,N_14886,N_14824);
nor U15501 (N_15501,N_14880,N_15159);
nand U15502 (N_15502,N_14929,N_14807);
and U15503 (N_15503,N_15019,N_15010);
nand U15504 (N_15504,N_15154,N_15125);
nand U15505 (N_15505,N_15011,N_15070);
nor U15506 (N_15506,N_14942,N_15160);
or U15507 (N_15507,N_14867,N_14923);
nand U15508 (N_15508,N_15096,N_14983);
nor U15509 (N_15509,N_14818,N_14993);
nor U15510 (N_15510,N_14854,N_15093);
nand U15511 (N_15511,N_14961,N_15079);
or U15512 (N_15512,N_15140,N_14851);
nor U15513 (N_15513,N_15061,N_14903);
nand U15514 (N_15514,N_15012,N_14844);
nand U15515 (N_15515,N_14975,N_14888);
and U15516 (N_15516,N_15135,N_15176);
or U15517 (N_15517,N_14993,N_14857);
or U15518 (N_15518,N_14992,N_14868);
nor U15519 (N_15519,N_15172,N_15135);
and U15520 (N_15520,N_15112,N_15085);
nor U15521 (N_15521,N_15027,N_15137);
and U15522 (N_15522,N_14839,N_14837);
nand U15523 (N_15523,N_14968,N_14801);
nor U15524 (N_15524,N_14882,N_15005);
nor U15525 (N_15525,N_15156,N_15058);
nand U15526 (N_15526,N_15029,N_15058);
or U15527 (N_15527,N_14846,N_15112);
or U15528 (N_15528,N_15163,N_15112);
nor U15529 (N_15529,N_14830,N_14955);
and U15530 (N_15530,N_14969,N_15164);
and U15531 (N_15531,N_15032,N_14835);
or U15532 (N_15532,N_14847,N_15114);
nand U15533 (N_15533,N_14814,N_15154);
or U15534 (N_15534,N_14874,N_15005);
and U15535 (N_15535,N_14986,N_14923);
nor U15536 (N_15536,N_14868,N_15059);
nand U15537 (N_15537,N_14849,N_15182);
nand U15538 (N_15538,N_15029,N_14935);
nand U15539 (N_15539,N_15158,N_14924);
and U15540 (N_15540,N_14841,N_15056);
nand U15541 (N_15541,N_14810,N_15037);
and U15542 (N_15542,N_15167,N_14896);
nand U15543 (N_15543,N_15074,N_14974);
nor U15544 (N_15544,N_14806,N_14918);
or U15545 (N_15545,N_15165,N_15135);
nand U15546 (N_15546,N_15173,N_14905);
and U15547 (N_15547,N_15125,N_15182);
nand U15548 (N_15548,N_15187,N_14885);
or U15549 (N_15549,N_14894,N_15037);
or U15550 (N_15550,N_15058,N_14979);
nor U15551 (N_15551,N_15028,N_14834);
nand U15552 (N_15552,N_14870,N_14849);
or U15553 (N_15553,N_15033,N_14937);
nor U15554 (N_15554,N_15012,N_15151);
nand U15555 (N_15555,N_15155,N_15098);
or U15556 (N_15556,N_14846,N_14897);
and U15557 (N_15557,N_15060,N_14933);
and U15558 (N_15558,N_14824,N_15161);
and U15559 (N_15559,N_14923,N_14840);
and U15560 (N_15560,N_15154,N_15169);
nand U15561 (N_15561,N_14852,N_14920);
nand U15562 (N_15562,N_15061,N_15170);
or U15563 (N_15563,N_15198,N_14974);
nor U15564 (N_15564,N_15160,N_15132);
or U15565 (N_15565,N_15080,N_15039);
nand U15566 (N_15566,N_15121,N_15019);
and U15567 (N_15567,N_14824,N_15086);
or U15568 (N_15568,N_15001,N_15175);
and U15569 (N_15569,N_15174,N_14893);
nand U15570 (N_15570,N_15038,N_15101);
or U15571 (N_15571,N_14929,N_14839);
nand U15572 (N_15572,N_15177,N_15023);
and U15573 (N_15573,N_14865,N_15051);
nand U15574 (N_15574,N_15122,N_14809);
nand U15575 (N_15575,N_15049,N_15003);
xor U15576 (N_15576,N_15130,N_14928);
nand U15577 (N_15577,N_15175,N_14849);
and U15578 (N_15578,N_15189,N_14951);
and U15579 (N_15579,N_14803,N_14813);
nand U15580 (N_15580,N_15196,N_15150);
nand U15581 (N_15581,N_15154,N_14865);
or U15582 (N_15582,N_14926,N_15133);
nand U15583 (N_15583,N_15092,N_15016);
or U15584 (N_15584,N_15135,N_15170);
or U15585 (N_15585,N_14874,N_15078);
and U15586 (N_15586,N_14810,N_15116);
and U15587 (N_15587,N_15111,N_14867);
or U15588 (N_15588,N_14972,N_15186);
or U15589 (N_15589,N_15186,N_15038);
nand U15590 (N_15590,N_14955,N_15030);
or U15591 (N_15591,N_14822,N_14827);
nand U15592 (N_15592,N_15076,N_14882);
nor U15593 (N_15593,N_15045,N_14848);
and U15594 (N_15594,N_14909,N_15114);
nor U15595 (N_15595,N_15074,N_15015);
or U15596 (N_15596,N_14925,N_15142);
nand U15597 (N_15597,N_14983,N_14927);
nor U15598 (N_15598,N_14928,N_14816);
nand U15599 (N_15599,N_15032,N_15045);
and U15600 (N_15600,N_15541,N_15335);
nor U15601 (N_15601,N_15207,N_15416);
nand U15602 (N_15602,N_15204,N_15361);
and U15603 (N_15603,N_15514,N_15376);
and U15604 (N_15604,N_15559,N_15371);
nand U15605 (N_15605,N_15283,N_15262);
or U15606 (N_15606,N_15302,N_15467);
nor U15607 (N_15607,N_15585,N_15385);
nor U15608 (N_15608,N_15466,N_15445);
or U15609 (N_15609,N_15243,N_15575);
and U15610 (N_15610,N_15460,N_15334);
and U15611 (N_15611,N_15530,N_15473);
or U15612 (N_15612,N_15446,N_15494);
nand U15613 (N_15613,N_15411,N_15496);
nand U15614 (N_15614,N_15309,N_15599);
nor U15615 (N_15615,N_15324,N_15367);
xnor U15616 (N_15616,N_15421,N_15456);
or U15617 (N_15617,N_15295,N_15423);
or U15618 (N_15618,N_15407,N_15241);
nor U15619 (N_15619,N_15248,N_15429);
and U15620 (N_15620,N_15595,N_15435);
xnor U15621 (N_15621,N_15223,N_15228);
nor U15622 (N_15622,N_15568,N_15327);
nor U15623 (N_15623,N_15201,N_15574);
nand U15624 (N_15624,N_15458,N_15234);
or U15625 (N_15625,N_15570,N_15409);
and U15626 (N_15626,N_15434,N_15364);
nand U15627 (N_15627,N_15260,N_15566);
nand U15628 (N_15628,N_15214,N_15529);
and U15629 (N_15629,N_15224,N_15239);
and U15630 (N_15630,N_15598,N_15455);
nand U15631 (N_15631,N_15386,N_15534);
nand U15632 (N_15632,N_15323,N_15488);
nand U15633 (N_15633,N_15545,N_15457);
nand U15634 (N_15634,N_15512,N_15352);
nand U15635 (N_15635,N_15205,N_15443);
and U15636 (N_15636,N_15450,N_15439);
or U15637 (N_15637,N_15313,N_15237);
or U15638 (N_15638,N_15451,N_15558);
nand U15639 (N_15639,N_15543,N_15348);
and U15640 (N_15640,N_15502,N_15479);
or U15641 (N_15641,N_15261,N_15221);
and U15642 (N_15642,N_15259,N_15249);
nor U15643 (N_15643,N_15572,N_15372);
and U15644 (N_15644,N_15393,N_15480);
nor U15645 (N_15645,N_15342,N_15490);
and U15646 (N_15646,N_15483,N_15252);
and U15647 (N_15647,N_15481,N_15404);
nor U15648 (N_15648,N_15509,N_15269);
or U15649 (N_15649,N_15402,N_15418);
nor U15650 (N_15650,N_15300,N_15245);
nand U15651 (N_15651,N_15307,N_15441);
nor U15652 (N_15652,N_15581,N_15485);
nand U15653 (N_15653,N_15553,N_15544);
nand U15654 (N_15654,N_15392,N_15338);
and U15655 (N_15655,N_15589,N_15403);
nor U15656 (N_15656,N_15329,N_15280);
and U15657 (N_15657,N_15408,N_15235);
or U15658 (N_15658,N_15288,N_15378);
nor U15659 (N_15659,N_15584,N_15586);
or U15660 (N_15660,N_15216,N_15384);
nor U15661 (N_15661,N_15561,N_15522);
nand U15662 (N_15662,N_15515,N_15444);
nor U15663 (N_15663,N_15231,N_15330);
nor U15664 (N_15664,N_15567,N_15463);
nor U15665 (N_15665,N_15311,N_15424);
nor U15666 (N_15666,N_15351,N_15286);
nor U15667 (N_15667,N_15346,N_15533);
nand U15668 (N_15668,N_15405,N_15263);
and U15669 (N_15669,N_15202,N_15347);
nand U15670 (N_15670,N_15316,N_15537);
nor U15671 (N_15671,N_15357,N_15208);
nor U15672 (N_15672,N_15301,N_15217);
nand U15673 (N_15673,N_15548,N_15218);
nor U15674 (N_15674,N_15555,N_15503);
nor U15675 (N_15675,N_15256,N_15505);
xnor U15676 (N_15676,N_15209,N_15410);
and U15677 (N_15677,N_15399,N_15588);
nor U15678 (N_15678,N_15491,N_15428);
or U15679 (N_15679,N_15356,N_15290);
and U15680 (N_15680,N_15577,N_15336);
or U15681 (N_15681,N_15229,N_15507);
or U15682 (N_15682,N_15226,N_15374);
or U15683 (N_15683,N_15486,N_15582);
nand U15684 (N_15684,N_15211,N_15268);
or U15685 (N_15685,N_15279,N_15487);
xnor U15686 (N_15686,N_15275,N_15213);
and U15687 (N_15687,N_15325,N_15292);
nor U15688 (N_15688,N_15244,N_15580);
and U15689 (N_15689,N_15412,N_15255);
nor U15690 (N_15690,N_15363,N_15546);
nor U15691 (N_15691,N_15369,N_15565);
nand U15692 (N_15692,N_15382,N_15390);
nand U15693 (N_15693,N_15344,N_15511);
and U15694 (N_15694,N_15508,N_15375);
or U15695 (N_15695,N_15227,N_15551);
nand U15696 (N_15696,N_15413,N_15321);
and U15697 (N_15697,N_15454,N_15383);
nor U15698 (N_15698,N_15556,N_15499);
nand U15699 (N_15699,N_15510,N_15562);
nand U15700 (N_15700,N_15563,N_15345);
nor U15701 (N_15701,N_15354,N_15471);
nand U15702 (N_15702,N_15587,N_15484);
nand U15703 (N_15703,N_15287,N_15477);
xor U15704 (N_15704,N_15339,N_15516);
or U15705 (N_15705,N_15319,N_15525);
and U15706 (N_15706,N_15225,N_15440);
and U15707 (N_15707,N_15519,N_15521);
and U15708 (N_15708,N_15297,N_15276);
or U15709 (N_15709,N_15539,N_15293);
and U15710 (N_15710,N_15258,N_15266);
or U15711 (N_15711,N_15219,N_15353);
nand U15712 (N_15712,N_15337,N_15314);
nor U15713 (N_15713,N_15554,N_15448);
and U15714 (N_15714,N_15267,N_15569);
nor U15715 (N_15715,N_15583,N_15236);
or U15716 (N_15716,N_15538,N_15447);
or U15717 (N_15717,N_15513,N_15366);
nand U15718 (N_15718,N_15482,N_15594);
or U15719 (N_15719,N_15419,N_15305);
nor U15720 (N_15720,N_15282,N_15349);
nor U15721 (N_15721,N_15426,N_15401);
and U15722 (N_15722,N_15417,N_15406);
xnor U15723 (N_15723,N_15355,N_15273);
nand U15724 (N_15724,N_15452,N_15571);
nand U15725 (N_15725,N_15462,N_15535);
or U15726 (N_15726,N_15497,N_15272);
and U15727 (N_15727,N_15230,N_15464);
nand U15728 (N_15728,N_15475,N_15359);
or U15729 (N_15729,N_15246,N_15453);
nor U15730 (N_15730,N_15527,N_15542);
or U15731 (N_15731,N_15328,N_15425);
nand U15732 (N_15732,N_15238,N_15493);
nor U15733 (N_15733,N_15389,N_15536);
nand U15734 (N_15734,N_15242,N_15492);
nor U15735 (N_15735,N_15550,N_15251);
and U15736 (N_15736,N_15552,N_15564);
and U15737 (N_15737,N_15310,N_15506);
or U15738 (N_15738,N_15304,N_15518);
nor U15739 (N_15739,N_15277,N_15540);
and U15740 (N_15740,N_15358,N_15391);
nor U15741 (N_15741,N_15470,N_15365);
nor U15742 (N_15742,N_15222,N_15442);
nor U15743 (N_15743,N_15247,N_15461);
nor U15744 (N_15744,N_15362,N_15296);
or U15745 (N_15745,N_15596,N_15233);
nor U15746 (N_15746,N_15591,N_15579);
and U15747 (N_15747,N_15590,N_15289);
nor U15748 (N_15748,N_15210,N_15432);
or U15749 (N_15749,N_15489,N_15332);
and U15750 (N_15750,N_15315,N_15308);
nand U15751 (N_15751,N_15379,N_15547);
and U15752 (N_15752,N_15560,N_15526);
nand U15753 (N_15753,N_15250,N_15531);
nand U15754 (N_15754,N_15472,N_15415);
nor U15755 (N_15755,N_15422,N_15253);
or U15756 (N_15756,N_15387,N_15215);
and U15757 (N_15757,N_15427,N_15320);
nor U15758 (N_15758,N_15593,N_15341);
and U15759 (N_15759,N_15438,N_15370);
nor U15760 (N_15760,N_15524,N_15326);
and U15761 (N_15761,N_15278,N_15431);
and U15762 (N_15762,N_15257,N_15517);
or U15763 (N_15763,N_15343,N_15557);
and U15764 (N_15764,N_15200,N_15285);
or U15765 (N_15765,N_15264,N_15420);
or U15766 (N_15766,N_15294,N_15576);
nand U15767 (N_15767,N_15318,N_15592);
nor U15768 (N_15768,N_15433,N_15270);
and U15769 (N_15769,N_15469,N_15437);
or U15770 (N_15770,N_15265,N_15232);
nor U15771 (N_15771,N_15436,N_15573);
or U15772 (N_15772,N_15254,N_15377);
or U15773 (N_15773,N_15274,N_15360);
and U15774 (N_15774,N_15465,N_15271);
nor U15775 (N_15775,N_15212,N_15203);
and U15776 (N_15776,N_15501,N_15549);
and U15777 (N_15777,N_15306,N_15373);
nand U15778 (N_15778,N_15500,N_15206);
nand U15779 (N_15779,N_15532,N_15394);
and U15780 (N_15780,N_15504,N_15388);
and U15781 (N_15781,N_15523,N_15520);
and U15782 (N_15782,N_15281,N_15414);
nor U15783 (N_15783,N_15528,N_15468);
nor U15784 (N_15784,N_15578,N_15299);
nor U15785 (N_15785,N_15340,N_15396);
nor U15786 (N_15786,N_15380,N_15298);
nand U15787 (N_15787,N_15381,N_15476);
or U15788 (N_15788,N_15597,N_15498);
nand U15789 (N_15789,N_15291,N_15398);
nor U15790 (N_15790,N_15459,N_15430);
or U15791 (N_15791,N_15333,N_15317);
and U15792 (N_15792,N_15284,N_15303);
and U15793 (N_15793,N_15449,N_15220);
nor U15794 (N_15794,N_15368,N_15331);
or U15795 (N_15795,N_15322,N_15474);
nand U15796 (N_15796,N_15312,N_15478);
nand U15797 (N_15797,N_15397,N_15240);
nor U15798 (N_15798,N_15395,N_15400);
xnor U15799 (N_15799,N_15495,N_15350);
or U15800 (N_15800,N_15485,N_15489);
nand U15801 (N_15801,N_15389,N_15237);
or U15802 (N_15802,N_15252,N_15382);
and U15803 (N_15803,N_15596,N_15446);
nand U15804 (N_15804,N_15551,N_15406);
nand U15805 (N_15805,N_15556,N_15219);
nand U15806 (N_15806,N_15456,N_15329);
nand U15807 (N_15807,N_15441,N_15241);
nor U15808 (N_15808,N_15488,N_15351);
and U15809 (N_15809,N_15513,N_15294);
or U15810 (N_15810,N_15478,N_15364);
and U15811 (N_15811,N_15204,N_15372);
nand U15812 (N_15812,N_15422,N_15366);
nand U15813 (N_15813,N_15465,N_15315);
or U15814 (N_15814,N_15446,N_15384);
nand U15815 (N_15815,N_15444,N_15485);
nand U15816 (N_15816,N_15372,N_15298);
nor U15817 (N_15817,N_15315,N_15346);
or U15818 (N_15818,N_15297,N_15235);
and U15819 (N_15819,N_15586,N_15267);
nor U15820 (N_15820,N_15210,N_15362);
and U15821 (N_15821,N_15297,N_15532);
and U15822 (N_15822,N_15467,N_15205);
nand U15823 (N_15823,N_15404,N_15362);
or U15824 (N_15824,N_15419,N_15301);
and U15825 (N_15825,N_15495,N_15255);
nor U15826 (N_15826,N_15337,N_15510);
or U15827 (N_15827,N_15320,N_15339);
or U15828 (N_15828,N_15320,N_15480);
or U15829 (N_15829,N_15479,N_15572);
nor U15830 (N_15830,N_15380,N_15502);
nand U15831 (N_15831,N_15505,N_15361);
nor U15832 (N_15832,N_15523,N_15472);
nand U15833 (N_15833,N_15552,N_15548);
nand U15834 (N_15834,N_15423,N_15452);
and U15835 (N_15835,N_15478,N_15218);
nor U15836 (N_15836,N_15312,N_15421);
nor U15837 (N_15837,N_15359,N_15422);
nand U15838 (N_15838,N_15581,N_15451);
or U15839 (N_15839,N_15508,N_15301);
and U15840 (N_15840,N_15356,N_15474);
xnor U15841 (N_15841,N_15583,N_15506);
and U15842 (N_15842,N_15468,N_15332);
nand U15843 (N_15843,N_15599,N_15521);
nor U15844 (N_15844,N_15295,N_15470);
and U15845 (N_15845,N_15503,N_15262);
and U15846 (N_15846,N_15586,N_15555);
nand U15847 (N_15847,N_15513,N_15563);
nand U15848 (N_15848,N_15515,N_15359);
or U15849 (N_15849,N_15304,N_15447);
nand U15850 (N_15850,N_15328,N_15325);
nand U15851 (N_15851,N_15560,N_15328);
nand U15852 (N_15852,N_15214,N_15555);
nor U15853 (N_15853,N_15321,N_15275);
nor U15854 (N_15854,N_15419,N_15307);
nand U15855 (N_15855,N_15342,N_15209);
or U15856 (N_15856,N_15569,N_15572);
and U15857 (N_15857,N_15210,N_15563);
nor U15858 (N_15858,N_15537,N_15224);
and U15859 (N_15859,N_15354,N_15405);
or U15860 (N_15860,N_15544,N_15522);
nor U15861 (N_15861,N_15524,N_15246);
nand U15862 (N_15862,N_15272,N_15440);
nand U15863 (N_15863,N_15328,N_15307);
nor U15864 (N_15864,N_15256,N_15257);
and U15865 (N_15865,N_15355,N_15306);
nand U15866 (N_15866,N_15403,N_15431);
or U15867 (N_15867,N_15269,N_15577);
nand U15868 (N_15868,N_15375,N_15293);
nor U15869 (N_15869,N_15432,N_15248);
and U15870 (N_15870,N_15497,N_15540);
or U15871 (N_15871,N_15530,N_15592);
nor U15872 (N_15872,N_15339,N_15315);
nand U15873 (N_15873,N_15579,N_15544);
nand U15874 (N_15874,N_15578,N_15300);
and U15875 (N_15875,N_15429,N_15543);
or U15876 (N_15876,N_15414,N_15412);
and U15877 (N_15877,N_15580,N_15231);
or U15878 (N_15878,N_15561,N_15421);
or U15879 (N_15879,N_15570,N_15371);
or U15880 (N_15880,N_15505,N_15492);
nor U15881 (N_15881,N_15364,N_15333);
or U15882 (N_15882,N_15581,N_15421);
and U15883 (N_15883,N_15364,N_15428);
or U15884 (N_15884,N_15533,N_15271);
nand U15885 (N_15885,N_15281,N_15253);
or U15886 (N_15886,N_15588,N_15381);
or U15887 (N_15887,N_15351,N_15382);
nand U15888 (N_15888,N_15538,N_15315);
nand U15889 (N_15889,N_15291,N_15568);
nor U15890 (N_15890,N_15378,N_15535);
or U15891 (N_15891,N_15304,N_15399);
nand U15892 (N_15892,N_15242,N_15267);
nand U15893 (N_15893,N_15408,N_15312);
or U15894 (N_15894,N_15289,N_15313);
or U15895 (N_15895,N_15244,N_15390);
nand U15896 (N_15896,N_15311,N_15277);
and U15897 (N_15897,N_15558,N_15260);
nand U15898 (N_15898,N_15396,N_15538);
and U15899 (N_15899,N_15456,N_15535);
nand U15900 (N_15900,N_15466,N_15471);
nand U15901 (N_15901,N_15253,N_15271);
nor U15902 (N_15902,N_15355,N_15559);
or U15903 (N_15903,N_15588,N_15425);
or U15904 (N_15904,N_15518,N_15575);
nor U15905 (N_15905,N_15486,N_15363);
and U15906 (N_15906,N_15530,N_15224);
nor U15907 (N_15907,N_15280,N_15452);
or U15908 (N_15908,N_15256,N_15495);
nor U15909 (N_15909,N_15223,N_15458);
or U15910 (N_15910,N_15302,N_15365);
nand U15911 (N_15911,N_15238,N_15598);
nor U15912 (N_15912,N_15514,N_15271);
nand U15913 (N_15913,N_15295,N_15460);
and U15914 (N_15914,N_15503,N_15352);
nor U15915 (N_15915,N_15278,N_15465);
nor U15916 (N_15916,N_15433,N_15366);
or U15917 (N_15917,N_15317,N_15479);
nand U15918 (N_15918,N_15599,N_15382);
nand U15919 (N_15919,N_15455,N_15349);
nor U15920 (N_15920,N_15401,N_15451);
and U15921 (N_15921,N_15253,N_15532);
nor U15922 (N_15922,N_15218,N_15266);
nand U15923 (N_15923,N_15256,N_15278);
nand U15924 (N_15924,N_15504,N_15424);
nor U15925 (N_15925,N_15530,N_15463);
and U15926 (N_15926,N_15553,N_15479);
nand U15927 (N_15927,N_15349,N_15229);
or U15928 (N_15928,N_15281,N_15369);
and U15929 (N_15929,N_15523,N_15373);
or U15930 (N_15930,N_15397,N_15416);
nand U15931 (N_15931,N_15388,N_15557);
or U15932 (N_15932,N_15486,N_15326);
and U15933 (N_15933,N_15567,N_15231);
and U15934 (N_15934,N_15547,N_15375);
and U15935 (N_15935,N_15529,N_15224);
and U15936 (N_15936,N_15350,N_15593);
and U15937 (N_15937,N_15368,N_15205);
nor U15938 (N_15938,N_15343,N_15477);
or U15939 (N_15939,N_15576,N_15375);
nor U15940 (N_15940,N_15377,N_15553);
nand U15941 (N_15941,N_15251,N_15331);
nand U15942 (N_15942,N_15319,N_15418);
nand U15943 (N_15943,N_15517,N_15378);
and U15944 (N_15944,N_15236,N_15560);
nand U15945 (N_15945,N_15400,N_15313);
and U15946 (N_15946,N_15460,N_15287);
nand U15947 (N_15947,N_15320,N_15550);
or U15948 (N_15948,N_15280,N_15332);
nor U15949 (N_15949,N_15258,N_15253);
nor U15950 (N_15950,N_15207,N_15378);
and U15951 (N_15951,N_15264,N_15316);
nand U15952 (N_15952,N_15598,N_15492);
nor U15953 (N_15953,N_15218,N_15394);
or U15954 (N_15954,N_15582,N_15502);
nor U15955 (N_15955,N_15524,N_15492);
and U15956 (N_15956,N_15348,N_15589);
nand U15957 (N_15957,N_15266,N_15574);
or U15958 (N_15958,N_15599,N_15296);
and U15959 (N_15959,N_15434,N_15282);
and U15960 (N_15960,N_15593,N_15499);
and U15961 (N_15961,N_15545,N_15517);
nand U15962 (N_15962,N_15379,N_15208);
or U15963 (N_15963,N_15454,N_15306);
or U15964 (N_15964,N_15291,N_15373);
nor U15965 (N_15965,N_15545,N_15376);
and U15966 (N_15966,N_15398,N_15325);
or U15967 (N_15967,N_15208,N_15498);
nor U15968 (N_15968,N_15242,N_15539);
and U15969 (N_15969,N_15432,N_15369);
or U15970 (N_15970,N_15595,N_15221);
and U15971 (N_15971,N_15286,N_15220);
or U15972 (N_15972,N_15317,N_15222);
and U15973 (N_15973,N_15427,N_15583);
nand U15974 (N_15974,N_15435,N_15278);
or U15975 (N_15975,N_15574,N_15332);
xnor U15976 (N_15976,N_15353,N_15554);
nor U15977 (N_15977,N_15557,N_15471);
nor U15978 (N_15978,N_15382,N_15212);
and U15979 (N_15979,N_15264,N_15516);
or U15980 (N_15980,N_15472,N_15243);
nor U15981 (N_15981,N_15582,N_15480);
and U15982 (N_15982,N_15483,N_15278);
and U15983 (N_15983,N_15256,N_15425);
and U15984 (N_15984,N_15469,N_15548);
and U15985 (N_15985,N_15237,N_15445);
or U15986 (N_15986,N_15238,N_15223);
or U15987 (N_15987,N_15244,N_15449);
or U15988 (N_15988,N_15477,N_15321);
and U15989 (N_15989,N_15224,N_15295);
nor U15990 (N_15990,N_15587,N_15227);
nor U15991 (N_15991,N_15547,N_15236);
and U15992 (N_15992,N_15223,N_15251);
and U15993 (N_15993,N_15202,N_15599);
and U15994 (N_15994,N_15335,N_15204);
nor U15995 (N_15995,N_15277,N_15547);
or U15996 (N_15996,N_15490,N_15228);
or U15997 (N_15997,N_15554,N_15384);
nand U15998 (N_15998,N_15321,N_15501);
and U15999 (N_15999,N_15518,N_15478);
nor U16000 (N_16000,N_15763,N_15841);
and U16001 (N_16001,N_15886,N_15725);
or U16002 (N_16002,N_15993,N_15897);
and U16003 (N_16003,N_15867,N_15907);
and U16004 (N_16004,N_15929,N_15925);
nand U16005 (N_16005,N_15856,N_15739);
and U16006 (N_16006,N_15774,N_15979);
and U16007 (N_16007,N_15687,N_15716);
and U16008 (N_16008,N_15669,N_15985);
and U16009 (N_16009,N_15924,N_15640);
or U16010 (N_16010,N_15805,N_15996);
and U16011 (N_16011,N_15697,N_15641);
and U16012 (N_16012,N_15633,N_15876);
or U16013 (N_16013,N_15807,N_15631);
nor U16014 (N_16014,N_15730,N_15748);
nand U16015 (N_16015,N_15652,N_15817);
and U16016 (N_16016,N_15982,N_15840);
and U16017 (N_16017,N_15857,N_15622);
and U16018 (N_16018,N_15849,N_15971);
nor U16019 (N_16019,N_15789,N_15884);
or U16020 (N_16020,N_15923,N_15629);
nand U16021 (N_16021,N_15727,N_15664);
nor U16022 (N_16022,N_15920,N_15607);
nor U16023 (N_16023,N_15699,N_15831);
or U16024 (N_16024,N_15832,N_15936);
or U16025 (N_16025,N_15975,N_15987);
nand U16026 (N_16026,N_15863,N_15812);
nand U16027 (N_16027,N_15684,N_15811);
or U16028 (N_16028,N_15715,N_15645);
and U16029 (N_16029,N_15802,N_15881);
or U16030 (N_16030,N_15628,N_15646);
nor U16031 (N_16031,N_15617,N_15708);
nand U16032 (N_16032,N_15816,N_15778);
nor U16033 (N_16033,N_15665,N_15614);
and U16034 (N_16034,N_15958,N_15685);
and U16035 (N_16035,N_15660,N_15951);
or U16036 (N_16036,N_15911,N_15829);
or U16037 (N_16037,N_15972,N_15657);
nor U16038 (N_16038,N_15843,N_15906);
nand U16039 (N_16039,N_15775,N_15674);
and U16040 (N_16040,N_15813,N_15711);
nor U16041 (N_16041,N_15950,N_15980);
and U16042 (N_16042,N_15720,N_15922);
nand U16043 (N_16043,N_15943,N_15693);
and U16044 (N_16044,N_15648,N_15865);
nor U16045 (N_16045,N_15998,N_15825);
and U16046 (N_16046,N_15990,N_15937);
nor U16047 (N_16047,N_15689,N_15655);
and U16048 (N_16048,N_15605,N_15848);
or U16049 (N_16049,N_15932,N_15814);
nor U16050 (N_16050,N_15735,N_15823);
nor U16051 (N_16051,N_15838,N_15928);
nor U16052 (N_16052,N_15703,N_15624);
or U16053 (N_16053,N_15760,N_15673);
nor U16054 (N_16054,N_15626,N_15706);
nand U16055 (N_16055,N_15968,N_15681);
nand U16056 (N_16056,N_15724,N_15839);
nor U16057 (N_16057,N_15926,N_15959);
nor U16058 (N_16058,N_15644,N_15885);
and U16059 (N_16059,N_15634,N_15905);
nand U16060 (N_16060,N_15873,N_15948);
nand U16061 (N_16061,N_15903,N_15977);
nand U16062 (N_16062,N_15757,N_15714);
nand U16063 (N_16063,N_15773,N_15654);
nor U16064 (N_16064,N_15868,N_15771);
and U16065 (N_16065,N_15870,N_15653);
and U16066 (N_16066,N_15675,N_15686);
and U16067 (N_16067,N_15600,N_15967);
nor U16068 (N_16068,N_15667,N_15830);
nor U16069 (N_16069,N_15759,N_15747);
nor U16070 (N_16070,N_15846,N_15888);
and U16071 (N_16071,N_15670,N_15909);
nor U16072 (N_16072,N_15808,N_15688);
and U16073 (N_16073,N_15637,N_15939);
or U16074 (N_16074,N_15707,N_15934);
or U16075 (N_16075,N_15753,N_15734);
and U16076 (N_16076,N_15676,N_15916);
or U16077 (N_16077,N_15917,N_15726);
nand U16078 (N_16078,N_15938,N_15851);
or U16079 (N_16079,N_15866,N_15902);
nor U16080 (N_16080,N_15784,N_15709);
nand U16081 (N_16081,N_15954,N_15860);
and U16082 (N_16082,N_15842,N_15723);
or U16083 (N_16083,N_15690,N_15961);
nor U16084 (N_16084,N_15649,N_15986);
or U16085 (N_16085,N_15780,N_15898);
and U16086 (N_16086,N_15671,N_15651);
nor U16087 (N_16087,N_15820,N_15696);
and U16088 (N_16088,N_15701,N_15764);
or U16089 (N_16089,N_15755,N_15683);
and U16090 (N_16090,N_15650,N_15766);
xor U16091 (N_16091,N_15722,N_15768);
xor U16092 (N_16092,N_15758,N_15694);
and U16093 (N_16093,N_15835,N_15964);
nand U16094 (N_16094,N_15658,N_15601);
nor U16095 (N_16095,N_15892,N_15705);
nor U16096 (N_16096,N_15604,N_15619);
and U16097 (N_16097,N_15743,N_15765);
or U16098 (N_16098,N_15988,N_15792);
or U16099 (N_16099,N_15862,N_15719);
and U16100 (N_16100,N_15608,N_15620);
or U16101 (N_16101,N_15994,N_15798);
or U16102 (N_16102,N_15736,N_15603);
nand U16103 (N_16103,N_15744,N_15894);
and U16104 (N_16104,N_15962,N_15844);
or U16105 (N_16105,N_15899,N_15983);
nor U16106 (N_16106,N_15908,N_15733);
or U16107 (N_16107,N_15606,N_15826);
nand U16108 (N_16108,N_15615,N_15946);
or U16109 (N_16109,N_15956,N_15861);
or U16110 (N_16110,N_15636,N_15761);
nor U16111 (N_16111,N_15869,N_15901);
or U16112 (N_16112,N_15957,N_15799);
or U16113 (N_16113,N_15889,N_15737);
nor U16114 (N_16114,N_15610,N_15661);
or U16115 (N_16115,N_15700,N_15879);
nor U16116 (N_16116,N_15679,N_15837);
nor U16117 (N_16117,N_15772,N_15893);
nor U16118 (N_16118,N_15989,N_15965);
nand U16119 (N_16119,N_15795,N_15611);
or U16120 (N_16120,N_15895,N_15969);
nand U16121 (N_16121,N_15625,N_15793);
nand U16122 (N_16122,N_15896,N_15621);
and U16123 (N_16123,N_15790,N_15921);
xnor U16124 (N_16124,N_15941,N_15995);
and U16125 (N_16125,N_15970,N_15642);
nor U16126 (N_16126,N_15635,N_15692);
and U16127 (N_16127,N_15992,N_15791);
nand U16128 (N_16128,N_15878,N_15618);
and U16129 (N_16129,N_15682,N_15632);
and U16130 (N_16130,N_15663,N_15949);
or U16131 (N_16131,N_15984,N_15827);
nor U16132 (N_16132,N_15847,N_15877);
nor U16133 (N_16133,N_15738,N_15776);
and U16134 (N_16134,N_15915,N_15821);
and U16135 (N_16135,N_15721,N_15769);
and U16136 (N_16136,N_15746,N_15612);
nand U16137 (N_16137,N_15656,N_15945);
or U16138 (N_16138,N_15672,N_15749);
nand U16139 (N_16139,N_15627,N_15616);
and U16140 (N_16140,N_15850,N_15787);
nand U16141 (N_16141,N_15864,N_15872);
nor U16142 (N_16142,N_15854,N_15930);
nor U16143 (N_16143,N_15940,N_15741);
or U16144 (N_16144,N_15942,N_15858);
nand U16145 (N_16145,N_15639,N_15638);
or U16146 (N_16146,N_15777,N_15887);
xor U16147 (N_16147,N_15800,N_15918);
nor U16148 (N_16148,N_15732,N_15974);
nor U16149 (N_16149,N_15677,N_15852);
nor U16150 (N_16150,N_15698,N_15904);
xor U16151 (N_16151,N_15643,N_15781);
nor U16152 (N_16152,N_15810,N_15731);
and U16153 (N_16153,N_15953,N_15871);
nor U16154 (N_16154,N_15824,N_15678);
nor U16155 (N_16155,N_15728,N_15931);
nor U16156 (N_16156,N_15900,N_15783);
or U16157 (N_16157,N_15702,N_15796);
nor U16158 (N_16158,N_15713,N_15752);
or U16159 (N_16159,N_15712,N_15801);
nor U16160 (N_16160,N_15828,N_15815);
nand U16161 (N_16161,N_15999,N_15819);
or U16162 (N_16162,N_15740,N_15797);
or U16163 (N_16163,N_15874,N_15880);
or U16164 (N_16164,N_15630,N_15859);
nor U16165 (N_16165,N_15704,N_15890);
or U16166 (N_16166,N_15602,N_15834);
or U16167 (N_16167,N_15845,N_15875);
nor U16168 (N_16168,N_15767,N_15933);
or U16169 (N_16169,N_15717,N_15853);
or U16170 (N_16170,N_15891,N_15609);
and U16171 (N_16171,N_15912,N_15751);
or U16172 (N_16172,N_15822,N_15788);
nor U16173 (N_16173,N_15613,N_15659);
nand U16174 (N_16174,N_15779,N_15770);
nor U16175 (N_16175,N_15960,N_15978);
nor U16176 (N_16176,N_15680,N_15750);
and U16177 (N_16177,N_15785,N_15662);
or U16178 (N_16178,N_15833,N_15809);
or U16179 (N_16179,N_15745,N_15910);
or U16180 (N_16180,N_15666,N_15976);
and U16181 (N_16181,N_15804,N_15710);
and U16182 (N_16182,N_15973,N_15955);
and U16183 (N_16183,N_15818,N_15794);
or U16184 (N_16184,N_15782,N_15691);
or U16185 (N_16185,N_15668,N_15997);
or U16186 (N_16186,N_15695,N_15913);
or U16187 (N_16187,N_15718,N_15981);
nand U16188 (N_16188,N_15729,N_15952);
and U16189 (N_16189,N_15762,N_15963);
nand U16190 (N_16190,N_15927,N_15883);
nand U16191 (N_16191,N_15623,N_15966);
nor U16192 (N_16192,N_15803,N_15914);
or U16193 (N_16193,N_15944,N_15991);
and U16194 (N_16194,N_15855,N_15919);
or U16195 (N_16195,N_15756,N_15935);
nor U16196 (N_16196,N_15754,N_15742);
and U16197 (N_16197,N_15806,N_15836);
and U16198 (N_16198,N_15947,N_15882);
or U16199 (N_16199,N_15786,N_15647);
or U16200 (N_16200,N_15709,N_15704);
nand U16201 (N_16201,N_15652,N_15852);
and U16202 (N_16202,N_15902,N_15933);
nor U16203 (N_16203,N_15921,N_15696);
and U16204 (N_16204,N_15733,N_15915);
nand U16205 (N_16205,N_15841,N_15772);
nor U16206 (N_16206,N_15914,N_15969);
nand U16207 (N_16207,N_15993,N_15750);
nand U16208 (N_16208,N_15792,N_15677);
nor U16209 (N_16209,N_15879,N_15661);
nand U16210 (N_16210,N_15924,N_15651);
nor U16211 (N_16211,N_15839,N_15675);
or U16212 (N_16212,N_15971,N_15744);
or U16213 (N_16213,N_15632,N_15916);
nand U16214 (N_16214,N_15742,N_15906);
and U16215 (N_16215,N_15892,N_15688);
nor U16216 (N_16216,N_15669,N_15863);
nand U16217 (N_16217,N_15846,N_15936);
nand U16218 (N_16218,N_15726,N_15659);
nand U16219 (N_16219,N_15861,N_15828);
nand U16220 (N_16220,N_15823,N_15916);
or U16221 (N_16221,N_15649,N_15758);
nor U16222 (N_16222,N_15904,N_15814);
nand U16223 (N_16223,N_15833,N_15871);
or U16224 (N_16224,N_15915,N_15852);
nand U16225 (N_16225,N_15731,N_15985);
nand U16226 (N_16226,N_15745,N_15679);
or U16227 (N_16227,N_15804,N_15719);
and U16228 (N_16228,N_15651,N_15913);
and U16229 (N_16229,N_15630,N_15647);
nor U16230 (N_16230,N_15664,N_15882);
nor U16231 (N_16231,N_15948,N_15724);
nand U16232 (N_16232,N_15660,N_15821);
nand U16233 (N_16233,N_15626,N_15817);
nor U16234 (N_16234,N_15872,N_15648);
and U16235 (N_16235,N_15758,N_15772);
or U16236 (N_16236,N_15688,N_15846);
and U16237 (N_16237,N_15734,N_15771);
and U16238 (N_16238,N_15870,N_15623);
or U16239 (N_16239,N_15735,N_15955);
xor U16240 (N_16240,N_15695,N_15772);
nor U16241 (N_16241,N_15815,N_15865);
nor U16242 (N_16242,N_15909,N_15698);
xor U16243 (N_16243,N_15696,N_15841);
nand U16244 (N_16244,N_15769,N_15609);
nor U16245 (N_16245,N_15687,N_15740);
nand U16246 (N_16246,N_15843,N_15817);
or U16247 (N_16247,N_15653,N_15656);
nand U16248 (N_16248,N_15955,N_15794);
nand U16249 (N_16249,N_15899,N_15914);
or U16250 (N_16250,N_15894,N_15925);
nor U16251 (N_16251,N_15640,N_15622);
or U16252 (N_16252,N_15682,N_15962);
nor U16253 (N_16253,N_15720,N_15864);
and U16254 (N_16254,N_15775,N_15665);
and U16255 (N_16255,N_15827,N_15705);
nand U16256 (N_16256,N_15852,N_15786);
or U16257 (N_16257,N_15926,N_15832);
xnor U16258 (N_16258,N_15717,N_15686);
nor U16259 (N_16259,N_15830,N_15860);
nand U16260 (N_16260,N_15613,N_15806);
and U16261 (N_16261,N_15772,N_15686);
or U16262 (N_16262,N_15712,N_15880);
or U16263 (N_16263,N_15759,N_15929);
or U16264 (N_16264,N_15976,N_15833);
nor U16265 (N_16265,N_15812,N_15852);
nand U16266 (N_16266,N_15741,N_15962);
or U16267 (N_16267,N_15647,N_15950);
nor U16268 (N_16268,N_15894,N_15765);
nand U16269 (N_16269,N_15872,N_15669);
or U16270 (N_16270,N_15742,N_15827);
nor U16271 (N_16271,N_15761,N_15609);
nand U16272 (N_16272,N_15813,N_15759);
nor U16273 (N_16273,N_15632,N_15828);
or U16274 (N_16274,N_15623,N_15866);
and U16275 (N_16275,N_15933,N_15728);
or U16276 (N_16276,N_15620,N_15938);
nand U16277 (N_16277,N_15992,N_15740);
nor U16278 (N_16278,N_15950,N_15848);
or U16279 (N_16279,N_15803,N_15792);
and U16280 (N_16280,N_15981,N_15845);
and U16281 (N_16281,N_15911,N_15888);
or U16282 (N_16282,N_15762,N_15719);
and U16283 (N_16283,N_15747,N_15750);
or U16284 (N_16284,N_15870,N_15929);
nor U16285 (N_16285,N_15891,N_15921);
or U16286 (N_16286,N_15940,N_15745);
and U16287 (N_16287,N_15741,N_15810);
or U16288 (N_16288,N_15634,N_15886);
or U16289 (N_16289,N_15909,N_15933);
xor U16290 (N_16290,N_15786,N_15893);
and U16291 (N_16291,N_15776,N_15924);
and U16292 (N_16292,N_15876,N_15753);
or U16293 (N_16293,N_15757,N_15694);
and U16294 (N_16294,N_15986,N_15965);
and U16295 (N_16295,N_15605,N_15648);
nor U16296 (N_16296,N_15931,N_15916);
nor U16297 (N_16297,N_15616,N_15953);
nor U16298 (N_16298,N_15651,N_15818);
nand U16299 (N_16299,N_15922,N_15612);
nor U16300 (N_16300,N_15843,N_15800);
nor U16301 (N_16301,N_15831,N_15647);
and U16302 (N_16302,N_15819,N_15646);
and U16303 (N_16303,N_15857,N_15618);
nand U16304 (N_16304,N_15716,N_15702);
nand U16305 (N_16305,N_15738,N_15944);
nor U16306 (N_16306,N_15614,N_15948);
xnor U16307 (N_16307,N_15863,N_15679);
and U16308 (N_16308,N_15842,N_15674);
nor U16309 (N_16309,N_15785,N_15864);
nor U16310 (N_16310,N_15708,N_15997);
nor U16311 (N_16311,N_15736,N_15683);
and U16312 (N_16312,N_15879,N_15849);
nand U16313 (N_16313,N_15906,N_15834);
or U16314 (N_16314,N_15953,N_15918);
nor U16315 (N_16315,N_15841,N_15721);
and U16316 (N_16316,N_15737,N_15948);
nor U16317 (N_16317,N_15820,N_15817);
nor U16318 (N_16318,N_15623,N_15815);
and U16319 (N_16319,N_15650,N_15623);
nand U16320 (N_16320,N_15722,N_15950);
or U16321 (N_16321,N_15925,N_15835);
or U16322 (N_16322,N_15848,N_15925);
nand U16323 (N_16323,N_15676,N_15638);
nor U16324 (N_16324,N_15808,N_15950);
and U16325 (N_16325,N_15865,N_15716);
or U16326 (N_16326,N_15698,N_15873);
nor U16327 (N_16327,N_15857,N_15802);
nand U16328 (N_16328,N_15889,N_15728);
nor U16329 (N_16329,N_15855,N_15802);
or U16330 (N_16330,N_15828,N_15930);
nand U16331 (N_16331,N_15927,N_15740);
or U16332 (N_16332,N_15867,N_15861);
nand U16333 (N_16333,N_15735,N_15716);
and U16334 (N_16334,N_15760,N_15946);
nand U16335 (N_16335,N_15755,N_15719);
and U16336 (N_16336,N_15715,N_15697);
nor U16337 (N_16337,N_15952,N_15794);
or U16338 (N_16338,N_15950,N_15771);
nand U16339 (N_16339,N_15834,N_15664);
and U16340 (N_16340,N_15730,N_15631);
nor U16341 (N_16341,N_15786,N_15869);
nand U16342 (N_16342,N_15761,N_15831);
nand U16343 (N_16343,N_15769,N_15915);
nand U16344 (N_16344,N_15631,N_15798);
nor U16345 (N_16345,N_15730,N_15998);
nand U16346 (N_16346,N_15816,N_15827);
nand U16347 (N_16347,N_15647,N_15690);
nor U16348 (N_16348,N_15629,N_15614);
nand U16349 (N_16349,N_15801,N_15858);
nor U16350 (N_16350,N_15696,N_15946);
or U16351 (N_16351,N_15888,N_15832);
nor U16352 (N_16352,N_15853,N_15743);
nor U16353 (N_16353,N_15733,N_15787);
or U16354 (N_16354,N_15687,N_15739);
nand U16355 (N_16355,N_15624,N_15792);
and U16356 (N_16356,N_15943,N_15833);
nor U16357 (N_16357,N_15611,N_15750);
nand U16358 (N_16358,N_15937,N_15655);
and U16359 (N_16359,N_15923,N_15958);
nor U16360 (N_16360,N_15929,N_15672);
nand U16361 (N_16361,N_15789,N_15762);
or U16362 (N_16362,N_15841,N_15995);
nand U16363 (N_16363,N_15662,N_15879);
nand U16364 (N_16364,N_15721,N_15982);
nand U16365 (N_16365,N_15777,N_15799);
nand U16366 (N_16366,N_15758,N_15678);
or U16367 (N_16367,N_15895,N_15612);
nor U16368 (N_16368,N_15640,N_15651);
nand U16369 (N_16369,N_15688,N_15638);
nor U16370 (N_16370,N_15800,N_15730);
and U16371 (N_16371,N_15869,N_15824);
nand U16372 (N_16372,N_15949,N_15840);
and U16373 (N_16373,N_15986,N_15610);
nand U16374 (N_16374,N_15976,N_15746);
or U16375 (N_16375,N_15879,N_15965);
nor U16376 (N_16376,N_15656,N_15965);
or U16377 (N_16377,N_15959,N_15668);
and U16378 (N_16378,N_15686,N_15770);
or U16379 (N_16379,N_15662,N_15709);
nor U16380 (N_16380,N_15837,N_15778);
or U16381 (N_16381,N_15865,N_15600);
or U16382 (N_16382,N_15621,N_15760);
nor U16383 (N_16383,N_15801,N_15674);
or U16384 (N_16384,N_15662,N_15839);
and U16385 (N_16385,N_15791,N_15824);
nand U16386 (N_16386,N_15747,N_15907);
or U16387 (N_16387,N_15717,N_15910);
and U16388 (N_16388,N_15669,N_15836);
nand U16389 (N_16389,N_15614,N_15719);
and U16390 (N_16390,N_15655,N_15972);
and U16391 (N_16391,N_15787,N_15915);
and U16392 (N_16392,N_15884,N_15826);
nand U16393 (N_16393,N_15943,N_15617);
nor U16394 (N_16394,N_15724,N_15661);
nand U16395 (N_16395,N_15622,N_15652);
or U16396 (N_16396,N_15805,N_15678);
nor U16397 (N_16397,N_15620,N_15684);
and U16398 (N_16398,N_15653,N_15991);
nor U16399 (N_16399,N_15706,N_15836);
nor U16400 (N_16400,N_16012,N_16039);
and U16401 (N_16401,N_16303,N_16097);
nand U16402 (N_16402,N_16105,N_16094);
and U16403 (N_16403,N_16369,N_16395);
nand U16404 (N_16404,N_16175,N_16291);
nand U16405 (N_16405,N_16252,N_16214);
or U16406 (N_16406,N_16196,N_16030);
nor U16407 (N_16407,N_16298,N_16217);
and U16408 (N_16408,N_16006,N_16248);
and U16409 (N_16409,N_16100,N_16269);
and U16410 (N_16410,N_16378,N_16087);
nor U16411 (N_16411,N_16274,N_16372);
nand U16412 (N_16412,N_16076,N_16180);
or U16413 (N_16413,N_16223,N_16146);
nor U16414 (N_16414,N_16238,N_16268);
nand U16415 (N_16415,N_16185,N_16201);
nand U16416 (N_16416,N_16163,N_16153);
or U16417 (N_16417,N_16391,N_16392);
and U16418 (N_16418,N_16042,N_16074);
nand U16419 (N_16419,N_16330,N_16229);
and U16420 (N_16420,N_16383,N_16237);
or U16421 (N_16421,N_16243,N_16205);
nand U16422 (N_16422,N_16216,N_16352);
or U16423 (N_16423,N_16353,N_16145);
and U16424 (N_16424,N_16359,N_16317);
nand U16425 (N_16425,N_16056,N_16133);
or U16426 (N_16426,N_16040,N_16013);
and U16427 (N_16427,N_16092,N_16150);
nand U16428 (N_16428,N_16376,N_16308);
or U16429 (N_16429,N_16025,N_16109);
nor U16430 (N_16430,N_16335,N_16301);
or U16431 (N_16431,N_16231,N_16351);
nor U16432 (N_16432,N_16363,N_16050);
or U16433 (N_16433,N_16136,N_16388);
nor U16434 (N_16434,N_16350,N_16270);
nand U16435 (N_16435,N_16179,N_16354);
and U16436 (N_16436,N_16021,N_16202);
or U16437 (N_16437,N_16278,N_16059);
and U16438 (N_16438,N_16336,N_16297);
and U16439 (N_16439,N_16287,N_16296);
and U16440 (N_16440,N_16257,N_16347);
and U16441 (N_16441,N_16272,N_16055);
nand U16442 (N_16442,N_16325,N_16144);
nor U16443 (N_16443,N_16398,N_16151);
or U16444 (N_16444,N_16079,N_16188);
or U16445 (N_16445,N_16191,N_16022);
nor U16446 (N_16446,N_16183,N_16159);
nand U16447 (N_16447,N_16187,N_16311);
nor U16448 (N_16448,N_16096,N_16137);
or U16449 (N_16449,N_16121,N_16209);
nand U16450 (N_16450,N_16332,N_16210);
xnor U16451 (N_16451,N_16104,N_16259);
nor U16452 (N_16452,N_16043,N_16171);
or U16453 (N_16453,N_16091,N_16095);
or U16454 (N_16454,N_16283,N_16184);
nand U16455 (N_16455,N_16067,N_16240);
and U16456 (N_16456,N_16305,N_16318);
and U16457 (N_16457,N_16256,N_16307);
nor U16458 (N_16458,N_16023,N_16235);
nor U16459 (N_16459,N_16340,N_16176);
nand U16460 (N_16460,N_16134,N_16054);
and U16461 (N_16461,N_16062,N_16281);
or U16462 (N_16462,N_16027,N_16379);
nor U16463 (N_16463,N_16186,N_16098);
and U16464 (N_16464,N_16199,N_16182);
nor U16465 (N_16465,N_16010,N_16009);
and U16466 (N_16466,N_16385,N_16085);
or U16467 (N_16467,N_16315,N_16215);
nand U16468 (N_16468,N_16066,N_16265);
nor U16469 (N_16469,N_16211,N_16036);
nor U16470 (N_16470,N_16049,N_16143);
and U16471 (N_16471,N_16266,N_16247);
and U16472 (N_16472,N_16005,N_16194);
or U16473 (N_16473,N_16310,N_16344);
nand U16474 (N_16474,N_16371,N_16213);
nor U16475 (N_16475,N_16386,N_16168);
nor U16476 (N_16476,N_16355,N_16293);
and U16477 (N_16477,N_16129,N_16299);
nor U16478 (N_16478,N_16292,N_16008);
and U16479 (N_16479,N_16033,N_16206);
nand U16480 (N_16480,N_16173,N_16140);
nor U16481 (N_16481,N_16032,N_16069);
and U16482 (N_16482,N_16192,N_16341);
and U16483 (N_16483,N_16128,N_16000);
or U16484 (N_16484,N_16280,N_16364);
or U16485 (N_16485,N_16068,N_16086);
or U16486 (N_16486,N_16241,N_16261);
and U16487 (N_16487,N_16246,N_16189);
and U16488 (N_16488,N_16115,N_16255);
and U16489 (N_16489,N_16116,N_16323);
nor U16490 (N_16490,N_16029,N_16250);
or U16491 (N_16491,N_16276,N_16155);
and U16492 (N_16492,N_16224,N_16031);
and U16493 (N_16493,N_16160,N_16393);
xor U16494 (N_16494,N_16164,N_16058);
nand U16495 (N_16495,N_16161,N_16181);
or U16496 (N_16496,N_16290,N_16028);
or U16497 (N_16497,N_16239,N_16198);
and U16498 (N_16498,N_16396,N_16367);
and U16499 (N_16499,N_16333,N_16156);
nand U16500 (N_16500,N_16390,N_16234);
and U16501 (N_16501,N_16356,N_16294);
nor U16502 (N_16502,N_16349,N_16226);
and U16503 (N_16503,N_16177,N_16316);
and U16504 (N_16504,N_16002,N_16288);
or U16505 (N_16505,N_16289,N_16120);
nand U16506 (N_16506,N_16020,N_16319);
nand U16507 (N_16507,N_16382,N_16320);
nor U16508 (N_16508,N_16001,N_16394);
nand U16509 (N_16509,N_16061,N_16254);
or U16510 (N_16510,N_16152,N_16195);
nand U16511 (N_16511,N_16380,N_16070);
nor U16512 (N_16512,N_16242,N_16147);
and U16513 (N_16513,N_16112,N_16381);
nand U16514 (N_16514,N_16167,N_16063);
nand U16515 (N_16515,N_16375,N_16174);
nand U16516 (N_16516,N_16071,N_16065);
nand U16517 (N_16517,N_16119,N_16111);
and U16518 (N_16518,N_16267,N_16387);
nand U16519 (N_16519,N_16329,N_16014);
nor U16520 (N_16520,N_16142,N_16221);
nand U16521 (N_16521,N_16222,N_16172);
and U16522 (N_16522,N_16314,N_16374);
nor U16523 (N_16523,N_16130,N_16309);
nor U16524 (N_16524,N_16135,N_16038);
or U16525 (N_16525,N_16282,N_16011);
or U16526 (N_16526,N_16236,N_16080);
or U16527 (N_16527,N_16228,N_16017);
nor U16528 (N_16528,N_16377,N_16232);
and U16529 (N_16529,N_16007,N_16273);
and U16530 (N_16530,N_16004,N_16060);
and U16531 (N_16531,N_16117,N_16016);
or U16532 (N_16532,N_16334,N_16384);
nand U16533 (N_16533,N_16126,N_16026);
nor U16534 (N_16534,N_16107,N_16053);
and U16535 (N_16535,N_16338,N_16075);
and U16536 (N_16536,N_16102,N_16088);
nand U16537 (N_16537,N_16346,N_16295);
or U16538 (N_16538,N_16113,N_16122);
nand U16539 (N_16539,N_16108,N_16219);
or U16540 (N_16540,N_16342,N_16162);
or U16541 (N_16541,N_16397,N_16337);
nand U16542 (N_16542,N_16077,N_16244);
nand U16543 (N_16543,N_16052,N_16233);
or U16544 (N_16544,N_16141,N_16037);
nand U16545 (N_16545,N_16362,N_16200);
nor U16546 (N_16546,N_16131,N_16207);
or U16547 (N_16547,N_16348,N_16360);
nor U16548 (N_16548,N_16227,N_16082);
and U16549 (N_16549,N_16304,N_16157);
nand U16550 (N_16550,N_16279,N_16099);
or U16551 (N_16551,N_16165,N_16399);
or U16552 (N_16552,N_16044,N_16103);
or U16553 (N_16553,N_16313,N_16190);
nand U16554 (N_16554,N_16230,N_16170);
or U16555 (N_16555,N_16101,N_16262);
nand U16556 (N_16556,N_16015,N_16114);
and U16557 (N_16557,N_16327,N_16193);
nor U16558 (N_16558,N_16045,N_16300);
nand U16559 (N_16559,N_16132,N_16218);
and U16560 (N_16560,N_16245,N_16041);
and U16561 (N_16561,N_16258,N_16083);
and U16562 (N_16562,N_16048,N_16148);
and U16563 (N_16563,N_16034,N_16263);
nor U16564 (N_16564,N_16345,N_16249);
nand U16565 (N_16565,N_16073,N_16220);
or U16566 (N_16566,N_16158,N_16264);
and U16567 (N_16567,N_16139,N_16123);
or U16568 (N_16568,N_16064,N_16169);
or U16569 (N_16569,N_16138,N_16322);
or U16570 (N_16570,N_16125,N_16324);
nand U16571 (N_16571,N_16024,N_16284);
and U16572 (N_16572,N_16271,N_16110);
nand U16573 (N_16573,N_16357,N_16057);
nor U16574 (N_16574,N_16124,N_16343);
nor U16575 (N_16575,N_16361,N_16035);
nand U16576 (N_16576,N_16078,N_16306);
xnor U16577 (N_16577,N_16260,N_16328);
or U16578 (N_16578,N_16018,N_16312);
and U16579 (N_16579,N_16339,N_16326);
and U16580 (N_16580,N_16225,N_16208);
and U16581 (N_16581,N_16389,N_16149);
and U16582 (N_16582,N_16072,N_16373);
nand U16583 (N_16583,N_16321,N_16093);
nor U16584 (N_16584,N_16197,N_16204);
and U16585 (N_16585,N_16368,N_16277);
and U16586 (N_16586,N_16154,N_16046);
or U16587 (N_16587,N_16275,N_16358);
or U16588 (N_16588,N_16118,N_16253);
nand U16589 (N_16589,N_16019,N_16166);
and U16590 (N_16590,N_16331,N_16302);
or U16591 (N_16591,N_16212,N_16003);
nor U16592 (N_16592,N_16106,N_16370);
and U16593 (N_16593,N_16089,N_16366);
and U16594 (N_16594,N_16090,N_16081);
or U16595 (N_16595,N_16051,N_16178);
nand U16596 (N_16596,N_16203,N_16047);
nand U16597 (N_16597,N_16127,N_16285);
nor U16598 (N_16598,N_16286,N_16365);
nand U16599 (N_16599,N_16084,N_16251);
nor U16600 (N_16600,N_16075,N_16174);
or U16601 (N_16601,N_16040,N_16319);
and U16602 (N_16602,N_16134,N_16272);
nor U16603 (N_16603,N_16387,N_16154);
or U16604 (N_16604,N_16379,N_16368);
nand U16605 (N_16605,N_16097,N_16041);
or U16606 (N_16606,N_16293,N_16324);
or U16607 (N_16607,N_16320,N_16175);
nor U16608 (N_16608,N_16394,N_16352);
nand U16609 (N_16609,N_16224,N_16223);
nand U16610 (N_16610,N_16114,N_16026);
nor U16611 (N_16611,N_16318,N_16078);
nor U16612 (N_16612,N_16398,N_16373);
nor U16613 (N_16613,N_16224,N_16368);
nand U16614 (N_16614,N_16129,N_16154);
or U16615 (N_16615,N_16195,N_16061);
nor U16616 (N_16616,N_16359,N_16017);
and U16617 (N_16617,N_16195,N_16288);
nand U16618 (N_16618,N_16110,N_16070);
and U16619 (N_16619,N_16129,N_16328);
nor U16620 (N_16620,N_16112,N_16111);
nand U16621 (N_16621,N_16138,N_16378);
nand U16622 (N_16622,N_16114,N_16395);
nand U16623 (N_16623,N_16272,N_16186);
or U16624 (N_16624,N_16022,N_16300);
nor U16625 (N_16625,N_16017,N_16383);
nand U16626 (N_16626,N_16374,N_16262);
or U16627 (N_16627,N_16374,N_16275);
nand U16628 (N_16628,N_16112,N_16189);
or U16629 (N_16629,N_16274,N_16046);
or U16630 (N_16630,N_16071,N_16061);
nand U16631 (N_16631,N_16071,N_16255);
and U16632 (N_16632,N_16180,N_16067);
nand U16633 (N_16633,N_16282,N_16168);
or U16634 (N_16634,N_16073,N_16346);
or U16635 (N_16635,N_16386,N_16165);
and U16636 (N_16636,N_16090,N_16169);
or U16637 (N_16637,N_16154,N_16146);
or U16638 (N_16638,N_16397,N_16096);
or U16639 (N_16639,N_16359,N_16008);
nor U16640 (N_16640,N_16298,N_16207);
nand U16641 (N_16641,N_16325,N_16028);
nor U16642 (N_16642,N_16031,N_16061);
nor U16643 (N_16643,N_16088,N_16232);
nor U16644 (N_16644,N_16093,N_16085);
or U16645 (N_16645,N_16254,N_16078);
or U16646 (N_16646,N_16127,N_16089);
or U16647 (N_16647,N_16209,N_16017);
nand U16648 (N_16648,N_16261,N_16379);
nor U16649 (N_16649,N_16192,N_16285);
nand U16650 (N_16650,N_16069,N_16061);
and U16651 (N_16651,N_16136,N_16128);
or U16652 (N_16652,N_16311,N_16261);
nor U16653 (N_16653,N_16276,N_16349);
nor U16654 (N_16654,N_16374,N_16029);
or U16655 (N_16655,N_16391,N_16105);
nor U16656 (N_16656,N_16184,N_16282);
or U16657 (N_16657,N_16193,N_16161);
nor U16658 (N_16658,N_16027,N_16391);
nand U16659 (N_16659,N_16321,N_16251);
and U16660 (N_16660,N_16370,N_16091);
xor U16661 (N_16661,N_16157,N_16229);
and U16662 (N_16662,N_16119,N_16353);
nor U16663 (N_16663,N_16061,N_16179);
nor U16664 (N_16664,N_16248,N_16216);
nand U16665 (N_16665,N_16123,N_16358);
or U16666 (N_16666,N_16076,N_16236);
or U16667 (N_16667,N_16116,N_16240);
nand U16668 (N_16668,N_16161,N_16237);
nand U16669 (N_16669,N_16072,N_16364);
and U16670 (N_16670,N_16182,N_16133);
nand U16671 (N_16671,N_16137,N_16122);
nor U16672 (N_16672,N_16246,N_16114);
and U16673 (N_16673,N_16072,N_16067);
or U16674 (N_16674,N_16265,N_16361);
or U16675 (N_16675,N_16029,N_16082);
or U16676 (N_16676,N_16298,N_16021);
nor U16677 (N_16677,N_16112,N_16192);
or U16678 (N_16678,N_16044,N_16118);
or U16679 (N_16679,N_16108,N_16120);
nand U16680 (N_16680,N_16342,N_16074);
nand U16681 (N_16681,N_16316,N_16001);
or U16682 (N_16682,N_16351,N_16210);
nor U16683 (N_16683,N_16057,N_16029);
nor U16684 (N_16684,N_16315,N_16358);
or U16685 (N_16685,N_16388,N_16397);
and U16686 (N_16686,N_16020,N_16061);
nor U16687 (N_16687,N_16058,N_16090);
nand U16688 (N_16688,N_16036,N_16243);
and U16689 (N_16689,N_16048,N_16353);
and U16690 (N_16690,N_16332,N_16080);
and U16691 (N_16691,N_16282,N_16073);
nand U16692 (N_16692,N_16084,N_16144);
or U16693 (N_16693,N_16326,N_16006);
nand U16694 (N_16694,N_16223,N_16015);
xnor U16695 (N_16695,N_16013,N_16370);
nor U16696 (N_16696,N_16261,N_16000);
and U16697 (N_16697,N_16079,N_16171);
nor U16698 (N_16698,N_16099,N_16053);
nand U16699 (N_16699,N_16373,N_16280);
nor U16700 (N_16700,N_16130,N_16228);
and U16701 (N_16701,N_16193,N_16055);
or U16702 (N_16702,N_16094,N_16153);
nor U16703 (N_16703,N_16025,N_16058);
and U16704 (N_16704,N_16038,N_16065);
or U16705 (N_16705,N_16360,N_16253);
and U16706 (N_16706,N_16301,N_16148);
nand U16707 (N_16707,N_16383,N_16106);
nand U16708 (N_16708,N_16306,N_16137);
nor U16709 (N_16709,N_16300,N_16207);
or U16710 (N_16710,N_16017,N_16030);
nor U16711 (N_16711,N_16141,N_16210);
nor U16712 (N_16712,N_16140,N_16022);
nor U16713 (N_16713,N_16318,N_16273);
and U16714 (N_16714,N_16276,N_16018);
nor U16715 (N_16715,N_16195,N_16054);
nor U16716 (N_16716,N_16273,N_16102);
xor U16717 (N_16717,N_16067,N_16053);
nor U16718 (N_16718,N_16158,N_16181);
and U16719 (N_16719,N_16163,N_16390);
nand U16720 (N_16720,N_16304,N_16126);
and U16721 (N_16721,N_16141,N_16332);
nor U16722 (N_16722,N_16196,N_16302);
or U16723 (N_16723,N_16331,N_16152);
nor U16724 (N_16724,N_16382,N_16272);
and U16725 (N_16725,N_16053,N_16100);
and U16726 (N_16726,N_16171,N_16333);
nor U16727 (N_16727,N_16269,N_16231);
or U16728 (N_16728,N_16073,N_16321);
and U16729 (N_16729,N_16182,N_16135);
nand U16730 (N_16730,N_16311,N_16249);
and U16731 (N_16731,N_16387,N_16046);
and U16732 (N_16732,N_16230,N_16279);
and U16733 (N_16733,N_16040,N_16130);
nand U16734 (N_16734,N_16399,N_16298);
or U16735 (N_16735,N_16218,N_16373);
nor U16736 (N_16736,N_16283,N_16026);
nand U16737 (N_16737,N_16146,N_16264);
and U16738 (N_16738,N_16121,N_16108);
and U16739 (N_16739,N_16026,N_16028);
or U16740 (N_16740,N_16300,N_16344);
or U16741 (N_16741,N_16350,N_16020);
and U16742 (N_16742,N_16273,N_16027);
or U16743 (N_16743,N_16244,N_16203);
nand U16744 (N_16744,N_16126,N_16281);
nor U16745 (N_16745,N_16363,N_16030);
nand U16746 (N_16746,N_16334,N_16164);
nand U16747 (N_16747,N_16011,N_16175);
and U16748 (N_16748,N_16180,N_16227);
and U16749 (N_16749,N_16376,N_16127);
and U16750 (N_16750,N_16271,N_16293);
nand U16751 (N_16751,N_16297,N_16277);
nor U16752 (N_16752,N_16168,N_16361);
or U16753 (N_16753,N_16115,N_16241);
or U16754 (N_16754,N_16217,N_16225);
and U16755 (N_16755,N_16365,N_16027);
nor U16756 (N_16756,N_16136,N_16245);
and U16757 (N_16757,N_16327,N_16319);
nand U16758 (N_16758,N_16275,N_16165);
and U16759 (N_16759,N_16240,N_16203);
or U16760 (N_16760,N_16114,N_16350);
nand U16761 (N_16761,N_16292,N_16285);
nor U16762 (N_16762,N_16071,N_16325);
nand U16763 (N_16763,N_16035,N_16198);
nand U16764 (N_16764,N_16126,N_16023);
or U16765 (N_16765,N_16020,N_16128);
and U16766 (N_16766,N_16100,N_16126);
or U16767 (N_16767,N_16300,N_16369);
nor U16768 (N_16768,N_16047,N_16114);
nor U16769 (N_16769,N_16318,N_16043);
nand U16770 (N_16770,N_16034,N_16319);
nand U16771 (N_16771,N_16005,N_16310);
or U16772 (N_16772,N_16140,N_16353);
and U16773 (N_16773,N_16219,N_16290);
nor U16774 (N_16774,N_16013,N_16293);
and U16775 (N_16775,N_16043,N_16117);
nor U16776 (N_16776,N_16262,N_16209);
nor U16777 (N_16777,N_16378,N_16050);
nand U16778 (N_16778,N_16221,N_16318);
nand U16779 (N_16779,N_16251,N_16294);
and U16780 (N_16780,N_16182,N_16122);
or U16781 (N_16781,N_16389,N_16394);
and U16782 (N_16782,N_16199,N_16188);
and U16783 (N_16783,N_16177,N_16350);
and U16784 (N_16784,N_16386,N_16045);
nor U16785 (N_16785,N_16017,N_16303);
nand U16786 (N_16786,N_16082,N_16360);
nor U16787 (N_16787,N_16158,N_16398);
or U16788 (N_16788,N_16043,N_16235);
nand U16789 (N_16789,N_16041,N_16131);
and U16790 (N_16790,N_16218,N_16351);
or U16791 (N_16791,N_16348,N_16329);
and U16792 (N_16792,N_16072,N_16088);
or U16793 (N_16793,N_16029,N_16257);
nor U16794 (N_16794,N_16146,N_16020);
nor U16795 (N_16795,N_16301,N_16394);
nor U16796 (N_16796,N_16279,N_16105);
and U16797 (N_16797,N_16197,N_16335);
or U16798 (N_16798,N_16207,N_16176);
and U16799 (N_16799,N_16266,N_16335);
or U16800 (N_16800,N_16535,N_16430);
nand U16801 (N_16801,N_16603,N_16687);
or U16802 (N_16802,N_16481,N_16634);
and U16803 (N_16803,N_16538,N_16589);
or U16804 (N_16804,N_16762,N_16774);
nand U16805 (N_16805,N_16661,N_16401);
and U16806 (N_16806,N_16614,N_16644);
and U16807 (N_16807,N_16722,N_16460);
and U16808 (N_16808,N_16699,N_16599);
and U16809 (N_16809,N_16658,N_16587);
and U16810 (N_16810,N_16709,N_16609);
or U16811 (N_16811,N_16767,N_16412);
or U16812 (N_16812,N_16441,N_16453);
and U16813 (N_16813,N_16763,N_16531);
nand U16814 (N_16814,N_16575,N_16542);
nor U16815 (N_16815,N_16653,N_16488);
and U16816 (N_16816,N_16546,N_16469);
nor U16817 (N_16817,N_16734,N_16438);
nand U16818 (N_16818,N_16465,N_16655);
nand U16819 (N_16819,N_16704,N_16640);
nor U16820 (N_16820,N_16731,N_16627);
nand U16821 (N_16821,N_16549,N_16406);
and U16822 (N_16822,N_16606,N_16632);
and U16823 (N_16823,N_16418,N_16678);
nor U16824 (N_16824,N_16682,N_16543);
and U16825 (N_16825,N_16563,N_16751);
or U16826 (N_16826,N_16732,N_16552);
nand U16827 (N_16827,N_16663,N_16649);
and U16828 (N_16828,N_16548,N_16689);
or U16829 (N_16829,N_16679,N_16659);
nand U16830 (N_16830,N_16404,N_16623);
nor U16831 (N_16831,N_16684,N_16555);
nor U16832 (N_16832,N_16757,N_16509);
or U16833 (N_16833,N_16675,N_16502);
nand U16834 (N_16834,N_16739,N_16760);
or U16835 (N_16835,N_16773,N_16437);
nand U16836 (N_16836,N_16786,N_16781);
or U16837 (N_16837,N_16500,N_16586);
nor U16838 (N_16838,N_16748,N_16654);
and U16839 (N_16839,N_16780,N_16499);
or U16840 (N_16840,N_16651,N_16671);
or U16841 (N_16841,N_16428,N_16667);
or U16842 (N_16842,N_16424,N_16777);
xnor U16843 (N_16843,N_16512,N_16723);
and U16844 (N_16844,N_16440,N_16436);
nor U16845 (N_16845,N_16683,N_16419);
or U16846 (N_16846,N_16420,N_16733);
or U16847 (N_16847,N_16685,N_16525);
nor U16848 (N_16848,N_16592,N_16454);
or U16849 (N_16849,N_16426,N_16539);
nand U16850 (N_16850,N_16666,N_16434);
and U16851 (N_16851,N_16585,N_16456);
and U16852 (N_16852,N_16580,N_16700);
nor U16853 (N_16853,N_16544,N_16583);
nand U16854 (N_16854,N_16743,N_16520);
or U16855 (N_16855,N_16421,N_16506);
or U16856 (N_16856,N_16534,N_16533);
nand U16857 (N_16857,N_16630,N_16772);
and U16858 (N_16858,N_16501,N_16672);
and U16859 (N_16859,N_16680,N_16571);
and U16860 (N_16860,N_16598,N_16676);
or U16861 (N_16861,N_16726,N_16519);
and U16862 (N_16862,N_16411,N_16513);
nor U16863 (N_16863,N_16686,N_16590);
nor U16864 (N_16864,N_16656,N_16776);
or U16865 (N_16865,N_16737,N_16769);
nor U16866 (N_16866,N_16712,N_16507);
nor U16867 (N_16867,N_16641,N_16629);
or U16868 (N_16868,N_16466,N_16615);
or U16869 (N_16869,N_16462,N_16472);
nand U16870 (N_16870,N_16783,N_16574);
nand U16871 (N_16871,N_16435,N_16558);
nand U16872 (N_16872,N_16797,N_16711);
and U16873 (N_16873,N_16573,N_16607);
or U16874 (N_16874,N_16497,N_16619);
nand U16875 (N_16875,N_16638,N_16715);
nor U16876 (N_16876,N_16639,N_16647);
nor U16877 (N_16877,N_16601,N_16668);
or U16878 (N_16878,N_16727,N_16681);
or U16879 (N_16879,N_16511,N_16725);
nor U16880 (N_16880,N_16556,N_16514);
nand U16881 (N_16881,N_16554,N_16405);
nand U16882 (N_16882,N_16622,N_16528);
nand U16883 (N_16883,N_16596,N_16621);
and U16884 (N_16884,N_16439,N_16738);
nand U16885 (N_16885,N_16650,N_16487);
nand U16886 (N_16886,N_16610,N_16728);
nand U16887 (N_16887,N_16402,N_16518);
nor U16888 (N_16888,N_16477,N_16444);
or U16889 (N_16889,N_16799,N_16787);
xor U16890 (N_16890,N_16720,N_16673);
nor U16891 (N_16891,N_16692,N_16597);
or U16892 (N_16892,N_16407,N_16752);
and U16893 (N_16893,N_16642,N_16457);
nand U16894 (N_16894,N_16625,N_16527);
nand U16895 (N_16895,N_16648,N_16522);
nor U16896 (N_16896,N_16532,N_16761);
nor U16897 (N_16897,N_16482,N_16714);
or U16898 (N_16898,N_16459,N_16403);
xnor U16899 (N_16899,N_16551,N_16793);
or U16900 (N_16900,N_16701,N_16505);
and U16901 (N_16901,N_16479,N_16474);
nor U16902 (N_16902,N_16576,N_16643);
and U16903 (N_16903,N_16768,N_16717);
and U16904 (N_16904,N_16478,N_16451);
xnor U16905 (N_16905,N_16766,N_16624);
or U16906 (N_16906,N_16788,N_16742);
or U16907 (N_16907,N_16600,N_16657);
and U16908 (N_16908,N_16785,N_16702);
and U16909 (N_16909,N_16521,N_16662);
nor U16910 (N_16910,N_16559,N_16794);
or U16911 (N_16911,N_16461,N_16495);
nand U16912 (N_16912,N_16694,N_16594);
or U16913 (N_16913,N_16703,N_16526);
nand U16914 (N_16914,N_16753,N_16557);
nand U16915 (N_16915,N_16631,N_16523);
nor U16916 (N_16916,N_16540,N_16705);
nand U16917 (N_16917,N_16747,N_16645);
and U16918 (N_16918,N_16413,N_16605);
nor U16919 (N_16919,N_16423,N_16503);
xor U16920 (N_16920,N_16758,N_16467);
nor U16921 (N_16921,N_16579,N_16541);
nand U16922 (N_16922,N_16798,N_16612);
nor U16923 (N_16923,N_16568,N_16566);
nor U16924 (N_16924,N_16664,N_16468);
or U16925 (N_16925,N_16516,N_16431);
nor U16926 (N_16926,N_16789,N_16792);
or U16927 (N_16927,N_16670,N_16446);
or U16928 (N_16928,N_16425,N_16724);
or U16929 (N_16929,N_16448,N_16635);
and U16930 (N_16930,N_16791,N_16409);
nor U16931 (N_16931,N_16464,N_16782);
or U16932 (N_16932,N_16442,N_16691);
nand U16933 (N_16933,N_16674,N_16765);
nor U16934 (N_16934,N_16569,N_16553);
nand U16935 (N_16935,N_16713,N_16484);
and U16936 (N_16936,N_16494,N_16755);
nor U16937 (N_16937,N_16562,N_16779);
nand U16938 (N_16938,N_16473,N_16633);
or U16939 (N_16939,N_16618,N_16617);
xnor U16940 (N_16940,N_16449,N_16480);
nand U16941 (N_16941,N_16524,N_16616);
nand U16942 (N_16942,N_16749,N_16508);
nor U16943 (N_16943,N_16690,N_16486);
or U16944 (N_16944,N_16536,N_16578);
nand U16945 (N_16945,N_16537,N_16417);
nor U16946 (N_16946,N_16608,N_16447);
and U16947 (N_16947,N_16470,N_16445);
or U16948 (N_16948,N_16652,N_16577);
nand U16949 (N_16949,N_16795,N_16471);
nor U16950 (N_16950,N_16570,N_16410);
and U16951 (N_16951,N_16707,N_16408);
nand U16952 (N_16952,N_16626,N_16730);
nor U16953 (N_16953,N_16427,N_16744);
nand U16954 (N_16954,N_16771,N_16591);
nand U16955 (N_16955,N_16665,N_16669);
or U16956 (N_16956,N_16491,N_16706);
nor U16957 (N_16957,N_16565,N_16493);
and U16958 (N_16958,N_16604,N_16452);
nand U16959 (N_16959,N_16510,N_16595);
nand U16960 (N_16960,N_16564,N_16490);
nand U16961 (N_16961,N_16611,N_16517);
nor U16962 (N_16962,N_16560,N_16400);
and U16963 (N_16963,N_16778,N_16588);
nand U16964 (N_16964,N_16475,N_16593);
or U16965 (N_16965,N_16489,N_16740);
nand U16966 (N_16966,N_16756,N_16415);
or U16967 (N_16967,N_16504,N_16572);
and U16968 (N_16968,N_16476,N_16677);
nor U16969 (N_16969,N_16414,N_16567);
nor U16970 (N_16970,N_16628,N_16498);
or U16971 (N_16971,N_16416,N_16746);
or U16972 (N_16972,N_16429,N_16710);
or U16973 (N_16973,N_16796,N_16530);
nor U16974 (N_16974,N_16637,N_16721);
and U16975 (N_16975,N_16547,N_16492);
nand U16976 (N_16976,N_16695,N_16697);
nor U16977 (N_16977,N_16708,N_16581);
nand U16978 (N_16978,N_16485,N_16775);
and U16979 (N_16979,N_16432,N_16443);
nor U16980 (N_16980,N_16584,N_16602);
nor U16981 (N_16981,N_16745,N_16550);
xor U16982 (N_16982,N_16741,N_16688);
nand U16983 (N_16983,N_16463,N_16693);
xor U16984 (N_16984,N_16458,N_16716);
nor U16985 (N_16985,N_16515,N_16784);
nor U16986 (N_16986,N_16764,N_16698);
nand U16987 (N_16987,N_16433,N_16660);
nor U16988 (N_16988,N_16561,N_16735);
or U16989 (N_16989,N_16529,N_16620);
and U16990 (N_16990,N_16545,N_16750);
or U16991 (N_16991,N_16770,N_16759);
nand U16992 (N_16992,N_16736,N_16483);
nor U16993 (N_16993,N_16719,N_16582);
nor U16994 (N_16994,N_16790,N_16646);
nand U16995 (N_16995,N_16696,N_16422);
nand U16996 (N_16996,N_16613,N_16636);
nor U16997 (N_16997,N_16496,N_16450);
or U16998 (N_16998,N_16718,N_16754);
nor U16999 (N_16999,N_16729,N_16455);
or U17000 (N_17000,N_16614,N_16641);
nor U17001 (N_17001,N_16483,N_16573);
or U17002 (N_17002,N_16577,N_16784);
or U17003 (N_17003,N_16734,N_16490);
nor U17004 (N_17004,N_16628,N_16458);
or U17005 (N_17005,N_16408,N_16621);
nand U17006 (N_17006,N_16558,N_16750);
and U17007 (N_17007,N_16481,N_16758);
nand U17008 (N_17008,N_16743,N_16423);
nand U17009 (N_17009,N_16665,N_16641);
nor U17010 (N_17010,N_16789,N_16684);
nand U17011 (N_17011,N_16707,N_16738);
nand U17012 (N_17012,N_16717,N_16611);
or U17013 (N_17013,N_16539,N_16415);
and U17014 (N_17014,N_16655,N_16425);
nand U17015 (N_17015,N_16727,N_16534);
nand U17016 (N_17016,N_16538,N_16610);
nor U17017 (N_17017,N_16521,N_16520);
or U17018 (N_17018,N_16608,N_16568);
and U17019 (N_17019,N_16545,N_16556);
nand U17020 (N_17020,N_16583,N_16730);
or U17021 (N_17021,N_16747,N_16544);
nand U17022 (N_17022,N_16693,N_16590);
and U17023 (N_17023,N_16490,N_16433);
nand U17024 (N_17024,N_16607,N_16650);
nand U17025 (N_17025,N_16662,N_16528);
nand U17026 (N_17026,N_16667,N_16406);
nor U17027 (N_17027,N_16798,N_16779);
or U17028 (N_17028,N_16752,N_16428);
nor U17029 (N_17029,N_16793,N_16785);
or U17030 (N_17030,N_16491,N_16786);
nor U17031 (N_17031,N_16696,N_16615);
nor U17032 (N_17032,N_16601,N_16776);
nor U17033 (N_17033,N_16654,N_16671);
and U17034 (N_17034,N_16453,N_16655);
nor U17035 (N_17035,N_16778,N_16748);
xnor U17036 (N_17036,N_16624,N_16534);
or U17037 (N_17037,N_16798,N_16724);
and U17038 (N_17038,N_16766,N_16703);
and U17039 (N_17039,N_16507,N_16761);
xnor U17040 (N_17040,N_16671,N_16772);
or U17041 (N_17041,N_16751,N_16645);
nor U17042 (N_17042,N_16468,N_16632);
or U17043 (N_17043,N_16794,N_16494);
nand U17044 (N_17044,N_16404,N_16539);
or U17045 (N_17045,N_16484,N_16430);
and U17046 (N_17046,N_16768,N_16574);
nor U17047 (N_17047,N_16416,N_16715);
or U17048 (N_17048,N_16648,N_16770);
and U17049 (N_17049,N_16644,N_16521);
nor U17050 (N_17050,N_16513,N_16652);
nand U17051 (N_17051,N_16529,N_16677);
nor U17052 (N_17052,N_16731,N_16422);
nand U17053 (N_17053,N_16720,N_16647);
nand U17054 (N_17054,N_16451,N_16458);
or U17055 (N_17055,N_16762,N_16674);
nor U17056 (N_17056,N_16703,N_16679);
and U17057 (N_17057,N_16556,N_16711);
nor U17058 (N_17058,N_16530,N_16456);
nor U17059 (N_17059,N_16439,N_16621);
nand U17060 (N_17060,N_16535,N_16781);
or U17061 (N_17061,N_16573,N_16605);
or U17062 (N_17062,N_16505,N_16459);
nor U17063 (N_17063,N_16538,N_16687);
or U17064 (N_17064,N_16491,N_16601);
or U17065 (N_17065,N_16691,N_16648);
and U17066 (N_17066,N_16577,N_16523);
nor U17067 (N_17067,N_16754,N_16473);
or U17068 (N_17068,N_16645,N_16703);
nand U17069 (N_17069,N_16506,N_16412);
nand U17070 (N_17070,N_16592,N_16516);
nor U17071 (N_17071,N_16580,N_16776);
nor U17072 (N_17072,N_16644,N_16795);
and U17073 (N_17073,N_16765,N_16477);
and U17074 (N_17074,N_16753,N_16679);
and U17075 (N_17075,N_16631,N_16569);
and U17076 (N_17076,N_16456,N_16529);
and U17077 (N_17077,N_16608,N_16787);
nor U17078 (N_17078,N_16419,N_16648);
or U17079 (N_17079,N_16624,N_16622);
nand U17080 (N_17080,N_16433,N_16454);
nor U17081 (N_17081,N_16465,N_16756);
nor U17082 (N_17082,N_16697,N_16706);
nand U17083 (N_17083,N_16630,N_16415);
nor U17084 (N_17084,N_16447,N_16647);
and U17085 (N_17085,N_16724,N_16740);
or U17086 (N_17086,N_16411,N_16555);
nor U17087 (N_17087,N_16708,N_16772);
or U17088 (N_17088,N_16798,N_16511);
nor U17089 (N_17089,N_16743,N_16518);
and U17090 (N_17090,N_16520,N_16497);
or U17091 (N_17091,N_16744,N_16629);
nand U17092 (N_17092,N_16495,N_16427);
nand U17093 (N_17093,N_16484,N_16620);
nand U17094 (N_17094,N_16419,N_16531);
and U17095 (N_17095,N_16436,N_16421);
nand U17096 (N_17096,N_16771,N_16558);
nor U17097 (N_17097,N_16569,N_16566);
or U17098 (N_17098,N_16720,N_16577);
or U17099 (N_17099,N_16635,N_16594);
or U17100 (N_17100,N_16539,N_16685);
and U17101 (N_17101,N_16790,N_16691);
nand U17102 (N_17102,N_16654,N_16784);
nand U17103 (N_17103,N_16751,N_16442);
or U17104 (N_17104,N_16432,N_16609);
nand U17105 (N_17105,N_16618,N_16581);
and U17106 (N_17106,N_16601,N_16617);
nor U17107 (N_17107,N_16480,N_16551);
nand U17108 (N_17108,N_16487,N_16547);
or U17109 (N_17109,N_16667,N_16771);
or U17110 (N_17110,N_16422,N_16417);
nor U17111 (N_17111,N_16709,N_16684);
or U17112 (N_17112,N_16684,N_16626);
nand U17113 (N_17113,N_16438,N_16758);
nand U17114 (N_17114,N_16730,N_16657);
nand U17115 (N_17115,N_16468,N_16636);
or U17116 (N_17116,N_16680,N_16626);
or U17117 (N_17117,N_16601,N_16744);
and U17118 (N_17118,N_16758,N_16733);
and U17119 (N_17119,N_16639,N_16454);
nand U17120 (N_17120,N_16516,N_16594);
nand U17121 (N_17121,N_16657,N_16781);
nand U17122 (N_17122,N_16601,N_16789);
and U17123 (N_17123,N_16620,N_16785);
nor U17124 (N_17124,N_16730,N_16782);
nand U17125 (N_17125,N_16654,N_16582);
nor U17126 (N_17126,N_16448,N_16695);
and U17127 (N_17127,N_16400,N_16436);
and U17128 (N_17128,N_16602,N_16720);
or U17129 (N_17129,N_16603,N_16677);
nor U17130 (N_17130,N_16484,N_16697);
nand U17131 (N_17131,N_16550,N_16770);
or U17132 (N_17132,N_16681,N_16722);
nand U17133 (N_17133,N_16529,N_16480);
or U17134 (N_17134,N_16478,N_16658);
and U17135 (N_17135,N_16587,N_16475);
or U17136 (N_17136,N_16661,N_16498);
nor U17137 (N_17137,N_16486,N_16618);
and U17138 (N_17138,N_16744,N_16726);
or U17139 (N_17139,N_16723,N_16651);
nand U17140 (N_17140,N_16757,N_16688);
nor U17141 (N_17141,N_16696,N_16748);
nand U17142 (N_17142,N_16784,N_16555);
nand U17143 (N_17143,N_16786,N_16656);
and U17144 (N_17144,N_16726,N_16428);
nor U17145 (N_17145,N_16795,N_16758);
nor U17146 (N_17146,N_16713,N_16743);
nand U17147 (N_17147,N_16647,N_16497);
nor U17148 (N_17148,N_16682,N_16638);
or U17149 (N_17149,N_16594,N_16459);
nand U17150 (N_17150,N_16590,N_16513);
nand U17151 (N_17151,N_16580,N_16450);
nor U17152 (N_17152,N_16703,N_16509);
nand U17153 (N_17153,N_16636,N_16459);
nor U17154 (N_17154,N_16759,N_16688);
and U17155 (N_17155,N_16518,N_16522);
nor U17156 (N_17156,N_16521,N_16535);
or U17157 (N_17157,N_16644,N_16608);
or U17158 (N_17158,N_16548,N_16463);
or U17159 (N_17159,N_16708,N_16780);
and U17160 (N_17160,N_16468,N_16494);
nand U17161 (N_17161,N_16743,N_16680);
nor U17162 (N_17162,N_16656,N_16447);
nand U17163 (N_17163,N_16642,N_16413);
nor U17164 (N_17164,N_16665,N_16427);
nor U17165 (N_17165,N_16731,N_16733);
nor U17166 (N_17166,N_16600,N_16539);
nand U17167 (N_17167,N_16410,N_16601);
nand U17168 (N_17168,N_16458,N_16578);
or U17169 (N_17169,N_16705,N_16529);
and U17170 (N_17170,N_16643,N_16471);
nor U17171 (N_17171,N_16556,N_16692);
or U17172 (N_17172,N_16682,N_16477);
or U17173 (N_17173,N_16486,N_16470);
and U17174 (N_17174,N_16713,N_16731);
nor U17175 (N_17175,N_16517,N_16647);
and U17176 (N_17176,N_16534,N_16782);
nand U17177 (N_17177,N_16408,N_16629);
or U17178 (N_17178,N_16649,N_16494);
or U17179 (N_17179,N_16779,N_16422);
nand U17180 (N_17180,N_16481,N_16599);
and U17181 (N_17181,N_16705,N_16791);
or U17182 (N_17182,N_16585,N_16554);
nand U17183 (N_17183,N_16644,N_16783);
nand U17184 (N_17184,N_16511,N_16585);
nand U17185 (N_17185,N_16661,N_16667);
nand U17186 (N_17186,N_16553,N_16596);
or U17187 (N_17187,N_16639,N_16767);
nor U17188 (N_17188,N_16544,N_16596);
nand U17189 (N_17189,N_16569,N_16635);
nand U17190 (N_17190,N_16414,N_16795);
or U17191 (N_17191,N_16773,N_16642);
or U17192 (N_17192,N_16707,N_16737);
and U17193 (N_17193,N_16456,N_16498);
and U17194 (N_17194,N_16578,N_16512);
nor U17195 (N_17195,N_16567,N_16772);
nand U17196 (N_17196,N_16583,N_16712);
nand U17197 (N_17197,N_16611,N_16751);
nand U17198 (N_17198,N_16608,N_16672);
or U17199 (N_17199,N_16682,N_16575);
nand U17200 (N_17200,N_17179,N_17106);
or U17201 (N_17201,N_17021,N_16844);
nand U17202 (N_17202,N_17126,N_16816);
nor U17203 (N_17203,N_17031,N_17045);
nor U17204 (N_17204,N_17092,N_16826);
nand U17205 (N_17205,N_17034,N_17038);
and U17206 (N_17206,N_17145,N_17057);
nor U17207 (N_17207,N_16980,N_17164);
nor U17208 (N_17208,N_17067,N_16891);
nor U17209 (N_17209,N_17152,N_17079);
and U17210 (N_17210,N_17195,N_16962);
nor U17211 (N_17211,N_16943,N_17119);
xor U17212 (N_17212,N_17018,N_16992);
and U17213 (N_17213,N_16807,N_16843);
nor U17214 (N_17214,N_16839,N_17107);
nand U17215 (N_17215,N_17069,N_17175);
and U17216 (N_17216,N_16964,N_17177);
nor U17217 (N_17217,N_16921,N_16824);
nor U17218 (N_17218,N_17178,N_16919);
or U17219 (N_17219,N_16995,N_16814);
and U17220 (N_17220,N_16979,N_16915);
or U17221 (N_17221,N_17003,N_16867);
nor U17222 (N_17222,N_16856,N_16961);
or U17223 (N_17223,N_17155,N_16848);
nor U17224 (N_17224,N_16847,N_17176);
xor U17225 (N_17225,N_16935,N_16914);
and U17226 (N_17226,N_17037,N_17080);
nand U17227 (N_17227,N_16803,N_17082);
nor U17228 (N_17228,N_17011,N_17174);
or U17229 (N_17229,N_17066,N_16969);
or U17230 (N_17230,N_16936,N_16916);
or U17231 (N_17231,N_17188,N_17138);
or U17232 (N_17232,N_16859,N_16972);
nor U17233 (N_17233,N_17049,N_17035);
or U17234 (N_17234,N_17120,N_17058);
nor U17235 (N_17235,N_17137,N_16925);
nor U17236 (N_17236,N_17091,N_16905);
nor U17237 (N_17237,N_17148,N_16813);
or U17238 (N_17238,N_16850,N_17173);
nor U17239 (N_17239,N_17022,N_17103);
nand U17240 (N_17240,N_17167,N_17004);
or U17241 (N_17241,N_17059,N_17019);
or U17242 (N_17242,N_17190,N_16868);
or U17243 (N_17243,N_16892,N_17189);
or U17244 (N_17244,N_17054,N_16896);
and U17245 (N_17245,N_16895,N_16874);
and U17246 (N_17246,N_17182,N_17109);
and U17247 (N_17247,N_17196,N_17063);
nand U17248 (N_17248,N_16959,N_16990);
nor U17249 (N_17249,N_16886,N_16815);
or U17250 (N_17250,N_17170,N_16893);
nor U17251 (N_17251,N_16955,N_17186);
or U17252 (N_17252,N_17072,N_16897);
or U17253 (N_17253,N_16952,N_16842);
nor U17254 (N_17254,N_16997,N_17132);
nor U17255 (N_17255,N_17005,N_16909);
nand U17256 (N_17256,N_17023,N_16951);
nor U17257 (N_17257,N_17141,N_17007);
nand U17258 (N_17258,N_17042,N_16911);
nor U17259 (N_17259,N_17012,N_16864);
nand U17260 (N_17260,N_16827,N_17181);
nor U17261 (N_17261,N_17168,N_17036);
or U17262 (N_17262,N_16821,N_16890);
nand U17263 (N_17263,N_16963,N_16883);
and U17264 (N_17264,N_17117,N_16945);
nand U17265 (N_17265,N_17051,N_17029);
or U17266 (N_17266,N_17169,N_17136);
and U17267 (N_17267,N_17151,N_17146);
and U17268 (N_17268,N_16900,N_17127);
nand U17269 (N_17269,N_17135,N_16889);
nor U17270 (N_17270,N_17076,N_17013);
and U17271 (N_17271,N_16913,N_16817);
and U17272 (N_17272,N_17028,N_16818);
and U17273 (N_17273,N_16907,N_17194);
or U17274 (N_17274,N_16903,N_17165);
or U17275 (N_17275,N_16869,N_17143);
nor U17276 (N_17276,N_17184,N_17001);
or U17277 (N_17277,N_16993,N_16872);
nand U17278 (N_17278,N_17077,N_17187);
or U17279 (N_17279,N_17162,N_16879);
or U17280 (N_17280,N_17095,N_16970);
or U17281 (N_17281,N_17071,N_16941);
and U17282 (N_17282,N_17123,N_16823);
nor U17283 (N_17283,N_17033,N_16923);
or U17284 (N_17284,N_16860,N_16965);
nor U17285 (N_17285,N_17040,N_17070);
nor U17286 (N_17286,N_17147,N_17180);
or U17287 (N_17287,N_16849,N_16950);
nor U17288 (N_17288,N_16940,N_17133);
or U17289 (N_17289,N_17122,N_16924);
and U17290 (N_17290,N_16953,N_16967);
and U17291 (N_17291,N_16804,N_16899);
or U17292 (N_17292,N_16948,N_17192);
nand U17293 (N_17293,N_17010,N_17044);
xnor U17294 (N_17294,N_16881,N_17097);
nand U17295 (N_17295,N_16926,N_17084);
or U17296 (N_17296,N_17183,N_16981);
or U17297 (N_17297,N_17124,N_16986);
xnor U17298 (N_17298,N_16910,N_17006);
nor U17299 (N_17299,N_17197,N_16946);
nand U17300 (N_17300,N_16831,N_16938);
or U17301 (N_17301,N_16837,N_17089);
xor U17302 (N_17302,N_16838,N_16810);
nor U17303 (N_17303,N_16876,N_16819);
nor U17304 (N_17304,N_17199,N_17000);
nand U17305 (N_17305,N_16968,N_17157);
nor U17306 (N_17306,N_17093,N_17101);
nor U17307 (N_17307,N_16862,N_17185);
or U17308 (N_17308,N_17088,N_16882);
and U17309 (N_17309,N_17144,N_17128);
nor U17310 (N_17310,N_17161,N_17171);
and U17311 (N_17311,N_17149,N_17191);
or U17312 (N_17312,N_17061,N_17140);
or U17313 (N_17313,N_17153,N_16822);
and U17314 (N_17314,N_17163,N_16870);
nand U17315 (N_17315,N_17159,N_16989);
and U17316 (N_17316,N_16987,N_17015);
nand U17317 (N_17317,N_16853,N_17008);
or U17318 (N_17318,N_17074,N_17098);
and U17319 (N_17319,N_16937,N_17087);
nor U17320 (N_17320,N_16801,N_16858);
or U17321 (N_17321,N_17048,N_17024);
and U17322 (N_17322,N_16912,N_17125);
nor U17323 (N_17323,N_16960,N_17016);
nand U17324 (N_17324,N_17052,N_16825);
nor U17325 (N_17325,N_16851,N_17114);
nor U17326 (N_17326,N_17115,N_16939);
and U17327 (N_17327,N_16840,N_16894);
or U17328 (N_17328,N_17130,N_17154);
nand U17329 (N_17329,N_16871,N_16944);
or U17330 (N_17330,N_16977,N_16836);
and U17331 (N_17331,N_16934,N_17139);
nand U17332 (N_17332,N_16854,N_16855);
and U17333 (N_17333,N_16954,N_17172);
nand U17334 (N_17334,N_16957,N_16878);
nor U17335 (N_17335,N_17043,N_16920);
and U17336 (N_17336,N_16830,N_17198);
and U17337 (N_17337,N_17083,N_16829);
nand U17338 (N_17338,N_16861,N_17090);
or U17339 (N_17339,N_16863,N_17121);
or U17340 (N_17340,N_16976,N_16991);
nor U17341 (N_17341,N_17116,N_17050);
or U17342 (N_17342,N_17073,N_17158);
or U17343 (N_17343,N_16835,N_16994);
and U17344 (N_17344,N_17105,N_16802);
and U17345 (N_17345,N_16973,N_17002);
and U17346 (N_17346,N_17102,N_16978);
nand U17347 (N_17347,N_17150,N_17094);
nor U17348 (N_17348,N_16932,N_16820);
xor U17349 (N_17349,N_16996,N_17131);
nand U17350 (N_17350,N_17030,N_16885);
or U17351 (N_17351,N_16806,N_16949);
and U17352 (N_17352,N_17041,N_16873);
nor U17353 (N_17353,N_16956,N_17020);
and U17354 (N_17354,N_17075,N_16884);
or U17355 (N_17355,N_17065,N_16933);
nor U17356 (N_17356,N_16832,N_16984);
nor U17357 (N_17357,N_16811,N_17113);
nand U17358 (N_17358,N_17156,N_17142);
nor U17359 (N_17359,N_17055,N_17104);
nor U17360 (N_17360,N_16888,N_17160);
nor U17361 (N_17361,N_16812,N_17026);
nand U17362 (N_17362,N_16846,N_17009);
nand U17363 (N_17363,N_17100,N_16922);
nand U17364 (N_17364,N_17060,N_17062);
or U17365 (N_17365,N_17046,N_17129);
and U17366 (N_17366,N_17068,N_17081);
nor U17367 (N_17367,N_17099,N_16898);
nand U17368 (N_17368,N_17032,N_16975);
nor U17369 (N_17369,N_16971,N_16908);
and U17370 (N_17370,N_16947,N_16805);
and U17371 (N_17371,N_16800,N_17039);
and U17372 (N_17372,N_16904,N_17064);
or U17373 (N_17373,N_17086,N_17056);
or U17374 (N_17374,N_17118,N_16877);
or U17375 (N_17375,N_16931,N_17110);
nand U17376 (N_17376,N_16966,N_17112);
and U17377 (N_17377,N_16841,N_16828);
or U17378 (N_17378,N_16942,N_17085);
or U17379 (N_17379,N_16902,N_16930);
or U17380 (N_17380,N_16917,N_16808);
or U17381 (N_17381,N_17111,N_17096);
xnor U17382 (N_17382,N_17025,N_17166);
nand U17383 (N_17383,N_16834,N_17017);
or U17384 (N_17384,N_16866,N_16985);
or U17385 (N_17385,N_16833,N_16958);
and U17386 (N_17386,N_16974,N_16928);
nor U17387 (N_17387,N_16845,N_16865);
nand U17388 (N_17388,N_16988,N_17134);
nand U17389 (N_17389,N_17027,N_16929);
nor U17390 (N_17390,N_17047,N_16983);
nand U17391 (N_17391,N_17193,N_16880);
or U17392 (N_17392,N_17108,N_16901);
nor U17393 (N_17393,N_16887,N_16999);
nor U17394 (N_17394,N_16918,N_16857);
nor U17395 (N_17395,N_17014,N_17078);
and U17396 (N_17396,N_16809,N_16982);
and U17397 (N_17397,N_16906,N_16875);
and U17398 (N_17398,N_17053,N_16852);
and U17399 (N_17399,N_16927,N_16998);
or U17400 (N_17400,N_16893,N_17155);
nor U17401 (N_17401,N_17130,N_17074);
nor U17402 (N_17402,N_16888,N_17104);
or U17403 (N_17403,N_17106,N_16918);
or U17404 (N_17404,N_16911,N_17193);
nor U17405 (N_17405,N_17123,N_16811);
and U17406 (N_17406,N_16904,N_17076);
nand U17407 (N_17407,N_16844,N_17149);
and U17408 (N_17408,N_17113,N_16906);
or U17409 (N_17409,N_17127,N_16986);
nand U17410 (N_17410,N_17156,N_17122);
and U17411 (N_17411,N_16941,N_17129);
and U17412 (N_17412,N_17064,N_17061);
or U17413 (N_17413,N_17151,N_17098);
or U17414 (N_17414,N_17100,N_16948);
or U17415 (N_17415,N_16878,N_17092);
or U17416 (N_17416,N_16843,N_17141);
nand U17417 (N_17417,N_16893,N_16952);
and U17418 (N_17418,N_17044,N_16806);
and U17419 (N_17419,N_16920,N_16919);
nand U17420 (N_17420,N_16848,N_17190);
and U17421 (N_17421,N_16970,N_17102);
nand U17422 (N_17422,N_17182,N_16820);
and U17423 (N_17423,N_16933,N_16974);
nor U17424 (N_17424,N_16903,N_17166);
or U17425 (N_17425,N_16889,N_16883);
nor U17426 (N_17426,N_16997,N_16882);
nor U17427 (N_17427,N_16973,N_17065);
or U17428 (N_17428,N_17197,N_17106);
nor U17429 (N_17429,N_16878,N_16803);
nand U17430 (N_17430,N_16816,N_17194);
or U17431 (N_17431,N_17072,N_16935);
nor U17432 (N_17432,N_17056,N_17197);
or U17433 (N_17433,N_16971,N_16932);
or U17434 (N_17434,N_16935,N_17132);
nor U17435 (N_17435,N_16890,N_17027);
nor U17436 (N_17436,N_17078,N_16904);
or U17437 (N_17437,N_16818,N_16885);
or U17438 (N_17438,N_17005,N_16961);
nand U17439 (N_17439,N_16961,N_16841);
nand U17440 (N_17440,N_16824,N_17191);
and U17441 (N_17441,N_17114,N_17038);
nor U17442 (N_17442,N_17152,N_16824);
nand U17443 (N_17443,N_17163,N_16858);
nor U17444 (N_17444,N_17047,N_16879);
or U17445 (N_17445,N_16864,N_16997);
and U17446 (N_17446,N_17010,N_17159);
or U17447 (N_17447,N_17034,N_17033);
nand U17448 (N_17448,N_17056,N_16800);
and U17449 (N_17449,N_17120,N_17022);
or U17450 (N_17450,N_16940,N_16918);
or U17451 (N_17451,N_17156,N_17019);
and U17452 (N_17452,N_17176,N_17106);
nor U17453 (N_17453,N_17008,N_16945);
nor U17454 (N_17454,N_17157,N_16825);
nand U17455 (N_17455,N_16957,N_16994);
and U17456 (N_17456,N_16810,N_16922);
nand U17457 (N_17457,N_16889,N_17065);
or U17458 (N_17458,N_17079,N_16957);
or U17459 (N_17459,N_16856,N_17123);
nand U17460 (N_17460,N_16992,N_17000);
nor U17461 (N_17461,N_17139,N_17144);
and U17462 (N_17462,N_17077,N_16848);
xnor U17463 (N_17463,N_16934,N_17120);
or U17464 (N_17464,N_17158,N_17008);
nand U17465 (N_17465,N_17197,N_16833);
or U17466 (N_17466,N_17181,N_16803);
or U17467 (N_17467,N_17127,N_17078);
and U17468 (N_17468,N_16926,N_16818);
nand U17469 (N_17469,N_16983,N_17026);
and U17470 (N_17470,N_16888,N_16987);
xor U17471 (N_17471,N_16906,N_16917);
nand U17472 (N_17472,N_16853,N_17157);
or U17473 (N_17473,N_17072,N_16968);
or U17474 (N_17474,N_16998,N_17168);
nand U17475 (N_17475,N_16910,N_16836);
and U17476 (N_17476,N_16989,N_16944);
nor U17477 (N_17477,N_16876,N_16955);
and U17478 (N_17478,N_16850,N_16917);
and U17479 (N_17479,N_17100,N_16999);
nand U17480 (N_17480,N_17046,N_17108);
nand U17481 (N_17481,N_16900,N_17088);
nor U17482 (N_17482,N_16914,N_17027);
or U17483 (N_17483,N_17026,N_16841);
and U17484 (N_17484,N_16829,N_17066);
nor U17485 (N_17485,N_16957,N_17119);
or U17486 (N_17486,N_17121,N_17030);
and U17487 (N_17487,N_17018,N_17147);
and U17488 (N_17488,N_17105,N_16867);
nor U17489 (N_17489,N_16895,N_17181);
and U17490 (N_17490,N_17170,N_17123);
or U17491 (N_17491,N_17174,N_16999);
or U17492 (N_17492,N_16824,N_16811);
or U17493 (N_17493,N_16904,N_16846);
and U17494 (N_17494,N_16946,N_17044);
nand U17495 (N_17495,N_16855,N_16896);
or U17496 (N_17496,N_16814,N_17001);
and U17497 (N_17497,N_16993,N_16889);
and U17498 (N_17498,N_17045,N_16874);
nor U17499 (N_17499,N_17089,N_17046);
nor U17500 (N_17500,N_17178,N_17053);
or U17501 (N_17501,N_16838,N_16997);
or U17502 (N_17502,N_17089,N_17131);
nor U17503 (N_17503,N_17036,N_17038);
nor U17504 (N_17504,N_17028,N_16917);
nand U17505 (N_17505,N_17198,N_16985);
and U17506 (N_17506,N_16873,N_17079);
and U17507 (N_17507,N_17092,N_16951);
or U17508 (N_17508,N_16902,N_17110);
nor U17509 (N_17509,N_16872,N_16852);
or U17510 (N_17510,N_17113,N_16967);
nand U17511 (N_17511,N_17189,N_17088);
or U17512 (N_17512,N_16911,N_17121);
nand U17513 (N_17513,N_17142,N_17113);
nand U17514 (N_17514,N_17000,N_16851);
or U17515 (N_17515,N_17084,N_17060);
nand U17516 (N_17516,N_17106,N_17086);
nand U17517 (N_17517,N_17099,N_17111);
and U17518 (N_17518,N_16898,N_17051);
nand U17519 (N_17519,N_17049,N_16898);
nand U17520 (N_17520,N_16980,N_17065);
and U17521 (N_17521,N_17188,N_16836);
or U17522 (N_17522,N_16923,N_16936);
and U17523 (N_17523,N_16908,N_17135);
nand U17524 (N_17524,N_16914,N_17178);
nor U17525 (N_17525,N_16923,N_16895);
nand U17526 (N_17526,N_16830,N_16972);
or U17527 (N_17527,N_17151,N_17015);
nor U17528 (N_17528,N_16912,N_16985);
or U17529 (N_17529,N_17071,N_16886);
nor U17530 (N_17530,N_17043,N_17041);
nor U17531 (N_17531,N_17153,N_16947);
or U17532 (N_17532,N_17129,N_17113);
or U17533 (N_17533,N_16953,N_17064);
or U17534 (N_17534,N_16830,N_17070);
or U17535 (N_17535,N_17163,N_16900);
nor U17536 (N_17536,N_16882,N_17040);
nor U17537 (N_17537,N_16947,N_17119);
nand U17538 (N_17538,N_16826,N_16989);
nand U17539 (N_17539,N_17184,N_16893);
and U17540 (N_17540,N_16847,N_17124);
or U17541 (N_17541,N_17052,N_16957);
and U17542 (N_17542,N_16813,N_16859);
nand U17543 (N_17543,N_17088,N_16975);
nand U17544 (N_17544,N_16988,N_17096);
or U17545 (N_17545,N_16849,N_17041);
nand U17546 (N_17546,N_17024,N_17180);
nor U17547 (N_17547,N_16926,N_17058);
nor U17548 (N_17548,N_16970,N_16807);
nand U17549 (N_17549,N_16898,N_16983);
nand U17550 (N_17550,N_17073,N_17061);
nor U17551 (N_17551,N_16805,N_16816);
and U17552 (N_17552,N_17046,N_17132);
and U17553 (N_17553,N_17123,N_17193);
nor U17554 (N_17554,N_17175,N_17177);
nand U17555 (N_17555,N_17054,N_16970);
nand U17556 (N_17556,N_16997,N_16989);
nand U17557 (N_17557,N_16994,N_16904);
or U17558 (N_17558,N_16870,N_16988);
or U17559 (N_17559,N_16984,N_16888);
and U17560 (N_17560,N_16994,N_17014);
nand U17561 (N_17561,N_17164,N_17012);
or U17562 (N_17562,N_16936,N_16893);
nand U17563 (N_17563,N_16815,N_16923);
and U17564 (N_17564,N_16890,N_17089);
and U17565 (N_17565,N_16931,N_17002);
and U17566 (N_17566,N_16876,N_17104);
and U17567 (N_17567,N_17016,N_17141);
or U17568 (N_17568,N_17114,N_17042);
and U17569 (N_17569,N_17133,N_16894);
or U17570 (N_17570,N_16930,N_17144);
and U17571 (N_17571,N_16902,N_16817);
and U17572 (N_17572,N_16843,N_17003);
nor U17573 (N_17573,N_17025,N_16853);
or U17574 (N_17574,N_17068,N_16962);
nand U17575 (N_17575,N_17067,N_17199);
nor U17576 (N_17576,N_16972,N_17096);
and U17577 (N_17577,N_17150,N_17120);
and U17578 (N_17578,N_16872,N_16830);
or U17579 (N_17579,N_17122,N_17028);
and U17580 (N_17580,N_17168,N_16850);
or U17581 (N_17581,N_16857,N_17014);
or U17582 (N_17582,N_17185,N_17186);
and U17583 (N_17583,N_16994,N_17071);
or U17584 (N_17584,N_17157,N_16908);
and U17585 (N_17585,N_16884,N_17071);
nand U17586 (N_17586,N_17015,N_17164);
nor U17587 (N_17587,N_16823,N_17073);
nand U17588 (N_17588,N_16989,N_16942);
nand U17589 (N_17589,N_17006,N_17135);
nor U17590 (N_17590,N_16856,N_16985);
and U17591 (N_17591,N_17070,N_17089);
nor U17592 (N_17592,N_16838,N_16915);
nor U17593 (N_17593,N_17197,N_17119);
nand U17594 (N_17594,N_16810,N_17108);
nor U17595 (N_17595,N_17028,N_16924);
and U17596 (N_17596,N_16848,N_17056);
or U17597 (N_17597,N_16914,N_16961);
and U17598 (N_17598,N_17134,N_16833);
nand U17599 (N_17599,N_16842,N_16849);
nand U17600 (N_17600,N_17348,N_17429);
and U17601 (N_17601,N_17545,N_17587);
and U17602 (N_17602,N_17302,N_17365);
nand U17603 (N_17603,N_17237,N_17398);
nor U17604 (N_17604,N_17564,N_17327);
xnor U17605 (N_17605,N_17571,N_17406);
and U17606 (N_17606,N_17464,N_17479);
or U17607 (N_17607,N_17596,N_17289);
nor U17608 (N_17608,N_17534,N_17377);
nand U17609 (N_17609,N_17450,N_17583);
nand U17610 (N_17610,N_17238,N_17259);
nand U17611 (N_17611,N_17514,N_17345);
and U17612 (N_17612,N_17267,N_17498);
nand U17613 (N_17613,N_17561,N_17355);
nor U17614 (N_17614,N_17559,N_17414);
and U17615 (N_17615,N_17352,N_17445);
and U17616 (N_17616,N_17402,N_17469);
nand U17617 (N_17617,N_17536,N_17550);
nand U17618 (N_17618,N_17547,N_17428);
or U17619 (N_17619,N_17552,N_17364);
or U17620 (N_17620,N_17509,N_17463);
or U17621 (N_17621,N_17217,N_17490);
or U17622 (N_17622,N_17443,N_17255);
nand U17623 (N_17623,N_17439,N_17412);
nand U17624 (N_17624,N_17314,N_17307);
nand U17625 (N_17625,N_17465,N_17395);
nor U17626 (N_17626,N_17310,N_17529);
nor U17627 (N_17627,N_17320,N_17366);
or U17628 (N_17628,N_17535,N_17339);
and U17629 (N_17629,N_17495,N_17342);
nor U17630 (N_17630,N_17591,N_17388);
and U17631 (N_17631,N_17321,N_17408);
or U17632 (N_17632,N_17472,N_17375);
and U17633 (N_17633,N_17417,N_17525);
or U17634 (N_17634,N_17542,N_17353);
nand U17635 (N_17635,N_17354,N_17248);
and U17636 (N_17636,N_17523,N_17367);
and U17637 (N_17637,N_17585,N_17549);
and U17638 (N_17638,N_17218,N_17383);
nor U17639 (N_17639,N_17319,N_17329);
and U17640 (N_17640,N_17462,N_17501);
or U17641 (N_17641,N_17249,N_17309);
nor U17642 (N_17642,N_17566,N_17347);
or U17643 (N_17643,N_17568,N_17297);
nand U17644 (N_17644,N_17234,N_17210);
or U17645 (N_17645,N_17468,N_17291);
nor U17646 (N_17646,N_17563,N_17477);
nor U17647 (N_17647,N_17504,N_17203);
and U17648 (N_17648,N_17569,N_17332);
or U17649 (N_17649,N_17376,N_17539);
and U17650 (N_17650,N_17546,N_17356);
nor U17651 (N_17651,N_17260,N_17500);
or U17652 (N_17652,N_17494,N_17308);
nor U17653 (N_17653,N_17460,N_17499);
and U17654 (N_17654,N_17516,N_17415);
or U17655 (N_17655,N_17251,N_17598);
or U17656 (N_17656,N_17374,N_17244);
nor U17657 (N_17657,N_17437,N_17225);
nor U17658 (N_17658,N_17577,N_17593);
nor U17659 (N_17659,N_17502,N_17432);
and U17660 (N_17660,N_17590,N_17470);
and U17661 (N_17661,N_17527,N_17278);
and U17662 (N_17662,N_17396,N_17215);
nand U17663 (N_17663,N_17394,N_17294);
or U17664 (N_17664,N_17341,N_17497);
and U17665 (N_17665,N_17492,N_17584);
nor U17666 (N_17666,N_17474,N_17457);
nand U17667 (N_17667,N_17452,N_17228);
nand U17668 (N_17668,N_17476,N_17390);
or U17669 (N_17669,N_17288,N_17455);
nand U17670 (N_17670,N_17325,N_17493);
nor U17671 (N_17671,N_17287,N_17524);
or U17672 (N_17672,N_17243,N_17200);
and U17673 (N_17673,N_17335,N_17570);
or U17674 (N_17674,N_17360,N_17491);
nor U17675 (N_17675,N_17338,N_17592);
nor U17676 (N_17676,N_17433,N_17544);
and U17677 (N_17677,N_17232,N_17485);
nand U17678 (N_17678,N_17382,N_17481);
and U17679 (N_17679,N_17368,N_17370);
nor U17680 (N_17680,N_17265,N_17580);
and U17681 (N_17681,N_17480,N_17317);
nand U17682 (N_17682,N_17451,N_17594);
nor U17683 (N_17683,N_17206,N_17252);
and U17684 (N_17684,N_17286,N_17582);
nand U17685 (N_17685,N_17540,N_17576);
and U17686 (N_17686,N_17344,N_17334);
nor U17687 (N_17687,N_17373,N_17358);
and U17688 (N_17688,N_17558,N_17475);
nor U17689 (N_17689,N_17586,N_17386);
nand U17690 (N_17690,N_17236,N_17211);
and U17691 (N_17691,N_17467,N_17221);
nand U17692 (N_17692,N_17471,N_17579);
nor U17693 (N_17693,N_17324,N_17446);
or U17694 (N_17694,N_17240,N_17487);
nor U17695 (N_17695,N_17220,N_17515);
nand U17696 (N_17696,N_17254,N_17283);
nor U17697 (N_17697,N_17336,N_17279);
nor U17698 (N_17698,N_17262,N_17526);
nor U17699 (N_17699,N_17424,N_17557);
nor U17700 (N_17700,N_17316,N_17213);
nor U17701 (N_17701,N_17548,N_17397);
nand U17702 (N_17702,N_17410,N_17484);
xor U17703 (N_17703,N_17303,N_17538);
or U17704 (N_17704,N_17298,N_17513);
or U17705 (N_17705,N_17226,N_17407);
and U17706 (N_17706,N_17510,N_17223);
nor U17707 (N_17707,N_17507,N_17253);
nand U17708 (N_17708,N_17290,N_17459);
nor U17709 (N_17709,N_17263,N_17567);
and U17710 (N_17710,N_17553,N_17519);
and U17711 (N_17711,N_17378,N_17266);
or U17712 (N_17712,N_17456,N_17560);
and U17713 (N_17713,N_17400,N_17436);
or U17714 (N_17714,N_17554,N_17482);
nor U17715 (N_17715,N_17242,N_17430);
nor U17716 (N_17716,N_17207,N_17573);
or U17717 (N_17717,N_17268,N_17328);
nor U17718 (N_17718,N_17361,N_17280);
and U17719 (N_17719,N_17276,N_17293);
xnor U17720 (N_17720,N_17209,N_17421);
nor U17721 (N_17721,N_17229,N_17512);
or U17722 (N_17722,N_17532,N_17247);
nand U17723 (N_17723,N_17274,N_17387);
nand U17724 (N_17724,N_17305,N_17322);
or U17725 (N_17725,N_17277,N_17447);
nand U17726 (N_17726,N_17261,N_17216);
nand U17727 (N_17727,N_17426,N_17438);
nand U17728 (N_17728,N_17311,N_17299);
nor U17729 (N_17729,N_17541,N_17588);
nand U17730 (N_17730,N_17312,N_17363);
nand U17731 (N_17731,N_17423,N_17343);
or U17732 (N_17732,N_17489,N_17401);
nor U17733 (N_17733,N_17359,N_17533);
and U17734 (N_17734,N_17454,N_17440);
nand U17735 (N_17735,N_17503,N_17201);
nand U17736 (N_17736,N_17292,N_17449);
or U17737 (N_17737,N_17425,N_17420);
and U17738 (N_17738,N_17511,N_17337);
or U17739 (N_17739,N_17372,N_17530);
nor U17740 (N_17740,N_17486,N_17441);
nand U17741 (N_17741,N_17369,N_17349);
nor U17742 (N_17742,N_17304,N_17257);
or U17743 (N_17743,N_17380,N_17589);
nand U17744 (N_17744,N_17379,N_17371);
nor U17745 (N_17745,N_17250,N_17435);
nand U17746 (N_17746,N_17381,N_17416);
nor U17747 (N_17747,N_17403,N_17224);
nor U17748 (N_17748,N_17434,N_17409);
nor U17749 (N_17749,N_17208,N_17281);
or U17750 (N_17750,N_17340,N_17357);
or U17751 (N_17751,N_17442,N_17362);
nor U17752 (N_17752,N_17230,N_17419);
or U17753 (N_17753,N_17543,N_17488);
nor U17754 (N_17754,N_17574,N_17405);
nand U17755 (N_17755,N_17264,N_17528);
nor U17756 (N_17756,N_17326,N_17385);
nor U17757 (N_17757,N_17202,N_17306);
nor U17758 (N_17758,N_17595,N_17296);
or U17759 (N_17759,N_17205,N_17565);
or U17760 (N_17760,N_17246,N_17496);
or U17761 (N_17761,N_17575,N_17453);
and U17762 (N_17762,N_17473,N_17521);
nor U17763 (N_17763,N_17422,N_17241);
nor U17764 (N_17764,N_17517,N_17413);
nand U17765 (N_17765,N_17418,N_17214);
nor U17766 (N_17766,N_17458,N_17531);
nand U17767 (N_17767,N_17331,N_17333);
nor U17768 (N_17768,N_17384,N_17391);
nor U17769 (N_17769,N_17204,N_17245);
nor U17770 (N_17770,N_17285,N_17346);
or U17771 (N_17771,N_17555,N_17315);
xor U17772 (N_17772,N_17508,N_17404);
nand U17773 (N_17773,N_17227,N_17239);
or U17774 (N_17774,N_17284,N_17448);
nand U17775 (N_17775,N_17295,N_17258);
and U17776 (N_17776,N_17212,N_17269);
nor U17777 (N_17777,N_17222,N_17466);
or U17778 (N_17778,N_17256,N_17578);
and U17779 (N_17779,N_17461,N_17444);
and U17780 (N_17780,N_17478,N_17551);
or U17781 (N_17781,N_17505,N_17483);
nand U17782 (N_17782,N_17520,N_17597);
nor U17783 (N_17783,N_17282,N_17537);
nor U17784 (N_17784,N_17522,N_17351);
and U17785 (N_17785,N_17330,N_17411);
or U17786 (N_17786,N_17270,N_17273);
nand U17787 (N_17787,N_17318,N_17572);
or U17788 (N_17788,N_17389,N_17300);
nand U17789 (N_17789,N_17233,N_17350);
or U17790 (N_17790,N_17581,N_17323);
xor U17791 (N_17791,N_17393,N_17271);
or U17792 (N_17792,N_17313,N_17431);
nor U17793 (N_17793,N_17556,N_17301);
nor U17794 (N_17794,N_17599,N_17562);
nor U17795 (N_17795,N_17399,N_17275);
nor U17796 (N_17796,N_17235,N_17518);
nand U17797 (N_17797,N_17506,N_17427);
or U17798 (N_17798,N_17392,N_17272);
nor U17799 (N_17799,N_17231,N_17219);
xor U17800 (N_17800,N_17532,N_17374);
nand U17801 (N_17801,N_17522,N_17354);
and U17802 (N_17802,N_17390,N_17598);
nor U17803 (N_17803,N_17438,N_17332);
nand U17804 (N_17804,N_17430,N_17414);
nand U17805 (N_17805,N_17325,N_17336);
or U17806 (N_17806,N_17310,N_17493);
and U17807 (N_17807,N_17315,N_17422);
nand U17808 (N_17808,N_17430,N_17483);
or U17809 (N_17809,N_17588,N_17413);
and U17810 (N_17810,N_17480,N_17590);
nand U17811 (N_17811,N_17307,N_17312);
and U17812 (N_17812,N_17223,N_17394);
and U17813 (N_17813,N_17541,N_17524);
or U17814 (N_17814,N_17307,N_17519);
nor U17815 (N_17815,N_17348,N_17322);
nor U17816 (N_17816,N_17496,N_17432);
nor U17817 (N_17817,N_17471,N_17415);
and U17818 (N_17818,N_17485,N_17468);
and U17819 (N_17819,N_17288,N_17219);
nor U17820 (N_17820,N_17467,N_17264);
nand U17821 (N_17821,N_17493,N_17574);
nor U17822 (N_17822,N_17225,N_17204);
and U17823 (N_17823,N_17483,N_17401);
or U17824 (N_17824,N_17394,N_17308);
nor U17825 (N_17825,N_17310,N_17484);
and U17826 (N_17826,N_17375,N_17541);
nor U17827 (N_17827,N_17461,N_17357);
and U17828 (N_17828,N_17405,N_17450);
nand U17829 (N_17829,N_17559,N_17260);
nand U17830 (N_17830,N_17232,N_17482);
nand U17831 (N_17831,N_17307,N_17551);
nor U17832 (N_17832,N_17530,N_17569);
nor U17833 (N_17833,N_17560,N_17570);
and U17834 (N_17834,N_17323,N_17282);
nand U17835 (N_17835,N_17440,N_17340);
nor U17836 (N_17836,N_17596,N_17283);
or U17837 (N_17837,N_17245,N_17390);
and U17838 (N_17838,N_17215,N_17498);
and U17839 (N_17839,N_17443,N_17547);
or U17840 (N_17840,N_17240,N_17349);
or U17841 (N_17841,N_17216,N_17408);
nor U17842 (N_17842,N_17333,N_17229);
nor U17843 (N_17843,N_17442,N_17204);
nor U17844 (N_17844,N_17358,N_17507);
and U17845 (N_17845,N_17297,N_17356);
nand U17846 (N_17846,N_17481,N_17350);
nand U17847 (N_17847,N_17235,N_17230);
nand U17848 (N_17848,N_17408,N_17591);
or U17849 (N_17849,N_17506,N_17369);
or U17850 (N_17850,N_17258,N_17450);
nor U17851 (N_17851,N_17329,N_17546);
and U17852 (N_17852,N_17557,N_17497);
and U17853 (N_17853,N_17322,N_17331);
nor U17854 (N_17854,N_17213,N_17384);
or U17855 (N_17855,N_17209,N_17215);
or U17856 (N_17856,N_17480,N_17415);
nor U17857 (N_17857,N_17596,N_17243);
or U17858 (N_17858,N_17251,N_17445);
and U17859 (N_17859,N_17515,N_17510);
nor U17860 (N_17860,N_17433,N_17591);
and U17861 (N_17861,N_17267,N_17306);
nor U17862 (N_17862,N_17410,N_17214);
nor U17863 (N_17863,N_17401,N_17351);
or U17864 (N_17864,N_17450,N_17508);
or U17865 (N_17865,N_17550,N_17369);
xor U17866 (N_17866,N_17219,N_17277);
or U17867 (N_17867,N_17552,N_17492);
nand U17868 (N_17868,N_17449,N_17374);
or U17869 (N_17869,N_17274,N_17351);
or U17870 (N_17870,N_17265,N_17371);
or U17871 (N_17871,N_17237,N_17463);
and U17872 (N_17872,N_17338,N_17535);
nor U17873 (N_17873,N_17322,N_17430);
or U17874 (N_17874,N_17455,N_17468);
and U17875 (N_17875,N_17209,N_17236);
nor U17876 (N_17876,N_17470,N_17500);
or U17877 (N_17877,N_17397,N_17336);
nor U17878 (N_17878,N_17588,N_17437);
and U17879 (N_17879,N_17559,N_17360);
or U17880 (N_17880,N_17450,N_17482);
nor U17881 (N_17881,N_17434,N_17483);
and U17882 (N_17882,N_17447,N_17305);
nor U17883 (N_17883,N_17490,N_17267);
nand U17884 (N_17884,N_17228,N_17201);
or U17885 (N_17885,N_17235,N_17569);
or U17886 (N_17886,N_17295,N_17347);
nor U17887 (N_17887,N_17534,N_17384);
or U17888 (N_17888,N_17283,N_17301);
and U17889 (N_17889,N_17292,N_17387);
and U17890 (N_17890,N_17401,N_17588);
or U17891 (N_17891,N_17359,N_17409);
nor U17892 (N_17892,N_17506,N_17334);
nor U17893 (N_17893,N_17530,N_17538);
and U17894 (N_17894,N_17267,N_17477);
nor U17895 (N_17895,N_17571,N_17216);
nand U17896 (N_17896,N_17206,N_17336);
and U17897 (N_17897,N_17442,N_17488);
or U17898 (N_17898,N_17311,N_17340);
or U17899 (N_17899,N_17304,N_17560);
nor U17900 (N_17900,N_17518,N_17254);
or U17901 (N_17901,N_17266,N_17315);
or U17902 (N_17902,N_17560,N_17384);
or U17903 (N_17903,N_17501,N_17546);
or U17904 (N_17904,N_17206,N_17544);
xnor U17905 (N_17905,N_17491,N_17523);
or U17906 (N_17906,N_17549,N_17357);
nor U17907 (N_17907,N_17224,N_17584);
and U17908 (N_17908,N_17417,N_17212);
nor U17909 (N_17909,N_17595,N_17500);
nor U17910 (N_17910,N_17255,N_17519);
or U17911 (N_17911,N_17278,N_17234);
or U17912 (N_17912,N_17428,N_17350);
and U17913 (N_17913,N_17465,N_17581);
nor U17914 (N_17914,N_17484,N_17255);
or U17915 (N_17915,N_17295,N_17266);
nand U17916 (N_17916,N_17413,N_17572);
and U17917 (N_17917,N_17316,N_17553);
and U17918 (N_17918,N_17537,N_17272);
nand U17919 (N_17919,N_17553,N_17472);
nand U17920 (N_17920,N_17261,N_17457);
and U17921 (N_17921,N_17278,N_17480);
or U17922 (N_17922,N_17337,N_17462);
nand U17923 (N_17923,N_17263,N_17301);
xnor U17924 (N_17924,N_17531,N_17295);
or U17925 (N_17925,N_17532,N_17275);
nand U17926 (N_17926,N_17528,N_17237);
nor U17927 (N_17927,N_17397,N_17532);
and U17928 (N_17928,N_17403,N_17222);
nand U17929 (N_17929,N_17566,N_17440);
and U17930 (N_17930,N_17357,N_17365);
nor U17931 (N_17931,N_17400,N_17576);
and U17932 (N_17932,N_17366,N_17297);
or U17933 (N_17933,N_17491,N_17552);
nor U17934 (N_17934,N_17258,N_17332);
nand U17935 (N_17935,N_17427,N_17531);
nor U17936 (N_17936,N_17382,N_17507);
or U17937 (N_17937,N_17249,N_17507);
and U17938 (N_17938,N_17248,N_17576);
nand U17939 (N_17939,N_17217,N_17524);
nand U17940 (N_17940,N_17292,N_17259);
and U17941 (N_17941,N_17400,N_17524);
and U17942 (N_17942,N_17280,N_17552);
and U17943 (N_17943,N_17380,N_17284);
or U17944 (N_17944,N_17480,N_17533);
nand U17945 (N_17945,N_17331,N_17381);
and U17946 (N_17946,N_17204,N_17327);
nor U17947 (N_17947,N_17303,N_17427);
nand U17948 (N_17948,N_17256,N_17553);
and U17949 (N_17949,N_17308,N_17252);
nand U17950 (N_17950,N_17396,N_17392);
nor U17951 (N_17951,N_17295,N_17298);
and U17952 (N_17952,N_17422,N_17283);
nor U17953 (N_17953,N_17325,N_17429);
or U17954 (N_17954,N_17394,N_17257);
and U17955 (N_17955,N_17492,N_17290);
nor U17956 (N_17956,N_17567,N_17278);
nand U17957 (N_17957,N_17366,N_17313);
or U17958 (N_17958,N_17415,N_17200);
nor U17959 (N_17959,N_17441,N_17211);
nor U17960 (N_17960,N_17596,N_17360);
or U17961 (N_17961,N_17323,N_17435);
and U17962 (N_17962,N_17393,N_17562);
or U17963 (N_17963,N_17387,N_17205);
or U17964 (N_17964,N_17366,N_17432);
and U17965 (N_17965,N_17215,N_17574);
nor U17966 (N_17966,N_17328,N_17249);
and U17967 (N_17967,N_17449,N_17430);
or U17968 (N_17968,N_17408,N_17362);
or U17969 (N_17969,N_17277,N_17304);
nor U17970 (N_17970,N_17379,N_17370);
nor U17971 (N_17971,N_17352,N_17334);
and U17972 (N_17972,N_17293,N_17587);
and U17973 (N_17973,N_17577,N_17564);
or U17974 (N_17974,N_17535,N_17491);
nor U17975 (N_17975,N_17212,N_17346);
and U17976 (N_17976,N_17220,N_17504);
nor U17977 (N_17977,N_17371,N_17217);
nand U17978 (N_17978,N_17343,N_17379);
nand U17979 (N_17979,N_17379,N_17447);
and U17980 (N_17980,N_17436,N_17264);
or U17981 (N_17981,N_17437,N_17507);
or U17982 (N_17982,N_17455,N_17249);
nand U17983 (N_17983,N_17222,N_17211);
nand U17984 (N_17984,N_17348,N_17236);
nor U17985 (N_17985,N_17411,N_17299);
nand U17986 (N_17986,N_17298,N_17269);
xor U17987 (N_17987,N_17317,N_17411);
nor U17988 (N_17988,N_17245,N_17243);
or U17989 (N_17989,N_17281,N_17569);
or U17990 (N_17990,N_17522,N_17591);
nor U17991 (N_17991,N_17444,N_17532);
nor U17992 (N_17992,N_17470,N_17369);
nand U17993 (N_17993,N_17408,N_17499);
nor U17994 (N_17994,N_17434,N_17347);
or U17995 (N_17995,N_17308,N_17336);
and U17996 (N_17996,N_17315,N_17551);
nor U17997 (N_17997,N_17217,N_17408);
nor U17998 (N_17998,N_17597,N_17499);
nor U17999 (N_17999,N_17226,N_17228);
or U18000 (N_18000,N_17652,N_17782);
nor U18001 (N_18001,N_17962,N_17663);
and U18002 (N_18002,N_17786,N_17928);
nand U18003 (N_18003,N_17708,N_17628);
nand U18004 (N_18004,N_17697,N_17722);
or U18005 (N_18005,N_17727,N_17830);
or U18006 (N_18006,N_17760,N_17668);
nor U18007 (N_18007,N_17993,N_17709);
or U18008 (N_18008,N_17702,N_17989);
and U18009 (N_18009,N_17891,N_17968);
or U18010 (N_18010,N_17673,N_17689);
and U18011 (N_18011,N_17634,N_17821);
nor U18012 (N_18012,N_17649,N_17792);
or U18013 (N_18013,N_17600,N_17864);
nand U18014 (N_18014,N_17982,N_17753);
nand U18015 (N_18015,N_17909,N_17633);
nand U18016 (N_18016,N_17677,N_17806);
nor U18017 (N_18017,N_17808,N_17761);
or U18018 (N_18018,N_17882,N_17904);
or U18019 (N_18019,N_17738,N_17755);
and U18020 (N_18020,N_17720,N_17903);
nor U18021 (N_18021,N_17701,N_17953);
nand U18022 (N_18022,N_17839,N_17878);
nor U18023 (N_18023,N_17818,N_17721);
xnor U18024 (N_18024,N_17898,N_17840);
or U18025 (N_18025,N_17921,N_17960);
nor U18026 (N_18026,N_17790,N_17667);
nand U18027 (N_18027,N_17674,N_17912);
nor U18028 (N_18028,N_17813,N_17876);
and U18029 (N_18029,N_17712,N_17682);
and U18030 (N_18030,N_17672,N_17883);
nor U18031 (N_18031,N_17774,N_17662);
nand U18032 (N_18032,N_17926,N_17620);
nor U18033 (N_18033,N_17841,N_17857);
and U18034 (N_18034,N_17829,N_17935);
and U18035 (N_18035,N_17804,N_17739);
and U18036 (N_18036,N_17811,N_17743);
nor U18037 (N_18037,N_17868,N_17884);
and U18038 (N_18038,N_17779,N_17713);
or U18039 (N_18039,N_17601,N_17836);
or U18040 (N_18040,N_17852,N_17759);
nor U18041 (N_18041,N_17837,N_17966);
nand U18042 (N_18042,N_17951,N_17723);
nor U18043 (N_18043,N_17687,N_17715);
nand U18044 (N_18044,N_17606,N_17870);
nor U18045 (N_18045,N_17736,N_17660);
and U18046 (N_18046,N_17608,N_17783);
nand U18047 (N_18047,N_17793,N_17819);
or U18048 (N_18048,N_17932,N_17843);
nand U18049 (N_18049,N_17825,N_17653);
and U18050 (N_18050,N_17860,N_17645);
nand U18051 (N_18051,N_17627,N_17844);
and U18052 (N_18052,N_17916,N_17820);
or U18053 (N_18053,N_17970,N_17719);
or U18054 (N_18054,N_17675,N_17958);
nand U18055 (N_18055,N_17855,N_17861);
and U18056 (N_18056,N_17906,N_17805);
or U18057 (N_18057,N_17763,N_17975);
or U18058 (N_18058,N_17936,N_17987);
or U18059 (N_18059,N_17748,N_17872);
nand U18060 (N_18060,N_17914,N_17895);
nand U18061 (N_18061,N_17991,N_17661);
and U18062 (N_18062,N_17611,N_17940);
nand U18063 (N_18063,N_17803,N_17671);
nor U18064 (N_18064,N_17937,N_17776);
or U18065 (N_18065,N_17901,N_17961);
and U18066 (N_18066,N_17828,N_17886);
and U18067 (N_18067,N_17616,N_17703);
and U18068 (N_18068,N_17866,N_17648);
or U18069 (N_18069,N_17605,N_17724);
nand U18070 (N_18070,N_17874,N_17758);
or U18071 (N_18071,N_17983,N_17676);
nor U18072 (N_18072,N_17955,N_17918);
and U18073 (N_18073,N_17642,N_17771);
nor U18074 (N_18074,N_17740,N_17757);
and U18075 (N_18075,N_17607,N_17623);
or U18076 (N_18076,N_17698,N_17964);
nor U18077 (N_18077,N_17917,N_17665);
nand U18078 (N_18078,N_17603,N_17777);
or U18079 (N_18079,N_17969,N_17859);
and U18080 (N_18080,N_17899,N_17659);
and U18081 (N_18081,N_17988,N_17832);
nor U18082 (N_18082,N_17833,N_17907);
nor U18083 (N_18083,N_17683,N_17746);
nor U18084 (N_18084,N_17822,N_17920);
and U18085 (N_18085,N_17716,N_17871);
nand U18086 (N_18086,N_17831,N_17775);
nand U18087 (N_18087,N_17944,N_17690);
nand U18088 (N_18088,N_17826,N_17700);
or U18089 (N_18089,N_17963,N_17930);
nor U18090 (N_18090,N_17824,N_17629);
nor U18091 (N_18091,N_17744,N_17880);
and U18092 (N_18092,N_17950,N_17934);
nor U18093 (N_18093,N_17990,N_17902);
nand U18094 (N_18094,N_17992,N_17887);
and U18095 (N_18095,N_17796,N_17762);
and U18096 (N_18096,N_17637,N_17794);
or U18097 (N_18097,N_17952,N_17905);
or U18098 (N_18098,N_17994,N_17681);
or U18099 (N_18099,N_17823,N_17881);
or U18100 (N_18100,N_17625,N_17707);
nand U18101 (N_18101,N_17609,N_17965);
or U18102 (N_18102,N_17849,N_17893);
or U18103 (N_18103,N_17696,N_17635);
nor U18104 (N_18104,N_17730,N_17706);
nor U18105 (N_18105,N_17945,N_17853);
nor U18106 (N_18106,N_17725,N_17985);
nor U18107 (N_18107,N_17984,N_17734);
nand U18108 (N_18108,N_17630,N_17910);
nand U18109 (N_18109,N_17741,N_17834);
nand U18110 (N_18110,N_17956,N_17856);
nand U18111 (N_18111,N_17613,N_17612);
nor U18112 (N_18112,N_17638,N_17997);
nand U18113 (N_18113,N_17971,N_17919);
and U18114 (N_18114,N_17655,N_17657);
nand U18115 (N_18115,N_17685,N_17737);
nor U18116 (N_18116,N_17892,N_17717);
and U18117 (N_18117,N_17908,N_17654);
nor U18118 (N_18118,N_17631,N_17924);
nand U18119 (N_18119,N_17889,N_17764);
nand U18120 (N_18120,N_17646,N_17851);
or U18121 (N_18121,N_17827,N_17810);
or U18122 (N_18122,N_17943,N_17797);
or U18123 (N_18123,N_17941,N_17888);
and U18124 (N_18124,N_17948,N_17896);
and U18125 (N_18125,N_17778,N_17981);
and U18126 (N_18126,N_17699,N_17614);
or U18127 (N_18127,N_17604,N_17694);
and U18128 (N_18128,N_17704,N_17858);
nand U18129 (N_18129,N_17789,N_17767);
nor U18130 (N_18130,N_17729,N_17726);
nor U18131 (N_18131,N_17766,N_17626);
and U18132 (N_18132,N_17974,N_17897);
nor U18133 (N_18133,N_17747,N_17666);
nand U18134 (N_18134,N_17817,N_17848);
nand U18135 (N_18135,N_17765,N_17754);
nand U18136 (N_18136,N_17877,N_17954);
nor U18137 (N_18137,N_17756,N_17807);
nor U18138 (N_18138,N_17610,N_17996);
nor U18139 (N_18139,N_17885,N_17732);
nand U18140 (N_18140,N_17618,N_17742);
and U18141 (N_18141,N_17647,N_17999);
or U18142 (N_18142,N_17927,N_17802);
nor U18143 (N_18143,N_17768,N_17800);
and U18144 (N_18144,N_17602,N_17879);
nor U18145 (N_18145,N_17938,N_17693);
nor U18146 (N_18146,N_17745,N_17711);
and U18147 (N_18147,N_17890,N_17986);
or U18148 (N_18148,N_17644,N_17735);
nor U18149 (N_18149,N_17731,N_17939);
nand U18150 (N_18150,N_17998,N_17769);
and U18151 (N_18151,N_17773,N_17925);
nor U18152 (N_18152,N_17845,N_17816);
nor U18153 (N_18153,N_17695,N_17842);
nor U18154 (N_18154,N_17915,N_17619);
nand U18155 (N_18155,N_17705,N_17641);
or U18156 (N_18156,N_17894,N_17976);
and U18157 (N_18157,N_17809,N_17980);
or U18158 (N_18158,N_17733,N_17664);
and U18159 (N_18159,N_17617,N_17632);
nand U18160 (N_18160,N_17781,N_17650);
and U18161 (N_18161,N_17995,N_17780);
nand U18162 (N_18162,N_17949,N_17639);
nor U18163 (N_18163,N_17622,N_17656);
and U18164 (N_18164,N_17798,N_17770);
or U18165 (N_18165,N_17752,N_17847);
and U18166 (N_18166,N_17815,N_17791);
nand U18167 (N_18167,N_17913,N_17801);
nor U18168 (N_18168,N_17692,N_17863);
or U18169 (N_18169,N_17957,N_17850);
or U18170 (N_18170,N_17710,N_17787);
and U18171 (N_18171,N_17688,N_17788);
or U18172 (N_18172,N_17862,N_17942);
or U18173 (N_18173,N_17749,N_17865);
nor U18174 (N_18174,N_17947,N_17691);
or U18175 (N_18175,N_17911,N_17799);
nand U18176 (N_18176,N_17679,N_17669);
nor U18177 (N_18177,N_17651,N_17977);
and U18178 (N_18178,N_17978,N_17873);
and U18179 (N_18179,N_17838,N_17875);
nor U18180 (N_18180,N_17624,N_17946);
or U18181 (N_18181,N_17785,N_17686);
nand U18182 (N_18182,N_17922,N_17979);
and U18183 (N_18183,N_17636,N_17795);
nand U18184 (N_18184,N_17973,N_17714);
and U18185 (N_18185,N_17835,N_17929);
or U18186 (N_18186,N_17923,N_17670);
or U18187 (N_18187,N_17728,N_17854);
nand U18188 (N_18188,N_17621,N_17684);
and U18189 (N_18189,N_17750,N_17846);
nand U18190 (N_18190,N_17972,N_17643);
nand U18191 (N_18191,N_17967,N_17718);
nor U18192 (N_18192,N_17812,N_17867);
and U18193 (N_18193,N_17933,N_17640);
nand U18194 (N_18194,N_17931,N_17900);
nor U18195 (N_18195,N_17772,N_17680);
nand U18196 (N_18196,N_17814,N_17678);
or U18197 (N_18197,N_17869,N_17959);
nor U18198 (N_18198,N_17784,N_17751);
and U18199 (N_18199,N_17658,N_17615);
and U18200 (N_18200,N_17815,N_17713);
and U18201 (N_18201,N_17756,N_17641);
nand U18202 (N_18202,N_17906,N_17708);
nor U18203 (N_18203,N_17719,N_17936);
nor U18204 (N_18204,N_17975,N_17848);
and U18205 (N_18205,N_17835,N_17666);
nor U18206 (N_18206,N_17651,N_17690);
nand U18207 (N_18207,N_17787,N_17650);
nand U18208 (N_18208,N_17606,N_17897);
nand U18209 (N_18209,N_17628,N_17926);
and U18210 (N_18210,N_17911,N_17661);
and U18211 (N_18211,N_17638,N_17813);
nor U18212 (N_18212,N_17815,N_17968);
and U18213 (N_18213,N_17648,N_17610);
and U18214 (N_18214,N_17869,N_17779);
nand U18215 (N_18215,N_17841,N_17720);
nor U18216 (N_18216,N_17946,N_17824);
or U18217 (N_18217,N_17739,N_17802);
nor U18218 (N_18218,N_17693,N_17645);
or U18219 (N_18219,N_17747,N_17681);
or U18220 (N_18220,N_17738,N_17832);
nand U18221 (N_18221,N_17781,N_17633);
or U18222 (N_18222,N_17863,N_17641);
nand U18223 (N_18223,N_17692,N_17678);
nor U18224 (N_18224,N_17905,N_17887);
nor U18225 (N_18225,N_17912,N_17808);
nor U18226 (N_18226,N_17607,N_17863);
and U18227 (N_18227,N_17980,N_17647);
and U18228 (N_18228,N_17843,N_17604);
or U18229 (N_18229,N_17728,N_17680);
nand U18230 (N_18230,N_17634,N_17921);
nand U18231 (N_18231,N_17674,N_17672);
or U18232 (N_18232,N_17941,N_17875);
nor U18233 (N_18233,N_17971,N_17967);
nand U18234 (N_18234,N_17769,N_17745);
nor U18235 (N_18235,N_17896,N_17964);
nor U18236 (N_18236,N_17682,N_17678);
nor U18237 (N_18237,N_17863,N_17892);
nand U18238 (N_18238,N_17668,N_17624);
nand U18239 (N_18239,N_17625,N_17626);
and U18240 (N_18240,N_17752,N_17907);
and U18241 (N_18241,N_17919,N_17946);
or U18242 (N_18242,N_17713,N_17756);
nand U18243 (N_18243,N_17752,N_17987);
nor U18244 (N_18244,N_17980,N_17699);
or U18245 (N_18245,N_17928,N_17935);
nor U18246 (N_18246,N_17888,N_17815);
nor U18247 (N_18247,N_17628,N_17904);
and U18248 (N_18248,N_17624,N_17688);
or U18249 (N_18249,N_17765,N_17648);
nand U18250 (N_18250,N_17824,N_17627);
nand U18251 (N_18251,N_17634,N_17612);
and U18252 (N_18252,N_17808,N_17703);
or U18253 (N_18253,N_17669,N_17883);
or U18254 (N_18254,N_17818,N_17840);
or U18255 (N_18255,N_17621,N_17971);
and U18256 (N_18256,N_17766,N_17882);
and U18257 (N_18257,N_17662,N_17959);
and U18258 (N_18258,N_17964,N_17880);
and U18259 (N_18259,N_17902,N_17985);
nand U18260 (N_18260,N_17603,N_17697);
and U18261 (N_18261,N_17985,N_17745);
or U18262 (N_18262,N_17763,N_17605);
nand U18263 (N_18263,N_17857,N_17723);
and U18264 (N_18264,N_17819,N_17614);
nand U18265 (N_18265,N_17926,N_17799);
and U18266 (N_18266,N_17952,N_17668);
or U18267 (N_18267,N_17858,N_17968);
nor U18268 (N_18268,N_17927,N_17934);
nand U18269 (N_18269,N_17846,N_17635);
nand U18270 (N_18270,N_17815,N_17842);
nand U18271 (N_18271,N_17635,N_17795);
nor U18272 (N_18272,N_17644,N_17957);
nor U18273 (N_18273,N_17995,N_17683);
nand U18274 (N_18274,N_17716,N_17897);
nor U18275 (N_18275,N_17984,N_17992);
or U18276 (N_18276,N_17847,N_17893);
or U18277 (N_18277,N_17898,N_17659);
nand U18278 (N_18278,N_17971,N_17922);
nand U18279 (N_18279,N_17813,N_17981);
nor U18280 (N_18280,N_17874,N_17614);
or U18281 (N_18281,N_17620,N_17928);
nand U18282 (N_18282,N_17879,N_17856);
nor U18283 (N_18283,N_17968,N_17913);
or U18284 (N_18284,N_17640,N_17998);
nand U18285 (N_18285,N_17960,N_17876);
and U18286 (N_18286,N_17720,N_17881);
nor U18287 (N_18287,N_17608,N_17729);
and U18288 (N_18288,N_17857,N_17839);
nor U18289 (N_18289,N_17701,N_17784);
or U18290 (N_18290,N_17792,N_17914);
nor U18291 (N_18291,N_17956,N_17732);
nor U18292 (N_18292,N_17795,N_17756);
or U18293 (N_18293,N_17751,N_17798);
nand U18294 (N_18294,N_17792,N_17628);
and U18295 (N_18295,N_17774,N_17976);
nor U18296 (N_18296,N_17938,N_17782);
and U18297 (N_18297,N_17677,N_17611);
nor U18298 (N_18298,N_17625,N_17781);
or U18299 (N_18299,N_17673,N_17908);
or U18300 (N_18300,N_17867,N_17821);
or U18301 (N_18301,N_17745,N_17720);
nor U18302 (N_18302,N_17873,N_17966);
nor U18303 (N_18303,N_17775,N_17663);
or U18304 (N_18304,N_17886,N_17682);
nor U18305 (N_18305,N_17669,N_17831);
nor U18306 (N_18306,N_17851,N_17672);
and U18307 (N_18307,N_17733,N_17886);
nand U18308 (N_18308,N_17793,N_17668);
xnor U18309 (N_18309,N_17774,N_17654);
and U18310 (N_18310,N_17733,N_17632);
and U18311 (N_18311,N_17775,N_17758);
or U18312 (N_18312,N_17631,N_17673);
nor U18313 (N_18313,N_17809,N_17975);
nor U18314 (N_18314,N_17645,N_17912);
and U18315 (N_18315,N_17847,N_17795);
or U18316 (N_18316,N_17925,N_17755);
or U18317 (N_18317,N_17757,N_17822);
nor U18318 (N_18318,N_17905,N_17769);
and U18319 (N_18319,N_17840,N_17843);
nand U18320 (N_18320,N_17816,N_17620);
nand U18321 (N_18321,N_17892,N_17899);
xnor U18322 (N_18322,N_17714,N_17854);
nor U18323 (N_18323,N_17979,N_17810);
nor U18324 (N_18324,N_17611,N_17659);
or U18325 (N_18325,N_17832,N_17927);
nor U18326 (N_18326,N_17610,N_17932);
and U18327 (N_18327,N_17831,N_17845);
nand U18328 (N_18328,N_17748,N_17643);
nor U18329 (N_18329,N_17993,N_17706);
and U18330 (N_18330,N_17679,N_17645);
or U18331 (N_18331,N_17783,N_17944);
or U18332 (N_18332,N_17872,N_17916);
nand U18333 (N_18333,N_17670,N_17759);
nand U18334 (N_18334,N_17822,N_17712);
or U18335 (N_18335,N_17621,N_17788);
or U18336 (N_18336,N_17966,N_17714);
nand U18337 (N_18337,N_17990,N_17826);
and U18338 (N_18338,N_17988,N_17624);
and U18339 (N_18339,N_17960,N_17679);
and U18340 (N_18340,N_17603,N_17713);
or U18341 (N_18341,N_17633,N_17699);
and U18342 (N_18342,N_17937,N_17849);
and U18343 (N_18343,N_17687,N_17825);
nand U18344 (N_18344,N_17970,N_17677);
and U18345 (N_18345,N_17786,N_17930);
nor U18346 (N_18346,N_17880,N_17941);
nor U18347 (N_18347,N_17987,N_17604);
nand U18348 (N_18348,N_17657,N_17777);
and U18349 (N_18349,N_17896,N_17894);
nand U18350 (N_18350,N_17650,N_17880);
nand U18351 (N_18351,N_17895,N_17821);
nand U18352 (N_18352,N_17804,N_17915);
nor U18353 (N_18353,N_17689,N_17888);
nor U18354 (N_18354,N_17954,N_17838);
nor U18355 (N_18355,N_17743,N_17646);
nand U18356 (N_18356,N_17749,N_17800);
nor U18357 (N_18357,N_17833,N_17617);
or U18358 (N_18358,N_17919,N_17893);
and U18359 (N_18359,N_17988,N_17987);
nor U18360 (N_18360,N_17639,N_17662);
and U18361 (N_18361,N_17966,N_17826);
nor U18362 (N_18362,N_17643,N_17998);
xor U18363 (N_18363,N_17870,N_17628);
nor U18364 (N_18364,N_17834,N_17692);
or U18365 (N_18365,N_17908,N_17918);
nor U18366 (N_18366,N_17804,N_17647);
nand U18367 (N_18367,N_17909,N_17689);
nand U18368 (N_18368,N_17936,N_17868);
nor U18369 (N_18369,N_17858,N_17725);
nor U18370 (N_18370,N_17848,N_17831);
nor U18371 (N_18371,N_17613,N_17667);
nand U18372 (N_18372,N_17654,N_17943);
or U18373 (N_18373,N_17847,N_17933);
nor U18374 (N_18374,N_17758,N_17937);
or U18375 (N_18375,N_17616,N_17774);
xor U18376 (N_18376,N_17751,N_17806);
nand U18377 (N_18377,N_17929,N_17937);
or U18378 (N_18378,N_17934,N_17683);
and U18379 (N_18379,N_17841,N_17782);
or U18380 (N_18380,N_17766,N_17643);
nor U18381 (N_18381,N_17696,N_17885);
and U18382 (N_18382,N_17921,N_17988);
or U18383 (N_18383,N_17697,N_17653);
and U18384 (N_18384,N_17648,N_17842);
nand U18385 (N_18385,N_17627,N_17836);
or U18386 (N_18386,N_17684,N_17715);
and U18387 (N_18387,N_17878,N_17851);
or U18388 (N_18388,N_17860,N_17715);
nor U18389 (N_18389,N_17770,N_17935);
nand U18390 (N_18390,N_17917,N_17602);
and U18391 (N_18391,N_17922,N_17751);
nand U18392 (N_18392,N_17869,N_17875);
or U18393 (N_18393,N_17735,N_17976);
nand U18394 (N_18394,N_17819,N_17655);
nor U18395 (N_18395,N_17861,N_17989);
nand U18396 (N_18396,N_17788,N_17707);
or U18397 (N_18397,N_17756,N_17851);
nor U18398 (N_18398,N_17997,N_17680);
nand U18399 (N_18399,N_17609,N_17927);
nor U18400 (N_18400,N_18326,N_18209);
nand U18401 (N_18401,N_18039,N_18134);
and U18402 (N_18402,N_18100,N_18375);
nor U18403 (N_18403,N_18170,N_18069);
and U18404 (N_18404,N_18009,N_18362);
nor U18405 (N_18405,N_18080,N_18276);
and U18406 (N_18406,N_18171,N_18353);
or U18407 (N_18407,N_18366,N_18393);
nand U18408 (N_18408,N_18186,N_18245);
nand U18409 (N_18409,N_18242,N_18260);
nand U18410 (N_18410,N_18157,N_18236);
nor U18411 (N_18411,N_18004,N_18056);
nand U18412 (N_18412,N_18101,N_18371);
and U18413 (N_18413,N_18088,N_18113);
or U18414 (N_18414,N_18002,N_18399);
and U18415 (N_18415,N_18062,N_18099);
or U18416 (N_18416,N_18051,N_18094);
nand U18417 (N_18417,N_18067,N_18047);
or U18418 (N_18418,N_18241,N_18279);
nor U18419 (N_18419,N_18141,N_18177);
or U18420 (N_18420,N_18304,N_18104);
and U18421 (N_18421,N_18087,N_18060);
nor U18422 (N_18422,N_18125,N_18078);
or U18423 (N_18423,N_18187,N_18312);
or U18424 (N_18424,N_18015,N_18131);
and U18425 (N_18425,N_18129,N_18194);
and U18426 (N_18426,N_18050,N_18331);
nor U18427 (N_18427,N_18149,N_18109);
and U18428 (N_18428,N_18003,N_18359);
and U18429 (N_18429,N_18289,N_18382);
and U18430 (N_18430,N_18354,N_18226);
nor U18431 (N_18431,N_18044,N_18280);
nand U18432 (N_18432,N_18302,N_18182);
nor U18433 (N_18433,N_18300,N_18019);
nor U18434 (N_18434,N_18085,N_18025);
nor U18435 (N_18435,N_18152,N_18268);
or U18436 (N_18436,N_18369,N_18398);
or U18437 (N_18437,N_18223,N_18073);
and U18438 (N_18438,N_18159,N_18224);
nor U18439 (N_18439,N_18204,N_18107);
nor U18440 (N_18440,N_18063,N_18328);
nor U18441 (N_18441,N_18266,N_18197);
nor U18442 (N_18442,N_18074,N_18017);
nand U18443 (N_18443,N_18330,N_18077);
nor U18444 (N_18444,N_18337,N_18255);
nor U18445 (N_18445,N_18325,N_18285);
and U18446 (N_18446,N_18365,N_18263);
and U18447 (N_18447,N_18052,N_18161);
or U18448 (N_18448,N_18158,N_18195);
xnor U18449 (N_18449,N_18291,N_18035);
or U18450 (N_18450,N_18167,N_18173);
nor U18451 (N_18451,N_18207,N_18090);
nand U18452 (N_18452,N_18251,N_18225);
and U18453 (N_18453,N_18007,N_18174);
nand U18454 (N_18454,N_18306,N_18023);
or U18455 (N_18455,N_18299,N_18054);
or U18456 (N_18456,N_18313,N_18228);
or U18457 (N_18457,N_18361,N_18321);
nor U18458 (N_18458,N_18165,N_18079);
or U18459 (N_18459,N_18234,N_18189);
nand U18460 (N_18460,N_18130,N_18388);
nand U18461 (N_18461,N_18114,N_18033);
nor U18462 (N_18462,N_18272,N_18075);
nor U18463 (N_18463,N_18363,N_18091);
nand U18464 (N_18464,N_18380,N_18386);
or U18465 (N_18465,N_18309,N_18335);
or U18466 (N_18466,N_18132,N_18348);
nor U18467 (N_18467,N_18217,N_18237);
or U18468 (N_18468,N_18083,N_18200);
and U18469 (N_18469,N_18316,N_18305);
nor U18470 (N_18470,N_18324,N_18274);
or U18471 (N_18471,N_18180,N_18253);
nor U18472 (N_18472,N_18258,N_18153);
nor U18473 (N_18473,N_18288,N_18095);
nand U18474 (N_18474,N_18367,N_18198);
nor U18475 (N_18475,N_18344,N_18112);
and U18476 (N_18476,N_18277,N_18061);
or U18477 (N_18477,N_18168,N_18201);
nand U18478 (N_18478,N_18093,N_18188);
or U18479 (N_18479,N_18036,N_18137);
nor U18480 (N_18480,N_18133,N_18127);
or U18481 (N_18481,N_18227,N_18357);
or U18482 (N_18482,N_18287,N_18249);
or U18483 (N_18483,N_18281,N_18084);
nor U18484 (N_18484,N_18065,N_18105);
nand U18485 (N_18485,N_18163,N_18071);
nand U18486 (N_18486,N_18038,N_18257);
and U18487 (N_18487,N_18292,N_18097);
nand U18488 (N_18488,N_18142,N_18081);
and U18489 (N_18489,N_18164,N_18179);
nor U18490 (N_18490,N_18111,N_18233);
or U18491 (N_18491,N_18307,N_18252);
and U18492 (N_18492,N_18058,N_18117);
or U18493 (N_18493,N_18203,N_18322);
nand U18494 (N_18494,N_18246,N_18191);
nand U18495 (N_18495,N_18301,N_18356);
or U18496 (N_18496,N_18351,N_18219);
or U18497 (N_18497,N_18270,N_18028);
nand U18498 (N_18498,N_18368,N_18243);
nand U18499 (N_18499,N_18218,N_18310);
nand U18500 (N_18500,N_18064,N_18210);
nor U18501 (N_18501,N_18381,N_18118);
nand U18502 (N_18502,N_18096,N_18121);
nand U18503 (N_18503,N_18024,N_18010);
nand U18504 (N_18504,N_18333,N_18184);
nand U18505 (N_18505,N_18394,N_18146);
or U18506 (N_18506,N_18046,N_18384);
nor U18507 (N_18507,N_18372,N_18072);
nor U18508 (N_18508,N_18150,N_18254);
nor U18509 (N_18509,N_18396,N_18021);
nand U18510 (N_18510,N_18139,N_18001);
or U18511 (N_18511,N_18323,N_18123);
nand U18512 (N_18512,N_18031,N_18042);
and U18513 (N_18513,N_18190,N_18145);
nand U18514 (N_18514,N_18136,N_18143);
and U18515 (N_18515,N_18032,N_18378);
nand U18516 (N_18516,N_18278,N_18317);
nor U18517 (N_18517,N_18108,N_18314);
or U18518 (N_18518,N_18346,N_18284);
xnor U18519 (N_18519,N_18259,N_18140);
nand U18520 (N_18520,N_18012,N_18379);
or U18521 (N_18521,N_18162,N_18048);
and U18522 (N_18522,N_18208,N_18282);
nor U18523 (N_18523,N_18205,N_18053);
and U18524 (N_18524,N_18068,N_18193);
or U18525 (N_18525,N_18026,N_18397);
nor U18526 (N_18526,N_18342,N_18119);
and U18527 (N_18527,N_18387,N_18202);
nor U18528 (N_18528,N_18269,N_18120);
or U18529 (N_18529,N_18235,N_18247);
nand U18530 (N_18530,N_18290,N_18156);
nand U18531 (N_18531,N_18338,N_18350);
nand U18532 (N_18532,N_18320,N_18057);
or U18533 (N_18533,N_18041,N_18347);
or U18534 (N_18534,N_18303,N_18006);
nor U18535 (N_18535,N_18261,N_18176);
nand U18536 (N_18536,N_18192,N_18030);
or U18537 (N_18537,N_18345,N_18102);
xnor U18538 (N_18538,N_18395,N_18206);
or U18539 (N_18539,N_18144,N_18358);
nor U18540 (N_18540,N_18327,N_18373);
nor U18541 (N_18541,N_18391,N_18339);
xor U18542 (N_18542,N_18390,N_18374);
and U18543 (N_18543,N_18016,N_18283);
and U18544 (N_18544,N_18175,N_18089);
or U18545 (N_18545,N_18250,N_18213);
nor U18546 (N_18546,N_18154,N_18298);
nor U18547 (N_18547,N_18264,N_18181);
nor U18548 (N_18548,N_18221,N_18018);
or U18549 (N_18549,N_18138,N_18318);
and U18550 (N_18550,N_18238,N_18011);
nor U18551 (N_18551,N_18066,N_18037);
nor U18552 (N_18552,N_18343,N_18240);
nand U18553 (N_18553,N_18352,N_18020);
nand U18554 (N_18554,N_18349,N_18148);
or U18555 (N_18555,N_18022,N_18248);
nand U18556 (N_18556,N_18124,N_18212);
nand U18557 (N_18557,N_18014,N_18059);
and U18558 (N_18558,N_18286,N_18049);
or U18559 (N_18559,N_18329,N_18392);
nor U18560 (N_18560,N_18055,N_18334);
nand U18561 (N_18561,N_18000,N_18256);
nand U18562 (N_18562,N_18013,N_18332);
or U18563 (N_18563,N_18377,N_18043);
nand U18564 (N_18564,N_18040,N_18103);
nand U18565 (N_18565,N_18360,N_18106);
or U18566 (N_18566,N_18244,N_18172);
and U18567 (N_18567,N_18222,N_18151);
nand U18568 (N_18568,N_18383,N_18385);
and U18569 (N_18569,N_18370,N_18045);
and U18570 (N_18570,N_18389,N_18265);
nand U18571 (N_18571,N_18214,N_18110);
nand U18572 (N_18572,N_18147,N_18216);
and U18573 (N_18573,N_18178,N_18169);
nand U18574 (N_18574,N_18271,N_18295);
and U18575 (N_18575,N_18092,N_18294);
nand U18576 (N_18576,N_18308,N_18376);
nand U18577 (N_18577,N_18355,N_18166);
or U18578 (N_18578,N_18183,N_18275);
and U18579 (N_18579,N_18199,N_18341);
nand U18580 (N_18580,N_18315,N_18070);
nand U18581 (N_18581,N_18196,N_18160);
nand U18582 (N_18582,N_18034,N_18311);
nor U18583 (N_18583,N_18293,N_18116);
nand U18584 (N_18584,N_18336,N_18082);
nor U18585 (N_18585,N_18267,N_18220);
or U18586 (N_18586,N_18364,N_18005);
nor U18587 (N_18587,N_18122,N_18231);
nand U18588 (N_18588,N_18296,N_18076);
nor U18589 (N_18589,N_18230,N_18297);
or U18590 (N_18590,N_18098,N_18155);
or U18591 (N_18591,N_18185,N_18008);
nor U18592 (N_18592,N_18029,N_18239);
nand U18593 (N_18593,N_18115,N_18215);
nand U18594 (N_18594,N_18126,N_18229);
or U18595 (N_18595,N_18211,N_18128);
nand U18596 (N_18596,N_18027,N_18232);
nand U18597 (N_18597,N_18273,N_18319);
or U18598 (N_18598,N_18135,N_18340);
and U18599 (N_18599,N_18086,N_18262);
nor U18600 (N_18600,N_18347,N_18214);
nor U18601 (N_18601,N_18089,N_18058);
nor U18602 (N_18602,N_18247,N_18136);
nand U18603 (N_18603,N_18393,N_18200);
nand U18604 (N_18604,N_18134,N_18056);
and U18605 (N_18605,N_18215,N_18394);
nor U18606 (N_18606,N_18056,N_18026);
or U18607 (N_18607,N_18094,N_18289);
and U18608 (N_18608,N_18396,N_18052);
and U18609 (N_18609,N_18058,N_18294);
nand U18610 (N_18610,N_18244,N_18248);
nor U18611 (N_18611,N_18342,N_18009);
nor U18612 (N_18612,N_18186,N_18238);
nor U18613 (N_18613,N_18333,N_18221);
and U18614 (N_18614,N_18321,N_18181);
and U18615 (N_18615,N_18148,N_18165);
and U18616 (N_18616,N_18137,N_18076);
nand U18617 (N_18617,N_18360,N_18036);
nand U18618 (N_18618,N_18261,N_18154);
nand U18619 (N_18619,N_18065,N_18388);
or U18620 (N_18620,N_18209,N_18293);
and U18621 (N_18621,N_18026,N_18036);
nand U18622 (N_18622,N_18260,N_18107);
or U18623 (N_18623,N_18064,N_18233);
nand U18624 (N_18624,N_18158,N_18179);
nor U18625 (N_18625,N_18283,N_18093);
or U18626 (N_18626,N_18292,N_18399);
xor U18627 (N_18627,N_18187,N_18151);
nand U18628 (N_18628,N_18113,N_18381);
nand U18629 (N_18629,N_18275,N_18145);
nand U18630 (N_18630,N_18053,N_18027);
nand U18631 (N_18631,N_18310,N_18292);
nand U18632 (N_18632,N_18044,N_18301);
nor U18633 (N_18633,N_18125,N_18155);
nor U18634 (N_18634,N_18053,N_18200);
or U18635 (N_18635,N_18220,N_18297);
nand U18636 (N_18636,N_18072,N_18125);
or U18637 (N_18637,N_18342,N_18168);
and U18638 (N_18638,N_18206,N_18174);
and U18639 (N_18639,N_18342,N_18366);
or U18640 (N_18640,N_18307,N_18232);
or U18641 (N_18641,N_18354,N_18134);
or U18642 (N_18642,N_18201,N_18131);
or U18643 (N_18643,N_18019,N_18326);
nand U18644 (N_18644,N_18017,N_18131);
nand U18645 (N_18645,N_18365,N_18177);
nor U18646 (N_18646,N_18169,N_18002);
or U18647 (N_18647,N_18193,N_18039);
nor U18648 (N_18648,N_18362,N_18231);
or U18649 (N_18649,N_18392,N_18238);
nand U18650 (N_18650,N_18286,N_18111);
or U18651 (N_18651,N_18078,N_18301);
nor U18652 (N_18652,N_18127,N_18088);
nor U18653 (N_18653,N_18010,N_18133);
nor U18654 (N_18654,N_18187,N_18321);
and U18655 (N_18655,N_18358,N_18189);
nor U18656 (N_18656,N_18173,N_18241);
nand U18657 (N_18657,N_18023,N_18006);
and U18658 (N_18658,N_18042,N_18268);
nand U18659 (N_18659,N_18268,N_18002);
nand U18660 (N_18660,N_18183,N_18058);
and U18661 (N_18661,N_18091,N_18383);
nor U18662 (N_18662,N_18172,N_18175);
and U18663 (N_18663,N_18033,N_18198);
nand U18664 (N_18664,N_18180,N_18313);
nor U18665 (N_18665,N_18347,N_18189);
nand U18666 (N_18666,N_18054,N_18053);
nand U18667 (N_18667,N_18004,N_18326);
nand U18668 (N_18668,N_18060,N_18088);
nor U18669 (N_18669,N_18250,N_18078);
xor U18670 (N_18670,N_18203,N_18275);
or U18671 (N_18671,N_18072,N_18325);
nand U18672 (N_18672,N_18037,N_18223);
and U18673 (N_18673,N_18369,N_18206);
and U18674 (N_18674,N_18298,N_18358);
or U18675 (N_18675,N_18383,N_18374);
nor U18676 (N_18676,N_18124,N_18274);
or U18677 (N_18677,N_18148,N_18357);
nor U18678 (N_18678,N_18296,N_18151);
nand U18679 (N_18679,N_18321,N_18371);
nor U18680 (N_18680,N_18083,N_18134);
and U18681 (N_18681,N_18189,N_18259);
and U18682 (N_18682,N_18347,N_18202);
nand U18683 (N_18683,N_18113,N_18234);
xnor U18684 (N_18684,N_18297,N_18068);
nor U18685 (N_18685,N_18290,N_18074);
nand U18686 (N_18686,N_18317,N_18359);
and U18687 (N_18687,N_18038,N_18085);
nand U18688 (N_18688,N_18373,N_18323);
and U18689 (N_18689,N_18285,N_18089);
or U18690 (N_18690,N_18095,N_18326);
nor U18691 (N_18691,N_18111,N_18121);
nand U18692 (N_18692,N_18359,N_18309);
and U18693 (N_18693,N_18142,N_18271);
and U18694 (N_18694,N_18398,N_18056);
nor U18695 (N_18695,N_18204,N_18329);
and U18696 (N_18696,N_18267,N_18043);
and U18697 (N_18697,N_18251,N_18044);
nor U18698 (N_18698,N_18007,N_18044);
nand U18699 (N_18699,N_18140,N_18020);
and U18700 (N_18700,N_18235,N_18180);
nor U18701 (N_18701,N_18363,N_18312);
and U18702 (N_18702,N_18233,N_18114);
nor U18703 (N_18703,N_18155,N_18048);
or U18704 (N_18704,N_18363,N_18196);
nand U18705 (N_18705,N_18167,N_18377);
and U18706 (N_18706,N_18385,N_18324);
nand U18707 (N_18707,N_18155,N_18180);
and U18708 (N_18708,N_18233,N_18065);
and U18709 (N_18709,N_18346,N_18331);
nor U18710 (N_18710,N_18079,N_18160);
nor U18711 (N_18711,N_18352,N_18024);
or U18712 (N_18712,N_18266,N_18198);
nand U18713 (N_18713,N_18164,N_18188);
or U18714 (N_18714,N_18037,N_18200);
nor U18715 (N_18715,N_18180,N_18244);
nor U18716 (N_18716,N_18214,N_18367);
or U18717 (N_18717,N_18239,N_18032);
or U18718 (N_18718,N_18179,N_18010);
nand U18719 (N_18719,N_18139,N_18026);
and U18720 (N_18720,N_18019,N_18373);
and U18721 (N_18721,N_18324,N_18122);
nand U18722 (N_18722,N_18184,N_18381);
or U18723 (N_18723,N_18352,N_18281);
nand U18724 (N_18724,N_18101,N_18004);
nand U18725 (N_18725,N_18184,N_18003);
nor U18726 (N_18726,N_18353,N_18106);
nor U18727 (N_18727,N_18371,N_18207);
or U18728 (N_18728,N_18204,N_18076);
nand U18729 (N_18729,N_18233,N_18272);
nor U18730 (N_18730,N_18326,N_18180);
nor U18731 (N_18731,N_18332,N_18204);
or U18732 (N_18732,N_18256,N_18138);
or U18733 (N_18733,N_18029,N_18191);
and U18734 (N_18734,N_18227,N_18326);
nand U18735 (N_18735,N_18244,N_18336);
nor U18736 (N_18736,N_18191,N_18042);
or U18737 (N_18737,N_18101,N_18130);
nor U18738 (N_18738,N_18120,N_18349);
nand U18739 (N_18739,N_18048,N_18043);
or U18740 (N_18740,N_18347,N_18343);
nor U18741 (N_18741,N_18161,N_18275);
nand U18742 (N_18742,N_18229,N_18360);
or U18743 (N_18743,N_18168,N_18226);
or U18744 (N_18744,N_18186,N_18284);
and U18745 (N_18745,N_18349,N_18295);
or U18746 (N_18746,N_18116,N_18095);
nand U18747 (N_18747,N_18321,N_18383);
and U18748 (N_18748,N_18021,N_18305);
nor U18749 (N_18749,N_18114,N_18398);
nor U18750 (N_18750,N_18221,N_18269);
or U18751 (N_18751,N_18103,N_18189);
and U18752 (N_18752,N_18155,N_18005);
nor U18753 (N_18753,N_18393,N_18182);
nand U18754 (N_18754,N_18019,N_18231);
nor U18755 (N_18755,N_18182,N_18312);
and U18756 (N_18756,N_18044,N_18330);
or U18757 (N_18757,N_18268,N_18107);
nand U18758 (N_18758,N_18223,N_18270);
nand U18759 (N_18759,N_18370,N_18157);
nor U18760 (N_18760,N_18388,N_18103);
xor U18761 (N_18761,N_18296,N_18320);
nor U18762 (N_18762,N_18302,N_18107);
and U18763 (N_18763,N_18138,N_18281);
or U18764 (N_18764,N_18285,N_18094);
nand U18765 (N_18765,N_18019,N_18122);
and U18766 (N_18766,N_18134,N_18125);
nand U18767 (N_18767,N_18194,N_18115);
nor U18768 (N_18768,N_18017,N_18309);
nand U18769 (N_18769,N_18257,N_18078);
nand U18770 (N_18770,N_18077,N_18396);
nor U18771 (N_18771,N_18134,N_18350);
nor U18772 (N_18772,N_18248,N_18075);
nor U18773 (N_18773,N_18059,N_18308);
or U18774 (N_18774,N_18181,N_18157);
nand U18775 (N_18775,N_18099,N_18037);
nor U18776 (N_18776,N_18233,N_18298);
and U18777 (N_18777,N_18184,N_18203);
and U18778 (N_18778,N_18353,N_18390);
or U18779 (N_18779,N_18299,N_18194);
nand U18780 (N_18780,N_18378,N_18109);
nand U18781 (N_18781,N_18278,N_18041);
and U18782 (N_18782,N_18097,N_18074);
and U18783 (N_18783,N_18006,N_18182);
nand U18784 (N_18784,N_18313,N_18164);
nor U18785 (N_18785,N_18333,N_18385);
nor U18786 (N_18786,N_18344,N_18045);
nand U18787 (N_18787,N_18355,N_18033);
or U18788 (N_18788,N_18315,N_18021);
nor U18789 (N_18789,N_18192,N_18281);
or U18790 (N_18790,N_18194,N_18144);
and U18791 (N_18791,N_18135,N_18010);
or U18792 (N_18792,N_18121,N_18244);
nand U18793 (N_18793,N_18366,N_18026);
and U18794 (N_18794,N_18265,N_18339);
nor U18795 (N_18795,N_18132,N_18258);
or U18796 (N_18796,N_18346,N_18326);
or U18797 (N_18797,N_18101,N_18344);
and U18798 (N_18798,N_18238,N_18385);
nor U18799 (N_18799,N_18115,N_18331);
nor U18800 (N_18800,N_18557,N_18493);
and U18801 (N_18801,N_18500,N_18470);
nor U18802 (N_18802,N_18647,N_18583);
or U18803 (N_18803,N_18764,N_18789);
or U18804 (N_18804,N_18637,N_18618);
nand U18805 (N_18805,N_18515,N_18722);
nand U18806 (N_18806,N_18437,N_18741);
and U18807 (N_18807,N_18656,N_18589);
nor U18808 (N_18808,N_18550,N_18695);
nand U18809 (N_18809,N_18621,N_18723);
and U18810 (N_18810,N_18428,N_18790);
or U18811 (N_18811,N_18766,N_18607);
and U18812 (N_18812,N_18592,N_18691);
or U18813 (N_18813,N_18672,N_18799);
nand U18814 (N_18814,N_18655,N_18420);
nor U18815 (N_18815,N_18675,N_18775);
and U18816 (N_18816,N_18599,N_18432);
and U18817 (N_18817,N_18536,N_18451);
nand U18818 (N_18818,N_18457,N_18732);
nor U18819 (N_18819,N_18733,N_18768);
nand U18820 (N_18820,N_18452,N_18664);
nand U18821 (N_18821,N_18495,N_18575);
nand U18822 (N_18822,N_18636,N_18702);
nor U18823 (N_18823,N_18716,N_18794);
or U18824 (N_18824,N_18605,N_18441);
and U18825 (N_18825,N_18415,N_18706);
nand U18826 (N_18826,N_18724,N_18552);
nand U18827 (N_18827,N_18458,N_18658);
nand U18828 (N_18828,N_18549,N_18507);
nor U18829 (N_18829,N_18701,N_18459);
or U18830 (N_18830,N_18753,N_18727);
nor U18831 (N_18831,N_18566,N_18491);
and U18832 (N_18832,N_18438,N_18760);
and U18833 (N_18833,N_18796,N_18631);
nand U18834 (N_18834,N_18523,N_18609);
and U18835 (N_18835,N_18781,N_18413);
nand U18836 (N_18836,N_18759,N_18795);
and U18837 (N_18837,N_18522,N_18612);
nand U18838 (N_18838,N_18628,N_18614);
or U18839 (N_18839,N_18496,N_18453);
and U18840 (N_18840,N_18662,N_18524);
and U18841 (N_18841,N_18471,N_18638);
or U18842 (N_18842,N_18719,N_18411);
or U18843 (N_18843,N_18676,N_18797);
or U18844 (N_18844,N_18551,N_18450);
or U18845 (N_18845,N_18418,N_18782);
or U18846 (N_18846,N_18620,N_18783);
nand U18847 (N_18847,N_18712,N_18624);
or U18848 (N_18848,N_18565,N_18731);
and U18849 (N_18849,N_18529,N_18689);
or U18850 (N_18850,N_18460,N_18475);
or U18851 (N_18851,N_18476,N_18761);
nand U18852 (N_18852,N_18544,N_18682);
or U18853 (N_18853,N_18641,N_18560);
or U18854 (N_18854,N_18633,N_18520);
and U18855 (N_18855,N_18651,N_18553);
nand U18856 (N_18856,N_18587,N_18663);
or U18857 (N_18857,N_18581,N_18506);
or U18858 (N_18858,N_18713,N_18464);
nor U18859 (N_18859,N_18516,N_18659);
and U18860 (N_18860,N_18585,N_18772);
nand U18861 (N_18861,N_18720,N_18499);
nand U18862 (N_18862,N_18410,N_18742);
and U18863 (N_18863,N_18472,N_18538);
nand U18864 (N_18864,N_18696,N_18674);
or U18865 (N_18865,N_18579,N_18673);
or U18866 (N_18866,N_18677,N_18517);
nor U18867 (N_18867,N_18617,N_18690);
or U18868 (N_18868,N_18700,N_18639);
and U18869 (N_18869,N_18632,N_18705);
nand U18870 (N_18870,N_18652,N_18462);
nor U18871 (N_18871,N_18660,N_18685);
and U18872 (N_18872,N_18667,N_18466);
or U18873 (N_18873,N_18449,N_18704);
nor U18874 (N_18874,N_18521,N_18447);
or U18875 (N_18875,N_18698,N_18755);
nand U18876 (N_18876,N_18431,N_18440);
nand U18877 (N_18877,N_18683,N_18433);
nand U18878 (N_18878,N_18519,N_18779);
and U18879 (N_18879,N_18750,N_18409);
nand U18880 (N_18880,N_18564,N_18444);
and U18881 (N_18881,N_18541,N_18773);
xor U18882 (N_18882,N_18613,N_18417);
and U18883 (N_18883,N_18518,N_18487);
nor U18884 (N_18884,N_18709,N_18615);
or U18885 (N_18885,N_18503,N_18535);
nor U18886 (N_18886,N_18558,N_18419);
and U18887 (N_18887,N_18545,N_18703);
nor U18888 (N_18888,N_18717,N_18527);
or U18889 (N_18889,N_18494,N_18769);
or U18890 (N_18890,N_18473,N_18714);
nand U18891 (N_18891,N_18665,N_18596);
xor U18892 (N_18892,N_18563,N_18534);
and U18893 (N_18893,N_18436,N_18569);
or U18894 (N_18894,N_18735,N_18671);
nor U18895 (N_18895,N_18505,N_18711);
nor U18896 (N_18896,N_18502,N_18467);
nor U18897 (N_18897,N_18582,N_18435);
and U18898 (N_18898,N_18559,N_18603);
and U18899 (N_18899,N_18679,N_18590);
nand U18900 (N_18900,N_18721,N_18478);
and U18901 (N_18901,N_18501,N_18424);
nand U18902 (N_18902,N_18623,N_18416);
or U18903 (N_18903,N_18758,N_18622);
nor U18904 (N_18904,N_18484,N_18481);
nand U18905 (N_18905,N_18606,N_18770);
nor U18906 (N_18906,N_18543,N_18497);
nand U18907 (N_18907,N_18403,N_18430);
nor U18908 (N_18908,N_18739,N_18412);
or U18909 (N_18909,N_18490,N_18697);
or U18910 (N_18910,N_18680,N_18454);
and U18911 (N_18911,N_18729,N_18474);
nor U18912 (N_18912,N_18530,N_18580);
or U18913 (N_18913,N_18743,N_18539);
or U18914 (N_18914,N_18602,N_18414);
or U18915 (N_18915,N_18608,N_18456);
and U18916 (N_18916,N_18598,N_18514);
or U18917 (N_18917,N_18600,N_18512);
or U18918 (N_18918,N_18648,N_18793);
nand U18919 (N_18919,N_18687,N_18640);
and U18920 (N_18920,N_18455,N_18747);
nand U18921 (N_18921,N_18528,N_18480);
or U18922 (N_18922,N_18445,N_18601);
or U18923 (N_18923,N_18771,N_18469);
nand U18924 (N_18924,N_18567,N_18798);
nor U18925 (N_18925,N_18785,N_18584);
and U18926 (N_18926,N_18571,N_18791);
and U18927 (N_18927,N_18461,N_18526);
or U18928 (N_18928,N_18692,N_18402);
nand U18929 (N_18929,N_18776,N_18630);
or U18930 (N_18930,N_18483,N_18562);
nand U18931 (N_18931,N_18792,N_18654);
or U18932 (N_18932,N_18588,N_18678);
and U18933 (N_18933,N_18407,N_18533);
or U18934 (N_18934,N_18572,N_18547);
or U18935 (N_18935,N_18684,N_18578);
nor U18936 (N_18936,N_18554,N_18477);
and U18937 (N_18937,N_18737,N_18668);
or U18938 (N_18938,N_18510,N_18486);
or U18939 (N_18939,N_18504,N_18763);
nor U18940 (N_18940,N_18446,N_18787);
nand U18941 (N_18941,N_18594,N_18754);
nor U18942 (N_18942,N_18540,N_18548);
or U18943 (N_18943,N_18670,N_18626);
nand U18944 (N_18944,N_18400,N_18492);
or U18945 (N_18945,N_18718,N_18489);
or U18946 (N_18946,N_18757,N_18784);
and U18947 (N_18947,N_18744,N_18734);
nor U18948 (N_18948,N_18650,N_18745);
or U18949 (N_18949,N_18555,N_18568);
and U18950 (N_18950,N_18644,N_18408);
nand U18951 (N_18951,N_18681,N_18710);
nand U18952 (N_18952,N_18748,N_18509);
nand U18953 (N_18953,N_18511,N_18715);
nor U18954 (N_18954,N_18746,N_18777);
xor U18955 (N_18955,N_18762,N_18767);
nand U18956 (N_18956,N_18556,N_18642);
and U18957 (N_18957,N_18405,N_18574);
nor U18958 (N_18958,N_18726,N_18422);
nor U18959 (N_18959,N_18774,N_18625);
nand U18960 (N_18960,N_18597,N_18669);
nor U18961 (N_18961,N_18423,N_18699);
nand U18962 (N_18962,N_18468,N_18482);
nor U18963 (N_18963,N_18661,N_18604);
nor U18964 (N_18964,N_18780,N_18573);
and U18965 (N_18965,N_18740,N_18421);
or U18966 (N_18966,N_18708,N_18629);
nand U18967 (N_18967,N_18646,N_18610);
and U18968 (N_18968,N_18751,N_18666);
or U18969 (N_18969,N_18593,N_18479);
nor U18970 (N_18970,N_18465,N_18730);
nand U18971 (N_18971,N_18765,N_18485);
nor U18972 (N_18972,N_18645,N_18439);
and U18973 (N_18973,N_18532,N_18649);
nand U18974 (N_18974,N_18404,N_18595);
nor U18975 (N_18975,N_18778,N_18756);
and U18976 (N_18976,N_18488,N_18707);
and U18977 (N_18977,N_18508,N_18448);
nor U18978 (N_18978,N_18738,N_18576);
or U18979 (N_18979,N_18643,N_18463);
or U18980 (N_18980,N_18694,N_18736);
or U18981 (N_18981,N_18611,N_18442);
or U18982 (N_18982,N_18786,N_18427);
nand U18983 (N_18983,N_18635,N_18443);
or U18984 (N_18984,N_18426,N_18513);
nand U18985 (N_18985,N_18725,N_18406);
nor U18986 (N_18986,N_18686,N_18570);
nor U18987 (N_18987,N_18619,N_18634);
or U18988 (N_18988,N_18591,N_18693);
or U18989 (N_18989,N_18429,N_18657);
or U18990 (N_18990,N_18728,N_18561);
nor U18991 (N_18991,N_18537,N_18788);
and U18992 (N_18992,N_18688,N_18425);
or U18993 (N_18993,N_18531,N_18542);
nand U18994 (N_18994,N_18586,N_18752);
xor U18995 (N_18995,N_18653,N_18546);
and U18996 (N_18996,N_18525,N_18616);
or U18997 (N_18997,N_18498,N_18401);
or U18998 (N_18998,N_18577,N_18749);
nand U18999 (N_18999,N_18434,N_18627);
nor U19000 (N_19000,N_18534,N_18642);
nand U19001 (N_19001,N_18499,N_18701);
or U19002 (N_19002,N_18743,N_18552);
nand U19003 (N_19003,N_18661,N_18578);
nor U19004 (N_19004,N_18781,N_18632);
nor U19005 (N_19005,N_18591,N_18466);
nor U19006 (N_19006,N_18743,N_18541);
or U19007 (N_19007,N_18776,N_18474);
nor U19008 (N_19008,N_18710,N_18421);
nand U19009 (N_19009,N_18686,N_18584);
or U19010 (N_19010,N_18696,N_18650);
nor U19011 (N_19011,N_18651,N_18610);
or U19012 (N_19012,N_18537,N_18576);
nand U19013 (N_19013,N_18443,N_18608);
or U19014 (N_19014,N_18572,N_18544);
or U19015 (N_19015,N_18506,N_18512);
nand U19016 (N_19016,N_18443,N_18469);
or U19017 (N_19017,N_18769,N_18644);
nand U19018 (N_19018,N_18738,N_18607);
and U19019 (N_19019,N_18573,N_18681);
nand U19020 (N_19020,N_18467,N_18622);
nand U19021 (N_19021,N_18739,N_18786);
or U19022 (N_19022,N_18744,N_18560);
nor U19023 (N_19023,N_18765,N_18650);
nand U19024 (N_19024,N_18552,N_18775);
and U19025 (N_19025,N_18746,N_18624);
nand U19026 (N_19026,N_18770,N_18443);
nand U19027 (N_19027,N_18687,N_18446);
and U19028 (N_19028,N_18470,N_18677);
or U19029 (N_19029,N_18513,N_18505);
nand U19030 (N_19030,N_18710,N_18587);
nand U19031 (N_19031,N_18581,N_18694);
or U19032 (N_19032,N_18485,N_18725);
or U19033 (N_19033,N_18634,N_18668);
and U19034 (N_19034,N_18447,N_18703);
or U19035 (N_19035,N_18605,N_18737);
or U19036 (N_19036,N_18758,N_18773);
or U19037 (N_19037,N_18703,N_18503);
nand U19038 (N_19038,N_18462,N_18749);
and U19039 (N_19039,N_18463,N_18674);
nor U19040 (N_19040,N_18733,N_18649);
nor U19041 (N_19041,N_18587,N_18688);
and U19042 (N_19042,N_18781,N_18663);
nor U19043 (N_19043,N_18690,N_18460);
nor U19044 (N_19044,N_18577,N_18786);
or U19045 (N_19045,N_18786,N_18524);
nor U19046 (N_19046,N_18775,N_18525);
or U19047 (N_19047,N_18630,N_18621);
nor U19048 (N_19048,N_18510,N_18533);
or U19049 (N_19049,N_18783,N_18472);
and U19050 (N_19050,N_18473,N_18539);
and U19051 (N_19051,N_18589,N_18684);
or U19052 (N_19052,N_18515,N_18429);
and U19053 (N_19053,N_18534,N_18654);
or U19054 (N_19054,N_18644,N_18666);
nand U19055 (N_19055,N_18690,N_18545);
or U19056 (N_19056,N_18689,N_18575);
and U19057 (N_19057,N_18759,N_18695);
and U19058 (N_19058,N_18488,N_18747);
nor U19059 (N_19059,N_18410,N_18535);
or U19060 (N_19060,N_18474,N_18645);
or U19061 (N_19061,N_18744,N_18426);
nand U19062 (N_19062,N_18797,N_18559);
and U19063 (N_19063,N_18633,N_18524);
nand U19064 (N_19064,N_18784,N_18609);
and U19065 (N_19065,N_18619,N_18756);
or U19066 (N_19066,N_18582,N_18790);
nand U19067 (N_19067,N_18475,N_18456);
or U19068 (N_19068,N_18412,N_18464);
nand U19069 (N_19069,N_18605,N_18683);
nand U19070 (N_19070,N_18486,N_18727);
nand U19071 (N_19071,N_18420,N_18553);
nor U19072 (N_19072,N_18591,N_18745);
nor U19073 (N_19073,N_18573,N_18586);
and U19074 (N_19074,N_18530,N_18402);
and U19075 (N_19075,N_18624,N_18718);
nor U19076 (N_19076,N_18511,N_18439);
nor U19077 (N_19077,N_18735,N_18652);
nand U19078 (N_19078,N_18690,N_18414);
nor U19079 (N_19079,N_18647,N_18694);
nor U19080 (N_19080,N_18628,N_18510);
nand U19081 (N_19081,N_18536,N_18760);
or U19082 (N_19082,N_18724,N_18670);
and U19083 (N_19083,N_18752,N_18680);
nand U19084 (N_19084,N_18646,N_18450);
and U19085 (N_19085,N_18527,N_18621);
nand U19086 (N_19086,N_18453,N_18745);
or U19087 (N_19087,N_18717,N_18611);
and U19088 (N_19088,N_18441,N_18470);
nor U19089 (N_19089,N_18563,N_18437);
and U19090 (N_19090,N_18620,N_18419);
nor U19091 (N_19091,N_18489,N_18746);
nor U19092 (N_19092,N_18665,N_18638);
or U19093 (N_19093,N_18653,N_18679);
nor U19094 (N_19094,N_18459,N_18575);
or U19095 (N_19095,N_18577,N_18591);
and U19096 (N_19096,N_18689,N_18486);
or U19097 (N_19097,N_18478,N_18524);
nand U19098 (N_19098,N_18602,N_18468);
nor U19099 (N_19099,N_18482,N_18444);
nand U19100 (N_19100,N_18654,N_18777);
nor U19101 (N_19101,N_18612,N_18705);
nor U19102 (N_19102,N_18527,N_18740);
nand U19103 (N_19103,N_18412,N_18666);
nand U19104 (N_19104,N_18786,N_18645);
nor U19105 (N_19105,N_18703,N_18543);
and U19106 (N_19106,N_18576,N_18485);
nand U19107 (N_19107,N_18462,N_18769);
nor U19108 (N_19108,N_18477,N_18416);
nand U19109 (N_19109,N_18413,N_18613);
or U19110 (N_19110,N_18678,N_18431);
nand U19111 (N_19111,N_18416,N_18439);
nand U19112 (N_19112,N_18605,N_18422);
xnor U19113 (N_19113,N_18708,N_18452);
xnor U19114 (N_19114,N_18717,N_18469);
or U19115 (N_19115,N_18603,N_18771);
nor U19116 (N_19116,N_18517,N_18595);
and U19117 (N_19117,N_18638,N_18718);
nor U19118 (N_19118,N_18549,N_18798);
nand U19119 (N_19119,N_18468,N_18494);
or U19120 (N_19120,N_18530,N_18536);
and U19121 (N_19121,N_18459,N_18753);
or U19122 (N_19122,N_18699,N_18593);
and U19123 (N_19123,N_18694,N_18661);
and U19124 (N_19124,N_18474,N_18439);
nand U19125 (N_19125,N_18536,N_18586);
nor U19126 (N_19126,N_18448,N_18400);
or U19127 (N_19127,N_18726,N_18667);
and U19128 (N_19128,N_18667,N_18658);
nor U19129 (N_19129,N_18569,N_18531);
nor U19130 (N_19130,N_18465,N_18587);
nor U19131 (N_19131,N_18555,N_18511);
nor U19132 (N_19132,N_18691,N_18427);
or U19133 (N_19133,N_18401,N_18766);
and U19134 (N_19134,N_18648,N_18677);
nor U19135 (N_19135,N_18671,N_18711);
nand U19136 (N_19136,N_18579,N_18545);
or U19137 (N_19137,N_18661,N_18642);
nand U19138 (N_19138,N_18416,N_18540);
or U19139 (N_19139,N_18758,N_18703);
and U19140 (N_19140,N_18721,N_18593);
or U19141 (N_19141,N_18757,N_18741);
nor U19142 (N_19142,N_18609,N_18619);
xor U19143 (N_19143,N_18631,N_18499);
nor U19144 (N_19144,N_18436,N_18613);
nand U19145 (N_19145,N_18615,N_18749);
nand U19146 (N_19146,N_18733,N_18556);
nand U19147 (N_19147,N_18624,N_18621);
nor U19148 (N_19148,N_18756,N_18493);
or U19149 (N_19149,N_18664,N_18551);
nand U19150 (N_19150,N_18768,N_18710);
nand U19151 (N_19151,N_18705,N_18684);
nor U19152 (N_19152,N_18684,N_18704);
and U19153 (N_19153,N_18718,N_18600);
nand U19154 (N_19154,N_18644,N_18720);
and U19155 (N_19155,N_18701,N_18559);
or U19156 (N_19156,N_18533,N_18599);
nand U19157 (N_19157,N_18418,N_18463);
nor U19158 (N_19158,N_18662,N_18502);
nand U19159 (N_19159,N_18445,N_18516);
or U19160 (N_19160,N_18544,N_18708);
and U19161 (N_19161,N_18615,N_18402);
nor U19162 (N_19162,N_18569,N_18592);
nand U19163 (N_19163,N_18463,N_18452);
and U19164 (N_19164,N_18787,N_18793);
nor U19165 (N_19165,N_18649,N_18589);
nand U19166 (N_19166,N_18681,N_18709);
and U19167 (N_19167,N_18526,N_18456);
nand U19168 (N_19168,N_18504,N_18450);
nand U19169 (N_19169,N_18535,N_18550);
nand U19170 (N_19170,N_18409,N_18505);
or U19171 (N_19171,N_18641,N_18672);
nor U19172 (N_19172,N_18763,N_18615);
nor U19173 (N_19173,N_18757,N_18732);
and U19174 (N_19174,N_18781,N_18571);
or U19175 (N_19175,N_18578,N_18778);
nand U19176 (N_19176,N_18689,N_18597);
nand U19177 (N_19177,N_18556,N_18741);
or U19178 (N_19178,N_18644,N_18401);
nor U19179 (N_19179,N_18681,N_18402);
nand U19180 (N_19180,N_18676,N_18519);
and U19181 (N_19181,N_18638,N_18409);
nand U19182 (N_19182,N_18531,N_18660);
and U19183 (N_19183,N_18526,N_18776);
or U19184 (N_19184,N_18590,N_18788);
or U19185 (N_19185,N_18647,N_18715);
and U19186 (N_19186,N_18423,N_18564);
nand U19187 (N_19187,N_18451,N_18771);
or U19188 (N_19188,N_18796,N_18740);
and U19189 (N_19189,N_18658,N_18759);
nand U19190 (N_19190,N_18494,N_18694);
nor U19191 (N_19191,N_18799,N_18594);
nor U19192 (N_19192,N_18724,N_18772);
or U19193 (N_19193,N_18781,N_18614);
nor U19194 (N_19194,N_18747,N_18637);
and U19195 (N_19195,N_18628,N_18737);
or U19196 (N_19196,N_18593,N_18701);
nor U19197 (N_19197,N_18427,N_18409);
or U19198 (N_19198,N_18643,N_18414);
or U19199 (N_19199,N_18675,N_18460);
or U19200 (N_19200,N_18916,N_18929);
nand U19201 (N_19201,N_18808,N_18823);
xor U19202 (N_19202,N_18947,N_19093);
and U19203 (N_19203,N_19025,N_19000);
nand U19204 (N_19204,N_19165,N_18937);
nand U19205 (N_19205,N_18858,N_18821);
and U19206 (N_19206,N_19113,N_18851);
and U19207 (N_19207,N_18822,N_18862);
and U19208 (N_19208,N_19037,N_19094);
or U19209 (N_19209,N_19177,N_18838);
nand U19210 (N_19210,N_18941,N_19073);
nand U19211 (N_19211,N_19072,N_19131);
nand U19212 (N_19212,N_19164,N_18870);
nand U19213 (N_19213,N_18807,N_19029);
nor U19214 (N_19214,N_18846,N_18918);
and U19215 (N_19215,N_19076,N_18969);
and U19216 (N_19216,N_18889,N_19035);
nand U19217 (N_19217,N_18897,N_18844);
or U19218 (N_19218,N_18886,N_18950);
nor U19219 (N_19219,N_18881,N_18917);
nand U19220 (N_19220,N_19122,N_19186);
and U19221 (N_19221,N_19124,N_19003);
nor U19222 (N_19222,N_18802,N_19013);
nor U19223 (N_19223,N_19097,N_19028);
nor U19224 (N_19224,N_19018,N_18824);
nor U19225 (N_19225,N_19087,N_19066);
and U19226 (N_19226,N_19085,N_18909);
or U19227 (N_19227,N_19022,N_18901);
xor U19228 (N_19228,N_19173,N_18925);
xnor U19229 (N_19229,N_18880,N_18884);
nor U19230 (N_19230,N_19128,N_18961);
nand U19231 (N_19231,N_18800,N_19106);
nand U19232 (N_19232,N_18922,N_18826);
nor U19233 (N_19233,N_19084,N_19154);
nor U19234 (N_19234,N_19100,N_18914);
and U19235 (N_19235,N_19050,N_19160);
and U19236 (N_19236,N_18811,N_18833);
nand U19237 (N_19237,N_19019,N_19112);
and U19238 (N_19238,N_19143,N_18908);
and U19239 (N_19239,N_19041,N_19105);
nand U19240 (N_19240,N_18907,N_19082);
or U19241 (N_19241,N_18899,N_18840);
nand U19242 (N_19242,N_19167,N_18995);
nor U19243 (N_19243,N_18836,N_19129);
or U19244 (N_19244,N_18970,N_18968);
and U19245 (N_19245,N_18841,N_19153);
or U19246 (N_19246,N_19139,N_19063);
nand U19247 (N_19247,N_18819,N_18866);
nor U19248 (N_19248,N_18935,N_18905);
nand U19249 (N_19249,N_19006,N_18818);
nor U19250 (N_19250,N_19055,N_19161);
nand U19251 (N_19251,N_19107,N_19194);
nand U19252 (N_19252,N_18878,N_19046);
nor U19253 (N_19253,N_19089,N_18949);
nand U19254 (N_19254,N_18816,N_19034);
nor U19255 (N_19255,N_19104,N_19101);
nor U19256 (N_19256,N_19032,N_19140);
or U19257 (N_19257,N_18997,N_18834);
and U19258 (N_19258,N_19008,N_19155);
and U19259 (N_19259,N_18988,N_18959);
or U19260 (N_19260,N_19189,N_18888);
nand U19261 (N_19261,N_19135,N_19075);
or U19262 (N_19262,N_18953,N_18892);
nor U19263 (N_19263,N_18952,N_18853);
nand U19264 (N_19264,N_19118,N_19133);
nand U19265 (N_19265,N_18837,N_18946);
and U19266 (N_19266,N_18923,N_18965);
and U19267 (N_19267,N_19145,N_18887);
nand U19268 (N_19268,N_18810,N_19051);
xor U19269 (N_19269,N_18976,N_19011);
and U19270 (N_19270,N_19020,N_19081);
nand U19271 (N_19271,N_18857,N_19168);
nor U19272 (N_19272,N_18924,N_18872);
and U19273 (N_19273,N_18933,N_19036);
and U19274 (N_19274,N_19103,N_19064);
or U19275 (N_19275,N_19062,N_19117);
or U19276 (N_19276,N_19110,N_18806);
nor U19277 (N_19277,N_19150,N_18913);
nand U19278 (N_19278,N_18904,N_19125);
and U19279 (N_19279,N_18876,N_19195);
and U19280 (N_19280,N_19114,N_19183);
or U19281 (N_19281,N_18948,N_18813);
and U19282 (N_19282,N_18996,N_18891);
and U19283 (N_19283,N_18864,N_18874);
or U19284 (N_19284,N_18859,N_19079);
or U19285 (N_19285,N_19121,N_18812);
and U19286 (N_19286,N_18954,N_19061);
and U19287 (N_19287,N_18999,N_18932);
nand U19288 (N_19288,N_18977,N_19067);
nand U19289 (N_19289,N_18860,N_19198);
nand U19290 (N_19290,N_19180,N_19136);
or U19291 (N_19291,N_19132,N_19060);
and U19292 (N_19292,N_18987,N_18980);
nand U19293 (N_19293,N_19152,N_18903);
or U19294 (N_19294,N_19175,N_18825);
and U19295 (N_19295,N_19141,N_18981);
nor U19296 (N_19296,N_19111,N_19159);
and U19297 (N_19297,N_18936,N_19007);
and U19298 (N_19298,N_18957,N_18877);
nand U19299 (N_19299,N_18985,N_19127);
and U19300 (N_19300,N_18894,N_18958);
and U19301 (N_19301,N_19123,N_19040);
or U19302 (N_19302,N_18854,N_18911);
and U19303 (N_19303,N_19109,N_19069);
nor U19304 (N_19304,N_19002,N_19039);
nor U19305 (N_19305,N_19172,N_19197);
and U19306 (N_19306,N_19014,N_18962);
or U19307 (N_19307,N_18882,N_19095);
or U19308 (N_19308,N_18982,N_18960);
nor U19309 (N_19309,N_18898,N_19166);
nand U19310 (N_19310,N_18852,N_19056);
nand U19311 (N_19311,N_18963,N_19030);
nand U19312 (N_19312,N_18895,N_19009);
and U19313 (N_19313,N_18972,N_18865);
nand U19314 (N_19314,N_19042,N_18817);
or U19315 (N_19315,N_18990,N_19090);
nand U19316 (N_19316,N_19017,N_18839);
and U19317 (N_19317,N_18993,N_18873);
nor U19318 (N_19318,N_19043,N_18931);
or U19319 (N_19319,N_18978,N_18934);
nor U19320 (N_19320,N_18998,N_19188);
or U19321 (N_19321,N_19120,N_19102);
nor U19322 (N_19322,N_19144,N_19016);
and U19323 (N_19323,N_18938,N_19187);
nand U19324 (N_19324,N_19047,N_18831);
nor U19325 (N_19325,N_18919,N_19181);
and U19326 (N_19326,N_19059,N_19169);
nand U19327 (N_19327,N_18805,N_19191);
or U19328 (N_19328,N_19156,N_19057);
and U19329 (N_19329,N_18991,N_18885);
or U19330 (N_19330,N_18845,N_18912);
nor U19331 (N_19331,N_19170,N_18832);
and U19332 (N_19332,N_18902,N_19048);
nand U19333 (N_19333,N_19171,N_19163);
and U19334 (N_19334,N_19053,N_18939);
and U19335 (N_19335,N_19147,N_18994);
nand U19336 (N_19336,N_19024,N_19126);
and U19337 (N_19337,N_18944,N_18966);
and U19338 (N_19338,N_19026,N_19074);
nand U19339 (N_19339,N_19031,N_19080);
or U19340 (N_19340,N_19096,N_18809);
nand U19341 (N_19341,N_18979,N_19092);
or U19342 (N_19342,N_19138,N_19091);
and U19343 (N_19343,N_18974,N_18986);
nor U19344 (N_19344,N_18875,N_19158);
nand U19345 (N_19345,N_18971,N_18955);
nand U19346 (N_19346,N_19182,N_19179);
nand U19347 (N_19347,N_19088,N_18879);
nor U19348 (N_19348,N_18921,N_18893);
or U19349 (N_19349,N_18868,N_19071);
nor U19350 (N_19350,N_18835,N_18945);
nand U19351 (N_19351,N_18984,N_19142);
or U19352 (N_19352,N_19116,N_19192);
nor U19353 (N_19353,N_18942,N_19086);
or U19354 (N_19354,N_19070,N_18927);
nor U19355 (N_19355,N_18801,N_18842);
xnor U19356 (N_19356,N_19049,N_19068);
nor U19357 (N_19357,N_19052,N_18964);
and U19358 (N_19358,N_18983,N_19157);
nand U19359 (N_19359,N_19099,N_19115);
and U19360 (N_19360,N_18951,N_19190);
nor U19361 (N_19361,N_19149,N_18804);
nand U19362 (N_19362,N_18975,N_18848);
nor U19363 (N_19363,N_19199,N_18973);
or U19364 (N_19364,N_18830,N_19010);
nand U19365 (N_19365,N_19038,N_18910);
and U19366 (N_19366,N_18956,N_19083);
nor U19367 (N_19367,N_18920,N_19045);
xor U19368 (N_19368,N_18900,N_18883);
and U19369 (N_19369,N_18869,N_18850);
nand U19370 (N_19370,N_18896,N_18926);
nand U19371 (N_19371,N_18928,N_19137);
nor U19372 (N_19372,N_18815,N_19001);
nand U19373 (N_19373,N_19058,N_19193);
nor U19374 (N_19374,N_19044,N_19174);
or U19375 (N_19375,N_18863,N_18967);
nand U19376 (N_19376,N_18906,N_18855);
nand U19377 (N_19377,N_19184,N_19065);
and U19378 (N_19378,N_18915,N_19185);
nor U19379 (N_19379,N_19151,N_18930);
or U19380 (N_19380,N_19027,N_18871);
nand U19381 (N_19381,N_19077,N_18890);
or U19382 (N_19382,N_18814,N_18820);
nor U19383 (N_19383,N_19148,N_19146);
and U19384 (N_19384,N_19015,N_19119);
and U19385 (N_19385,N_19196,N_19054);
xnor U19386 (N_19386,N_19033,N_19130);
nor U19387 (N_19387,N_18940,N_19178);
or U19388 (N_19388,N_18827,N_19078);
nor U19389 (N_19389,N_18828,N_18989);
nor U19390 (N_19390,N_18803,N_18867);
nor U19391 (N_19391,N_19012,N_18856);
and U19392 (N_19392,N_18843,N_18829);
or U19393 (N_19393,N_19098,N_18992);
nor U19394 (N_19394,N_18849,N_19162);
nand U19395 (N_19395,N_19108,N_19004);
or U19396 (N_19396,N_19134,N_19021);
and U19397 (N_19397,N_18861,N_18847);
and U19398 (N_19398,N_19023,N_19005);
nor U19399 (N_19399,N_18943,N_19176);
or U19400 (N_19400,N_19069,N_18964);
nor U19401 (N_19401,N_18928,N_19060);
or U19402 (N_19402,N_19054,N_19044);
nand U19403 (N_19403,N_18869,N_19000);
and U19404 (N_19404,N_19171,N_18944);
nor U19405 (N_19405,N_18993,N_18963);
or U19406 (N_19406,N_18844,N_18913);
and U19407 (N_19407,N_19056,N_18969);
nand U19408 (N_19408,N_18902,N_19167);
nor U19409 (N_19409,N_18842,N_19020);
and U19410 (N_19410,N_18829,N_19193);
nand U19411 (N_19411,N_19154,N_19191);
or U19412 (N_19412,N_19161,N_19057);
nand U19413 (N_19413,N_19103,N_19138);
or U19414 (N_19414,N_19027,N_18936);
or U19415 (N_19415,N_18960,N_18939);
nand U19416 (N_19416,N_18969,N_19114);
nor U19417 (N_19417,N_18824,N_19099);
and U19418 (N_19418,N_19157,N_18974);
nand U19419 (N_19419,N_18838,N_19036);
nor U19420 (N_19420,N_19039,N_18822);
nand U19421 (N_19421,N_18865,N_19080);
and U19422 (N_19422,N_19134,N_18935);
and U19423 (N_19423,N_19095,N_18913);
nand U19424 (N_19424,N_18995,N_19089);
or U19425 (N_19425,N_18961,N_19178);
nand U19426 (N_19426,N_18902,N_18905);
or U19427 (N_19427,N_19120,N_18870);
nor U19428 (N_19428,N_19140,N_19024);
nor U19429 (N_19429,N_19167,N_18905);
nor U19430 (N_19430,N_19082,N_19144);
or U19431 (N_19431,N_18850,N_18872);
and U19432 (N_19432,N_18861,N_19097);
nand U19433 (N_19433,N_18995,N_18848);
nand U19434 (N_19434,N_19110,N_18957);
nor U19435 (N_19435,N_19177,N_19184);
nand U19436 (N_19436,N_19043,N_18861);
nand U19437 (N_19437,N_19016,N_18905);
xnor U19438 (N_19438,N_18823,N_19126);
nor U19439 (N_19439,N_19088,N_18963);
or U19440 (N_19440,N_19147,N_19049);
nand U19441 (N_19441,N_19112,N_18858);
nand U19442 (N_19442,N_19169,N_19036);
or U19443 (N_19443,N_18863,N_18937);
nor U19444 (N_19444,N_19174,N_18868);
or U19445 (N_19445,N_19006,N_18865);
nor U19446 (N_19446,N_18904,N_18809);
or U19447 (N_19447,N_19125,N_18951);
and U19448 (N_19448,N_19110,N_18922);
or U19449 (N_19449,N_18853,N_19144);
and U19450 (N_19450,N_18840,N_18975);
or U19451 (N_19451,N_18900,N_19152);
nand U19452 (N_19452,N_18867,N_18930);
nor U19453 (N_19453,N_18823,N_18915);
nand U19454 (N_19454,N_19110,N_19079);
nor U19455 (N_19455,N_18901,N_19154);
nor U19456 (N_19456,N_19021,N_18890);
or U19457 (N_19457,N_18858,N_19166);
nand U19458 (N_19458,N_18837,N_18996);
nand U19459 (N_19459,N_19014,N_18810);
nor U19460 (N_19460,N_19114,N_18824);
or U19461 (N_19461,N_19036,N_18977);
nand U19462 (N_19462,N_18873,N_19019);
and U19463 (N_19463,N_19001,N_19022);
nand U19464 (N_19464,N_18955,N_19075);
and U19465 (N_19465,N_19029,N_18987);
or U19466 (N_19466,N_19008,N_18959);
nand U19467 (N_19467,N_18884,N_18904);
nand U19468 (N_19468,N_19093,N_19117);
nor U19469 (N_19469,N_18945,N_19007);
nand U19470 (N_19470,N_19062,N_18963);
nand U19471 (N_19471,N_18879,N_18906);
nand U19472 (N_19472,N_19051,N_18877);
nor U19473 (N_19473,N_18847,N_19154);
and U19474 (N_19474,N_19040,N_19100);
and U19475 (N_19475,N_19076,N_18889);
nor U19476 (N_19476,N_18854,N_19050);
or U19477 (N_19477,N_18937,N_18940);
nand U19478 (N_19478,N_19151,N_18986);
or U19479 (N_19479,N_19048,N_19168);
nand U19480 (N_19480,N_18949,N_18942);
nand U19481 (N_19481,N_19186,N_19019);
nor U19482 (N_19482,N_19185,N_18859);
or U19483 (N_19483,N_18866,N_18947);
xnor U19484 (N_19484,N_18948,N_19148);
and U19485 (N_19485,N_18981,N_19065);
nor U19486 (N_19486,N_19120,N_18803);
nand U19487 (N_19487,N_19195,N_18853);
nor U19488 (N_19488,N_19175,N_18862);
nor U19489 (N_19489,N_19183,N_18986);
nor U19490 (N_19490,N_18889,N_19172);
and U19491 (N_19491,N_18889,N_19054);
xor U19492 (N_19492,N_18814,N_18870);
nor U19493 (N_19493,N_18847,N_19114);
and U19494 (N_19494,N_19180,N_19097);
or U19495 (N_19495,N_18861,N_18982);
or U19496 (N_19496,N_18919,N_19031);
nor U19497 (N_19497,N_18956,N_18932);
or U19498 (N_19498,N_19041,N_18927);
nor U19499 (N_19499,N_18996,N_18961);
and U19500 (N_19500,N_18952,N_19073);
and U19501 (N_19501,N_19028,N_19171);
nand U19502 (N_19502,N_18938,N_18910);
nor U19503 (N_19503,N_18952,N_18912);
nor U19504 (N_19504,N_19145,N_18868);
or U19505 (N_19505,N_18964,N_18989);
nor U19506 (N_19506,N_19060,N_18987);
or U19507 (N_19507,N_18806,N_19060);
nor U19508 (N_19508,N_18980,N_18902);
nand U19509 (N_19509,N_19006,N_19196);
or U19510 (N_19510,N_18931,N_19056);
nor U19511 (N_19511,N_18916,N_18814);
nor U19512 (N_19512,N_18953,N_18980);
or U19513 (N_19513,N_18835,N_18839);
nor U19514 (N_19514,N_18976,N_18833);
nand U19515 (N_19515,N_18856,N_18939);
nor U19516 (N_19516,N_19176,N_18965);
nand U19517 (N_19517,N_18934,N_18926);
nor U19518 (N_19518,N_19116,N_19150);
or U19519 (N_19519,N_19065,N_19099);
nor U19520 (N_19520,N_19174,N_18943);
nand U19521 (N_19521,N_19064,N_18851);
or U19522 (N_19522,N_19172,N_19016);
nor U19523 (N_19523,N_18899,N_18824);
or U19524 (N_19524,N_18955,N_18976);
nand U19525 (N_19525,N_18864,N_19003);
nand U19526 (N_19526,N_18825,N_19036);
or U19527 (N_19527,N_19153,N_19121);
nor U19528 (N_19528,N_18962,N_19109);
nor U19529 (N_19529,N_18932,N_18955);
or U19530 (N_19530,N_18868,N_18938);
or U19531 (N_19531,N_19155,N_18966);
nor U19532 (N_19532,N_19183,N_19097);
nor U19533 (N_19533,N_19033,N_18983);
nor U19534 (N_19534,N_18957,N_19044);
and U19535 (N_19535,N_19070,N_19082);
and U19536 (N_19536,N_18894,N_18949);
nor U19537 (N_19537,N_19043,N_19173);
or U19538 (N_19538,N_19018,N_19073);
nor U19539 (N_19539,N_18956,N_19135);
nand U19540 (N_19540,N_18965,N_19193);
nand U19541 (N_19541,N_19027,N_18921);
nand U19542 (N_19542,N_18892,N_18912);
or U19543 (N_19543,N_18818,N_19105);
and U19544 (N_19544,N_19130,N_19049);
nand U19545 (N_19545,N_18964,N_18978);
and U19546 (N_19546,N_18902,N_19109);
and U19547 (N_19547,N_19045,N_18919);
and U19548 (N_19548,N_19096,N_19193);
and U19549 (N_19549,N_18892,N_18940);
or U19550 (N_19550,N_18893,N_18895);
nand U19551 (N_19551,N_19155,N_18875);
nand U19552 (N_19552,N_19131,N_19034);
or U19553 (N_19553,N_19071,N_18840);
nor U19554 (N_19554,N_19119,N_18973);
nand U19555 (N_19555,N_18837,N_18885);
nor U19556 (N_19556,N_19110,N_19147);
and U19557 (N_19557,N_18998,N_18975);
nand U19558 (N_19558,N_18853,N_18951);
nand U19559 (N_19559,N_19090,N_19176);
nand U19560 (N_19560,N_18913,N_18889);
and U19561 (N_19561,N_18875,N_19037);
nor U19562 (N_19562,N_19132,N_18865);
and U19563 (N_19563,N_18802,N_19066);
nor U19564 (N_19564,N_19057,N_19008);
nor U19565 (N_19565,N_18936,N_18927);
or U19566 (N_19566,N_18893,N_19175);
or U19567 (N_19567,N_18893,N_19014);
and U19568 (N_19568,N_19081,N_18914);
or U19569 (N_19569,N_18892,N_18811);
and U19570 (N_19570,N_19099,N_19126);
and U19571 (N_19571,N_19040,N_19172);
and U19572 (N_19572,N_19114,N_18997);
and U19573 (N_19573,N_19088,N_18902);
or U19574 (N_19574,N_19145,N_19101);
or U19575 (N_19575,N_18908,N_19037);
or U19576 (N_19576,N_18976,N_18901);
or U19577 (N_19577,N_19020,N_19025);
or U19578 (N_19578,N_19182,N_19060);
or U19579 (N_19579,N_18901,N_18855);
nand U19580 (N_19580,N_19018,N_19096);
nand U19581 (N_19581,N_18998,N_18961);
or U19582 (N_19582,N_18865,N_18827);
or U19583 (N_19583,N_18869,N_19019);
nand U19584 (N_19584,N_18842,N_19189);
nor U19585 (N_19585,N_19098,N_19007);
and U19586 (N_19586,N_19094,N_19172);
nor U19587 (N_19587,N_19054,N_19163);
or U19588 (N_19588,N_18893,N_18878);
and U19589 (N_19589,N_19066,N_19092);
nor U19590 (N_19590,N_19052,N_18857);
and U19591 (N_19591,N_18952,N_19118);
nor U19592 (N_19592,N_19189,N_18959);
and U19593 (N_19593,N_19048,N_19139);
nand U19594 (N_19594,N_19147,N_19051);
nand U19595 (N_19595,N_19100,N_19185);
nor U19596 (N_19596,N_19002,N_19183);
nor U19597 (N_19597,N_18949,N_19062);
and U19598 (N_19598,N_19166,N_19155);
nand U19599 (N_19599,N_19181,N_19056);
or U19600 (N_19600,N_19209,N_19366);
nor U19601 (N_19601,N_19267,N_19427);
nand U19602 (N_19602,N_19308,N_19493);
nor U19603 (N_19603,N_19322,N_19241);
and U19604 (N_19604,N_19595,N_19357);
nor U19605 (N_19605,N_19349,N_19499);
or U19606 (N_19606,N_19354,N_19553);
or U19607 (N_19607,N_19356,N_19491);
nand U19608 (N_19608,N_19251,N_19237);
and U19609 (N_19609,N_19232,N_19541);
nand U19610 (N_19610,N_19546,N_19299);
nor U19611 (N_19611,N_19304,N_19408);
or U19612 (N_19612,N_19524,N_19351);
nor U19613 (N_19613,N_19216,N_19453);
or U19614 (N_19614,N_19501,N_19570);
or U19615 (N_19615,N_19221,N_19328);
nor U19616 (N_19616,N_19573,N_19447);
nor U19617 (N_19617,N_19201,N_19314);
and U19618 (N_19618,N_19440,N_19548);
and U19619 (N_19619,N_19327,N_19426);
and U19620 (N_19620,N_19466,N_19297);
nor U19621 (N_19621,N_19487,N_19464);
or U19622 (N_19622,N_19584,N_19536);
and U19623 (N_19623,N_19436,N_19222);
or U19624 (N_19624,N_19326,N_19259);
and U19625 (N_19625,N_19270,N_19332);
or U19626 (N_19626,N_19391,N_19264);
nor U19627 (N_19627,N_19517,N_19262);
or U19628 (N_19628,N_19204,N_19579);
and U19629 (N_19629,N_19463,N_19286);
nor U19630 (N_19630,N_19520,N_19420);
nand U19631 (N_19631,N_19557,N_19476);
nor U19632 (N_19632,N_19335,N_19465);
nand U19633 (N_19633,N_19210,N_19376);
and U19634 (N_19634,N_19361,N_19223);
and U19635 (N_19635,N_19323,N_19559);
or U19636 (N_19636,N_19229,N_19431);
nor U19637 (N_19637,N_19249,N_19468);
or U19638 (N_19638,N_19537,N_19333);
or U19639 (N_19639,N_19258,N_19534);
nand U19640 (N_19640,N_19254,N_19490);
nor U19641 (N_19641,N_19371,N_19578);
nand U19642 (N_19642,N_19377,N_19280);
nand U19643 (N_19643,N_19485,N_19581);
nand U19644 (N_19644,N_19279,N_19471);
nor U19645 (N_19645,N_19217,N_19244);
nor U19646 (N_19646,N_19211,N_19511);
or U19647 (N_19647,N_19393,N_19392);
nand U19648 (N_19648,N_19302,N_19418);
or U19649 (N_19649,N_19292,N_19576);
or U19650 (N_19650,N_19489,N_19274);
nor U19651 (N_19651,N_19288,N_19394);
and U19652 (N_19652,N_19290,N_19320);
nor U19653 (N_19653,N_19372,N_19321);
nor U19654 (N_19654,N_19535,N_19564);
nor U19655 (N_19655,N_19345,N_19514);
nor U19656 (N_19656,N_19448,N_19383);
nor U19657 (N_19657,N_19592,N_19437);
nand U19658 (N_19658,N_19594,N_19213);
nor U19659 (N_19659,N_19227,N_19449);
or U19660 (N_19660,N_19398,N_19325);
nand U19661 (N_19661,N_19593,N_19563);
and U19662 (N_19662,N_19482,N_19363);
and U19663 (N_19663,N_19291,N_19329);
xnor U19664 (N_19664,N_19336,N_19547);
or U19665 (N_19665,N_19273,N_19247);
or U19666 (N_19666,N_19386,N_19462);
and U19667 (N_19667,N_19240,N_19331);
and U19668 (N_19668,N_19330,N_19246);
nand U19669 (N_19669,N_19544,N_19384);
and U19670 (N_19670,N_19538,N_19340);
xnor U19671 (N_19671,N_19375,N_19575);
nand U19672 (N_19672,N_19528,N_19307);
or U19673 (N_19673,N_19556,N_19589);
xnor U19674 (N_19674,N_19586,N_19219);
nor U19675 (N_19675,N_19269,N_19452);
nand U19676 (N_19676,N_19587,N_19532);
or U19677 (N_19677,N_19255,N_19470);
and U19678 (N_19678,N_19577,N_19225);
nor U19679 (N_19679,N_19206,N_19226);
nand U19680 (N_19680,N_19303,N_19294);
nor U19681 (N_19681,N_19425,N_19224);
and U19682 (N_19682,N_19261,N_19359);
nor U19683 (N_19683,N_19282,N_19272);
or U19684 (N_19684,N_19390,N_19271);
and U19685 (N_19685,N_19413,N_19539);
or U19686 (N_19686,N_19498,N_19389);
and U19687 (N_19687,N_19342,N_19549);
nor U19688 (N_19688,N_19341,N_19545);
and U19689 (N_19689,N_19234,N_19504);
nand U19690 (N_19690,N_19405,N_19521);
and U19691 (N_19691,N_19347,N_19287);
nor U19692 (N_19692,N_19355,N_19250);
or U19693 (N_19693,N_19235,N_19560);
and U19694 (N_19694,N_19457,N_19571);
nor U19695 (N_19695,N_19407,N_19414);
nor U19696 (N_19696,N_19515,N_19367);
or U19697 (N_19697,N_19481,N_19551);
or U19698 (N_19698,N_19508,N_19590);
nand U19699 (N_19699,N_19358,N_19301);
and U19700 (N_19700,N_19236,N_19439);
nand U19701 (N_19701,N_19572,N_19554);
and U19702 (N_19702,N_19523,N_19474);
and U19703 (N_19703,N_19374,N_19239);
xnor U19704 (N_19704,N_19380,N_19442);
nand U19705 (N_19705,N_19555,N_19315);
and U19706 (N_19706,N_19588,N_19284);
nand U19707 (N_19707,N_19566,N_19403);
nand U19708 (N_19708,N_19215,N_19519);
and U19709 (N_19709,N_19467,N_19568);
nor U19710 (N_19710,N_19387,N_19253);
nand U19711 (N_19711,N_19552,N_19458);
nor U19712 (N_19712,N_19339,N_19218);
nor U19713 (N_19713,N_19343,N_19574);
or U19714 (N_19714,N_19260,N_19472);
and U19715 (N_19715,N_19446,N_19283);
nand U19716 (N_19716,N_19451,N_19207);
and U19717 (N_19717,N_19510,N_19205);
nor U19718 (N_19718,N_19319,N_19382);
nand U19719 (N_19719,N_19434,N_19395);
and U19720 (N_19720,N_19245,N_19561);
nand U19721 (N_19721,N_19518,N_19399);
or U19722 (N_19722,N_19404,N_19542);
nor U19723 (N_19723,N_19500,N_19344);
nor U19724 (N_19724,N_19311,N_19317);
or U19725 (N_19725,N_19483,N_19379);
or U19726 (N_19726,N_19443,N_19432);
nor U19727 (N_19727,N_19582,N_19313);
and U19728 (N_19728,N_19373,N_19248);
nor U19729 (N_19729,N_19369,N_19334);
and U19730 (N_19730,N_19479,N_19461);
and U19731 (N_19731,N_19475,N_19370);
or U19732 (N_19732,N_19348,N_19296);
or U19733 (N_19733,N_19591,N_19435);
nor U19734 (N_19734,N_19455,N_19202);
nor U19735 (N_19735,N_19353,N_19421);
and U19736 (N_19736,N_19423,N_19480);
nor U19737 (N_19737,N_19486,N_19505);
nor U19738 (N_19738,N_19506,N_19502);
nand U19739 (N_19739,N_19306,N_19459);
nor U19740 (N_19740,N_19200,N_19309);
nand U19741 (N_19741,N_19295,N_19265);
or U19742 (N_19742,N_19208,N_19550);
nand U19743 (N_19743,N_19415,N_19424);
nor U19744 (N_19744,N_19428,N_19278);
nand U19745 (N_19745,N_19238,N_19396);
xor U19746 (N_19746,N_19212,N_19233);
nand U19747 (N_19747,N_19312,N_19350);
or U19748 (N_19748,N_19360,N_19569);
nand U19749 (N_19749,N_19530,N_19598);
nor U19750 (N_19750,N_19531,N_19507);
and U19751 (N_19751,N_19512,N_19364);
or U19752 (N_19752,N_19289,N_19324);
nand U19753 (N_19753,N_19441,N_19516);
nand U19754 (N_19754,N_19565,N_19597);
nor U19755 (N_19755,N_19585,N_19580);
nand U19756 (N_19756,N_19275,N_19495);
nor U19757 (N_19757,N_19526,N_19484);
or U19758 (N_19758,N_19263,N_19362);
nor U19759 (N_19759,N_19316,N_19293);
nor U19760 (N_19760,N_19228,N_19558);
nor U19761 (N_19761,N_19281,N_19397);
nor U19762 (N_19762,N_19477,N_19402);
nor U19763 (N_19763,N_19417,N_19444);
nor U19764 (N_19764,N_19496,N_19522);
or U19765 (N_19765,N_19266,N_19406);
or U19766 (N_19766,N_19368,N_19540);
nor U19767 (N_19767,N_19346,N_19252);
or U19768 (N_19768,N_19378,N_19460);
nand U19769 (N_19769,N_19438,N_19409);
and U19770 (N_19770,N_19419,N_19220);
and U19771 (N_19771,N_19445,N_19318);
nand U19772 (N_19772,N_19567,N_19529);
and U19773 (N_19773,N_19300,N_19429);
nor U19774 (N_19774,N_19385,N_19381);
or U19775 (N_19775,N_19422,N_19388);
or U19776 (N_19776,N_19285,N_19243);
and U19777 (N_19777,N_19203,N_19562);
and U19778 (N_19778,N_19513,N_19256);
nand U19779 (N_19779,N_19543,N_19410);
or U19780 (N_19780,N_19492,N_19411);
and U19781 (N_19781,N_19214,N_19583);
nand U19782 (N_19782,N_19412,N_19527);
nor U19783 (N_19783,N_19503,N_19365);
or U19784 (N_19784,N_19599,N_19298);
or U19785 (N_19785,N_19488,N_19257);
and U19786 (N_19786,N_19430,N_19242);
nand U19787 (N_19787,N_19596,N_19338);
or U19788 (N_19788,N_19450,N_19509);
and U19789 (N_19789,N_19433,N_19469);
and U19790 (N_19790,N_19277,N_19305);
nor U19791 (N_19791,N_19231,N_19276);
nand U19792 (N_19792,N_19416,N_19400);
nand U19793 (N_19793,N_19494,N_19401);
nand U19794 (N_19794,N_19497,N_19473);
or U19795 (N_19795,N_19310,N_19533);
nor U19796 (N_19796,N_19454,N_19352);
nor U19797 (N_19797,N_19337,N_19478);
nor U19798 (N_19798,N_19456,N_19268);
nor U19799 (N_19799,N_19525,N_19230);
nor U19800 (N_19800,N_19393,N_19308);
nor U19801 (N_19801,N_19357,N_19587);
or U19802 (N_19802,N_19325,N_19510);
and U19803 (N_19803,N_19542,N_19330);
nand U19804 (N_19804,N_19448,N_19431);
nor U19805 (N_19805,N_19590,N_19364);
or U19806 (N_19806,N_19563,N_19448);
and U19807 (N_19807,N_19388,N_19236);
nand U19808 (N_19808,N_19204,N_19525);
nand U19809 (N_19809,N_19500,N_19278);
and U19810 (N_19810,N_19373,N_19211);
nor U19811 (N_19811,N_19271,N_19430);
nand U19812 (N_19812,N_19486,N_19489);
nand U19813 (N_19813,N_19330,N_19250);
or U19814 (N_19814,N_19543,N_19552);
nand U19815 (N_19815,N_19379,N_19358);
or U19816 (N_19816,N_19261,N_19494);
and U19817 (N_19817,N_19201,N_19214);
or U19818 (N_19818,N_19370,N_19376);
nand U19819 (N_19819,N_19419,N_19267);
or U19820 (N_19820,N_19220,N_19575);
nand U19821 (N_19821,N_19281,N_19301);
nand U19822 (N_19822,N_19538,N_19415);
and U19823 (N_19823,N_19463,N_19544);
nand U19824 (N_19824,N_19454,N_19324);
nor U19825 (N_19825,N_19290,N_19548);
or U19826 (N_19826,N_19249,N_19411);
and U19827 (N_19827,N_19557,N_19590);
or U19828 (N_19828,N_19422,N_19551);
and U19829 (N_19829,N_19330,N_19257);
or U19830 (N_19830,N_19293,N_19251);
nor U19831 (N_19831,N_19249,N_19421);
and U19832 (N_19832,N_19510,N_19458);
and U19833 (N_19833,N_19277,N_19588);
nor U19834 (N_19834,N_19408,N_19434);
nor U19835 (N_19835,N_19445,N_19372);
nor U19836 (N_19836,N_19225,N_19319);
or U19837 (N_19837,N_19564,N_19416);
nor U19838 (N_19838,N_19470,N_19293);
nand U19839 (N_19839,N_19546,N_19579);
nor U19840 (N_19840,N_19409,N_19419);
and U19841 (N_19841,N_19249,N_19536);
and U19842 (N_19842,N_19416,N_19548);
nand U19843 (N_19843,N_19513,N_19452);
or U19844 (N_19844,N_19558,N_19436);
or U19845 (N_19845,N_19250,N_19474);
or U19846 (N_19846,N_19216,N_19480);
nand U19847 (N_19847,N_19425,N_19512);
and U19848 (N_19848,N_19478,N_19506);
and U19849 (N_19849,N_19426,N_19219);
and U19850 (N_19850,N_19447,N_19222);
nor U19851 (N_19851,N_19309,N_19418);
and U19852 (N_19852,N_19230,N_19274);
and U19853 (N_19853,N_19255,N_19308);
nor U19854 (N_19854,N_19480,N_19425);
and U19855 (N_19855,N_19390,N_19250);
nand U19856 (N_19856,N_19292,N_19462);
or U19857 (N_19857,N_19519,N_19301);
nand U19858 (N_19858,N_19362,N_19508);
or U19859 (N_19859,N_19435,N_19529);
nor U19860 (N_19860,N_19324,N_19235);
or U19861 (N_19861,N_19481,N_19253);
nor U19862 (N_19862,N_19257,N_19379);
nor U19863 (N_19863,N_19444,N_19569);
or U19864 (N_19864,N_19215,N_19418);
and U19865 (N_19865,N_19351,N_19264);
and U19866 (N_19866,N_19542,N_19372);
nand U19867 (N_19867,N_19329,N_19218);
nand U19868 (N_19868,N_19342,N_19250);
nor U19869 (N_19869,N_19479,N_19433);
nand U19870 (N_19870,N_19586,N_19334);
or U19871 (N_19871,N_19201,N_19356);
nor U19872 (N_19872,N_19231,N_19306);
and U19873 (N_19873,N_19321,N_19351);
or U19874 (N_19874,N_19210,N_19399);
and U19875 (N_19875,N_19504,N_19577);
nand U19876 (N_19876,N_19335,N_19469);
and U19877 (N_19877,N_19260,N_19532);
and U19878 (N_19878,N_19271,N_19235);
nor U19879 (N_19879,N_19504,N_19386);
or U19880 (N_19880,N_19553,N_19530);
nor U19881 (N_19881,N_19443,N_19215);
or U19882 (N_19882,N_19330,N_19559);
or U19883 (N_19883,N_19386,N_19231);
and U19884 (N_19884,N_19350,N_19517);
and U19885 (N_19885,N_19508,N_19455);
and U19886 (N_19886,N_19243,N_19273);
and U19887 (N_19887,N_19553,N_19335);
and U19888 (N_19888,N_19314,N_19587);
and U19889 (N_19889,N_19200,N_19460);
nor U19890 (N_19890,N_19479,N_19397);
nor U19891 (N_19891,N_19386,N_19258);
and U19892 (N_19892,N_19547,N_19394);
and U19893 (N_19893,N_19510,N_19250);
nor U19894 (N_19894,N_19448,N_19577);
or U19895 (N_19895,N_19262,N_19424);
and U19896 (N_19896,N_19389,N_19274);
nand U19897 (N_19897,N_19486,N_19229);
or U19898 (N_19898,N_19363,N_19247);
nor U19899 (N_19899,N_19360,N_19365);
nand U19900 (N_19900,N_19478,N_19319);
nand U19901 (N_19901,N_19412,N_19599);
nor U19902 (N_19902,N_19493,N_19436);
or U19903 (N_19903,N_19263,N_19568);
nor U19904 (N_19904,N_19271,N_19508);
nor U19905 (N_19905,N_19480,N_19545);
nand U19906 (N_19906,N_19286,N_19452);
or U19907 (N_19907,N_19320,N_19596);
nand U19908 (N_19908,N_19257,N_19520);
nand U19909 (N_19909,N_19244,N_19400);
nor U19910 (N_19910,N_19372,N_19285);
nor U19911 (N_19911,N_19357,N_19247);
nand U19912 (N_19912,N_19494,N_19373);
and U19913 (N_19913,N_19373,N_19512);
nor U19914 (N_19914,N_19494,N_19295);
and U19915 (N_19915,N_19262,N_19240);
and U19916 (N_19916,N_19517,N_19210);
nand U19917 (N_19917,N_19444,N_19591);
or U19918 (N_19918,N_19591,N_19527);
nand U19919 (N_19919,N_19290,N_19442);
nand U19920 (N_19920,N_19205,N_19280);
or U19921 (N_19921,N_19401,N_19567);
or U19922 (N_19922,N_19549,N_19214);
and U19923 (N_19923,N_19481,N_19439);
nor U19924 (N_19924,N_19471,N_19315);
nand U19925 (N_19925,N_19549,N_19531);
and U19926 (N_19926,N_19473,N_19375);
nor U19927 (N_19927,N_19219,N_19338);
nand U19928 (N_19928,N_19399,N_19297);
and U19929 (N_19929,N_19337,N_19299);
and U19930 (N_19930,N_19289,N_19591);
or U19931 (N_19931,N_19480,N_19562);
nor U19932 (N_19932,N_19260,N_19488);
or U19933 (N_19933,N_19370,N_19280);
or U19934 (N_19934,N_19314,N_19440);
and U19935 (N_19935,N_19503,N_19578);
nor U19936 (N_19936,N_19500,N_19464);
or U19937 (N_19937,N_19202,N_19304);
or U19938 (N_19938,N_19245,N_19469);
nor U19939 (N_19939,N_19520,N_19518);
nand U19940 (N_19940,N_19372,N_19202);
nor U19941 (N_19941,N_19271,N_19416);
and U19942 (N_19942,N_19298,N_19472);
or U19943 (N_19943,N_19385,N_19548);
or U19944 (N_19944,N_19590,N_19581);
nor U19945 (N_19945,N_19202,N_19413);
and U19946 (N_19946,N_19289,N_19387);
and U19947 (N_19947,N_19563,N_19238);
or U19948 (N_19948,N_19588,N_19414);
nor U19949 (N_19949,N_19562,N_19355);
or U19950 (N_19950,N_19557,N_19446);
nor U19951 (N_19951,N_19571,N_19248);
nand U19952 (N_19952,N_19494,N_19366);
and U19953 (N_19953,N_19584,N_19238);
and U19954 (N_19954,N_19451,N_19546);
nand U19955 (N_19955,N_19233,N_19344);
nor U19956 (N_19956,N_19328,N_19338);
nand U19957 (N_19957,N_19214,N_19364);
and U19958 (N_19958,N_19331,N_19569);
and U19959 (N_19959,N_19461,N_19431);
nand U19960 (N_19960,N_19436,N_19580);
nor U19961 (N_19961,N_19350,N_19265);
and U19962 (N_19962,N_19235,N_19285);
nand U19963 (N_19963,N_19424,N_19444);
or U19964 (N_19964,N_19395,N_19574);
and U19965 (N_19965,N_19532,N_19229);
nand U19966 (N_19966,N_19337,N_19530);
nor U19967 (N_19967,N_19499,N_19255);
or U19968 (N_19968,N_19486,N_19230);
nor U19969 (N_19969,N_19280,N_19458);
nor U19970 (N_19970,N_19305,N_19477);
nand U19971 (N_19971,N_19232,N_19264);
or U19972 (N_19972,N_19371,N_19238);
nor U19973 (N_19973,N_19258,N_19565);
and U19974 (N_19974,N_19411,N_19420);
nor U19975 (N_19975,N_19574,N_19315);
nor U19976 (N_19976,N_19303,N_19362);
and U19977 (N_19977,N_19458,N_19431);
and U19978 (N_19978,N_19526,N_19494);
and U19979 (N_19979,N_19536,N_19241);
or U19980 (N_19980,N_19379,N_19517);
nor U19981 (N_19981,N_19476,N_19321);
or U19982 (N_19982,N_19251,N_19289);
or U19983 (N_19983,N_19246,N_19207);
nand U19984 (N_19984,N_19218,N_19543);
nand U19985 (N_19985,N_19531,N_19236);
nor U19986 (N_19986,N_19531,N_19408);
nor U19987 (N_19987,N_19270,N_19340);
nor U19988 (N_19988,N_19275,N_19432);
and U19989 (N_19989,N_19338,N_19562);
or U19990 (N_19990,N_19409,N_19441);
and U19991 (N_19991,N_19321,N_19568);
nor U19992 (N_19992,N_19475,N_19391);
nor U19993 (N_19993,N_19560,N_19543);
nand U19994 (N_19994,N_19559,N_19290);
nor U19995 (N_19995,N_19537,N_19270);
or U19996 (N_19996,N_19513,N_19510);
nor U19997 (N_19997,N_19420,N_19200);
and U19998 (N_19998,N_19228,N_19512);
nor U19999 (N_19999,N_19293,N_19447);
and UO_0 (O_0,N_19612,N_19706);
nor UO_1 (O_1,N_19946,N_19750);
nand UO_2 (O_2,N_19951,N_19967);
nand UO_3 (O_3,N_19836,N_19714);
or UO_4 (O_4,N_19776,N_19662);
and UO_5 (O_5,N_19827,N_19793);
nand UO_6 (O_6,N_19938,N_19957);
nand UO_7 (O_7,N_19870,N_19780);
nand UO_8 (O_8,N_19752,N_19751);
and UO_9 (O_9,N_19701,N_19925);
and UO_10 (O_10,N_19647,N_19990);
and UO_11 (O_11,N_19964,N_19656);
nor UO_12 (O_12,N_19815,N_19670);
nand UO_13 (O_13,N_19866,N_19959);
and UO_14 (O_14,N_19893,N_19829);
nor UO_15 (O_15,N_19619,N_19687);
nand UO_16 (O_16,N_19824,N_19673);
xor UO_17 (O_17,N_19853,N_19801);
and UO_18 (O_18,N_19861,N_19920);
and UO_19 (O_19,N_19688,N_19728);
nor UO_20 (O_20,N_19930,N_19678);
or UO_21 (O_21,N_19718,N_19999);
or UO_22 (O_22,N_19826,N_19790);
and UO_23 (O_23,N_19624,N_19653);
and UO_24 (O_24,N_19939,N_19926);
nand UO_25 (O_25,N_19969,N_19680);
and UO_26 (O_26,N_19772,N_19982);
and UO_27 (O_27,N_19807,N_19702);
and UO_28 (O_28,N_19968,N_19880);
and UO_29 (O_29,N_19984,N_19667);
and UO_30 (O_30,N_19844,N_19769);
or UO_31 (O_31,N_19983,N_19710);
nor UO_32 (O_32,N_19980,N_19846);
nor UO_33 (O_33,N_19734,N_19633);
or UO_34 (O_34,N_19813,N_19794);
nand UO_35 (O_35,N_19778,N_19655);
nor UO_36 (O_36,N_19877,N_19909);
nand UO_37 (O_37,N_19860,N_19935);
and UO_38 (O_38,N_19966,N_19689);
or UO_39 (O_39,N_19685,N_19927);
and UO_40 (O_40,N_19858,N_19819);
nand UO_41 (O_41,N_19806,N_19742);
or UO_42 (O_42,N_19623,N_19631);
or UO_43 (O_43,N_19975,N_19894);
nand UO_44 (O_44,N_19683,N_19977);
or UO_45 (O_45,N_19901,N_19757);
nor UO_46 (O_46,N_19717,N_19989);
nand UO_47 (O_47,N_19630,N_19625);
and UO_48 (O_48,N_19998,N_19665);
nand UO_49 (O_49,N_19690,N_19922);
nand UO_50 (O_50,N_19889,N_19876);
nand UO_51 (O_51,N_19740,N_19981);
nor UO_52 (O_52,N_19875,N_19614);
or UO_53 (O_53,N_19764,N_19708);
or UO_54 (O_54,N_19945,N_19747);
nand UO_55 (O_55,N_19638,N_19944);
and UO_56 (O_56,N_19885,N_19672);
nand UO_57 (O_57,N_19960,N_19881);
nor UO_58 (O_58,N_19765,N_19973);
or UO_59 (O_59,N_19737,N_19715);
or UO_60 (O_60,N_19629,N_19917);
nand UO_61 (O_61,N_19779,N_19912);
or UO_62 (O_62,N_19635,N_19963);
nand UO_63 (O_63,N_19664,N_19962);
and UO_64 (O_64,N_19906,N_19642);
xor UO_65 (O_65,N_19895,N_19732);
or UO_66 (O_66,N_19652,N_19684);
or UO_67 (O_67,N_19785,N_19992);
or UO_68 (O_68,N_19755,N_19654);
nand UO_69 (O_69,N_19756,N_19608);
nand UO_70 (O_70,N_19798,N_19822);
or UO_71 (O_71,N_19784,N_19682);
nand UO_72 (O_72,N_19848,N_19847);
or UO_73 (O_73,N_19816,N_19695);
nor UO_74 (O_74,N_19676,N_19852);
nand UO_75 (O_75,N_19952,N_19716);
and UO_76 (O_76,N_19868,N_19943);
nand UO_77 (O_77,N_19767,N_19928);
and UO_78 (O_78,N_19735,N_19805);
and UO_79 (O_79,N_19646,N_19660);
and UO_80 (O_80,N_19803,N_19703);
and UO_81 (O_81,N_19726,N_19995);
or UO_82 (O_82,N_19965,N_19797);
nand UO_83 (O_83,N_19787,N_19753);
nand UO_84 (O_84,N_19843,N_19993);
and UO_85 (O_85,N_19712,N_19804);
and UO_86 (O_86,N_19615,N_19659);
and UO_87 (O_87,N_19634,N_19788);
nand UO_88 (O_88,N_19955,N_19621);
and UO_89 (O_89,N_19949,N_19723);
nor UO_90 (O_90,N_19934,N_19869);
or UO_91 (O_91,N_19919,N_19611);
xor UO_92 (O_92,N_19762,N_19763);
nor UO_93 (O_93,N_19768,N_19746);
and UO_94 (O_94,N_19617,N_19907);
nand UO_95 (O_95,N_19613,N_19872);
or UO_96 (O_96,N_19627,N_19773);
and UO_97 (O_97,N_19626,N_19771);
nor UO_98 (O_98,N_19650,N_19668);
or UO_99 (O_99,N_19792,N_19908);
nand UO_100 (O_100,N_19834,N_19727);
or UO_101 (O_101,N_19645,N_19748);
or UO_102 (O_102,N_19758,N_19905);
or UO_103 (O_103,N_19759,N_19622);
and UO_104 (O_104,N_19979,N_19825);
or UO_105 (O_105,N_19675,N_19602);
nand UO_106 (O_106,N_19741,N_19958);
or UO_107 (O_107,N_19810,N_19867);
nand UO_108 (O_108,N_19855,N_19641);
or UO_109 (O_109,N_19692,N_19986);
or UO_110 (O_110,N_19904,N_19738);
nor UO_111 (O_111,N_19796,N_19677);
and UO_112 (O_112,N_19828,N_19637);
or UO_113 (O_113,N_19809,N_19818);
and UO_114 (O_114,N_19820,N_19886);
nand UO_115 (O_115,N_19823,N_19971);
or UO_116 (O_116,N_19812,N_19976);
nor UO_117 (O_117,N_19942,N_19863);
nor UO_118 (O_118,N_19865,N_19658);
or UO_119 (O_119,N_19814,N_19657);
or UO_120 (O_120,N_19666,N_19648);
or UO_121 (O_121,N_19839,N_19761);
nand UO_122 (O_122,N_19704,N_19760);
nor UO_123 (O_123,N_19775,N_19719);
nor UO_124 (O_124,N_19879,N_19897);
or UO_125 (O_125,N_19850,N_19639);
nor UO_126 (O_126,N_19896,N_19974);
and UO_127 (O_127,N_19817,N_19857);
nand UO_128 (O_128,N_19749,N_19936);
and UO_129 (O_129,N_19941,N_19700);
nand UO_130 (O_130,N_19720,N_19661);
nor UO_131 (O_131,N_19808,N_19671);
and UO_132 (O_132,N_19953,N_19996);
nor UO_133 (O_133,N_19831,N_19838);
or UO_134 (O_134,N_19699,N_19777);
or UO_135 (O_135,N_19725,N_19864);
nand UO_136 (O_136,N_19910,N_19988);
and UO_137 (O_137,N_19892,N_19915);
nand UO_138 (O_138,N_19709,N_19947);
and UO_139 (O_139,N_19698,N_19991);
and UO_140 (O_140,N_19950,N_19610);
nor UO_141 (O_141,N_19888,N_19837);
and UO_142 (O_142,N_19651,N_19849);
or UO_143 (O_143,N_19636,N_19916);
nor UO_144 (O_144,N_19911,N_19891);
nand UO_145 (O_145,N_19724,N_19851);
nand UO_146 (O_146,N_19733,N_19628);
nand UO_147 (O_147,N_19603,N_19620);
or UO_148 (O_148,N_19994,N_19795);
and UO_149 (O_149,N_19640,N_19663);
and UO_150 (O_150,N_19900,N_19845);
and UO_151 (O_151,N_19743,N_19832);
or UO_152 (O_152,N_19821,N_19800);
or UO_153 (O_153,N_19609,N_19887);
or UO_154 (O_154,N_19841,N_19697);
and UO_155 (O_155,N_19978,N_19883);
nand UO_156 (O_156,N_19691,N_19929);
nor UO_157 (O_157,N_19948,N_19791);
nor UO_158 (O_158,N_19729,N_19713);
nand UO_159 (O_159,N_19890,N_19882);
nor UO_160 (O_160,N_19931,N_19711);
nor UO_161 (O_161,N_19679,N_19707);
nand UO_162 (O_162,N_19766,N_19921);
nor UO_163 (O_163,N_19937,N_19669);
and UO_164 (O_164,N_19924,N_19693);
or UO_165 (O_165,N_19722,N_19754);
or UO_166 (O_166,N_19874,N_19811);
nor UO_167 (O_167,N_19783,N_19644);
or UO_168 (O_168,N_19898,N_19607);
nor UO_169 (O_169,N_19961,N_19903);
nand UO_170 (O_170,N_19744,N_19681);
and UO_171 (O_171,N_19840,N_19730);
nor UO_172 (O_172,N_19601,N_19954);
or UO_173 (O_173,N_19830,N_19873);
nor UO_174 (O_174,N_19854,N_19856);
nand UO_175 (O_175,N_19745,N_19782);
and UO_176 (O_176,N_19739,N_19731);
and UO_177 (O_177,N_19605,N_19970);
nand UO_178 (O_178,N_19972,N_19932);
nand UO_179 (O_179,N_19923,N_19770);
nor UO_180 (O_180,N_19899,N_19616);
or UO_181 (O_181,N_19781,N_19600);
or UO_182 (O_182,N_19884,N_19902);
or UO_183 (O_183,N_19774,N_19786);
nor UO_184 (O_184,N_19649,N_19987);
nor UO_185 (O_185,N_19632,N_19859);
nor UO_186 (O_186,N_19940,N_19913);
and UO_187 (O_187,N_19878,N_19835);
nor UO_188 (O_188,N_19674,N_19705);
nor UO_189 (O_189,N_19871,N_19606);
nand UO_190 (O_190,N_19799,N_19918);
nor UO_191 (O_191,N_19604,N_19802);
nor UO_192 (O_192,N_19789,N_19736);
nand UO_193 (O_193,N_19842,N_19862);
nor UO_194 (O_194,N_19686,N_19914);
nor UO_195 (O_195,N_19933,N_19618);
nor UO_196 (O_196,N_19694,N_19985);
nor UO_197 (O_197,N_19696,N_19643);
xnor UO_198 (O_198,N_19956,N_19833);
nor UO_199 (O_199,N_19721,N_19997);
nand UO_200 (O_200,N_19935,N_19757);
and UO_201 (O_201,N_19995,N_19647);
nor UO_202 (O_202,N_19680,N_19835);
or UO_203 (O_203,N_19969,N_19743);
or UO_204 (O_204,N_19969,N_19705);
nand UO_205 (O_205,N_19879,N_19764);
or UO_206 (O_206,N_19943,N_19789);
nor UO_207 (O_207,N_19779,N_19959);
nor UO_208 (O_208,N_19876,N_19921);
nand UO_209 (O_209,N_19849,N_19986);
or UO_210 (O_210,N_19762,N_19656);
and UO_211 (O_211,N_19612,N_19841);
nand UO_212 (O_212,N_19933,N_19795);
or UO_213 (O_213,N_19721,N_19632);
and UO_214 (O_214,N_19779,N_19915);
or UO_215 (O_215,N_19663,N_19890);
nand UO_216 (O_216,N_19830,N_19660);
xnor UO_217 (O_217,N_19817,N_19907);
nor UO_218 (O_218,N_19942,N_19806);
nand UO_219 (O_219,N_19853,N_19866);
nor UO_220 (O_220,N_19736,N_19611);
and UO_221 (O_221,N_19957,N_19863);
and UO_222 (O_222,N_19788,N_19903);
or UO_223 (O_223,N_19830,N_19683);
or UO_224 (O_224,N_19700,N_19854);
and UO_225 (O_225,N_19618,N_19606);
nor UO_226 (O_226,N_19681,N_19888);
xnor UO_227 (O_227,N_19641,N_19906);
nor UO_228 (O_228,N_19767,N_19941);
nor UO_229 (O_229,N_19796,N_19951);
and UO_230 (O_230,N_19863,N_19695);
nand UO_231 (O_231,N_19792,N_19922);
and UO_232 (O_232,N_19701,N_19853);
and UO_233 (O_233,N_19766,N_19756);
nor UO_234 (O_234,N_19798,N_19780);
xor UO_235 (O_235,N_19966,N_19735);
nor UO_236 (O_236,N_19833,N_19807);
nand UO_237 (O_237,N_19612,N_19806);
nor UO_238 (O_238,N_19745,N_19885);
and UO_239 (O_239,N_19792,N_19752);
nand UO_240 (O_240,N_19632,N_19806);
or UO_241 (O_241,N_19781,N_19995);
nand UO_242 (O_242,N_19821,N_19855);
and UO_243 (O_243,N_19618,N_19689);
nand UO_244 (O_244,N_19602,N_19906);
or UO_245 (O_245,N_19637,N_19825);
nand UO_246 (O_246,N_19771,N_19844);
nand UO_247 (O_247,N_19610,N_19904);
and UO_248 (O_248,N_19749,N_19908);
or UO_249 (O_249,N_19745,N_19842);
or UO_250 (O_250,N_19649,N_19754);
nor UO_251 (O_251,N_19610,N_19827);
nor UO_252 (O_252,N_19759,N_19697);
nor UO_253 (O_253,N_19938,N_19908);
and UO_254 (O_254,N_19819,N_19878);
and UO_255 (O_255,N_19707,N_19911);
or UO_256 (O_256,N_19629,N_19950);
nor UO_257 (O_257,N_19711,N_19696);
nor UO_258 (O_258,N_19860,N_19946);
nor UO_259 (O_259,N_19629,N_19657);
nor UO_260 (O_260,N_19763,N_19850);
nand UO_261 (O_261,N_19773,N_19763);
nand UO_262 (O_262,N_19638,N_19686);
nand UO_263 (O_263,N_19960,N_19880);
and UO_264 (O_264,N_19769,N_19838);
and UO_265 (O_265,N_19633,N_19876);
and UO_266 (O_266,N_19655,N_19989);
or UO_267 (O_267,N_19719,N_19711);
and UO_268 (O_268,N_19656,N_19805);
nor UO_269 (O_269,N_19881,N_19943);
and UO_270 (O_270,N_19907,N_19701);
nor UO_271 (O_271,N_19637,N_19740);
or UO_272 (O_272,N_19904,N_19694);
and UO_273 (O_273,N_19839,N_19917);
nor UO_274 (O_274,N_19720,N_19839);
and UO_275 (O_275,N_19882,N_19631);
nor UO_276 (O_276,N_19673,N_19699);
nand UO_277 (O_277,N_19748,N_19729);
or UO_278 (O_278,N_19841,N_19657);
nor UO_279 (O_279,N_19922,N_19828);
nand UO_280 (O_280,N_19989,N_19958);
nand UO_281 (O_281,N_19714,N_19957);
and UO_282 (O_282,N_19703,N_19855);
and UO_283 (O_283,N_19822,N_19969);
nand UO_284 (O_284,N_19782,N_19971);
or UO_285 (O_285,N_19955,N_19679);
or UO_286 (O_286,N_19790,N_19969);
or UO_287 (O_287,N_19828,N_19858);
xor UO_288 (O_288,N_19893,N_19614);
and UO_289 (O_289,N_19653,N_19789);
and UO_290 (O_290,N_19657,N_19649);
or UO_291 (O_291,N_19789,N_19641);
nand UO_292 (O_292,N_19646,N_19718);
or UO_293 (O_293,N_19699,N_19805);
and UO_294 (O_294,N_19990,N_19976);
nor UO_295 (O_295,N_19998,N_19749);
nand UO_296 (O_296,N_19669,N_19844);
or UO_297 (O_297,N_19787,N_19724);
nand UO_298 (O_298,N_19654,N_19768);
nor UO_299 (O_299,N_19873,N_19657);
xor UO_300 (O_300,N_19799,N_19970);
and UO_301 (O_301,N_19844,N_19682);
and UO_302 (O_302,N_19884,N_19900);
nor UO_303 (O_303,N_19683,N_19978);
nor UO_304 (O_304,N_19666,N_19966);
and UO_305 (O_305,N_19604,N_19652);
nor UO_306 (O_306,N_19895,N_19893);
nand UO_307 (O_307,N_19778,N_19800);
nor UO_308 (O_308,N_19641,N_19626);
nand UO_309 (O_309,N_19679,N_19807);
and UO_310 (O_310,N_19710,N_19714);
nor UO_311 (O_311,N_19753,N_19759);
nor UO_312 (O_312,N_19855,N_19688);
and UO_313 (O_313,N_19767,N_19653);
nand UO_314 (O_314,N_19754,N_19614);
or UO_315 (O_315,N_19664,N_19948);
nor UO_316 (O_316,N_19829,N_19928);
or UO_317 (O_317,N_19732,N_19814);
nor UO_318 (O_318,N_19764,N_19716);
nor UO_319 (O_319,N_19881,N_19928);
nor UO_320 (O_320,N_19845,N_19876);
nand UO_321 (O_321,N_19992,N_19782);
or UO_322 (O_322,N_19774,N_19930);
and UO_323 (O_323,N_19680,N_19740);
or UO_324 (O_324,N_19922,N_19975);
nor UO_325 (O_325,N_19764,N_19857);
or UO_326 (O_326,N_19844,N_19890);
nor UO_327 (O_327,N_19909,N_19908);
and UO_328 (O_328,N_19806,N_19973);
nor UO_329 (O_329,N_19633,N_19786);
or UO_330 (O_330,N_19914,N_19665);
nand UO_331 (O_331,N_19694,N_19657);
nand UO_332 (O_332,N_19688,N_19790);
nand UO_333 (O_333,N_19607,N_19635);
or UO_334 (O_334,N_19938,N_19879);
nor UO_335 (O_335,N_19975,N_19606);
and UO_336 (O_336,N_19885,N_19862);
nor UO_337 (O_337,N_19920,N_19881);
nor UO_338 (O_338,N_19846,N_19997);
or UO_339 (O_339,N_19956,N_19891);
and UO_340 (O_340,N_19881,N_19699);
nand UO_341 (O_341,N_19718,N_19736);
and UO_342 (O_342,N_19631,N_19841);
nand UO_343 (O_343,N_19644,N_19873);
nor UO_344 (O_344,N_19684,N_19961);
or UO_345 (O_345,N_19911,N_19890);
nor UO_346 (O_346,N_19748,N_19943);
and UO_347 (O_347,N_19698,N_19607);
nor UO_348 (O_348,N_19606,N_19826);
and UO_349 (O_349,N_19725,N_19672);
or UO_350 (O_350,N_19894,N_19628);
or UO_351 (O_351,N_19998,N_19949);
or UO_352 (O_352,N_19710,N_19716);
nor UO_353 (O_353,N_19712,N_19954);
nand UO_354 (O_354,N_19980,N_19705);
nand UO_355 (O_355,N_19979,N_19757);
nor UO_356 (O_356,N_19634,N_19619);
nor UO_357 (O_357,N_19651,N_19694);
nor UO_358 (O_358,N_19835,N_19911);
and UO_359 (O_359,N_19840,N_19838);
and UO_360 (O_360,N_19676,N_19762);
xnor UO_361 (O_361,N_19923,N_19940);
or UO_362 (O_362,N_19991,N_19937);
or UO_363 (O_363,N_19858,N_19854);
nor UO_364 (O_364,N_19724,N_19799);
or UO_365 (O_365,N_19913,N_19875);
nor UO_366 (O_366,N_19717,N_19754);
and UO_367 (O_367,N_19955,N_19627);
nand UO_368 (O_368,N_19904,N_19772);
or UO_369 (O_369,N_19959,N_19756);
or UO_370 (O_370,N_19626,N_19921);
nor UO_371 (O_371,N_19848,N_19953);
nand UO_372 (O_372,N_19831,N_19671);
and UO_373 (O_373,N_19735,N_19904);
nor UO_374 (O_374,N_19755,N_19849);
and UO_375 (O_375,N_19904,N_19618);
and UO_376 (O_376,N_19980,N_19812);
or UO_377 (O_377,N_19935,N_19678);
or UO_378 (O_378,N_19889,N_19610);
and UO_379 (O_379,N_19695,N_19657);
nor UO_380 (O_380,N_19770,N_19933);
and UO_381 (O_381,N_19940,N_19997);
or UO_382 (O_382,N_19643,N_19681);
nand UO_383 (O_383,N_19755,N_19778);
or UO_384 (O_384,N_19899,N_19606);
and UO_385 (O_385,N_19929,N_19943);
nor UO_386 (O_386,N_19874,N_19902);
nor UO_387 (O_387,N_19830,N_19975);
and UO_388 (O_388,N_19829,N_19728);
or UO_389 (O_389,N_19997,N_19906);
or UO_390 (O_390,N_19902,N_19814);
and UO_391 (O_391,N_19613,N_19625);
or UO_392 (O_392,N_19613,N_19683);
nor UO_393 (O_393,N_19889,N_19617);
nand UO_394 (O_394,N_19836,N_19899);
nor UO_395 (O_395,N_19814,N_19747);
and UO_396 (O_396,N_19676,N_19631);
nand UO_397 (O_397,N_19742,N_19657);
nor UO_398 (O_398,N_19610,N_19653);
nand UO_399 (O_399,N_19671,N_19676);
and UO_400 (O_400,N_19667,N_19705);
or UO_401 (O_401,N_19687,N_19985);
nor UO_402 (O_402,N_19726,N_19750);
nand UO_403 (O_403,N_19969,N_19877);
and UO_404 (O_404,N_19769,N_19780);
nand UO_405 (O_405,N_19685,N_19671);
and UO_406 (O_406,N_19689,N_19625);
nand UO_407 (O_407,N_19925,N_19613);
or UO_408 (O_408,N_19785,N_19606);
and UO_409 (O_409,N_19788,N_19765);
nand UO_410 (O_410,N_19683,N_19886);
nand UO_411 (O_411,N_19931,N_19650);
and UO_412 (O_412,N_19707,N_19671);
nor UO_413 (O_413,N_19905,N_19610);
xor UO_414 (O_414,N_19917,N_19947);
or UO_415 (O_415,N_19796,N_19606);
or UO_416 (O_416,N_19612,N_19604);
nor UO_417 (O_417,N_19653,N_19991);
and UO_418 (O_418,N_19872,N_19654);
or UO_419 (O_419,N_19993,N_19858);
or UO_420 (O_420,N_19620,N_19619);
or UO_421 (O_421,N_19933,N_19940);
nand UO_422 (O_422,N_19725,N_19809);
nor UO_423 (O_423,N_19761,N_19987);
and UO_424 (O_424,N_19760,N_19974);
nand UO_425 (O_425,N_19803,N_19715);
nand UO_426 (O_426,N_19927,N_19681);
nand UO_427 (O_427,N_19670,N_19608);
nor UO_428 (O_428,N_19985,N_19628);
and UO_429 (O_429,N_19908,N_19687);
and UO_430 (O_430,N_19952,N_19863);
nand UO_431 (O_431,N_19965,N_19747);
nor UO_432 (O_432,N_19680,N_19736);
nand UO_433 (O_433,N_19792,N_19801);
nor UO_434 (O_434,N_19754,N_19817);
or UO_435 (O_435,N_19641,N_19619);
and UO_436 (O_436,N_19608,N_19964);
nand UO_437 (O_437,N_19725,N_19791);
and UO_438 (O_438,N_19673,N_19927);
nor UO_439 (O_439,N_19670,N_19892);
or UO_440 (O_440,N_19614,N_19872);
or UO_441 (O_441,N_19942,N_19670);
or UO_442 (O_442,N_19684,N_19975);
nand UO_443 (O_443,N_19980,N_19637);
nand UO_444 (O_444,N_19665,N_19869);
nand UO_445 (O_445,N_19818,N_19613);
xor UO_446 (O_446,N_19864,N_19743);
and UO_447 (O_447,N_19913,N_19822);
nand UO_448 (O_448,N_19850,N_19886);
nand UO_449 (O_449,N_19778,N_19824);
or UO_450 (O_450,N_19798,N_19923);
and UO_451 (O_451,N_19701,N_19825);
nor UO_452 (O_452,N_19859,N_19919);
or UO_453 (O_453,N_19896,N_19690);
nand UO_454 (O_454,N_19981,N_19758);
or UO_455 (O_455,N_19645,N_19610);
nand UO_456 (O_456,N_19703,N_19951);
and UO_457 (O_457,N_19679,N_19646);
nor UO_458 (O_458,N_19979,N_19874);
nand UO_459 (O_459,N_19762,N_19871);
and UO_460 (O_460,N_19828,N_19654);
or UO_461 (O_461,N_19739,N_19695);
nor UO_462 (O_462,N_19836,N_19795);
nand UO_463 (O_463,N_19748,N_19828);
and UO_464 (O_464,N_19681,N_19799);
nor UO_465 (O_465,N_19728,N_19938);
nand UO_466 (O_466,N_19951,N_19808);
and UO_467 (O_467,N_19954,N_19988);
and UO_468 (O_468,N_19669,N_19728);
or UO_469 (O_469,N_19882,N_19801);
nor UO_470 (O_470,N_19889,N_19953);
or UO_471 (O_471,N_19652,N_19781);
nor UO_472 (O_472,N_19681,N_19836);
xnor UO_473 (O_473,N_19663,N_19947);
or UO_474 (O_474,N_19922,N_19638);
nand UO_475 (O_475,N_19983,N_19671);
nor UO_476 (O_476,N_19604,N_19869);
and UO_477 (O_477,N_19732,N_19677);
or UO_478 (O_478,N_19681,N_19873);
and UO_479 (O_479,N_19886,N_19984);
nand UO_480 (O_480,N_19773,N_19945);
or UO_481 (O_481,N_19669,N_19905);
nor UO_482 (O_482,N_19760,N_19810);
and UO_483 (O_483,N_19669,N_19924);
nand UO_484 (O_484,N_19652,N_19760);
nand UO_485 (O_485,N_19749,N_19728);
nand UO_486 (O_486,N_19768,N_19903);
nor UO_487 (O_487,N_19904,N_19740);
nor UO_488 (O_488,N_19826,N_19966);
and UO_489 (O_489,N_19868,N_19972);
nor UO_490 (O_490,N_19995,N_19771);
or UO_491 (O_491,N_19809,N_19904);
nor UO_492 (O_492,N_19884,N_19714);
nand UO_493 (O_493,N_19805,N_19927);
nand UO_494 (O_494,N_19766,N_19620);
or UO_495 (O_495,N_19646,N_19973);
nor UO_496 (O_496,N_19808,N_19853);
nor UO_497 (O_497,N_19859,N_19760);
nor UO_498 (O_498,N_19933,N_19792);
xor UO_499 (O_499,N_19996,N_19662);
nand UO_500 (O_500,N_19661,N_19943);
and UO_501 (O_501,N_19735,N_19996);
or UO_502 (O_502,N_19997,N_19622);
nor UO_503 (O_503,N_19600,N_19805);
and UO_504 (O_504,N_19811,N_19621);
nand UO_505 (O_505,N_19822,N_19880);
nand UO_506 (O_506,N_19623,N_19765);
or UO_507 (O_507,N_19854,N_19851);
or UO_508 (O_508,N_19714,N_19888);
nand UO_509 (O_509,N_19808,N_19980);
and UO_510 (O_510,N_19739,N_19957);
nand UO_511 (O_511,N_19938,N_19724);
nor UO_512 (O_512,N_19962,N_19940);
or UO_513 (O_513,N_19702,N_19673);
or UO_514 (O_514,N_19924,N_19611);
nand UO_515 (O_515,N_19997,N_19746);
nor UO_516 (O_516,N_19928,N_19748);
and UO_517 (O_517,N_19605,N_19802);
and UO_518 (O_518,N_19616,N_19631);
nor UO_519 (O_519,N_19972,N_19606);
nor UO_520 (O_520,N_19741,N_19620);
nand UO_521 (O_521,N_19851,N_19970);
nand UO_522 (O_522,N_19859,N_19645);
nand UO_523 (O_523,N_19863,N_19824);
nand UO_524 (O_524,N_19746,N_19636);
and UO_525 (O_525,N_19783,N_19767);
nor UO_526 (O_526,N_19690,N_19810);
and UO_527 (O_527,N_19616,N_19736);
nor UO_528 (O_528,N_19914,N_19610);
nand UO_529 (O_529,N_19640,N_19795);
nor UO_530 (O_530,N_19664,N_19614);
and UO_531 (O_531,N_19689,N_19797);
nand UO_532 (O_532,N_19811,N_19656);
and UO_533 (O_533,N_19749,N_19732);
and UO_534 (O_534,N_19984,N_19977);
nand UO_535 (O_535,N_19832,N_19655);
nor UO_536 (O_536,N_19847,N_19866);
or UO_537 (O_537,N_19660,N_19620);
nand UO_538 (O_538,N_19848,N_19791);
and UO_539 (O_539,N_19615,N_19890);
nand UO_540 (O_540,N_19719,N_19666);
or UO_541 (O_541,N_19928,N_19963);
nor UO_542 (O_542,N_19932,N_19918);
or UO_543 (O_543,N_19668,N_19826);
nor UO_544 (O_544,N_19900,N_19801);
and UO_545 (O_545,N_19785,N_19780);
or UO_546 (O_546,N_19739,N_19871);
and UO_547 (O_547,N_19856,N_19880);
or UO_548 (O_548,N_19653,N_19915);
nand UO_549 (O_549,N_19611,N_19616);
nor UO_550 (O_550,N_19985,N_19888);
nand UO_551 (O_551,N_19899,N_19623);
nand UO_552 (O_552,N_19683,N_19807);
or UO_553 (O_553,N_19951,N_19770);
nand UO_554 (O_554,N_19629,N_19966);
nor UO_555 (O_555,N_19911,N_19715);
nor UO_556 (O_556,N_19850,N_19853);
or UO_557 (O_557,N_19898,N_19863);
or UO_558 (O_558,N_19916,N_19900);
and UO_559 (O_559,N_19978,N_19761);
or UO_560 (O_560,N_19893,N_19900);
nor UO_561 (O_561,N_19968,N_19821);
nand UO_562 (O_562,N_19911,N_19651);
nand UO_563 (O_563,N_19625,N_19874);
xor UO_564 (O_564,N_19911,N_19698);
and UO_565 (O_565,N_19661,N_19761);
and UO_566 (O_566,N_19628,N_19915);
and UO_567 (O_567,N_19758,N_19665);
or UO_568 (O_568,N_19643,N_19717);
or UO_569 (O_569,N_19984,N_19839);
nand UO_570 (O_570,N_19629,N_19901);
and UO_571 (O_571,N_19804,N_19886);
nor UO_572 (O_572,N_19932,N_19855);
and UO_573 (O_573,N_19698,N_19725);
nor UO_574 (O_574,N_19726,N_19899);
nor UO_575 (O_575,N_19946,N_19851);
nand UO_576 (O_576,N_19871,N_19897);
nand UO_577 (O_577,N_19641,N_19925);
nand UO_578 (O_578,N_19763,N_19614);
or UO_579 (O_579,N_19817,N_19964);
nand UO_580 (O_580,N_19928,N_19783);
nand UO_581 (O_581,N_19775,N_19738);
nor UO_582 (O_582,N_19753,N_19826);
or UO_583 (O_583,N_19828,N_19733);
nor UO_584 (O_584,N_19941,N_19720);
nand UO_585 (O_585,N_19661,N_19611);
or UO_586 (O_586,N_19828,N_19628);
and UO_587 (O_587,N_19856,N_19897);
nand UO_588 (O_588,N_19671,N_19900);
nand UO_589 (O_589,N_19990,N_19690);
nor UO_590 (O_590,N_19932,N_19610);
nor UO_591 (O_591,N_19870,N_19892);
or UO_592 (O_592,N_19799,N_19965);
or UO_593 (O_593,N_19864,N_19682);
or UO_594 (O_594,N_19672,N_19666);
nand UO_595 (O_595,N_19864,N_19961);
nand UO_596 (O_596,N_19670,N_19718);
nand UO_597 (O_597,N_19988,N_19745);
or UO_598 (O_598,N_19769,N_19619);
nor UO_599 (O_599,N_19911,N_19923);
nand UO_600 (O_600,N_19729,N_19837);
or UO_601 (O_601,N_19603,N_19803);
nor UO_602 (O_602,N_19849,N_19932);
nand UO_603 (O_603,N_19680,N_19815);
nor UO_604 (O_604,N_19830,N_19689);
and UO_605 (O_605,N_19798,N_19699);
nand UO_606 (O_606,N_19819,N_19646);
or UO_607 (O_607,N_19886,N_19888);
and UO_608 (O_608,N_19891,N_19941);
nand UO_609 (O_609,N_19702,N_19846);
nor UO_610 (O_610,N_19671,N_19626);
and UO_611 (O_611,N_19920,N_19853);
nand UO_612 (O_612,N_19780,N_19936);
nor UO_613 (O_613,N_19721,N_19915);
and UO_614 (O_614,N_19915,N_19670);
and UO_615 (O_615,N_19742,N_19785);
nor UO_616 (O_616,N_19667,N_19771);
nor UO_617 (O_617,N_19698,N_19890);
and UO_618 (O_618,N_19604,N_19864);
nand UO_619 (O_619,N_19963,N_19651);
or UO_620 (O_620,N_19675,N_19674);
nor UO_621 (O_621,N_19654,N_19661);
nor UO_622 (O_622,N_19676,N_19860);
nor UO_623 (O_623,N_19968,N_19675);
nand UO_624 (O_624,N_19739,N_19855);
nor UO_625 (O_625,N_19815,N_19814);
nor UO_626 (O_626,N_19694,N_19945);
and UO_627 (O_627,N_19648,N_19841);
and UO_628 (O_628,N_19699,N_19695);
and UO_629 (O_629,N_19606,N_19878);
and UO_630 (O_630,N_19979,N_19789);
nand UO_631 (O_631,N_19606,N_19981);
nand UO_632 (O_632,N_19620,N_19864);
or UO_633 (O_633,N_19662,N_19925);
or UO_634 (O_634,N_19778,N_19650);
and UO_635 (O_635,N_19874,N_19914);
or UO_636 (O_636,N_19812,N_19975);
and UO_637 (O_637,N_19643,N_19638);
nor UO_638 (O_638,N_19732,N_19896);
nor UO_639 (O_639,N_19913,N_19784);
or UO_640 (O_640,N_19682,N_19785);
nand UO_641 (O_641,N_19701,N_19877);
and UO_642 (O_642,N_19885,N_19889);
and UO_643 (O_643,N_19649,N_19666);
nor UO_644 (O_644,N_19654,N_19762);
nand UO_645 (O_645,N_19989,N_19797);
or UO_646 (O_646,N_19643,N_19713);
nor UO_647 (O_647,N_19784,N_19701);
nand UO_648 (O_648,N_19638,N_19805);
nor UO_649 (O_649,N_19600,N_19817);
nor UO_650 (O_650,N_19659,N_19997);
and UO_651 (O_651,N_19848,N_19664);
xnor UO_652 (O_652,N_19998,N_19880);
and UO_653 (O_653,N_19946,N_19691);
or UO_654 (O_654,N_19638,N_19659);
nor UO_655 (O_655,N_19956,N_19781);
nor UO_656 (O_656,N_19993,N_19997);
nand UO_657 (O_657,N_19604,N_19984);
nand UO_658 (O_658,N_19669,N_19625);
and UO_659 (O_659,N_19708,N_19642);
or UO_660 (O_660,N_19968,N_19663);
nand UO_661 (O_661,N_19936,N_19664);
nand UO_662 (O_662,N_19660,N_19650);
nand UO_663 (O_663,N_19963,N_19724);
nand UO_664 (O_664,N_19853,N_19675);
and UO_665 (O_665,N_19836,N_19832);
or UO_666 (O_666,N_19669,N_19705);
nand UO_667 (O_667,N_19851,N_19941);
and UO_668 (O_668,N_19861,N_19794);
or UO_669 (O_669,N_19661,N_19651);
or UO_670 (O_670,N_19765,N_19618);
or UO_671 (O_671,N_19813,N_19675);
and UO_672 (O_672,N_19648,N_19967);
and UO_673 (O_673,N_19884,N_19645);
nor UO_674 (O_674,N_19888,N_19665);
nor UO_675 (O_675,N_19953,N_19816);
and UO_676 (O_676,N_19741,N_19952);
and UO_677 (O_677,N_19939,N_19990);
nand UO_678 (O_678,N_19608,N_19647);
nand UO_679 (O_679,N_19815,N_19856);
nand UO_680 (O_680,N_19638,N_19656);
nand UO_681 (O_681,N_19984,N_19988);
nor UO_682 (O_682,N_19743,N_19904);
nor UO_683 (O_683,N_19638,N_19965);
nand UO_684 (O_684,N_19978,N_19843);
nor UO_685 (O_685,N_19823,N_19672);
nor UO_686 (O_686,N_19748,N_19960);
and UO_687 (O_687,N_19938,N_19714);
nand UO_688 (O_688,N_19817,N_19866);
and UO_689 (O_689,N_19637,N_19874);
and UO_690 (O_690,N_19628,N_19944);
and UO_691 (O_691,N_19693,N_19708);
and UO_692 (O_692,N_19972,N_19971);
nor UO_693 (O_693,N_19837,N_19685);
nand UO_694 (O_694,N_19747,N_19925);
nand UO_695 (O_695,N_19716,N_19645);
nor UO_696 (O_696,N_19852,N_19642);
nand UO_697 (O_697,N_19719,N_19627);
nand UO_698 (O_698,N_19936,N_19725);
nor UO_699 (O_699,N_19948,N_19900);
nand UO_700 (O_700,N_19946,N_19846);
or UO_701 (O_701,N_19742,N_19949);
xor UO_702 (O_702,N_19683,N_19967);
nor UO_703 (O_703,N_19938,N_19734);
and UO_704 (O_704,N_19995,N_19605);
or UO_705 (O_705,N_19782,N_19956);
and UO_706 (O_706,N_19922,N_19980);
nand UO_707 (O_707,N_19621,N_19605);
and UO_708 (O_708,N_19913,N_19871);
or UO_709 (O_709,N_19999,N_19804);
nor UO_710 (O_710,N_19885,N_19777);
and UO_711 (O_711,N_19657,N_19914);
and UO_712 (O_712,N_19760,N_19973);
and UO_713 (O_713,N_19724,N_19858);
nor UO_714 (O_714,N_19626,N_19822);
nand UO_715 (O_715,N_19897,N_19847);
or UO_716 (O_716,N_19740,N_19885);
nand UO_717 (O_717,N_19805,N_19760);
nor UO_718 (O_718,N_19810,N_19836);
nand UO_719 (O_719,N_19979,N_19669);
and UO_720 (O_720,N_19616,N_19648);
nor UO_721 (O_721,N_19614,N_19922);
or UO_722 (O_722,N_19869,N_19916);
xor UO_723 (O_723,N_19974,N_19992);
nand UO_724 (O_724,N_19621,N_19645);
or UO_725 (O_725,N_19659,N_19709);
and UO_726 (O_726,N_19709,N_19937);
nor UO_727 (O_727,N_19829,N_19920);
or UO_728 (O_728,N_19752,N_19935);
and UO_729 (O_729,N_19944,N_19903);
or UO_730 (O_730,N_19889,N_19982);
and UO_731 (O_731,N_19687,N_19689);
xor UO_732 (O_732,N_19719,N_19768);
nand UO_733 (O_733,N_19978,N_19910);
and UO_734 (O_734,N_19974,N_19912);
or UO_735 (O_735,N_19912,N_19799);
nor UO_736 (O_736,N_19846,N_19781);
nor UO_737 (O_737,N_19634,N_19754);
nand UO_738 (O_738,N_19951,N_19655);
nor UO_739 (O_739,N_19632,N_19670);
and UO_740 (O_740,N_19606,N_19932);
nor UO_741 (O_741,N_19839,N_19866);
nor UO_742 (O_742,N_19937,N_19625);
nand UO_743 (O_743,N_19973,N_19849);
and UO_744 (O_744,N_19776,N_19810);
nand UO_745 (O_745,N_19785,N_19782);
nand UO_746 (O_746,N_19671,N_19834);
and UO_747 (O_747,N_19997,N_19756);
or UO_748 (O_748,N_19694,N_19704);
and UO_749 (O_749,N_19892,N_19612);
nor UO_750 (O_750,N_19882,N_19742);
nand UO_751 (O_751,N_19622,N_19820);
and UO_752 (O_752,N_19843,N_19872);
nor UO_753 (O_753,N_19762,N_19907);
or UO_754 (O_754,N_19969,N_19750);
and UO_755 (O_755,N_19951,N_19986);
nor UO_756 (O_756,N_19638,N_19772);
and UO_757 (O_757,N_19759,N_19818);
nand UO_758 (O_758,N_19679,N_19717);
and UO_759 (O_759,N_19751,N_19908);
and UO_760 (O_760,N_19803,N_19806);
nand UO_761 (O_761,N_19869,N_19931);
or UO_762 (O_762,N_19979,N_19953);
nor UO_763 (O_763,N_19775,N_19869);
nand UO_764 (O_764,N_19828,N_19736);
or UO_765 (O_765,N_19695,N_19837);
nand UO_766 (O_766,N_19793,N_19768);
or UO_767 (O_767,N_19743,N_19911);
or UO_768 (O_768,N_19618,N_19759);
or UO_769 (O_769,N_19615,N_19683);
or UO_770 (O_770,N_19622,N_19951);
and UO_771 (O_771,N_19660,N_19688);
or UO_772 (O_772,N_19758,N_19792);
nand UO_773 (O_773,N_19667,N_19929);
nor UO_774 (O_774,N_19834,N_19708);
or UO_775 (O_775,N_19823,N_19810);
nor UO_776 (O_776,N_19823,N_19709);
and UO_777 (O_777,N_19648,N_19984);
nand UO_778 (O_778,N_19728,N_19735);
nor UO_779 (O_779,N_19781,N_19726);
nand UO_780 (O_780,N_19759,N_19606);
nand UO_781 (O_781,N_19676,N_19638);
or UO_782 (O_782,N_19818,N_19602);
or UO_783 (O_783,N_19883,N_19713);
nor UO_784 (O_784,N_19903,N_19917);
nor UO_785 (O_785,N_19988,N_19671);
and UO_786 (O_786,N_19627,N_19893);
nand UO_787 (O_787,N_19705,N_19784);
and UO_788 (O_788,N_19775,N_19770);
nand UO_789 (O_789,N_19956,N_19737);
nor UO_790 (O_790,N_19856,N_19789);
and UO_791 (O_791,N_19809,N_19827);
nor UO_792 (O_792,N_19792,N_19693);
or UO_793 (O_793,N_19671,N_19923);
nor UO_794 (O_794,N_19973,N_19926);
and UO_795 (O_795,N_19917,N_19875);
nand UO_796 (O_796,N_19687,N_19751);
and UO_797 (O_797,N_19796,N_19683);
and UO_798 (O_798,N_19627,N_19976);
or UO_799 (O_799,N_19989,N_19763);
and UO_800 (O_800,N_19836,N_19671);
nand UO_801 (O_801,N_19739,N_19780);
or UO_802 (O_802,N_19708,N_19813);
nand UO_803 (O_803,N_19871,N_19610);
nand UO_804 (O_804,N_19765,N_19881);
or UO_805 (O_805,N_19925,N_19815);
nand UO_806 (O_806,N_19607,N_19954);
or UO_807 (O_807,N_19986,N_19910);
or UO_808 (O_808,N_19880,N_19626);
xnor UO_809 (O_809,N_19963,N_19801);
nor UO_810 (O_810,N_19704,N_19785);
xor UO_811 (O_811,N_19746,N_19941);
and UO_812 (O_812,N_19999,N_19883);
or UO_813 (O_813,N_19971,N_19900);
nand UO_814 (O_814,N_19778,N_19749);
nor UO_815 (O_815,N_19647,N_19674);
and UO_816 (O_816,N_19914,N_19689);
or UO_817 (O_817,N_19726,N_19893);
nor UO_818 (O_818,N_19614,N_19799);
and UO_819 (O_819,N_19644,N_19986);
and UO_820 (O_820,N_19640,N_19688);
nand UO_821 (O_821,N_19822,N_19991);
or UO_822 (O_822,N_19953,N_19944);
nand UO_823 (O_823,N_19780,N_19812);
and UO_824 (O_824,N_19936,N_19921);
or UO_825 (O_825,N_19966,N_19615);
or UO_826 (O_826,N_19935,N_19742);
nor UO_827 (O_827,N_19838,N_19772);
and UO_828 (O_828,N_19703,N_19957);
or UO_829 (O_829,N_19761,N_19758);
nor UO_830 (O_830,N_19665,N_19887);
and UO_831 (O_831,N_19666,N_19791);
and UO_832 (O_832,N_19738,N_19812);
and UO_833 (O_833,N_19870,N_19967);
nand UO_834 (O_834,N_19921,N_19892);
and UO_835 (O_835,N_19633,N_19725);
or UO_836 (O_836,N_19824,N_19713);
and UO_837 (O_837,N_19618,N_19736);
and UO_838 (O_838,N_19625,N_19887);
or UO_839 (O_839,N_19981,N_19676);
or UO_840 (O_840,N_19908,N_19789);
or UO_841 (O_841,N_19788,N_19662);
or UO_842 (O_842,N_19643,N_19811);
and UO_843 (O_843,N_19613,N_19782);
and UO_844 (O_844,N_19769,N_19820);
or UO_845 (O_845,N_19971,N_19650);
or UO_846 (O_846,N_19971,N_19994);
and UO_847 (O_847,N_19764,N_19956);
and UO_848 (O_848,N_19863,N_19742);
nor UO_849 (O_849,N_19740,N_19908);
nand UO_850 (O_850,N_19758,N_19679);
nor UO_851 (O_851,N_19909,N_19741);
nand UO_852 (O_852,N_19790,N_19867);
and UO_853 (O_853,N_19888,N_19659);
or UO_854 (O_854,N_19951,N_19965);
nor UO_855 (O_855,N_19894,N_19942);
nor UO_856 (O_856,N_19811,N_19870);
nor UO_857 (O_857,N_19720,N_19844);
nor UO_858 (O_858,N_19924,N_19681);
nor UO_859 (O_859,N_19743,N_19967);
nand UO_860 (O_860,N_19803,N_19902);
or UO_861 (O_861,N_19945,N_19744);
and UO_862 (O_862,N_19903,N_19821);
nor UO_863 (O_863,N_19758,N_19802);
nand UO_864 (O_864,N_19884,N_19809);
xnor UO_865 (O_865,N_19784,N_19903);
nand UO_866 (O_866,N_19686,N_19920);
nand UO_867 (O_867,N_19942,N_19719);
and UO_868 (O_868,N_19862,N_19929);
and UO_869 (O_869,N_19851,N_19886);
nor UO_870 (O_870,N_19630,N_19725);
and UO_871 (O_871,N_19673,N_19711);
nand UO_872 (O_872,N_19708,N_19775);
and UO_873 (O_873,N_19935,N_19899);
and UO_874 (O_874,N_19828,N_19740);
nor UO_875 (O_875,N_19846,N_19817);
nor UO_876 (O_876,N_19838,N_19876);
nand UO_877 (O_877,N_19820,N_19631);
or UO_878 (O_878,N_19674,N_19915);
nor UO_879 (O_879,N_19944,N_19669);
nand UO_880 (O_880,N_19680,N_19899);
nor UO_881 (O_881,N_19693,N_19874);
nand UO_882 (O_882,N_19737,N_19778);
nor UO_883 (O_883,N_19930,N_19974);
nor UO_884 (O_884,N_19796,N_19870);
nor UO_885 (O_885,N_19789,N_19719);
or UO_886 (O_886,N_19972,N_19818);
nand UO_887 (O_887,N_19816,N_19692);
or UO_888 (O_888,N_19660,N_19711);
or UO_889 (O_889,N_19827,N_19947);
nand UO_890 (O_890,N_19624,N_19686);
nor UO_891 (O_891,N_19988,N_19746);
xor UO_892 (O_892,N_19994,N_19693);
xnor UO_893 (O_893,N_19822,N_19623);
or UO_894 (O_894,N_19879,N_19662);
xnor UO_895 (O_895,N_19906,N_19774);
nor UO_896 (O_896,N_19825,N_19931);
nor UO_897 (O_897,N_19844,N_19731);
and UO_898 (O_898,N_19872,N_19780);
nand UO_899 (O_899,N_19713,N_19960);
and UO_900 (O_900,N_19972,N_19663);
or UO_901 (O_901,N_19862,N_19772);
nor UO_902 (O_902,N_19707,N_19808);
and UO_903 (O_903,N_19891,N_19650);
nor UO_904 (O_904,N_19831,N_19982);
nor UO_905 (O_905,N_19663,N_19603);
and UO_906 (O_906,N_19930,N_19862);
nor UO_907 (O_907,N_19615,N_19769);
nand UO_908 (O_908,N_19672,N_19997);
and UO_909 (O_909,N_19711,N_19800);
or UO_910 (O_910,N_19944,N_19710);
and UO_911 (O_911,N_19799,N_19978);
nor UO_912 (O_912,N_19718,N_19600);
nor UO_913 (O_913,N_19820,N_19815);
nand UO_914 (O_914,N_19870,N_19915);
nand UO_915 (O_915,N_19899,N_19676);
nand UO_916 (O_916,N_19608,N_19828);
and UO_917 (O_917,N_19700,N_19900);
or UO_918 (O_918,N_19664,N_19670);
and UO_919 (O_919,N_19771,N_19627);
and UO_920 (O_920,N_19696,N_19603);
nand UO_921 (O_921,N_19749,N_19792);
nand UO_922 (O_922,N_19928,N_19651);
and UO_923 (O_923,N_19817,N_19956);
nand UO_924 (O_924,N_19880,N_19940);
and UO_925 (O_925,N_19800,N_19773);
nor UO_926 (O_926,N_19875,N_19967);
and UO_927 (O_927,N_19998,N_19858);
nand UO_928 (O_928,N_19692,N_19957);
nand UO_929 (O_929,N_19770,N_19898);
and UO_930 (O_930,N_19644,N_19908);
and UO_931 (O_931,N_19835,N_19649);
nor UO_932 (O_932,N_19917,N_19974);
nor UO_933 (O_933,N_19880,N_19874);
nand UO_934 (O_934,N_19916,N_19689);
and UO_935 (O_935,N_19914,N_19802);
and UO_936 (O_936,N_19894,N_19926);
nand UO_937 (O_937,N_19676,N_19793);
and UO_938 (O_938,N_19820,N_19969);
nand UO_939 (O_939,N_19725,N_19908);
or UO_940 (O_940,N_19838,N_19922);
or UO_941 (O_941,N_19665,N_19651);
and UO_942 (O_942,N_19998,N_19788);
and UO_943 (O_943,N_19913,N_19789);
and UO_944 (O_944,N_19703,N_19832);
or UO_945 (O_945,N_19726,N_19870);
and UO_946 (O_946,N_19749,N_19995);
nand UO_947 (O_947,N_19706,N_19614);
or UO_948 (O_948,N_19662,N_19617);
nand UO_949 (O_949,N_19812,N_19686);
and UO_950 (O_950,N_19709,N_19983);
and UO_951 (O_951,N_19635,N_19698);
and UO_952 (O_952,N_19883,N_19712);
and UO_953 (O_953,N_19855,N_19966);
and UO_954 (O_954,N_19873,N_19828);
and UO_955 (O_955,N_19627,N_19718);
or UO_956 (O_956,N_19930,N_19728);
and UO_957 (O_957,N_19696,N_19894);
or UO_958 (O_958,N_19736,N_19964);
and UO_959 (O_959,N_19747,N_19803);
or UO_960 (O_960,N_19699,N_19954);
nand UO_961 (O_961,N_19768,N_19811);
nand UO_962 (O_962,N_19740,N_19910);
nor UO_963 (O_963,N_19655,N_19886);
or UO_964 (O_964,N_19761,N_19871);
nand UO_965 (O_965,N_19909,N_19836);
and UO_966 (O_966,N_19741,N_19781);
nor UO_967 (O_967,N_19852,N_19860);
and UO_968 (O_968,N_19841,N_19815);
and UO_969 (O_969,N_19669,N_19863);
nor UO_970 (O_970,N_19688,N_19745);
nor UO_971 (O_971,N_19669,N_19965);
or UO_972 (O_972,N_19780,N_19881);
or UO_973 (O_973,N_19634,N_19942);
and UO_974 (O_974,N_19832,N_19945);
nand UO_975 (O_975,N_19954,N_19675);
or UO_976 (O_976,N_19747,N_19749);
or UO_977 (O_977,N_19663,N_19651);
nor UO_978 (O_978,N_19893,N_19991);
or UO_979 (O_979,N_19724,N_19882);
and UO_980 (O_980,N_19621,N_19979);
nor UO_981 (O_981,N_19804,N_19600);
and UO_982 (O_982,N_19717,N_19945);
nor UO_983 (O_983,N_19804,N_19991);
or UO_984 (O_984,N_19802,N_19934);
and UO_985 (O_985,N_19708,N_19763);
or UO_986 (O_986,N_19682,N_19749);
and UO_987 (O_987,N_19735,N_19989);
nor UO_988 (O_988,N_19909,N_19693);
nor UO_989 (O_989,N_19843,N_19874);
and UO_990 (O_990,N_19723,N_19676);
nor UO_991 (O_991,N_19846,N_19924);
nand UO_992 (O_992,N_19757,N_19671);
nor UO_993 (O_993,N_19879,N_19737);
nand UO_994 (O_994,N_19735,N_19806);
nor UO_995 (O_995,N_19921,N_19661);
or UO_996 (O_996,N_19982,N_19636);
nand UO_997 (O_997,N_19765,N_19992);
nor UO_998 (O_998,N_19789,N_19704);
and UO_999 (O_999,N_19687,N_19909);
or UO_1000 (O_1000,N_19885,N_19902);
and UO_1001 (O_1001,N_19619,N_19719);
or UO_1002 (O_1002,N_19799,N_19762);
or UO_1003 (O_1003,N_19636,N_19863);
or UO_1004 (O_1004,N_19834,N_19920);
nor UO_1005 (O_1005,N_19658,N_19872);
or UO_1006 (O_1006,N_19657,N_19913);
or UO_1007 (O_1007,N_19898,N_19667);
or UO_1008 (O_1008,N_19794,N_19612);
or UO_1009 (O_1009,N_19753,N_19652);
or UO_1010 (O_1010,N_19812,N_19915);
and UO_1011 (O_1011,N_19746,N_19771);
or UO_1012 (O_1012,N_19795,N_19867);
or UO_1013 (O_1013,N_19753,N_19883);
nor UO_1014 (O_1014,N_19983,N_19770);
or UO_1015 (O_1015,N_19870,N_19909);
or UO_1016 (O_1016,N_19973,N_19846);
and UO_1017 (O_1017,N_19729,N_19814);
nand UO_1018 (O_1018,N_19792,N_19877);
and UO_1019 (O_1019,N_19687,N_19812);
or UO_1020 (O_1020,N_19854,N_19617);
nor UO_1021 (O_1021,N_19793,N_19754);
or UO_1022 (O_1022,N_19924,N_19890);
and UO_1023 (O_1023,N_19886,N_19866);
and UO_1024 (O_1024,N_19976,N_19735);
nor UO_1025 (O_1025,N_19930,N_19834);
or UO_1026 (O_1026,N_19603,N_19732);
or UO_1027 (O_1027,N_19849,N_19735);
nand UO_1028 (O_1028,N_19635,N_19705);
and UO_1029 (O_1029,N_19994,N_19992);
nand UO_1030 (O_1030,N_19705,N_19803);
nor UO_1031 (O_1031,N_19898,N_19987);
nor UO_1032 (O_1032,N_19639,N_19640);
nand UO_1033 (O_1033,N_19936,N_19826);
nor UO_1034 (O_1034,N_19649,N_19781);
nor UO_1035 (O_1035,N_19832,N_19782);
nand UO_1036 (O_1036,N_19718,N_19974);
nand UO_1037 (O_1037,N_19944,N_19956);
or UO_1038 (O_1038,N_19874,N_19965);
and UO_1039 (O_1039,N_19774,N_19771);
nor UO_1040 (O_1040,N_19710,N_19779);
or UO_1041 (O_1041,N_19883,N_19635);
nor UO_1042 (O_1042,N_19800,N_19919);
or UO_1043 (O_1043,N_19819,N_19949);
or UO_1044 (O_1044,N_19625,N_19876);
nor UO_1045 (O_1045,N_19847,N_19780);
nor UO_1046 (O_1046,N_19624,N_19679);
or UO_1047 (O_1047,N_19962,N_19971);
and UO_1048 (O_1048,N_19657,N_19613);
nor UO_1049 (O_1049,N_19954,N_19882);
or UO_1050 (O_1050,N_19756,N_19901);
nand UO_1051 (O_1051,N_19880,N_19797);
and UO_1052 (O_1052,N_19611,N_19861);
and UO_1053 (O_1053,N_19669,N_19731);
or UO_1054 (O_1054,N_19711,N_19830);
nor UO_1055 (O_1055,N_19771,N_19983);
nand UO_1056 (O_1056,N_19889,N_19629);
and UO_1057 (O_1057,N_19830,N_19871);
nand UO_1058 (O_1058,N_19629,N_19748);
and UO_1059 (O_1059,N_19748,N_19953);
and UO_1060 (O_1060,N_19794,N_19620);
and UO_1061 (O_1061,N_19652,N_19669);
nand UO_1062 (O_1062,N_19665,N_19920);
nand UO_1063 (O_1063,N_19928,N_19697);
and UO_1064 (O_1064,N_19793,N_19954);
nor UO_1065 (O_1065,N_19755,N_19723);
nor UO_1066 (O_1066,N_19900,N_19903);
nand UO_1067 (O_1067,N_19648,N_19777);
nor UO_1068 (O_1068,N_19977,N_19780);
and UO_1069 (O_1069,N_19769,N_19639);
or UO_1070 (O_1070,N_19790,N_19623);
nor UO_1071 (O_1071,N_19896,N_19811);
and UO_1072 (O_1072,N_19627,N_19729);
nor UO_1073 (O_1073,N_19918,N_19751);
nor UO_1074 (O_1074,N_19734,N_19656);
nand UO_1075 (O_1075,N_19839,N_19620);
and UO_1076 (O_1076,N_19738,N_19654);
and UO_1077 (O_1077,N_19707,N_19841);
nand UO_1078 (O_1078,N_19718,N_19979);
nand UO_1079 (O_1079,N_19928,N_19887);
nand UO_1080 (O_1080,N_19907,N_19802);
and UO_1081 (O_1081,N_19963,N_19961);
or UO_1082 (O_1082,N_19840,N_19645);
nor UO_1083 (O_1083,N_19784,N_19678);
and UO_1084 (O_1084,N_19747,N_19742);
nor UO_1085 (O_1085,N_19742,N_19957);
and UO_1086 (O_1086,N_19951,N_19998);
or UO_1087 (O_1087,N_19616,N_19749);
nand UO_1088 (O_1088,N_19850,N_19611);
nor UO_1089 (O_1089,N_19666,N_19742);
or UO_1090 (O_1090,N_19828,N_19774);
and UO_1091 (O_1091,N_19934,N_19836);
and UO_1092 (O_1092,N_19854,N_19661);
nand UO_1093 (O_1093,N_19827,N_19644);
or UO_1094 (O_1094,N_19935,N_19859);
and UO_1095 (O_1095,N_19994,N_19949);
or UO_1096 (O_1096,N_19769,N_19646);
nor UO_1097 (O_1097,N_19881,N_19804);
nand UO_1098 (O_1098,N_19755,N_19721);
nand UO_1099 (O_1099,N_19836,N_19931);
nor UO_1100 (O_1100,N_19820,N_19714);
nand UO_1101 (O_1101,N_19914,N_19804);
nor UO_1102 (O_1102,N_19968,N_19775);
nor UO_1103 (O_1103,N_19661,N_19954);
nor UO_1104 (O_1104,N_19971,N_19865);
or UO_1105 (O_1105,N_19657,N_19852);
nor UO_1106 (O_1106,N_19710,N_19742);
nor UO_1107 (O_1107,N_19851,N_19629);
and UO_1108 (O_1108,N_19745,N_19723);
nor UO_1109 (O_1109,N_19730,N_19754);
nand UO_1110 (O_1110,N_19980,N_19757);
or UO_1111 (O_1111,N_19628,N_19606);
nand UO_1112 (O_1112,N_19820,N_19789);
nor UO_1113 (O_1113,N_19692,N_19776);
nor UO_1114 (O_1114,N_19991,N_19680);
nor UO_1115 (O_1115,N_19894,N_19609);
nor UO_1116 (O_1116,N_19907,N_19635);
nand UO_1117 (O_1117,N_19745,N_19886);
nand UO_1118 (O_1118,N_19908,N_19897);
or UO_1119 (O_1119,N_19930,N_19735);
nor UO_1120 (O_1120,N_19670,N_19821);
nand UO_1121 (O_1121,N_19925,N_19645);
and UO_1122 (O_1122,N_19906,N_19674);
and UO_1123 (O_1123,N_19696,N_19997);
nor UO_1124 (O_1124,N_19638,N_19663);
nand UO_1125 (O_1125,N_19720,N_19723);
nor UO_1126 (O_1126,N_19934,N_19972);
nand UO_1127 (O_1127,N_19979,N_19792);
nand UO_1128 (O_1128,N_19602,N_19622);
and UO_1129 (O_1129,N_19662,N_19831);
and UO_1130 (O_1130,N_19922,N_19953);
nand UO_1131 (O_1131,N_19717,N_19811);
nand UO_1132 (O_1132,N_19741,N_19641);
nor UO_1133 (O_1133,N_19785,N_19903);
nor UO_1134 (O_1134,N_19810,N_19848);
nor UO_1135 (O_1135,N_19845,N_19840);
and UO_1136 (O_1136,N_19824,N_19716);
nor UO_1137 (O_1137,N_19847,N_19972);
nor UO_1138 (O_1138,N_19915,N_19874);
nand UO_1139 (O_1139,N_19721,N_19883);
or UO_1140 (O_1140,N_19953,N_19885);
and UO_1141 (O_1141,N_19762,N_19981);
nor UO_1142 (O_1142,N_19812,N_19749);
nor UO_1143 (O_1143,N_19736,N_19842);
nor UO_1144 (O_1144,N_19846,N_19809);
nand UO_1145 (O_1145,N_19711,N_19930);
or UO_1146 (O_1146,N_19887,N_19800);
nor UO_1147 (O_1147,N_19841,N_19916);
or UO_1148 (O_1148,N_19712,N_19890);
and UO_1149 (O_1149,N_19994,N_19819);
or UO_1150 (O_1150,N_19623,N_19932);
nor UO_1151 (O_1151,N_19891,N_19928);
nand UO_1152 (O_1152,N_19865,N_19624);
or UO_1153 (O_1153,N_19660,N_19899);
nand UO_1154 (O_1154,N_19647,N_19966);
nand UO_1155 (O_1155,N_19942,N_19845);
or UO_1156 (O_1156,N_19699,N_19643);
and UO_1157 (O_1157,N_19728,N_19744);
and UO_1158 (O_1158,N_19944,N_19845);
nor UO_1159 (O_1159,N_19965,N_19633);
or UO_1160 (O_1160,N_19933,N_19929);
nand UO_1161 (O_1161,N_19890,N_19976);
nor UO_1162 (O_1162,N_19964,N_19888);
nor UO_1163 (O_1163,N_19620,N_19657);
nor UO_1164 (O_1164,N_19985,N_19899);
nand UO_1165 (O_1165,N_19707,N_19761);
nor UO_1166 (O_1166,N_19912,N_19650);
nand UO_1167 (O_1167,N_19723,N_19828);
nand UO_1168 (O_1168,N_19664,N_19751);
nor UO_1169 (O_1169,N_19924,N_19848);
and UO_1170 (O_1170,N_19937,N_19752);
nor UO_1171 (O_1171,N_19758,N_19888);
or UO_1172 (O_1172,N_19808,N_19756);
and UO_1173 (O_1173,N_19647,N_19936);
nor UO_1174 (O_1174,N_19636,N_19796);
and UO_1175 (O_1175,N_19974,N_19621);
nor UO_1176 (O_1176,N_19688,N_19823);
nor UO_1177 (O_1177,N_19981,N_19750);
and UO_1178 (O_1178,N_19805,N_19976);
or UO_1179 (O_1179,N_19855,N_19997);
and UO_1180 (O_1180,N_19941,N_19992);
nor UO_1181 (O_1181,N_19957,N_19695);
nand UO_1182 (O_1182,N_19608,N_19881);
nand UO_1183 (O_1183,N_19817,N_19655);
and UO_1184 (O_1184,N_19847,N_19744);
or UO_1185 (O_1185,N_19993,N_19871);
nor UO_1186 (O_1186,N_19813,N_19895);
nor UO_1187 (O_1187,N_19853,N_19852);
and UO_1188 (O_1188,N_19952,N_19740);
and UO_1189 (O_1189,N_19803,N_19771);
and UO_1190 (O_1190,N_19630,N_19995);
nand UO_1191 (O_1191,N_19966,N_19650);
nor UO_1192 (O_1192,N_19793,N_19772);
nor UO_1193 (O_1193,N_19634,N_19821);
nor UO_1194 (O_1194,N_19895,N_19770);
and UO_1195 (O_1195,N_19620,N_19956);
nor UO_1196 (O_1196,N_19655,N_19664);
and UO_1197 (O_1197,N_19974,N_19869);
nor UO_1198 (O_1198,N_19753,N_19945);
nand UO_1199 (O_1199,N_19633,N_19913);
nor UO_1200 (O_1200,N_19937,N_19740);
or UO_1201 (O_1201,N_19860,N_19954);
nor UO_1202 (O_1202,N_19994,N_19613);
and UO_1203 (O_1203,N_19922,N_19783);
or UO_1204 (O_1204,N_19689,N_19601);
and UO_1205 (O_1205,N_19841,N_19722);
nor UO_1206 (O_1206,N_19986,N_19911);
or UO_1207 (O_1207,N_19730,N_19834);
and UO_1208 (O_1208,N_19939,N_19707);
and UO_1209 (O_1209,N_19733,N_19639);
and UO_1210 (O_1210,N_19736,N_19601);
and UO_1211 (O_1211,N_19649,N_19753);
nor UO_1212 (O_1212,N_19710,N_19605);
nor UO_1213 (O_1213,N_19875,N_19933);
nor UO_1214 (O_1214,N_19626,N_19604);
nor UO_1215 (O_1215,N_19870,N_19858);
nor UO_1216 (O_1216,N_19645,N_19995);
nand UO_1217 (O_1217,N_19668,N_19961);
nand UO_1218 (O_1218,N_19781,N_19795);
nand UO_1219 (O_1219,N_19972,N_19963);
and UO_1220 (O_1220,N_19859,N_19774);
nor UO_1221 (O_1221,N_19685,N_19640);
or UO_1222 (O_1222,N_19809,N_19784);
or UO_1223 (O_1223,N_19801,N_19971);
and UO_1224 (O_1224,N_19794,N_19982);
nand UO_1225 (O_1225,N_19749,N_19624);
or UO_1226 (O_1226,N_19898,N_19900);
or UO_1227 (O_1227,N_19777,N_19830);
nand UO_1228 (O_1228,N_19632,N_19885);
nand UO_1229 (O_1229,N_19635,N_19802);
nor UO_1230 (O_1230,N_19831,N_19930);
nand UO_1231 (O_1231,N_19673,N_19828);
and UO_1232 (O_1232,N_19866,N_19999);
nor UO_1233 (O_1233,N_19946,N_19765);
nand UO_1234 (O_1234,N_19648,N_19974);
nor UO_1235 (O_1235,N_19767,N_19921);
and UO_1236 (O_1236,N_19814,N_19816);
nor UO_1237 (O_1237,N_19887,N_19900);
and UO_1238 (O_1238,N_19632,N_19802);
xnor UO_1239 (O_1239,N_19686,N_19795);
and UO_1240 (O_1240,N_19739,N_19735);
and UO_1241 (O_1241,N_19866,N_19650);
nor UO_1242 (O_1242,N_19791,N_19728);
or UO_1243 (O_1243,N_19838,N_19627);
and UO_1244 (O_1244,N_19953,N_19756);
nor UO_1245 (O_1245,N_19669,N_19626);
or UO_1246 (O_1246,N_19948,N_19985);
nand UO_1247 (O_1247,N_19819,N_19727);
and UO_1248 (O_1248,N_19953,N_19860);
or UO_1249 (O_1249,N_19615,N_19965);
nor UO_1250 (O_1250,N_19723,N_19713);
nor UO_1251 (O_1251,N_19602,N_19651);
nand UO_1252 (O_1252,N_19838,N_19927);
or UO_1253 (O_1253,N_19727,N_19768);
or UO_1254 (O_1254,N_19714,N_19690);
nand UO_1255 (O_1255,N_19602,N_19816);
or UO_1256 (O_1256,N_19808,N_19836);
or UO_1257 (O_1257,N_19722,N_19844);
nand UO_1258 (O_1258,N_19815,N_19893);
nor UO_1259 (O_1259,N_19778,N_19852);
or UO_1260 (O_1260,N_19971,N_19745);
nand UO_1261 (O_1261,N_19713,N_19658);
nand UO_1262 (O_1262,N_19954,N_19899);
nor UO_1263 (O_1263,N_19809,N_19797);
nor UO_1264 (O_1264,N_19779,N_19935);
and UO_1265 (O_1265,N_19682,N_19653);
and UO_1266 (O_1266,N_19743,N_19650);
nor UO_1267 (O_1267,N_19601,N_19919);
or UO_1268 (O_1268,N_19691,N_19673);
or UO_1269 (O_1269,N_19862,N_19964);
nor UO_1270 (O_1270,N_19869,N_19669);
or UO_1271 (O_1271,N_19777,N_19854);
nor UO_1272 (O_1272,N_19919,N_19857);
nand UO_1273 (O_1273,N_19725,N_19645);
nor UO_1274 (O_1274,N_19910,N_19941);
nor UO_1275 (O_1275,N_19715,N_19702);
and UO_1276 (O_1276,N_19976,N_19915);
nand UO_1277 (O_1277,N_19744,N_19832);
and UO_1278 (O_1278,N_19833,N_19941);
or UO_1279 (O_1279,N_19638,N_19711);
or UO_1280 (O_1280,N_19917,N_19749);
nor UO_1281 (O_1281,N_19653,N_19930);
or UO_1282 (O_1282,N_19907,N_19611);
nand UO_1283 (O_1283,N_19676,N_19712);
or UO_1284 (O_1284,N_19638,N_19630);
nor UO_1285 (O_1285,N_19812,N_19833);
or UO_1286 (O_1286,N_19842,N_19639);
and UO_1287 (O_1287,N_19614,N_19887);
nand UO_1288 (O_1288,N_19695,N_19933);
and UO_1289 (O_1289,N_19862,N_19770);
nand UO_1290 (O_1290,N_19678,N_19878);
and UO_1291 (O_1291,N_19774,N_19972);
nand UO_1292 (O_1292,N_19882,N_19601);
nand UO_1293 (O_1293,N_19659,N_19701);
nor UO_1294 (O_1294,N_19680,N_19657);
and UO_1295 (O_1295,N_19652,N_19639);
nor UO_1296 (O_1296,N_19977,N_19720);
nand UO_1297 (O_1297,N_19672,N_19698);
nand UO_1298 (O_1298,N_19918,N_19841);
or UO_1299 (O_1299,N_19614,N_19715);
or UO_1300 (O_1300,N_19907,N_19746);
nand UO_1301 (O_1301,N_19608,N_19965);
and UO_1302 (O_1302,N_19968,N_19830);
or UO_1303 (O_1303,N_19888,N_19605);
nand UO_1304 (O_1304,N_19808,N_19899);
and UO_1305 (O_1305,N_19671,N_19958);
or UO_1306 (O_1306,N_19997,N_19888);
nor UO_1307 (O_1307,N_19604,N_19702);
and UO_1308 (O_1308,N_19875,N_19634);
nor UO_1309 (O_1309,N_19817,N_19918);
or UO_1310 (O_1310,N_19669,N_19709);
and UO_1311 (O_1311,N_19899,N_19753);
or UO_1312 (O_1312,N_19963,N_19712);
and UO_1313 (O_1313,N_19967,N_19618);
nor UO_1314 (O_1314,N_19902,N_19658);
nand UO_1315 (O_1315,N_19652,N_19901);
nand UO_1316 (O_1316,N_19873,N_19703);
nor UO_1317 (O_1317,N_19659,N_19825);
and UO_1318 (O_1318,N_19680,N_19864);
or UO_1319 (O_1319,N_19862,N_19744);
or UO_1320 (O_1320,N_19745,N_19866);
nand UO_1321 (O_1321,N_19925,N_19637);
nor UO_1322 (O_1322,N_19670,N_19943);
or UO_1323 (O_1323,N_19695,N_19868);
xnor UO_1324 (O_1324,N_19685,N_19864);
or UO_1325 (O_1325,N_19660,N_19920);
and UO_1326 (O_1326,N_19820,N_19968);
nand UO_1327 (O_1327,N_19794,N_19712);
and UO_1328 (O_1328,N_19865,N_19828);
or UO_1329 (O_1329,N_19909,N_19665);
nand UO_1330 (O_1330,N_19806,N_19996);
and UO_1331 (O_1331,N_19831,N_19837);
nand UO_1332 (O_1332,N_19935,N_19932);
nor UO_1333 (O_1333,N_19637,N_19943);
nor UO_1334 (O_1334,N_19797,N_19712);
and UO_1335 (O_1335,N_19940,N_19908);
nor UO_1336 (O_1336,N_19905,N_19802);
nor UO_1337 (O_1337,N_19662,N_19806);
nor UO_1338 (O_1338,N_19690,N_19768);
nand UO_1339 (O_1339,N_19696,N_19691);
xnor UO_1340 (O_1340,N_19825,N_19746);
nand UO_1341 (O_1341,N_19954,N_19673);
and UO_1342 (O_1342,N_19813,N_19875);
nand UO_1343 (O_1343,N_19603,N_19797);
and UO_1344 (O_1344,N_19954,N_19605);
or UO_1345 (O_1345,N_19821,N_19955);
nor UO_1346 (O_1346,N_19658,N_19617);
nand UO_1347 (O_1347,N_19752,N_19682);
or UO_1348 (O_1348,N_19610,N_19978);
and UO_1349 (O_1349,N_19938,N_19851);
or UO_1350 (O_1350,N_19682,N_19787);
xnor UO_1351 (O_1351,N_19791,N_19636);
nand UO_1352 (O_1352,N_19828,N_19888);
nand UO_1353 (O_1353,N_19776,N_19971);
or UO_1354 (O_1354,N_19604,N_19619);
or UO_1355 (O_1355,N_19918,N_19649);
and UO_1356 (O_1356,N_19751,N_19673);
nor UO_1357 (O_1357,N_19800,N_19679);
or UO_1358 (O_1358,N_19968,N_19847);
nand UO_1359 (O_1359,N_19858,N_19820);
nor UO_1360 (O_1360,N_19748,N_19689);
nor UO_1361 (O_1361,N_19819,N_19957);
nor UO_1362 (O_1362,N_19678,N_19793);
or UO_1363 (O_1363,N_19726,N_19814);
nor UO_1364 (O_1364,N_19989,N_19862);
and UO_1365 (O_1365,N_19898,N_19635);
nand UO_1366 (O_1366,N_19689,N_19910);
or UO_1367 (O_1367,N_19830,N_19877);
and UO_1368 (O_1368,N_19999,N_19600);
nor UO_1369 (O_1369,N_19843,N_19971);
nand UO_1370 (O_1370,N_19760,N_19961);
or UO_1371 (O_1371,N_19975,N_19823);
nor UO_1372 (O_1372,N_19828,N_19976);
and UO_1373 (O_1373,N_19743,N_19826);
or UO_1374 (O_1374,N_19990,N_19605);
nand UO_1375 (O_1375,N_19826,N_19796);
nand UO_1376 (O_1376,N_19732,N_19629);
and UO_1377 (O_1377,N_19755,N_19904);
or UO_1378 (O_1378,N_19891,N_19682);
nor UO_1379 (O_1379,N_19730,N_19798);
nor UO_1380 (O_1380,N_19832,N_19692);
and UO_1381 (O_1381,N_19718,N_19679);
nor UO_1382 (O_1382,N_19873,N_19853);
or UO_1383 (O_1383,N_19614,N_19895);
nor UO_1384 (O_1384,N_19871,N_19986);
or UO_1385 (O_1385,N_19802,N_19775);
nor UO_1386 (O_1386,N_19669,N_19852);
nand UO_1387 (O_1387,N_19688,N_19657);
and UO_1388 (O_1388,N_19862,N_19868);
or UO_1389 (O_1389,N_19888,N_19759);
nand UO_1390 (O_1390,N_19885,N_19933);
and UO_1391 (O_1391,N_19725,N_19784);
or UO_1392 (O_1392,N_19885,N_19710);
and UO_1393 (O_1393,N_19874,N_19823);
nand UO_1394 (O_1394,N_19967,N_19907);
and UO_1395 (O_1395,N_19687,N_19928);
nor UO_1396 (O_1396,N_19952,N_19817);
and UO_1397 (O_1397,N_19730,N_19884);
or UO_1398 (O_1398,N_19833,N_19954);
and UO_1399 (O_1399,N_19645,N_19677);
and UO_1400 (O_1400,N_19789,N_19737);
nand UO_1401 (O_1401,N_19974,N_19752);
and UO_1402 (O_1402,N_19628,N_19852);
nor UO_1403 (O_1403,N_19957,N_19888);
nand UO_1404 (O_1404,N_19708,N_19613);
or UO_1405 (O_1405,N_19614,N_19767);
and UO_1406 (O_1406,N_19646,N_19868);
or UO_1407 (O_1407,N_19652,N_19834);
and UO_1408 (O_1408,N_19908,N_19866);
or UO_1409 (O_1409,N_19740,N_19975);
and UO_1410 (O_1410,N_19978,N_19946);
or UO_1411 (O_1411,N_19944,N_19633);
nand UO_1412 (O_1412,N_19931,N_19670);
and UO_1413 (O_1413,N_19681,N_19657);
and UO_1414 (O_1414,N_19818,N_19650);
or UO_1415 (O_1415,N_19684,N_19949);
nand UO_1416 (O_1416,N_19736,N_19742);
nand UO_1417 (O_1417,N_19675,N_19750);
nand UO_1418 (O_1418,N_19878,N_19917);
nand UO_1419 (O_1419,N_19711,N_19840);
or UO_1420 (O_1420,N_19973,N_19766);
and UO_1421 (O_1421,N_19863,N_19996);
nand UO_1422 (O_1422,N_19777,N_19786);
or UO_1423 (O_1423,N_19700,N_19911);
nor UO_1424 (O_1424,N_19864,N_19742);
or UO_1425 (O_1425,N_19849,N_19908);
nand UO_1426 (O_1426,N_19893,N_19631);
nor UO_1427 (O_1427,N_19832,N_19821);
or UO_1428 (O_1428,N_19759,N_19909);
nor UO_1429 (O_1429,N_19750,N_19621);
and UO_1430 (O_1430,N_19719,N_19953);
nand UO_1431 (O_1431,N_19802,N_19768);
or UO_1432 (O_1432,N_19873,N_19608);
or UO_1433 (O_1433,N_19792,N_19903);
and UO_1434 (O_1434,N_19676,N_19985);
or UO_1435 (O_1435,N_19635,N_19822);
nand UO_1436 (O_1436,N_19708,N_19784);
nand UO_1437 (O_1437,N_19898,N_19787);
nand UO_1438 (O_1438,N_19877,N_19754);
nor UO_1439 (O_1439,N_19972,N_19874);
nor UO_1440 (O_1440,N_19696,N_19690);
nand UO_1441 (O_1441,N_19948,N_19667);
nor UO_1442 (O_1442,N_19904,N_19794);
or UO_1443 (O_1443,N_19925,N_19626);
and UO_1444 (O_1444,N_19787,N_19981);
nand UO_1445 (O_1445,N_19864,N_19937);
and UO_1446 (O_1446,N_19826,N_19926);
nor UO_1447 (O_1447,N_19701,N_19767);
nand UO_1448 (O_1448,N_19869,N_19993);
nor UO_1449 (O_1449,N_19994,N_19804);
nor UO_1450 (O_1450,N_19655,N_19719);
nor UO_1451 (O_1451,N_19769,N_19727);
xnor UO_1452 (O_1452,N_19952,N_19990);
and UO_1453 (O_1453,N_19898,N_19836);
nor UO_1454 (O_1454,N_19992,N_19949);
and UO_1455 (O_1455,N_19930,N_19702);
or UO_1456 (O_1456,N_19771,N_19889);
nand UO_1457 (O_1457,N_19620,N_19786);
nor UO_1458 (O_1458,N_19840,N_19774);
nand UO_1459 (O_1459,N_19777,N_19789);
nor UO_1460 (O_1460,N_19709,N_19605);
and UO_1461 (O_1461,N_19873,N_19946);
or UO_1462 (O_1462,N_19902,N_19671);
or UO_1463 (O_1463,N_19763,N_19670);
or UO_1464 (O_1464,N_19938,N_19864);
nand UO_1465 (O_1465,N_19748,N_19736);
or UO_1466 (O_1466,N_19815,N_19632);
nor UO_1467 (O_1467,N_19835,N_19836);
and UO_1468 (O_1468,N_19629,N_19844);
nor UO_1469 (O_1469,N_19999,N_19945);
or UO_1470 (O_1470,N_19910,N_19932);
nor UO_1471 (O_1471,N_19661,N_19638);
nor UO_1472 (O_1472,N_19712,N_19636);
or UO_1473 (O_1473,N_19912,N_19824);
nor UO_1474 (O_1474,N_19707,N_19637);
nand UO_1475 (O_1475,N_19915,N_19636);
and UO_1476 (O_1476,N_19886,N_19855);
nand UO_1477 (O_1477,N_19677,N_19799);
nand UO_1478 (O_1478,N_19792,N_19876);
nor UO_1479 (O_1479,N_19964,N_19980);
or UO_1480 (O_1480,N_19775,N_19970);
or UO_1481 (O_1481,N_19937,N_19905);
and UO_1482 (O_1482,N_19780,N_19770);
nand UO_1483 (O_1483,N_19897,N_19813);
or UO_1484 (O_1484,N_19994,N_19765);
nor UO_1485 (O_1485,N_19945,N_19904);
or UO_1486 (O_1486,N_19882,N_19660);
and UO_1487 (O_1487,N_19872,N_19694);
nor UO_1488 (O_1488,N_19996,N_19867);
xor UO_1489 (O_1489,N_19997,N_19773);
and UO_1490 (O_1490,N_19996,N_19870);
xor UO_1491 (O_1491,N_19709,N_19688);
nor UO_1492 (O_1492,N_19902,N_19845);
and UO_1493 (O_1493,N_19754,N_19731);
and UO_1494 (O_1494,N_19934,N_19951);
nor UO_1495 (O_1495,N_19844,N_19994);
and UO_1496 (O_1496,N_19915,N_19754);
nor UO_1497 (O_1497,N_19787,N_19937);
nor UO_1498 (O_1498,N_19630,N_19695);
xor UO_1499 (O_1499,N_19778,N_19676);
nand UO_1500 (O_1500,N_19639,N_19772);
nand UO_1501 (O_1501,N_19771,N_19930);
nor UO_1502 (O_1502,N_19620,N_19706);
nand UO_1503 (O_1503,N_19788,N_19751);
and UO_1504 (O_1504,N_19641,N_19613);
nand UO_1505 (O_1505,N_19703,N_19637);
nand UO_1506 (O_1506,N_19938,N_19892);
or UO_1507 (O_1507,N_19767,N_19758);
and UO_1508 (O_1508,N_19745,N_19817);
and UO_1509 (O_1509,N_19831,N_19730);
and UO_1510 (O_1510,N_19894,N_19909);
nor UO_1511 (O_1511,N_19820,N_19650);
and UO_1512 (O_1512,N_19936,N_19977);
nand UO_1513 (O_1513,N_19813,N_19724);
xor UO_1514 (O_1514,N_19605,N_19800);
or UO_1515 (O_1515,N_19656,N_19695);
or UO_1516 (O_1516,N_19611,N_19917);
nand UO_1517 (O_1517,N_19674,N_19924);
nand UO_1518 (O_1518,N_19881,N_19696);
or UO_1519 (O_1519,N_19707,N_19616);
or UO_1520 (O_1520,N_19921,N_19610);
and UO_1521 (O_1521,N_19800,N_19812);
or UO_1522 (O_1522,N_19825,N_19662);
nor UO_1523 (O_1523,N_19850,N_19941);
nor UO_1524 (O_1524,N_19951,N_19725);
nand UO_1525 (O_1525,N_19703,N_19670);
nor UO_1526 (O_1526,N_19893,N_19904);
nor UO_1527 (O_1527,N_19671,N_19950);
or UO_1528 (O_1528,N_19944,N_19744);
and UO_1529 (O_1529,N_19847,N_19699);
or UO_1530 (O_1530,N_19719,N_19689);
and UO_1531 (O_1531,N_19648,N_19897);
and UO_1532 (O_1532,N_19771,N_19761);
nor UO_1533 (O_1533,N_19891,N_19729);
nor UO_1534 (O_1534,N_19859,N_19784);
or UO_1535 (O_1535,N_19771,N_19915);
and UO_1536 (O_1536,N_19832,N_19823);
and UO_1537 (O_1537,N_19972,N_19935);
or UO_1538 (O_1538,N_19730,N_19913);
or UO_1539 (O_1539,N_19601,N_19804);
and UO_1540 (O_1540,N_19967,N_19649);
nand UO_1541 (O_1541,N_19748,N_19667);
and UO_1542 (O_1542,N_19740,N_19687);
or UO_1543 (O_1543,N_19876,N_19977);
nor UO_1544 (O_1544,N_19718,N_19995);
nor UO_1545 (O_1545,N_19673,N_19767);
and UO_1546 (O_1546,N_19854,N_19913);
and UO_1547 (O_1547,N_19950,N_19905);
nor UO_1548 (O_1548,N_19857,N_19807);
and UO_1549 (O_1549,N_19688,N_19763);
nand UO_1550 (O_1550,N_19851,N_19844);
or UO_1551 (O_1551,N_19948,N_19706);
nand UO_1552 (O_1552,N_19943,N_19851);
nor UO_1553 (O_1553,N_19902,N_19903);
or UO_1554 (O_1554,N_19791,N_19965);
nor UO_1555 (O_1555,N_19735,N_19649);
and UO_1556 (O_1556,N_19714,N_19733);
or UO_1557 (O_1557,N_19872,N_19882);
nand UO_1558 (O_1558,N_19662,N_19856);
nand UO_1559 (O_1559,N_19949,N_19716);
nand UO_1560 (O_1560,N_19929,N_19706);
or UO_1561 (O_1561,N_19821,N_19887);
or UO_1562 (O_1562,N_19654,N_19801);
nand UO_1563 (O_1563,N_19735,N_19763);
and UO_1564 (O_1564,N_19818,N_19876);
xnor UO_1565 (O_1565,N_19691,N_19922);
xor UO_1566 (O_1566,N_19736,N_19690);
nor UO_1567 (O_1567,N_19830,N_19978);
and UO_1568 (O_1568,N_19614,N_19679);
and UO_1569 (O_1569,N_19627,N_19968);
or UO_1570 (O_1570,N_19915,N_19861);
nand UO_1571 (O_1571,N_19742,N_19689);
and UO_1572 (O_1572,N_19704,N_19941);
and UO_1573 (O_1573,N_19657,N_19612);
nor UO_1574 (O_1574,N_19979,N_19760);
nand UO_1575 (O_1575,N_19785,N_19890);
and UO_1576 (O_1576,N_19704,N_19722);
or UO_1577 (O_1577,N_19738,N_19862);
nand UO_1578 (O_1578,N_19812,N_19950);
nand UO_1579 (O_1579,N_19769,N_19873);
and UO_1580 (O_1580,N_19622,N_19702);
nor UO_1581 (O_1581,N_19718,N_19801);
nand UO_1582 (O_1582,N_19940,N_19781);
and UO_1583 (O_1583,N_19938,N_19738);
nor UO_1584 (O_1584,N_19735,N_19729);
or UO_1585 (O_1585,N_19732,N_19661);
nor UO_1586 (O_1586,N_19842,N_19976);
and UO_1587 (O_1587,N_19782,N_19732);
xor UO_1588 (O_1588,N_19757,N_19822);
nand UO_1589 (O_1589,N_19812,N_19798);
nand UO_1590 (O_1590,N_19870,N_19993);
and UO_1591 (O_1591,N_19607,N_19871);
nor UO_1592 (O_1592,N_19722,N_19919);
or UO_1593 (O_1593,N_19987,N_19888);
nor UO_1594 (O_1594,N_19925,N_19889);
or UO_1595 (O_1595,N_19812,N_19656);
nor UO_1596 (O_1596,N_19645,N_19945);
nor UO_1597 (O_1597,N_19774,N_19991);
nor UO_1598 (O_1598,N_19894,N_19915);
nor UO_1599 (O_1599,N_19986,N_19778);
or UO_1600 (O_1600,N_19831,N_19720);
or UO_1601 (O_1601,N_19897,N_19703);
and UO_1602 (O_1602,N_19777,N_19732);
or UO_1603 (O_1603,N_19887,N_19613);
nand UO_1604 (O_1604,N_19944,N_19879);
and UO_1605 (O_1605,N_19878,N_19944);
nand UO_1606 (O_1606,N_19698,N_19851);
nand UO_1607 (O_1607,N_19925,N_19920);
nand UO_1608 (O_1608,N_19794,N_19899);
and UO_1609 (O_1609,N_19948,N_19962);
nand UO_1610 (O_1610,N_19964,N_19757);
nand UO_1611 (O_1611,N_19931,N_19774);
nor UO_1612 (O_1612,N_19932,N_19921);
nor UO_1613 (O_1613,N_19625,N_19631);
nor UO_1614 (O_1614,N_19734,N_19705);
nor UO_1615 (O_1615,N_19690,N_19637);
nor UO_1616 (O_1616,N_19914,N_19620);
nand UO_1617 (O_1617,N_19993,N_19773);
nand UO_1618 (O_1618,N_19733,N_19718);
and UO_1619 (O_1619,N_19834,N_19944);
and UO_1620 (O_1620,N_19737,N_19832);
nor UO_1621 (O_1621,N_19693,N_19769);
or UO_1622 (O_1622,N_19907,N_19848);
and UO_1623 (O_1623,N_19875,N_19776);
nand UO_1624 (O_1624,N_19920,N_19724);
nand UO_1625 (O_1625,N_19927,N_19795);
nand UO_1626 (O_1626,N_19840,N_19869);
nand UO_1627 (O_1627,N_19776,N_19766);
nand UO_1628 (O_1628,N_19867,N_19838);
nor UO_1629 (O_1629,N_19930,N_19609);
nor UO_1630 (O_1630,N_19707,N_19746);
nor UO_1631 (O_1631,N_19822,N_19717);
or UO_1632 (O_1632,N_19636,N_19708);
or UO_1633 (O_1633,N_19794,N_19829);
nor UO_1634 (O_1634,N_19999,N_19932);
nor UO_1635 (O_1635,N_19871,N_19943);
nand UO_1636 (O_1636,N_19611,N_19971);
nor UO_1637 (O_1637,N_19935,N_19730);
nand UO_1638 (O_1638,N_19675,N_19640);
and UO_1639 (O_1639,N_19799,N_19990);
nor UO_1640 (O_1640,N_19607,N_19673);
nor UO_1641 (O_1641,N_19874,N_19856);
and UO_1642 (O_1642,N_19920,N_19805);
and UO_1643 (O_1643,N_19821,N_19653);
and UO_1644 (O_1644,N_19689,N_19871);
nor UO_1645 (O_1645,N_19986,N_19645);
and UO_1646 (O_1646,N_19909,N_19613);
nand UO_1647 (O_1647,N_19678,N_19721);
nor UO_1648 (O_1648,N_19820,N_19659);
nor UO_1649 (O_1649,N_19730,N_19648);
and UO_1650 (O_1650,N_19706,N_19667);
or UO_1651 (O_1651,N_19688,N_19674);
or UO_1652 (O_1652,N_19728,N_19890);
and UO_1653 (O_1653,N_19672,N_19601);
nor UO_1654 (O_1654,N_19755,N_19875);
and UO_1655 (O_1655,N_19812,N_19635);
nand UO_1656 (O_1656,N_19824,N_19770);
or UO_1657 (O_1657,N_19907,N_19663);
nor UO_1658 (O_1658,N_19981,N_19903);
nor UO_1659 (O_1659,N_19825,N_19912);
or UO_1660 (O_1660,N_19952,N_19865);
and UO_1661 (O_1661,N_19974,N_19645);
or UO_1662 (O_1662,N_19940,N_19907);
nand UO_1663 (O_1663,N_19795,N_19850);
nor UO_1664 (O_1664,N_19659,N_19796);
nand UO_1665 (O_1665,N_19688,N_19883);
nand UO_1666 (O_1666,N_19660,N_19996);
nor UO_1667 (O_1667,N_19785,N_19779);
or UO_1668 (O_1668,N_19847,N_19797);
nor UO_1669 (O_1669,N_19867,N_19835);
nand UO_1670 (O_1670,N_19694,N_19720);
nor UO_1671 (O_1671,N_19801,N_19852);
xor UO_1672 (O_1672,N_19609,N_19657);
or UO_1673 (O_1673,N_19737,N_19669);
or UO_1674 (O_1674,N_19902,N_19677);
nor UO_1675 (O_1675,N_19890,N_19880);
nand UO_1676 (O_1676,N_19791,N_19886);
and UO_1677 (O_1677,N_19936,N_19779);
and UO_1678 (O_1678,N_19747,N_19738);
nand UO_1679 (O_1679,N_19991,N_19923);
or UO_1680 (O_1680,N_19693,N_19948);
nor UO_1681 (O_1681,N_19646,N_19629);
or UO_1682 (O_1682,N_19696,N_19870);
and UO_1683 (O_1683,N_19764,N_19808);
nand UO_1684 (O_1684,N_19878,N_19733);
and UO_1685 (O_1685,N_19923,N_19984);
xnor UO_1686 (O_1686,N_19735,N_19761);
and UO_1687 (O_1687,N_19917,N_19814);
nand UO_1688 (O_1688,N_19951,N_19615);
and UO_1689 (O_1689,N_19627,N_19901);
nand UO_1690 (O_1690,N_19846,N_19748);
or UO_1691 (O_1691,N_19691,N_19630);
and UO_1692 (O_1692,N_19663,N_19937);
nor UO_1693 (O_1693,N_19656,N_19623);
or UO_1694 (O_1694,N_19894,N_19819);
or UO_1695 (O_1695,N_19726,N_19765);
and UO_1696 (O_1696,N_19921,N_19780);
nand UO_1697 (O_1697,N_19767,N_19611);
and UO_1698 (O_1698,N_19809,N_19712);
or UO_1699 (O_1699,N_19699,N_19700);
nor UO_1700 (O_1700,N_19755,N_19783);
nand UO_1701 (O_1701,N_19659,N_19699);
nand UO_1702 (O_1702,N_19966,N_19883);
nor UO_1703 (O_1703,N_19789,N_19832);
and UO_1704 (O_1704,N_19699,N_19786);
nand UO_1705 (O_1705,N_19860,N_19760);
nand UO_1706 (O_1706,N_19643,N_19967);
and UO_1707 (O_1707,N_19948,N_19772);
nand UO_1708 (O_1708,N_19741,N_19759);
nand UO_1709 (O_1709,N_19929,N_19814);
and UO_1710 (O_1710,N_19858,N_19853);
nand UO_1711 (O_1711,N_19881,N_19980);
nand UO_1712 (O_1712,N_19900,N_19661);
nor UO_1713 (O_1713,N_19686,N_19845);
nor UO_1714 (O_1714,N_19654,N_19986);
or UO_1715 (O_1715,N_19649,N_19623);
nand UO_1716 (O_1716,N_19870,N_19924);
nor UO_1717 (O_1717,N_19898,N_19908);
nor UO_1718 (O_1718,N_19859,N_19733);
nor UO_1719 (O_1719,N_19775,N_19894);
or UO_1720 (O_1720,N_19643,N_19839);
or UO_1721 (O_1721,N_19777,N_19618);
nand UO_1722 (O_1722,N_19820,N_19717);
or UO_1723 (O_1723,N_19620,N_19872);
and UO_1724 (O_1724,N_19624,N_19933);
nand UO_1725 (O_1725,N_19891,N_19985);
nand UO_1726 (O_1726,N_19987,N_19751);
or UO_1727 (O_1727,N_19755,N_19690);
nor UO_1728 (O_1728,N_19720,N_19920);
nand UO_1729 (O_1729,N_19804,N_19814);
nor UO_1730 (O_1730,N_19810,N_19743);
or UO_1731 (O_1731,N_19893,N_19650);
and UO_1732 (O_1732,N_19657,N_19816);
nand UO_1733 (O_1733,N_19878,N_19741);
nand UO_1734 (O_1734,N_19931,N_19954);
and UO_1735 (O_1735,N_19904,N_19714);
nor UO_1736 (O_1736,N_19744,N_19948);
or UO_1737 (O_1737,N_19849,N_19637);
and UO_1738 (O_1738,N_19957,N_19629);
nand UO_1739 (O_1739,N_19797,N_19690);
and UO_1740 (O_1740,N_19741,N_19911);
and UO_1741 (O_1741,N_19965,N_19846);
nor UO_1742 (O_1742,N_19812,N_19717);
and UO_1743 (O_1743,N_19876,N_19835);
nand UO_1744 (O_1744,N_19716,N_19818);
or UO_1745 (O_1745,N_19765,N_19921);
or UO_1746 (O_1746,N_19950,N_19912);
and UO_1747 (O_1747,N_19727,N_19829);
nand UO_1748 (O_1748,N_19812,N_19801);
nor UO_1749 (O_1749,N_19624,N_19827);
and UO_1750 (O_1750,N_19711,N_19668);
or UO_1751 (O_1751,N_19779,N_19860);
or UO_1752 (O_1752,N_19865,N_19683);
nor UO_1753 (O_1753,N_19723,N_19874);
nor UO_1754 (O_1754,N_19947,N_19677);
or UO_1755 (O_1755,N_19761,N_19606);
nand UO_1756 (O_1756,N_19896,N_19946);
and UO_1757 (O_1757,N_19750,N_19669);
and UO_1758 (O_1758,N_19773,N_19765);
nor UO_1759 (O_1759,N_19949,N_19838);
or UO_1760 (O_1760,N_19736,N_19740);
or UO_1761 (O_1761,N_19944,N_19894);
nand UO_1762 (O_1762,N_19654,N_19714);
and UO_1763 (O_1763,N_19659,N_19996);
nor UO_1764 (O_1764,N_19733,N_19937);
or UO_1765 (O_1765,N_19724,N_19951);
xor UO_1766 (O_1766,N_19929,N_19861);
nand UO_1767 (O_1767,N_19816,N_19669);
or UO_1768 (O_1768,N_19951,N_19698);
nor UO_1769 (O_1769,N_19841,N_19873);
xnor UO_1770 (O_1770,N_19972,N_19795);
nand UO_1771 (O_1771,N_19765,N_19798);
and UO_1772 (O_1772,N_19863,N_19762);
and UO_1773 (O_1773,N_19616,N_19686);
and UO_1774 (O_1774,N_19912,N_19840);
nor UO_1775 (O_1775,N_19997,N_19886);
nor UO_1776 (O_1776,N_19800,N_19735);
or UO_1777 (O_1777,N_19659,N_19734);
and UO_1778 (O_1778,N_19710,N_19712);
nor UO_1779 (O_1779,N_19663,N_19904);
nor UO_1780 (O_1780,N_19945,N_19777);
and UO_1781 (O_1781,N_19901,N_19604);
nor UO_1782 (O_1782,N_19933,N_19771);
or UO_1783 (O_1783,N_19663,N_19934);
nor UO_1784 (O_1784,N_19653,N_19968);
nand UO_1785 (O_1785,N_19634,N_19779);
nor UO_1786 (O_1786,N_19925,N_19941);
nor UO_1787 (O_1787,N_19951,N_19712);
and UO_1788 (O_1788,N_19861,N_19760);
nand UO_1789 (O_1789,N_19928,N_19711);
and UO_1790 (O_1790,N_19634,N_19752);
and UO_1791 (O_1791,N_19602,N_19703);
nor UO_1792 (O_1792,N_19831,N_19834);
or UO_1793 (O_1793,N_19755,N_19836);
xnor UO_1794 (O_1794,N_19817,N_19675);
nand UO_1795 (O_1795,N_19606,N_19960);
or UO_1796 (O_1796,N_19720,N_19746);
or UO_1797 (O_1797,N_19850,N_19851);
nand UO_1798 (O_1798,N_19924,N_19887);
nor UO_1799 (O_1799,N_19977,N_19667);
nand UO_1800 (O_1800,N_19826,N_19795);
or UO_1801 (O_1801,N_19784,N_19646);
and UO_1802 (O_1802,N_19657,N_19970);
nand UO_1803 (O_1803,N_19995,N_19848);
or UO_1804 (O_1804,N_19852,N_19813);
and UO_1805 (O_1805,N_19649,N_19904);
or UO_1806 (O_1806,N_19623,N_19994);
nand UO_1807 (O_1807,N_19757,N_19657);
nand UO_1808 (O_1808,N_19911,N_19901);
nor UO_1809 (O_1809,N_19867,N_19738);
nand UO_1810 (O_1810,N_19896,N_19852);
nand UO_1811 (O_1811,N_19861,N_19792);
nand UO_1812 (O_1812,N_19817,N_19760);
and UO_1813 (O_1813,N_19956,N_19648);
nand UO_1814 (O_1814,N_19644,N_19738);
and UO_1815 (O_1815,N_19910,N_19608);
and UO_1816 (O_1816,N_19753,N_19999);
xor UO_1817 (O_1817,N_19895,N_19783);
or UO_1818 (O_1818,N_19731,N_19875);
nand UO_1819 (O_1819,N_19861,N_19784);
or UO_1820 (O_1820,N_19948,N_19750);
nand UO_1821 (O_1821,N_19927,N_19704);
nor UO_1822 (O_1822,N_19656,N_19897);
nand UO_1823 (O_1823,N_19907,N_19675);
and UO_1824 (O_1824,N_19988,N_19723);
or UO_1825 (O_1825,N_19613,N_19720);
or UO_1826 (O_1826,N_19969,N_19868);
and UO_1827 (O_1827,N_19651,N_19739);
or UO_1828 (O_1828,N_19795,N_19830);
and UO_1829 (O_1829,N_19753,N_19615);
and UO_1830 (O_1830,N_19640,N_19887);
xnor UO_1831 (O_1831,N_19938,N_19828);
nand UO_1832 (O_1832,N_19753,N_19908);
or UO_1833 (O_1833,N_19787,N_19969);
and UO_1834 (O_1834,N_19965,N_19760);
or UO_1835 (O_1835,N_19734,N_19724);
or UO_1836 (O_1836,N_19602,N_19921);
and UO_1837 (O_1837,N_19985,N_19611);
and UO_1838 (O_1838,N_19808,N_19708);
nand UO_1839 (O_1839,N_19840,N_19860);
nand UO_1840 (O_1840,N_19967,N_19946);
nand UO_1841 (O_1841,N_19647,N_19613);
nand UO_1842 (O_1842,N_19837,N_19958);
or UO_1843 (O_1843,N_19990,N_19937);
nand UO_1844 (O_1844,N_19984,N_19924);
nand UO_1845 (O_1845,N_19685,N_19706);
and UO_1846 (O_1846,N_19794,N_19998);
and UO_1847 (O_1847,N_19770,N_19826);
nor UO_1848 (O_1848,N_19811,N_19641);
and UO_1849 (O_1849,N_19855,N_19629);
and UO_1850 (O_1850,N_19843,N_19868);
and UO_1851 (O_1851,N_19991,N_19999);
and UO_1852 (O_1852,N_19651,N_19890);
nand UO_1853 (O_1853,N_19736,N_19783);
and UO_1854 (O_1854,N_19997,N_19669);
or UO_1855 (O_1855,N_19860,N_19694);
or UO_1856 (O_1856,N_19635,N_19799);
or UO_1857 (O_1857,N_19746,N_19676);
nor UO_1858 (O_1858,N_19826,N_19858);
nand UO_1859 (O_1859,N_19730,N_19632);
and UO_1860 (O_1860,N_19896,N_19947);
nor UO_1861 (O_1861,N_19937,N_19961);
nor UO_1862 (O_1862,N_19745,N_19717);
or UO_1863 (O_1863,N_19761,N_19859);
and UO_1864 (O_1864,N_19763,N_19961);
and UO_1865 (O_1865,N_19695,N_19661);
nand UO_1866 (O_1866,N_19611,N_19716);
nor UO_1867 (O_1867,N_19642,N_19858);
nand UO_1868 (O_1868,N_19901,N_19812);
nor UO_1869 (O_1869,N_19993,N_19760);
or UO_1870 (O_1870,N_19613,N_19979);
nand UO_1871 (O_1871,N_19712,N_19635);
nor UO_1872 (O_1872,N_19930,N_19754);
and UO_1873 (O_1873,N_19860,N_19634);
nand UO_1874 (O_1874,N_19910,N_19626);
nand UO_1875 (O_1875,N_19971,N_19797);
or UO_1876 (O_1876,N_19655,N_19633);
or UO_1877 (O_1877,N_19674,N_19827);
nand UO_1878 (O_1878,N_19729,N_19606);
or UO_1879 (O_1879,N_19880,N_19747);
or UO_1880 (O_1880,N_19901,N_19733);
xnor UO_1881 (O_1881,N_19905,N_19709);
and UO_1882 (O_1882,N_19675,N_19844);
or UO_1883 (O_1883,N_19702,N_19886);
nor UO_1884 (O_1884,N_19898,N_19656);
nand UO_1885 (O_1885,N_19749,N_19898);
or UO_1886 (O_1886,N_19975,N_19625);
and UO_1887 (O_1887,N_19976,N_19886);
or UO_1888 (O_1888,N_19823,N_19725);
or UO_1889 (O_1889,N_19776,N_19654);
and UO_1890 (O_1890,N_19983,N_19911);
and UO_1891 (O_1891,N_19743,N_19778);
nor UO_1892 (O_1892,N_19967,N_19966);
or UO_1893 (O_1893,N_19797,N_19786);
or UO_1894 (O_1894,N_19793,N_19648);
and UO_1895 (O_1895,N_19681,N_19812);
nor UO_1896 (O_1896,N_19724,N_19763);
and UO_1897 (O_1897,N_19847,N_19773);
nand UO_1898 (O_1898,N_19786,N_19750);
nor UO_1899 (O_1899,N_19902,N_19855);
or UO_1900 (O_1900,N_19766,N_19845);
or UO_1901 (O_1901,N_19976,N_19756);
or UO_1902 (O_1902,N_19728,N_19988);
and UO_1903 (O_1903,N_19871,N_19779);
nor UO_1904 (O_1904,N_19705,N_19879);
xnor UO_1905 (O_1905,N_19753,N_19978);
or UO_1906 (O_1906,N_19773,N_19750);
nor UO_1907 (O_1907,N_19722,N_19970);
nand UO_1908 (O_1908,N_19632,N_19694);
or UO_1909 (O_1909,N_19877,N_19981);
and UO_1910 (O_1910,N_19890,N_19962);
and UO_1911 (O_1911,N_19721,N_19905);
nor UO_1912 (O_1912,N_19881,N_19994);
and UO_1913 (O_1913,N_19908,N_19809);
nor UO_1914 (O_1914,N_19895,N_19654);
or UO_1915 (O_1915,N_19859,N_19978);
nand UO_1916 (O_1916,N_19701,N_19829);
nor UO_1917 (O_1917,N_19882,N_19639);
nand UO_1918 (O_1918,N_19617,N_19956);
nor UO_1919 (O_1919,N_19744,N_19682);
and UO_1920 (O_1920,N_19739,N_19725);
or UO_1921 (O_1921,N_19606,N_19845);
and UO_1922 (O_1922,N_19860,N_19707);
nand UO_1923 (O_1923,N_19900,N_19937);
nand UO_1924 (O_1924,N_19747,N_19941);
or UO_1925 (O_1925,N_19848,N_19849);
nor UO_1926 (O_1926,N_19961,N_19737);
nor UO_1927 (O_1927,N_19851,N_19867);
nor UO_1928 (O_1928,N_19645,N_19876);
nand UO_1929 (O_1929,N_19903,N_19729);
nor UO_1930 (O_1930,N_19757,N_19827);
nand UO_1931 (O_1931,N_19865,N_19728);
or UO_1932 (O_1932,N_19807,N_19605);
nor UO_1933 (O_1933,N_19890,N_19706);
or UO_1934 (O_1934,N_19619,N_19902);
and UO_1935 (O_1935,N_19693,N_19676);
and UO_1936 (O_1936,N_19750,N_19627);
and UO_1937 (O_1937,N_19618,N_19802);
and UO_1938 (O_1938,N_19953,N_19986);
and UO_1939 (O_1939,N_19946,N_19828);
and UO_1940 (O_1940,N_19759,N_19676);
nor UO_1941 (O_1941,N_19601,N_19832);
and UO_1942 (O_1942,N_19690,N_19841);
nand UO_1943 (O_1943,N_19911,N_19996);
nor UO_1944 (O_1944,N_19975,N_19777);
or UO_1945 (O_1945,N_19795,N_19604);
nand UO_1946 (O_1946,N_19875,N_19856);
nor UO_1947 (O_1947,N_19770,N_19897);
nand UO_1948 (O_1948,N_19994,N_19617);
and UO_1949 (O_1949,N_19996,N_19720);
or UO_1950 (O_1950,N_19876,N_19669);
or UO_1951 (O_1951,N_19890,N_19654);
and UO_1952 (O_1952,N_19705,N_19944);
and UO_1953 (O_1953,N_19687,N_19959);
nand UO_1954 (O_1954,N_19783,N_19905);
and UO_1955 (O_1955,N_19755,N_19697);
and UO_1956 (O_1956,N_19877,N_19827);
nor UO_1957 (O_1957,N_19966,N_19705);
nand UO_1958 (O_1958,N_19814,N_19718);
or UO_1959 (O_1959,N_19683,N_19797);
and UO_1960 (O_1960,N_19735,N_19771);
nor UO_1961 (O_1961,N_19995,N_19988);
and UO_1962 (O_1962,N_19683,N_19853);
or UO_1963 (O_1963,N_19925,N_19736);
nand UO_1964 (O_1964,N_19966,N_19642);
nor UO_1965 (O_1965,N_19931,N_19682);
nor UO_1966 (O_1966,N_19924,N_19747);
or UO_1967 (O_1967,N_19962,N_19645);
or UO_1968 (O_1968,N_19641,N_19653);
nand UO_1969 (O_1969,N_19975,N_19622);
nor UO_1970 (O_1970,N_19797,N_19726);
nand UO_1971 (O_1971,N_19754,N_19714);
and UO_1972 (O_1972,N_19765,N_19655);
nand UO_1973 (O_1973,N_19803,N_19842);
nor UO_1974 (O_1974,N_19848,N_19797);
xnor UO_1975 (O_1975,N_19800,N_19710);
xor UO_1976 (O_1976,N_19908,N_19887);
and UO_1977 (O_1977,N_19906,N_19887);
nor UO_1978 (O_1978,N_19994,N_19751);
and UO_1979 (O_1979,N_19672,N_19908);
or UO_1980 (O_1980,N_19678,N_19645);
or UO_1981 (O_1981,N_19649,N_19644);
or UO_1982 (O_1982,N_19817,N_19883);
nand UO_1983 (O_1983,N_19986,N_19664);
and UO_1984 (O_1984,N_19704,N_19801);
nand UO_1985 (O_1985,N_19896,N_19924);
and UO_1986 (O_1986,N_19926,N_19948);
nor UO_1987 (O_1987,N_19694,N_19912);
nor UO_1988 (O_1988,N_19896,N_19855);
nand UO_1989 (O_1989,N_19934,N_19604);
and UO_1990 (O_1990,N_19718,N_19623);
or UO_1991 (O_1991,N_19759,N_19788);
and UO_1992 (O_1992,N_19662,N_19697);
nand UO_1993 (O_1993,N_19830,N_19653);
or UO_1994 (O_1994,N_19723,N_19969);
nor UO_1995 (O_1995,N_19702,N_19617);
nor UO_1996 (O_1996,N_19824,N_19695);
and UO_1997 (O_1997,N_19657,N_19645);
or UO_1998 (O_1998,N_19952,N_19655);
or UO_1999 (O_1999,N_19891,N_19932);
and UO_2000 (O_2000,N_19660,N_19801);
or UO_2001 (O_2001,N_19740,N_19725);
or UO_2002 (O_2002,N_19669,N_19699);
nand UO_2003 (O_2003,N_19745,N_19916);
nor UO_2004 (O_2004,N_19833,N_19899);
or UO_2005 (O_2005,N_19958,N_19823);
nor UO_2006 (O_2006,N_19706,N_19888);
nor UO_2007 (O_2007,N_19634,N_19719);
or UO_2008 (O_2008,N_19834,N_19777);
nor UO_2009 (O_2009,N_19972,N_19648);
nand UO_2010 (O_2010,N_19954,N_19809);
or UO_2011 (O_2011,N_19712,N_19806);
nor UO_2012 (O_2012,N_19653,N_19897);
nor UO_2013 (O_2013,N_19809,N_19789);
nand UO_2014 (O_2014,N_19778,N_19949);
or UO_2015 (O_2015,N_19939,N_19669);
nor UO_2016 (O_2016,N_19834,N_19600);
or UO_2017 (O_2017,N_19949,N_19708);
nor UO_2018 (O_2018,N_19716,N_19901);
and UO_2019 (O_2019,N_19742,N_19778);
and UO_2020 (O_2020,N_19688,N_19955);
or UO_2021 (O_2021,N_19608,N_19602);
or UO_2022 (O_2022,N_19908,N_19828);
nor UO_2023 (O_2023,N_19851,N_19823);
nor UO_2024 (O_2024,N_19949,N_19846);
nor UO_2025 (O_2025,N_19625,N_19717);
and UO_2026 (O_2026,N_19605,N_19751);
or UO_2027 (O_2027,N_19862,N_19959);
nor UO_2028 (O_2028,N_19812,N_19827);
nand UO_2029 (O_2029,N_19955,N_19616);
and UO_2030 (O_2030,N_19931,N_19949);
or UO_2031 (O_2031,N_19819,N_19788);
or UO_2032 (O_2032,N_19619,N_19891);
and UO_2033 (O_2033,N_19907,N_19609);
nor UO_2034 (O_2034,N_19890,N_19776);
nor UO_2035 (O_2035,N_19826,N_19775);
or UO_2036 (O_2036,N_19883,N_19918);
and UO_2037 (O_2037,N_19605,N_19996);
and UO_2038 (O_2038,N_19698,N_19844);
nor UO_2039 (O_2039,N_19933,N_19808);
and UO_2040 (O_2040,N_19946,N_19635);
nor UO_2041 (O_2041,N_19994,N_19637);
nor UO_2042 (O_2042,N_19619,N_19603);
nor UO_2043 (O_2043,N_19676,N_19925);
nand UO_2044 (O_2044,N_19764,N_19673);
nand UO_2045 (O_2045,N_19962,N_19696);
and UO_2046 (O_2046,N_19603,N_19886);
nand UO_2047 (O_2047,N_19640,N_19912);
nor UO_2048 (O_2048,N_19859,N_19909);
nor UO_2049 (O_2049,N_19955,N_19778);
or UO_2050 (O_2050,N_19652,N_19791);
or UO_2051 (O_2051,N_19911,N_19769);
and UO_2052 (O_2052,N_19884,N_19913);
nor UO_2053 (O_2053,N_19639,N_19859);
or UO_2054 (O_2054,N_19697,N_19829);
nor UO_2055 (O_2055,N_19616,N_19702);
and UO_2056 (O_2056,N_19738,N_19920);
nor UO_2057 (O_2057,N_19600,N_19672);
nor UO_2058 (O_2058,N_19813,N_19909);
or UO_2059 (O_2059,N_19761,N_19807);
nor UO_2060 (O_2060,N_19744,N_19894);
and UO_2061 (O_2061,N_19751,N_19950);
or UO_2062 (O_2062,N_19885,N_19813);
and UO_2063 (O_2063,N_19829,N_19857);
nand UO_2064 (O_2064,N_19848,N_19764);
and UO_2065 (O_2065,N_19729,N_19769);
and UO_2066 (O_2066,N_19946,N_19673);
nand UO_2067 (O_2067,N_19756,N_19978);
or UO_2068 (O_2068,N_19630,N_19948);
and UO_2069 (O_2069,N_19890,N_19638);
or UO_2070 (O_2070,N_19671,N_19894);
nor UO_2071 (O_2071,N_19890,N_19696);
or UO_2072 (O_2072,N_19923,N_19831);
or UO_2073 (O_2073,N_19975,N_19635);
and UO_2074 (O_2074,N_19894,N_19855);
nor UO_2075 (O_2075,N_19719,N_19816);
or UO_2076 (O_2076,N_19999,N_19844);
or UO_2077 (O_2077,N_19811,N_19946);
nor UO_2078 (O_2078,N_19673,N_19982);
and UO_2079 (O_2079,N_19606,N_19986);
and UO_2080 (O_2080,N_19648,N_19929);
or UO_2081 (O_2081,N_19948,N_19651);
xnor UO_2082 (O_2082,N_19656,N_19630);
nor UO_2083 (O_2083,N_19865,N_19758);
or UO_2084 (O_2084,N_19931,N_19918);
or UO_2085 (O_2085,N_19905,N_19760);
nor UO_2086 (O_2086,N_19789,N_19757);
and UO_2087 (O_2087,N_19921,N_19880);
and UO_2088 (O_2088,N_19637,N_19746);
nand UO_2089 (O_2089,N_19650,N_19851);
or UO_2090 (O_2090,N_19605,N_19846);
nor UO_2091 (O_2091,N_19746,N_19967);
or UO_2092 (O_2092,N_19759,N_19934);
nand UO_2093 (O_2093,N_19976,N_19928);
nor UO_2094 (O_2094,N_19731,N_19828);
nor UO_2095 (O_2095,N_19824,N_19730);
or UO_2096 (O_2096,N_19785,N_19790);
nand UO_2097 (O_2097,N_19667,N_19978);
nor UO_2098 (O_2098,N_19697,N_19979);
or UO_2099 (O_2099,N_19616,N_19744);
or UO_2100 (O_2100,N_19870,N_19844);
nand UO_2101 (O_2101,N_19783,N_19913);
and UO_2102 (O_2102,N_19890,N_19974);
and UO_2103 (O_2103,N_19674,N_19716);
nand UO_2104 (O_2104,N_19917,N_19661);
or UO_2105 (O_2105,N_19812,N_19906);
or UO_2106 (O_2106,N_19687,N_19862);
or UO_2107 (O_2107,N_19999,N_19951);
nor UO_2108 (O_2108,N_19832,N_19686);
or UO_2109 (O_2109,N_19605,N_19610);
nand UO_2110 (O_2110,N_19987,N_19840);
nand UO_2111 (O_2111,N_19810,N_19622);
and UO_2112 (O_2112,N_19656,N_19701);
nor UO_2113 (O_2113,N_19926,N_19660);
nor UO_2114 (O_2114,N_19760,N_19924);
nor UO_2115 (O_2115,N_19781,N_19791);
and UO_2116 (O_2116,N_19632,N_19958);
or UO_2117 (O_2117,N_19711,N_19720);
or UO_2118 (O_2118,N_19830,N_19974);
nor UO_2119 (O_2119,N_19683,N_19768);
nand UO_2120 (O_2120,N_19897,N_19782);
nor UO_2121 (O_2121,N_19671,N_19714);
and UO_2122 (O_2122,N_19943,N_19965);
or UO_2123 (O_2123,N_19772,N_19601);
nor UO_2124 (O_2124,N_19702,N_19910);
or UO_2125 (O_2125,N_19944,N_19614);
nor UO_2126 (O_2126,N_19631,N_19737);
and UO_2127 (O_2127,N_19763,N_19866);
or UO_2128 (O_2128,N_19865,N_19707);
nand UO_2129 (O_2129,N_19715,N_19707);
and UO_2130 (O_2130,N_19854,N_19967);
nor UO_2131 (O_2131,N_19962,N_19975);
nor UO_2132 (O_2132,N_19991,N_19617);
nor UO_2133 (O_2133,N_19833,N_19995);
nor UO_2134 (O_2134,N_19963,N_19731);
nor UO_2135 (O_2135,N_19674,N_19659);
and UO_2136 (O_2136,N_19632,N_19738);
nand UO_2137 (O_2137,N_19696,N_19830);
and UO_2138 (O_2138,N_19915,N_19701);
or UO_2139 (O_2139,N_19676,N_19933);
or UO_2140 (O_2140,N_19627,N_19953);
nor UO_2141 (O_2141,N_19865,N_19743);
nand UO_2142 (O_2142,N_19645,N_19911);
nand UO_2143 (O_2143,N_19837,N_19681);
nor UO_2144 (O_2144,N_19928,N_19706);
nor UO_2145 (O_2145,N_19811,N_19966);
or UO_2146 (O_2146,N_19950,N_19683);
and UO_2147 (O_2147,N_19889,N_19693);
and UO_2148 (O_2148,N_19994,N_19600);
and UO_2149 (O_2149,N_19941,N_19958);
nor UO_2150 (O_2150,N_19968,N_19885);
and UO_2151 (O_2151,N_19745,N_19794);
and UO_2152 (O_2152,N_19776,N_19614);
or UO_2153 (O_2153,N_19631,N_19658);
nand UO_2154 (O_2154,N_19895,N_19961);
nor UO_2155 (O_2155,N_19873,N_19667);
and UO_2156 (O_2156,N_19807,N_19924);
nor UO_2157 (O_2157,N_19747,N_19990);
and UO_2158 (O_2158,N_19992,N_19676);
and UO_2159 (O_2159,N_19638,N_19603);
nand UO_2160 (O_2160,N_19794,N_19646);
and UO_2161 (O_2161,N_19794,N_19779);
and UO_2162 (O_2162,N_19812,N_19967);
or UO_2163 (O_2163,N_19660,N_19758);
and UO_2164 (O_2164,N_19753,N_19796);
or UO_2165 (O_2165,N_19818,N_19772);
or UO_2166 (O_2166,N_19602,N_19807);
nand UO_2167 (O_2167,N_19982,N_19818);
or UO_2168 (O_2168,N_19630,N_19848);
xor UO_2169 (O_2169,N_19931,N_19627);
or UO_2170 (O_2170,N_19734,N_19966);
nand UO_2171 (O_2171,N_19997,N_19998);
nor UO_2172 (O_2172,N_19696,N_19663);
nor UO_2173 (O_2173,N_19922,N_19815);
or UO_2174 (O_2174,N_19666,N_19953);
nor UO_2175 (O_2175,N_19627,N_19748);
and UO_2176 (O_2176,N_19856,N_19718);
nor UO_2177 (O_2177,N_19934,N_19674);
nand UO_2178 (O_2178,N_19790,N_19663);
nor UO_2179 (O_2179,N_19632,N_19696);
and UO_2180 (O_2180,N_19953,N_19770);
nand UO_2181 (O_2181,N_19886,N_19714);
nand UO_2182 (O_2182,N_19769,N_19996);
nor UO_2183 (O_2183,N_19805,N_19633);
or UO_2184 (O_2184,N_19807,N_19936);
nand UO_2185 (O_2185,N_19832,N_19763);
and UO_2186 (O_2186,N_19981,N_19947);
and UO_2187 (O_2187,N_19939,N_19744);
or UO_2188 (O_2188,N_19674,N_19900);
or UO_2189 (O_2189,N_19878,N_19729);
xnor UO_2190 (O_2190,N_19996,N_19937);
or UO_2191 (O_2191,N_19690,N_19964);
nand UO_2192 (O_2192,N_19662,N_19730);
nor UO_2193 (O_2193,N_19769,N_19607);
nand UO_2194 (O_2194,N_19614,N_19925);
or UO_2195 (O_2195,N_19663,N_19852);
nor UO_2196 (O_2196,N_19820,N_19807);
and UO_2197 (O_2197,N_19928,N_19626);
or UO_2198 (O_2198,N_19639,N_19742);
nand UO_2199 (O_2199,N_19862,N_19719);
and UO_2200 (O_2200,N_19632,N_19642);
nand UO_2201 (O_2201,N_19905,N_19779);
nand UO_2202 (O_2202,N_19712,N_19787);
or UO_2203 (O_2203,N_19624,N_19633);
nor UO_2204 (O_2204,N_19990,N_19843);
nor UO_2205 (O_2205,N_19807,N_19872);
and UO_2206 (O_2206,N_19648,N_19632);
nand UO_2207 (O_2207,N_19611,N_19730);
nand UO_2208 (O_2208,N_19859,N_19959);
nand UO_2209 (O_2209,N_19729,N_19845);
or UO_2210 (O_2210,N_19979,N_19908);
and UO_2211 (O_2211,N_19851,N_19989);
nand UO_2212 (O_2212,N_19943,N_19689);
and UO_2213 (O_2213,N_19657,N_19753);
nor UO_2214 (O_2214,N_19660,N_19727);
or UO_2215 (O_2215,N_19706,N_19898);
nor UO_2216 (O_2216,N_19774,N_19791);
or UO_2217 (O_2217,N_19760,N_19804);
and UO_2218 (O_2218,N_19945,N_19643);
nor UO_2219 (O_2219,N_19644,N_19678);
and UO_2220 (O_2220,N_19701,N_19934);
nand UO_2221 (O_2221,N_19697,N_19747);
nand UO_2222 (O_2222,N_19616,N_19775);
or UO_2223 (O_2223,N_19676,N_19752);
or UO_2224 (O_2224,N_19904,N_19619);
and UO_2225 (O_2225,N_19947,N_19697);
nand UO_2226 (O_2226,N_19600,N_19785);
nor UO_2227 (O_2227,N_19697,N_19890);
nand UO_2228 (O_2228,N_19790,N_19988);
or UO_2229 (O_2229,N_19923,N_19829);
nand UO_2230 (O_2230,N_19617,N_19683);
and UO_2231 (O_2231,N_19700,N_19804);
nand UO_2232 (O_2232,N_19792,N_19662);
nand UO_2233 (O_2233,N_19782,N_19705);
nand UO_2234 (O_2234,N_19742,N_19691);
nor UO_2235 (O_2235,N_19880,N_19805);
xor UO_2236 (O_2236,N_19803,N_19996);
and UO_2237 (O_2237,N_19889,N_19611);
or UO_2238 (O_2238,N_19607,N_19851);
nor UO_2239 (O_2239,N_19680,N_19973);
nand UO_2240 (O_2240,N_19738,N_19616);
nand UO_2241 (O_2241,N_19742,N_19817);
and UO_2242 (O_2242,N_19970,N_19752);
or UO_2243 (O_2243,N_19773,N_19711);
or UO_2244 (O_2244,N_19875,N_19722);
or UO_2245 (O_2245,N_19638,N_19612);
or UO_2246 (O_2246,N_19686,N_19661);
or UO_2247 (O_2247,N_19716,N_19873);
nor UO_2248 (O_2248,N_19991,N_19733);
nand UO_2249 (O_2249,N_19712,N_19628);
and UO_2250 (O_2250,N_19719,N_19947);
nand UO_2251 (O_2251,N_19758,N_19729);
nor UO_2252 (O_2252,N_19926,N_19603);
nor UO_2253 (O_2253,N_19981,N_19994);
or UO_2254 (O_2254,N_19798,N_19715);
nor UO_2255 (O_2255,N_19677,N_19746);
and UO_2256 (O_2256,N_19970,N_19717);
nor UO_2257 (O_2257,N_19685,N_19804);
xnor UO_2258 (O_2258,N_19990,N_19927);
nand UO_2259 (O_2259,N_19766,N_19816);
and UO_2260 (O_2260,N_19939,N_19860);
and UO_2261 (O_2261,N_19942,N_19772);
nor UO_2262 (O_2262,N_19655,N_19815);
nand UO_2263 (O_2263,N_19762,N_19858);
and UO_2264 (O_2264,N_19956,N_19769);
and UO_2265 (O_2265,N_19974,N_19660);
nand UO_2266 (O_2266,N_19916,N_19908);
nor UO_2267 (O_2267,N_19661,N_19867);
nor UO_2268 (O_2268,N_19950,N_19883);
or UO_2269 (O_2269,N_19634,N_19716);
nand UO_2270 (O_2270,N_19929,N_19870);
nand UO_2271 (O_2271,N_19906,N_19784);
or UO_2272 (O_2272,N_19785,N_19787);
and UO_2273 (O_2273,N_19799,N_19661);
and UO_2274 (O_2274,N_19833,N_19851);
nor UO_2275 (O_2275,N_19850,N_19797);
nor UO_2276 (O_2276,N_19721,N_19717);
or UO_2277 (O_2277,N_19697,N_19999);
nand UO_2278 (O_2278,N_19893,N_19949);
and UO_2279 (O_2279,N_19776,N_19826);
or UO_2280 (O_2280,N_19644,N_19713);
and UO_2281 (O_2281,N_19646,N_19712);
or UO_2282 (O_2282,N_19704,N_19916);
or UO_2283 (O_2283,N_19670,N_19646);
or UO_2284 (O_2284,N_19915,N_19882);
xor UO_2285 (O_2285,N_19677,N_19816);
nor UO_2286 (O_2286,N_19671,N_19722);
and UO_2287 (O_2287,N_19633,N_19993);
nand UO_2288 (O_2288,N_19729,N_19784);
and UO_2289 (O_2289,N_19724,N_19892);
nor UO_2290 (O_2290,N_19682,N_19965);
and UO_2291 (O_2291,N_19789,N_19661);
nand UO_2292 (O_2292,N_19658,N_19705);
or UO_2293 (O_2293,N_19833,N_19707);
and UO_2294 (O_2294,N_19971,N_19623);
or UO_2295 (O_2295,N_19601,N_19735);
nand UO_2296 (O_2296,N_19645,N_19611);
nor UO_2297 (O_2297,N_19854,N_19677);
and UO_2298 (O_2298,N_19790,N_19613);
or UO_2299 (O_2299,N_19910,N_19959);
nand UO_2300 (O_2300,N_19954,N_19836);
or UO_2301 (O_2301,N_19763,N_19652);
nor UO_2302 (O_2302,N_19952,N_19602);
nor UO_2303 (O_2303,N_19729,N_19650);
or UO_2304 (O_2304,N_19643,N_19732);
or UO_2305 (O_2305,N_19910,N_19682);
nand UO_2306 (O_2306,N_19746,N_19711);
nand UO_2307 (O_2307,N_19787,N_19608);
or UO_2308 (O_2308,N_19799,N_19980);
and UO_2309 (O_2309,N_19844,N_19749);
nand UO_2310 (O_2310,N_19873,N_19709);
and UO_2311 (O_2311,N_19916,N_19673);
and UO_2312 (O_2312,N_19669,N_19690);
and UO_2313 (O_2313,N_19647,N_19622);
or UO_2314 (O_2314,N_19937,N_19632);
nor UO_2315 (O_2315,N_19946,N_19858);
nand UO_2316 (O_2316,N_19854,N_19646);
xor UO_2317 (O_2317,N_19651,N_19604);
or UO_2318 (O_2318,N_19970,N_19740);
nor UO_2319 (O_2319,N_19660,N_19929);
or UO_2320 (O_2320,N_19784,N_19825);
nand UO_2321 (O_2321,N_19788,N_19729);
nand UO_2322 (O_2322,N_19943,N_19696);
nand UO_2323 (O_2323,N_19762,N_19894);
nand UO_2324 (O_2324,N_19665,N_19634);
and UO_2325 (O_2325,N_19764,N_19782);
nor UO_2326 (O_2326,N_19786,N_19805);
nor UO_2327 (O_2327,N_19673,N_19984);
nand UO_2328 (O_2328,N_19633,N_19684);
nor UO_2329 (O_2329,N_19842,N_19972);
xnor UO_2330 (O_2330,N_19749,N_19784);
nand UO_2331 (O_2331,N_19957,N_19704);
nand UO_2332 (O_2332,N_19907,N_19935);
and UO_2333 (O_2333,N_19910,N_19606);
and UO_2334 (O_2334,N_19786,N_19865);
and UO_2335 (O_2335,N_19844,N_19706);
nor UO_2336 (O_2336,N_19886,N_19940);
and UO_2337 (O_2337,N_19826,N_19605);
nor UO_2338 (O_2338,N_19810,N_19745);
nand UO_2339 (O_2339,N_19783,N_19692);
nand UO_2340 (O_2340,N_19943,N_19817);
and UO_2341 (O_2341,N_19837,N_19824);
or UO_2342 (O_2342,N_19651,N_19953);
and UO_2343 (O_2343,N_19673,N_19975);
or UO_2344 (O_2344,N_19633,N_19800);
nor UO_2345 (O_2345,N_19811,N_19843);
or UO_2346 (O_2346,N_19946,N_19895);
or UO_2347 (O_2347,N_19794,N_19972);
nand UO_2348 (O_2348,N_19860,N_19851);
nand UO_2349 (O_2349,N_19761,N_19997);
or UO_2350 (O_2350,N_19695,N_19770);
or UO_2351 (O_2351,N_19771,N_19880);
nand UO_2352 (O_2352,N_19903,N_19674);
nand UO_2353 (O_2353,N_19808,N_19912);
nor UO_2354 (O_2354,N_19708,N_19801);
nand UO_2355 (O_2355,N_19897,N_19783);
nand UO_2356 (O_2356,N_19703,N_19829);
nand UO_2357 (O_2357,N_19627,N_19829);
nand UO_2358 (O_2358,N_19934,N_19742);
nor UO_2359 (O_2359,N_19783,N_19763);
and UO_2360 (O_2360,N_19654,N_19698);
nor UO_2361 (O_2361,N_19636,N_19716);
nand UO_2362 (O_2362,N_19631,N_19990);
and UO_2363 (O_2363,N_19611,N_19802);
nor UO_2364 (O_2364,N_19771,N_19607);
nor UO_2365 (O_2365,N_19751,N_19850);
xor UO_2366 (O_2366,N_19978,N_19765);
nor UO_2367 (O_2367,N_19947,N_19785);
nor UO_2368 (O_2368,N_19603,N_19715);
or UO_2369 (O_2369,N_19741,N_19917);
or UO_2370 (O_2370,N_19816,N_19796);
and UO_2371 (O_2371,N_19797,N_19710);
nor UO_2372 (O_2372,N_19797,N_19773);
and UO_2373 (O_2373,N_19651,N_19671);
nor UO_2374 (O_2374,N_19979,N_19913);
or UO_2375 (O_2375,N_19773,N_19893);
and UO_2376 (O_2376,N_19958,N_19623);
or UO_2377 (O_2377,N_19638,N_19832);
or UO_2378 (O_2378,N_19934,N_19614);
or UO_2379 (O_2379,N_19652,N_19940);
or UO_2380 (O_2380,N_19981,N_19873);
and UO_2381 (O_2381,N_19842,N_19965);
nand UO_2382 (O_2382,N_19646,N_19701);
nand UO_2383 (O_2383,N_19995,N_19636);
nor UO_2384 (O_2384,N_19671,N_19761);
nor UO_2385 (O_2385,N_19644,N_19971);
nor UO_2386 (O_2386,N_19809,N_19696);
and UO_2387 (O_2387,N_19771,N_19811);
nor UO_2388 (O_2388,N_19943,N_19995);
nand UO_2389 (O_2389,N_19980,N_19967);
and UO_2390 (O_2390,N_19731,N_19857);
nand UO_2391 (O_2391,N_19912,N_19874);
nand UO_2392 (O_2392,N_19840,N_19960);
nor UO_2393 (O_2393,N_19926,N_19802);
and UO_2394 (O_2394,N_19903,N_19977);
or UO_2395 (O_2395,N_19979,N_19617);
or UO_2396 (O_2396,N_19646,N_19911);
or UO_2397 (O_2397,N_19741,N_19833);
and UO_2398 (O_2398,N_19688,N_19838);
nor UO_2399 (O_2399,N_19722,N_19611);
nor UO_2400 (O_2400,N_19617,N_19857);
and UO_2401 (O_2401,N_19717,N_19954);
or UO_2402 (O_2402,N_19625,N_19732);
nand UO_2403 (O_2403,N_19600,N_19978);
and UO_2404 (O_2404,N_19604,N_19727);
and UO_2405 (O_2405,N_19713,N_19711);
nor UO_2406 (O_2406,N_19912,N_19617);
or UO_2407 (O_2407,N_19968,N_19786);
nor UO_2408 (O_2408,N_19919,N_19906);
nor UO_2409 (O_2409,N_19768,N_19815);
or UO_2410 (O_2410,N_19749,N_19903);
nand UO_2411 (O_2411,N_19759,N_19754);
or UO_2412 (O_2412,N_19984,N_19626);
nand UO_2413 (O_2413,N_19879,N_19722);
nor UO_2414 (O_2414,N_19958,N_19618);
and UO_2415 (O_2415,N_19658,N_19765);
nor UO_2416 (O_2416,N_19864,N_19608);
and UO_2417 (O_2417,N_19981,N_19719);
or UO_2418 (O_2418,N_19625,N_19755);
or UO_2419 (O_2419,N_19809,N_19857);
nand UO_2420 (O_2420,N_19883,N_19932);
and UO_2421 (O_2421,N_19781,N_19774);
nor UO_2422 (O_2422,N_19808,N_19732);
nor UO_2423 (O_2423,N_19779,N_19993);
nor UO_2424 (O_2424,N_19730,N_19664);
and UO_2425 (O_2425,N_19946,N_19824);
nor UO_2426 (O_2426,N_19695,N_19830);
and UO_2427 (O_2427,N_19608,N_19809);
nand UO_2428 (O_2428,N_19898,N_19673);
nor UO_2429 (O_2429,N_19660,N_19908);
nand UO_2430 (O_2430,N_19766,N_19829);
nor UO_2431 (O_2431,N_19939,N_19819);
nor UO_2432 (O_2432,N_19872,N_19686);
nand UO_2433 (O_2433,N_19801,N_19783);
nand UO_2434 (O_2434,N_19689,N_19881);
and UO_2435 (O_2435,N_19898,N_19717);
or UO_2436 (O_2436,N_19916,N_19844);
and UO_2437 (O_2437,N_19903,N_19980);
or UO_2438 (O_2438,N_19734,N_19984);
nand UO_2439 (O_2439,N_19746,N_19895);
and UO_2440 (O_2440,N_19941,N_19649);
nand UO_2441 (O_2441,N_19702,N_19857);
or UO_2442 (O_2442,N_19734,N_19914);
nand UO_2443 (O_2443,N_19798,N_19802);
nand UO_2444 (O_2444,N_19861,N_19701);
nand UO_2445 (O_2445,N_19676,N_19769);
nand UO_2446 (O_2446,N_19816,N_19951);
nand UO_2447 (O_2447,N_19803,N_19626);
and UO_2448 (O_2448,N_19750,N_19638);
or UO_2449 (O_2449,N_19707,N_19863);
nor UO_2450 (O_2450,N_19804,N_19646);
or UO_2451 (O_2451,N_19715,N_19648);
and UO_2452 (O_2452,N_19663,N_19945);
or UO_2453 (O_2453,N_19998,N_19631);
nor UO_2454 (O_2454,N_19827,N_19636);
nand UO_2455 (O_2455,N_19661,N_19884);
and UO_2456 (O_2456,N_19904,N_19661);
nand UO_2457 (O_2457,N_19985,N_19610);
or UO_2458 (O_2458,N_19819,N_19963);
nand UO_2459 (O_2459,N_19793,N_19786);
or UO_2460 (O_2460,N_19933,N_19882);
or UO_2461 (O_2461,N_19967,N_19849);
nand UO_2462 (O_2462,N_19753,N_19814);
nor UO_2463 (O_2463,N_19740,N_19873);
nand UO_2464 (O_2464,N_19986,N_19683);
nor UO_2465 (O_2465,N_19694,N_19909);
nand UO_2466 (O_2466,N_19797,N_19737);
and UO_2467 (O_2467,N_19940,N_19646);
or UO_2468 (O_2468,N_19749,N_19887);
and UO_2469 (O_2469,N_19893,N_19891);
nand UO_2470 (O_2470,N_19737,N_19756);
nand UO_2471 (O_2471,N_19742,N_19745);
or UO_2472 (O_2472,N_19799,N_19744);
or UO_2473 (O_2473,N_19770,N_19967);
nor UO_2474 (O_2474,N_19881,N_19888);
or UO_2475 (O_2475,N_19763,N_19680);
nor UO_2476 (O_2476,N_19744,N_19903);
nand UO_2477 (O_2477,N_19693,N_19805);
nor UO_2478 (O_2478,N_19898,N_19682);
and UO_2479 (O_2479,N_19829,N_19711);
nor UO_2480 (O_2480,N_19725,N_19708);
or UO_2481 (O_2481,N_19840,N_19894);
nand UO_2482 (O_2482,N_19712,N_19992);
and UO_2483 (O_2483,N_19783,N_19936);
and UO_2484 (O_2484,N_19722,N_19926);
nand UO_2485 (O_2485,N_19768,N_19850);
or UO_2486 (O_2486,N_19726,N_19926);
nor UO_2487 (O_2487,N_19665,N_19930);
or UO_2488 (O_2488,N_19779,N_19854);
nor UO_2489 (O_2489,N_19628,N_19691);
nand UO_2490 (O_2490,N_19949,N_19917);
or UO_2491 (O_2491,N_19854,N_19751);
and UO_2492 (O_2492,N_19639,N_19849);
and UO_2493 (O_2493,N_19918,N_19856);
nand UO_2494 (O_2494,N_19851,N_19845);
and UO_2495 (O_2495,N_19604,N_19996);
nor UO_2496 (O_2496,N_19954,N_19947);
or UO_2497 (O_2497,N_19820,N_19943);
or UO_2498 (O_2498,N_19681,N_19782);
or UO_2499 (O_2499,N_19938,N_19744);
endmodule