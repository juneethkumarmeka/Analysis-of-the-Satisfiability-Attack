module basic_1000_10000_1500_10_levels_1xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_449,In_43);
nor U1 (N_1,In_644,In_261);
and U2 (N_2,In_357,In_486);
or U3 (N_3,In_199,In_390);
nand U4 (N_4,In_899,In_334);
or U5 (N_5,In_281,In_673);
nor U6 (N_6,In_597,In_428);
nand U7 (N_7,In_285,In_313);
nor U8 (N_8,In_102,In_595);
or U9 (N_9,In_405,In_493);
nand U10 (N_10,In_373,In_750);
and U11 (N_11,In_648,In_84);
and U12 (N_12,In_946,In_478);
or U13 (N_13,In_156,In_631);
nor U14 (N_14,In_919,In_875);
nor U15 (N_15,In_747,In_839);
nor U16 (N_16,In_621,In_850);
nand U17 (N_17,In_793,In_136);
and U18 (N_18,In_705,In_387);
and U19 (N_19,In_430,In_212);
or U20 (N_20,In_820,In_776);
and U21 (N_21,In_95,In_828);
nand U22 (N_22,In_520,In_368);
and U23 (N_23,In_836,In_221);
or U24 (N_24,In_718,In_929);
nor U25 (N_25,In_286,In_532);
and U26 (N_26,In_344,In_164);
xor U27 (N_27,In_564,In_33);
or U28 (N_28,In_814,In_441);
nand U29 (N_29,In_15,In_259);
xor U30 (N_30,In_667,In_413);
nand U31 (N_31,In_751,In_873);
nor U32 (N_32,In_897,In_533);
and U33 (N_33,In_124,In_603);
nor U34 (N_34,In_420,In_243);
nand U35 (N_35,In_927,In_152);
or U36 (N_36,In_548,In_816);
and U37 (N_37,In_588,In_476);
nor U38 (N_38,In_865,In_176);
and U39 (N_39,In_332,In_193);
nand U40 (N_40,In_426,In_958);
or U41 (N_41,In_3,In_862);
nor U42 (N_42,In_52,In_643);
or U43 (N_43,In_492,In_184);
nand U44 (N_44,In_504,In_0);
nand U45 (N_45,In_687,In_108);
or U46 (N_46,In_146,In_926);
and U47 (N_47,In_216,In_561);
nand U48 (N_48,In_525,In_696);
or U49 (N_49,In_998,In_876);
nor U50 (N_50,In_309,In_479);
and U51 (N_51,In_396,In_801);
and U52 (N_52,In_275,In_560);
nand U53 (N_53,In_681,In_634);
or U54 (N_54,In_397,In_122);
and U55 (N_55,In_767,In_635);
or U56 (N_56,In_765,In_386);
nand U57 (N_57,In_361,In_855);
nor U58 (N_58,In_14,In_534);
and U59 (N_59,In_408,In_203);
and U60 (N_60,In_66,In_996);
or U61 (N_61,In_717,In_779);
and U62 (N_62,In_975,In_999);
and U63 (N_63,In_117,In_672);
nor U64 (N_64,In_42,In_893);
nor U65 (N_65,In_94,In_527);
or U66 (N_66,In_759,In_220);
nand U67 (N_67,In_498,In_213);
nand U68 (N_68,In_686,In_73);
xor U69 (N_69,In_715,In_445);
and U70 (N_70,In_518,In_783);
nand U71 (N_71,In_811,In_650);
and U72 (N_72,In_263,In_264);
or U73 (N_73,In_257,In_412);
and U74 (N_74,In_542,In_448);
or U75 (N_75,In_180,In_74);
and U76 (N_76,In_495,In_83);
nor U77 (N_77,In_436,In_961);
nor U78 (N_78,In_364,In_986);
and U79 (N_79,In_198,In_976);
nand U80 (N_80,In_740,In_699);
or U81 (N_81,In_487,In_802);
and U82 (N_82,In_840,In_21);
nand U83 (N_83,In_771,In_79);
or U84 (N_84,In_982,In_222);
nand U85 (N_85,In_63,In_950);
xnor U86 (N_86,In_292,In_728);
nand U87 (N_87,In_886,In_210);
nor U88 (N_88,In_928,In_111);
nand U89 (N_89,In_228,In_121);
nor U90 (N_90,In_105,In_513);
nand U91 (N_91,In_626,In_166);
or U92 (N_92,In_918,In_295);
or U93 (N_93,In_760,In_677);
and U94 (N_94,In_889,In_107);
or U95 (N_95,In_116,In_719);
nand U96 (N_96,In_558,In_517);
nor U97 (N_97,In_125,In_155);
or U98 (N_98,In_662,In_992);
and U99 (N_99,In_847,In_211);
and U100 (N_100,In_887,In_114);
nand U101 (N_101,In_819,In_985);
or U102 (N_102,In_379,In_591);
nor U103 (N_103,In_885,In_274);
or U104 (N_104,In_674,In_713);
nor U105 (N_105,In_823,In_853);
nor U106 (N_106,In_165,In_741);
nor U107 (N_107,In_419,In_129);
nor U108 (N_108,In_80,In_53);
nand U109 (N_109,In_407,In_777);
nand U110 (N_110,In_25,In_629);
and U111 (N_111,In_39,In_726);
nor U112 (N_112,In_153,In_645);
nor U113 (N_113,In_730,In_916);
and U114 (N_114,In_201,In_47);
nor U115 (N_115,In_872,In_485);
or U116 (N_116,In_908,In_447);
or U117 (N_117,In_797,In_181);
or U118 (N_118,In_133,In_370);
nor U119 (N_119,In_796,In_265);
or U120 (N_120,In_290,In_563);
nor U121 (N_121,In_911,In_651);
and U122 (N_122,In_331,In_774);
or U123 (N_123,In_659,In_362);
or U124 (N_124,In_963,In_308);
or U125 (N_125,In_177,In_112);
nand U126 (N_126,In_45,In_974);
nand U127 (N_127,In_115,In_318);
nand U128 (N_128,In_247,In_914);
nand U129 (N_129,In_197,In_615);
nor U130 (N_130,In_287,In_838);
or U131 (N_131,In_160,In_406);
or U132 (N_132,In_240,In_296);
nor U133 (N_133,In_670,In_342);
and U134 (N_134,In_27,In_143);
or U135 (N_135,In_846,In_398);
nand U136 (N_136,In_113,In_130);
nand U137 (N_137,In_903,In_64);
or U138 (N_138,In_972,In_784);
nor U139 (N_139,In_231,In_549);
and U140 (N_140,In_22,In_402);
nand U141 (N_141,In_764,In_748);
nand U142 (N_142,In_586,In_328);
and U143 (N_143,In_410,In_454);
and U144 (N_144,In_34,In_183);
and U145 (N_145,In_383,In_907);
or U146 (N_146,In_56,In_161);
or U147 (N_147,In_427,In_382);
and U148 (N_148,In_890,In_729);
nor U149 (N_149,In_572,In_957);
or U150 (N_150,In_30,In_954);
and U151 (N_151,In_709,In_949);
and U152 (N_152,In_786,In_967);
or U153 (N_153,In_460,In_551);
and U154 (N_154,In_790,In_131);
nand U155 (N_155,In_434,In_947);
nand U156 (N_156,In_763,In_140);
and U157 (N_157,In_191,In_754);
or U158 (N_158,In_721,In_293);
nand U159 (N_159,In_791,In_809);
nand U160 (N_160,In_550,In_28);
nand U161 (N_161,In_703,In_612);
or U162 (N_162,In_794,In_343);
or U163 (N_163,In_49,In_753);
nand U164 (N_164,In_554,In_339);
or U165 (N_165,In_16,In_11);
nand U166 (N_166,In_276,In_529);
and U167 (N_167,In_422,In_848);
nand U168 (N_168,In_277,In_241);
and U169 (N_169,In_269,In_898);
nand U170 (N_170,In_71,In_637);
and U171 (N_171,In_51,In_400);
nor U172 (N_172,In_358,In_864);
nand U173 (N_173,In_812,In_36);
or U174 (N_174,In_727,In_623);
nand U175 (N_175,In_266,In_252);
and U176 (N_176,In_69,In_145);
and U177 (N_177,In_6,In_639);
and U178 (N_178,In_189,In_636);
nor U179 (N_179,In_452,In_700);
or U180 (N_180,In_473,In_792);
nand U181 (N_181,In_280,In_157);
nor U182 (N_182,In_208,In_900);
and U183 (N_183,In_675,In_355);
or U184 (N_184,In_716,In_804);
or U185 (N_185,In_19,In_505);
nand U186 (N_186,In_607,In_20);
nor U187 (N_187,In_168,In_708);
or U188 (N_188,In_547,In_519);
nand U189 (N_189,In_614,In_137);
nor U190 (N_190,In_345,In_403);
and U191 (N_191,In_399,In_821);
nand U192 (N_192,In_321,In_943);
or U193 (N_193,In_239,In_769);
nand U194 (N_194,In_455,In_103);
or U195 (N_195,In_725,In_437);
or U196 (N_196,In_689,In_800);
nand U197 (N_197,In_394,In_314);
nand U198 (N_198,In_326,In_214);
and U199 (N_199,In_268,In_870);
and U200 (N_200,In_226,In_24);
nand U201 (N_201,In_638,In_465);
nand U202 (N_202,In_569,In_450);
nor U203 (N_203,In_141,In_543);
nand U204 (N_204,In_35,In_86);
and U205 (N_205,In_965,In_724);
or U206 (N_206,In_401,In_539);
nor U207 (N_207,In_323,In_90);
and U208 (N_208,In_660,In_249);
nand U209 (N_209,In_7,In_834);
or U210 (N_210,In_305,In_678);
and U211 (N_211,In_187,In_302);
nand U212 (N_212,In_509,In_149);
nand U213 (N_213,In_244,In_360);
or U214 (N_214,In_50,In_431);
nor U215 (N_215,In_977,In_581);
nor U216 (N_216,In_664,In_722);
nor U217 (N_217,In_444,In_340);
or U218 (N_218,In_494,In_200);
or U219 (N_219,In_54,In_844);
nand U220 (N_220,In_489,In_310);
or U221 (N_221,In_515,In_59);
nor U222 (N_222,In_271,In_471);
and U223 (N_223,In_127,In_766);
nand U224 (N_224,In_583,In_497);
and U225 (N_225,In_604,In_235);
nor U226 (N_226,In_710,In_579);
nand U227 (N_227,In_878,In_971);
nand U228 (N_228,In_657,In_555);
xor U229 (N_229,In_596,In_333);
nand U230 (N_230,In_500,In_474);
or U231 (N_231,In_956,In_807);
and U232 (N_232,In_537,In_393);
nor U233 (N_233,In_425,In_92);
nor U234 (N_234,In_162,In_805);
nand U235 (N_235,In_913,In_464);
nand U236 (N_236,In_756,In_646);
and U237 (N_237,In_990,In_737);
or U238 (N_238,In_938,In_869);
nor U239 (N_239,In_409,In_466);
and U240 (N_240,In_902,In_467);
xnor U241 (N_241,In_685,In_852);
nor U242 (N_242,In_566,In_327);
and U243 (N_243,In_883,In_311);
nand U244 (N_244,In_380,In_278);
nor U245 (N_245,In_817,In_679);
or U246 (N_246,In_225,In_780);
or U247 (N_247,In_251,In_808);
or U248 (N_248,In_788,In_171);
or U249 (N_249,In_933,In_714);
nand U250 (N_250,In_443,In_978);
nor U251 (N_251,In_468,In_854);
or U252 (N_252,In_421,In_580);
or U253 (N_253,In_507,In_138);
and U254 (N_254,In_306,In_458);
nor U255 (N_255,In_895,In_910);
nand U256 (N_256,In_2,In_952);
and U257 (N_257,In_559,In_438);
or U258 (N_258,In_882,In_562);
and U259 (N_259,In_540,In_363);
or U260 (N_260,In_435,In_411);
and U261 (N_261,In_142,In_608);
nor U262 (N_262,In_186,In_365);
and U263 (N_263,In_423,In_205);
and U264 (N_264,In_841,In_973);
and U265 (N_265,In_369,In_526);
or U266 (N_266,In_372,In_731);
and U267 (N_267,In_206,In_192);
nand U268 (N_268,In_154,In_881);
nor U269 (N_269,In_611,In_704);
and U270 (N_270,In_88,In_97);
nand U271 (N_271,In_46,In_463);
nor U272 (N_272,In_538,In_234);
nand U273 (N_273,In_948,In_366);
and U274 (N_274,In_322,In_217);
and U275 (N_275,In_905,In_598);
nand U276 (N_276,In_782,In_9);
nor U277 (N_277,In_496,In_502);
nand U278 (N_278,In_139,In_574);
and U279 (N_279,In_917,In_613);
and U280 (N_280,In_457,In_477);
or U281 (N_281,In_250,In_641);
nor U282 (N_282,In_723,In_906);
xnor U283 (N_283,In_236,In_842);
nor U284 (N_284,In_335,In_446);
or U285 (N_285,In_770,In_172);
or U286 (N_286,In_619,In_936);
nand U287 (N_287,In_484,In_768);
nor U288 (N_288,In_680,In_248);
nor U289 (N_289,In_432,In_338);
or U290 (N_290,In_934,In_483);
and U291 (N_291,In_110,In_632);
and U292 (N_292,In_215,In_147);
and U293 (N_293,In_691,In_652);
and U294 (N_294,In_698,In_93);
nor U295 (N_295,In_418,In_755);
nand U296 (N_296,In_545,In_324);
nand U297 (N_297,In_453,In_229);
and U298 (N_298,In_582,In_860);
or U299 (N_299,In_58,In_578);
nand U300 (N_300,In_351,In_70);
nand U301 (N_301,In_300,In_940);
and U302 (N_302,In_993,In_803);
or U303 (N_303,In_599,In_194);
or U304 (N_304,In_294,In_856);
nor U305 (N_305,In_589,In_253);
and U306 (N_306,In_592,In_416);
nand U307 (N_307,In_795,In_944);
or U308 (N_308,In_374,In_273);
and U309 (N_309,In_158,In_245);
and U310 (N_310,In_818,In_697);
or U311 (N_311,In_224,In_553);
or U312 (N_312,In_922,In_395);
nand U313 (N_313,In_602,In_896);
nand U314 (N_314,In_81,In_706);
or U315 (N_315,In_789,In_695);
and U316 (N_316,In_544,In_516);
and U317 (N_317,In_254,In_849);
and U318 (N_318,In_964,In_590);
nor U319 (N_319,In_462,In_96);
or U320 (N_320,In_874,In_227);
nand U321 (N_321,In_316,In_966);
or U322 (N_322,In_772,In_707);
nand U323 (N_323,In_825,In_546);
or U324 (N_324,In_12,In_330);
nand U325 (N_325,In_298,In_392);
and U326 (N_326,In_414,In_204);
nor U327 (N_327,In_829,In_151);
or U328 (N_328,In_858,In_337);
nand U329 (N_329,In_491,In_676);
or U330 (N_330,In_931,In_523);
nand U331 (N_331,In_530,In_404);
or U332 (N_332,In_758,In_238);
nor U333 (N_333,In_388,In_833);
or U334 (N_334,In_57,In_743);
nor U335 (N_335,In_951,In_984);
and U336 (N_336,In_778,In_867);
nor U337 (N_337,In_356,In_739);
and U338 (N_338,In_174,In_469);
and U339 (N_339,In_932,In_969);
and U340 (N_340,In_150,In_991);
or U341 (N_341,In_979,In_955);
or U342 (N_342,In_610,In_348);
nand U343 (N_343,In_488,In_503);
nor U344 (N_344,In_859,In_618);
and U345 (N_345,In_761,In_880);
nand U346 (N_346,In_541,In_733);
or U347 (N_347,In_381,In_304);
nor U348 (N_348,In_209,In_901);
and U349 (N_349,In_188,In_255);
and U350 (N_350,In_260,In_668);
nand U351 (N_351,In_10,In_319);
or U352 (N_352,In_350,In_26);
and U353 (N_353,In_745,In_371);
and U354 (N_354,In_267,In_822);
nor U355 (N_355,In_720,In_354);
and U356 (N_356,In_378,In_170);
nor U357 (N_357,In_568,In_995);
nand U358 (N_358,In_242,In_202);
and U359 (N_359,In_522,In_232);
and U360 (N_360,In_994,In_959);
nor U361 (N_361,In_23,In_835);
or U362 (N_362,In_456,In_702);
or U363 (N_363,In_148,In_37);
nor U364 (N_364,In_482,In_630);
nand U365 (N_365,In_647,In_207);
and U366 (N_366,In_106,In_871);
nor U367 (N_367,In_415,In_29);
and U368 (N_368,In_863,In_470);
nand U369 (N_369,In_417,In_65);
and U370 (N_370,In_892,In_18);
and U371 (N_371,In_924,In_690);
nand U372 (N_372,In_506,In_62);
nand U373 (N_373,In_459,In_785);
or U374 (N_374,In_594,In_101);
nor U375 (N_375,In_576,In_297);
and U376 (N_376,In_442,In_606);
nor U377 (N_377,In_104,In_806);
nor U378 (N_378,In_490,In_1);
or U379 (N_379,In_346,In_159);
nor U380 (N_380,In_570,In_601);
or U381 (N_381,In_781,In_461);
nor U382 (N_382,In_282,In_514);
nor U383 (N_383,In_144,In_480);
nand U384 (N_384,In_915,In_375);
nand U385 (N_385,In_256,In_762);
and U386 (N_386,In_953,In_389);
nand U387 (N_387,In_997,In_67);
nor U388 (N_388,In_89,In_535);
or U389 (N_389,In_798,In_830);
and U390 (N_390,In_831,In_303);
nand U391 (N_391,In_312,In_178);
nor U392 (N_392,In_653,In_552);
nand U393 (N_393,In_799,In_38);
nor U394 (N_394,In_605,In_521);
nand U395 (N_395,In_627,In_921);
nor U396 (N_396,In_752,In_923);
or U397 (N_397,In_120,In_237);
and U398 (N_398,In_861,In_499);
and U399 (N_399,In_665,In_937);
nor U400 (N_400,In_970,In_48);
or U401 (N_401,In_60,In_567);
nand U402 (N_402,In_288,In_987);
or U403 (N_403,In_787,In_877);
nor U404 (N_404,In_968,In_565);
nand U405 (N_405,In_654,In_884);
nand U406 (N_406,In_962,In_669);
nor U407 (N_407,In_40,In_894);
nand U408 (N_408,In_307,In_688);
nand U409 (N_409,In_989,In_195);
or U410 (N_410,In_100,In_301);
nand U411 (N_411,In_5,In_945);
or U412 (N_412,In_429,In_942);
or U413 (N_413,In_223,In_299);
or U414 (N_414,In_960,In_732);
nor U415 (N_415,In_868,In_891);
nor U416 (N_416,In_622,In_904);
nor U417 (N_417,In_930,In_391);
and U418 (N_418,In_190,In_329);
and U419 (N_419,In_620,In_649);
or U420 (N_420,In_433,In_72);
or U421 (N_421,In_616,In_624);
or U422 (N_422,In_501,In_983);
and U423 (N_423,In_82,In_377);
and U424 (N_424,In_17,In_711);
and U425 (N_425,In_219,In_175);
or U426 (N_426,In_557,In_55);
nand U427 (N_427,In_167,In_315);
nor U428 (N_428,In_134,In_283);
xor U429 (N_429,In_556,In_600);
and U430 (N_430,In_738,In_701);
or U431 (N_431,In_76,In_424);
nor U432 (N_432,In_118,In_683);
nand U433 (N_433,In_341,In_749);
and U434 (N_434,In_376,In_585);
nor U435 (N_435,In_218,In_41);
nand U436 (N_436,In_119,In_941);
nand U437 (N_437,In_179,In_640);
and U438 (N_438,In_91,In_185);
or U439 (N_439,In_512,In_352);
nand U440 (N_440,In_272,In_472);
nor U441 (N_441,In_531,In_75);
nor U442 (N_442,In_573,In_291);
nor U443 (N_443,In_815,In_481);
and U444 (N_444,In_775,In_68);
nor U445 (N_445,In_230,In_810);
and U446 (N_446,In_528,In_912);
nand U447 (N_447,In_879,In_524);
or U448 (N_448,In_920,In_385);
nand U449 (N_449,In_128,In_734);
or U450 (N_450,In_666,In_78);
and U451 (N_451,In_99,In_980);
nor U452 (N_452,In_87,In_284);
nand U453 (N_453,In_988,In_317);
and U454 (N_454,In_359,In_625);
and U455 (N_455,In_837,In_336);
nor U456 (N_456,In_289,In_832);
nand U457 (N_457,In_85,In_367);
or U458 (N_458,In_61,In_536);
and U459 (N_459,In_349,In_353);
nand U460 (N_460,In_888,In_735);
nand U461 (N_461,In_813,In_233);
nand U462 (N_462,In_135,In_246);
nand U463 (N_463,In_439,In_8);
and U464 (N_464,In_656,In_757);
or U465 (N_465,In_98,In_694);
nand U466 (N_466,In_658,In_866);
or U467 (N_467,In_826,In_320);
nor U468 (N_468,In_475,In_857);
nand U469 (N_469,In_935,In_577);
or U470 (N_470,In_824,In_981);
nand U471 (N_471,In_169,In_663);
and U472 (N_472,In_671,In_628);
nand U473 (N_473,In_742,In_270);
nor U474 (N_474,In_661,In_258);
or U475 (N_475,In_196,In_132);
or U476 (N_476,In_325,In_451);
and U477 (N_477,In_617,In_925);
and U478 (N_478,In_684,In_939);
xor U479 (N_479,In_712,In_508);
or U480 (N_480,In_571,In_692);
or U481 (N_481,In_633,In_642);
nor U482 (N_482,In_109,In_262);
nor U483 (N_483,In_587,In_347);
or U484 (N_484,In_440,In_13);
and U485 (N_485,In_693,In_32);
nand U486 (N_486,In_182,In_746);
and U487 (N_487,In_511,In_827);
nand U488 (N_488,In_851,In_909);
nand U489 (N_489,In_123,In_4);
nor U490 (N_490,In_593,In_173);
nand U491 (N_491,In_163,In_744);
or U492 (N_492,In_77,In_584);
nor U493 (N_493,In_31,In_773);
nand U494 (N_494,In_655,In_609);
nand U495 (N_495,In_44,In_510);
or U496 (N_496,In_126,In_575);
nand U497 (N_497,In_843,In_682);
and U498 (N_498,In_736,In_279);
nand U499 (N_499,In_845,In_384);
and U500 (N_500,In_173,In_196);
and U501 (N_501,In_78,In_214);
nand U502 (N_502,In_399,In_891);
nand U503 (N_503,In_899,In_442);
nor U504 (N_504,In_878,In_807);
xor U505 (N_505,In_467,In_372);
nor U506 (N_506,In_979,In_605);
nor U507 (N_507,In_331,In_946);
and U508 (N_508,In_838,In_216);
and U509 (N_509,In_191,In_806);
nand U510 (N_510,In_683,In_288);
and U511 (N_511,In_867,In_911);
nand U512 (N_512,In_57,In_706);
or U513 (N_513,In_385,In_425);
or U514 (N_514,In_112,In_398);
nand U515 (N_515,In_486,In_923);
or U516 (N_516,In_349,In_779);
and U517 (N_517,In_496,In_895);
or U518 (N_518,In_628,In_928);
and U519 (N_519,In_121,In_190);
and U520 (N_520,In_783,In_796);
nand U521 (N_521,In_180,In_296);
and U522 (N_522,In_547,In_356);
and U523 (N_523,In_8,In_416);
and U524 (N_524,In_780,In_430);
or U525 (N_525,In_875,In_620);
xnor U526 (N_526,In_994,In_32);
nand U527 (N_527,In_9,In_351);
nand U528 (N_528,In_743,In_600);
nand U529 (N_529,In_835,In_422);
nand U530 (N_530,In_142,In_983);
and U531 (N_531,In_509,In_260);
nor U532 (N_532,In_225,In_659);
and U533 (N_533,In_222,In_94);
or U534 (N_534,In_359,In_770);
nand U535 (N_535,In_900,In_416);
or U536 (N_536,In_32,In_189);
nor U537 (N_537,In_628,In_291);
or U538 (N_538,In_427,In_811);
and U539 (N_539,In_290,In_308);
nor U540 (N_540,In_613,In_71);
nand U541 (N_541,In_971,In_324);
nand U542 (N_542,In_540,In_131);
nand U543 (N_543,In_25,In_496);
nand U544 (N_544,In_956,In_925);
and U545 (N_545,In_632,In_402);
or U546 (N_546,In_835,In_464);
nand U547 (N_547,In_739,In_212);
and U548 (N_548,In_148,In_301);
nand U549 (N_549,In_806,In_775);
nor U550 (N_550,In_164,In_393);
nand U551 (N_551,In_171,In_281);
nand U552 (N_552,In_832,In_446);
nor U553 (N_553,In_317,In_360);
nand U554 (N_554,In_980,In_215);
or U555 (N_555,In_950,In_887);
and U556 (N_556,In_924,In_65);
or U557 (N_557,In_147,In_720);
or U558 (N_558,In_762,In_909);
or U559 (N_559,In_595,In_747);
nand U560 (N_560,In_565,In_981);
nand U561 (N_561,In_362,In_425);
or U562 (N_562,In_511,In_942);
and U563 (N_563,In_96,In_606);
nand U564 (N_564,In_955,In_499);
nand U565 (N_565,In_879,In_767);
and U566 (N_566,In_641,In_976);
nor U567 (N_567,In_309,In_24);
or U568 (N_568,In_685,In_935);
or U569 (N_569,In_512,In_2);
nor U570 (N_570,In_58,In_994);
nand U571 (N_571,In_446,In_674);
nand U572 (N_572,In_792,In_993);
or U573 (N_573,In_709,In_807);
or U574 (N_574,In_387,In_943);
and U575 (N_575,In_788,In_97);
nand U576 (N_576,In_142,In_284);
and U577 (N_577,In_778,In_97);
nand U578 (N_578,In_1,In_580);
or U579 (N_579,In_584,In_500);
or U580 (N_580,In_93,In_122);
nand U581 (N_581,In_994,In_339);
nor U582 (N_582,In_81,In_478);
or U583 (N_583,In_687,In_605);
and U584 (N_584,In_755,In_323);
or U585 (N_585,In_294,In_641);
or U586 (N_586,In_440,In_456);
nor U587 (N_587,In_232,In_813);
and U588 (N_588,In_689,In_304);
nand U589 (N_589,In_596,In_385);
nand U590 (N_590,In_181,In_552);
nor U591 (N_591,In_23,In_826);
and U592 (N_592,In_856,In_896);
nand U593 (N_593,In_831,In_76);
and U594 (N_594,In_915,In_183);
and U595 (N_595,In_416,In_922);
or U596 (N_596,In_130,In_207);
or U597 (N_597,In_937,In_621);
or U598 (N_598,In_237,In_693);
nand U599 (N_599,In_916,In_761);
and U600 (N_600,In_943,In_373);
xor U601 (N_601,In_125,In_99);
and U602 (N_602,In_315,In_693);
or U603 (N_603,In_779,In_431);
and U604 (N_604,In_86,In_199);
nand U605 (N_605,In_579,In_298);
nor U606 (N_606,In_140,In_930);
and U607 (N_607,In_167,In_966);
or U608 (N_608,In_244,In_193);
nand U609 (N_609,In_749,In_295);
nand U610 (N_610,In_170,In_303);
or U611 (N_611,In_156,In_722);
nand U612 (N_612,In_623,In_183);
or U613 (N_613,In_783,In_667);
nand U614 (N_614,In_829,In_122);
and U615 (N_615,In_830,In_718);
xnor U616 (N_616,In_186,In_422);
nand U617 (N_617,In_871,In_104);
nand U618 (N_618,In_265,In_719);
and U619 (N_619,In_788,In_554);
or U620 (N_620,In_28,In_676);
nand U621 (N_621,In_480,In_520);
nor U622 (N_622,In_618,In_792);
or U623 (N_623,In_576,In_706);
xnor U624 (N_624,In_145,In_728);
nand U625 (N_625,In_83,In_416);
nor U626 (N_626,In_134,In_235);
nor U627 (N_627,In_881,In_294);
and U628 (N_628,In_429,In_298);
and U629 (N_629,In_705,In_684);
nand U630 (N_630,In_338,In_200);
and U631 (N_631,In_882,In_787);
nor U632 (N_632,In_400,In_265);
nand U633 (N_633,In_169,In_601);
nor U634 (N_634,In_685,In_469);
and U635 (N_635,In_562,In_580);
nand U636 (N_636,In_313,In_29);
nor U637 (N_637,In_605,In_123);
or U638 (N_638,In_431,In_38);
nand U639 (N_639,In_234,In_901);
or U640 (N_640,In_864,In_120);
nand U641 (N_641,In_12,In_38);
or U642 (N_642,In_516,In_811);
and U643 (N_643,In_424,In_689);
or U644 (N_644,In_552,In_104);
or U645 (N_645,In_215,In_636);
and U646 (N_646,In_900,In_920);
nand U647 (N_647,In_60,In_754);
nand U648 (N_648,In_650,In_175);
or U649 (N_649,In_559,In_567);
or U650 (N_650,In_78,In_730);
or U651 (N_651,In_897,In_674);
and U652 (N_652,In_80,In_967);
xnor U653 (N_653,In_547,In_749);
and U654 (N_654,In_774,In_863);
nand U655 (N_655,In_339,In_261);
or U656 (N_656,In_978,In_202);
or U657 (N_657,In_958,In_568);
nor U658 (N_658,In_839,In_409);
or U659 (N_659,In_191,In_162);
nor U660 (N_660,In_724,In_728);
nand U661 (N_661,In_19,In_480);
or U662 (N_662,In_912,In_891);
or U663 (N_663,In_866,In_750);
nor U664 (N_664,In_843,In_271);
nor U665 (N_665,In_333,In_730);
nand U666 (N_666,In_893,In_870);
and U667 (N_667,In_653,In_42);
nor U668 (N_668,In_459,In_395);
or U669 (N_669,In_621,In_87);
nand U670 (N_670,In_398,In_424);
or U671 (N_671,In_598,In_783);
or U672 (N_672,In_634,In_151);
nand U673 (N_673,In_734,In_952);
nand U674 (N_674,In_97,In_952);
nand U675 (N_675,In_258,In_948);
nand U676 (N_676,In_13,In_268);
and U677 (N_677,In_275,In_980);
or U678 (N_678,In_103,In_41);
nand U679 (N_679,In_221,In_126);
or U680 (N_680,In_794,In_492);
and U681 (N_681,In_266,In_713);
or U682 (N_682,In_101,In_188);
or U683 (N_683,In_468,In_575);
and U684 (N_684,In_296,In_399);
nand U685 (N_685,In_327,In_17);
nor U686 (N_686,In_417,In_370);
and U687 (N_687,In_116,In_395);
and U688 (N_688,In_286,In_268);
nor U689 (N_689,In_658,In_939);
nand U690 (N_690,In_279,In_801);
nand U691 (N_691,In_840,In_283);
and U692 (N_692,In_850,In_650);
or U693 (N_693,In_769,In_93);
nand U694 (N_694,In_473,In_993);
and U695 (N_695,In_694,In_58);
and U696 (N_696,In_822,In_779);
xnor U697 (N_697,In_301,In_269);
nand U698 (N_698,In_332,In_969);
nor U699 (N_699,In_531,In_197);
xnor U700 (N_700,In_909,In_955);
and U701 (N_701,In_781,In_218);
and U702 (N_702,In_807,In_330);
and U703 (N_703,In_387,In_734);
or U704 (N_704,In_430,In_80);
nand U705 (N_705,In_984,In_236);
and U706 (N_706,In_333,In_951);
xnor U707 (N_707,In_526,In_628);
or U708 (N_708,In_395,In_904);
and U709 (N_709,In_752,In_66);
nand U710 (N_710,In_693,In_842);
or U711 (N_711,In_891,In_179);
nor U712 (N_712,In_911,In_918);
and U713 (N_713,In_46,In_237);
nor U714 (N_714,In_461,In_614);
nor U715 (N_715,In_572,In_242);
nand U716 (N_716,In_265,In_419);
nor U717 (N_717,In_535,In_182);
nand U718 (N_718,In_504,In_723);
nor U719 (N_719,In_941,In_95);
nor U720 (N_720,In_768,In_572);
nand U721 (N_721,In_452,In_737);
xor U722 (N_722,In_821,In_738);
and U723 (N_723,In_110,In_304);
nor U724 (N_724,In_407,In_228);
nor U725 (N_725,In_238,In_797);
nor U726 (N_726,In_208,In_583);
and U727 (N_727,In_100,In_411);
and U728 (N_728,In_129,In_408);
nor U729 (N_729,In_642,In_273);
xnor U730 (N_730,In_985,In_419);
nor U731 (N_731,In_72,In_147);
nor U732 (N_732,In_109,In_792);
nand U733 (N_733,In_150,In_964);
and U734 (N_734,In_782,In_741);
and U735 (N_735,In_187,In_311);
and U736 (N_736,In_879,In_475);
and U737 (N_737,In_826,In_80);
nand U738 (N_738,In_948,In_200);
nand U739 (N_739,In_828,In_117);
nor U740 (N_740,In_262,In_309);
nand U741 (N_741,In_677,In_11);
nor U742 (N_742,In_344,In_851);
or U743 (N_743,In_112,In_290);
nand U744 (N_744,In_591,In_540);
or U745 (N_745,In_183,In_917);
nor U746 (N_746,In_28,In_621);
and U747 (N_747,In_194,In_958);
nand U748 (N_748,In_484,In_13);
nor U749 (N_749,In_308,In_950);
and U750 (N_750,In_958,In_939);
nor U751 (N_751,In_614,In_581);
nor U752 (N_752,In_83,In_391);
and U753 (N_753,In_436,In_219);
or U754 (N_754,In_610,In_228);
and U755 (N_755,In_668,In_982);
nor U756 (N_756,In_150,In_200);
nand U757 (N_757,In_84,In_680);
nor U758 (N_758,In_964,In_469);
nor U759 (N_759,In_256,In_908);
nor U760 (N_760,In_627,In_636);
nor U761 (N_761,In_934,In_305);
xor U762 (N_762,In_392,In_262);
nand U763 (N_763,In_331,In_199);
and U764 (N_764,In_91,In_993);
or U765 (N_765,In_501,In_203);
and U766 (N_766,In_452,In_284);
or U767 (N_767,In_871,In_309);
and U768 (N_768,In_137,In_332);
or U769 (N_769,In_328,In_514);
nor U770 (N_770,In_570,In_93);
and U771 (N_771,In_864,In_781);
or U772 (N_772,In_849,In_933);
or U773 (N_773,In_23,In_828);
and U774 (N_774,In_52,In_645);
or U775 (N_775,In_680,In_383);
nand U776 (N_776,In_903,In_350);
nand U777 (N_777,In_802,In_217);
nand U778 (N_778,In_65,In_704);
or U779 (N_779,In_473,In_560);
and U780 (N_780,In_697,In_496);
and U781 (N_781,In_961,In_258);
nand U782 (N_782,In_64,In_315);
nor U783 (N_783,In_94,In_977);
or U784 (N_784,In_328,In_868);
nor U785 (N_785,In_103,In_846);
or U786 (N_786,In_210,In_18);
or U787 (N_787,In_207,In_858);
and U788 (N_788,In_88,In_773);
and U789 (N_789,In_848,In_453);
and U790 (N_790,In_283,In_810);
nor U791 (N_791,In_298,In_802);
xnor U792 (N_792,In_47,In_614);
nand U793 (N_793,In_252,In_347);
and U794 (N_794,In_368,In_718);
nand U795 (N_795,In_593,In_681);
or U796 (N_796,In_331,In_979);
or U797 (N_797,In_131,In_832);
nand U798 (N_798,In_440,In_482);
and U799 (N_799,In_617,In_299);
and U800 (N_800,In_464,In_568);
and U801 (N_801,In_848,In_497);
and U802 (N_802,In_679,In_27);
nand U803 (N_803,In_714,In_944);
nand U804 (N_804,In_117,In_583);
nand U805 (N_805,In_564,In_596);
or U806 (N_806,In_742,In_565);
or U807 (N_807,In_343,In_525);
nand U808 (N_808,In_193,In_960);
or U809 (N_809,In_938,In_857);
or U810 (N_810,In_460,In_876);
or U811 (N_811,In_329,In_535);
and U812 (N_812,In_966,In_224);
and U813 (N_813,In_557,In_696);
or U814 (N_814,In_45,In_582);
nand U815 (N_815,In_63,In_369);
nor U816 (N_816,In_356,In_748);
or U817 (N_817,In_256,In_176);
nand U818 (N_818,In_408,In_425);
and U819 (N_819,In_117,In_873);
or U820 (N_820,In_41,In_631);
nand U821 (N_821,In_442,In_184);
nand U822 (N_822,In_53,In_744);
and U823 (N_823,In_851,In_904);
nor U824 (N_824,In_810,In_582);
nor U825 (N_825,In_464,In_978);
and U826 (N_826,In_302,In_249);
nand U827 (N_827,In_596,In_379);
and U828 (N_828,In_835,In_785);
or U829 (N_829,In_274,In_669);
nor U830 (N_830,In_411,In_552);
nand U831 (N_831,In_102,In_361);
and U832 (N_832,In_75,In_550);
nand U833 (N_833,In_448,In_301);
nand U834 (N_834,In_631,In_422);
or U835 (N_835,In_93,In_500);
nor U836 (N_836,In_112,In_47);
nand U837 (N_837,In_207,In_51);
and U838 (N_838,In_932,In_974);
and U839 (N_839,In_922,In_274);
nor U840 (N_840,In_687,In_51);
and U841 (N_841,In_587,In_252);
or U842 (N_842,In_694,In_41);
nor U843 (N_843,In_740,In_697);
nor U844 (N_844,In_456,In_215);
nor U845 (N_845,In_260,In_972);
and U846 (N_846,In_395,In_884);
and U847 (N_847,In_547,In_75);
or U848 (N_848,In_13,In_382);
and U849 (N_849,In_577,In_525);
and U850 (N_850,In_362,In_663);
or U851 (N_851,In_77,In_964);
and U852 (N_852,In_725,In_831);
or U853 (N_853,In_500,In_783);
nor U854 (N_854,In_179,In_994);
nor U855 (N_855,In_477,In_70);
and U856 (N_856,In_774,In_664);
nand U857 (N_857,In_886,In_145);
nor U858 (N_858,In_112,In_909);
nor U859 (N_859,In_84,In_63);
nand U860 (N_860,In_155,In_748);
nor U861 (N_861,In_501,In_534);
xor U862 (N_862,In_507,In_543);
or U863 (N_863,In_145,In_834);
nand U864 (N_864,In_86,In_411);
and U865 (N_865,In_311,In_756);
and U866 (N_866,In_661,In_677);
or U867 (N_867,In_132,In_531);
nor U868 (N_868,In_246,In_929);
or U869 (N_869,In_888,In_149);
or U870 (N_870,In_790,In_89);
nand U871 (N_871,In_359,In_163);
nor U872 (N_872,In_698,In_770);
and U873 (N_873,In_533,In_428);
or U874 (N_874,In_427,In_112);
and U875 (N_875,In_996,In_991);
nand U876 (N_876,In_522,In_649);
and U877 (N_877,In_522,In_241);
or U878 (N_878,In_21,In_359);
or U879 (N_879,In_700,In_297);
or U880 (N_880,In_236,In_632);
and U881 (N_881,In_6,In_615);
nor U882 (N_882,In_501,In_498);
nor U883 (N_883,In_881,In_309);
or U884 (N_884,In_139,In_838);
or U885 (N_885,In_569,In_36);
nand U886 (N_886,In_210,In_317);
nor U887 (N_887,In_378,In_55);
or U888 (N_888,In_737,In_476);
and U889 (N_889,In_270,In_909);
nand U890 (N_890,In_84,In_705);
xor U891 (N_891,In_127,In_504);
and U892 (N_892,In_410,In_729);
nand U893 (N_893,In_401,In_983);
and U894 (N_894,In_51,In_853);
or U895 (N_895,In_102,In_16);
or U896 (N_896,In_99,In_765);
nand U897 (N_897,In_519,In_550);
and U898 (N_898,In_158,In_566);
nor U899 (N_899,In_572,In_718);
or U900 (N_900,In_536,In_325);
or U901 (N_901,In_199,In_381);
or U902 (N_902,In_337,In_730);
and U903 (N_903,In_335,In_320);
xor U904 (N_904,In_910,In_785);
and U905 (N_905,In_137,In_236);
and U906 (N_906,In_68,In_438);
xnor U907 (N_907,In_54,In_682);
or U908 (N_908,In_482,In_891);
and U909 (N_909,In_685,In_853);
or U910 (N_910,In_756,In_395);
or U911 (N_911,In_278,In_52);
nand U912 (N_912,In_248,In_837);
nand U913 (N_913,In_136,In_62);
or U914 (N_914,In_233,In_724);
and U915 (N_915,In_51,In_237);
or U916 (N_916,In_173,In_421);
nor U917 (N_917,In_426,In_434);
or U918 (N_918,In_887,In_301);
or U919 (N_919,In_257,In_492);
xnor U920 (N_920,In_715,In_333);
nor U921 (N_921,In_464,In_130);
or U922 (N_922,In_83,In_573);
and U923 (N_923,In_270,In_142);
nand U924 (N_924,In_131,In_564);
or U925 (N_925,In_570,In_477);
and U926 (N_926,In_872,In_927);
and U927 (N_927,In_192,In_829);
nor U928 (N_928,In_526,In_959);
or U929 (N_929,In_774,In_482);
nor U930 (N_930,In_791,In_463);
and U931 (N_931,In_259,In_723);
nand U932 (N_932,In_888,In_419);
or U933 (N_933,In_334,In_624);
and U934 (N_934,In_833,In_416);
nand U935 (N_935,In_317,In_679);
nor U936 (N_936,In_757,In_349);
nand U937 (N_937,In_418,In_357);
nand U938 (N_938,In_730,In_434);
nor U939 (N_939,In_154,In_440);
and U940 (N_940,In_775,In_397);
nor U941 (N_941,In_751,In_693);
or U942 (N_942,In_833,In_887);
and U943 (N_943,In_751,In_929);
and U944 (N_944,In_863,In_577);
nand U945 (N_945,In_96,In_457);
nand U946 (N_946,In_947,In_433);
nand U947 (N_947,In_106,In_786);
and U948 (N_948,In_798,In_406);
nor U949 (N_949,In_542,In_1);
and U950 (N_950,In_676,In_919);
or U951 (N_951,In_371,In_792);
nand U952 (N_952,In_491,In_874);
nor U953 (N_953,In_991,In_334);
and U954 (N_954,In_974,In_730);
nand U955 (N_955,In_355,In_324);
nor U956 (N_956,In_30,In_354);
or U957 (N_957,In_881,In_815);
or U958 (N_958,In_517,In_191);
nand U959 (N_959,In_721,In_552);
or U960 (N_960,In_566,In_587);
and U961 (N_961,In_970,In_702);
nor U962 (N_962,In_762,In_223);
and U963 (N_963,In_167,In_225);
or U964 (N_964,In_712,In_983);
nor U965 (N_965,In_932,In_95);
nand U966 (N_966,In_690,In_559);
and U967 (N_967,In_337,In_756);
nand U968 (N_968,In_343,In_922);
and U969 (N_969,In_829,In_76);
nand U970 (N_970,In_761,In_456);
nor U971 (N_971,In_979,In_18);
nand U972 (N_972,In_205,In_851);
nor U973 (N_973,In_375,In_405);
nand U974 (N_974,In_740,In_815);
nor U975 (N_975,In_14,In_854);
nand U976 (N_976,In_922,In_317);
xor U977 (N_977,In_69,In_177);
and U978 (N_978,In_725,In_574);
nor U979 (N_979,In_640,In_393);
nor U980 (N_980,In_183,In_459);
nor U981 (N_981,In_461,In_736);
and U982 (N_982,In_656,In_786);
or U983 (N_983,In_953,In_763);
nand U984 (N_984,In_176,In_153);
nor U985 (N_985,In_401,In_824);
and U986 (N_986,In_858,In_234);
and U987 (N_987,In_811,In_789);
nor U988 (N_988,In_576,In_283);
nor U989 (N_989,In_571,In_767);
or U990 (N_990,In_897,In_940);
nor U991 (N_991,In_48,In_401);
nand U992 (N_992,In_766,In_493);
and U993 (N_993,In_753,In_126);
nand U994 (N_994,In_599,In_757);
nand U995 (N_995,In_742,In_76);
and U996 (N_996,In_193,In_219);
nor U997 (N_997,In_315,In_265);
and U998 (N_998,In_531,In_427);
nand U999 (N_999,In_690,In_909);
or U1000 (N_1000,N_57,N_34);
nor U1001 (N_1001,N_310,N_2);
or U1002 (N_1002,N_198,N_317);
and U1003 (N_1003,N_155,N_214);
nand U1004 (N_1004,N_363,N_845);
or U1005 (N_1005,N_351,N_466);
or U1006 (N_1006,N_809,N_19);
nor U1007 (N_1007,N_407,N_801);
nor U1008 (N_1008,N_725,N_773);
nand U1009 (N_1009,N_192,N_373);
or U1010 (N_1010,N_0,N_425);
or U1011 (N_1011,N_322,N_319);
nor U1012 (N_1012,N_247,N_877);
nor U1013 (N_1013,N_372,N_481);
nand U1014 (N_1014,N_14,N_768);
nand U1015 (N_1015,N_510,N_259);
or U1016 (N_1016,N_131,N_978);
or U1017 (N_1017,N_638,N_513);
and U1018 (N_1018,N_691,N_541);
nor U1019 (N_1019,N_552,N_222);
and U1020 (N_1020,N_1,N_819);
and U1021 (N_1021,N_187,N_128);
nor U1022 (N_1022,N_227,N_955);
nand U1023 (N_1023,N_665,N_921);
nand U1024 (N_1024,N_124,N_353);
and U1025 (N_1025,N_190,N_29);
xor U1026 (N_1026,N_677,N_284);
nand U1027 (N_1027,N_778,N_365);
nor U1028 (N_1028,N_200,N_573);
nor U1029 (N_1029,N_603,N_436);
and U1030 (N_1030,N_199,N_586);
or U1031 (N_1031,N_428,N_554);
or U1032 (N_1032,N_35,N_566);
nor U1033 (N_1033,N_663,N_143);
and U1034 (N_1034,N_637,N_672);
and U1035 (N_1035,N_551,N_450);
nor U1036 (N_1036,N_816,N_742);
and U1037 (N_1037,N_972,N_864);
or U1038 (N_1038,N_21,N_460);
and U1039 (N_1039,N_485,N_430);
or U1040 (N_1040,N_984,N_895);
nor U1041 (N_1041,N_10,N_257);
and U1042 (N_1042,N_25,N_901);
xnor U1043 (N_1043,N_426,N_91);
nor U1044 (N_1044,N_60,N_817);
or U1045 (N_1045,N_17,N_100);
and U1046 (N_1046,N_869,N_431);
nor U1047 (N_1047,N_120,N_255);
and U1048 (N_1048,N_797,N_508);
or U1049 (N_1049,N_735,N_888);
and U1050 (N_1050,N_467,N_754);
nor U1051 (N_1051,N_746,N_115);
or U1052 (N_1052,N_195,N_739);
or U1053 (N_1053,N_612,N_770);
or U1054 (N_1054,N_920,N_592);
and U1055 (N_1055,N_313,N_463);
or U1056 (N_1056,N_579,N_610);
or U1057 (N_1057,N_223,N_653);
or U1058 (N_1058,N_82,N_681);
and U1059 (N_1059,N_418,N_49);
nand U1060 (N_1060,N_881,N_46);
and U1061 (N_1061,N_170,N_557);
or U1062 (N_1062,N_7,N_184);
nand U1063 (N_1063,N_364,N_772);
nand U1064 (N_1064,N_549,N_102);
or U1065 (N_1065,N_687,N_133);
and U1066 (N_1066,N_647,N_333);
nor U1067 (N_1067,N_890,N_639);
nor U1068 (N_1068,N_504,N_759);
or U1069 (N_1069,N_400,N_537);
and U1070 (N_1070,N_235,N_3);
or U1071 (N_1071,N_420,N_655);
nor U1072 (N_1072,N_138,N_590);
and U1073 (N_1073,N_849,N_623);
and U1074 (N_1074,N_501,N_453);
or U1075 (N_1075,N_862,N_747);
nand U1076 (N_1076,N_445,N_959);
nor U1077 (N_1077,N_424,N_990);
or U1078 (N_1078,N_52,N_185);
nor U1079 (N_1079,N_926,N_547);
nor U1080 (N_1080,N_705,N_375);
and U1081 (N_1081,N_873,N_381);
nand U1082 (N_1082,N_753,N_38);
or U1083 (N_1083,N_414,N_531);
nor U1084 (N_1084,N_497,N_615);
nand U1085 (N_1085,N_847,N_749);
or U1086 (N_1086,N_44,N_838);
nand U1087 (N_1087,N_345,N_848);
and U1088 (N_1088,N_927,N_871);
nor U1089 (N_1089,N_833,N_237);
and U1090 (N_1090,N_93,N_514);
and U1091 (N_1091,N_495,N_65);
nand U1092 (N_1092,N_795,N_904);
nor U1093 (N_1093,N_201,N_180);
or U1094 (N_1094,N_477,N_852);
nand U1095 (N_1095,N_347,N_692);
or U1096 (N_1096,N_587,N_708);
nor U1097 (N_1097,N_490,N_12);
nor U1098 (N_1098,N_397,N_814);
or U1099 (N_1099,N_661,N_51);
and U1100 (N_1100,N_188,N_225);
nand U1101 (N_1101,N_776,N_412);
or U1102 (N_1102,N_475,N_202);
or U1103 (N_1103,N_876,N_197);
nor U1104 (N_1104,N_265,N_24);
nand U1105 (N_1105,N_534,N_89);
or U1106 (N_1106,N_962,N_470);
or U1107 (N_1107,N_50,N_516);
and U1108 (N_1108,N_289,N_238);
nand U1109 (N_1109,N_448,N_897);
and U1110 (N_1110,N_973,N_713);
or U1111 (N_1111,N_951,N_218);
or U1112 (N_1112,N_991,N_480);
nand U1113 (N_1113,N_230,N_8);
nand U1114 (N_1114,N_368,N_168);
nor U1115 (N_1115,N_611,N_521);
nor U1116 (N_1116,N_454,N_285);
and U1117 (N_1117,N_686,N_792);
nand U1118 (N_1118,N_99,N_244);
and U1119 (N_1119,N_787,N_800);
and U1120 (N_1120,N_483,N_828);
and U1121 (N_1121,N_58,N_731);
or U1122 (N_1122,N_613,N_757);
nor U1123 (N_1123,N_429,N_164);
nand U1124 (N_1124,N_829,N_179);
nor U1125 (N_1125,N_473,N_633);
nand U1126 (N_1126,N_376,N_660);
or U1127 (N_1127,N_857,N_494);
or U1128 (N_1128,N_206,N_277);
or U1129 (N_1129,N_616,N_90);
or U1130 (N_1130,N_918,N_191);
nand U1131 (N_1131,N_174,N_346);
and U1132 (N_1132,N_335,N_872);
nor U1133 (N_1133,N_894,N_181);
and U1134 (N_1134,N_961,N_156);
and U1135 (N_1135,N_362,N_323);
or U1136 (N_1136,N_134,N_506);
nor U1137 (N_1137,N_818,N_628);
nor U1138 (N_1138,N_246,N_59);
nor U1139 (N_1139,N_387,N_752);
nor U1140 (N_1140,N_404,N_956);
nor U1141 (N_1141,N_261,N_964);
nand U1142 (N_1142,N_940,N_5);
nand U1143 (N_1143,N_356,N_437);
nor U1144 (N_1144,N_953,N_491);
nand U1145 (N_1145,N_204,N_925);
or U1146 (N_1146,N_875,N_777);
nand U1147 (N_1147,N_807,N_502);
nor U1148 (N_1148,N_6,N_699);
or U1149 (N_1149,N_329,N_975);
and U1150 (N_1150,N_910,N_331);
nor U1151 (N_1151,N_600,N_841);
nand U1152 (N_1152,N_283,N_813);
nor U1153 (N_1153,N_576,N_649);
nor U1154 (N_1154,N_83,N_127);
and U1155 (N_1155,N_249,N_636);
nor U1156 (N_1156,N_402,N_118);
nor U1157 (N_1157,N_574,N_824);
nand U1158 (N_1158,N_923,N_339);
or U1159 (N_1159,N_169,N_462);
nor U1160 (N_1160,N_342,N_76);
and U1161 (N_1161,N_733,N_891);
nor U1162 (N_1162,N_427,N_966);
and U1163 (N_1163,N_555,N_384);
or U1164 (N_1164,N_33,N_258);
nor U1165 (N_1165,N_468,N_388);
nand U1166 (N_1166,N_389,N_784);
or U1167 (N_1167,N_658,N_609);
nand U1168 (N_1168,N_79,N_417);
nor U1169 (N_1169,N_144,N_654);
nand U1170 (N_1170,N_666,N_619);
and U1171 (N_1171,N_657,N_520);
or U1172 (N_1172,N_606,N_906);
or U1173 (N_1173,N_523,N_446);
or U1174 (N_1174,N_294,N_464);
and U1175 (N_1175,N_30,N_648);
nor U1176 (N_1176,N_160,N_87);
nand U1177 (N_1177,N_720,N_775);
and U1178 (N_1178,N_456,N_64);
and U1179 (N_1179,N_908,N_769);
nor U1180 (N_1180,N_511,N_844);
nand U1181 (N_1181,N_86,N_561);
and U1182 (N_1182,N_267,N_126);
nand U1183 (N_1183,N_799,N_780);
nor U1184 (N_1184,N_765,N_444);
nand U1185 (N_1185,N_183,N_315);
nand U1186 (N_1186,N_545,N_148);
nor U1187 (N_1187,N_309,N_320);
nand U1188 (N_1188,N_915,N_23);
nor U1189 (N_1189,N_26,N_789);
nor U1190 (N_1190,N_682,N_321);
nor U1191 (N_1191,N_909,N_167);
or U1192 (N_1192,N_885,N_78);
nand U1193 (N_1193,N_843,N_994);
or U1194 (N_1194,N_938,N_583);
or U1195 (N_1195,N_934,N_960);
and U1196 (N_1196,N_624,N_211);
or U1197 (N_1197,N_336,N_620);
nor U1198 (N_1198,N_117,N_919);
and U1199 (N_1199,N_738,N_499);
or U1200 (N_1200,N_842,N_865);
nor U1201 (N_1201,N_465,N_945);
nand U1202 (N_1202,N_602,N_782);
nand U1203 (N_1203,N_965,N_748);
or U1204 (N_1204,N_358,N_532);
nor U1205 (N_1205,N_233,N_861);
and U1206 (N_1206,N_348,N_986);
nand U1207 (N_1207,N_745,N_860);
nand U1208 (N_1208,N_589,N_998);
and U1209 (N_1209,N_729,N_39);
nand U1210 (N_1210,N_874,N_288);
or U1211 (N_1211,N_297,N_601);
and U1212 (N_1212,N_379,N_312);
and U1213 (N_1213,N_264,N_162);
and U1214 (N_1214,N_883,N_292);
nand U1215 (N_1215,N_675,N_300);
nor U1216 (N_1216,N_367,N_736);
and U1217 (N_1217,N_689,N_798);
and U1218 (N_1218,N_559,N_643);
and U1219 (N_1219,N_219,N_4);
or U1220 (N_1220,N_413,N_922);
nand U1221 (N_1221,N_604,N_526);
or U1222 (N_1222,N_318,N_421);
and U1223 (N_1223,N_101,N_868);
nand U1224 (N_1224,N_125,N_434);
nor U1225 (N_1225,N_617,N_669);
nor U1226 (N_1226,N_811,N_271);
nand U1227 (N_1227,N_498,N_152);
nand U1228 (N_1228,N_147,N_54);
nor U1229 (N_1229,N_301,N_108);
and U1230 (N_1230,N_471,N_145);
or U1231 (N_1231,N_382,N_361);
nor U1232 (N_1232,N_716,N_154);
nand U1233 (N_1233,N_251,N_110);
or U1234 (N_1234,N_298,N_571);
nand U1235 (N_1235,N_762,N_136);
or U1236 (N_1236,N_596,N_567);
or U1237 (N_1237,N_366,N_478);
nand U1238 (N_1238,N_970,N_774);
and U1239 (N_1239,N_761,N_245);
or U1240 (N_1240,N_410,N_812);
and U1241 (N_1241,N_900,N_791);
nand U1242 (N_1242,N_538,N_393);
nand U1243 (N_1243,N_31,N_979);
and U1244 (N_1244,N_597,N_703);
nand U1245 (N_1245,N_176,N_296);
nand U1246 (N_1246,N_827,N_548);
nor U1247 (N_1247,N_539,N_435);
and U1248 (N_1248,N_546,N_898);
xnor U1249 (N_1249,N_482,N_931);
or U1250 (N_1250,N_77,N_447);
or U1251 (N_1251,N_73,N_664);
nor U1252 (N_1252,N_291,N_710);
nor U1253 (N_1253,N_305,N_751);
nand U1254 (N_1254,N_679,N_378);
nand U1255 (N_1255,N_268,N_27);
nor U1256 (N_1256,N_805,N_338);
or U1257 (N_1257,N_667,N_702);
nor U1258 (N_1258,N_493,N_455);
nor U1259 (N_1259,N_142,N_943);
nand U1260 (N_1260,N_999,N_693);
or U1261 (N_1261,N_273,N_887);
and U1262 (N_1262,N_451,N_71);
or U1263 (N_1263,N_582,N_670);
nor U1264 (N_1264,N_967,N_377);
nand U1265 (N_1265,N_47,N_210);
or U1266 (N_1266,N_70,N_61);
or U1267 (N_1267,N_422,N_879);
nand U1268 (N_1268,N_240,N_936);
nor U1269 (N_1269,N_216,N_645);
nor U1270 (N_1270,N_355,N_568);
or U1271 (N_1271,N_157,N_28);
nor U1272 (N_1272,N_260,N_280);
nand U1273 (N_1273,N_607,N_826);
nand U1274 (N_1274,N_831,N_734);
or U1275 (N_1275,N_153,N_969);
and U1276 (N_1276,N_928,N_439);
or U1277 (N_1277,N_149,N_275);
nor U1278 (N_1278,N_656,N_189);
or U1279 (N_1279,N_272,N_109);
and U1280 (N_1280,N_698,N_618);
nor U1281 (N_1281,N_785,N_977);
or U1282 (N_1282,N_405,N_282);
or U1283 (N_1283,N_253,N_53);
nand U1284 (N_1284,N_553,N_987);
nand U1285 (N_1285,N_727,N_263);
or U1286 (N_1286,N_760,N_853);
or U1287 (N_1287,N_239,N_942);
or U1288 (N_1288,N_644,N_886);
or U1289 (N_1289,N_578,N_349);
nand U1290 (N_1290,N_113,N_182);
nand U1291 (N_1291,N_903,N_171);
or U1292 (N_1292,N_562,N_194);
and U1293 (N_1293,N_242,N_896);
nand U1294 (N_1294,N_40,N_486);
nand U1295 (N_1295,N_254,N_146);
and U1296 (N_1296,N_88,N_905);
or U1297 (N_1297,N_764,N_755);
nand U1298 (N_1298,N_767,N_403);
or U1299 (N_1299,N_357,N_719);
nor U1300 (N_1300,N_515,N_139);
nor U1301 (N_1301,N_850,N_302);
and U1302 (N_1302,N_593,N_457);
or U1303 (N_1303,N_166,N_43);
nor U1304 (N_1304,N_196,N_779);
nand U1305 (N_1305,N_121,N_981);
nand U1306 (N_1306,N_803,N_438);
and U1307 (N_1307,N_411,N_947);
or U1308 (N_1308,N_172,N_856);
and U1309 (N_1309,N_808,N_458);
nor U1310 (N_1310,N_794,N_671);
and U1311 (N_1311,N_415,N_311);
nand U1312 (N_1312,N_867,N_524);
or U1313 (N_1313,N_804,N_634);
or U1314 (N_1314,N_581,N_983);
and U1315 (N_1315,N_328,N_392);
or U1316 (N_1316,N_723,N_252);
or U1317 (N_1317,N_825,N_533);
and U1318 (N_1318,N_766,N_122);
or U1319 (N_1319,N_878,N_893);
xor U1320 (N_1320,N_806,N_229);
and U1321 (N_1321,N_85,N_996);
nand U1322 (N_1322,N_750,N_371);
nor U1323 (N_1323,N_509,N_16);
and U1324 (N_1324,N_846,N_714);
or U1325 (N_1325,N_62,N_783);
or U1326 (N_1326,N_651,N_324);
nor U1327 (N_1327,N_67,N_32);
xor U1328 (N_1328,N_650,N_395);
nor U1329 (N_1329,N_209,N_221);
nand U1330 (N_1330,N_68,N_870);
nand U1331 (N_1331,N_408,N_13);
nand U1332 (N_1332,N_659,N_530);
nand U1333 (N_1333,N_112,N_383);
nand U1334 (N_1334,N_614,N_917);
and U1335 (N_1335,N_540,N_158);
and U1336 (N_1336,N_550,N_711);
nand U1337 (N_1337,N_695,N_224);
nor U1338 (N_1338,N_461,N_832);
and U1339 (N_1339,N_688,N_274);
and U1340 (N_1340,N_884,N_758);
nand U1341 (N_1341,N_55,N_406);
nor U1342 (N_1342,N_823,N_243);
nand U1343 (N_1343,N_810,N_95);
or U1344 (N_1344,N_307,N_880);
nand U1345 (N_1345,N_902,N_565);
or U1346 (N_1346,N_343,N_584);
nor U1347 (N_1347,N_968,N_81);
or U1348 (N_1348,N_939,N_678);
nor U1349 (N_1349,N_858,N_443);
nor U1350 (N_1350,N_132,N_74);
or U1351 (N_1351,N_982,N_684);
and U1352 (N_1352,N_341,N_855);
nor U1353 (N_1353,N_866,N_354);
nand U1354 (N_1354,N_360,N_327);
or U1355 (N_1355,N_18,N_889);
or U1356 (N_1356,N_899,N_840);
nand U1357 (N_1357,N_863,N_525);
nor U1358 (N_1358,N_588,N_488);
and U1359 (N_1359,N_56,N_957);
xnor U1360 (N_1360,N_69,N_84);
nand U1361 (N_1361,N_627,N_701);
nor U1362 (N_1362,N_911,N_625);
or U1363 (N_1363,N_944,N_706);
and U1364 (N_1364,N_116,N_226);
and U1365 (N_1365,N_177,N_646);
or U1366 (N_1366,N_286,N_790);
nand U1367 (N_1367,N_950,N_788);
and U1368 (N_1368,N_212,N_22);
nand U1369 (N_1369,N_141,N_15);
and U1370 (N_1370,N_217,N_270);
and U1371 (N_1371,N_709,N_203);
nand U1372 (N_1372,N_556,N_935);
nand U1373 (N_1373,N_985,N_63);
nand U1374 (N_1374,N_835,N_48);
and U1375 (N_1375,N_92,N_266);
and U1376 (N_1376,N_11,N_220);
or U1377 (N_1377,N_963,N_111);
or U1378 (N_1378,N_952,N_449);
xor U1379 (N_1379,N_815,N_304);
or U1380 (N_1380,N_173,N_676);
and U1381 (N_1381,N_186,N_924);
nand U1382 (N_1382,N_42,N_390);
nor U1383 (N_1383,N_741,N_949);
or U1384 (N_1384,N_907,N_522);
nand U1385 (N_1385,N_279,N_380);
xor U1386 (N_1386,N_718,N_20);
or U1387 (N_1387,N_932,N_995);
nand U1388 (N_1388,N_72,N_80);
or U1389 (N_1389,N_228,N_107);
and U1390 (N_1390,N_370,N_974);
nand U1391 (N_1391,N_631,N_241);
or U1392 (N_1392,N_756,N_575);
nor U1393 (N_1393,N_572,N_822);
and U1394 (N_1394,N_635,N_930);
and U1395 (N_1395,N_299,N_642);
or U1396 (N_1396,N_640,N_599);
nor U1397 (N_1397,N_316,N_690);
and U1398 (N_1398,N_560,N_401);
or U1399 (N_1399,N_771,N_276);
and U1400 (N_1400,N_912,N_459);
and U1401 (N_1401,N_326,N_595);
and U1402 (N_1402,N_608,N_442);
and U1403 (N_1403,N_704,N_859);
nand U1404 (N_1404,N_992,N_674);
and U1405 (N_1405,N_489,N_834);
or U1406 (N_1406,N_854,N_913);
and U1407 (N_1407,N_350,N_452);
and U1408 (N_1408,N_668,N_839);
and U1409 (N_1409,N_487,N_9);
nand U1410 (N_1410,N_632,N_662);
and U1411 (N_1411,N_989,N_802);
nand U1412 (N_1412,N_96,N_45);
or U1413 (N_1413,N_507,N_256);
or U1414 (N_1414,N_558,N_399);
or U1415 (N_1415,N_193,N_993);
and U1416 (N_1416,N_290,N_94);
nand U1417 (N_1417,N_104,N_916);
nor U1418 (N_1418,N_937,N_505);
nor U1419 (N_1419,N_208,N_744);
nand U1420 (N_1420,N_369,N_432);
and U1421 (N_1421,N_793,N_732);
or U1422 (N_1422,N_106,N_398);
or U1423 (N_1423,N_374,N_715);
and U1424 (N_1424,N_536,N_278);
xnor U1425 (N_1425,N_626,N_352);
or U1426 (N_1426,N_135,N_591);
or U1427 (N_1427,N_717,N_503);
or U1428 (N_1428,N_409,N_41);
or U1429 (N_1429,N_287,N_781);
nor U1430 (N_1430,N_696,N_476);
or U1431 (N_1431,N_416,N_997);
or U1432 (N_1432,N_712,N_700);
nor U1433 (N_1433,N_137,N_123);
nor U1434 (N_1434,N_441,N_165);
nor U1435 (N_1435,N_580,N_652);
or U1436 (N_1436,N_178,N_114);
and U1437 (N_1437,N_948,N_570);
and U1438 (N_1438,N_543,N_492);
nor U1439 (N_1439,N_474,N_308);
and U1440 (N_1440,N_103,N_37);
nand U1441 (N_1441,N_330,N_232);
nand U1442 (N_1442,N_234,N_215);
nor U1443 (N_1443,N_621,N_391);
nor U1444 (N_1444,N_707,N_694);
and U1445 (N_1445,N_728,N_914);
or U1446 (N_1446,N_518,N_231);
or U1447 (N_1447,N_75,N_622);
nand U1448 (N_1448,N_958,N_564);
nor U1449 (N_1449,N_344,N_269);
nor U1450 (N_1450,N_97,N_281);
and U1451 (N_1451,N_527,N_293);
nor U1452 (N_1452,N_433,N_954);
and U1453 (N_1453,N_594,N_685);
nand U1454 (N_1454,N_248,N_66);
nor U1455 (N_1455,N_236,N_314);
nor U1456 (N_1456,N_820,N_512);
nand U1457 (N_1457,N_569,N_500);
nor U1458 (N_1458,N_519,N_325);
and U1459 (N_1459,N_929,N_737);
and U1460 (N_1460,N_697,N_743);
and U1461 (N_1461,N_535,N_721);
or U1462 (N_1462,N_933,N_306);
and U1463 (N_1463,N_213,N_971);
nand U1464 (N_1464,N_150,N_517);
and U1465 (N_1465,N_821,N_359);
and U1466 (N_1466,N_641,N_337);
nand U1467 (N_1467,N_161,N_119);
nor U1468 (N_1468,N_976,N_207);
nor U1469 (N_1469,N_605,N_151);
nor U1470 (N_1470,N_340,N_730);
nand U1471 (N_1471,N_542,N_334);
nor U1472 (N_1472,N_683,N_528);
nor U1473 (N_1473,N_386,N_740);
nand U1474 (N_1474,N_763,N_577);
and U1475 (N_1475,N_303,N_726);
nand U1476 (N_1476,N_205,N_105);
and U1477 (N_1477,N_796,N_496);
nor U1478 (N_1478,N_159,N_484);
and U1479 (N_1479,N_722,N_36);
or U1480 (N_1480,N_988,N_673);
nand U1481 (N_1481,N_529,N_786);
nor U1482 (N_1482,N_385,N_396);
and U1483 (N_1483,N_472,N_140);
and U1484 (N_1484,N_423,N_630);
or U1485 (N_1485,N_129,N_98);
nor U1486 (N_1486,N_941,N_250);
nor U1487 (N_1487,N_469,N_130);
nor U1488 (N_1488,N_563,N_598);
and U1489 (N_1489,N_836,N_419);
and U1490 (N_1490,N_332,N_440);
and U1491 (N_1491,N_980,N_629);
nand U1492 (N_1492,N_295,N_724);
or U1493 (N_1493,N_394,N_680);
or U1494 (N_1494,N_882,N_851);
nand U1495 (N_1495,N_837,N_830);
or U1496 (N_1496,N_479,N_544);
nand U1497 (N_1497,N_892,N_946);
nand U1498 (N_1498,N_163,N_585);
nor U1499 (N_1499,N_262,N_175);
nor U1500 (N_1500,N_915,N_130);
and U1501 (N_1501,N_663,N_61);
or U1502 (N_1502,N_849,N_375);
nor U1503 (N_1503,N_604,N_927);
nor U1504 (N_1504,N_232,N_195);
and U1505 (N_1505,N_149,N_448);
and U1506 (N_1506,N_833,N_911);
or U1507 (N_1507,N_272,N_502);
or U1508 (N_1508,N_595,N_208);
nand U1509 (N_1509,N_178,N_331);
and U1510 (N_1510,N_276,N_728);
nand U1511 (N_1511,N_186,N_48);
nor U1512 (N_1512,N_476,N_868);
nand U1513 (N_1513,N_760,N_277);
or U1514 (N_1514,N_353,N_178);
nand U1515 (N_1515,N_872,N_26);
and U1516 (N_1516,N_367,N_169);
or U1517 (N_1517,N_61,N_412);
or U1518 (N_1518,N_467,N_937);
and U1519 (N_1519,N_741,N_360);
and U1520 (N_1520,N_545,N_436);
nand U1521 (N_1521,N_347,N_132);
nor U1522 (N_1522,N_398,N_688);
xnor U1523 (N_1523,N_870,N_169);
and U1524 (N_1524,N_193,N_472);
and U1525 (N_1525,N_827,N_820);
nand U1526 (N_1526,N_395,N_183);
or U1527 (N_1527,N_802,N_583);
nor U1528 (N_1528,N_3,N_277);
nand U1529 (N_1529,N_505,N_480);
and U1530 (N_1530,N_139,N_547);
and U1531 (N_1531,N_879,N_798);
nor U1532 (N_1532,N_537,N_245);
and U1533 (N_1533,N_185,N_546);
nand U1534 (N_1534,N_172,N_609);
nand U1535 (N_1535,N_763,N_195);
or U1536 (N_1536,N_610,N_17);
nand U1537 (N_1537,N_317,N_106);
or U1538 (N_1538,N_313,N_732);
or U1539 (N_1539,N_258,N_485);
and U1540 (N_1540,N_512,N_406);
nor U1541 (N_1541,N_645,N_962);
or U1542 (N_1542,N_283,N_52);
and U1543 (N_1543,N_320,N_815);
nor U1544 (N_1544,N_389,N_208);
or U1545 (N_1545,N_495,N_333);
and U1546 (N_1546,N_900,N_308);
nand U1547 (N_1547,N_443,N_823);
nor U1548 (N_1548,N_803,N_123);
xnor U1549 (N_1549,N_28,N_954);
nand U1550 (N_1550,N_726,N_162);
or U1551 (N_1551,N_200,N_120);
nor U1552 (N_1552,N_458,N_32);
and U1553 (N_1553,N_473,N_604);
and U1554 (N_1554,N_482,N_967);
nor U1555 (N_1555,N_387,N_769);
nor U1556 (N_1556,N_575,N_272);
nor U1557 (N_1557,N_211,N_319);
and U1558 (N_1558,N_992,N_598);
nand U1559 (N_1559,N_885,N_118);
and U1560 (N_1560,N_69,N_444);
and U1561 (N_1561,N_179,N_705);
and U1562 (N_1562,N_256,N_750);
nand U1563 (N_1563,N_406,N_601);
nor U1564 (N_1564,N_477,N_823);
or U1565 (N_1565,N_96,N_840);
nand U1566 (N_1566,N_577,N_278);
nor U1567 (N_1567,N_624,N_253);
nor U1568 (N_1568,N_669,N_48);
and U1569 (N_1569,N_91,N_679);
nand U1570 (N_1570,N_320,N_906);
and U1571 (N_1571,N_855,N_246);
and U1572 (N_1572,N_165,N_614);
and U1573 (N_1573,N_374,N_733);
nand U1574 (N_1574,N_784,N_772);
and U1575 (N_1575,N_934,N_353);
and U1576 (N_1576,N_673,N_55);
or U1577 (N_1577,N_299,N_772);
nand U1578 (N_1578,N_129,N_124);
nand U1579 (N_1579,N_523,N_351);
nand U1580 (N_1580,N_39,N_611);
or U1581 (N_1581,N_607,N_734);
nor U1582 (N_1582,N_357,N_260);
or U1583 (N_1583,N_865,N_338);
and U1584 (N_1584,N_314,N_938);
or U1585 (N_1585,N_711,N_579);
nand U1586 (N_1586,N_549,N_145);
or U1587 (N_1587,N_287,N_462);
nor U1588 (N_1588,N_840,N_374);
and U1589 (N_1589,N_486,N_579);
and U1590 (N_1590,N_461,N_201);
and U1591 (N_1591,N_356,N_880);
nand U1592 (N_1592,N_609,N_486);
nor U1593 (N_1593,N_778,N_674);
or U1594 (N_1594,N_514,N_449);
nor U1595 (N_1595,N_212,N_579);
and U1596 (N_1596,N_203,N_737);
or U1597 (N_1597,N_320,N_354);
nor U1598 (N_1598,N_655,N_705);
and U1599 (N_1599,N_283,N_688);
or U1600 (N_1600,N_777,N_601);
nor U1601 (N_1601,N_165,N_482);
nor U1602 (N_1602,N_933,N_651);
nor U1603 (N_1603,N_768,N_670);
and U1604 (N_1604,N_142,N_268);
or U1605 (N_1605,N_72,N_2);
and U1606 (N_1606,N_583,N_150);
nand U1607 (N_1607,N_920,N_858);
nand U1608 (N_1608,N_743,N_53);
nor U1609 (N_1609,N_158,N_200);
nand U1610 (N_1610,N_321,N_668);
or U1611 (N_1611,N_276,N_991);
or U1612 (N_1612,N_89,N_706);
and U1613 (N_1613,N_603,N_194);
and U1614 (N_1614,N_142,N_724);
and U1615 (N_1615,N_289,N_761);
nor U1616 (N_1616,N_419,N_867);
nand U1617 (N_1617,N_682,N_634);
or U1618 (N_1618,N_522,N_385);
and U1619 (N_1619,N_514,N_407);
xor U1620 (N_1620,N_441,N_704);
nand U1621 (N_1621,N_584,N_843);
nor U1622 (N_1622,N_242,N_923);
and U1623 (N_1623,N_429,N_385);
and U1624 (N_1624,N_272,N_683);
and U1625 (N_1625,N_764,N_497);
and U1626 (N_1626,N_164,N_401);
and U1627 (N_1627,N_225,N_128);
nand U1628 (N_1628,N_641,N_108);
nor U1629 (N_1629,N_913,N_104);
nand U1630 (N_1630,N_346,N_395);
nand U1631 (N_1631,N_750,N_589);
nand U1632 (N_1632,N_578,N_316);
or U1633 (N_1633,N_632,N_762);
nor U1634 (N_1634,N_29,N_747);
or U1635 (N_1635,N_370,N_56);
or U1636 (N_1636,N_567,N_299);
xor U1637 (N_1637,N_100,N_903);
xor U1638 (N_1638,N_902,N_521);
or U1639 (N_1639,N_652,N_683);
nor U1640 (N_1640,N_101,N_808);
nor U1641 (N_1641,N_486,N_599);
nand U1642 (N_1642,N_211,N_869);
nor U1643 (N_1643,N_52,N_39);
or U1644 (N_1644,N_511,N_207);
nand U1645 (N_1645,N_109,N_254);
or U1646 (N_1646,N_553,N_815);
or U1647 (N_1647,N_751,N_888);
nor U1648 (N_1648,N_548,N_883);
or U1649 (N_1649,N_447,N_630);
nand U1650 (N_1650,N_157,N_942);
nand U1651 (N_1651,N_575,N_535);
or U1652 (N_1652,N_734,N_294);
and U1653 (N_1653,N_586,N_474);
nand U1654 (N_1654,N_649,N_899);
nor U1655 (N_1655,N_283,N_37);
nor U1656 (N_1656,N_239,N_835);
and U1657 (N_1657,N_134,N_853);
nor U1658 (N_1658,N_691,N_595);
nor U1659 (N_1659,N_674,N_896);
and U1660 (N_1660,N_826,N_292);
and U1661 (N_1661,N_682,N_539);
or U1662 (N_1662,N_375,N_547);
or U1663 (N_1663,N_501,N_487);
nand U1664 (N_1664,N_837,N_399);
or U1665 (N_1665,N_697,N_467);
nand U1666 (N_1666,N_839,N_819);
nand U1667 (N_1667,N_195,N_703);
or U1668 (N_1668,N_239,N_219);
and U1669 (N_1669,N_134,N_367);
and U1670 (N_1670,N_802,N_861);
nor U1671 (N_1671,N_652,N_165);
nor U1672 (N_1672,N_885,N_577);
or U1673 (N_1673,N_196,N_413);
nor U1674 (N_1674,N_776,N_69);
nor U1675 (N_1675,N_760,N_912);
nand U1676 (N_1676,N_941,N_202);
nand U1677 (N_1677,N_206,N_784);
or U1678 (N_1678,N_285,N_193);
nand U1679 (N_1679,N_637,N_449);
and U1680 (N_1680,N_620,N_203);
nor U1681 (N_1681,N_419,N_369);
and U1682 (N_1682,N_47,N_277);
nand U1683 (N_1683,N_566,N_327);
nor U1684 (N_1684,N_27,N_963);
or U1685 (N_1685,N_856,N_927);
and U1686 (N_1686,N_268,N_716);
or U1687 (N_1687,N_641,N_359);
xor U1688 (N_1688,N_562,N_342);
or U1689 (N_1689,N_467,N_568);
or U1690 (N_1690,N_505,N_62);
and U1691 (N_1691,N_800,N_773);
and U1692 (N_1692,N_906,N_67);
nand U1693 (N_1693,N_654,N_995);
or U1694 (N_1694,N_609,N_952);
and U1695 (N_1695,N_592,N_137);
nand U1696 (N_1696,N_697,N_856);
nor U1697 (N_1697,N_454,N_712);
nand U1698 (N_1698,N_509,N_563);
nand U1699 (N_1699,N_289,N_903);
or U1700 (N_1700,N_396,N_838);
nor U1701 (N_1701,N_52,N_854);
nor U1702 (N_1702,N_255,N_868);
nand U1703 (N_1703,N_380,N_585);
nand U1704 (N_1704,N_687,N_951);
and U1705 (N_1705,N_561,N_877);
nor U1706 (N_1706,N_483,N_244);
or U1707 (N_1707,N_383,N_743);
nand U1708 (N_1708,N_135,N_666);
nor U1709 (N_1709,N_682,N_754);
and U1710 (N_1710,N_798,N_360);
nor U1711 (N_1711,N_21,N_792);
nand U1712 (N_1712,N_77,N_330);
and U1713 (N_1713,N_317,N_807);
and U1714 (N_1714,N_319,N_774);
and U1715 (N_1715,N_903,N_776);
nor U1716 (N_1716,N_114,N_332);
nand U1717 (N_1717,N_699,N_296);
nor U1718 (N_1718,N_387,N_243);
nand U1719 (N_1719,N_961,N_598);
and U1720 (N_1720,N_742,N_751);
nor U1721 (N_1721,N_70,N_56);
and U1722 (N_1722,N_35,N_388);
nand U1723 (N_1723,N_635,N_875);
nand U1724 (N_1724,N_566,N_535);
nand U1725 (N_1725,N_22,N_475);
or U1726 (N_1726,N_291,N_256);
nand U1727 (N_1727,N_640,N_797);
nor U1728 (N_1728,N_945,N_944);
or U1729 (N_1729,N_668,N_806);
nor U1730 (N_1730,N_863,N_688);
or U1731 (N_1731,N_314,N_569);
and U1732 (N_1732,N_553,N_254);
nor U1733 (N_1733,N_876,N_395);
and U1734 (N_1734,N_603,N_832);
and U1735 (N_1735,N_30,N_263);
and U1736 (N_1736,N_829,N_765);
nand U1737 (N_1737,N_80,N_613);
or U1738 (N_1738,N_41,N_701);
and U1739 (N_1739,N_534,N_995);
nor U1740 (N_1740,N_206,N_183);
xor U1741 (N_1741,N_327,N_163);
nor U1742 (N_1742,N_573,N_872);
and U1743 (N_1743,N_454,N_189);
and U1744 (N_1744,N_916,N_515);
nand U1745 (N_1745,N_63,N_204);
and U1746 (N_1746,N_596,N_790);
and U1747 (N_1747,N_500,N_873);
nor U1748 (N_1748,N_311,N_178);
or U1749 (N_1749,N_327,N_609);
nor U1750 (N_1750,N_530,N_215);
nor U1751 (N_1751,N_368,N_847);
and U1752 (N_1752,N_508,N_96);
xnor U1753 (N_1753,N_657,N_427);
nand U1754 (N_1754,N_172,N_322);
and U1755 (N_1755,N_418,N_137);
nand U1756 (N_1756,N_166,N_393);
or U1757 (N_1757,N_894,N_702);
and U1758 (N_1758,N_699,N_219);
or U1759 (N_1759,N_925,N_155);
or U1760 (N_1760,N_212,N_503);
and U1761 (N_1761,N_203,N_684);
or U1762 (N_1762,N_823,N_435);
or U1763 (N_1763,N_598,N_348);
or U1764 (N_1764,N_468,N_364);
nor U1765 (N_1765,N_411,N_88);
and U1766 (N_1766,N_334,N_39);
or U1767 (N_1767,N_61,N_241);
nor U1768 (N_1768,N_603,N_788);
or U1769 (N_1769,N_696,N_358);
or U1770 (N_1770,N_766,N_394);
or U1771 (N_1771,N_824,N_346);
nor U1772 (N_1772,N_498,N_391);
nor U1773 (N_1773,N_905,N_330);
nand U1774 (N_1774,N_770,N_385);
and U1775 (N_1775,N_936,N_413);
nor U1776 (N_1776,N_815,N_12);
and U1777 (N_1777,N_61,N_705);
and U1778 (N_1778,N_557,N_321);
xnor U1779 (N_1779,N_430,N_789);
nand U1780 (N_1780,N_52,N_152);
or U1781 (N_1781,N_765,N_367);
nor U1782 (N_1782,N_836,N_538);
xnor U1783 (N_1783,N_646,N_944);
or U1784 (N_1784,N_412,N_546);
nor U1785 (N_1785,N_617,N_16);
and U1786 (N_1786,N_378,N_66);
nand U1787 (N_1787,N_528,N_430);
or U1788 (N_1788,N_202,N_648);
xnor U1789 (N_1789,N_866,N_242);
nor U1790 (N_1790,N_355,N_927);
or U1791 (N_1791,N_981,N_907);
nor U1792 (N_1792,N_255,N_786);
nor U1793 (N_1793,N_530,N_948);
and U1794 (N_1794,N_917,N_327);
and U1795 (N_1795,N_827,N_186);
nor U1796 (N_1796,N_387,N_643);
nand U1797 (N_1797,N_25,N_27);
nor U1798 (N_1798,N_941,N_860);
and U1799 (N_1799,N_23,N_359);
nor U1800 (N_1800,N_945,N_712);
and U1801 (N_1801,N_98,N_81);
nand U1802 (N_1802,N_531,N_372);
and U1803 (N_1803,N_903,N_912);
and U1804 (N_1804,N_595,N_743);
or U1805 (N_1805,N_124,N_957);
and U1806 (N_1806,N_632,N_657);
nor U1807 (N_1807,N_317,N_704);
or U1808 (N_1808,N_432,N_10);
and U1809 (N_1809,N_692,N_839);
nor U1810 (N_1810,N_668,N_631);
nor U1811 (N_1811,N_73,N_509);
nand U1812 (N_1812,N_134,N_877);
or U1813 (N_1813,N_455,N_502);
nor U1814 (N_1814,N_977,N_550);
nor U1815 (N_1815,N_645,N_250);
or U1816 (N_1816,N_367,N_432);
and U1817 (N_1817,N_749,N_582);
nand U1818 (N_1818,N_907,N_780);
or U1819 (N_1819,N_742,N_100);
nand U1820 (N_1820,N_919,N_969);
nor U1821 (N_1821,N_697,N_313);
nand U1822 (N_1822,N_438,N_243);
or U1823 (N_1823,N_278,N_216);
or U1824 (N_1824,N_754,N_351);
nor U1825 (N_1825,N_98,N_384);
and U1826 (N_1826,N_798,N_577);
and U1827 (N_1827,N_145,N_148);
nand U1828 (N_1828,N_448,N_642);
nand U1829 (N_1829,N_78,N_74);
and U1830 (N_1830,N_375,N_649);
nand U1831 (N_1831,N_311,N_891);
or U1832 (N_1832,N_597,N_606);
nand U1833 (N_1833,N_42,N_896);
nand U1834 (N_1834,N_657,N_578);
and U1835 (N_1835,N_469,N_775);
nand U1836 (N_1836,N_748,N_449);
or U1837 (N_1837,N_48,N_123);
and U1838 (N_1838,N_820,N_280);
nor U1839 (N_1839,N_689,N_895);
nand U1840 (N_1840,N_65,N_875);
and U1841 (N_1841,N_744,N_997);
and U1842 (N_1842,N_767,N_94);
or U1843 (N_1843,N_562,N_907);
or U1844 (N_1844,N_285,N_602);
nand U1845 (N_1845,N_192,N_791);
nor U1846 (N_1846,N_767,N_83);
nand U1847 (N_1847,N_472,N_744);
and U1848 (N_1848,N_23,N_951);
nand U1849 (N_1849,N_923,N_857);
nor U1850 (N_1850,N_658,N_464);
nand U1851 (N_1851,N_296,N_20);
nand U1852 (N_1852,N_505,N_974);
nor U1853 (N_1853,N_834,N_911);
nor U1854 (N_1854,N_225,N_77);
and U1855 (N_1855,N_714,N_392);
or U1856 (N_1856,N_907,N_320);
nand U1857 (N_1857,N_16,N_553);
or U1858 (N_1858,N_898,N_971);
nor U1859 (N_1859,N_456,N_671);
nand U1860 (N_1860,N_580,N_687);
nor U1861 (N_1861,N_628,N_392);
nand U1862 (N_1862,N_427,N_455);
or U1863 (N_1863,N_650,N_335);
and U1864 (N_1864,N_19,N_749);
or U1865 (N_1865,N_455,N_679);
and U1866 (N_1866,N_850,N_846);
nand U1867 (N_1867,N_120,N_32);
nor U1868 (N_1868,N_377,N_27);
or U1869 (N_1869,N_746,N_27);
or U1870 (N_1870,N_881,N_304);
nor U1871 (N_1871,N_346,N_804);
or U1872 (N_1872,N_699,N_232);
nand U1873 (N_1873,N_531,N_705);
or U1874 (N_1874,N_120,N_607);
and U1875 (N_1875,N_55,N_272);
nand U1876 (N_1876,N_56,N_787);
or U1877 (N_1877,N_339,N_48);
nor U1878 (N_1878,N_586,N_976);
and U1879 (N_1879,N_248,N_204);
or U1880 (N_1880,N_551,N_378);
or U1881 (N_1881,N_118,N_911);
nor U1882 (N_1882,N_852,N_530);
or U1883 (N_1883,N_395,N_391);
nand U1884 (N_1884,N_128,N_568);
and U1885 (N_1885,N_762,N_682);
or U1886 (N_1886,N_474,N_221);
nor U1887 (N_1887,N_509,N_663);
and U1888 (N_1888,N_132,N_958);
or U1889 (N_1889,N_70,N_986);
or U1890 (N_1890,N_699,N_21);
or U1891 (N_1891,N_629,N_242);
or U1892 (N_1892,N_350,N_339);
nor U1893 (N_1893,N_208,N_51);
or U1894 (N_1894,N_149,N_669);
and U1895 (N_1895,N_781,N_627);
nor U1896 (N_1896,N_13,N_708);
and U1897 (N_1897,N_113,N_628);
and U1898 (N_1898,N_509,N_158);
or U1899 (N_1899,N_679,N_117);
and U1900 (N_1900,N_761,N_363);
or U1901 (N_1901,N_977,N_309);
and U1902 (N_1902,N_514,N_785);
nand U1903 (N_1903,N_522,N_330);
or U1904 (N_1904,N_320,N_382);
nand U1905 (N_1905,N_692,N_949);
and U1906 (N_1906,N_878,N_352);
or U1907 (N_1907,N_547,N_897);
nor U1908 (N_1908,N_206,N_53);
and U1909 (N_1909,N_496,N_479);
nand U1910 (N_1910,N_234,N_718);
nor U1911 (N_1911,N_227,N_626);
and U1912 (N_1912,N_51,N_717);
or U1913 (N_1913,N_239,N_185);
nand U1914 (N_1914,N_601,N_757);
or U1915 (N_1915,N_947,N_985);
nor U1916 (N_1916,N_780,N_906);
nor U1917 (N_1917,N_928,N_508);
nand U1918 (N_1918,N_500,N_392);
or U1919 (N_1919,N_590,N_480);
or U1920 (N_1920,N_932,N_973);
or U1921 (N_1921,N_520,N_785);
and U1922 (N_1922,N_343,N_37);
nand U1923 (N_1923,N_28,N_607);
nor U1924 (N_1924,N_244,N_475);
nand U1925 (N_1925,N_153,N_388);
or U1926 (N_1926,N_879,N_736);
nor U1927 (N_1927,N_46,N_317);
or U1928 (N_1928,N_689,N_863);
nor U1929 (N_1929,N_234,N_787);
or U1930 (N_1930,N_893,N_758);
and U1931 (N_1931,N_116,N_418);
nand U1932 (N_1932,N_182,N_507);
xor U1933 (N_1933,N_559,N_134);
nand U1934 (N_1934,N_785,N_699);
nand U1935 (N_1935,N_556,N_674);
nor U1936 (N_1936,N_846,N_868);
or U1937 (N_1937,N_890,N_813);
or U1938 (N_1938,N_757,N_120);
nand U1939 (N_1939,N_162,N_200);
nand U1940 (N_1940,N_720,N_106);
nand U1941 (N_1941,N_485,N_275);
or U1942 (N_1942,N_998,N_379);
nand U1943 (N_1943,N_840,N_639);
or U1944 (N_1944,N_241,N_110);
or U1945 (N_1945,N_485,N_858);
nor U1946 (N_1946,N_967,N_90);
nor U1947 (N_1947,N_947,N_329);
nor U1948 (N_1948,N_719,N_842);
or U1949 (N_1949,N_163,N_246);
or U1950 (N_1950,N_205,N_186);
nor U1951 (N_1951,N_295,N_831);
and U1952 (N_1952,N_876,N_388);
nor U1953 (N_1953,N_588,N_961);
and U1954 (N_1954,N_560,N_928);
nor U1955 (N_1955,N_603,N_707);
nand U1956 (N_1956,N_977,N_530);
nand U1957 (N_1957,N_594,N_412);
nor U1958 (N_1958,N_295,N_914);
or U1959 (N_1959,N_766,N_52);
or U1960 (N_1960,N_610,N_979);
or U1961 (N_1961,N_826,N_362);
or U1962 (N_1962,N_995,N_748);
and U1963 (N_1963,N_469,N_339);
nor U1964 (N_1964,N_599,N_616);
or U1965 (N_1965,N_797,N_292);
or U1966 (N_1966,N_725,N_534);
or U1967 (N_1967,N_376,N_926);
nand U1968 (N_1968,N_8,N_703);
and U1969 (N_1969,N_108,N_544);
nor U1970 (N_1970,N_263,N_13);
or U1971 (N_1971,N_362,N_99);
or U1972 (N_1972,N_546,N_100);
or U1973 (N_1973,N_295,N_141);
nor U1974 (N_1974,N_96,N_744);
nand U1975 (N_1975,N_519,N_380);
nor U1976 (N_1976,N_676,N_698);
nand U1977 (N_1977,N_552,N_156);
nor U1978 (N_1978,N_936,N_571);
nand U1979 (N_1979,N_92,N_157);
and U1980 (N_1980,N_877,N_871);
or U1981 (N_1981,N_879,N_584);
nor U1982 (N_1982,N_408,N_247);
nand U1983 (N_1983,N_691,N_401);
xor U1984 (N_1984,N_625,N_1);
and U1985 (N_1985,N_251,N_991);
nor U1986 (N_1986,N_380,N_118);
or U1987 (N_1987,N_127,N_986);
or U1988 (N_1988,N_379,N_475);
and U1989 (N_1989,N_924,N_469);
nor U1990 (N_1990,N_713,N_914);
or U1991 (N_1991,N_781,N_161);
nor U1992 (N_1992,N_703,N_682);
and U1993 (N_1993,N_956,N_922);
nor U1994 (N_1994,N_846,N_702);
and U1995 (N_1995,N_989,N_618);
nand U1996 (N_1996,N_65,N_693);
or U1997 (N_1997,N_564,N_683);
nand U1998 (N_1998,N_486,N_21);
or U1999 (N_1999,N_736,N_691);
nor U2000 (N_2000,N_1118,N_1756);
and U2001 (N_2001,N_1899,N_1987);
nand U2002 (N_2002,N_1026,N_1128);
nand U2003 (N_2003,N_1690,N_1373);
and U2004 (N_2004,N_1417,N_1673);
nor U2005 (N_2005,N_1038,N_1172);
and U2006 (N_2006,N_1149,N_1372);
and U2007 (N_2007,N_1667,N_1918);
or U2008 (N_2008,N_1312,N_1794);
or U2009 (N_2009,N_1743,N_1747);
nand U2010 (N_2010,N_1279,N_1754);
nor U2011 (N_2011,N_1330,N_1167);
nand U2012 (N_2012,N_1993,N_1805);
and U2013 (N_2013,N_1711,N_1979);
or U2014 (N_2014,N_1737,N_1908);
or U2015 (N_2015,N_1543,N_1764);
nand U2016 (N_2016,N_1284,N_1553);
nor U2017 (N_2017,N_1657,N_1988);
nor U2018 (N_2018,N_1045,N_1307);
or U2019 (N_2019,N_1071,N_1566);
and U2020 (N_2020,N_1051,N_1913);
or U2021 (N_2021,N_1075,N_1391);
and U2022 (N_2022,N_1871,N_1792);
nor U2023 (N_2023,N_1121,N_1145);
nand U2024 (N_2024,N_1019,N_1466);
and U2025 (N_2025,N_1403,N_1724);
nand U2026 (N_2026,N_1322,N_1855);
nand U2027 (N_2027,N_1893,N_1483);
xor U2028 (N_2028,N_1909,N_1056);
nand U2029 (N_2029,N_1895,N_1361);
and U2030 (N_2030,N_1206,N_1867);
nor U2031 (N_2031,N_1286,N_1348);
nor U2032 (N_2032,N_1544,N_1649);
and U2033 (N_2033,N_1992,N_1691);
nand U2034 (N_2034,N_1961,N_1059);
nor U2035 (N_2035,N_1161,N_1933);
nand U2036 (N_2036,N_1249,N_1827);
nor U2037 (N_2037,N_1437,N_1453);
or U2038 (N_2038,N_1624,N_1584);
nor U2039 (N_2039,N_1801,N_1050);
and U2040 (N_2040,N_1707,N_1920);
and U2041 (N_2041,N_1628,N_1213);
and U2042 (N_2042,N_1314,N_1105);
or U2043 (N_2043,N_1454,N_1469);
or U2044 (N_2044,N_1804,N_1795);
and U2045 (N_2045,N_1338,N_1672);
and U2046 (N_2046,N_1491,N_1100);
or U2047 (N_2047,N_1418,N_1364);
nand U2048 (N_2048,N_1263,N_1168);
nor U2049 (N_2049,N_1502,N_1040);
nor U2050 (N_2050,N_1571,N_1254);
and U2051 (N_2051,N_1677,N_1549);
and U2052 (N_2052,N_1822,N_1237);
nor U2053 (N_2053,N_1610,N_1209);
nor U2054 (N_2054,N_1425,N_1394);
nor U2055 (N_2055,N_1715,N_1116);
nor U2056 (N_2056,N_1255,N_1024);
nand U2057 (N_2057,N_1017,N_1450);
or U2058 (N_2058,N_1346,N_1052);
nor U2059 (N_2059,N_1999,N_1949);
nand U2060 (N_2060,N_1318,N_1305);
or U2061 (N_2061,N_1151,N_1402);
and U2062 (N_2062,N_1477,N_1938);
or U2063 (N_2063,N_1400,N_1865);
and U2064 (N_2064,N_1309,N_1496);
xnor U2065 (N_2065,N_1319,N_1081);
or U2066 (N_2066,N_1212,N_1970);
or U2067 (N_2067,N_1775,N_1660);
nand U2068 (N_2068,N_1223,N_1790);
and U2069 (N_2069,N_1759,N_1746);
or U2070 (N_2070,N_1510,N_1587);
or U2071 (N_2071,N_1296,N_1260);
nor U2072 (N_2072,N_1273,N_1640);
or U2073 (N_2073,N_1383,N_1839);
or U2074 (N_2074,N_1902,N_1655);
nand U2075 (N_2075,N_1718,N_1749);
or U2076 (N_2076,N_1973,N_1243);
or U2077 (N_2077,N_1604,N_1879);
or U2078 (N_2078,N_1097,N_1262);
and U2079 (N_2079,N_1456,N_1658);
nand U2080 (N_2080,N_1609,N_1041);
nand U2081 (N_2081,N_1726,N_1411);
nor U2082 (N_2082,N_1981,N_1951);
nor U2083 (N_2083,N_1798,N_1803);
nor U2084 (N_2084,N_1634,N_1295);
and U2085 (N_2085,N_1144,N_1773);
and U2086 (N_2086,N_1107,N_1004);
and U2087 (N_2087,N_1449,N_1680);
nor U2088 (N_2088,N_1072,N_1969);
and U2089 (N_2089,N_1165,N_1397);
nand U2090 (N_2090,N_1520,N_1872);
and U2091 (N_2091,N_1304,N_1084);
nand U2092 (N_2092,N_1245,N_1122);
nand U2093 (N_2093,N_1142,N_1717);
and U2094 (N_2094,N_1772,N_1113);
or U2095 (N_2095,N_1635,N_1952);
and U2096 (N_2096,N_1575,N_1321);
and U2097 (N_2097,N_1174,N_1217);
nor U2098 (N_2098,N_1336,N_1170);
xor U2099 (N_2099,N_1214,N_1508);
or U2100 (N_2100,N_1340,N_1796);
and U2101 (N_2101,N_1222,N_1617);
or U2102 (N_2102,N_1415,N_1405);
and U2103 (N_2103,N_1028,N_1110);
or U2104 (N_2104,N_1499,N_1712);
nor U2105 (N_2105,N_1727,N_1386);
nor U2106 (N_2106,N_1016,N_1457);
and U2107 (N_2107,N_1080,N_1581);
or U2108 (N_2108,N_1461,N_1079);
or U2109 (N_2109,N_1830,N_1375);
nand U2110 (N_2110,N_1009,N_1602);
and U2111 (N_2111,N_1007,N_1094);
and U2112 (N_2112,N_1720,N_1897);
nor U2113 (N_2113,N_1676,N_1941);
nor U2114 (N_2114,N_1384,N_1064);
nand U2115 (N_2115,N_1177,N_1152);
and U2116 (N_2116,N_1848,N_1432);
and U2117 (N_2117,N_1275,N_1408);
or U2118 (N_2118,N_1721,N_1476);
nor U2119 (N_2119,N_1641,N_1387);
nand U2120 (N_2120,N_1367,N_1236);
xor U2121 (N_2121,N_1991,N_1083);
nor U2122 (N_2122,N_1734,N_1960);
and U2123 (N_2123,N_1027,N_1687);
or U2124 (N_2124,N_1115,N_1579);
and U2125 (N_2125,N_1374,N_1250);
or U2126 (N_2126,N_1333,N_1003);
and U2127 (N_2127,N_1272,N_1732);
and U2128 (N_2128,N_1120,N_1376);
nand U2129 (N_2129,N_1215,N_1911);
and U2130 (N_2130,N_1967,N_1932);
or U2131 (N_2131,N_1274,N_1129);
and U2132 (N_2132,N_1102,N_1328);
nor U2133 (N_2133,N_1576,N_1613);
or U2134 (N_2134,N_1661,N_1430);
and U2135 (N_2135,N_1465,N_1564);
or U2136 (N_2136,N_1958,N_1092);
nand U2137 (N_2137,N_1204,N_1504);
and U2138 (N_2138,N_1946,N_1585);
or U2139 (N_2139,N_1751,N_1123);
nor U2140 (N_2140,N_1696,N_1515);
and U2141 (N_2141,N_1234,N_1820);
nor U2142 (N_2142,N_1533,N_1605);
or U2143 (N_2143,N_1621,N_1183);
nand U2144 (N_2144,N_1968,N_1345);
and U2145 (N_2145,N_1745,N_1020);
and U2146 (N_2146,N_1664,N_1414);
and U2147 (N_2147,N_1875,N_1195);
and U2148 (N_2148,N_1114,N_1870);
nand U2149 (N_2149,N_1627,N_1943);
or U2150 (N_2150,N_1399,N_1324);
nor U2151 (N_2151,N_1208,N_1423);
nand U2152 (N_2152,N_1448,N_1668);
nor U2153 (N_2153,N_1767,N_1440);
or U2154 (N_2154,N_1599,N_1833);
nand U2155 (N_2155,N_1269,N_1265);
or U2156 (N_2156,N_1555,N_1858);
and U2157 (N_2157,N_1244,N_1828);
or U2158 (N_2158,N_1002,N_1488);
nand U2159 (N_2159,N_1252,N_1140);
nor U2160 (N_2160,N_1686,N_1860);
nand U2161 (N_2161,N_1439,N_1436);
or U2162 (N_2162,N_1203,N_1445);
nor U2163 (N_2163,N_1906,N_1021);
or U2164 (N_2164,N_1847,N_1280);
and U2165 (N_2165,N_1401,N_1350);
nor U2166 (N_2166,N_1138,N_1577);
or U2167 (N_2167,N_1153,N_1843);
nor U2168 (N_2168,N_1886,N_1482);
nor U2169 (N_2169,N_1331,N_1070);
nor U2170 (N_2170,N_1342,N_1154);
or U2171 (N_2171,N_1451,N_1662);
or U2172 (N_2172,N_1950,N_1963);
nand U2173 (N_2173,N_1325,N_1352);
and U2174 (N_2174,N_1065,N_1823);
nand U2175 (N_2175,N_1486,N_1939);
and U2176 (N_2176,N_1228,N_1306);
and U2177 (N_2177,N_1651,N_1883);
nand U2178 (N_2178,N_1853,N_1166);
or U2179 (N_2179,N_1537,N_1251);
and U2180 (N_2180,N_1890,N_1347);
nand U2181 (N_2181,N_1173,N_1701);
nor U2182 (N_2182,N_1196,N_1479);
nor U2183 (N_2183,N_1904,N_1859);
and U2184 (N_2184,N_1903,N_1665);
nand U2185 (N_2185,N_1888,N_1066);
nand U2186 (N_2186,N_1956,N_1355);
nand U2187 (N_2187,N_1616,N_1485);
and U2188 (N_2188,N_1467,N_1229);
or U2189 (N_2189,N_1238,N_1689);
nor U2190 (N_2190,N_1735,N_1516);
and U2191 (N_2191,N_1971,N_1335);
or U2192 (N_2192,N_1629,N_1039);
nand U2193 (N_2193,N_1901,N_1877);
nand U2194 (N_2194,N_1339,N_1940);
or U2195 (N_2195,N_1219,N_1438);
and U2196 (N_2196,N_1512,N_1791);
nand U2197 (N_2197,N_1876,N_1099);
or U2198 (N_2198,N_1054,N_1766);
or U2199 (N_2199,N_1974,N_1527);
and U2200 (N_2200,N_1101,N_1648);
nand U2201 (N_2201,N_1817,N_1601);
nand U2202 (N_2202,N_1567,N_1679);
nor U2203 (N_2203,N_1313,N_1193);
nor U2204 (N_2204,N_1854,N_1589);
nor U2205 (N_2205,N_1595,N_1380);
and U2206 (N_2206,N_1921,N_1618);
nand U2207 (N_2207,N_1211,N_1731);
nor U2208 (N_2208,N_1954,N_1704);
nor U2209 (N_2209,N_1643,N_1106);
or U2210 (N_2210,N_1659,N_1714);
and U2211 (N_2211,N_1344,N_1022);
and U2212 (N_2212,N_1639,N_1710);
nor U2213 (N_2213,N_1093,N_1620);
nand U2214 (N_2214,N_1137,N_1750);
nor U2215 (N_2215,N_1568,N_1010);
nor U2216 (N_2216,N_1558,N_1239);
or U2217 (N_2217,N_1363,N_1055);
nand U2218 (N_2218,N_1044,N_1852);
nand U2219 (N_2219,N_1034,N_1936);
nor U2220 (N_2220,N_1670,N_1594);
nor U2221 (N_2221,N_1163,N_1242);
nor U2222 (N_2222,N_1422,N_1266);
and U2223 (N_2223,N_1884,N_1836);
and U2224 (N_2224,N_1135,N_1300);
and U2225 (N_2225,N_1557,N_1642);
and U2226 (N_2226,N_1320,N_1162);
nor U2227 (N_2227,N_1914,N_1907);
nor U2228 (N_2228,N_1126,N_1753);
or U2229 (N_2229,N_1569,N_1292);
and U2230 (N_2230,N_1089,N_1261);
and U2231 (N_2231,N_1542,N_1600);
nor U2232 (N_2232,N_1232,N_1849);
or U2233 (N_2233,N_1471,N_1316);
nor U2234 (N_2234,N_1755,N_1287);
and U2235 (N_2235,N_1785,N_1591);
or U2236 (N_2236,N_1258,N_1741);
or U2237 (N_2237,N_1521,N_1518);
nor U2238 (N_2238,N_1646,N_1574);
nand U2239 (N_2239,N_1838,N_1233);
nand U2240 (N_2240,N_1290,N_1141);
and U2241 (N_2241,N_1861,N_1562);
and U2242 (N_2242,N_1636,N_1580);
or U2243 (N_2243,N_1277,N_1494);
or U2244 (N_2244,N_1606,N_1014);
or U2245 (N_2245,N_1930,N_1484);
nor U2246 (N_2246,N_1674,N_1500);
nor U2247 (N_2247,N_1783,N_1682);
nand U2248 (N_2248,N_1117,N_1788);
nor U2249 (N_2249,N_1612,N_1150);
nor U2250 (N_2250,N_1087,N_1001);
or U2251 (N_2251,N_1986,N_1736);
and U2252 (N_2252,N_1559,N_1507);
and U2253 (N_2253,N_1841,N_1327);
and U2254 (N_2254,N_1011,N_1942);
nor U2255 (N_2255,N_1199,N_1104);
and U2256 (N_2256,N_1545,N_1497);
nand U2257 (N_2257,N_1288,N_1389);
nor U2258 (N_2258,N_1271,N_1898);
or U2259 (N_2259,N_1308,N_1810);
and U2260 (N_2260,N_1207,N_1326);
or U2261 (N_2261,N_1431,N_1495);
nor U2262 (N_2262,N_1959,N_1663);
nand U2263 (N_2263,N_1998,N_1057);
and U2264 (N_2264,N_1377,N_1966);
nor U2265 (N_2265,N_1529,N_1480);
nor U2266 (N_2266,N_1124,N_1030);
or U2267 (N_2267,N_1758,N_1354);
and U2268 (N_2268,N_1873,N_1298);
nand U2269 (N_2269,N_1846,N_1937);
nor U2270 (N_2270,N_1807,N_1637);
or U2271 (N_2271,N_1825,N_1538);
xor U2272 (N_2272,N_1536,N_1460);
and U2273 (N_2273,N_1722,N_1977);
nand U2274 (N_2274,N_1370,N_1656);
nand U2275 (N_2275,N_1511,N_1996);
nand U2276 (N_2276,N_1230,N_1257);
and U2277 (N_2277,N_1994,N_1808);
and U2278 (N_2278,N_1005,N_1623);
nand U2279 (N_2279,N_1730,N_1984);
or U2280 (N_2280,N_1813,N_1225);
and U2281 (N_2281,N_1334,N_1443);
and U2282 (N_2282,N_1427,N_1832);
xor U2283 (N_2283,N_1688,N_1851);
nand U2284 (N_2284,N_1844,N_1492);
and U2285 (N_2285,N_1834,N_1698);
and U2286 (N_2286,N_1410,N_1935);
or U2287 (N_2287,N_1200,N_1761);
nor U2288 (N_2288,N_1894,N_1561);
or U2289 (N_2289,N_1353,N_1519);
nand U2290 (N_2290,N_1980,N_1548);
nand U2291 (N_2291,N_1366,N_1159);
nor U2292 (N_2292,N_1713,N_1915);
and U2293 (N_2293,N_1112,N_1428);
or U2294 (N_2294,N_1925,N_1446);
or U2295 (N_2295,N_1419,N_1098);
or U2296 (N_2296,N_1535,N_1809);
and U2297 (N_2297,N_1311,N_1806);
nor U2298 (N_2298,N_1652,N_1990);
nor U2299 (N_2299,N_1146,N_1725);
nand U2300 (N_2300,N_1824,N_1390);
nand U2301 (N_2301,N_1085,N_1171);
nand U2302 (N_2302,N_1835,N_1708);
nand U2303 (N_2303,N_1259,N_1205);
nor U2304 (N_2304,N_1184,N_1046);
and U2305 (N_2305,N_1049,N_1404);
nor U2306 (N_2306,N_1771,N_1797);
nor U2307 (N_2307,N_1995,N_1076);
nand U2308 (N_2308,N_1095,N_1799);
and U2309 (N_2309,N_1882,N_1845);
nor U2310 (N_2310,N_1033,N_1444);
and U2311 (N_2311,N_1692,N_1393);
nor U2312 (N_2312,N_1119,N_1694);
and U2313 (N_2313,N_1916,N_1596);
or U2314 (N_2314,N_1025,N_1365);
and U2315 (N_2315,N_1442,N_1435);
or U2316 (N_2316,N_1955,N_1493);
or U2317 (N_2317,N_1945,N_1647);
or U2318 (N_2318,N_1829,N_1187);
nor U2319 (N_2319,N_1598,N_1297);
or U2320 (N_2320,N_1189,N_1246);
nor U2321 (N_2321,N_1294,N_1550);
nor U2322 (N_2322,N_1359,N_1744);
and U2323 (N_2323,N_1586,N_1774);
nor U2324 (N_2324,N_1819,N_1474);
or U2325 (N_2325,N_1776,N_1818);
nand U2326 (N_2326,N_1626,N_1551);
and U2327 (N_2327,N_1175,N_1654);
nor U2328 (N_2328,N_1748,N_1927);
nand U2329 (N_2329,N_1198,N_1323);
xnor U2330 (N_2330,N_1880,N_1638);
or U2331 (N_2331,N_1928,N_1302);
or U2332 (N_2332,N_1392,N_1015);
or U2333 (N_2333,N_1289,N_1369);
nand U2334 (N_2334,N_1139,N_1702);
or U2335 (N_2335,N_1815,N_1357);
and U2336 (N_2336,N_1248,N_1891);
nand U2337 (N_2337,N_1912,N_1910);
nor U2338 (N_2338,N_1455,N_1784);
nor U2339 (N_2339,N_1088,N_1190);
nand U2340 (N_2340,N_1887,N_1630);
and U2341 (N_2341,N_1892,N_1182);
and U2342 (N_2342,N_1681,N_1191);
nor U2343 (N_2343,N_1247,N_1765);
nand U2344 (N_2344,N_1957,N_1625);
nor U2345 (N_2345,N_1475,N_1343);
nand U2346 (N_2346,N_1573,N_1157);
nand U2347 (N_2347,N_1517,N_1420);
and U2348 (N_2348,N_1278,N_1043);
nand U2349 (N_2349,N_1762,N_1134);
xor U2350 (N_2350,N_1133,N_1434);
nand U2351 (N_2351,N_1757,N_1096);
nor U2352 (N_2352,N_1983,N_1513);
nand U2353 (N_2353,N_1220,N_1006);
nand U2354 (N_2354,N_1351,N_1090);
and U2355 (N_2355,N_1077,N_1814);
and U2356 (N_2356,N_1035,N_1224);
nand U2357 (N_2357,N_1180,N_1752);
nor U2358 (N_2358,N_1881,N_1685);
and U2359 (N_2359,N_1074,N_1256);
and U2360 (N_2360,N_1866,N_1768);
nor U2361 (N_2361,N_1082,N_1885);
and U2362 (N_2362,N_1831,N_1179);
nor U2363 (N_2363,N_1395,N_1644);
nor U2364 (N_2364,N_1723,N_1862);
nand U2365 (N_2365,N_1147,N_1036);
and U2366 (N_2366,N_1560,N_1413);
or U2367 (N_2367,N_1127,N_1282);
nor U2368 (N_2368,N_1086,N_1675);
nor U2369 (N_2369,N_1706,N_1315);
xor U2370 (N_2370,N_1109,N_1058);
nor U2371 (N_2371,N_1053,N_1582);
or U2372 (N_2372,N_1607,N_1490);
or U2373 (N_2373,N_1412,N_1965);
nand U2374 (N_2374,N_1683,N_1012);
nor U2375 (N_2375,N_1148,N_1802);
nor U2376 (N_2376,N_1032,N_1962);
nor U2377 (N_2377,N_1556,N_1632);
nand U2378 (N_2378,N_1498,N_1650);
or U2379 (N_2379,N_1565,N_1760);
or U2380 (N_2380,N_1023,N_1285);
nand U2381 (N_2381,N_1793,N_1976);
nor U2382 (N_2382,N_1889,N_1633);
or U2383 (N_2383,N_1763,N_1329);
nand U2384 (N_2384,N_1132,N_1522);
nand U2385 (N_2385,N_1666,N_1473);
and U2386 (N_2386,N_1864,N_1780);
and U2387 (N_2387,N_1944,N_1381);
or U2388 (N_2388,N_1464,N_1964);
and U2389 (N_2389,N_1530,N_1164);
or U2390 (N_2390,N_1356,N_1563);
nand U2391 (N_2391,N_1441,N_1593);
and U2392 (N_2392,N_1406,N_1917);
and U2393 (N_2393,N_1842,N_1878);
and U2394 (N_2394,N_1900,N_1358);
nor U2395 (N_2395,N_1188,N_1934);
and U2396 (N_2396,N_1856,N_1197);
nor U2397 (N_2397,N_1291,N_1777);
or U2398 (N_2398,N_1919,N_1421);
nor U2399 (N_2399,N_1201,N_1705);
nand U2400 (N_2400,N_1018,N_1470);
nor U2401 (N_2401,N_1905,N_1501);
xor U2402 (N_2402,N_1837,N_1067);
or U2403 (N_2403,N_1826,N_1953);
and U2404 (N_2404,N_1235,N_1332);
nand U2405 (N_2405,N_1653,N_1534);
and U2406 (N_2406,N_1210,N_1409);
nand U2407 (N_2407,N_1740,N_1130);
and U2408 (N_2408,N_1226,N_1787);
nor U2409 (N_2409,N_1037,N_1989);
and U2410 (N_2410,N_1293,N_1281);
nand U2411 (N_2411,N_1812,N_1985);
nand U2412 (N_2412,N_1216,N_1301);
nand U2413 (N_2413,N_1253,N_1947);
nand U2414 (N_2414,N_1669,N_1388);
nor U2415 (N_2415,N_1742,N_1531);
or U2416 (N_2416,N_1136,N_1013);
nor U2417 (N_2417,N_1310,N_1231);
nand U2418 (N_2418,N_1462,N_1614);
nor U2419 (N_2419,N_1608,N_1382);
nand U2420 (N_2420,N_1779,N_1433);
or U2421 (N_2421,N_1398,N_1769);
nand U2422 (N_2422,N_1948,N_1506);
nor U2423 (N_2423,N_1029,N_1111);
and U2424 (N_2424,N_1221,N_1489);
nor U2425 (N_2425,N_1816,N_1671);
or U2426 (N_2426,N_1181,N_1583);
and U2427 (N_2427,N_1341,N_1202);
nand U2428 (N_2428,N_1929,N_1592);
and U2429 (N_2429,N_1103,N_1570);
and U2430 (N_2430,N_1611,N_1997);
and U2431 (N_2431,N_1061,N_1972);
or U2432 (N_2432,N_1468,N_1487);
and U2433 (N_2433,N_1378,N_1267);
nand U2434 (N_2434,N_1385,N_1709);
or U2435 (N_2435,N_1982,N_1588);
nor U2436 (N_2436,N_1268,N_1176);
and U2437 (N_2437,N_1227,N_1424);
or U2438 (N_2438,N_1552,N_1108);
and U2439 (N_2439,N_1684,N_1695);
nand U2440 (N_2440,N_1458,N_1619);
and U2441 (N_2441,N_1526,N_1240);
and U2442 (N_2442,N_1185,N_1615);
and U2443 (N_2443,N_1459,N_1603);
and U2444 (N_2444,N_1811,N_1194);
or U2445 (N_2445,N_1699,N_1703);
and U2446 (N_2446,N_1218,N_1645);
and U2447 (N_2447,N_1368,N_1078);
and U2448 (N_2448,N_1697,N_1733);
nand U2449 (N_2449,N_1523,N_1371);
nand U2450 (N_2450,N_1091,N_1738);
and U2451 (N_2451,N_1192,N_1868);
and U2452 (N_2452,N_1186,N_1360);
and U2453 (N_2453,N_1975,N_1155);
nor U2454 (N_2454,N_1008,N_1525);
nor U2455 (N_2455,N_1800,N_1283);
nor U2456 (N_2456,N_1063,N_1728);
nand U2457 (N_2457,N_1048,N_1156);
and U2458 (N_2458,N_1540,N_1396);
nand U2459 (N_2459,N_1869,N_1317);
nor U2460 (N_2460,N_1578,N_1926);
nor U2461 (N_2461,N_1276,N_1426);
and U2462 (N_2462,N_1923,N_1739);
and U2463 (N_2463,N_1524,N_1539);
or U2464 (N_2464,N_1060,N_1478);
nand U2465 (N_2465,N_1069,N_1857);
and U2466 (N_2466,N_1622,N_1874);
nor U2467 (N_2467,N_1678,N_1782);
or U2468 (N_2468,N_1590,N_1447);
nand U2469 (N_2469,N_1178,N_1978);
nor U2470 (N_2470,N_1031,N_1264);
nor U2471 (N_2471,N_1716,N_1693);
or U2472 (N_2472,N_1700,N_1509);
nand U2473 (N_2473,N_1481,N_1532);
and U2474 (N_2474,N_1472,N_1546);
or U2475 (N_2475,N_1299,N_1160);
nor U2476 (N_2476,N_1407,N_1597);
nand U2477 (N_2477,N_1778,N_1789);
or U2478 (N_2478,N_1303,N_1047);
or U2479 (N_2479,N_1541,N_1131);
or U2480 (N_2480,N_1514,N_1631);
nand U2481 (N_2481,N_1781,N_1379);
nand U2482 (N_2482,N_1850,N_1042);
or U2483 (N_2483,N_1924,N_1840);
or U2484 (N_2484,N_1062,N_1241);
nand U2485 (N_2485,N_1429,N_1547);
and U2486 (N_2486,N_1922,N_1073);
nor U2487 (N_2487,N_1863,N_1143);
or U2488 (N_2488,N_1896,N_1000);
or U2489 (N_2489,N_1270,N_1169);
nor U2490 (N_2490,N_1505,N_1125);
or U2491 (N_2491,N_1068,N_1416);
or U2492 (N_2492,N_1770,N_1554);
nand U2493 (N_2493,N_1452,N_1158);
nand U2494 (N_2494,N_1503,N_1337);
or U2495 (N_2495,N_1572,N_1786);
and U2496 (N_2496,N_1463,N_1729);
or U2497 (N_2497,N_1528,N_1821);
nand U2498 (N_2498,N_1719,N_1349);
nand U2499 (N_2499,N_1362,N_1931);
or U2500 (N_2500,N_1638,N_1343);
nand U2501 (N_2501,N_1374,N_1078);
nor U2502 (N_2502,N_1557,N_1524);
nand U2503 (N_2503,N_1464,N_1978);
and U2504 (N_2504,N_1019,N_1993);
or U2505 (N_2505,N_1917,N_1872);
nor U2506 (N_2506,N_1614,N_1925);
nor U2507 (N_2507,N_1061,N_1790);
nor U2508 (N_2508,N_1498,N_1500);
nand U2509 (N_2509,N_1665,N_1643);
and U2510 (N_2510,N_1063,N_1830);
and U2511 (N_2511,N_1694,N_1815);
or U2512 (N_2512,N_1974,N_1844);
and U2513 (N_2513,N_1903,N_1336);
nor U2514 (N_2514,N_1988,N_1777);
nand U2515 (N_2515,N_1646,N_1283);
and U2516 (N_2516,N_1203,N_1281);
nand U2517 (N_2517,N_1985,N_1429);
nand U2518 (N_2518,N_1129,N_1372);
nand U2519 (N_2519,N_1238,N_1639);
or U2520 (N_2520,N_1366,N_1765);
and U2521 (N_2521,N_1036,N_1500);
nand U2522 (N_2522,N_1954,N_1484);
xor U2523 (N_2523,N_1343,N_1450);
nand U2524 (N_2524,N_1248,N_1674);
nor U2525 (N_2525,N_1391,N_1057);
nand U2526 (N_2526,N_1395,N_1880);
nor U2527 (N_2527,N_1006,N_1162);
or U2528 (N_2528,N_1941,N_1910);
nand U2529 (N_2529,N_1544,N_1827);
nor U2530 (N_2530,N_1176,N_1061);
nor U2531 (N_2531,N_1322,N_1097);
nor U2532 (N_2532,N_1399,N_1130);
nor U2533 (N_2533,N_1906,N_1333);
or U2534 (N_2534,N_1056,N_1183);
nor U2535 (N_2535,N_1049,N_1561);
and U2536 (N_2536,N_1629,N_1102);
or U2537 (N_2537,N_1868,N_1950);
or U2538 (N_2538,N_1711,N_1401);
nand U2539 (N_2539,N_1768,N_1333);
nor U2540 (N_2540,N_1243,N_1874);
nor U2541 (N_2541,N_1057,N_1646);
or U2542 (N_2542,N_1324,N_1010);
and U2543 (N_2543,N_1318,N_1927);
or U2544 (N_2544,N_1581,N_1576);
nor U2545 (N_2545,N_1158,N_1873);
nor U2546 (N_2546,N_1534,N_1982);
nor U2547 (N_2547,N_1421,N_1960);
nor U2548 (N_2548,N_1320,N_1853);
or U2549 (N_2549,N_1798,N_1141);
and U2550 (N_2550,N_1617,N_1748);
and U2551 (N_2551,N_1569,N_1147);
and U2552 (N_2552,N_1933,N_1869);
nand U2553 (N_2553,N_1302,N_1242);
xnor U2554 (N_2554,N_1401,N_1999);
and U2555 (N_2555,N_1987,N_1567);
nand U2556 (N_2556,N_1142,N_1301);
nor U2557 (N_2557,N_1526,N_1441);
nand U2558 (N_2558,N_1645,N_1423);
nor U2559 (N_2559,N_1682,N_1909);
nand U2560 (N_2560,N_1583,N_1064);
or U2561 (N_2561,N_1347,N_1449);
nand U2562 (N_2562,N_1812,N_1749);
and U2563 (N_2563,N_1808,N_1702);
nand U2564 (N_2564,N_1306,N_1040);
nor U2565 (N_2565,N_1328,N_1411);
and U2566 (N_2566,N_1302,N_1218);
and U2567 (N_2567,N_1698,N_1410);
or U2568 (N_2568,N_1330,N_1078);
or U2569 (N_2569,N_1071,N_1579);
or U2570 (N_2570,N_1402,N_1125);
and U2571 (N_2571,N_1840,N_1504);
nor U2572 (N_2572,N_1631,N_1445);
and U2573 (N_2573,N_1196,N_1050);
and U2574 (N_2574,N_1392,N_1849);
nand U2575 (N_2575,N_1022,N_1346);
and U2576 (N_2576,N_1610,N_1944);
and U2577 (N_2577,N_1273,N_1816);
and U2578 (N_2578,N_1694,N_1492);
nor U2579 (N_2579,N_1494,N_1319);
nor U2580 (N_2580,N_1384,N_1939);
nand U2581 (N_2581,N_1188,N_1770);
and U2582 (N_2582,N_1522,N_1810);
or U2583 (N_2583,N_1076,N_1514);
xor U2584 (N_2584,N_1861,N_1875);
nand U2585 (N_2585,N_1028,N_1043);
nand U2586 (N_2586,N_1948,N_1545);
nor U2587 (N_2587,N_1277,N_1664);
nor U2588 (N_2588,N_1373,N_1765);
or U2589 (N_2589,N_1941,N_1283);
or U2590 (N_2590,N_1438,N_1495);
nand U2591 (N_2591,N_1213,N_1449);
or U2592 (N_2592,N_1995,N_1674);
or U2593 (N_2593,N_1026,N_1066);
and U2594 (N_2594,N_1807,N_1741);
and U2595 (N_2595,N_1415,N_1317);
or U2596 (N_2596,N_1985,N_1510);
nor U2597 (N_2597,N_1156,N_1745);
and U2598 (N_2598,N_1743,N_1615);
or U2599 (N_2599,N_1945,N_1767);
and U2600 (N_2600,N_1634,N_1149);
and U2601 (N_2601,N_1319,N_1159);
or U2602 (N_2602,N_1937,N_1605);
or U2603 (N_2603,N_1411,N_1880);
nand U2604 (N_2604,N_1122,N_1397);
nand U2605 (N_2605,N_1779,N_1530);
nor U2606 (N_2606,N_1960,N_1212);
nor U2607 (N_2607,N_1803,N_1072);
nand U2608 (N_2608,N_1436,N_1798);
or U2609 (N_2609,N_1547,N_1999);
nor U2610 (N_2610,N_1041,N_1433);
nor U2611 (N_2611,N_1082,N_1117);
and U2612 (N_2612,N_1299,N_1744);
xor U2613 (N_2613,N_1709,N_1364);
and U2614 (N_2614,N_1932,N_1177);
nor U2615 (N_2615,N_1578,N_1288);
or U2616 (N_2616,N_1799,N_1776);
nand U2617 (N_2617,N_1269,N_1920);
nand U2618 (N_2618,N_1180,N_1111);
or U2619 (N_2619,N_1479,N_1938);
nor U2620 (N_2620,N_1040,N_1641);
nand U2621 (N_2621,N_1973,N_1336);
or U2622 (N_2622,N_1434,N_1964);
nand U2623 (N_2623,N_1125,N_1458);
nor U2624 (N_2624,N_1405,N_1837);
or U2625 (N_2625,N_1193,N_1385);
nor U2626 (N_2626,N_1976,N_1063);
or U2627 (N_2627,N_1141,N_1500);
nand U2628 (N_2628,N_1837,N_1528);
and U2629 (N_2629,N_1100,N_1886);
and U2630 (N_2630,N_1807,N_1325);
nor U2631 (N_2631,N_1897,N_1849);
nand U2632 (N_2632,N_1918,N_1578);
nand U2633 (N_2633,N_1659,N_1587);
nor U2634 (N_2634,N_1205,N_1919);
or U2635 (N_2635,N_1676,N_1689);
nor U2636 (N_2636,N_1039,N_1137);
or U2637 (N_2637,N_1261,N_1406);
nand U2638 (N_2638,N_1557,N_1088);
and U2639 (N_2639,N_1189,N_1599);
nor U2640 (N_2640,N_1484,N_1430);
and U2641 (N_2641,N_1221,N_1940);
nand U2642 (N_2642,N_1075,N_1847);
and U2643 (N_2643,N_1837,N_1543);
nor U2644 (N_2644,N_1113,N_1448);
or U2645 (N_2645,N_1904,N_1837);
nor U2646 (N_2646,N_1120,N_1512);
nor U2647 (N_2647,N_1070,N_1630);
nand U2648 (N_2648,N_1243,N_1493);
and U2649 (N_2649,N_1601,N_1815);
nor U2650 (N_2650,N_1814,N_1850);
nand U2651 (N_2651,N_1267,N_1216);
or U2652 (N_2652,N_1991,N_1656);
xnor U2653 (N_2653,N_1811,N_1132);
nor U2654 (N_2654,N_1157,N_1191);
and U2655 (N_2655,N_1929,N_1693);
nand U2656 (N_2656,N_1098,N_1881);
and U2657 (N_2657,N_1455,N_1334);
and U2658 (N_2658,N_1981,N_1260);
nor U2659 (N_2659,N_1331,N_1162);
and U2660 (N_2660,N_1920,N_1447);
and U2661 (N_2661,N_1395,N_1531);
and U2662 (N_2662,N_1813,N_1835);
and U2663 (N_2663,N_1501,N_1553);
or U2664 (N_2664,N_1667,N_1909);
and U2665 (N_2665,N_1488,N_1185);
nand U2666 (N_2666,N_1519,N_1317);
nor U2667 (N_2667,N_1100,N_1254);
nand U2668 (N_2668,N_1929,N_1230);
nor U2669 (N_2669,N_1766,N_1330);
xnor U2670 (N_2670,N_1674,N_1605);
and U2671 (N_2671,N_1389,N_1151);
nor U2672 (N_2672,N_1127,N_1520);
or U2673 (N_2673,N_1940,N_1640);
xor U2674 (N_2674,N_1456,N_1355);
nand U2675 (N_2675,N_1406,N_1611);
nand U2676 (N_2676,N_1910,N_1642);
nand U2677 (N_2677,N_1243,N_1081);
nand U2678 (N_2678,N_1345,N_1478);
nor U2679 (N_2679,N_1236,N_1792);
and U2680 (N_2680,N_1642,N_1183);
and U2681 (N_2681,N_1658,N_1780);
nand U2682 (N_2682,N_1962,N_1044);
and U2683 (N_2683,N_1910,N_1485);
or U2684 (N_2684,N_1626,N_1744);
or U2685 (N_2685,N_1068,N_1800);
or U2686 (N_2686,N_1981,N_1875);
nor U2687 (N_2687,N_1470,N_1004);
nor U2688 (N_2688,N_1052,N_1448);
and U2689 (N_2689,N_1605,N_1929);
nand U2690 (N_2690,N_1954,N_1946);
nor U2691 (N_2691,N_1344,N_1962);
and U2692 (N_2692,N_1184,N_1236);
nand U2693 (N_2693,N_1046,N_1121);
nor U2694 (N_2694,N_1910,N_1337);
or U2695 (N_2695,N_1856,N_1512);
and U2696 (N_2696,N_1162,N_1554);
nor U2697 (N_2697,N_1270,N_1517);
nand U2698 (N_2698,N_1896,N_1359);
nand U2699 (N_2699,N_1993,N_1391);
or U2700 (N_2700,N_1663,N_1439);
nand U2701 (N_2701,N_1925,N_1095);
and U2702 (N_2702,N_1147,N_1944);
nor U2703 (N_2703,N_1233,N_1562);
or U2704 (N_2704,N_1248,N_1010);
nand U2705 (N_2705,N_1668,N_1401);
nand U2706 (N_2706,N_1671,N_1423);
and U2707 (N_2707,N_1124,N_1063);
or U2708 (N_2708,N_1129,N_1067);
and U2709 (N_2709,N_1041,N_1838);
nand U2710 (N_2710,N_1660,N_1429);
xor U2711 (N_2711,N_1358,N_1447);
nor U2712 (N_2712,N_1046,N_1643);
and U2713 (N_2713,N_1492,N_1028);
nor U2714 (N_2714,N_1017,N_1581);
nand U2715 (N_2715,N_1130,N_1642);
and U2716 (N_2716,N_1615,N_1484);
nor U2717 (N_2717,N_1066,N_1783);
nand U2718 (N_2718,N_1238,N_1487);
nor U2719 (N_2719,N_1747,N_1781);
nand U2720 (N_2720,N_1055,N_1551);
nor U2721 (N_2721,N_1557,N_1001);
nand U2722 (N_2722,N_1395,N_1423);
nor U2723 (N_2723,N_1703,N_1115);
nand U2724 (N_2724,N_1590,N_1163);
nor U2725 (N_2725,N_1372,N_1247);
nand U2726 (N_2726,N_1228,N_1131);
nor U2727 (N_2727,N_1196,N_1890);
nor U2728 (N_2728,N_1912,N_1734);
and U2729 (N_2729,N_1112,N_1917);
nand U2730 (N_2730,N_1709,N_1554);
nor U2731 (N_2731,N_1345,N_1670);
and U2732 (N_2732,N_1074,N_1842);
and U2733 (N_2733,N_1762,N_1988);
nor U2734 (N_2734,N_1427,N_1949);
nor U2735 (N_2735,N_1644,N_1727);
and U2736 (N_2736,N_1234,N_1357);
or U2737 (N_2737,N_1340,N_1124);
nor U2738 (N_2738,N_1877,N_1935);
or U2739 (N_2739,N_1110,N_1146);
or U2740 (N_2740,N_1688,N_1481);
or U2741 (N_2741,N_1147,N_1720);
xnor U2742 (N_2742,N_1768,N_1772);
nand U2743 (N_2743,N_1018,N_1134);
and U2744 (N_2744,N_1116,N_1326);
or U2745 (N_2745,N_1744,N_1163);
or U2746 (N_2746,N_1888,N_1372);
and U2747 (N_2747,N_1581,N_1768);
nand U2748 (N_2748,N_1196,N_1757);
or U2749 (N_2749,N_1182,N_1545);
or U2750 (N_2750,N_1440,N_1115);
nor U2751 (N_2751,N_1614,N_1023);
nor U2752 (N_2752,N_1397,N_1766);
or U2753 (N_2753,N_1800,N_1021);
nand U2754 (N_2754,N_1180,N_1573);
nand U2755 (N_2755,N_1616,N_1101);
and U2756 (N_2756,N_1604,N_1982);
nand U2757 (N_2757,N_1484,N_1590);
nor U2758 (N_2758,N_1446,N_1964);
or U2759 (N_2759,N_1384,N_1476);
and U2760 (N_2760,N_1231,N_1434);
nand U2761 (N_2761,N_1704,N_1702);
and U2762 (N_2762,N_1656,N_1006);
nor U2763 (N_2763,N_1242,N_1733);
and U2764 (N_2764,N_1233,N_1313);
nor U2765 (N_2765,N_1580,N_1673);
and U2766 (N_2766,N_1519,N_1636);
and U2767 (N_2767,N_1485,N_1202);
nor U2768 (N_2768,N_1206,N_1299);
nand U2769 (N_2769,N_1072,N_1115);
or U2770 (N_2770,N_1594,N_1411);
nand U2771 (N_2771,N_1332,N_1639);
and U2772 (N_2772,N_1986,N_1955);
or U2773 (N_2773,N_1132,N_1773);
and U2774 (N_2774,N_1064,N_1999);
and U2775 (N_2775,N_1704,N_1005);
or U2776 (N_2776,N_1978,N_1694);
nor U2777 (N_2777,N_1453,N_1005);
nor U2778 (N_2778,N_1606,N_1085);
nand U2779 (N_2779,N_1357,N_1051);
nor U2780 (N_2780,N_1551,N_1573);
and U2781 (N_2781,N_1858,N_1714);
nand U2782 (N_2782,N_1629,N_1466);
nand U2783 (N_2783,N_1374,N_1299);
nor U2784 (N_2784,N_1339,N_1201);
nor U2785 (N_2785,N_1234,N_1409);
nand U2786 (N_2786,N_1301,N_1327);
or U2787 (N_2787,N_1642,N_1667);
nand U2788 (N_2788,N_1959,N_1989);
xnor U2789 (N_2789,N_1482,N_1612);
nand U2790 (N_2790,N_1478,N_1580);
or U2791 (N_2791,N_1739,N_1066);
or U2792 (N_2792,N_1344,N_1910);
and U2793 (N_2793,N_1966,N_1073);
or U2794 (N_2794,N_1563,N_1054);
nand U2795 (N_2795,N_1789,N_1724);
nand U2796 (N_2796,N_1880,N_1469);
nand U2797 (N_2797,N_1821,N_1622);
nand U2798 (N_2798,N_1960,N_1689);
or U2799 (N_2799,N_1838,N_1660);
nand U2800 (N_2800,N_1330,N_1437);
nand U2801 (N_2801,N_1661,N_1377);
and U2802 (N_2802,N_1152,N_1331);
or U2803 (N_2803,N_1095,N_1828);
nand U2804 (N_2804,N_1565,N_1934);
nor U2805 (N_2805,N_1027,N_1444);
and U2806 (N_2806,N_1411,N_1109);
nor U2807 (N_2807,N_1106,N_1742);
and U2808 (N_2808,N_1828,N_1204);
nor U2809 (N_2809,N_1357,N_1869);
or U2810 (N_2810,N_1306,N_1830);
and U2811 (N_2811,N_1540,N_1980);
and U2812 (N_2812,N_1562,N_1592);
and U2813 (N_2813,N_1237,N_1633);
nor U2814 (N_2814,N_1035,N_1118);
nor U2815 (N_2815,N_1562,N_1173);
and U2816 (N_2816,N_1361,N_1555);
nand U2817 (N_2817,N_1622,N_1735);
and U2818 (N_2818,N_1514,N_1625);
nand U2819 (N_2819,N_1558,N_1950);
or U2820 (N_2820,N_1151,N_1142);
nand U2821 (N_2821,N_1288,N_1148);
nand U2822 (N_2822,N_1464,N_1663);
nand U2823 (N_2823,N_1591,N_1737);
or U2824 (N_2824,N_1869,N_1199);
nand U2825 (N_2825,N_1112,N_1908);
or U2826 (N_2826,N_1177,N_1430);
nor U2827 (N_2827,N_1618,N_1676);
and U2828 (N_2828,N_1782,N_1424);
or U2829 (N_2829,N_1437,N_1075);
and U2830 (N_2830,N_1941,N_1658);
nand U2831 (N_2831,N_1213,N_1665);
and U2832 (N_2832,N_1615,N_1747);
nand U2833 (N_2833,N_1297,N_1573);
xnor U2834 (N_2834,N_1053,N_1307);
and U2835 (N_2835,N_1547,N_1789);
or U2836 (N_2836,N_1348,N_1916);
and U2837 (N_2837,N_1949,N_1455);
or U2838 (N_2838,N_1679,N_1615);
nor U2839 (N_2839,N_1118,N_1358);
nand U2840 (N_2840,N_1240,N_1388);
nor U2841 (N_2841,N_1856,N_1183);
or U2842 (N_2842,N_1734,N_1371);
nor U2843 (N_2843,N_1310,N_1017);
nand U2844 (N_2844,N_1331,N_1119);
and U2845 (N_2845,N_1336,N_1613);
or U2846 (N_2846,N_1942,N_1993);
or U2847 (N_2847,N_1512,N_1618);
nand U2848 (N_2848,N_1688,N_1834);
nand U2849 (N_2849,N_1736,N_1687);
or U2850 (N_2850,N_1790,N_1682);
nor U2851 (N_2851,N_1176,N_1409);
or U2852 (N_2852,N_1607,N_1071);
nor U2853 (N_2853,N_1978,N_1144);
nand U2854 (N_2854,N_1939,N_1719);
and U2855 (N_2855,N_1213,N_1077);
nor U2856 (N_2856,N_1514,N_1248);
or U2857 (N_2857,N_1080,N_1145);
or U2858 (N_2858,N_1176,N_1844);
or U2859 (N_2859,N_1885,N_1955);
nand U2860 (N_2860,N_1926,N_1860);
and U2861 (N_2861,N_1185,N_1029);
and U2862 (N_2862,N_1251,N_1862);
nand U2863 (N_2863,N_1092,N_1155);
and U2864 (N_2864,N_1052,N_1294);
nand U2865 (N_2865,N_1365,N_1626);
and U2866 (N_2866,N_1632,N_1610);
and U2867 (N_2867,N_1896,N_1180);
or U2868 (N_2868,N_1580,N_1633);
nand U2869 (N_2869,N_1689,N_1008);
nor U2870 (N_2870,N_1528,N_1922);
nand U2871 (N_2871,N_1924,N_1861);
nand U2872 (N_2872,N_1217,N_1873);
nand U2873 (N_2873,N_1186,N_1088);
or U2874 (N_2874,N_1366,N_1848);
and U2875 (N_2875,N_1285,N_1126);
and U2876 (N_2876,N_1539,N_1467);
and U2877 (N_2877,N_1588,N_1645);
and U2878 (N_2878,N_1589,N_1927);
or U2879 (N_2879,N_1120,N_1603);
nor U2880 (N_2880,N_1745,N_1021);
and U2881 (N_2881,N_1293,N_1311);
nor U2882 (N_2882,N_1246,N_1334);
or U2883 (N_2883,N_1700,N_1007);
and U2884 (N_2884,N_1754,N_1225);
nor U2885 (N_2885,N_1055,N_1748);
and U2886 (N_2886,N_1151,N_1649);
or U2887 (N_2887,N_1221,N_1231);
or U2888 (N_2888,N_1658,N_1513);
nand U2889 (N_2889,N_1761,N_1067);
and U2890 (N_2890,N_1804,N_1771);
or U2891 (N_2891,N_1836,N_1809);
nand U2892 (N_2892,N_1250,N_1881);
nor U2893 (N_2893,N_1367,N_1839);
and U2894 (N_2894,N_1847,N_1946);
or U2895 (N_2895,N_1664,N_1653);
nor U2896 (N_2896,N_1750,N_1204);
and U2897 (N_2897,N_1839,N_1059);
or U2898 (N_2898,N_1307,N_1491);
or U2899 (N_2899,N_1530,N_1048);
and U2900 (N_2900,N_1223,N_1920);
nand U2901 (N_2901,N_1511,N_1227);
and U2902 (N_2902,N_1173,N_1517);
nand U2903 (N_2903,N_1173,N_1925);
or U2904 (N_2904,N_1686,N_1386);
and U2905 (N_2905,N_1376,N_1984);
nor U2906 (N_2906,N_1049,N_1692);
or U2907 (N_2907,N_1250,N_1754);
nand U2908 (N_2908,N_1901,N_1590);
or U2909 (N_2909,N_1902,N_1026);
nor U2910 (N_2910,N_1850,N_1318);
nand U2911 (N_2911,N_1785,N_1083);
nor U2912 (N_2912,N_1930,N_1890);
or U2913 (N_2913,N_1216,N_1450);
nand U2914 (N_2914,N_1504,N_1442);
or U2915 (N_2915,N_1545,N_1133);
and U2916 (N_2916,N_1735,N_1985);
nand U2917 (N_2917,N_1419,N_1637);
or U2918 (N_2918,N_1387,N_1346);
or U2919 (N_2919,N_1340,N_1636);
or U2920 (N_2920,N_1439,N_1850);
nor U2921 (N_2921,N_1955,N_1322);
and U2922 (N_2922,N_1336,N_1965);
nor U2923 (N_2923,N_1541,N_1614);
nand U2924 (N_2924,N_1929,N_1790);
nor U2925 (N_2925,N_1522,N_1660);
and U2926 (N_2926,N_1805,N_1031);
xor U2927 (N_2927,N_1621,N_1852);
or U2928 (N_2928,N_1316,N_1972);
nor U2929 (N_2929,N_1698,N_1626);
nor U2930 (N_2930,N_1110,N_1354);
and U2931 (N_2931,N_1722,N_1281);
nand U2932 (N_2932,N_1489,N_1844);
nand U2933 (N_2933,N_1828,N_1767);
and U2934 (N_2934,N_1546,N_1450);
nand U2935 (N_2935,N_1310,N_1860);
nor U2936 (N_2936,N_1600,N_1746);
and U2937 (N_2937,N_1858,N_1441);
nor U2938 (N_2938,N_1849,N_1794);
and U2939 (N_2939,N_1514,N_1498);
or U2940 (N_2940,N_1173,N_1882);
nor U2941 (N_2941,N_1318,N_1158);
nand U2942 (N_2942,N_1298,N_1426);
nor U2943 (N_2943,N_1495,N_1538);
and U2944 (N_2944,N_1778,N_1972);
nor U2945 (N_2945,N_1173,N_1337);
or U2946 (N_2946,N_1417,N_1178);
and U2947 (N_2947,N_1362,N_1535);
nand U2948 (N_2948,N_1580,N_1890);
and U2949 (N_2949,N_1842,N_1021);
nand U2950 (N_2950,N_1809,N_1597);
nor U2951 (N_2951,N_1162,N_1928);
nor U2952 (N_2952,N_1954,N_1786);
nor U2953 (N_2953,N_1717,N_1667);
and U2954 (N_2954,N_1251,N_1794);
nand U2955 (N_2955,N_1973,N_1239);
nor U2956 (N_2956,N_1429,N_1221);
and U2957 (N_2957,N_1268,N_1120);
and U2958 (N_2958,N_1239,N_1939);
and U2959 (N_2959,N_1696,N_1611);
or U2960 (N_2960,N_1401,N_1452);
and U2961 (N_2961,N_1012,N_1466);
and U2962 (N_2962,N_1584,N_1538);
and U2963 (N_2963,N_1923,N_1139);
and U2964 (N_2964,N_1767,N_1696);
and U2965 (N_2965,N_1115,N_1734);
nor U2966 (N_2966,N_1551,N_1769);
nor U2967 (N_2967,N_1624,N_1015);
and U2968 (N_2968,N_1130,N_1869);
and U2969 (N_2969,N_1440,N_1972);
and U2970 (N_2970,N_1589,N_1291);
and U2971 (N_2971,N_1316,N_1357);
and U2972 (N_2972,N_1906,N_1326);
nor U2973 (N_2973,N_1333,N_1642);
nand U2974 (N_2974,N_1868,N_1645);
or U2975 (N_2975,N_1421,N_1907);
and U2976 (N_2976,N_1274,N_1328);
nand U2977 (N_2977,N_1490,N_1773);
or U2978 (N_2978,N_1371,N_1792);
nand U2979 (N_2979,N_1500,N_1565);
or U2980 (N_2980,N_1124,N_1345);
or U2981 (N_2981,N_1478,N_1084);
nor U2982 (N_2982,N_1483,N_1829);
and U2983 (N_2983,N_1722,N_1266);
nand U2984 (N_2984,N_1912,N_1919);
and U2985 (N_2985,N_1623,N_1928);
nor U2986 (N_2986,N_1812,N_1349);
and U2987 (N_2987,N_1100,N_1261);
and U2988 (N_2988,N_1175,N_1994);
and U2989 (N_2989,N_1664,N_1204);
nor U2990 (N_2990,N_1342,N_1952);
nand U2991 (N_2991,N_1939,N_1741);
nand U2992 (N_2992,N_1327,N_1069);
and U2993 (N_2993,N_1326,N_1902);
or U2994 (N_2994,N_1754,N_1870);
and U2995 (N_2995,N_1701,N_1905);
or U2996 (N_2996,N_1973,N_1498);
and U2997 (N_2997,N_1547,N_1336);
or U2998 (N_2998,N_1173,N_1614);
nor U2999 (N_2999,N_1120,N_1232);
nand U3000 (N_3000,N_2259,N_2724);
and U3001 (N_3001,N_2386,N_2780);
nor U3002 (N_3002,N_2102,N_2237);
and U3003 (N_3003,N_2223,N_2045);
and U3004 (N_3004,N_2631,N_2271);
and U3005 (N_3005,N_2784,N_2994);
nor U3006 (N_3006,N_2949,N_2554);
or U3007 (N_3007,N_2912,N_2123);
nand U3008 (N_3008,N_2312,N_2461);
or U3009 (N_3009,N_2925,N_2566);
nor U3010 (N_3010,N_2786,N_2677);
or U3011 (N_3011,N_2194,N_2487);
nor U3012 (N_3012,N_2068,N_2836);
or U3013 (N_3013,N_2191,N_2519);
and U3014 (N_3014,N_2426,N_2051);
nand U3015 (N_3015,N_2336,N_2712);
and U3016 (N_3016,N_2470,N_2409);
nor U3017 (N_3017,N_2553,N_2720);
or U3018 (N_3018,N_2258,N_2290);
or U3019 (N_3019,N_2961,N_2615);
nand U3020 (N_3020,N_2438,N_2732);
nand U3021 (N_3021,N_2681,N_2176);
and U3022 (N_3022,N_2061,N_2083);
and U3023 (N_3023,N_2413,N_2215);
nor U3024 (N_3024,N_2182,N_2991);
and U3025 (N_3025,N_2486,N_2457);
and U3026 (N_3026,N_2520,N_2451);
nand U3027 (N_3027,N_2391,N_2735);
nor U3028 (N_3028,N_2659,N_2888);
nand U3029 (N_3029,N_2620,N_2455);
nor U3030 (N_3030,N_2179,N_2710);
and U3031 (N_3031,N_2129,N_2639);
nand U3032 (N_3032,N_2465,N_2142);
or U3033 (N_3033,N_2227,N_2035);
and U3034 (N_3034,N_2221,N_2698);
or U3035 (N_3035,N_2313,N_2351);
and U3036 (N_3036,N_2376,N_2481);
and U3037 (N_3037,N_2892,N_2324);
or U3038 (N_3038,N_2610,N_2901);
nor U3039 (N_3039,N_2619,N_2573);
and U3040 (N_3040,N_2740,N_2785);
nor U3041 (N_3041,N_2604,N_2136);
and U3042 (N_3042,N_2776,N_2704);
nor U3043 (N_3043,N_2502,N_2262);
or U3044 (N_3044,N_2467,N_2371);
xnor U3045 (N_3045,N_2529,N_2331);
and U3046 (N_3046,N_2781,N_2415);
nor U3047 (N_3047,N_2877,N_2468);
nor U3048 (N_3048,N_2446,N_2008);
nor U3049 (N_3049,N_2010,N_2178);
nor U3050 (N_3050,N_2791,N_2950);
nor U3051 (N_3051,N_2322,N_2755);
nor U3052 (N_3052,N_2841,N_2066);
or U3053 (N_3053,N_2072,N_2640);
or U3054 (N_3054,N_2004,N_2301);
nor U3055 (N_3055,N_2354,N_2396);
nor U3056 (N_3056,N_2911,N_2863);
or U3057 (N_3057,N_2975,N_2434);
or U3058 (N_3058,N_2431,N_2500);
nand U3059 (N_3059,N_2655,N_2666);
or U3060 (N_3060,N_2978,N_2582);
nand U3061 (N_3061,N_2071,N_2183);
nor U3062 (N_3062,N_2737,N_2211);
nor U3063 (N_3063,N_2144,N_2496);
and U3064 (N_3064,N_2809,N_2074);
and U3065 (N_3065,N_2593,N_2253);
or U3066 (N_3066,N_2318,N_2942);
and U3067 (N_3067,N_2319,N_2694);
or U3068 (N_3068,N_2377,N_2646);
and U3069 (N_3069,N_2518,N_2944);
nor U3070 (N_3070,N_2130,N_2343);
nor U3071 (N_3071,N_2335,N_2374);
and U3072 (N_3072,N_2098,N_2663);
nand U3073 (N_3073,N_2344,N_2804);
or U3074 (N_3074,N_2450,N_2839);
and U3075 (N_3075,N_2011,N_2418);
nor U3076 (N_3076,N_2443,N_2998);
nand U3077 (N_3077,N_2169,N_2889);
nand U3078 (N_3078,N_2497,N_2628);
nor U3079 (N_3079,N_2736,N_2357);
nor U3080 (N_3080,N_2820,N_2229);
and U3081 (N_3081,N_2858,N_2452);
nand U3082 (N_3082,N_2430,N_2203);
nor U3083 (N_3083,N_2362,N_2078);
nor U3084 (N_3084,N_2972,N_2089);
nand U3085 (N_3085,N_2556,N_2760);
or U3086 (N_3086,N_2161,N_2128);
nand U3087 (N_3087,N_2289,N_2267);
nand U3088 (N_3088,N_2846,N_2095);
and U3089 (N_3089,N_2297,N_2032);
and U3090 (N_3090,N_2230,N_2635);
nor U3091 (N_3091,N_2742,N_2985);
xnor U3092 (N_3092,N_2600,N_2898);
nor U3093 (N_3093,N_2086,N_2674);
nand U3094 (N_3094,N_2580,N_2495);
nor U3095 (N_3095,N_2433,N_2204);
and U3096 (N_3096,N_2454,N_2423);
nand U3097 (N_3097,N_2904,N_2940);
nor U3098 (N_3098,N_2387,N_2762);
xor U3099 (N_3099,N_2545,N_2462);
nand U3100 (N_3100,N_2231,N_2225);
and U3101 (N_3101,N_2206,N_2918);
nor U3102 (N_3102,N_2798,N_2705);
or U3103 (N_3103,N_2234,N_2268);
nand U3104 (N_3104,N_2624,N_2516);
nand U3105 (N_3105,N_2778,N_2796);
nor U3106 (N_3106,N_2192,N_2326);
nor U3107 (N_3107,N_2350,N_2676);
nand U3108 (N_3108,N_2125,N_2936);
nor U3109 (N_3109,N_2018,N_2026);
nor U3110 (N_3110,N_2541,N_2700);
or U3111 (N_3111,N_2706,N_2616);
or U3112 (N_3112,N_2818,N_2341);
and U3113 (N_3113,N_2730,N_2356);
or U3114 (N_3114,N_2217,N_2260);
nand U3115 (N_3115,N_2550,N_2902);
or U3116 (N_3116,N_2243,N_2862);
or U3117 (N_3117,N_2759,N_2568);
nand U3118 (N_3118,N_2650,N_2772);
nand U3119 (N_3119,N_2005,N_2514);
or U3120 (N_3120,N_2840,N_2265);
and U3121 (N_3121,N_2441,N_2490);
and U3122 (N_3122,N_2075,N_2345);
or U3123 (N_3123,N_2928,N_2442);
or U3124 (N_3124,N_2276,N_2524);
nor U3125 (N_3125,N_2381,N_2625);
nor U3126 (N_3126,N_2421,N_2167);
nand U3127 (N_3127,N_2241,N_2743);
nand U3128 (N_3128,N_2948,N_2475);
or U3129 (N_3129,N_2453,N_2419);
or U3130 (N_3130,N_2521,N_2716);
and U3131 (N_3131,N_2166,N_2581);
or U3132 (N_3132,N_2645,N_2835);
nand U3133 (N_3133,N_2565,N_2627);
and U3134 (N_3134,N_2802,N_2432);
nand U3135 (N_3135,N_2091,N_2284);
nor U3136 (N_3136,N_2188,N_2049);
nand U3137 (N_3137,N_2968,N_2137);
nor U3138 (N_3138,N_2164,N_2210);
and U3139 (N_3139,N_2879,N_2375);
or U3140 (N_3140,N_2492,N_2153);
or U3141 (N_3141,N_2036,N_2812);
nand U3142 (N_3142,N_2272,N_2233);
nand U3143 (N_3143,N_2771,N_2919);
nor U3144 (N_3144,N_2544,N_2852);
nor U3145 (N_3145,N_2346,N_2797);
and U3146 (N_3146,N_2684,N_2559);
and U3147 (N_3147,N_2849,N_2685);
nor U3148 (N_3148,N_2993,N_2517);
and U3149 (N_3149,N_2597,N_2574);
nor U3150 (N_3150,N_2886,N_2117);
xnor U3151 (N_3151,N_2410,N_2151);
xor U3152 (N_3152,N_2913,N_2763);
and U3153 (N_3153,N_2388,N_2589);
nand U3154 (N_3154,N_2569,N_2965);
or U3155 (N_3155,N_2379,N_2917);
nor U3156 (N_3156,N_2941,N_2850);
nand U3157 (N_3157,N_2583,N_2408);
nor U3158 (N_3158,N_2810,N_2533);
nor U3159 (N_3159,N_2165,N_2945);
xor U3160 (N_3160,N_2017,N_2548);
nor U3161 (N_3161,N_2296,N_2093);
and U3162 (N_3162,N_2672,N_2708);
and U3163 (N_3163,N_2722,N_2025);
nand U3164 (N_3164,N_2857,N_2067);
or U3165 (N_3165,N_2177,N_2493);
and U3166 (N_3166,N_2920,N_2437);
nand U3167 (N_3167,N_2242,N_2404);
and U3168 (N_3168,N_2788,N_2294);
nand U3169 (N_3169,N_2361,N_2946);
nand U3170 (N_3170,N_2293,N_2277);
nand U3171 (N_3171,N_2711,N_2751);
and U3172 (N_3172,N_2629,N_2668);
nor U3173 (N_3173,N_2922,N_2428);
or U3174 (N_3174,N_2990,N_2828);
nand U3175 (N_3175,N_2585,N_2477);
nor U3176 (N_3176,N_2355,N_2526);
and U3177 (N_3177,N_2915,N_2534);
or U3178 (N_3178,N_2825,N_2956);
or U3179 (N_3179,N_2370,N_2607);
nor U3180 (N_3180,N_2831,N_2739);
or U3181 (N_3181,N_2555,N_2824);
nor U3182 (N_3182,N_2982,N_2218);
or U3183 (N_3183,N_2140,N_2564);
nand U3184 (N_3184,N_2546,N_2422);
nor U3185 (N_3185,N_2727,N_2342);
nor U3186 (N_3186,N_2082,N_2851);
nand U3187 (N_3187,N_2504,N_2133);
and U3188 (N_3188,N_2845,N_2463);
or U3189 (N_3189,N_2606,N_2283);
and U3190 (N_3190,N_2172,N_2329);
and U3191 (N_3191,N_2333,N_2959);
and U3192 (N_3192,N_2506,N_2984);
and U3193 (N_3193,N_2875,N_2733);
and U3194 (N_3194,N_2721,N_2270);
and U3195 (N_3195,N_2171,N_2561);
xnor U3196 (N_3196,N_2731,N_2819);
nor U3197 (N_3197,N_2671,N_2943);
and U3198 (N_3198,N_2661,N_2577);
nand U3199 (N_3199,N_2843,N_2557);
and U3200 (N_3200,N_2150,N_2367);
nand U3201 (N_3201,N_2981,N_2251);
xnor U3202 (N_3202,N_2339,N_2152);
nor U3203 (N_3203,N_2592,N_2000);
nor U3204 (N_3204,N_2603,N_2590);
nand U3205 (N_3205,N_2479,N_2031);
and U3206 (N_3206,N_2632,N_2837);
and U3207 (N_3207,N_2325,N_2139);
nand U3208 (N_3208,N_2833,N_2330);
and U3209 (N_3209,N_2114,N_2397);
and U3210 (N_3210,N_2013,N_2247);
nor U3211 (N_3211,N_2073,N_2586);
and U3212 (N_3212,N_2692,N_2910);
and U3213 (N_3213,N_2955,N_2807);
or U3214 (N_3214,N_2893,N_2108);
and U3215 (N_3215,N_2316,N_2750);
or U3216 (N_3216,N_2085,N_2808);
or U3217 (N_3217,N_2048,N_2682);
and U3218 (N_3218,N_2273,N_2449);
nand U3219 (N_3219,N_2488,N_2158);
and U3220 (N_3220,N_2947,N_2899);
and U3221 (N_3221,N_2505,N_2884);
nor U3222 (N_3222,N_2090,N_2199);
or U3223 (N_3223,N_2063,N_2480);
nand U3224 (N_3224,N_2257,N_2040);
nand U3225 (N_3225,N_2053,N_2088);
or U3226 (N_3226,N_2932,N_2281);
nand U3227 (N_3227,N_2044,N_2938);
nand U3228 (N_3228,N_2159,N_2216);
and U3229 (N_3229,N_2327,N_2195);
nor U3230 (N_3230,N_2775,N_2653);
nor U3231 (N_3231,N_2832,N_2099);
or U3232 (N_3232,N_2608,N_2077);
or U3233 (N_3233,N_2907,N_2767);
and U3234 (N_3234,N_2774,N_2359);
nand U3235 (N_3235,N_2236,N_2122);
nand U3236 (N_3236,N_2795,N_2429);
and U3237 (N_3237,N_2255,N_2952);
nand U3238 (N_3238,N_2538,N_2185);
or U3239 (N_3239,N_2363,N_2749);
nor U3240 (N_3240,N_2113,N_2707);
nand U3241 (N_3241,N_2773,N_2079);
nand U3242 (N_3242,N_2612,N_2880);
or U3243 (N_3243,N_2180,N_2485);
or U3244 (N_3244,N_2822,N_2552);
nand U3245 (N_3245,N_2537,N_2300);
nor U3246 (N_3246,N_2092,N_2829);
xor U3247 (N_3247,N_2060,N_2794);
or U3248 (N_3248,N_2378,N_2842);
xor U3249 (N_3249,N_2473,N_2623);
nor U3250 (N_3250,N_2870,N_2405);
nor U3251 (N_3251,N_2382,N_2679);
and U3252 (N_3252,N_2403,N_2637);
or U3253 (N_3253,N_2906,N_2864);
nor U3254 (N_3254,N_2718,N_2368);
or U3255 (N_3255,N_2799,N_2921);
or U3256 (N_3256,N_2156,N_2512);
or U3257 (N_3257,N_2530,N_2872);
nand U3258 (N_3258,N_2527,N_2935);
nand U3259 (N_3259,N_2197,N_2303);
nand U3260 (N_3260,N_2996,N_2372);
or U3261 (N_3261,N_2189,N_2069);
or U3262 (N_3262,N_2212,N_2278);
nand U3263 (N_3263,N_2636,N_2535);
or U3264 (N_3264,N_2638,N_2246);
nor U3265 (N_3265,N_2688,N_2908);
nand U3266 (N_3266,N_2364,N_2168);
nand U3267 (N_3267,N_2240,N_2869);
and U3268 (N_3268,N_2295,N_2957);
nand U3269 (N_3269,N_2205,N_2081);
nand U3270 (N_3270,N_2929,N_2207);
and U3271 (N_3271,N_2890,N_2777);
nand U3272 (N_3272,N_2758,N_2916);
nand U3273 (N_3273,N_2579,N_2369);
or U3274 (N_3274,N_2466,N_2914);
nor U3275 (N_3275,N_2058,N_2201);
and U3276 (N_3276,N_2232,N_2347);
or U3277 (N_3277,N_2334,N_2046);
nand U3278 (N_3278,N_2016,N_2726);
nor U3279 (N_3279,N_2562,N_2444);
and U3280 (N_3280,N_2811,N_2023);
nand U3281 (N_3281,N_2392,N_2245);
nor U3282 (N_3282,N_2588,N_2633);
or U3283 (N_3283,N_2332,N_2644);
nor U3284 (N_3284,N_2613,N_2385);
or U3285 (N_3285,N_2815,N_2252);
or U3286 (N_3286,N_2728,N_2966);
or U3287 (N_3287,N_2611,N_2744);
and U3288 (N_3288,N_2275,N_2539);
or U3289 (N_3289,N_2838,N_2503);
nor U3290 (N_3290,N_2003,N_2121);
and U3291 (N_3291,N_2037,N_2543);
and U3292 (N_3292,N_2126,N_2790);
or U3293 (N_3293,N_2630,N_2494);
or U3294 (N_3294,N_2274,N_2508);
xnor U3295 (N_3295,N_2399,N_2393);
or U3296 (N_3296,N_2039,N_2244);
and U3297 (N_3297,N_2891,N_2792);
nor U3298 (N_3298,N_2304,N_2106);
nand U3299 (N_3299,N_2691,N_2100);
or U3300 (N_3300,N_2525,N_2248);
or U3301 (N_3301,N_2305,N_2690);
nand U3302 (N_3302,N_2202,N_2697);
nor U3303 (N_3303,N_2686,N_2173);
nand U3304 (N_3304,N_2622,N_2859);
or U3305 (N_3305,N_2513,N_2400);
or U3306 (N_3306,N_2927,N_2980);
nand U3307 (N_3307,N_2406,N_2154);
and U3308 (N_3308,N_2407,N_2469);
nand U3309 (N_3309,N_2097,N_2311);
or U3310 (N_3310,N_2987,N_2900);
or U3311 (N_3311,N_2412,N_2286);
nor U3312 (N_3312,N_2033,N_2282);
or U3313 (N_3313,N_2220,N_2427);
or U3314 (N_3314,N_2747,N_2020);
and U3315 (N_3315,N_2848,N_2222);
or U3316 (N_3316,N_2971,N_2219);
nor U3317 (N_3317,N_2757,N_2522);
and U3318 (N_3318,N_2654,N_2417);
nand U3319 (N_3319,N_2181,N_2584);
nand U3320 (N_3320,N_2157,N_2816);
nor U3321 (N_3321,N_2658,N_2292);
nor U3322 (N_3322,N_2214,N_2977);
nand U3323 (N_3323,N_2782,N_2456);
and U3324 (N_3324,N_2547,N_2306);
xnor U3325 (N_3325,N_2034,N_2563);
and U3326 (N_3326,N_2976,N_2989);
nor U3327 (N_3327,N_2614,N_2349);
or U3328 (N_3328,N_2143,N_2052);
nand U3329 (N_3329,N_2643,N_2752);
nor U3330 (N_3330,N_2883,N_2315);
nand U3331 (N_3331,N_2992,N_2012);
and U3332 (N_3332,N_2155,N_2395);
nor U3333 (N_3333,N_2605,N_2963);
nand U3334 (N_3334,N_2933,N_2854);
nor U3335 (N_3335,N_2145,N_2373);
nand U3336 (N_3336,N_2873,N_2065);
and U3337 (N_3337,N_2340,N_2411);
and U3338 (N_3338,N_2055,N_2865);
or U3339 (N_3339,N_2196,N_2054);
and U3340 (N_3340,N_2254,N_2954);
nor U3341 (N_3341,N_2560,N_2856);
and U3342 (N_3342,N_2894,N_2476);
nand U3343 (N_3343,N_2734,N_2909);
nor U3344 (N_3344,N_2116,N_2308);
nor U3345 (N_3345,N_2056,N_2876);
nor U3346 (N_3346,N_2649,N_2022);
or U3347 (N_3347,N_2120,N_2621);
nor U3348 (N_3348,N_2200,N_2328);
and U3349 (N_3349,N_2101,N_2830);
nand U3350 (N_3350,N_2964,N_2360);
or U3351 (N_3351,N_2314,N_2986);
nor U3352 (N_3352,N_2024,N_2132);
or U3353 (N_3353,N_2641,N_2609);
and U3354 (N_3354,N_2670,N_2995);
nand U3355 (N_3355,N_2713,N_2683);
or U3356 (N_3356,N_2317,N_2261);
nor U3357 (N_3357,N_2198,N_2709);
nand U3358 (N_3358,N_2715,N_2703);
and U3359 (N_3359,N_2094,N_2353);
and U3360 (N_3360,N_2800,N_2887);
nand U3361 (N_3361,N_2787,N_2110);
nand U3362 (N_3362,N_2184,N_2107);
or U3363 (N_3363,N_2439,N_2471);
or U3364 (N_3364,N_2783,N_2238);
nor U3365 (N_3365,N_2748,N_2310);
and U3366 (N_3366,N_2511,N_2460);
and U3367 (N_3367,N_2489,N_2571);
and U3368 (N_3368,N_2660,N_2224);
nand U3369 (N_3369,N_2021,N_2309);
or U3370 (N_3370,N_2124,N_2885);
and U3371 (N_3371,N_2263,N_2498);
nand U3372 (N_3372,N_2515,N_2930);
nand U3373 (N_3373,N_2939,N_2664);
nand U3374 (N_3374,N_2983,N_2087);
or U3375 (N_3375,N_2626,N_2482);
or U3376 (N_3376,N_2905,N_2599);
and U3377 (N_3377,N_2702,N_2425);
nor U3378 (N_3378,N_2699,N_2440);
and U3379 (N_3379,N_2401,N_2424);
or U3380 (N_3380,N_2882,N_2162);
nand U3381 (N_3381,N_2866,N_2384);
nand U3382 (N_3382,N_2678,N_2366);
and U3383 (N_3383,N_2510,N_2027);
and U3384 (N_3384,N_2030,N_2050);
nand U3385 (N_3385,N_2134,N_2806);
nand U3386 (N_3386,N_2398,N_2484);
and U3387 (N_3387,N_2119,N_2029);
nand U3388 (N_3388,N_2501,N_2307);
nor U3389 (N_3389,N_2109,N_2104);
nand U3390 (N_3390,N_2299,N_2696);
or U3391 (N_3391,N_2951,N_2878);
nand U3392 (N_3392,N_2601,N_2765);
nor U3393 (N_3393,N_2667,N_2348);
or U3394 (N_3394,N_2595,N_2014);
nand U3395 (N_3395,N_2717,N_2970);
or U3396 (N_3396,N_2594,N_2239);
and U3397 (N_3397,N_2937,N_2805);
or U3398 (N_3398,N_2009,N_2163);
nor U3399 (N_3399,N_2567,N_2801);
nor U3400 (N_3400,N_2570,N_2953);
and U3401 (N_3401,N_2598,N_2076);
nor U3402 (N_3402,N_2834,N_2754);
or U3403 (N_3403,N_2320,N_2903);
and U3404 (N_3404,N_2298,N_2042);
nand U3405 (N_3405,N_2389,N_2148);
nand U3406 (N_3406,N_2847,N_2542);
nand U3407 (N_3407,N_2974,N_2714);
and U3408 (N_3408,N_2558,N_2007);
nand U3409 (N_3409,N_2115,N_2578);
nor U3410 (N_3410,N_2436,N_2602);
and U3411 (N_3411,N_2458,N_2175);
or U3412 (N_3412,N_2874,N_2096);
nor U3413 (N_3413,N_2186,N_2390);
or U3414 (N_3414,N_2070,N_2826);
nand U3415 (N_3415,N_2213,N_2687);
and U3416 (N_3416,N_2149,N_2587);
nor U3417 (N_3417,N_2228,N_2491);
nand U3418 (N_3418,N_2923,N_2729);
and U3419 (N_3419,N_2472,N_2745);
or U3420 (N_3420,N_2693,N_2483);
nor U3421 (N_3421,N_2931,N_2531);
nand U3422 (N_3422,N_2459,N_2394);
nand U3423 (N_3423,N_2651,N_2507);
or U3424 (N_3424,N_2019,N_2285);
or U3425 (N_3425,N_2634,N_2043);
nand U3426 (N_3426,N_2827,N_2973);
nand U3427 (N_3427,N_2768,N_2015);
nand U3428 (N_3428,N_2861,N_2689);
nand U3429 (N_3429,N_2028,N_2323);
nor U3430 (N_3430,N_2979,N_2435);
or U3431 (N_3431,N_2002,N_2761);
nand U3432 (N_3432,N_2118,N_2249);
nand U3433 (N_3433,N_2867,N_2793);
or U3434 (N_3434,N_2958,N_2445);
or U3435 (N_3435,N_2147,N_2725);
nand U3436 (N_3436,N_2291,N_2138);
and U3437 (N_3437,N_2665,N_2041);
nor U3438 (N_3438,N_2766,N_2648);
nor U3439 (N_3439,N_2814,N_2414);
and U3440 (N_3440,N_2821,N_2860);
and U3441 (N_3441,N_2652,N_2084);
nand U3442 (N_3442,N_2111,N_2135);
or U3443 (N_3443,N_2064,N_2001);
or U3444 (N_3444,N_2112,N_2823);
nand U3445 (N_3445,N_2723,N_2038);
and U3446 (N_3446,N_2895,N_2209);
nand U3447 (N_3447,N_2208,N_2057);
or U3448 (N_3448,N_2174,N_2591);
xnor U3449 (N_3449,N_2871,N_2738);
nor U3450 (N_3450,N_2962,N_2617);
xnor U3451 (N_3451,N_2287,N_2596);
and U3452 (N_3452,N_2402,N_2999);
or U3453 (N_3453,N_2146,N_2080);
and U3454 (N_3454,N_2352,N_2006);
or U3455 (N_3455,N_2881,N_2187);
nand U3456 (N_3456,N_2642,N_2779);
nand U3457 (N_3457,N_2288,N_2536);
nor U3458 (N_3458,N_2380,N_2509);
nand U3459 (N_3459,N_2764,N_2127);
nor U3460 (N_3460,N_2528,N_2926);
nand U3461 (N_3461,N_2540,N_2447);
or U3462 (N_3462,N_2160,N_2662);
nand U3463 (N_3463,N_2719,N_2549);
nor U3464 (N_3464,N_2817,N_2855);
and U3465 (N_3465,N_2969,N_2474);
or U3466 (N_3466,N_2280,N_2675);
nor U3467 (N_3467,N_2647,N_2673);
nand U3468 (N_3468,N_2868,N_2193);
nand U3469 (N_3469,N_2657,N_2448);
and U3470 (N_3470,N_2853,N_2813);
nor U3471 (N_3471,N_2756,N_2464);
nor U3472 (N_3472,N_2551,N_2264);
or U3473 (N_3473,N_2383,N_2059);
and U3474 (N_3474,N_2420,N_2656);
nor U3475 (N_3475,N_2321,N_2960);
or U3476 (N_3476,N_2103,N_2934);
and U3477 (N_3477,N_2741,N_2746);
and U3478 (N_3478,N_2576,N_2572);
nand U3479 (N_3479,N_2844,N_2499);
nand U3480 (N_3480,N_2226,N_2618);
and U3481 (N_3481,N_2141,N_2235);
or U3482 (N_3482,N_2988,N_2478);
or U3483 (N_3483,N_2190,N_2924);
nor U3484 (N_3484,N_2575,N_2695);
or U3485 (N_3485,N_2266,N_2105);
nand U3486 (N_3486,N_2256,N_2770);
nor U3487 (N_3487,N_2669,N_2897);
nor U3488 (N_3488,N_2523,N_2337);
nor U3489 (N_3489,N_2416,N_2338);
nor U3490 (N_3490,N_2358,N_2789);
xnor U3491 (N_3491,N_2302,N_2769);
nand U3492 (N_3492,N_2170,N_2269);
nand U3493 (N_3493,N_2997,N_2803);
nand U3494 (N_3494,N_2896,N_2062);
xnor U3495 (N_3495,N_2701,N_2753);
nand U3496 (N_3496,N_2047,N_2131);
nor U3497 (N_3497,N_2250,N_2365);
nor U3498 (N_3498,N_2680,N_2967);
nor U3499 (N_3499,N_2532,N_2279);
or U3500 (N_3500,N_2537,N_2966);
or U3501 (N_3501,N_2746,N_2027);
nand U3502 (N_3502,N_2404,N_2433);
and U3503 (N_3503,N_2259,N_2001);
and U3504 (N_3504,N_2024,N_2756);
nor U3505 (N_3505,N_2833,N_2118);
and U3506 (N_3506,N_2522,N_2923);
nor U3507 (N_3507,N_2990,N_2089);
nor U3508 (N_3508,N_2437,N_2383);
or U3509 (N_3509,N_2814,N_2717);
xnor U3510 (N_3510,N_2282,N_2308);
nor U3511 (N_3511,N_2204,N_2345);
nand U3512 (N_3512,N_2285,N_2333);
nor U3513 (N_3513,N_2812,N_2981);
nand U3514 (N_3514,N_2497,N_2407);
nand U3515 (N_3515,N_2730,N_2990);
nor U3516 (N_3516,N_2672,N_2075);
or U3517 (N_3517,N_2732,N_2334);
or U3518 (N_3518,N_2452,N_2249);
or U3519 (N_3519,N_2090,N_2642);
or U3520 (N_3520,N_2422,N_2945);
nand U3521 (N_3521,N_2622,N_2278);
and U3522 (N_3522,N_2919,N_2882);
or U3523 (N_3523,N_2644,N_2456);
nand U3524 (N_3524,N_2835,N_2961);
nor U3525 (N_3525,N_2504,N_2789);
and U3526 (N_3526,N_2475,N_2319);
nor U3527 (N_3527,N_2777,N_2595);
nor U3528 (N_3528,N_2942,N_2639);
or U3529 (N_3529,N_2215,N_2472);
nand U3530 (N_3530,N_2318,N_2288);
or U3531 (N_3531,N_2633,N_2859);
nor U3532 (N_3532,N_2397,N_2765);
nor U3533 (N_3533,N_2487,N_2729);
nand U3534 (N_3534,N_2677,N_2449);
and U3535 (N_3535,N_2010,N_2575);
or U3536 (N_3536,N_2166,N_2203);
and U3537 (N_3537,N_2135,N_2839);
nor U3538 (N_3538,N_2580,N_2594);
or U3539 (N_3539,N_2021,N_2203);
or U3540 (N_3540,N_2506,N_2664);
nand U3541 (N_3541,N_2385,N_2740);
and U3542 (N_3542,N_2855,N_2905);
nand U3543 (N_3543,N_2928,N_2400);
nor U3544 (N_3544,N_2417,N_2529);
and U3545 (N_3545,N_2136,N_2416);
nor U3546 (N_3546,N_2971,N_2943);
nand U3547 (N_3547,N_2712,N_2886);
and U3548 (N_3548,N_2881,N_2898);
nand U3549 (N_3549,N_2284,N_2655);
nor U3550 (N_3550,N_2779,N_2754);
nand U3551 (N_3551,N_2341,N_2658);
nand U3552 (N_3552,N_2119,N_2298);
nor U3553 (N_3553,N_2498,N_2400);
nor U3554 (N_3554,N_2435,N_2078);
nand U3555 (N_3555,N_2240,N_2406);
nor U3556 (N_3556,N_2399,N_2804);
nor U3557 (N_3557,N_2049,N_2075);
nand U3558 (N_3558,N_2091,N_2449);
or U3559 (N_3559,N_2599,N_2130);
or U3560 (N_3560,N_2669,N_2559);
nor U3561 (N_3561,N_2074,N_2860);
nand U3562 (N_3562,N_2660,N_2493);
or U3563 (N_3563,N_2925,N_2040);
and U3564 (N_3564,N_2657,N_2852);
or U3565 (N_3565,N_2764,N_2697);
and U3566 (N_3566,N_2777,N_2148);
or U3567 (N_3567,N_2467,N_2961);
xnor U3568 (N_3568,N_2109,N_2558);
nor U3569 (N_3569,N_2534,N_2266);
and U3570 (N_3570,N_2277,N_2213);
or U3571 (N_3571,N_2880,N_2092);
nor U3572 (N_3572,N_2159,N_2118);
nor U3573 (N_3573,N_2463,N_2188);
and U3574 (N_3574,N_2597,N_2339);
nand U3575 (N_3575,N_2012,N_2007);
or U3576 (N_3576,N_2264,N_2627);
nand U3577 (N_3577,N_2839,N_2497);
xnor U3578 (N_3578,N_2320,N_2224);
or U3579 (N_3579,N_2084,N_2419);
nand U3580 (N_3580,N_2697,N_2105);
and U3581 (N_3581,N_2866,N_2265);
or U3582 (N_3582,N_2296,N_2427);
and U3583 (N_3583,N_2858,N_2432);
nand U3584 (N_3584,N_2149,N_2092);
nand U3585 (N_3585,N_2464,N_2624);
or U3586 (N_3586,N_2165,N_2775);
nor U3587 (N_3587,N_2750,N_2799);
nand U3588 (N_3588,N_2726,N_2080);
or U3589 (N_3589,N_2332,N_2695);
nand U3590 (N_3590,N_2690,N_2397);
or U3591 (N_3591,N_2320,N_2095);
or U3592 (N_3592,N_2415,N_2346);
or U3593 (N_3593,N_2662,N_2636);
nand U3594 (N_3594,N_2384,N_2610);
nand U3595 (N_3595,N_2723,N_2607);
and U3596 (N_3596,N_2904,N_2270);
nand U3597 (N_3597,N_2615,N_2990);
or U3598 (N_3598,N_2452,N_2439);
nor U3599 (N_3599,N_2105,N_2623);
and U3600 (N_3600,N_2495,N_2736);
and U3601 (N_3601,N_2518,N_2583);
nor U3602 (N_3602,N_2518,N_2502);
nor U3603 (N_3603,N_2383,N_2163);
or U3604 (N_3604,N_2537,N_2384);
nor U3605 (N_3605,N_2124,N_2102);
xnor U3606 (N_3606,N_2592,N_2644);
and U3607 (N_3607,N_2589,N_2879);
nor U3608 (N_3608,N_2959,N_2929);
xnor U3609 (N_3609,N_2870,N_2828);
nand U3610 (N_3610,N_2604,N_2373);
and U3611 (N_3611,N_2792,N_2062);
and U3612 (N_3612,N_2614,N_2612);
nand U3613 (N_3613,N_2915,N_2335);
nor U3614 (N_3614,N_2542,N_2969);
nor U3615 (N_3615,N_2452,N_2936);
nor U3616 (N_3616,N_2754,N_2916);
or U3617 (N_3617,N_2236,N_2361);
or U3618 (N_3618,N_2372,N_2050);
nor U3619 (N_3619,N_2217,N_2204);
or U3620 (N_3620,N_2441,N_2578);
or U3621 (N_3621,N_2376,N_2887);
or U3622 (N_3622,N_2884,N_2470);
and U3623 (N_3623,N_2815,N_2128);
nand U3624 (N_3624,N_2439,N_2420);
nor U3625 (N_3625,N_2485,N_2733);
and U3626 (N_3626,N_2939,N_2404);
nand U3627 (N_3627,N_2864,N_2363);
nand U3628 (N_3628,N_2091,N_2160);
and U3629 (N_3629,N_2620,N_2019);
or U3630 (N_3630,N_2654,N_2083);
or U3631 (N_3631,N_2916,N_2902);
nand U3632 (N_3632,N_2609,N_2788);
nand U3633 (N_3633,N_2669,N_2272);
nand U3634 (N_3634,N_2865,N_2224);
nand U3635 (N_3635,N_2258,N_2796);
nor U3636 (N_3636,N_2962,N_2216);
or U3637 (N_3637,N_2098,N_2925);
nor U3638 (N_3638,N_2379,N_2548);
and U3639 (N_3639,N_2382,N_2994);
nand U3640 (N_3640,N_2405,N_2893);
and U3641 (N_3641,N_2022,N_2418);
nor U3642 (N_3642,N_2540,N_2773);
nor U3643 (N_3643,N_2926,N_2134);
and U3644 (N_3644,N_2905,N_2285);
nor U3645 (N_3645,N_2667,N_2551);
or U3646 (N_3646,N_2912,N_2261);
nor U3647 (N_3647,N_2183,N_2984);
or U3648 (N_3648,N_2424,N_2539);
or U3649 (N_3649,N_2533,N_2790);
nor U3650 (N_3650,N_2151,N_2821);
and U3651 (N_3651,N_2555,N_2780);
nand U3652 (N_3652,N_2058,N_2442);
nor U3653 (N_3653,N_2345,N_2073);
nand U3654 (N_3654,N_2648,N_2231);
nand U3655 (N_3655,N_2162,N_2827);
or U3656 (N_3656,N_2676,N_2269);
or U3657 (N_3657,N_2149,N_2700);
or U3658 (N_3658,N_2900,N_2015);
or U3659 (N_3659,N_2482,N_2104);
and U3660 (N_3660,N_2363,N_2955);
or U3661 (N_3661,N_2183,N_2952);
nor U3662 (N_3662,N_2002,N_2324);
nand U3663 (N_3663,N_2828,N_2535);
nor U3664 (N_3664,N_2065,N_2318);
nand U3665 (N_3665,N_2012,N_2374);
nor U3666 (N_3666,N_2067,N_2831);
nand U3667 (N_3667,N_2358,N_2079);
and U3668 (N_3668,N_2256,N_2931);
nand U3669 (N_3669,N_2011,N_2637);
nor U3670 (N_3670,N_2862,N_2695);
and U3671 (N_3671,N_2135,N_2952);
or U3672 (N_3672,N_2042,N_2287);
or U3673 (N_3673,N_2249,N_2207);
and U3674 (N_3674,N_2640,N_2004);
and U3675 (N_3675,N_2101,N_2429);
or U3676 (N_3676,N_2707,N_2901);
nand U3677 (N_3677,N_2298,N_2055);
nor U3678 (N_3678,N_2445,N_2036);
nor U3679 (N_3679,N_2077,N_2439);
and U3680 (N_3680,N_2569,N_2944);
nand U3681 (N_3681,N_2976,N_2466);
nor U3682 (N_3682,N_2412,N_2175);
nor U3683 (N_3683,N_2403,N_2755);
or U3684 (N_3684,N_2523,N_2081);
or U3685 (N_3685,N_2499,N_2911);
and U3686 (N_3686,N_2072,N_2404);
and U3687 (N_3687,N_2790,N_2629);
nor U3688 (N_3688,N_2508,N_2775);
or U3689 (N_3689,N_2210,N_2415);
nand U3690 (N_3690,N_2504,N_2498);
and U3691 (N_3691,N_2039,N_2263);
nand U3692 (N_3692,N_2500,N_2610);
and U3693 (N_3693,N_2559,N_2073);
nor U3694 (N_3694,N_2246,N_2259);
nor U3695 (N_3695,N_2047,N_2630);
and U3696 (N_3696,N_2303,N_2082);
nand U3697 (N_3697,N_2025,N_2841);
nand U3698 (N_3698,N_2134,N_2363);
or U3699 (N_3699,N_2368,N_2559);
nand U3700 (N_3700,N_2641,N_2988);
nand U3701 (N_3701,N_2344,N_2555);
nor U3702 (N_3702,N_2124,N_2616);
nor U3703 (N_3703,N_2908,N_2024);
and U3704 (N_3704,N_2988,N_2814);
or U3705 (N_3705,N_2172,N_2400);
nor U3706 (N_3706,N_2816,N_2670);
nor U3707 (N_3707,N_2305,N_2431);
and U3708 (N_3708,N_2164,N_2008);
nor U3709 (N_3709,N_2928,N_2557);
nor U3710 (N_3710,N_2067,N_2442);
nand U3711 (N_3711,N_2080,N_2359);
nand U3712 (N_3712,N_2429,N_2481);
nor U3713 (N_3713,N_2460,N_2666);
nor U3714 (N_3714,N_2029,N_2140);
nand U3715 (N_3715,N_2502,N_2897);
or U3716 (N_3716,N_2630,N_2950);
nand U3717 (N_3717,N_2245,N_2897);
nor U3718 (N_3718,N_2291,N_2170);
or U3719 (N_3719,N_2154,N_2263);
or U3720 (N_3720,N_2229,N_2152);
and U3721 (N_3721,N_2889,N_2704);
and U3722 (N_3722,N_2073,N_2931);
and U3723 (N_3723,N_2751,N_2290);
and U3724 (N_3724,N_2845,N_2678);
nand U3725 (N_3725,N_2546,N_2034);
or U3726 (N_3726,N_2546,N_2722);
nand U3727 (N_3727,N_2134,N_2215);
or U3728 (N_3728,N_2835,N_2182);
and U3729 (N_3729,N_2189,N_2339);
nor U3730 (N_3730,N_2673,N_2840);
nand U3731 (N_3731,N_2694,N_2451);
nor U3732 (N_3732,N_2865,N_2259);
or U3733 (N_3733,N_2298,N_2397);
and U3734 (N_3734,N_2216,N_2066);
nand U3735 (N_3735,N_2250,N_2105);
nand U3736 (N_3736,N_2053,N_2626);
nand U3737 (N_3737,N_2542,N_2872);
nor U3738 (N_3738,N_2099,N_2994);
and U3739 (N_3739,N_2611,N_2648);
nand U3740 (N_3740,N_2507,N_2616);
or U3741 (N_3741,N_2396,N_2426);
and U3742 (N_3742,N_2392,N_2408);
nor U3743 (N_3743,N_2284,N_2398);
and U3744 (N_3744,N_2071,N_2944);
nor U3745 (N_3745,N_2670,N_2722);
or U3746 (N_3746,N_2748,N_2918);
or U3747 (N_3747,N_2648,N_2065);
or U3748 (N_3748,N_2621,N_2578);
and U3749 (N_3749,N_2749,N_2640);
or U3750 (N_3750,N_2932,N_2453);
or U3751 (N_3751,N_2798,N_2800);
nand U3752 (N_3752,N_2851,N_2382);
and U3753 (N_3753,N_2945,N_2764);
or U3754 (N_3754,N_2205,N_2939);
or U3755 (N_3755,N_2385,N_2652);
nor U3756 (N_3756,N_2655,N_2887);
nor U3757 (N_3757,N_2068,N_2879);
and U3758 (N_3758,N_2708,N_2003);
or U3759 (N_3759,N_2041,N_2785);
nor U3760 (N_3760,N_2353,N_2570);
nor U3761 (N_3761,N_2694,N_2766);
nand U3762 (N_3762,N_2351,N_2525);
nor U3763 (N_3763,N_2649,N_2978);
nor U3764 (N_3764,N_2458,N_2815);
nand U3765 (N_3765,N_2195,N_2553);
or U3766 (N_3766,N_2545,N_2804);
or U3767 (N_3767,N_2639,N_2732);
nand U3768 (N_3768,N_2831,N_2323);
or U3769 (N_3769,N_2762,N_2527);
nand U3770 (N_3770,N_2183,N_2583);
and U3771 (N_3771,N_2583,N_2248);
nor U3772 (N_3772,N_2043,N_2905);
nand U3773 (N_3773,N_2073,N_2016);
and U3774 (N_3774,N_2163,N_2007);
or U3775 (N_3775,N_2878,N_2398);
nor U3776 (N_3776,N_2171,N_2824);
xor U3777 (N_3777,N_2462,N_2725);
nor U3778 (N_3778,N_2936,N_2056);
and U3779 (N_3779,N_2141,N_2778);
and U3780 (N_3780,N_2141,N_2596);
nand U3781 (N_3781,N_2518,N_2851);
or U3782 (N_3782,N_2463,N_2977);
and U3783 (N_3783,N_2381,N_2452);
nand U3784 (N_3784,N_2796,N_2839);
or U3785 (N_3785,N_2888,N_2353);
nand U3786 (N_3786,N_2516,N_2820);
nand U3787 (N_3787,N_2045,N_2486);
nand U3788 (N_3788,N_2068,N_2278);
or U3789 (N_3789,N_2353,N_2614);
or U3790 (N_3790,N_2094,N_2132);
or U3791 (N_3791,N_2837,N_2189);
nor U3792 (N_3792,N_2783,N_2152);
nor U3793 (N_3793,N_2334,N_2012);
and U3794 (N_3794,N_2713,N_2952);
and U3795 (N_3795,N_2431,N_2556);
nor U3796 (N_3796,N_2126,N_2666);
nor U3797 (N_3797,N_2518,N_2834);
or U3798 (N_3798,N_2602,N_2297);
nand U3799 (N_3799,N_2841,N_2604);
nor U3800 (N_3800,N_2506,N_2383);
nor U3801 (N_3801,N_2774,N_2558);
and U3802 (N_3802,N_2074,N_2453);
nor U3803 (N_3803,N_2038,N_2983);
nor U3804 (N_3804,N_2527,N_2540);
nor U3805 (N_3805,N_2430,N_2976);
nor U3806 (N_3806,N_2557,N_2908);
or U3807 (N_3807,N_2980,N_2450);
or U3808 (N_3808,N_2745,N_2788);
nor U3809 (N_3809,N_2040,N_2932);
nor U3810 (N_3810,N_2239,N_2690);
and U3811 (N_3811,N_2378,N_2829);
or U3812 (N_3812,N_2557,N_2942);
nor U3813 (N_3813,N_2058,N_2663);
or U3814 (N_3814,N_2367,N_2876);
or U3815 (N_3815,N_2347,N_2988);
nand U3816 (N_3816,N_2711,N_2572);
or U3817 (N_3817,N_2912,N_2008);
nor U3818 (N_3818,N_2784,N_2704);
and U3819 (N_3819,N_2026,N_2124);
or U3820 (N_3820,N_2994,N_2670);
and U3821 (N_3821,N_2771,N_2896);
or U3822 (N_3822,N_2472,N_2608);
and U3823 (N_3823,N_2593,N_2397);
or U3824 (N_3824,N_2144,N_2242);
and U3825 (N_3825,N_2525,N_2652);
nand U3826 (N_3826,N_2047,N_2077);
or U3827 (N_3827,N_2491,N_2846);
and U3828 (N_3828,N_2249,N_2545);
or U3829 (N_3829,N_2089,N_2693);
nand U3830 (N_3830,N_2826,N_2174);
and U3831 (N_3831,N_2426,N_2924);
nand U3832 (N_3832,N_2012,N_2473);
and U3833 (N_3833,N_2660,N_2612);
or U3834 (N_3834,N_2552,N_2660);
and U3835 (N_3835,N_2970,N_2046);
or U3836 (N_3836,N_2244,N_2402);
nor U3837 (N_3837,N_2761,N_2357);
xor U3838 (N_3838,N_2252,N_2876);
or U3839 (N_3839,N_2779,N_2882);
nor U3840 (N_3840,N_2209,N_2711);
or U3841 (N_3841,N_2039,N_2429);
and U3842 (N_3842,N_2800,N_2097);
or U3843 (N_3843,N_2533,N_2762);
or U3844 (N_3844,N_2597,N_2199);
or U3845 (N_3845,N_2609,N_2298);
and U3846 (N_3846,N_2148,N_2873);
and U3847 (N_3847,N_2431,N_2651);
and U3848 (N_3848,N_2101,N_2760);
and U3849 (N_3849,N_2258,N_2770);
nand U3850 (N_3850,N_2443,N_2670);
and U3851 (N_3851,N_2143,N_2272);
nor U3852 (N_3852,N_2974,N_2598);
nand U3853 (N_3853,N_2406,N_2782);
nor U3854 (N_3854,N_2729,N_2434);
and U3855 (N_3855,N_2215,N_2891);
nor U3856 (N_3856,N_2288,N_2369);
and U3857 (N_3857,N_2950,N_2031);
and U3858 (N_3858,N_2000,N_2670);
nor U3859 (N_3859,N_2814,N_2523);
nand U3860 (N_3860,N_2300,N_2228);
nor U3861 (N_3861,N_2285,N_2790);
nor U3862 (N_3862,N_2458,N_2528);
nand U3863 (N_3863,N_2387,N_2067);
nor U3864 (N_3864,N_2911,N_2443);
nand U3865 (N_3865,N_2737,N_2425);
nor U3866 (N_3866,N_2602,N_2151);
nor U3867 (N_3867,N_2469,N_2672);
and U3868 (N_3868,N_2339,N_2644);
nand U3869 (N_3869,N_2559,N_2953);
or U3870 (N_3870,N_2883,N_2595);
nor U3871 (N_3871,N_2706,N_2699);
nand U3872 (N_3872,N_2713,N_2673);
and U3873 (N_3873,N_2113,N_2078);
or U3874 (N_3874,N_2003,N_2817);
nand U3875 (N_3875,N_2339,N_2990);
or U3876 (N_3876,N_2337,N_2129);
nand U3877 (N_3877,N_2720,N_2933);
and U3878 (N_3878,N_2346,N_2398);
or U3879 (N_3879,N_2934,N_2836);
and U3880 (N_3880,N_2186,N_2286);
and U3881 (N_3881,N_2641,N_2784);
nand U3882 (N_3882,N_2653,N_2452);
or U3883 (N_3883,N_2445,N_2264);
or U3884 (N_3884,N_2804,N_2244);
or U3885 (N_3885,N_2041,N_2318);
or U3886 (N_3886,N_2723,N_2238);
and U3887 (N_3887,N_2469,N_2487);
nor U3888 (N_3888,N_2638,N_2853);
or U3889 (N_3889,N_2513,N_2346);
or U3890 (N_3890,N_2629,N_2154);
and U3891 (N_3891,N_2031,N_2361);
and U3892 (N_3892,N_2841,N_2458);
or U3893 (N_3893,N_2392,N_2005);
nor U3894 (N_3894,N_2728,N_2885);
nor U3895 (N_3895,N_2111,N_2521);
or U3896 (N_3896,N_2364,N_2198);
or U3897 (N_3897,N_2423,N_2023);
nand U3898 (N_3898,N_2174,N_2892);
nand U3899 (N_3899,N_2579,N_2287);
and U3900 (N_3900,N_2573,N_2450);
nand U3901 (N_3901,N_2440,N_2996);
nand U3902 (N_3902,N_2930,N_2801);
and U3903 (N_3903,N_2826,N_2400);
nand U3904 (N_3904,N_2113,N_2095);
nor U3905 (N_3905,N_2950,N_2982);
and U3906 (N_3906,N_2892,N_2893);
and U3907 (N_3907,N_2735,N_2541);
nand U3908 (N_3908,N_2783,N_2822);
nand U3909 (N_3909,N_2242,N_2152);
nand U3910 (N_3910,N_2262,N_2812);
and U3911 (N_3911,N_2383,N_2385);
or U3912 (N_3912,N_2839,N_2106);
and U3913 (N_3913,N_2730,N_2094);
and U3914 (N_3914,N_2502,N_2687);
nor U3915 (N_3915,N_2746,N_2072);
nand U3916 (N_3916,N_2053,N_2165);
nand U3917 (N_3917,N_2740,N_2421);
and U3918 (N_3918,N_2710,N_2891);
and U3919 (N_3919,N_2854,N_2609);
nand U3920 (N_3920,N_2607,N_2480);
and U3921 (N_3921,N_2297,N_2290);
nand U3922 (N_3922,N_2651,N_2353);
or U3923 (N_3923,N_2606,N_2544);
and U3924 (N_3924,N_2265,N_2454);
or U3925 (N_3925,N_2950,N_2101);
and U3926 (N_3926,N_2484,N_2282);
and U3927 (N_3927,N_2688,N_2716);
or U3928 (N_3928,N_2528,N_2759);
nor U3929 (N_3929,N_2803,N_2366);
nand U3930 (N_3930,N_2190,N_2041);
nor U3931 (N_3931,N_2977,N_2279);
and U3932 (N_3932,N_2884,N_2585);
or U3933 (N_3933,N_2017,N_2601);
nor U3934 (N_3934,N_2109,N_2514);
or U3935 (N_3935,N_2122,N_2588);
and U3936 (N_3936,N_2154,N_2442);
nor U3937 (N_3937,N_2706,N_2138);
or U3938 (N_3938,N_2155,N_2546);
or U3939 (N_3939,N_2972,N_2047);
and U3940 (N_3940,N_2379,N_2673);
and U3941 (N_3941,N_2804,N_2873);
and U3942 (N_3942,N_2248,N_2754);
and U3943 (N_3943,N_2610,N_2767);
nand U3944 (N_3944,N_2062,N_2390);
nor U3945 (N_3945,N_2393,N_2593);
or U3946 (N_3946,N_2720,N_2048);
xor U3947 (N_3947,N_2862,N_2586);
nor U3948 (N_3948,N_2682,N_2406);
and U3949 (N_3949,N_2673,N_2402);
or U3950 (N_3950,N_2003,N_2374);
nand U3951 (N_3951,N_2620,N_2832);
xor U3952 (N_3952,N_2296,N_2531);
and U3953 (N_3953,N_2521,N_2088);
nor U3954 (N_3954,N_2544,N_2304);
nor U3955 (N_3955,N_2626,N_2951);
nand U3956 (N_3956,N_2216,N_2705);
nor U3957 (N_3957,N_2444,N_2361);
or U3958 (N_3958,N_2581,N_2771);
and U3959 (N_3959,N_2691,N_2302);
and U3960 (N_3960,N_2289,N_2695);
xnor U3961 (N_3961,N_2991,N_2959);
or U3962 (N_3962,N_2108,N_2976);
and U3963 (N_3963,N_2327,N_2013);
nand U3964 (N_3964,N_2749,N_2975);
and U3965 (N_3965,N_2729,N_2762);
or U3966 (N_3966,N_2808,N_2516);
or U3967 (N_3967,N_2689,N_2920);
nand U3968 (N_3968,N_2594,N_2040);
or U3969 (N_3969,N_2948,N_2555);
nand U3970 (N_3970,N_2127,N_2666);
and U3971 (N_3971,N_2479,N_2662);
or U3972 (N_3972,N_2223,N_2420);
nor U3973 (N_3973,N_2627,N_2464);
and U3974 (N_3974,N_2256,N_2719);
and U3975 (N_3975,N_2617,N_2340);
nor U3976 (N_3976,N_2795,N_2933);
and U3977 (N_3977,N_2520,N_2869);
nand U3978 (N_3978,N_2441,N_2604);
nor U3979 (N_3979,N_2617,N_2800);
nor U3980 (N_3980,N_2379,N_2459);
nor U3981 (N_3981,N_2583,N_2337);
nand U3982 (N_3982,N_2034,N_2949);
nor U3983 (N_3983,N_2566,N_2404);
or U3984 (N_3984,N_2886,N_2473);
nand U3985 (N_3985,N_2730,N_2396);
nor U3986 (N_3986,N_2336,N_2239);
and U3987 (N_3987,N_2977,N_2814);
and U3988 (N_3988,N_2447,N_2282);
nor U3989 (N_3989,N_2377,N_2115);
nand U3990 (N_3990,N_2731,N_2317);
and U3991 (N_3991,N_2788,N_2930);
nand U3992 (N_3992,N_2582,N_2598);
nand U3993 (N_3993,N_2637,N_2473);
or U3994 (N_3994,N_2610,N_2736);
or U3995 (N_3995,N_2211,N_2768);
nand U3996 (N_3996,N_2419,N_2190);
and U3997 (N_3997,N_2143,N_2962);
and U3998 (N_3998,N_2590,N_2175);
or U3999 (N_3999,N_2962,N_2024);
and U4000 (N_4000,N_3731,N_3220);
nand U4001 (N_4001,N_3216,N_3133);
and U4002 (N_4002,N_3193,N_3494);
xor U4003 (N_4003,N_3088,N_3395);
nor U4004 (N_4004,N_3670,N_3944);
nor U4005 (N_4005,N_3111,N_3983);
and U4006 (N_4006,N_3744,N_3267);
or U4007 (N_4007,N_3376,N_3642);
or U4008 (N_4008,N_3257,N_3362);
and U4009 (N_4009,N_3072,N_3291);
nor U4010 (N_4010,N_3358,N_3471);
nor U4011 (N_4011,N_3755,N_3003);
nor U4012 (N_4012,N_3531,N_3977);
or U4013 (N_4013,N_3048,N_3852);
xnor U4014 (N_4014,N_3096,N_3971);
or U4015 (N_4015,N_3819,N_3951);
and U4016 (N_4016,N_3459,N_3488);
nor U4017 (N_4017,N_3209,N_3595);
or U4018 (N_4018,N_3312,N_3636);
nor U4019 (N_4019,N_3781,N_3136);
xnor U4020 (N_4020,N_3866,N_3876);
nor U4021 (N_4021,N_3094,N_3586);
nor U4022 (N_4022,N_3752,N_3184);
nand U4023 (N_4023,N_3310,N_3735);
nand U4024 (N_4024,N_3909,N_3380);
and U4025 (N_4025,N_3857,N_3101);
nand U4026 (N_4026,N_3299,N_3489);
nor U4027 (N_4027,N_3712,N_3198);
or U4028 (N_4028,N_3428,N_3192);
nor U4029 (N_4029,N_3073,N_3730);
or U4030 (N_4030,N_3972,N_3892);
and U4031 (N_4031,N_3577,N_3791);
and U4032 (N_4032,N_3848,N_3946);
and U4033 (N_4033,N_3913,N_3681);
and U4034 (N_4034,N_3068,N_3968);
and U4035 (N_4035,N_3254,N_3877);
or U4036 (N_4036,N_3130,N_3478);
nand U4037 (N_4037,N_3182,N_3527);
nor U4038 (N_4038,N_3979,N_3235);
or U4039 (N_4039,N_3328,N_3539);
and U4040 (N_4040,N_3483,N_3770);
or U4041 (N_4041,N_3701,N_3902);
xor U4042 (N_4042,N_3378,N_3695);
nand U4043 (N_4043,N_3637,N_3528);
nand U4044 (N_4044,N_3444,N_3896);
nor U4045 (N_4045,N_3274,N_3166);
or U4046 (N_4046,N_3202,N_3584);
nor U4047 (N_4047,N_3367,N_3954);
nand U4048 (N_4048,N_3861,N_3006);
or U4049 (N_4049,N_3596,N_3936);
or U4050 (N_4050,N_3980,N_3987);
nand U4051 (N_4051,N_3749,N_3524);
nand U4052 (N_4052,N_3967,N_3470);
nand U4053 (N_4053,N_3839,N_3827);
nor U4054 (N_4054,N_3425,N_3445);
or U4055 (N_4055,N_3141,N_3665);
and U4056 (N_4056,N_3052,N_3639);
and U4057 (N_4057,N_3806,N_3070);
nor U4058 (N_4058,N_3587,N_3846);
or U4059 (N_4059,N_3032,N_3122);
and U4060 (N_4060,N_3222,N_3423);
nor U4061 (N_4061,N_3958,N_3690);
nand U4062 (N_4062,N_3914,N_3700);
nor U4063 (N_4063,N_3903,N_3138);
xor U4064 (N_4064,N_3810,N_3245);
nor U4065 (N_4065,N_3982,N_3549);
and U4066 (N_4066,N_3789,N_3547);
and U4067 (N_4067,N_3939,N_3463);
nor U4068 (N_4068,N_3208,N_3104);
nor U4069 (N_4069,N_3634,N_3585);
nand U4070 (N_4070,N_3985,N_3994);
nor U4071 (N_4071,N_3809,N_3451);
or U4072 (N_4072,N_3273,N_3435);
nor U4073 (N_4073,N_3099,N_3760);
or U4074 (N_4074,N_3170,N_3793);
nand U4075 (N_4075,N_3575,N_3623);
nand U4076 (N_4076,N_3233,N_3414);
or U4077 (N_4077,N_3763,N_3685);
or U4078 (N_4078,N_3468,N_3895);
nand U4079 (N_4079,N_3777,N_3010);
or U4080 (N_4080,N_3128,N_3103);
nand U4081 (N_4081,N_3082,N_3662);
nor U4082 (N_4082,N_3276,N_3053);
or U4083 (N_4083,N_3785,N_3578);
and U4084 (N_4084,N_3106,N_3934);
and U4085 (N_4085,N_3297,N_3828);
nand U4086 (N_4086,N_3204,N_3616);
nor U4087 (N_4087,N_3945,N_3963);
nand U4088 (N_4088,N_3705,N_3013);
and U4089 (N_4089,N_3516,N_3338);
nand U4090 (N_4090,N_3645,N_3180);
or U4091 (N_4091,N_3379,N_3862);
nand U4092 (N_4092,N_3349,N_3869);
or U4093 (N_4093,N_3776,N_3477);
or U4094 (N_4094,N_3412,N_3237);
nand U4095 (N_4095,N_3829,N_3314);
and U4096 (N_4096,N_3692,N_3969);
and U4097 (N_4097,N_3990,N_3572);
and U4098 (N_4098,N_3837,N_3044);
nor U4099 (N_4099,N_3788,N_3309);
nand U4100 (N_4100,N_3461,N_3970);
nor U4101 (N_4101,N_3051,N_3105);
nand U4102 (N_4102,N_3600,N_3579);
and U4103 (N_4103,N_3456,N_3253);
nand U4104 (N_4104,N_3834,N_3455);
and U4105 (N_4105,N_3250,N_3519);
nand U4106 (N_4106,N_3300,N_3020);
and U4107 (N_4107,N_3880,N_3015);
and U4108 (N_4108,N_3200,N_3486);
and U4109 (N_4109,N_3675,N_3559);
and U4110 (N_4110,N_3065,N_3028);
and U4111 (N_4111,N_3038,N_3342);
nor U4112 (N_4112,N_3654,N_3322);
and U4113 (N_4113,N_3256,N_3050);
nor U4114 (N_4114,N_3437,N_3526);
and U4115 (N_4115,N_3707,N_3340);
nand U4116 (N_4116,N_3981,N_3125);
nor U4117 (N_4117,N_3782,N_3077);
nor U4118 (N_4118,N_3761,N_3074);
and U4119 (N_4119,N_3897,N_3404);
and U4120 (N_4120,N_3629,N_3830);
and U4121 (N_4121,N_3714,N_3567);
and U4122 (N_4122,N_3097,N_3541);
nor U4123 (N_4123,N_3239,N_3574);
or U4124 (N_4124,N_3870,N_3940);
and U4125 (N_4125,N_3917,N_3807);
and U4126 (N_4126,N_3368,N_3748);
nand U4127 (N_4127,N_3594,N_3004);
or U4128 (N_4128,N_3624,N_3668);
nand U4129 (N_4129,N_3792,N_3740);
and U4130 (N_4130,N_3049,N_3238);
nand U4131 (N_4131,N_3589,N_3509);
xor U4132 (N_4132,N_3382,N_3605);
nor U4133 (N_4133,N_3710,N_3150);
nand U4134 (N_4134,N_3635,N_3500);
and U4135 (N_4135,N_3953,N_3779);
nand U4136 (N_4136,N_3696,N_3446);
and U4137 (N_4137,N_3484,N_3080);
nand U4138 (N_4138,N_3139,N_3957);
nor U4139 (N_4139,N_3619,N_3821);
xnor U4140 (N_4140,N_3501,N_3568);
nor U4141 (N_4141,N_3177,N_3554);
or U4142 (N_4142,N_3986,N_3904);
nand U4143 (N_4143,N_3865,N_3129);
and U4144 (N_4144,N_3544,N_3910);
nor U4145 (N_4145,N_3132,N_3569);
nor U4146 (N_4146,N_3090,N_3984);
and U4147 (N_4147,N_3203,N_3289);
nand U4148 (N_4148,N_3001,N_3092);
nand U4149 (N_4149,N_3408,N_3115);
or U4150 (N_4150,N_3326,N_3534);
and U4151 (N_4151,N_3960,N_3604);
nand U4152 (N_4152,N_3964,N_3774);
nor U4153 (N_4153,N_3883,N_3346);
or U4154 (N_4154,N_3157,N_3306);
nor U4155 (N_4155,N_3186,N_3956);
and U4156 (N_4156,N_3337,N_3978);
nand U4157 (N_4157,N_3110,N_3504);
and U4158 (N_4158,N_3840,N_3523);
nand U4159 (N_4159,N_3369,N_3007);
and U4160 (N_4160,N_3440,N_3386);
or U4161 (N_4161,N_3113,N_3679);
nor U4162 (N_4162,N_3075,N_3796);
nor U4163 (N_4163,N_3268,N_3033);
and U4164 (N_4164,N_3330,N_3993);
nor U4165 (N_4165,N_3548,N_3421);
nor U4166 (N_4166,N_3264,N_3438);
and U4167 (N_4167,N_3546,N_3259);
or U4168 (N_4168,N_3609,N_3805);
or U4169 (N_4169,N_3581,N_3717);
or U4170 (N_4170,N_3027,N_3031);
or U4171 (N_4171,N_3000,N_3162);
or U4172 (N_4172,N_3699,N_3947);
nand U4173 (N_4173,N_3640,N_3304);
nand U4174 (N_4174,N_3089,N_3307);
or U4175 (N_4175,N_3244,N_3284);
or U4176 (N_4176,N_3508,N_3784);
or U4177 (N_4177,N_3801,N_3540);
nor U4178 (N_4178,N_3173,N_3511);
nand U4179 (N_4179,N_3148,N_3155);
nor U4180 (N_4180,N_3783,N_3227);
nand U4181 (N_4181,N_3551,N_3164);
nand U4182 (N_4182,N_3906,N_3171);
nand U4183 (N_4183,N_3773,N_3686);
or U4184 (N_4184,N_3641,N_3079);
nand U4185 (N_4185,N_3187,N_3556);
nor U4186 (N_4186,N_3364,N_3688);
nand U4187 (N_4187,N_3037,N_3287);
nor U4188 (N_4188,N_3948,N_3669);
nor U4189 (N_4189,N_3885,N_3725);
nand U4190 (N_4190,N_3659,N_3353);
and U4191 (N_4191,N_3067,N_3036);
nor U4192 (N_4192,N_3397,N_3413);
nand U4193 (N_4193,N_3905,N_3360);
nand U4194 (N_4194,N_3288,N_3281);
nor U4195 (N_4195,N_3927,N_3232);
nor U4196 (N_4196,N_3411,N_3592);
nor U4197 (N_4197,N_3429,N_3873);
or U4198 (N_4198,N_3814,N_3667);
or U4199 (N_4199,N_3453,N_3178);
nand U4200 (N_4200,N_3142,N_3794);
or U4201 (N_4201,N_3112,N_3974);
nand U4202 (N_4202,N_3197,N_3816);
nand U4203 (N_4203,N_3697,N_3263);
and U4204 (N_4204,N_3011,N_3343);
nand U4205 (N_4205,N_3201,N_3648);
nor U4206 (N_4206,N_3797,N_3618);
and U4207 (N_4207,N_3560,N_3406);
nor U4208 (N_4208,N_3709,N_3290);
nand U4209 (N_4209,N_3370,N_3884);
and U4210 (N_4210,N_3392,N_3998);
and U4211 (N_4211,N_3181,N_3098);
nor U4212 (N_4212,N_3599,N_3780);
or U4213 (N_4213,N_3704,N_3745);
nor U4214 (N_4214,N_3621,N_3510);
and U4215 (N_4215,N_3887,N_3506);
and U4216 (N_4216,N_3210,N_3664);
or U4217 (N_4217,N_3747,N_3179);
or U4218 (N_4218,N_3850,N_3331);
and U4219 (N_4219,N_3736,N_3039);
and U4220 (N_4220,N_3450,N_3663);
nand U4221 (N_4221,N_3499,N_3515);
nand U4222 (N_4222,N_3942,N_3924);
or U4223 (N_4223,N_3630,N_3485);
or U4224 (N_4224,N_3091,N_3283);
and U4225 (N_4225,N_3188,N_3348);
or U4226 (N_4226,N_3230,N_3441);
and U4227 (N_4227,N_3739,N_3085);
nand U4228 (N_4228,N_3512,N_3228);
or U4229 (N_4229,N_3847,N_3938);
and U4230 (N_4230,N_3661,N_3464);
and U4231 (N_4231,N_3279,N_3497);
nand U4232 (N_4232,N_3851,N_3107);
nor U4233 (N_4233,N_3992,N_3160);
nand U4234 (N_4234,N_3093,N_3633);
nor U4235 (N_4235,N_3874,N_3118);
nand U4236 (N_4236,N_3831,N_3625);
nor U4237 (N_4237,N_3009,N_3658);
or U4238 (N_4238,N_3260,N_3520);
or U4239 (N_4239,N_3632,N_3172);
and U4240 (N_4240,N_3057,N_3339);
nor U4241 (N_4241,N_3894,N_3466);
nand U4242 (N_4242,N_3900,N_3035);
nor U4243 (N_4243,N_3644,N_3550);
and U4244 (N_4244,N_3332,N_3126);
nand U4245 (N_4245,N_3682,N_3243);
or U4246 (N_4246,N_3590,N_3741);
and U4247 (N_4247,N_3860,N_3046);
nand U4248 (N_4248,N_3615,N_3071);
and U4249 (N_4249,N_3398,N_3858);
nand U4250 (N_4250,N_3918,N_3234);
and U4251 (N_4251,N_3875,N_3778);
nand U4252 (N_4252,N_3124,N_3989);
nand U4253 (N_4253,N_3365,N_3116);
or U4254 (N_4254,N_3651,N_3069);
or U4255 (N_4255,N_3350,N_3532);
nor U4256 (N_4256,N_3277,N_3389);
and U4257 (N_4257,N_3815,N_3347);
and U4258 (N_4258,N_3762,N_3912);
or U4259 (N_4259,N_3950,N_3812);
and U4260 (N_4260,N_3855,N_3649);
or U4261 (N_4261,N_3286,N_3390);
xnor U4262 (N_4262,N_3727,N_3562);
and U4263 (N_4263,N_3826,N_3418);
nand U4264 (N_4264,N_3147,N_3768);
or U4265 (N_4265,N_3564,N_3867);
nand U4266 (N_4266,N_3135,N_3465);
or U4267 (N_4267,N_3570,N_3481);
nand U4268 (N_4268,N_3375,N_3388);
nand U4269 (N_4269,N_3721,N_3236);
or U4270 (N_4270,N_3751,N_3996);
nand U4271 (N_4271,N_3156,N_3191);
nand U4272 (N_4272,N_3711,N_3282);
or U4273 (N_4273,N_3937,N_3545);
nand U4274 (N_4274,N_3305,N_3573);
nand U4275 (N_4275,N_3384,N_3225);
or U4276 (N_4276,N_3603,N_3034);
nor U4277 (N_4277,N_3008,N_3333);
nor U4278 (N_4278,N_3835,N_3566);
and U4279 (N_4279,N_3302,N_3943);
and U4280 (N_4280,N_3666,N_3716);
nand U4281 (N_4281,N_3401,N_3436);
or U4282 (N_4282,N_3657,N_3607);
nand U4283 (N_4283,N_3206,N_3507);
and U4284 (N_4284,N_3361,N_3928);
nand U4285 (N_4285,N_3026,N_3231);
nor U4286 (N_4286,N_3476,N_3102);
nor U4287 (N_4287,N_3647,N_3845);
and U4288 (N_4288,N_3643,N_3002);
or U4289 (N_4289,N_3726,N_3248);
nor U4290 (N_4290,N_3247,N_3355);
nor U4291 (N_4291,N_3680,N_3561);
nand U4292 (N_4292,N_3713,N_3315);
or U4293 (N_4293,N_3017,N_3399);
and U4294 (N_4294,N_3706,N_3676);
nand U4295 (N_4295,N_3822,N_3371);
or U4296 (N_4296,N_3285,N_3795);
nand U4297 (N_4297,N_3190,N_3652);
nor U4298 (N_4298,N_3498,N_3063);
nor U4299 (N_4299,N_3802,N_3757);
or U4300 (N_4300,N_3764,N_3759);
and U4301 (N_4301,N_3893,N_3134);
nor U4302 (N_4302,N_3374,N_3698);
and U4303 (N_4303,N_3854,N_3868);
nand U4304 (N_4304,N_3871,N_3505);
or U4305 (N_4305,N_3223,N_3872);
and U4306 (N_4306,N_3359,N_3750);
nand U4307 (N_4307,N_3167,N_3517);
and U4308 (N_4308,N_3813,N_3058);
or U4309 (N_4309,N_3427,N_3394);
xor U4310 (N_4310,N_3354,N_3023);
or U4311 (N_4311,N_3194,N_3426);
or U4312 (N_4312,N_3999,N_3321);
nand U4313 (N_4313,N_3415,N_3563);
nor U4314 (N_4314,N_3514,N_3765);
nand U4315 (N_4315,N_3753,N_3434);
or U4316 (N_4316,N_3448,N_3280);
or U4317 (N_4317,N_3976,N_3738);
nand U4318 (N_4318,N_3005,N_3258);
and U4319 (N_4319,N_3078,N_3702);
and U4320 (N_4320,N_3724,N_3732);
or U4321 (N_4321,N_3965,N_3055);
xor U4322 (N_4322,N_3327,N_3255);
and U4323 (N_4323,N_3215,N_3095);
or U4324 (N_4324,N_3195,N_3878);
nand U4325 (N_4325,N_3628,N_3811);
nand U4326 (N_4326,N_3149,N_3087);
nor U4327 (N_4327,N_3018,N_3185);
and U4328 (N_4328,N_3952,N_3703);
and U4329 (N_4329,N_3432,N_3298);
or U4330 (N_4330,N_3301,N_3966);
or U4331 (N_4331,N_3626,N_3422);
nor U4332 (N_4332,N_3121,N_3224);
or U4333 (N_4333,N_3317,N_3767);
and U4334 (N_4334,N_3955,N_3153);
and U4335 (N_4335,N_3061,N_3988);
nor U4336 (N_4336,N_3723,N_3932);
nor U4337 (N_4337,N_3059,N_3229);
nor U4338 (N_4338,N_3189,N_3687);
nand U4339 (N_4339,N_3165,N_3472);
nand U4340 (N_4340,N_3396,N_3933);
nand U4341 (N_4341,N_3901,N_3205);
nor U4342 (N_4342,N_3758,N_3041);
and U4343 (N_4343,N_3833,N_3271);
nor U4344 (N_4344,N_3296,N_3734);
and U4345 (N_4345,N_3601,N_3495);
nand U4346 (N_4346,N_3108,N_3842);
or U4347 (N_4347,N_3926,N_3949);
or U4348 (N_4348,N_3400,N_3799);
and U4349 (N_4349,N_3742,N_3292);
or U4350 (N_4350,N_3729,N_3487);
and U4351 (N_4351,N_3241,N_3683);
or U4352 (N_4352,N_3558,N_3424);
nand U4353 (N_4353,N_3145,N_3555);
nand U4354 (N_4354,N_3691,N_3114);
and U4355 (N_4355,N_3252,N_3995);
and U4356 (N_4356,N_3303,N_3460);
nor U4357 (N_4357,N_3503,N_3907);
nand U4358 (N_4358,N_3733,N_3293);
and U4359 (N_4359,N_3818,N_3475);
nor U4360 (N_4360,N_3019,N_3480);
nor U4361 (N_4361,N_3614,N_3931);
and U4362 (N_4362,N_3890,N_3174);
nand U4363 (N_4363,N_3045,N_3152);
nor U4364 (N_4364,N_3746,N_3673);
and U4365 (N_4365,N_3462,N_3457);
nor U4366 (N_4366,N_3602,N_3660);
or U4367 (N_4367,N_3529,N_3060);
nand U4368 (N_4368,N_3888,N_3617);
and U4369 (N_4369,N_3064,N_3720);
and U4370 (N_4370,N_3800,N_3054);
or U4371 (N_4371,N_3535,N_3492);
nand U4372 (N_4372,N_3620,N_3832);
or U4373 (N_4373,N_3442,N_3533);
or U4374 (N_4374,N_3217,N_3522);
nand U4375 (N_4375,N_3161,N_3922);
nor U4376 (N_4376,N_3168,N_3693);
nand U4377 (N_4377,N_3825,N_3372);
nor U4378 (N_4378,N_3859,N_3021);
and U4379 (N_4379,N_3351,N_3449);
nor U4380 (N_4380,N_3469,N_3084);
and U4381 (N_4381,N_3221,N_3775);
nand U4382 (N_4382,N_3804,N_3159);
and U4383 (N_4383,N_3593,N_3366);
and U4384 (N_4384,N_3684,N_3925);
and U4385 (N_4385,N_3029,N_3708);
nand U4386 (N_4386,N_3898,N_3219);
or U4387 (N_4387,N_3320,N_3606);
or U4388 (N_4388,N_3269,N_3308);
nor U4389 (N_4389,N_3419,N_3923);
and U4390 (N_4390,N_3610,N_3908);
nor U4391 (N_4391,N_3671,N_3588);
or U4392 (N_4392,N_3718,N_3385);
nand U4393 (N_4393,N_3175,N_3447);
or U4394 (N_4394,N_3325,N_3557);
nor U4395 (N_4395,N_3737,N_3324);
nor U4396 (N_4396,N_3576,N_3117);
nand U4397 (N_4397,N_3100,N_3226);
nor U4398 (N_4398,N_3334,N_3538);
or U4399 (N_4399,N_3158,N_3433);
or U4400 (N_4400,N_3319,N_3920);
nor U4401 (N_4401,N_3961,N_3743);
and U4402 (N_4402,N_3016,N_3479);
nand U4403 (N_4403,N_3656,N_3787);
nand U4404 (N_4404,N_3416,N_3915);
nor U4405 (N_4405,N_3482,N_3597);
and U4406 (N_4406,N_3886,N_3959);
and U4407 (N_4407,N_3653,N_3689);
and U4408 (N_4408,N_3323,N_3265);
or U4409 (N_4409,N_3631,N_3798);
nor U4410 (N_4410,N_3882,N_3803);
nor U4411 (N_4411,N_3542,N_3771);
nand U4412 (N_4412,N_3169,N_3318);
or U4413 (N_4413,N_3443,N_3405);
and U4414 (N_4414,N_3997,N_3377);
or U4415 (N_4415,N_3199,N_3454);
xnor U4416 (N_4416,N_3140,N_3373);
or U4417 (N_4417,N_3335,N_3565);
and U4418 (N_4418,N_3808,N_3154);
and U4419 (N_4419,N_3881,N_3344);
and U4420 (N_4420,N_3543,N_3790);
and U4421 (N_4421,N_3921,N_3772);
or U4422 (N_4422,N_3820,N_3537);
and U4423 (N_4423,N_3694,N_3137);
nand U4424 (N_4424,N_3530,N_3043);
nand U4425 (N_4425,N_3911,N_3608);
or U4426 (N_4426,N_3715,N_3083);
or U4427 (N_4427,N_3393,N_3127);
nand U4428 (N_4428,N_3719,N_3613);
nand U4429 (N_4429,N_3176,N_3975);
or U4430 (N_4430,N_3261,N_3973);
or U4431 (N_4431,N_3146,N_3844);
or U4432 (N_4432,N_3251,N_3278);
and U4433 (N_4433,N_3025,N_3383);
or U4434 (N_4434,N_3863,N_3467);
nand U4435 (N_4435,N_3240,N_3040);
nor U4436 (N_4436,N_3262,N_3430);
nand U4437 (N_4437,N_3329,N_3941);
nand U4438 (N_4438,N_3431,N_3196);
nand U4439 (N_4439,N_3493,N_3042);
nand U4440 (N_4440,N_3313,N_3722);
nand U4441 (N_4441,N_3756,N_3824);
nand U4442 (N_4442,N_3991,N_3582);
nand U4443 (N_4443,N_3109,N_3341);
nand U4444 (N_4444,N_3066,N_3491);
nand U4445 (N_4445,N_3270,N_3728);
or U4446 (N_4446,N_3218,N_3352);
or U4447 (N_4447,N_3536,N_3123);
and U4448 (N_4448,N_3316,N_3650);
nor U4449 (N_4449,N_3391,N_3056);
nand U4450 (N_4450,N_3357,N_3754);
nor U4451 (N_4451,N_3674,N_3611);
nor U4452 (N_4452,N_3212,N_3163);
xor U4453 (N_4453,N_3409,N_3246);
nand U4454 (N_4454,N_3513,N_3249);
and U4455 (N_4455,N_3345,N_3410);
or U4456 (N_4456,N_3836,N_3786);
or U4457 (N_4457,N_3211,N_3151);
nand U4458 (N_4458,N_3081,N_3417);
or U4459 (N_4459,N_3612,N_3916);
and U4460 (N_4460,N_3525,N_3521);
nor U4461 (N_4461,N_3183,N_3899);
or U4462 (N_4462,N_3919,N_3213);
or U4463 (N_4463,N_3571,N_3047);
nor U4464 (N_4464,N_3311,N_3766);
nor U4465 (N_4465,N_3214,N_3553);
nor U4466 (N_4466,N_3439,N_3420);
and U4467 (N_4467,N_3024,N_3962);
nor U4468 (N_4468,N_3014,N_3275);
nand U4469 (N_4469,N_3552,N_3929);
nand U4470 (N_4470,N_3062,N_3119);
nand U4471 (N_4471,N_3242,N_3490);
or U4472 (N_4472,N_3841,N_3144);
and U4473 (N_4473,N_3458,N_3843);
nand U4474 (N_4474,N_3823,N_3769);
nand U4475 (N_4475,N_3387,N_3879);
nand U4476 (N_4476,N_3891,N_3131);
and U4477 (N_4477,N_3935,N_3638);
or U4478 (N_4478,N_3646,N_3502);
or U4479 (N_4479,N_3583,N_3580);
nand U4480 (N_4480,N_3627,N_3381);
nand U4481 (N_4481,N_3086,N_3356);
or U4482 (N_4482,N_3677,N_3622);
and U4483 (N_4483,N_3518,N_3856);
nand U4484 (N_4484,N_3207,N_3678);
and U4485 (N_4485,N_3012,N_3672);
and U4486 (N_4486,N_3030,N_3403);
nand U4487 (N_4487,N_3655,N_3294);
or U4488 (N_4488,N_3266,N_3336);
or U4489 (N_4489,N_3817,N_3849);
nor U4490 (N_4490,N_3474,N_3295);
nor U4491 (N_4491,N_3272,N_3452);
nor U4492 (N_4492,N_3402,N_3363);
or U4493 (N_4493,N_3022,N_3598);
or U4494 (N_4494,N_3864,N_3889);
nand U4495 (N_4495,N_3143,N_3930);
nand U4496 (N_4496,N_3473,N_3407);
nand U4497 (N_4497,N_3591,N_3853);
and U4498 (N_4498,N_3496,N_3120);
or U4499 (N_4499,N_3076,N_3838);
nor U4500 (N_4500,N_3307,N_3241);
or U4501 (N_4501,N_3106,N_3738);
and U4502 (N_4502,N_3870,N_3978);
nand U4503 (N_4503,N_3672,N_3406);
nor U4504 (N_4504,N_3690,N_3784);
and U4505 (N_4505,N_3314,N_3997);
nand U4506 (N_4506,N_3813,N_3647);
or U4507 (N_4507,N_3806,N_3850);
nor U4508 (N_4508,N_3985,N_3871);
nor U4509 (N_4509,N_3517,N_3002);
or U4510 (N_4510,N_3537,N_3737);
nor U4511 (N_4511,N_3509,N_3880);
nand U4512 (N_4512,N_3665,N_3344);
or U4513 (N_4513,N_3233,N_3591);
or U4514 (N_4514,N_3839,N_3225);
or U4515 (N_4515,N_3099,N_3544);
or U4516 (N_4516,N_3095,N_3421);
nand U4517 (N_4517,N_3389,N_3756);
nor U4518 (N_4518,N_3216,N_3208);
nor U4519 (N_4519,N_3363,N_3646);
nand U4520 (N_4520,N_3597,N_3566);
nor U4521 (N_4521,N_3556,N_3283);
nand U4522 (N_4522,N_3015,N_3615);
and U4523 (N_4523,N_3053,N_3503);
and U4524 (N_4524,N_3548,N_3754);
nand U4525 (N_4525,N_3387,N_3332);
nor U4526 (N_4526,N_3949,N_3434);
and U4527 (N_4527,N_3365,N_3812);
nor U4528 (N_4528,N_3310,N_3723);
and U4529 (N_4529,N_3603,N_3163);
nand U4530 (N_4530,N_3064,N_3338);
and U4531 (N_4531,N_3335,N_3389);
or U4532 (N_4532,N_3742,N_3902);
nor U4533 (N_4533,N_3222,N_3170);
and U4534 (N_4534,N_3993,N_3032);
or U4535 (N_4535,N_3156,N_3482);
or U4536 (N_4536,N_3724,N_3885);
or U4537 (N_4537,N_3191,N_3888);
nand U4538 (N_4538,N_3922,N_3537);
nor U4539 (N_4539,N_3807,N_3464);
nor U4540 (N_4540,N_3662,N_3304);
and U4541 (N_4541,N_3989,N_3728);
or U4542 (N_4542,N_3913,N_3091);
xor U4543 (N_4543,N_3467,N_3720);
nand U4544 (N_4544,N_3133,N_3980);
or U4545 (N_4545,N_3528,N_3263);
and U4546 (N_4546,N_3941,N_3903);
nand U4547 (N_4547,N_3536,N_3583);
nor U4548 (N_4548,N_3609,N_3758);
or U4549 (N_4549,N_3062,N_3425);
nand U4550 (N_4550,N_3946,N_3154);
nor U4551 (N_4551,N_3146,N_3201);
nor U4552 (N_4552,N_3471,N_3910);
or U4553 (N_4553,N_3856,N_3689);
or U4554 (N_4554,N_3784,N_3065);
nand U4555 (N_4555,N_3218,N_3700);
or U4556 (N_4556,N_3708,N_3382);
nor U4557 (N_4557,N_3450,N_3699);
nand U4558 (N_4558,N_3380,N_3568);
or U4559 (N_4559,N_3032,N_3360);
or U4560 (N_4560,N_3322,N_3130);
and U4561 (N_4561,N_3801,N_3738);
nor U4562 (N_4562,N_3189,N_3785);
nand U4563 (N_4563,N_3011,N_3755);
or U4564 (N_4564,N_3303,N_3139);
and U4565 (N_4565,N_3120,N_3762);
and U4566 (N_4566,N_3770,N_3252);
or U4567 (N_4567,N_3414,N_3550);
nor U4568 (N_4568,N_3488,N_3662);
or U4569 (N_4569,N_3808,N_3315);
xnor U4570 (N_4570,N_3878,N_3509);
and U4571 (N_4571,N_3028,N_3251);
and U4572 (N_4572,N_3613,N_3162);
nand U4573 (N_4573,N_3196,N_3910);
nand U4574 (N_4574,N_3689,N_3275);
nor U4575 (N_4575,N_3769,N_3957);
nor U4576 (N_4576,N_3744,N_3471);
nor U4577 (N_4577,N_3699,N_3245);
or U4578 (N_4578,N_3236,N_3299);
or U4579 (N_4579,N_3530,N_3739);
nor U4580 (N_4580,N_3177,N_3440);
or U4581 (N_4581,N_3803,N_3115);
nand U4582 (N_4582,N_3709,N_3084);
nand U4583 (N_4583,N_3918,N_3026);
nor U4584 (N_4584,N_3579,N_3197);
and U4585 (N_4585,N_3445,N_3008);
and U4586 (N_4586,N_3288,N_3704);
nand U4587 (N_4587,N_3895,N_3869);
and U4588 (N_4588,N_3007,N_3173);
nand U4589 (N_4589,N_3740,N_3321);
nand U4590 (N_4590,N_3203,N_3401);
nand U4591 (N_4591,N_3033,N_3771);
or U4592 (N_4592,N_3385,N_3693);
and U4593 (N_4593,N_3348,N_3680);
nand U4594 (N_4594,N_3328,N_3593);
or U4595 (N_4595,N_3444,N_3390);
nor U4596 (N_4596,N_3613,N_3929);
nand U4597 (N_4597,N_3821,N_3612);
nand U4598 (N_4598,N_3071,N_3015);
or U4599 (N_4599,N_3342,N_3514);
or U4600 (N_4600,N_3421,N_3976);
nand U4601 (N_4601,N_3173,N_3448);
nor U4602 (N_4602,N_3459,N_3339);
and U4603 (N_4603,N_3757,N_3041);
or U4604 (N_4604,N_3538,N_3868);
nand U4605 (N_4605,N_3496,N_3287);
or U4606 (N_4606,N_3442,N_3238);
nor U4607 (N_4607,N_3809,N_3650);
and U4608 (N_4608,N_3669,N_3914);
nor U4609 (N_4609,N_3091,N_3105);
nor U4610 (N_4610,N_3493,N_3697);
nor U4611 (N_4611,N_3843,N_3609);
nand U4612 (N_4612,N_3864,N_3554);
nor U4613 (N_4613,N_3825,N_3918);
or U4614 (N_4614,N_3466,N_3323);
or U4615 (N_4615,N_3695,N_3194);
nor U4616 (N_4616,N_3666,N_3040);
nor U4617 (N_4617,N_3776,N_3165);
and U4618 (N_4618,N_3941,N_3449);
nor U4619 (N_4619,N_3772,N_3433);
or U4620 (N_4620,N_3393,N_3605);
and U4621 (N_4621,N_3765,N_3857);
or U4622 (N_4622,N_3223,N_3366);
nand U4623 (N_4623,N_3844,N_3297);
and U4624 (N_4624,N_3968,N_3731);
nor U4625 (N_4625,N_3040,N_3962);
nand U4626 (N_4626,N_3695,N_3856);
or U4627 (N_4627,N_3812,N_3142);
or U4628 (N_4628,N_3549,N_3469);
nand U4629 (N_4629,N_3547,N_3769);
and U4630 (N_4630,N_3842,N_3033);
nand U4631 (N_4631,N_3746,N_3989);
nor U4632 (N_4632,N_3493,N_3399);
nand U4633 (N_4633,N_3208,N_3337);
and U4634 (N_4634,N_3814,N_3162);
or U4635 (N_4635,N_3010,N_3846);
xor U4636 (N_4636,N_3399,N_3117);
nand U4637 (N_4637,N_3734,N_3162);
nand U4638 (N_4638,N_3027,N_3017);
or U4639 (N_4639,N_3181,N_3135);
nor U4640 (N_4640,N_3992,N_3540);
and U4641 (N_4641,N_3603,N_3440);
and U4642 (N_4642,N_3776,N_3298);
nor U4643 (N_4643,N_3094,N_3381);
nand U4644 (N_4644,N_3134,N_3094);
nor U4645 (N_4645,N_3714,N_3857);
xor U4646 (N_4646,N_3467,N_3818);
nand U4647 (N_4647,N_3543,N_3114);
nand U4648 (N_4648,N_3716,N_3079);
or U4649 (N_4649,N_3613,N_3823);
or U4650 (N_4650,N_3942,N_3027);
or U4651 (N_4651,N_3364,N_3896);
nand U4652 (N_4652,N_3108,N_3839);
nand U4653 (N_4653,N_3594,N_3605);
or U4654 (N_4654,N_3298,N_3904);
nand U4655 (N_4655,N_3368,N_3735);
nor U4656 (N_4656,N_3360,N_3962);
nor U4657 (N_4657,N_3081,N_3123);
nand U4658 (N_4658,N_3691,N_3715);
nand U4659 (N_4659,N_3074,N_3919);
and U4660 (N_4660,N_3276,N_3936);
nor U4661 (N_4661,N_3525,N_3762);
nand U4662 (N_4662,N_3568,N_3726);
or U4663 (N_4663,N_3403,N_3271);
and U4664 (N_4664,N_3441,N_3136);
nor U4665 (N_4665,N_3102,N_3998);
and U4666 (N_4666,N_3222,N_3781);
nand U4667 (N_4667,N_3020,N_3448);
and U4668 (N_4668,N_3442,N_3649);
or U4669 (N_4669,N_3878,N_3171);
or U4670 (N_4670,N_3954,N_3221);
or U4671 (N_4671,N_3305,N_3017);
nand U4672 (N_4672,N_3224,N_3951);
nand U4673 (N_4673,N_3336,N_3585);
or U4674 (N_4674,N_3214,N_3701);
and U4675 (N_4675,N_3927,N_3423);
nand U4676 (N_4676,N_3481,N_3940);
nand U4677 (N_4677,N_3002,N_3458);
and U4678 (N_4678,N_3530,N_3401);
or U4679 (N_4679,N_3686,N_3928);
nor U4680 (N_4680,N_3808,N_3517);
nand U4681 (N_4681,N_3639,N_3055);
nor U4682 (N_4682,N_3145,N_3504);
or U4683 (N_4683,N_3027,N_3458);
or U4684 (N_4684,N_3347,N_3419);
nand U4685 (N_4685,N_3355,N_3545);
nand U4686 (N_4686,N_3530,N_3497);
nor U4687 (N_4687,N_3426,N_3036);
or U4688 (N_4688,N_3837,N_3665);
nor U4689 (N_4689,N_3749,N_3010);
nand U4690 (N_4690,N_3188,N_3573);
and U4691 (N_4691,N_3036,N_3851);
or U4692 (N_4692,N_3427,N_3010);
nor U4693 (N_4693,N_3766,N_3959);
nand U4694 (N_4694,N_3447,N_3279);
or U4695 (N_4695,N_3667,N_3281);
nand U4696 (N_4696,N_3217,N_3288);
and U4697 (N_4697,N_3009,N_3281);
and U4698 (N_4698,N_3438,N_3940);
nor U4699 (N_4699,N_3964,N_3488);
nor U4700 (N_4700,N_3463,N_3764);
nand U4701 (N_4701,N_3693,N_3739);
or U4702 (N_4702,N_3743,N_3663);
and U4703 (N_4703,N_3681,N_3610);
nor U4704 (N_4704,N_3193,N_3200);
nand U4705 (N_4705,N_3932,N_3963);
nor U4706 (N_4706,N_3086,N_3990);
and U4707 (N_4707,N_3960,N_3199);
nor U4708 (N_4708,N_3697,N_3938);
or U4709 (N_4709,N_3953,N_3508);
nand U4710 (N_4710,N_3955,N_3178);
or U4711 (N_4711,N_3358,N_3713);
nand U4712 (N_4712,N_3794,N_3444);
nand U4713 (N_4713,N_3623,N_3443);
nand U4714 (N_4714,N_3400,N_3032);
and U4715 (N_4715,N_3025,N_3054);
nor U4716 (N_4716,N_3651,N_3999);
or U4717 (N_4717,N_3586,N_3522);
nor U4718 (N_4718,N_3566,N_3973);
or U4719 (N_4719,N_3820,N_3111);
and U4720 (N_4720,N_3534,N_3480);
or U4721 (N_4721,N_3755,N_3711);
and U4722 (N_4722,N_3747,N_3487);
and U4723 (N_4723,N_3534,N_3077);
or U4724 (N_4724,N_3085,N_3364);
nor U4725 (N_4725,N_3718,N_3086);
nor U4726 (N_4726,N_3152,N_3948);
nand U4727 (N_4727,N_3909,N_3969);
nand U4728 (N_4728,N_3932,N_3070);
or U4729 (N_4729,N_3283,N_3069);
nor U4730 (N_4730,N_3538,N_3415);
nand U4731 (N_4731,N_3751,N_3059);
nand U4732 (N_4732,N_3178,N_3614);
or U4733 (N_4733,N_3793,N_3610);
or U4734 (N_4734,N_3495,N_3941);
and U4735 (N_4735,N_3293,N_3185);
or U4736 (N_4736,N_3986,N_3334);
nand U4737 (N_4737,N_3506,N_3372);
or U4738 (N_4738,N_3391,N_3456);
or U4739 (N_4739,N_3587,N_3313);
nand U4740 (N_4740,N_3357,N_3019);
or U4741 (N_4741,N_3281,N_3299);
or U4742 (N_4742,N_3134,N_3298);
and U4743 (N_4743,N_3868,N_3351);
nand U4744 (N_4744,N_3817,N_3341);
and U4745 (N_4745,N_3706,N_3302);
and U4746 (N_4746,N_3248,N_3439);
nor U4747 (N_4747,N_3559,N_3925);
nand U4748 (N_4748,N_3854,N_3343);
or U4749 (N_4749,N_3446,N_3195);
nand U4750 (N_4750,N_3495,N_3170);
or U4751 (N_4751,N_3057,N_3864);
and U4752 (N_4752,N_3281,N_3961);
nor U4753 (N_4753,N_3205,N_3273);
or U4754 (N_4754,N_3902,N_3896);
and U4755 (N_4755,N_3741,N_3008);
nand U4756 (N_4756,N_3051,N_3097);
nor U4757 (N_4757,N_3380,N_3482);
nor U4758 (N_4758,N_3777,N_3586);
nor U4759 (N_4759,N_3059,N_3547);
nor U4760 (N_4760,N_3015,N_3810);
nor U4761 (N_4761,N_3432,N_3607);
or U4762 (N_4762,N_3326,N_3788);
nor U4763 (N_4763,N_3495,N_3463);
nand U4764 (N_4764,N_3135,N_3666);
and U4765 (N_4765,N_3135,N_3505);
or U4766 (N_4766,N_3604,N_3169);
nand U4767 (N_4767,N_3781,N_3576);
nor U4768 (N_4768,N_3749,N_3188);
nor U4769 (N_4769,N_3178,N_3660);
and U4770 (N_4770,N_3649,N_3451);
and U4771 (N_4771,N_3487,N_3087);
nor U4772 (N_4772,N_3271,N_3391);
nor U4773 (N_4773,N_3228,N_3762);
and U4774 (N_4774,N_3288,N_3518);
nand U4775 (N_4775,N_3964,N_3146);
nor U4776 (N_4776,N_3936,N_3983);
nand U4777 (N_4777,N_3174,N_3032);
nor U4778 (N_4778,N_3120,N_3505);
or U4779 (N_4779,N_3985,N_3211);
or U4780 (N_4780,N_3174,N_3562);
or U4781 (N_4781,N_3651,N_3361);
or U4782 (N_4782,N_3792,N_3080);
nand U4783 (N_4783,N_3889,N_3686);
nand U4784 (N_4784,N_3230,N_3290);
nor U4785 (N_4785,N_3661,N_3112);
nand U4786 (N_4786,N_3445,N_3263);
nand U4787 (N_4787,N_3416,N_3003);
and U4788 (N_4788,N_3993,N_3225);
nor U4789 (N_4789,N_3065,N_3638);
nand U4790 (N_4790,N_3122,N_3508);
and U4791 (N_4791,N_3493,N_3212);
and U4792 (N_4792,N_3768,N_3449);
and U4793 (N_4793,N_3536,N_3837);
and U4794 (N_4794,N_3748,N_3660);
or U4795 (N_4795,N_3416,N_3279);
and U4796 (N_4796,N_3699,N_3384);
and U4797 (N_4797,N_3913,N_3604);
and U4798 (N_4798,N_3921,N_3504);
and U4799 (N_4799,N_3458,N_3024);
nor U4800 (N_4800,N_3895,N_3326);
or U4801 (N_4801,N_3549,N_3327);
nor U4802 (N_4802,N_3099,N_3275);
and U4803 (N_4803,N_3860,N_3698);
nand U4804 (N_4804,N_3478,N_3054);
nand U4805 (N_4805,N_3415,N_3287);
nor U4806 (N_4806,N_3611,N_3907);
or U4807 (N_4807,N_3283,N_3125);
or U4808 (N_4808,N_3320,N_3281);
and U4809 (N_4809,N_3772,N_3440);
or U4810 (N_4810,N_3570,N_3000);
or U4811 (N_4811,N_3289,N_3716);
or U4812 (N_4812,N_3034,N_3583);
and U4813 (N_4813,N_3710,N_3420);
or U4814 (N_4814,N_3432,N_3685);
nand U4815 (N_4815,N_3754,N_3400);
or U4816 (N_4816,N_3289,N_3228);
and U4817 (N_4817,N_3362,N_3961);
or U4818 (N_4818,N_3203,N_3867);
nor U4819 (N_4819,N_3806,N_3667);
or U4820 (N_4820,N_3842,N_3120);
nor U4821 (N_4821,N_3001,N_3862);
and U4822 (N_4822,N_3215,N_3094);
nor U4823 (N_4823,N_3245,N_3841);
nor U4824 (N_4824,N_3333,N_3985);
nor U4825 (N_4825,N_3329,N_3992);
nor U4826 (N_4826,N_3647,N_3461);
and U4827 (N_4827,N_3201,N_3607);
and U4828 (N_4828,N_3503,N_3428);
nor U4829 (N_4829,N_3828,N_3243);
nand U4830 (N_4830,N_3092,N_3368);
nand U4831 (N_4831,N_3967,N_3524);
or U4832 (N_4832,N_3494,N_3268);
nor U4833 (N_4833,N_3734,N_3621);
nor U4834 (N_4834,N_3930,N_3067);
nand U4835 (N_4835,N_3900,N_3747);
nand U4836 (N_4836,N_3314,N_3841);
or U4837 (N_4837,N_3895,N_3056);
or U4838 (N_4838,N_3609,N_3149);
nand U4839 (N_4839,N_3026,N_3655);
and U4840 (N_4840,N_3124,N_3362);
nor U4841 (N_4841,N_3706,N_3027);
nor U4842 (N_4842,N_3693,N_3347);
or U4843 (N_4843,N_3421,N_3846);
and U4844 (N_4844,N_3771,N_3995);
or U4845 (N_4845,N_3669,N_3145);
xnor U4846 (N_4846,N_3955,N_3796);
or U4847 (N_4847,N_3743,N_3865);
or U4848 (N_4848,N_3056,N_3263);
or U4849 (N_4849,N_3881,N_3759);
nor U4850 (N_4850,N_3447,N_3348);
nor U4851 (N_4851,N_3540,N_3972);
and U4852 (N_4852,N_3307,N_3684);
nor U4853 (N_4853,N_3565,N_3222);
nand U4854 (N_4854,N_3260,N_3466);
nor U4855 (N_4855,N_3162,N_3184);
and U4856 (N_4856,N_3669,N_3469);
nand U4857 (N_4857,N_3323,N_3378);
nor U4858 (N_4858,N_3187,N_3233);
or U4859 (N_4859,N_3192,N_3599);
or U4860 (N_4860,N_3605,N_3158);
and U4861 (N_4861,N_3153,N_3851);
or U4862 (N_4862,N_3932,N_3429);
or U4863 (N_4863,N_3774,N_3190);
nand U4864 (N_4864,N_3985,N_3933);
or U4865 (N_4865,N_3798,N_3708);
and U4866 (N_4866,N_3839,N_3025);
nor U4867 (N_4867,N_3895,N_3749);
and U4868 (N_4868,N_3668,N_3666);
and U4869 (N_4869,N_3217,N_3935);
nand U4870 (N_4870,N_3709,N_3515);
and U4871 (N_4871,N_3033,N_3716);
and U4872 (N_4872,N_3985,N_3957);
or U4873 (N_4873,N_3898,N_3097);
xor U4874 (N_4874,N_3348,N_3897);
or U4875 (N_4875,N_3247,N_3971);
nor U4876 (N_4876,N_3456,N_3383);
nand U4877 (N_4877,N_3812,N_3250);
and U4878 (N_4878,N_3116,N_3275);
nor U4879 (N_4879,N_3742,N_3507);
nor U4880 (N_4880,N_3752,N_3557);
and U4881 (N_4881,N_3339,N_3279);
nor U4882 (N_4882,N_3717,N_3720);
or U4883 (N_4883,N_3430,N_3245);
or U4884 (N_4884,N_3183,N_3451);
and U4885 (N_4885,N_3334,N_3519);
nand U4886 (N_4886,N_3008,N_3761);
nor U4887 (N_4887,N_3871,N_3738);
nor U4888 (N_4888,N_3535,N_3334);
or U4889 (N_4889,N_3301,N_3263);
nor U4890 (N_4890,N_3186,N_3878);
or U4891 (N_4891,N_3104,N_3327);
nand U4892 (N_4892,N_3002,N_3728);
nand U4893 (N_4893,N_3220,N_3811);
nor U4894 (N_4894,N_3139,N_3207);
or U4895 (N_4895,N_3955,N_3308);
xor U4896 (N_4896,N_3371,N_3701);
and U4897 (N_4897,N_3997,N_3725);
nor U4898 (N_4898,N_3023,N_3085);
nand U4899 (N_4899,N_3669,N_3762);
nor U4900 (N_4900,N_3764,N_3868);
nor U4901 (N_4901,N_3859,N_3191);
or U4902 (N_4902,N_3526,N_3560);
nand U4903 (N_4903,N_3881,N_3827);
or U4904 (N_4904,N_3066,N_3882);
or U4905 (N_4905,N_3268,N_3991);
or U4906 (N_4906,N_3653,N_3771);
and U4907 (N_4907,N_3235,N_3280);
and U4908 (N_4908,N_3414,N_3625);
or U4909 (N_4909,N_3349,N_3835);
nor U4910 (N_4910,N_3811,N_3095);
nand U4911 (N_4911,N_3279,N_3737);
nand U4912 (N_4912,N_3950,N_3486);
or U4913 (N_4913,N_3634,N_3423);
or U4914 (N_4914,N_3008,N_3663);
nor U4915 (N_4915,N_3008,N_3652);
and U4916 (N_4916,N_3709,N_3800);
and U4917 (N_4917,N_3264,N_3015);
and U4918 (N_4918,N_3503,N_3522);
nand U4919 (N_4919,N_3630,N_3260);
and U4920 (N_4920,N_3228,N_3654);
and U4921 (N_4921,N_3184,N_3384);
and U4922 (N_4922,N_3121,N_3122);
or U4923 (N_4923,N_3586,N_3222);
and U4924 (N_4924,N_3525,N_3459);
nor U4925 (N_4925,N_3092,N_3237);
or U4926 (N_4926,N_3657,N_3926);
xor U4927 (N_4927,N_3766,N_3237);
or U4928 (N_4928,N_3037,N_3323);
nand U4929 (N_4929,N_3658,N_3405);
and U4930 (N_4930,N_3800,N_3285);
nor U4931 (N_4931,N_3686,N_3012);
nand U4932 (N_4932,N_3111,N_3631);
nand U4933 (N_4933,N_3971,N_3205);
nand U4934 (N_4934,N_3390,N_3313);
nor U4935 (N_4935,N_3782,N_3987);
or U4936 (N_4936,N_3629,N_3431);
and U4937 (N_4937,N_3963,N_3434);
or U4938 (N_4938,N_3433,N_3404);
and U4939 (N_4939,N_3834,N_3536);
nor U4940 (N_4940,N_3649,N_3337);
nand U4941 (N_4941,N_3411,N_3227);
nand U4942 (N_4942,N_3431,N_3321);
or U4943 (N_4943,N_3488,N_3223);
and U4944 (N_4944,N_3868,N_3362);
or U4945 (N_4945,N_3921,N_3155);
or U4946 (N_4946,N_3751,N_3229);
and U4947 (N_4947,N_3579,N_3540);
nor U4948 (N_4948,N_3694,N_3178);
nor U4949 (N_4949,N_3788,N_3720);
or U4950 (N_4950,N_3162,N_3562);
nand U4951 (N_4951,N_3292,N_3392);
or U4952 (N_4952,N_3421,N_3586);
and U4953 (N_4953,N_3513,N_3050);
and U4954 (N_4954,N_3535,N_3796);
nor U4955 (N_4955,N_3531,N_3721);
nand U4956 (N_4956,N_3825,N_3963);
or U4957 (N_4957,N_3345,N_3725);
or U4958 (N_4958,N_3229,N_3893);
or U4959 (N_4959,N_3335,N_3095);
or U4960 (N_4960,N_3782,N_3555);
or U4961 (N_4961,N_3629,N_3776);
nand U4962 (N_4962,N_3014,N_3642);
or U4963 (N_4963,N_3002,N_3251);
nor U4964 (N_4964,N_3191,N_3188);
nor U4965 (N_4965,N_3980,N_3141);
nand U4966 (N_4966,N_3443,N_3258);
and U4967 (N_4967,N_3959,N_3067);
and U4968 (N_4968,N_3329,N_3859);
nor U4969 (N_4969,N_3904,N_3583);
or U4970 (N_4970,N_3294,N_3616);
nor U4971 (N_4971,N_3227,N_3241);
nand U4972 (N_4972,N_3660,N_3225);
nand U4973 (N_4973,N_3923,N_3247);
and U4974 (N_4974,N_3965,N_3361);
and U4975 (N_4975,N_3066,N_3050);
nor U4976 (N_4976,N_3512,N_3237);
nor U4977 (N_4977,N_3402,N_3622);
and U4978 (N_4978,N_3393,N_3723);
and U4979 (N_4979,N_3958,N_3365);
nor U4980 (N_4980,N_3432,N_3012);
or U4981 (N_4981,N_3453,N_3935);
nand U4982 (N_4982,N_3520,N_3163);
or U4983 (N_4983,N_3124,N_3640);
nor U4984 (N_4984,N_3108,N_3829);
and U4985 (N_4985,N_3473,N_3915);
and U4986 (N_4986,N_3531,N_3790);
nand U4987 (N_4987,N_3821,N_3749);
xor U4988 (N_4988,N_3154,N_3518);
nor U4989 (N_4989,N_3315,N_3256);
or U4990 (N_4990,N_3895,N_3703);
nand U4991 (N_4991,N_3978,N_3685);
or U4992 (N_4992,N_3265,N_3293);
or U4993 (N_4993,N_3076,N_3562);
nand U4994 (N_4994,N_3609,N_3098);
and U4995 (N_4995,N_3048,N_3686);
nor U4996 (N_4996,N_3166,N_3286);
nor U4997 (N_4997,N_3729,N_3109);
nand U4998 (N_4998,N_3930,N_3632);
nor U4999 (N_4999,N_3383,N_3622);
or U5000 (N_5000,N_4399,N_4662);
nand U5001 (N_5001,N_4082,N_4079);
or U5002 (N_5002,N_4950,N_4222);
or U5003 (N_5003,N_4672,N_4324);
nor U5004 (N_5004,N_4437,N_4373);
nor U5005 (N_5005,N_4684,N_4893);
or U5006 (N_5006,N_4901,N_4622);
and U5007 (N_5007,N_4561,N_4003);
xor U5008 (N_5008,N_4503,N_4468);
nor U5009 (N_5009,N_4416,N_4525);
or U5010 (N_5010,N_4858,N_4822);
and U5011 (N_5011,N_4170,N_4095);
nor U5012 (N_5012,N_4466,N_4993);
nor U5013 (N_5013,N_4743,N_4796);
nor U5014 (N_5014,N_4763,N_4550);
or U5015 (N_5015,N_4517,N_4974);
nor U5016 (N_5016,N_4707,N_4855);
nor U5017 (N_5017,N_4012,N_4188);
or U5018 (N_5018,N_4345,N_4702);
nand U5019 (N_5019,N_4093,N_4395);
nor U5020 (N_5020,N_4911,N_4547);
and U5021 (N_5021,N_4654,N_4757);
nand U5022 (N_5022,N_4585,N_4570);
nand U5023 (N_5023,N_4758,N_4803);
nand U5024 (N_5024,N_4101,N_4545);
and U5025 (N_5025,N_4464,N_4669);
nand U5026 (N_5026,N_4594,N_4586);
nor U5027 (N_5027,N_4853,N_4411);
nor U5028 (N_5028,N_4535,N_4029);
nand U5029 (N_5029,N_4209,N_4904);
nand U5030 (N_5030,N_4938,N_4293);
and U5031 (N_5031,N_4750,N_4691);
nand U5032 (N_5032,N_4176,N_4870);
nand U5033 (N_5033,N_4818,N_4939);
nor U5034 (N_5034,N_4027,N_4231);
and U5035 (N_5035,N_4916,N_4582);
nor U5036 (N_5036,N_4753,N_4787);
or U5037 (N_5037,N_4652,N_4429);
or U5038 (N_5038,N_4329,N_4339);
or U5039 (N_5039,N_4191,N_4857);
nor U5040 (N_5040,N_4600,N_4267);
nand U5041 (N_5041,N_4184,N_4829);
xor U5042 (N_5042,N_4051,N_4747);
and U5043 (N_5043,N_4276,N_4733);
or U5044 (N_5044,N_4877,N_4167);
or U5045 (N_5045,N_4462,N_4777);
nand U5046 (N_5046,N_4283,N_4129);
nor U5047 (N_5047,N_4371,N_4103);
and U5048 (N_5048,N_4386,N_4649);
and U5049 (N_5049,N_4784,N_4775);
nor U5050 (N_5050,N_4348,N_4526);
nand U5051 (N_5051,N_4794,N_4761);
or U5052 (N_5052,N_4328,N_4618);
or U5053 (N_5053,N_4040,N_4154);
and U5054 (N_5054,N_4709,N_4984);
nor U5055 (N_5055,N_4491,N_4490);
nor U5056 (N_5056,N_4039,N_4971);
nand U5057 (N_5057,N_4512,N_4653);
nor U5058 (N_5058,N_4088,N_4797);
or U5059 (N_5059,N_4655,N_4241);
and U5060 (N_5060,N_4885,N_4495);
nand U5061 (N_5061,N_4420,N_4453);
nor U5062 (N_5062,N_4951,N_4224);
or U5063 (N_5063,N_4929,N_4456);
nor U5064 (N_5064,N_4712,N_4113);
or U5065 (N_5065,N_4940,N_4620);
nor U5066 (N_5066,N_4480,N_4615);
and U5067 (N_5067,N_4382,N_4350);
or U5068 (N_5068,N_4045,N_4683);
and U5069 (N_5069,N_4827,N_4041);
or U5070 (N_5070,N_4115,N_4835);
nor U5071 (N_5071,N_4770,N_4659);
or U5072 (N_5072,N_4201,N_4583);
nor U5073 (N_5073,N_4403,N_4694);
or U5074 (N_5074,N_4979,N_4821);
or U5075 (N_5075,N_4352,N_4776);
nor U5076 (N_5076,N_4643,N_4688);
nand U5077 (N_5077,N_4214,N_4319);
and U5078 (N_5078,N_4054,N_4160);
nor U5079 (N_5079,N_4919,N_4987);
nand U5080 (N_5080,N_4365,N_4566);
or U5081 (N_5081,N_4179,N_4445);
nand U5082 (N_5082,N_4174,N_4349);
nand U5083 (N_5083,N_4021,N_4237);
nand U5084 (N_5084,N_4754,N_4676);
nand U5085 (N_5085,N_4133,N_4675);
and U5086 (N_5086,N_4166,N_4623);
and U5087 (N_5087,N_4508,N_4959);
nor U5088 (N_5088,N_4047,N_4717);
nand U5089 (N_5089,N_4251,N_4142);
nor U5090 (N_5090,N_4791,N_4514);
nor U5091 (N_5091,N_4851,N_4700);
nand U5092 (N_5092,N_4457,N_4104);
or U5093 (N_5093,N_4628,N_4376);
nor U5094 (N_5094,N_4390,N_4367);
or U5095 (N_5095,N_4317,N_4217);
nor U5096 (N_5096,N_4132,N_4347);
nand U5097 (N_5097,N_4250,N_4891);
nor U5098 (N_5098,N_4286,N_4931);
and U5099 (N_5099,N_4605,N_4837);
nor U5100 (N_5100,N_4557,N_4579);
xor U5101 (N_5101,N_4478,N_4446);
or U5102 (N_5102,N_4368,N_4769);
nor U5103 (N_5103,N_4599,N_4022);
nor U5104 (N_5104,N_4455,N_4522);
nand U5105 (N_5105,N_4543,N_4363);
xnor U5106 (N_5106,N_4590,N_4255);
nor U5107 (N_5107,N_4482,N_4076);
nor U5108 (N_5108,N_4779,N_4894);
or U5109 (N_5109,N_4513,N_4812);
and U5110 (N_5110,N_4243,N_4888);
nor U5111 (N_5111,N_4872,N_4679);
or U5112 (N_5112,N_4606,N_4426);
and U5113 (N_5113,N_4704,N_4258);
or U5114 (N_5114,N_4074,N_4299);
nor U5115 (N_5115,N_4854,N_4555);
and U5116 (N_5116,N_4072,N_4660);
or U5117 (N_5117,N_4730,N_4573);
or U5118 (N_5118,N_4856,N_4266);
nand U5119 (N_5119,N_4591,N_4026);
nand U5120 (N_5120,N_4344,N_4504);
or U5121 (N_5121,N_4746,N_4354);
xnor U5122 (N_5122,N_4177,N_4533);
and U5123 (N_5123,N_4942,N_4033);
nor U5124 (N_5124,N_4137,N_4621);
and U5125 (N_5125,N_4603,N_4185);
nand U5126 (N_5126,N_4398,N_4239);
nor U5127 (N_5127,N_4346,N_4548);
nand U5128 (N_5128,N_4500,N_4969);
or U5129 (N_5129,N_4634,N_4007);
and U5130 (N_5130,N_4648,N_4719);
nor U5131 (N_5131,N_4430,N_4278);
nor U5132 (N_5132,N_4073,N_4646);
nand U5133 (N_5133,N_4682,N_4492);
or U5134 (N_5134,N_4014,N_4650);
nand U5135 (N_5135,N_4145,N_4277);
or U5136 (N_5136,N_4832,N_4874);
nor U5137 (N_5137,N_4943,N_4289);
xnor U5138 (N_5138,N_4604,N_4476);
nand U5139 (N_5139,N_4147,N_4415);
or U5140 (N_5140,N_4988,N_4954);
nor U5141 (N_5141,N_4926,N_4296);
or U5142 (N_5142,N_4238,N_4001);
and U5143 (N_5143,N_4795,N_4218);
and U5144 (N_5144,N_4062,N_4633);
and U5145 (N_5145,N_4509,N_4448);
or U5146 (N_5146,N_4272,N_4895);
nand U5147 (N_5147,N_4537,N_4510);
and U5148 (N_5148,N_4486,N_4117);
and U5149 (N_5149,N_4859,N_4203);
or U5150 (N_5150,N_4678,N_4925);
and U5151 (N_5151,N_4256,N_4994);
and U5152 (N_5152,N_4595,N_4778);
nor U5153 (N_5153,N_4301,N_4866);
nor U5154 (N_5154,N_4805,N_4574);
and U5155 (N_5155,N_4444,N_4069);
nor U5156 (N_5156,N_4802,N_4275);
nand U5157 (N_5157,N_4941,N_4240);
or U5158 (N_5158,N_4078,N_4090);
nor U5159 (N_5159,N_4693,N_4171);
and U5160 (N_5160,N_4413,N_4249);
nor U5161 (N_5161,N_4970,N_4519);
xor U5162 (N_5162,N_4362,N_4773);
xor U5163 (N_5163,N_4656,N_4718);
nor U5164 (N_5164,N_4781,N_4559);
nor U5165 (N_5165,N_4013,N_4521);
xnor U5166 (N_5166,N_4609,N_4479);
nor U5167 (N_5167,N_4640,N_4128);
and U5168 (N_5168,N_4303,N_4175);
nand U5169 (N_5169,N_4488,N_4635);
and U5170 (N_5170,N_4774,N_4493);
nand U5171 (N_5171,N_4551,N_4976);
or U5172 (N_5172,N_4116,N_4424);
and U5173 (N_5173,N_4112,N_4842);
nand U5174 (N_5174,N_4198,N_4536);
nor U5175 (N_5175,N_4019,N_4157);
and U5176 (N_5176,N_4358,N_4125);
nor U5177 (N_5177,N_4729,N_4703);
nand U5178 (N_5178,N_4048,N_4638);
nor U5179 (N_5179,N_4542,N_4527);
or U5180 (N_5180,N_4418,N_4783);
nand U5181 (N_5181,N_4765,N_4864);
nand U5182 (N_5182,N_4505,N_4828);
or U5183 (N_5183,N_4955,N_4965);
or U5184 (N_5184,N_4696,N_4883);
and U5185 (N_5185,N_4035,N_4316);
nand U5186 (N_5186,N_4685,N_4274);
nor U5187 (N_5187,N_4152,N_4641);
and U5188 (N_5188,N_4742,N_4793);
or U5189 (N_5189,N_4708,N_4215);
or U5190 (N_5190,N_4098,N_4569);
or U5191 (N_5191,N_4879,N_4120);
nand U5192 (N_5192,N_4515,N_4936);
nand U5193 (N_5193,N_4830,N_4681);
and U5194 (N_5194,N_4099,N_4106);
nor U5195 (N_5195,N_4980,N_4865);
or U5196 (N_5196,N_4930,N_4952);
and U5197 (N_5197,N_4204,N_4452);
nand U5198 (N_5198,N_4111,N_4211);
nand U5199 (N_5199,N_4917,N_4875);
or U5200 (N_5200,N_4244,N_4330);
nor U5201 (N_5201,N_4210,N_4253);
and U5202 (N_5202,N_4999,N_4982);
nand U5203 (N_5203,N_4847,N_4169);
or U5204 (N_5204,N_4905,N_4944);
and U5205 (N_5205,N_4320,N_4182);
nor U5206 (N_5206,N_4886,N_4017);
nand U5207 (N_5207,N_4973,N_4037);
or U5208 (N_5208,N_4817,N_4809);
and U5209 (N_5209,N_4902,N_4540);
or U5210 (N_5210,N_4036,N_4531);
nor U5211 (N_5211,N_4028,N_4247);
or U5212 (N_5212,N_4738,N_4394);
nor U5213 (N_5213,N_4226,N_4121);
nand U5214 (N_5214,N_4392,N_4325);
or U5215 (N_5215,N_4966,N_4617);
nand U5216 (N_5216,N_4884,N_4181);
and U5217 (N_5217,N_4260,N_4567);
xnor U5218 (N_5218,N_4998,N_4506);
or U5219 (N_5219,N_4862,N_4731);
nor U5220 (N_5220,N_4610,N_4340);
nand U5221 (N_5221,N_4789,N_4421);
or U5222 (N_5222,N_4706,N_4196);
and U5223 (N_5223,N_4501,N_4192);
and U5224 (N_5224,N_4219,N_4524);
nor U5225 (N_5225,N_4447,N_4183);
xnor U5226 (N_5226,N_4186,N_4587);
or U5227 (N_5227,N_4564,N_4080);
nand U5228 (N_5228,N_4962,N_4337);
and U5229 (N_5229,N_4661,N_4530);
nor U5230 (N_5230,N_4897,N_4923);
nor U5231 (N_5231,N_4589,N_4248);
and U5232 (N_5232,N_4701,N_4528);
or U5233 (N_5233,N_4387,N_4846);
nor U5234 (N_5234,N_4967,N_4910);
and U5235 (N_5235,N_4932,N_4168);
or U5236 (N_5236,N_4280,N_4126);
or U5237 (N_5237,N_4044,N_4496);
nor U5238 (N_5238,N_4372,N_4091);
or U5239 (N_5239,N_4711,N_4334);
nand U5240 (N_5240,N_4887,N_4849);
nand U5241 (N_5241,N_4443,N_4927);
nand U5242 (N_5242,N_4135,N_4451);
or U5243 (N_5243,N_4423,N_4996);
nor U5244 (N_5244,N_4458,N_4705);
xnor U5245 (N_5245,N_4100,N_4195);
nor U5246 (N_5246,N_4315,N_4245);
and U5247 (N_5247,N_4006,N_4002);
and U5248 (N_5248,N_4985,N_4302);
and U5249 (N_5249,N_4042,N_4066);
nor U5250 (N_5250,N_4232,N_4264);
nand U5251 (N_5251,N_4380,N_4651);
or U5252 (N_5252,N_4097,N_4355);
nand U5253 (N_5253,N_4223,N_4949);
nor U5254 (N_5254,N_4692,N_4841);
nor U5255 (N_5255,N_4406,N_4433);
nand U5256 (N_5256,N_4785,N_4052);
and U5257 (N_5257,N_4057,N_4477);
nor U5258 (N_5258,N_4084,N_4233);
and U5259 (N_5259,N_4336,N_4699);
or U5260 (N_5260,N_4305,N_4748);
and U5261 (N_5261,N_4808,N_4199);
or U5262 (N_5262,N_4351,N_4645);
and U5263 (N_5263,N_4804,N_4060);
xor U5264 (N_5264,N_4518,N_4228);
nand U5265 (N_5265,N_4307,N_4489);
and U5266 (N_5266,N_4295,N_4597);
and U5267 (N_5267,N_4193,N_4141);
or U5268 (N_5268,N_4736,N_4085);
and U5269 (N_5269,N_4983,N_4149);
nand U5270 (N_5270,N_4920,N_4529);
nor U5271 (N_5271,N_4374,N_4058);
nor U5272 (N_5272,N_4552,N_4740);
and U5273 (N_5273,N_4710,N_4046);
nor U5274 (N_5274,N_4667,N_4714);
and U5275 (N_5275,N_4234,N_4391);
nand U5276 (N_5276,N_4313,N_4471);
nand U5277 (N_5277,N_4083,N_4397);
nor U5278 (N_5278,N_4409,N_4206);
nand U5279 (N_5279,N_4127,N_4230);
or U5280 (N_5280,N_4790,N_4268);
nand U5281 (N_5281,N_4698,N_4216);
or U5282 (N_5282,N_4546,N_4294);
or U5283 (N_5283,N_4138,N_4136);
or U5284 (N_5284,N_4165,N_4227);
xnor U5285 (N_5285,N_4538,N_4997);
and U5286 (N_5286,N_4153,N_4860);
and U5287 (N_5287,N_4728,N_4913);
nor U5288 (N_5288,N_4207,N_4162);
nand U5289 (N_5289,N_4598,N_4146);
nor U5290 (N_5290,N_4134,N_4282);
and U5291 (N_5291,N_4637,N_4697);
or U5292 (N_5292,N_4321,N_4163);
and U5293 (N_5293,N_4739,N_4322);
or U5294 (N_5294,N_4318,N_4658);
nor U5295 (N_5295,N_4715,N_4148);
nor U5296 (N_5296,N_4194,N_4158);
nor U5297 (N_5297,N_4164,N_4800);
and U5298 (N_5298,N_4690,N_4049);
nand U5299 (N_5299,N_4364,N_4523);
nor U5300 (N_5300,N_4460,N_4089);
and U5301 (N_5301,N_4427,N_4908);
nor U5302 (N_5302,N_4831,N_4312);
or U5303 (N_5303,N_4991,N_4375);
and U5304 (N_5304,N_4792,N_4975);
and U5305 (N_5305,N_4686,N_4981);
or U5306 (N_5306,N_4122,N_4439);
and U5307 (N_5307,N_4619,N_4986);
nor U5308 (N_5308,N_4252,N_4086);
and U5309 (N_5309,N_4889,N_4903);
and U5310 (N_5310,N_4402,N_4438);
and U5311 (N_5311,N_4178,N_4945);
and U5312 (N_5312,N_4419,N_4922);
or U5313 (N_5313,N_4819,N_4532);
and U5314 (N_5314,N_4727,N_4326);
or U5315 (N_5315,N_4000,N_4405);
or U5316 (N_5316,N_4677,N_4937);
nor U5317 (N_5317,N_4881,N_4914);
nor U5318 (N_5318,N_4956,N_4011);
or U5319 (N_5319,N_4867,N_4311);
nor U5320 (N_5320,N_4636,N_4947);
or U5321 (N_5321,N_4139,N_4018);
or U5322 (N_5322,N_4273,N_4221);
and U5323 (N_5323,N_4338,N_4038);
or U5324 (N_5324,N_4150,N_4834);
or U5325 (N_5325,N_4071,N_4360);
nor U5326 (N_5326,N_4873,N_4465);
nand U5327 (N_5327,N_4670,N_4626);
nand U5328 (N_5328,N_4534,N_4843);
nor U5329 (N_5329,N_4494,N_4024);
and U5330 (N_5330,N_4357,N_4331);
and U5331 (N_5331,N_4671,N_4454);
nor U5332 (N_5332,N_4208,N_4200);
or U5333 (N_5333,N_4404,N_4788);
nor U5334 (N_5334,N_4899,N_4378);
and U5335 (N_5335,N_4554,N_4396);
and U5336 (N_5336,N_4824,N_4384);
and U5337 (N_5337,N_4377,N_4144);
nand U5338 (N_5338,N_4292,N_4553);
nand U5339 (N_5339,N_4657,N_4756);
or U5340 (N_5340,N_4580,N_4075);
nor U5341 (N_5341,N_4953,N_4664);
nand U5342 (N_5342,N_4385,N_4964);
and U5343 (N_5343,N_4483,N_4782);
nor U5344 (N_5344,N_4871,N_4300);
nor U5345 (N_5345,N_4156,N_4310);
nor U5346 (N_5346,N_4109,N_4716);
or U5347 (N_5347,N_4906,N_4124);
nand U5348 (N_5348,N_4995,N_4520);
or U5349 (N_5349,N_4823,N_4502);
nor U5350 (N_5350,N_4882,N_4972);
and U5351 (N_5351,N_4435,N_4766);
and U5352 (N_5352,N_4816,N_4306);
nor U5353 (N_5353,N_4432,N_4189);
or U5354 (N_5354,N_4839,N_4611);
or U5355 (N_5355,N_4845,N_4577);
or U5356 (N_5356,N_4050,N_4298);
nand U5357 (N_5357,N_4096,N_4815);
and U5358 (N_5358,N_4663,N_4863);
nor U5359 (N_5359,N_4484,N_4563);
and U5360 (N_5360,N_4401,N_4212);
nand U5361 (N_5361,N_4744,N_4053);
and U5362 (N_5362,N_4422,N_4838);
nand U5363 (N_5363,N_4487,N_4025);
and U5364 (N_5364,N_4912,N_4878);
nand U5365 (N_5365,N_4642,N_4497);
nor U5366 (N_5366,N_4065,N_4469);
nand U5367 (N_5367,N_4892,N_4467);
nand U5368 (N_5368,N_4549,N_4868);
or U5369 (N_5369,N_4631,N_4539);
xnor U5370 (N_5370,N_4630,N_4016);
or U5371 (N_5371,N_4370,N_4314);
nor U5372 (N_5372,N_4844,N_4989);
nand U5373 (N_5373,N_4159,N_4236);
xnor U5374 (N_5374,N_4449,N_4114);
and U5375 (N_5375,N_4110,N_4004);
nand U5376 (N_5376,N_4356,N_4576);
or U5377 (N_5377,N_4799,N_4246);
nor U5378 (N_5378,N_4880,N_4560);
nand U5379 (N_5379,N_4556,N_4934);
nand U5380 (N_5380,N_4814,N_4992);
xnor U5381 (N_5381,N_4584,N_4627);
or U5382 (N_5382,N_4647,N_4213);
nand U5383 (N_5383,N_4383,N_4190);
or U5384 (N_5384,N_4732,N_4768);
nor U5385 (N_5385,N_4607,N_4806);
nand U5386 (N_5386,N_4475,N_4909);
nor U5387 (N_5387,N_4713,N_4056);
and U5388 (N_5388,N_4265,N_4290);
and U5389 (N_5389,N_4151,N_4836);
or U5390 (N_5390,N_4481,N_4760);
nand U5391 (N_5391,N_4786,N_4673);
and U5392 (N_5392,N_4271,N_4608);
and U5393 (N_5393,N_4130,N_4131);
and U5394 (N_5394,N_4287,N_4107);
nand U5395 (N_5395,N_4850,N_4332);
xnor U5396 (N_5396,N_4616,N_4257);
or U5397 (N_5397,N_4741,N_4081);
nor U5398 (N_5398,N_4123,N_4327);
nand U5399 (N_5399,N_4840,N_4461);
and U5400 (N_5400,N_4474,N_4869);
nor U5401 (N_5401,N_4896,N_4825);
and U5402 (N_5402,N_4180,N_4279);
nand U5403 (N_5403,N_4541,N_4205);
nor U5404 (N_5404,N_4721,N_4063);
and U5405 (N_5405,N_4304,N_4833);
nor U5406 (N_5406,N_4291,N_4263);
nor U5407 (N_5407,N_4020,N_4262);
or U5408 (N_5408,N_4369,N_4023);
nand U5409 (N_5409,N_4359,N_4575);
and U5410 (N_5410,N_4343,N_4393);
nor U5411 (N_5411,N_4639,N_4695);
nand U5412 (N_5412,N_4612,N_4010);
or U5413 (N_5413,N_4285,N_4762);
nand U5414 (N_5414,N_4335,N_4087);
nand U5415 (N_5415,N_4119,N_4720);
and U5416 (N_5416,N_4558,N_4361);
nand U5417 (N_5417,N_4070,N_4751);
nor U5418 (N_5418,N_4507,N_4578);
or U5419 (N_5419,N_4725,N_4173);
or U5420 (N_5420,N_4408,N_4005);
or U5421 (N_5421,N_4470,N_4118);
and U5422 (N_5422,N_4068,N_4907);
and U5423 (N_5423,N_4723,N_4810);
nand U5424 (N_5424,N_4288,N_4472);
nand U5425 (N_5425,N_4102,N_4668);
nand U5426 (N_5426,N_4155,N_4961);
nand U5427 (N_5427,N_4094,N_4442);
nor U5428 (N_5428,N_4562,N_4499);
and U5429 (N_5429,N_4764,N_4724);
or U5430 (N_5430,N_4759,N_4333);
nor U5431 (N_5431,N_4254,N_4581);
or U5432 (N_5432,N_4407,N_4666);
nor U5433 (N_5433,N_4225,N_4958);
and U5434 (N_5434,N_4220,N_4933);
nor U5435 (N_5435,N_4172,N_4034);
nand U5436 (N_5436,N_4067,N_4077);
or U5437 (N_5437,N_4414,N_4852);
nor U5438 (N_5438,N_4032,N_4771);
nand U5439 (N_5439,N_4876,N_4459);
nor U5440 (N_5440,N_4436,N_4498);
nor U5441 (N_5441,N_4734,N_4450);
nand U5442 (N_5442,N_4284,N_4323);
and U5443 (N_5443,N_4772,N_4960);
nand U5444 (N_5444,N_4735,N_4516);
nand U5445 (N_5445,N_4918,N_4064);
nor U5446 (N_5446,N_4242,N_4202);
and U5447 (N_5447,N_4826,N_4798);
nand U5448 (N_5448,N_4473,N_4341);
nand U5449 (N_5449,N_4963,N_4737);
or U5450 (N_5450,N_4410,N_4614);
nand U5451 (N_5451,N_4625,N_4601);
and U5452 (N_5452,N_4921,N_4848);
or U5453 (N_5453,N_4425,N_4270);
nand U5454 (N_5454,N_4009,N_4968);
or U5455 (N_5455,N_4161,N_4689);
and U5456 (N_5456,N_4400,N_4412);
or U5457 (N_5457,N_4043,N_4593);
and U5458 (N_5458,N_4935,N_4485);
nor U5459 (N_5459,N_4572,N_4308);
nand U5460 (N_5460,N_4381,N_4915);
and U5461 (N_5461,N_4565,N_4342);
nor U5462 (N_5462,N_4990,N_4061);
or U5463 (N_5463,N_4632,N_4780);
nand U5464 (N_5464,N_4229,N_4031);
and U5465 (N_5465,N_4624,N_4108);
and U5466 (N_5466,N_4105,N_4568);
and U5467 (N_5467,N_4749,N_4309);
nand U5468 (N_5468,N_4767,N_4811);
and U5469 (N_5469,N_4745,N_4665);
and U5470 (N_5470,N_4752,N_4428);
and U5471 (N_5471,N_4269,N_4388);
nand U5472 (N_5472,N_4571,N_4687);
and U5473 (N_5473,N_4957,N_4613);
nand U5474 (N_5474,N_4511,N_4281);
or U5475 (N_5475,N_4680,N_4898);
nand U5476 (N_5476,N_4140,N_4379);
nor U5477 (N_5477,N_4629,N_4726);
nand U5478 (N_5478,N_4092,N_4861);
and U5479 (N_5479,N_4440,N_4417);
or U5480 (N_5480,N_4143,N_4801);
and U5481 (N_5481,N_4722,N_4596);
nand U5482 (N_5482,N_4820,N_4015);
nand U5483 (N_5483,N_4463,N_4924);
and U5484 (N_5484,N_4644,N_4259);
and U5485 (N_5485,N_4297,N_4890);
nand U5486 (N_5486,N_4008,N_4187);
nand U5487 (N_5487,N_4235,N_4059);
and U5488 (N_5488,N_4755,N_4389);
or U5489 (N_5489,N_4353,N_4261);
nor U5490 (N_5490,N_4813,N_4366);
or U5491 (N_5491,N_4928,N_4978);
nand U5492 (N_5492,N_4900,N_4592);
nand U5493 (N_5493,N_4544,N_4434);
or U5494 (N_5494,N_4674,N_4197);
and U5495 (N_5495,N_4588,N_4602);
and U5496 (N_5496,N_4431,N_4807);
xor U5497 (N_5497,N_4948,N_4441);
and U5498 (N_5498,N_4977,N_4055);
nand U5499 (N_5499,N_4030,N_4946);
nand U5500 (N_5500,N_4128,N_4552);
nor U5501 (N_5501,N_4081,N_4487);
and U5502 (N_5502,N_4773,N_4778);
nor U5503 (N_5503,N_4922,N_4354);
and U5504 (N_5504,N_4614,N_4227);
nor U5505 (N_5505,N_4919,N_4136);
and U5506 (N_5506,N_4963,N_4771);
nand U5507 (N_5507,N_4685,N_4511);
and U5508 (N_5508,N_4268,N_4538);
and U5509 (N_5509,N_4777,N_4505);
nor U5510 (N_5510,N_4627,N_4125);
nand U5511 (N_5511,N_4039,N_4033);
nor U5512 (N_5512,N_4182,N_4454);
or U5513 (N_5513,N_4438,N_4672);
nor U5514 (N_5514,N_4009,N_4530);
nand U5515 (N_5515,N_4693,N_4604);
and U5516 (N_5516,N_4401,N_4366);
or U5517 (N_5517,N_4918,N_4285);
and U5518 (N_5518,N_4580,N_4955);
nor U5519 (N_5519,N_4577,N_4522);
nor U5520 (N_5520,N_4267,N_4338);
nor U5521 (N_5521,N_4873,N_4308);
or U5522 (N_5522,N_4729,N_4261);
nor U5523 (N_5523,N_4586,N_4925);
and U5524 (N_5524,N_4683,N_4030);
nand U5525 (N_5525,N_4203,N_4772);
nand U5526 (N_5526,N_4191,N_4250);
and U5527 (N_5527,N_4958,N_4548);
nor U5528 (N_5528,N_4994,N_4749);
nor U5529 (N_5529,N_4541,N_4976);
nor U5530 (N_5530,N_4853,N_4477);
or U5531 (N_5531,N_4489,N_4513);
nand U5532 (N_5532,N_4131,N_4929);
nor U5533 (N_5533,N_4878,N_4686);
or U5534 (N_5534,N_4814,N_4114);
nor U5535 (N_5535,N_4465,N_4392);
nand U5536 (N_5536,N_4029,N_4473);
or U5537 (N_5537,N_4241,N_4097);
or U5538 (N_5538,N_4153,N_4729);
nand U5539 (N_5539,N_4772,N_4215);
nand U5540 (N_5540,N_4789,N_4487);
nor U5541 (N_5541,N_4473,N_4761);
nor U5542 (N_5542,N_4282,N_4541);
nand U5543 (N_5543,N_4140,N_4503);
nor U5544 (N_5544,N_4129,N_4602);
nand U5545 (N_5545,N_4931,N_4620);
nor U5546 (N_5546,N_4108,N_4883);
nand U5547 (N_5547,N_4923,N_4599);
nor U5548 (N_5548,N_4769,N_4094);
nand U5549 (N_5549,N_4804,N_4809);
nand U5550 (N_5550,N_4984,N_4927);
nand U5551 (N_5551,N_4940,N_4544);
and U5552 (N_5552,N_4476,N_4715);
or U5553 (N_5553,N_4769,N_4882);
nand U5554 (N_5554,N_4849,N_4153);
nand U5555 (N_5555,N_4068,N_4047);
or U5556 (N_5556,N_4685,N_4983);
or U5557 (N_5557,N_4297,N_4884);
nor U5558 (N_5558,N_4834,N_4781);
xnor U5559 (N_5559,N_4070,N_4861);
nor U5560 (N_5560,N_4589,N_4217);
and U5561 (N_5561,N_4673,N_4861);
and U5562 (N_5562,N_4872,N_4791);
nor U5563 (N_5563,N_4679,N_4843);
nor U5564 (N_5564,N_4162,N_4268);
and U5565 (N_5565,N_4708,N_4710);
and U5566 (N_5566,N_4520,N_4726);
nand U5567 (N_5567,N_4490,N_4029);
and U5568 (N_5568,N_4437,N_4449);
nor U5569 (N_5569,N_4990,N_4017);
and U5570 (N_5570,N_4946,N_4343);
nand U5571 (N_5571,N_4967,N_4659);
nand U5572 (N_5572,N_4439,N_4815);
or U5573 (N_5573,N_4985,N_4407);
nor U5574 (N_5574,N_4194,N_4497);
and U5575 (N_5575,N_4532,N_4729);
nor U5576 (N_5576,N_4761,N_4348);
nand U5577 (N_5577,N_4375,N_4497);
nor U5578 (N_5578,N_4608,N_4748);
or U5579 (N_5579,N_4321,N_4277);
or U5580 (N_5580,N_4810,N_4287);
or U5581 (N_5581,N_4306,N_4436);
nand U5582 (N_5582,N_4036,N_4136);
nand U5583 (N_5583,N_4461,N_4073);
or U5584 (N_5584,N_4136,N_4691);
and U5585 (N_5585,N_4508,N_4857);
or U5586 (N_5586,N_4136,N_4435);
and U5587 (N_5587,N_4008,N_4546);
nand U5588 (N_5588,N_4901,N_4441);
or U5589 (N_5589,N_4290,N_4053);
and U5590 (N_5590,N_4300,N_4868);
or U5591 (N_5591,N_4210,N_4009);
nor U5592 (N_5592,N_4579,N_4184);
nor U5593 (N_5593,N_4315,N_4288);
or U5594 (N_5594,N_4443,N_4026);
nand U5595 (N_5595,N_4314,N_4713);
nand U5596 (N_5596,N_4612,N_4941);
nand U5597 (N_5597,N_4387,N_4843);
or U5598 (N_5598,N_4117,N_4981);
or U5599 (N_5599,N_4223,N_4143);
and U5600 (N_5600,N_4563,N_4098);
nor U5601 (N_5601,N_4879,N_4814);
nand U5602 (N_5602,N_4402,N_4464);
or U5603 (N_5603,N_4339,N_4665);
and U5604 (N_5604,N_4143,N_4235);
nand U5605 (N_5605,N_4340,N_4259);
nand U5606 (N_5606,N_4497,N_4407);
and U5607 (N_5607,N_4802,N_4761);
xnor U5608 (N_5608,N_4862,N_4707);
nor U5609 (N_5609,N_4124,N_4688);
and U5610 (N_5610,N_4824,N_4635);
and U5611 (N_5611,N_4480,N_4463);
and U5612 (N_5612,N_4158,N_4439);
nor U5613 (N_5613,N_4766,N_4436);
nand U5614 (N_5614,N_4302,N_4955);
nand U5615 (N_5615,N_4503,N_4249);
and U5616 (N_5616,N_4965,N_4180);
or U5617 (N_5617,N_4614,N_4438);
nor U5618 (N_5618,N_4149,N_4930);
or U5619 (N_5619,N_4082,N_4785);
or U5620 (N_5620,N_4967,N_4004);
nor U5621 (N_5621,N_4140,N_4648);
xnor U5622 (N_5622,N_4623,N_4850);
nor U5623 (N_5623,N_4303,N_4893);
nand U5624 (N_5624,N_4697,N_4923);
nand U5625 (N_5625,N_4504,N_4584);
and U5626 (N_5626,N_4167,N_4314);
nand U5627 (N_5627,N_4562,N_4353);
and U5628 (N_5628,N_4951,N_4935);
nand U5629 (N_5629,N_4863,N_4488);
nor U5630 (N_5630,N_4136,N_4849);
and U5631 (N_5631,N_4038,N_4867);
and U5632 (N_5632,N_4414,N_4382);
and U5633 (N_5633,N_4637,N_4404);
or U5634 (N_5634,N_4940,N_4027);
and U5635 (N_5635,N_4038,N_4114);
nand U5636 (N_5636,N_4681,N_4927);
or U5637 (N_5637,N_4187,N_4534);
or U5638 (N_5638,N_4256,N_4472);
nand U5639 (N_5639,N_4069,N_4163);
or U5640 (N_5640,N_4331,N_4737);
nor U5641 (N_5641,N_4007,N_4855);
nor U5642 (N_5642,N_4874,N_4431);
and U5643 (N_5643,N_4682,N_4926);
and U5644 (N_5644,N_4012,N_4738);
nand U5645 (N_5645,N_4795,N_4048);
and U5646 (N_5646,N_4996,N_4550);
or U5647 (N_5647,N_4137,N_4129);
nor U5648 (N_5648,N_4270,N_4830);
xnor U5649 (N_5649,N_4788,N_4895);
nand U5650 (N_5650,N_4488,N_4063);
nand U5651 (N_5651,N_4372,N_4346);
and U5652 (N_5652,N_4858,N_4539);
and U5653 (N_5653,N_4493,N_4806);
or U5654 (N_5654,N_4311,N_4588);
nand U5655 (N_5655,N_4887,N_4745);
nand U5656 (N_5656,N_4935,N_4118);
and U5657 (N_5657,N_4003,N_4154);
nand U5658 (N_5658,N_4836,N_4558);
or U5659 (N_5659,N_4709,N_4756);
nand U5660 (N_5660,N_4343,N_4257);
nand U5661 (N_5661,N_4782,N_4706);
nor U5662 (N_5662,N_4995,N_4543);
nor U5663 (N_5663,N_4656,N_4697);
and U5664 (N_5664,N_4678,N_4206);
or U5665 (N_5665,N_4070,N_4626);
and U5666 (N_5666,N_4920,N_4549);
or U5667 (N_5667,N_4093,N_4964);
or U5668 (N_5668,N_4161,N_4223);
or U5669 (N_5669,N_4365,N_4319);
xnor U5670 (N_5670,N_4297,N_4639);
nor U5671 (N_5671,N_4014,N_4123);
and U5672 (N_5672,N_4680,N_4271);
or U5673 (N_5673,N_4456,N_4169);
nand U5674 (N_5674,N_4647,N_4508);
nor U5675 (N_5675,N_4230,N_4800);
nor U5676 (N_5676,N_4179,N_4679);
nor U5677 (N_5677,N_4771,N_4764);
and U5678 (N_5678,N_4081,N_4550);
or U5679 (N_5679,N_4145,N_4437);
nor U5680 (N_5680,N_4730,N_4145);
and U5681 (N_5681,N_4860,N_4623);
or U5682 (N_5682,N_4680,N_4836);
nor U5683 (N_5683,N_4170,N_4016);
nor U5684 (N_5684,N_4630,N_4939);
and U5685 (N_5685,N_4790,N_4109);
nand U5686 (N_5686,N_4713,N_4122);
and U5687 (N_5687,N_4483,N_4252);
nand U5688 (N_5688,N_4250,N_4170);
or U5689 (N_5689,N_4393,N_4768);
and U5690 (N_5690,N_4267,N_4554);
nand U5691 (N_5691,N_4290,N_4622);
or U5692 (N_5692,N_4491,N_4961);
or U5693 (N_5693,N_4273,N_4725);
or U5694 (N_5694,N_4525,N_4764);
and U5695 (N_5695,N_4959,N_4778);
nand U5696 (N_5696,N_4751,N_4185);
or U5697 (N_5697,N_4127,N_4539);
and U5698 (N_5698,N_4937,N_4599);
nand U5699 (N_5699,N_4252,N_4288);
nor U5700 (N_5700,N_4038,N_4805);
nand U5701 (N_5701,N_4217,N_4740);
or U5702 (N_5702,N_4944,N_4907);
nand U5703 (N_5703,N_4063,N_4263);
nand U5704 (N_5704,N_4158,N_4387);
nand U5705 (N_5705,N_4917,N_4066);
xnor U5706 (N_5706,N_4811,N_4141);
or U5707 (N_5707,N_4381,N_4600);
nand U5708 (N_5708,N_4496,N_4766);
nor U5709 (N_5709,N_4926,N_4694);
or U5710 (N_5710,N_4786,N_4232);
or U5711 (N_5711,N_4678,N_4886);
or U5712 (N_5712,N_4174,N_4097);
and U5713 (N_5713,N_4193,N_4798);
and U5714 (N_5714,N_4191,N_4242);
and U5715 (N_5715,N_4996,N_4140);
or U5716 (N_5716,N_4587,N_4350);
nand U5717 (N_5717,N_4065,N_4795);
or U5718 (N_5718,N_4029,N_4890);
or U5719 (N_5719,N_4836,N_4047);
or U5720 (N_5720,N_4744,N_4952);
nand U5721 (N_5721,N_4898,N_4424);
nand U5722 (N_5722,N_4562,N_4737);
nor U5723 (N_5723,N_4538,N_4641);
or U5724 (N_5724,N_4846,N_4670);
nor U5725 (N_5725,N_4500,N_4980);
xor U5726 (N_5726,N_4348,N_4587);
nor U5727 (N_5727,N_4727,N_4233);
and U5728 (N_5728,N_4341,N_4889);
and U5729 (N_5729,N_4387,N_4324);
or U5730 (N_5730,N_4449,N_4637);
nand U5731 (N_5731,N_4835,N_4779);
and U5732 (N_5732,N_4552,N_4441);
nand U5733 (N_5733,N_4855,N_4026);
nor U5734 (N_5734,N_4483,N_4070);
or U5735 (N_5735,N_4176,N_4623);
and U5736 (N_5736,N_4406,N_4031);
nand U5737 (N_5737,N_4021,N_4689);
nor U5738 (N_5738,N_4637,N_4761);
nor U5739 (N_5739,N_4209,N_4700);
nand U5740 (N_5740,N_4176,N_4638);
or U5741 (N_5741,N_4602,N_4950);
and U5742 (N_5742,N_4230,N_4174);
and U5743 (N_5743,N_4697,N_4179);
nor U5744 (N_5744,N_4003,N_4422);
nor U5745 (N_5745,N_4682,N_4382);
and U5746 (N_5746,N_4401,N_4111);
nor U5747 (N_5747,N_4345,N_4489);
nor U5748 (N_5748,N_4657,N_4141);
nor U5749 (N_5749,N_4527,N_4326);
nand U5750 (N_5750,N_4884,N_4803);
or U5751 (N_5751,N_4488,N_4396);
or U5752 (N_5752,N_4603,N_4043);
or U5753 (N_5753,N_4884,N_4377);
or U5754 (N_5754,N_4653,N_4683);
nor U5755 (N_5755,N_4081,N_4250);
and U5756 (N_5756,N_4105,N_4491);
and U5757 (N_5757,N_4575,N_4969);
and U5758 (N_5758,N_4622,N_4533);
or U5759 (N_5759,N_4981,N_4404);
and U5760 (N_5760,N_4092,N_4021);
nand U5761 (N_5761,N_4220,N_4084);
nand U5762 (N_5762,N_4043,N_4335);
nor U5763 (N_5763,N_4410,N_4947);
and U5764 (N_5764,N_4814,N_4231);
nand U5765 (N_5765,N_4971,N_4440);
or U5766 (N_5766,N_4484,N_4493);
nor U5767 (N_5767,N_4369,N_4391);
or U5768 (N_5768,N_4809,N_4805);
and U5769 (N_5769,N_4447,N_4844);
nor U5770 (N_5770,N_4575,N_4917);
xnor U5771 (N_5771,N_4524,N_4311);
or U5772 (N_5772,N_4228,N_4702);
nor U5773 (N_5773,N_4253,N_4127);
and U5774 (N_5774,N_4067,N_4580);
and U5775 (N_5775,N_4959,N_4554);
nand U5776 (N_5776,N_4955,N_4443);
and U5777 (N_5777,N_4761,N_4975);
and U5778 (N_5778,N_4882,N_4825);
and U5779 (N_5779,N_4340,N_4183);
nand U5780 (N_5780,N_4516,N_4705);
or U5781 (N_5781,N_4000,N_4276);
nor U5782 (N_5782,N_4326,N_4980);
and U5783 (N_5783,N_4091,N_4476);
nor U5784 (N_5784,N_4512,N_4697);
nor U5785 (N_5785,N_4378,N_4044);
and U5786 (N_5786,N_4555,N_4299);
nor U5787 (N_5787,N_4962,N_4305);
nand U5788 (N_5788,N_4923,N_4789);
or U5789 (N_5789,N_4181,N_4099);
nand U5790 (N_5790,N_4699,N_4980);
or U5791 (N_5791,N_4260,N_4162);
or U5792 (N_5792,N_4749,N_4561);
nor U5793 (N_5793,N_4309,N_4102);
nor U5794 (N_5794,N_4367,N_4178);
or U5795 (N_5795,N_4299,N_4545);
or U5796 (N_5796,N_4030,N_4773);
and U5797 (N_5797,N_4383,N_4835);
or U5798 (N_5798,N_4407,N_4270);
and U5799 (N_5799,N_4486,N_4966);
nor U5800 (N_5800,N_4963,N_4686);
nor U5801 (N_5801,N_4499,N_4736);
and U5802 (N_5802,N_4935,N_4686);
nor U5803 (N_5803,N_4112,N_4603);
or U5804 (N_5804,N_4995,N_4868);
nand U5805 (N_5805,N_4955,N_4095);
or U5806 (N_5806,N_4894,N_4194);
or U5807 (N_5807,N_4803,N_4324);
and U5808 (N_5808,N_4157,N_4011);
nand U5809 (N_5809,N_4037,N_4291);
nand U5810 (N_5810,N_4881,N_4903);
nand U5811 (N_5811,N_4419,N_4676);
nand U5812 (N_5812,N_4706,N_4636);
nor U5813 (N_5813,N_4001,N_4881);
nand U5814 (N_5814,N_4689,N_4187);
or U5815 (N_5815,N_4495,N_4709);
or U5816 (N_5816,N_4184,N_4434);
nand U5817 (N_5817,N_4211,N_4708);
and U5818 (N_5818,N_4539,N_4060);
nand U5819 (N_5819,N_4482,N_4055);
or U5820 (N_5820,N_4130,N_4812);
and U5821 (N_5821,N_4097,N_4292);
or U5822 (N_5822,N_4151,N_4512);
or U5823 (N_5823,N_4838,N_4910);
nor U5824 (N_5824,N_4542,N_4064);
nor U5825 (N_5825,N_4059,N_4653);
nand U5826 (N_5826,N_4280,N_4092);
nand U5827 (N_5827,N_4483,N_4104);
and U5828 (N_5828,N_4005,N_4911);
or U5829 (N_5829,N_4530,N_4110);
nand U5830 (N_5830,N_4894,N_4799);
nand U5831 (N_5831,N_4962,N_4975);
and U5832 (N_5832,N_4605,N_4345);
and U5833 (N_5833,N_4765,N_4194);
nor U5834 (N_5834,N_4512,N_4598);
xor U5835 (N_5835,N_4111,N_4101);
nor U5836 (N_5836,N_4217,N_4853);
and U5837 (N_5837,N_4555,N_4027);
or U5838 (N_5838,N_4656,N_4240);
or U5839 (N_5839,N_4126,N_4284);
nor U5840 (N_5840,N_4162,N_4602);
nand U5841 (N_5841,N_4624,N_4823);
nor U5842 (N_5842,N_4335,N_4784);
and U5843 (N_5843,N_4285,N_4150);
nand U5844 (N_5844,N_4235,N_4779);
nand U5845 (N_5845,N_4898,N_4651);
and U5846 (N_5846,N_4966,N_4762);
and U5847 (N_5847,N_4804,N_4664);
and U5848 (N_5848,N_4067,N_4908);
or U5849 (N_5849,N_4354,N_4182);
and U5850 (N_5850,N_4224,N_4025);
nand U5851 (N_5851,N_4045,N_4377);
and U5852 (N_5852,N_4033,N_4299);
xnor U5853 (N_5853,N_4068,N_4689);
nand U5854 (N_5854,N_4782,N_4542);
and U5855 (N_5855,N_4159,N_4190);
or U5856 (N_5856,N_4899,N_4420);
nor U5857 (N_5857,N_4121,N_4437);
or U5858 (N_5858,N_4465,N_4794);
nor U5859 (N_5859,N_4928,N_4004);
and U5860 (N_5860,N_4776,N_4585);
nand U5861 (N_5861,N_4375,N_4828);
and U5862 (N_5862,N_4557,N_4058);
and U5863 (N_5863,N_4051,N_4136);
and U5864 (N_5864,N_4337,N_4161);
and U5865 (N_5865,N_4737,N_4693);
or U5866 (N_5866,N_4594,N_4343);
nor U5867 (N_5867,N_4581,N_4543);
or U5868 (N_5868,N_4313,N_4865);
and U5869 (N_5869,N_4658,N_4379);
xor U5870 (N_5870,N_4496,N_4347);
nor U5871 (N_5871,N_4580,N_4950);
nand U5872 (N_5872,N_4046,N_4200);
and U5873 (N_5873,N_4823,N_4284);
nor U5874 (N_5874,N_4835,N_4522);
or U5875 (N_5875,N_4638,N_4778);
nor U5876 (N_5876,N_4931,N_4672);
nand U5877 (N_5877,N_4790,N_4394);
nand U5878 (N_5878,N_4336,N_4672);
nand U5879 (N_5879,N_4694,N_4621);
or U5880 (N_5880,N_4512,N_4733);
nor U5881 (N_5881,N_4676,N_4443);
nor U5882 (N_5882,N_4967,N_4786);
and U5883 (N_5883,N_4525,N_4376);
xnor U5884 (N_5884,N_4231,N_4153);
nor U5885 (N_5885,N_4907,N_4925);
or U5886 (N_5886,N_4582,N_4400);
and U5887 (N_5887,N_4361,N_4214);
nor U5888 (N_5888,N_4884,N_4861);
or U5889 (N_5889,N_4696,N_4011);
nand U5890 (N_5890,N_4520,N_4446);
nand U5891 (N_5891,N_4855,N_4439);
and U5892 (N_5892,N_4726,N_4064);
and U5893 (N_5893,N_4868,N_4915);
nor U5894 (N_5894,N_4225,N_4270);
nor U5895 (N_5895,N_4131,N_4047);
or U5896 (N_5896,N_4747,N_4420);
nor U5897 (N_5897,N_4594,N_4452);
or U5898 (N_5898,N_4729,N_4369);
nor U5899 (N_5899,N_4695,N_4039);
and U5900 (N_5900,N_4605,N_4560);
and U5901 (N_5901,N_4171,N_4639);
and U5902 (N_5902,N_4495,N_4844);
and U5903 (N_5903,N_4580,N_4442);
nand U5904 (N_5904,N_4194,N_4586);
and U5905 (N_5905,N_4143,N_4825);
or U5906 (N_5906,N_4918,N_4778);
and U5907 (N_5907,N_4470,N_4754);
or U5908 (N_5908,N_4870,N_4516);
nor U5909 (N_5909,N_4355,N_4509);
nor U5910 (N_5910,N_4491,N_4932);
and U5911 (N_5911,N_4585,N_4330);
nand U5912 (N_5912,N_4874,N_4737);
nor U5913 (N_5913,N_4220,N_4296);
nor U5914 (N_5914,N_4808,N_4175);
nor U5915 (N_5915,N_4934,N_4175);
and U5916 (N_5916,N_4126,N_4903);
nand U5917 (N_5917,N_4315,N_4028);
and U5918 (N_5918,N_4311,N_4509);
or U5919 (N_5919,N_4574,N_4712);
nor U5920 (N_5920,N_4950,N_4655);
or U5921 (N_5921,N_4405,N_4764);
or U5922 (N_5922,N_4893,N_4275);
or U5923 (N_5923,N_4953,N_4094);
nor U5924 (N_5924,N_4980,N_4183);
nand U5925 (N_5925,N_4614,N_4228);
nand U5926 (N_5926,N_4468,N_4779);
nor U5927 (N_5927,N_4565,N_4682);
or U5928 (N_5928,N_4523,N_4598);
and U5929 (N_5929,N_4297,N_4716);
nand U5930 (N_5930,N_4484,N_4198);
and U5931 (N_5931,N_4269,N_4370);
nand U5932 (N_5932,N_4430,N_4052);
and U5933 (N_5933,N_4854,N_4082);
nor U5934 (N_5934,N_4540,N_4843);
or U5935 (N_5935,N_4036,N_4753);
nor U5936 (N_5936,N_4094,N_4798);
nor U5937 (N_5937,N_4043,N_4972);
nand U5938 (N_5938,N_4978,N_4624);
nor U5939 (N_5939,N_4917,N_4127);
nand U5940 (N_5940,N_4897,N_4092);
nor U5941 (N_5941,N_4171,N_4628);
and U5942 (N_5942,N_4776,N_4349);
nand U5943 (N_5943,N_4850,N_4447);
nand U5944 (N_5944,N_4726,N_4960);
nand U5945 (N_5945,N_4085,N_4033);
nor U5946 (N_5946,N_4267,N_4772);
nor U5947 (N_5947,N_4768,N_4917);
and U5948 (N_5948,N_4151,N_4825);
and U5949 (N_5949,N_4668,N_4877);
nand U5950 (N_5950,N_4002,N_4139);
nand U5951 (N_5951,N_4050,N_4765);
and U5952 (N_5952,N_4080,N_4428);
nor U5953 (N_5953,N_4169,N_4572);
and U5954 (N_5954,N_4649,N_4887);
and U5955 (N_5955,N_4159,N_4089);
or U5956 (N_5956,N_4315,N_4117);
nand U5957 (N_5957,N_4297,N_4908);
and U5958 (N_5958,N_4320,N_4203);
xnor U5959 (N_5959,N_4813,N_4799);
and U5960 (N_5960,N_4519,N_4017);
and U5961 (N_5961,N_4024,N_4373);
nor U5962 (N_5962,N_4856,N_4699);
nand U5963 (N_5963,N_4578,N_4567);
xor U5964 (N_5964,N_4968,N_4973);
and U5965 (N_5965,N_4163,N_4565);
nand U5966 (N_5966,N_4818,N_4374);
nor U5967 (N_5967,N_4110,N_4702);
or U5968 (N_5968,N_4342,N_4137);
and U5969 (N_5969,N_4613,N_4181);
or U5970 (N_5970,N_4684,N_4223);
xnor U5971 (N_5971,N_4711,N_4167);
and U5972 (N_5972,N_4744,N_4715);
nor U5973 (N_5973,N_4648,N_4351);
or U5974 (N_5974,N_4553,N_4694);
or U5975 (N_5975,N_4463,N_4049);
nand U5976 (N_5976,N_4612,N_4766);
nand U5977 (N_5977,N_4748,N_4812);
or U5978 (N_5978,N_4627,N_4384);
or U5979 (N_5979,N_4671,N_4159);
or U5980 (N_5980,N_4301,N_4516);
or U5981 (N_5981,N_4116,N_4054);
nor U5982 (N_5982,N_4051,N_4646);
and U5983 (N_5983,N_4535,N_4496);
and U5984 (N_5984,N_4316,N_4351);
nand U5985 (N_5985,N_4192,N_4228);
or U5986 (N_5986,N_4964,N_4424);
nor U5987 (N_5987,N_4220,N_4026);
nand U5988 (N_5988,N_4625,N_4723);
nor U5989 (N_5989,N_4966,N_4201);
or U5990 (N_5990,N_4941,N_4916);
and U5991 (N_5991,N_4105,N_4040);
nor U5992 (N_5992,N_4665,N_4286);
xor U5993 (N_5993,N_4398,N_4918);
nand U5994 (N_5994,N_4032,N_4606);
nand U5995 (N_5995,N_4238,N_4668);
nand U5996 (N_5996,N_4783,N_4791);
nor U5997 (N_5997,N_4817,N_4405);
nand U5998 (N_5998,N_4498,N_4685);
and U5999 (N_5999,N_4168,N_4516);
nor U6000 (N_6000,N_5278,N_5690);
nand U6001 (N_6001,N_5955,N_5635);
and U6002 (N_6002,N_5454,N_5292);
and U6003 (N_6003,N_5648,N_5765);
and U6004 (N_6004,N_5423,N_5298);
nor U6005 (N_6005,N_5798,N_5311);
nor U6006 (N_6006,N_5343,N_5205);
nor U6007 (N_6007,N_5115,N_5669);
or U6008 (N_6008,N_5850,N_5450);
nand U6009 (N_6009,N_5312,N_5168);
nand U6010 (N_6010,N_5513,N_5891);
nand U6011 (N_6011,N_5439,N_5862);
nor U6012 (N_6012,N_5794,N_5724);
nand U6013 (N_6013,N_5252,N_5504);
and U6014 (N_6014,N_5321,N_5649);
and U6015 (N_6015,N_5553,N_5038);
and U6016 (N_6016,N_5296,N_5314);
nand U6017 (N_6017,N_5271,N_5385);
nor U6018 (N_6018,N_5554,N_5240);
and U6019 (N_6019,N_5814,N_5355);
and U6020 (N_6020,N_5297,N_5847);
nor U6021 (N_6021,N_5592,N_5490);
or U6022 (N_6022,N_5294,N_5566);
nand U6023 (N_6023,N_5942,N_5221);
or U6024 (N_6024,N_5101,N_5604);
and U6025 (N_6025,N_5744,N_5144);
nand U6026 (N_6026,N_5208,N_5791);
nand U6027 (N_6027,N_5920,N_5949);
nand U6028 (N_6028,N_5228,N_5611);
and U6029 (N_6029,N_5188,N_5515);
nand U6030 (N_6030,N_5393,N_5528);
and U6031 (N_6031,N_5280,N_5370);
or U6032 (N_6032,N_5526,N_5615);
nand U6033 (N_6033,N_5735,N_5276);
nand U6034 (N_6034,N_5756,N_5825);
or U6035 (N_6035,N_5728,N_5895);
nand U6036 (N_6036,N_5236,N_5265);
and U6037 (N_6037,N_5331,N_5054);
nor U6038 (N_6038,N_5471,N_5281);
and U6039 (N_6039,N_5667,N_5868);
nor U6040 (N_6040,N_5535,N_5532);
and U6041 (N_6041,N_5948,N_5935);
and U6042 (N_6042,N_5346,N_5788);
nor U6043 (N_6043,N_5670,N_5086);
nand U6044 (N_6044,N_5692,N_5557);
or U6045 (N_6045,N_5361,N_5016);
nor U6046 (N_6046,N_5516,N_5063);
or U6047 (N_6047,N_5755,N_5246);
nor U6048 (N_6048,N_5618,N_5636);
and U6049 (N_6049,N_5059,N_5448);
nand U6050 (N_6050,N_5770,N_5190);
and U6051 (N_6051,N_5123,N_5134);
and U6052 (N_6052,N_5107,N_5045);
and U6053 (N_6053,N_5926,N_5625);
nor U6054 (N_6054,N_5679,N_5778);
and U6055 (N_6055,N_5324,N_5646);
or U6056 (N_6056,N_5266,N_5198);
and U6057 (N_6057,N_5110,N_5033);
or U6058 (N_6058,N_5902,N_5395);
nand U6059 (N_6059,N_5588,N_5282);
or U6060 (N_6060,N_5180,N_5815);
nand U6061 (N_6061,N_5397,N_5118);
nand U6062 (N_6062,N_5167,N_5460);
and U6063 (N_6063,N_5351,N_5472);
or U6064 (N_6064,N_5170,N_5155);
nor U6065 (N_6065,N_5384,N_5512);
or U6066 (N_6066,N_5913,N_5817);
or U6067 (N_6067,N_5436,N_5438);
xnor U6068 (N_6068,N_5598,N_5412);
or U6069 (N_6069,N_5032,N_5995);
nor U6070 (N_6070,N_5863,N_5582);
nor U6071 (N_6071,N_5737,N_5521);
and U6072 (N_6072,N_5373,N_5947);
or U6073 (N_6073,N_5605,N_5458);
nand U6074 (N_6074,N_5142,N_5488);
nor U6075 (N_6075,N_5821,N_5199);
or U6076 (N_6076,N_5394,N_5042);
nor U6077 (N_6077,N_5225,N_5399);
and U6078 (N_6078,N_5507,N_5034);
xor U6079 (N_6079,N_5781,N_5166);
nand U6080 (N_6080,N_5174,N_5970);
nand U6081 (N_6081,N_5259,N_5882);
and U6082 (N_6082,N_5641,N_5435);
and U6083 (N_6083,N_5591,N_5991);
and U6084 (N_6084,N_5226,N_5456);
nor U6085 (N_6085,N_5733,N_5748);
or U6086 (N_6086,N_5322,N_5335);
nor U6087 (N_6087,N_5011,N_5017);
nor U6088 (N_6088,N_5015,N_5466);
and U6089 (N_6089,N_5342,N_5639);
nand U6090 (N_6090,N_5129,N_5723);
or U6091 (N_6091,N_5684,N_5631);
nor U6092 (N_6092,N_5905,N_5746);
or U6093 (N_6093,N_5884,N_5317);
and U6094 (N_6094,N_5579,N_5476);
nor U6095 (N_6095,N_5043,N_5302);
or U6096 (N_6096,N_5481,N_5119);
nor U6097 (N_6097,N_5090,N_5194);
and U6098 (N_6098,N_5382,N_5802);
nor U6099 (N_6099,N_5409,N_5457);
nor U6100 (N_6100,N_5116,N_5820);
or U6101 (N_6101,N_5900,N_5009);
nand U6102 (N_6102,N_5874,N_5293);
and U6103 (N_6103,N_5416,N_5067);
nand U6104 (N_6104,N_5734,N_5918);
nand U6105 (N_6105,N_5562,N_5289);
xor U6106 (N_6106,N_5889,N_5286);
nand U6107 (N_6107,N_5538,N_5068);
and U6108 (N_6108,N_5818,N_5697);
and U6109 (N_6109,N_5328,N_5517);
or U6110 (N_6110,N_5223,N_5131);
nor U6111 (N_6111,N_5376,N_5400);
or U6112 (N_6112,N_5719,N_5359);
nand U6113 (N_6113,N_5721,N_5089);
or U6114 (N_6114,N_5795,N_5607);
nor U6115 (N_6115,N_5944,N_5767);
nand U6116 (N_6116,N_5864,N_5299);
and U6117 (N_6117,N_5122,N_5430);
nor U6118 (N_6118,N_5994,N_5157);
or U6119 (N_6119,N_5374,N_5603);
and U6120 (N_6120,N_5128,N_5206);
and U6121 (N_6121,N_5903,N_5961);
or U6122 (N_6122,N_5686,N_5834);
and U6123 (N_6123,N_5921,N_5711);
nand U6124 (N_6124,N_5638,N_5838);
and U6125 (N_6125,N_5586,N_5567);
or U6126 (N_6126,N_5565,N_5674);
or U6127 (N_6127,N_5764,N_5845);
nand U6128 (N_6128,N_5387,N_5079);
nor U6129 (N_6129,N_5161,N_5685);
nand U6130 (N_6130,N_5572,N_5185);
nand U6131 (N_6131,N_5839,N_5852);
and U6132 (N_6132,N_5146,N_5957);
and U6133 (N_6133,N_5536,N_5258);
or U6134 (N_6134,N_5102,N_5487);
and U6135 (N_6135,N_5474,N_5621);
and U6136 (N_6136,N_5354,N_5912);
and U6137 (N_6137,N_5497,N_5887);
or U6138 (N_6138,N_5375,N_5774);
xnor U6139 (N_6139,N_5257,N_5277);
or U6140 (N_6140,N_5558,N_5828);
nor U6141 (N_6141,N_5007,N_5522);
or U6142 (N_6142,N_5150,N_5596);
and U6143 (N_6143,N_5360,N_5057);
nand U6144 (N_6144,N_5216,N_5717);
nand U6145 (N_6145,N_5514,N_5875);
nor U6146 (N_6146,N_5406,N_5181);
and U6147 (N_6147,N_5771,N_5836);
nor U6148 (N_6148,N_5851,N_5255);
or U6149 (N_6149,N_5837,N_5714);
nand U6150 (N_6150,N_5378,N_5111);
and U6151 (N_6151,N_5623,N_5696);
nand U6152 (N_6152,N_5563,N_5248);
and U6153 (N_6153,N_5928,N_5808);
nor U6154 (N_6154,N_5100,N_5888);
nor U6155 (N_6155,N_5530,N_5720);
or U6156 (N_6156,N_5801,N_5583);
and U6157 (N_6157,N_5632,N_5655);
or U6158 (N_6158,N_5945,N_5654);
nor U6159 (N_6159,N_5624,N_5492);
nand U6160 (N_6160,N_5407,N_5256);
nand U6161 (N_6161,N_5936,N_5643);
nor U6162 (N_6162,N_5062,N_5730);
nand U6163 (N_6163,N_5835,N_5442);
nand U6164 (N_6164,N_5018,N_5806);
xor U6165 (N_6165,N_5664,N_5822);
and U6166 (N_6166,N_5495,N_5657);
and U6167 (N_6167,N_5840,N_5590);
nand U6168 (N_6168,N_5477,N_5816);
nor U6169 (N_6169,N_5869,N_5447);
nand U6170 (N_6170,N_5196,N_5626);
or U6171 (N_6171,N_5824,N_5861);
and U6172 (N_6172,N_5511,N_5954);
nor U6173 (N_6173,N_5983,N_5092);
or U6174 (N_6174,N_5883,N_5362);
nand U6175 (N_6175,N_5803,N_5819);
or U6176 (N_6176,N_5358,N_5036);
nor U6177 (N_6177,N_5060,N_5812);
nand U6178 (N_6178,N_5204,N_5907);
nor U6179 (N_6179,N_5651,N_5391);
or U6180 (N_6180,N_5645,N_5543);
nor U6181 (N_6181,N_5178,N_5943);
and U6182 (N_6182,N_5113,N_5569);
and U6183 (N_6183,N_5908,N_5619);
and U6184 (N_6184,N_5041,N_5946);
or U6185 (N_6185,N_5212,N_5344);
nor U6186 (N_6186,N_5229,N_5489);
and U6187 (N_6187,N_5372,N_5073);
xnor U6188 (N_6188,N_5749,N_5666);
nor U6189 (N_6189,N_5811,N_5093);
or U6190 (N_6190,N_5233,N_5878);
and U6191 (N_6191,N_5989,N_5524);
nand U6192 (N_6192,N_5261,N_5750);
and U6193 (N_6193,N_5135,N_5827);
or U6194 (N_6194,N_5959,N_5540);
or U6195 (N_6195,N_5502,N_5929);
nor U6196 (N_6196,N_5046,N_5708);
nor U6197 (N_6197,N_5334,N_5760);
nor U6198 (N_6198,N_5831,N_5211);
and U6199 (N_6199,N_5885,N_5555);
and U6200 (N_6200,N_5209,N_5249);
nor U6201 (N_6201,N_5853,N_5491);
nor U6202 (N_6202,N_5333,N_5357);
nor U6203 (N_6203,N_5898,N_5176);
or U6204 (N_6204,N_5763,N_5189);
or U6205 (N_6205,N_5137,N_5201);
nor U6206 (N_6206,N_5419,N_5425);
or U6207 (N_6207,N_5743,N_5287);
nor U6208 (N_6208,N_5380,N_5222);
nor U6209 (N_6209,N_5077,N_5095);
nor U6210 (N_6210,N_5247,N_5753);
and U6211 (N_6211,N_5218,N_5859);
nor U6212 (N_6212,N_5318,N_5709);
nand U6213 (N_6213,N_5445,N_5584);
xor U6214 (N_6214,N_5600,N_5453);
and U6215 (N_6215,N_5061,N_5977);
or U6216 (N_6216,N_5958,N_5877);
nor U6217 (N_6217,N_5339,N_5316);
nor U6218 (N_6218,N_5576,N_5139);
and U6219 (N_6219,N_5025,N_5459);
xnor U6220 (N_6220,N_5421,N_5019);
and U6221 (N_6221,N_5024,N_5710);
and U6222 (N_6222,N_5106,N_5002);
nand U6223 (N_6223,N_5985,N_5608);
xor U6224 (N_6224,N_5589,N_5027);
and U6225 (N_6225,N_5581,N_5501);
or U6226 (N_6226,N_5356,N_5694);
and U6227 (N_6227,N_5633,N_5776);
xor U6228 (N_6228,N_5037,N_5577);
xor U6229 (N_6229,N_5706,N_5909);
or U6230 (N_6230,N_5200,N_5064);
nand U6231 (N_6231,N_5158,N_5049);
nor U6232 (N_6232,N_5148,N_5855);
xnor U6233 (N_6233,N_5953,N_5392);
nand U6234 (N_6234,N_5383,N_5715);
or U6235 (N_6235,N_5496,N_5005);
or U6236 (N_6236,N_5097,N_5133);
nor U6237 (N_6237,N_5580,N_5310);
and U6238 (N_6238,N_5288,N_5285);
and U6239 (N_6239,N_5799,N_5988);
nor U6240 (N_6240,N_5444,N_5021);
or U6241 (N_6241,N_5480,N_5230);
and U6242 (N_6242,N_5127,N_5768);
nand U6243 (N_6243,N_5052,N_5213);
and U6244 (N_6244,N_5677,N_5274);
or U6245 (N_6245,N_5126,N_5872);
nor U6246 (N_6246,N_5678,N_5069);
nand U6247 (N_6247,N_5854,N_5738);
nand U6248 (N_6248,N_5350,N_5044);
or U6249 (N_6249,N_5610,N_5780);
nand U6250 (N_6250,N_5616,N_5396);
and U6251 (N_6251,N_5703,N_5353);
nor U6252 (N_6252,N_5366,N_5518);
and U6253 (N_6253,N_5858,N_5125);
or U6254 (N_6254,N_5000,N_5132);
nor U6255 (N_6255,N_5388,N_5642);
or U6256 (N_6256,N_5072,N_5939);
nor U6257 (N_6257,N_5153,N_5571);
nor U6258 (N_6258,N_5637,N_5498);
and U6259 (N_6259,N_5702,N_5254);
nor U6260 (N_6260,N_5427,N_5108);
or U6261 (N_6261,N_5386,N_5413);
nor U6262 (N_6262,N_5873,N_5120);
and U6263 (N_6263,N_5162,N_5652);
nand U6264 (N_6264,N_5030,N_5217);
nor U6265 (N_6265,N_5849,N_5207);
and U6266 (N_6266,N_5237,N_5469);
or U6267 (N_6267,N_5922,N_5269);
nor U6268 (N_6268,N_5486,N_5440);
or U6269 (N_6269,N_5422,N_5932);
and U6270 (N_6270,N_5451,N_5475);
nor U6271 (N_6271,N_5154,N_5865);
nand U6272 (N_6272,N_5992,N_5896);
or U6273 (N_6273,N_5857,N_5974);
or U6274 (N_6274,N_5290,N_5964);
or U6275 (N_6275,N_5270,N_5634);
or U6276 (N_6276,N_5682,N_5319);
and U6277 (N_6277,N_5758,N_5175);
nor U6278 (N_6278,N_5088,N_5982);
and U6279 (N_6279,N_5751,N_5550);
or U6280 (N_6280,N_5345,N_5906);
nor U6281 (N_6281,N_5083,N_5473);
nor U6282 (N_6282,N_5681,N_5879);
and U6283 (N_6283,N_5091,N_5786);
or U6284 (N_6284,N_5081,N_5040);
nor U6285 (N_6285,N_5880,N_5109);
nand U6286 (N_6286,N_5202,N_5377);
nand U6287 (N_6287,N_5940,N_5006);
or U6288 (N_6288,N_5183,N_5337);
nand U6289 (N_6289,N_5892,N_5561);
or U6290 (N_6290,N_5508,N_5698);
nand U6291 (N_6291,N_5295,N_5578);
nor U6292 (N_6292,N_5722,N_5805);
nor U6293 (N_6293,N_5695,N_5143);
nor U6294 (N_6294,N_5465,N_5156);
nand U6295 (N_6295,N_5048,N_5593);
nand U6296 (N_6296,N_5004,N_5742);
or U6297 (N_6297,N_5449,N_5972);
nor U6298 (N_6298,N_5364,N_5160);
or U6299 (N_6299,N_5348,N_5700);
and U6300 (N_6300,N_5381,N_5503);
or U6301 (N_6301,N_5732,N_5661);
nand U6302 (N_6302,N_5673,N_5779);
and U6303 (N_6303,N_5745,N_5531);
and U6304 (N_6304,N_5739,N_5215);
nand U6305 (N_6305,N_5656,N_5647);
and U6306 (N_6306,N_5785,N_5860);
nor U6307 (N_6307,N_5833,N_5482);
nand U6308 (N_6308,N_5727,N_5573);
nand U6309 (N_6309,N_5028,N_5533);
and U6310 (N_6310,N_5956,N_5323);
nor U6311 (N_6311,N_5499,N_5379);
and U6312 (N_6312,N_5300,N_5415);
nor U6313 (N_6313,N_5164,N_5191);
or U6314 (N_6314,N_5537,N_5405);
and U6315 (N_6315,N_5901,N_5740);
and U6316 (N_6316,N_5980,N_5547);
nand U6317 (N_6317,N_5520,N_5149);
nor U6318 (N_6318,N_5979,N_5613);
nand U6319 (N_6319,N_5797,N_5338);
nor U6320 (N_6320,N_5446,N_5330);
xnor U6321 (N_6321,N_5716,N_5238);
nand U6322 (N_6322,N_5844,N_5870);
or U6323 (N_6323,N_5790,N_5663);
or U6324 (N_6324,N_5184,N_5494);
and U6325 (N_6325,N_5235,N_5975);
nand U6326 (N_6326,N_5683,N_5687);
nor U6327 (N_6327,N_5881,N_5529);
or U6328 (N_6328,N_5539,N_5053);
or U6329 (N_6329,N_5707,N_5915);
nor U6330 (N_6330,N_5124,N_5927);
or U6331 (N_6331,N_5899,N_5468);
nor U6332 (N_6332,N_5549,N_5332);
or U6333 (N_6333,N_5169,N_5741);
nand U6334 (N_6334,N_5597,N_5117);
or U6335 (N_6335,N_5479,N_5704);
or U6336 (N_6336,N_5644,N_5769);
nand U6337 (N_6337,N_5462,N_5484);
and U6338 (N_6338,N_5754,N_5757);
and U6339 (N_6339,N_5541,N_5390);
nor U6340 (N_6340,N_5078,N_5587);
or U6341 (N_6341,N_5919,N_5402);
nor U6342 (N_6342,N_5432,N_5241);
nand U6343 (N_6343,N_5999,N_5214);
nor U6344 (N_6344,N_5074,N_5519);
and U6345 (N_6345,N_5782,N_5483);
and U6346 (N_6346,N_5510,N_5418);
or U6347 (N_6347,N_5560,N_5309);
xor U6348 (N_6348,N_5931,N_5599);
nand U6349 (N_6349,N_5417,N_5762);
and U6350 (N_6350,N_5841,N_5609);
nand U6351 (N_6351,N_5308,N_5096);
nor U6352 (N_6352,N_5084,N_5147);
nand U6353 (N_6353,N_5012,N_5617);
nand U6354 (N_6354,N_5098,N_5094);
or U6355 (N_6355,N_5234,N_5056);
nor U6356 (N_6356,N_5910,N_5349);
nor U6357 (N_6357,N_5347,N_5242);
and U6358 (N_6358,N_5368,N_5930);
xor U6359 (N_6359,N_5960,N_5389);
or U6360 (N_6360,N_5141,N_5594);
nor U6361 (N_6361,N_5262,N_5253);
or U6362 (N_6362,N_5227,N_5231);
nor U6363 (N_6363,N_5614,N_5470);
nor U6364 (N_6364,N_5622,N_5726);
nand U6365 (N_6365,N_5705,N_5796);
and U6366 (N_6366,N_5568,N_5688);
nand U6367 (N_6367,N_5010,N_5570);
and U6368 (N_6368,N_5725,N_5452);
and U6369 (N_6369,N_5352,N_5284);
nor U6370 (N_6370,N_5485,N_5429);
nor U6371 (N_6371,N_5420,N_5545);
nand U6372 (N_6372,N_5401,N_5304);
nand U6373 (N_6373,N_5047,N_5219);
or U6374 (N_6374,N_5752,N_5969);
nand U6375 (N_6375,N_5966,N_5640);
and U6376 (N_6376,N_5013,N_5171);
nand U6377 (N_6377,N_5326,N_5203);
or U6378 (N_6378,N_5301,N_5431);
and U6379 (N_6379,N_5114,N_5998);
and U6380 (N_6380,N_5272,N_5990);
nor U6381 (N_6381,N_5434,N_5260);
nor U6382 (N_6382,N_5665,N_5291);
nand U6383 (N_6383,N_5244,N_5426);
nor U6384 (N_6384,N_5871,N_5173);
nand U6385 (N_6385,N_5993,N_5065);
or U6386 (N_6386,N_5658,N_5195);
and U6387 (N_6387,N_5414,N_5433);
and U6388 (N_6388,N_5672,N_5315);
or U6389 (N_6389,N_5085,N_5245);
or U6390 (N_6390,N_5029,N_5924);
nand U6391 (N_6391,N_5500,N_5601);
nand U6392 (N_6392,N_5058,N_5186);
nor U6393 (N_6393,N_5001,N_5856);
nand U6394 (N_6394,N_5145,N_5464);
xor U6395 (N_6395,N_5138,N_5787);
nor U6396 (N_6396,N_5220,N_5268);
or U6397 (N_6397,N_5224,N_5008);
nor U6398 (N_6398,N_5886,N_5976);
or U6399 (N_6399,N_5978,N_5986);
or U6400 (N_6400,N_5437,N_5112);
nand U6401 (N_6401,N_5239,N_5934);
and U6402 (N_6402,N_5014,N_5243);
nand U6403 (N_6403,N_5424,N_5306);
or U6404 (N_6404,N_5341,N_5283);
and U6405 (N_6405,N_5807,N_5693);
nand U6406 (N_6406,N_5398,N_5327);
or U6407 (N_6407,N_5267,N_5369);
or U6408 (N_6408,N_5534,N_5443);
nor U6409 (N_6409,N_5628,N_5968);
nand U6410 (N_6410,N_5546,N_5848);
nand U6411 (N_6411,N_5336,N_5165);
or U6412 (N_6412,N_5574,N_5867);
or U6413 (N_6413,N_5952,N_5428);
nand U6414 (N_6414,N_5938,N_5890);
or U6415 (N_6415,N_5897,N_5179);
nand U6416 (N_6416,N_5916,N_5800);
nor U6417 (N_6417,N_5140,N_5403);
and U6418 (N_6418,N_5793,N_5766);
nand U6419 (N_6419,N_5585,N_5055);
or U6420 (N_6420,N_5962,N_5441);
and U6421 (N_6421,N_5082,N_5772);
and U6422 (N_6422,N_5026,N_5263);
nand U6423 (N_6423,N_5971,N_5544);
or U6424 (N_6424,N_5668,N_5933);
and U6425 (N_6425,N_5813,N_5340);
nor U6426 (N_6426,N_5842,N_5659);
and U6427 (N_6427,N_5984,N_5320);
and U6428 (N_6428,N_5575,N_5210);
and U6429 (N_6429,N_5676,N_5963);
and U6430 (N_6430,N_5973,N_5784);
nand U6431 (N_6431,N_5411,N_5023);
or U6432 (N_6432,N_5792,N_5967);
nand U6433 (N_6433,N_5182,N_5675);
nor U6434 (N_6434,N_5050,N_5789);
and U6435 (N_6435,N_5662,N_5159);
nor U6436 (N_6436,N_5671,N_5163);
nor U6437 (N_6437,N_5996,N_5279);
or U6438 (N_6438,N_5893,N_5775);
and U6439 (N_6439,N_5950,N_5551);
nand U6440 (N_6440,N_5022,N_5691);
or U6441 (N_6441,N_5650,N_5612);
or U6442 (N_6442,N_5408,N_5251);
nor U6443 (N_6443,N_5542,N_5509);
nand U6444 (N_6444,N_5731,N_5325);
and U6445 (N_6445,N_5951,N_5556);
or U6446 (N_6446,N_5627,N_5777);
nor U6447 (N_6447,N_5564,N_5031);
nor U6448 (N_6448,N_5151,N_5699);
and U6449 (N_6449,N_5832,N_5804);
nor U6450 (N_6450,N_5066,N_5809);
and U6451 (N_6451,N_5917,N_5087);
or U6452 (N_6452,N_5275,N_5712);
nand U6453 (N_6453,N_5250,N_5136);
nor U6454 (N_6454,N_5177,N_5736);
nor U6455 (N_6455,N_5729,N_5404);
nor U6456 (N_6456,N_5506,N_5914);
or U6457 (N_6457,N_5747,N_5653);
nor U6458 (N_6458,N_5846,N_5620);
nor U6459 (N_6459,N_5076,N_5629);
and U6460 (N_6460,N_5761,N_5997);
nor U6461 (N_6461,N_5773,N_5104);
or U6462 (N_6462,N_5105,N_5329);
nand U6463 (N_6463,N_5783,N_5552);
nand U6464 (N_6464,N_5371,N_5467);
nand U6465 (N_6465,N_5904,N_5307);
and U6466 (N_6466,N_5925,N_5595);
nand U6467 (N_6467,N_5264,N_5701);
or U6468 (N_6468,N_5192,N_5051);
nand U6469 (N_6469,N_5039,N_5455);
nor U6470 (N_6470,N_5713,N_5810);
and U6471 (N_6471,N_5602,N_5193);
and U6472 (N_6472,N_5365,N_5099);
nor U6473 (N_6473,N_5478,N_5463);
and U6474 (N_6474,N_5829,N_5152);
nand U6475 (N_6475,N_5003,N_5718);
or U6476 (N_6476,N_5273,N_5313);
or U6477 (N_6477,N_5075,N_5172);
nand U6478 (N_6478,N_5525,N_5759);
nand U6479 (N_6479,N_5660,N_5923);
and U6480 (N_6480,N_5965,N_5876);
and U6481 (N_6481,N_5823,N_5527);
and U6482 (N_6482,N_5493,N_5937);
or U6483 (N_6483,N_5894,N_5866);
or U6484 (N_6484,N_5121,N_5363);
or U6485 (N_6485,N_5020,N_5071);
nor U6486 (N_6486,N_5367,N_5826);
and U6487 (N_6487,N_5523,N_5843);
and U6488 (N_6488,N_5303,N_5305);
xor U6489 (N_6489,N_5197,N_5232);
and U6490 (N_6490,N_5035,N_5103);
nand U6491 (N_6491,N_5680,N_5830);
nand U6492 (N_6492,N_5070,N_5505);
and U6493 (N_6493,N_5981,N_5911);
nor U6494 (N_6494,N_5606,N_5559);
or U6495 (N_6495,N_5630,N_5187);
and U6496 (N_6496,N_5130,N_5461);
and U6497 (N_6497,N_5941,N_5080);
nor U6498 (N_6498,N_5548,N_5987);
xor U6499 (N_6499,N_5410,N_5689);
nor U6500 (N_6500,N_5362,N_5175);
and U6501 (N_6501,N_5792,N_5899);
or U6502 (N_6502,N_5110,N_5559);
and U6503 (N_6503,N_5225,N_5713);
and U6504 (N_6504,N_5519,N_5870);
and U6505 (N_6505,N_5024,N_5291);
nor U6506 (N_6506,N_5681,N_5972);
or U6507 (N_6507,N_5417,N_5114);
and U6508 (N_6508,N_5408,N_5311);
nor U6509 (N_6509,N_5648,N_5499);
or U6510 (N_6510,N_5780,N_5981);
and U6511 (N_6511,N_5708,N_5562);
nand U6512 (N_6512,N_5762,N_5744);
nand U6513 (N_6513,N_5524,N_5425);
nor U6514 (N_6514,N_5288,N_5458);
nand U6515 (N_6515,N_5767,N_5381);
nand U6516 (N_6516,N_5068,N_5063);
nand U6517 (N_6517,N_5523,N_5897);
nor U6518 (N_6518,N_5444,N_5806);
nor U6519 (N_6519,N_5675,N_5890);
nor U6520 (N_6520,N_5616,N_5490);
nor U6521 (N_6521,N_5608,N_5136);
nand U6522 (N_6522,N_5060,N_5185);
and U6523 (N_6523,N_5832,N_5300);
nand U6524 (N_6524,N_5407,N_5801);
nor U6525 (N_6525,N_5224,N_5693);
nand U6526 (N_6526,N_5022,N_5925);
and U6527 (N_6527,N_5741,N_5349);
and U6528 (N_6528,N_5174,N_5807);
nor U6529 (N_6529,N_5168,N_5707);
or U6530 (N_6530,N_5229,N_5069);
nor U6531 (N_6531,N_5331,N_5465);
nand U6532 (N_6532,N_5105,N_5410);
and U6533 (N_6533,N_5793,N_5404);
or U6534 (N_6534,N_5778,N_5320);
nand U6535 (N_6535,N_5704,N_5674);
nand U6536 (N_6536,N_5737,N_5337);
or U6537 (N_6537,N_5204,N_5682);
nand U6538 (N_6538,N_5606,N_5414);
or U6539 (N_6539,N_5643,N_5802);
nor U6540 (N_6540,N_5450,N_5457);
or U6541 (N_6541,N_5784,N_5698);
nand U6542 (N_6542,N_5975,N_5950);
nor U6543 (N_6543,N_5073,N_5381);
or U6544 (N_6544,N_5119,N_5049);
nand U6545 (N_6545,N_5026,N_5315);
and U6546 (N_6546,N_5651,N_5993);
nand U6547 (N_6547,N_5808,N_5525);
nor U6548 (N_6548,N_5217,N_5705);
nor U6549 (N_6549,N_5318,N_5825);
or U6550 (N_6550,N_5597,N_5748);
or U6551 (N_6551,N_5344,N_5644);
nor U6552 (N_6552,N_5113,N_5509);
and U6553 (N_6553,N_5060,N_5221);
and U6554 (N_6554,N_5286,N_5291);
or U6555 (N_6555,N_5607,N_5667);
and U6556 (N_6556,N_5672,N_5868);
nand U6557 (N_6557,N_5659,N_5158);
nor U6558 (N_6558,N_5749,N_5475);
nand U6559 (N_6559,N_5368,N_5860);
nand U6560 (N_6560,N_5535,N_5568);
and U6561 (N_6561,N_5660,N_5744);
or U6562 (N_6562,N_5409,N_5621);
nand U6563 (N_6563,N_5634,N_5220);
nand U6564 (N_6564,N_5125,N_5228);
and U6565 (N_6565,N_5633,N_5758);
or U6566 (N_6566,N_5755,N_5066);
and U6567 (N_6567,N_5592,N_5581);
nand U6568 (N_6568,N_5434,N_5233);
and U6569 (N_6569,N_5046,N_5023);
or U6570 (N_6570,N_5222,N_5315);
and U6571 (N_6571,N_5898,N_5800);
or U6572 (N_6572,N_5116,N_5709);
nand U6573 (N_6573,N_5117,N_5796);
or U6574 (N_6574,N_5222,N_5620);
nand U6575 (N_6575,N_5140,N_5860);
and U6576 (N_6576,N_5500,N_5025);
or U6577 (N_6577,N_5134,N_5941);
nor U6578 (N_6578,N_5191,N_5812);
or U6579 (N_6579,N_5550,N_5730);
nor U6580 (N_6580,N_5771,N_5774);
nor U6581 (N_6581,N_5932,N_5452);
nor U6582 (N_6582,N_5430,N_5395);
nand U6583 (N_6583,N_5487,N_5353);
nand U6584 (N_6584,N_5582,N_5511);
nand U6585 (N_6585,N_5210,N_5679);
nor U6586 (N_6586,N_5154,N_5486);
nor U6587 (N_6587,N_5092,N_5941);
or U6588 (N_6588,N_5324,N_5803);
and U6589 (N_6589,N_5384,N_5398);
and U6590 (N_6590,N_5403,N_5982);
nand U6591 (N_6591,N_5254,N_5429);
nor U6592 (N_6592,N_5161,N_5538);
and U6593 (N_6593,N_5041,N_5222);
nor U6594 (N_6594,N_5841,N_5631);
or U6595 (N_6595,N_5994,N_5307);
and U6596 (N_6596,N_5123,N_5551);
and U6597 (N_6597,N_5713,N_5526);
nand U6598 (N_6598,N_5324,N_5047);
and U6599 (N_6599,N_5663,N_5935);
and U6600 (N_6600,N_5973,N_5621);
nand U6601 (N_6601,N_5268,N_5890);
nor U6602 (N_6602,N_5744,N_5152);
nor U6603 (N_6603,N_5337,N_5005);
nor U6604 (N_6604,N_5408,N_5874);
or U6605 (N_6605,N_5706,N_5170);
or U6606 (N_6606,N_5142,N_5859);
nand U6607 (N_6607,N_5340,N_5539);
and U6608 (N_6608,N_5003,N_5023);
or U6609 (N_6609,N_5418,N_5099);
nand U6610 (N_6610,N_5579,N_5518);
nor U6611 (N_6611,N_5845,N_5423);
nand U6612 (N_6612,N_5234,N_5544);
nand U6613 (N_6613,N_5112,N_5998);
and U6614 (N_6614,N_5268,N_5025);
nand U6615 (N_6615,N_5492,N_5082);
nor U6616 (N_6616,N_5358,N_5085);
or U6617 (N_6617,N_5089,N_5588);
and U6618 (N_6618,N_5730,N_5100);
nor U6619 (N_6619,N_5374,N_5031);
and U6620 (N_6620,N_5855,N_5415);
nor U6621 (N_6621,N_5859,N_5354);
or U6622 (N_6622,N_5618,N_5989);
and U6623 (N_6623,N_5620,N_5515);
and U6624 (N_6624,N_5541,N_5930);
or U6625 (N_6625,N_5508,N_5874);
and U6626 (N_6626,N_5184,N_5062);
nand U6627 (N_6627,N_5421,N_5339);
or U6628 (N_6628,N_5353,N_5812);
nor U6629 (N_6629,N_5322,N_5463);
nand U6630 (N_6630,N_5153,N_5207);
nor U6631 (N_6631,N_5759,N_5425);
nor U6632 (N_6632,N_5938,N_5548);
nand U6633 (N_6633,N_5180,N_5862);
or U6634 (N_6634,N_5684,N_5316);
nor U6635 (N_6635,N_5603,N_5276);
nand U6636 (N_6636,N_5292,N_5288);
or U6637 (N_6637,N_5083,N_5690);
or U6638 (N_6638,N_5433,N_5941);
and U6639 (N_6639,N_5636,N_5893);
nor U6640 (N_6640,N_5807,N_5753);
or U6641 (N_6641,N_5789,N_5341);
or U6642 (N_6642,N_5783,N_5965);
nand U6643 (N_6643,N_5294,N_5743);
nor U6644 (N_6644,N_5132,N_5158);
nand U6645 (N_6645,N_5836,N_5848);
or U6646 (N_6646,N_5701,N_5644);
and U6647 (N_6647,N_5613,N_5097);
nand U6648 (N_6648,N_5452,N_5443);
and U6649 (N_6649,N_5244,N_5566);
or U6650 (N_6650,N_5478,N_5169);
nand U6651 (N_6651,N_5068,N_5757);
or U6652 (N_6652,N_5098,N_5049);
nand U6653 (N_6653,N_5756,N_5262);
nor U6654 (N_6654,N_5805,N_5091);
nand U6655 (N_6655,N_5404,N_5630);
nor U6656 (N_6656,N_5118,N_5557);
or U6657 (N_6657,N_5769,N_5392);
nor U6658 (N_6658,N_5214,N_5796);
nor U6659 (N_6659,N_5059,N_5597);
or U6660 (N_6660,N_5907,N_5759);
and U6661 (N_6661,N_5530,N_5737);
nand U6662 (N_6662,N_5350,N_5420);
or U6663 (N_6663,N_5153,N_5568);
nor U6664 (N_6664,N_5013,N_5660);
nand U6665 (N_6665,N_5601,N_5176);
nor U6666 (N_6666,N_5706,N_5451);
nand U6667 (N_6667,N_5035,N_5260);
or U6668 (N_6668,N_5037,N_5435);
and U6669 (N_6669,N_5456,N_5592);
nor U6670 (N_6670,N_5758,N_5293);
nor U6671 (N_6671,N_5654,N_5800);
and U6672 (N_6672,N_5459,N_5425);
and U6673 (N_6673,N_5865,N_5744);
nor U6674 (N_6674,N_5921,N_5401);
and U6675 (N_6675,N_5617,N_5105);
and U6676 (N_6676,N_5888,N_5098);
or U6677 (N_6677,N_5758,N_5251);
nor U6678 (N_6678,N_5107,N_5093);
nor U6679 (N_6679,N_5257,N_5814);
nand U6680 (N_6680,N_5870,N_5557);
or U6681 (N_6681,N_5039,N_5149);
and U6682 (N_6682,N_5852,N_5163);
nor U6683 (N_6683,N_5859,N_5469);
nor U6684 (N_6684,N_5334,N_5014);
or U6685 (N_6685,N_5200,N_5264);
nand U6686 (N_6686,N_5102,N_5983);
or U6687 (N_6687,N_5629,N_5590);
or U6688 (N_6688,N_5727,N_5940);
or U6689 (N_6689,N_5502,N_5461);
or U6690 (N_6690,N_5253,N_5141);
or U6691 (N_6691,N_5446,N_5315);
and U6692 (N_6692,N_5006,N_5185);
nand U6693 (N_6693,N_5540,N_5775);
nand U6694 (N_6694,N_5023,N_5854);
nand U6695 (N_6695,N_5750,N_5427);
and U6696 (N_6696,N_5924,N_5713);
and U6697 (N_6697,N_5612,N_5405);
and U6698 (N_6698,N_5267,N_5758);
or U6699 (N_6699,N_5476,N_5769);
nand U6700 (N_6700,N_5863,N_5948);
nand U6701 (N_6701,N_5984,N_5913);
or U6702 (N_6702,N_5270,N_5679);
or U6703 (N_6703,N_5787,N_5285);
nand U6704 (N_6704,N_5660,N_5123);
nor U6705 (N_6705,N_5533,N_5873);
and U6706 (N_6706,N_5259,N_5864);
or U6707 (N_6707,N_5153,N_5609);
nor U6708 (N_6708,N_5612,N_5126);
or U6709 (N_6709,N_5596,N_5945);
and U6710 (N_6710,N_5053,N_5889);
and U6711 (N_6711,N_5331,N_5243);
and U6712 (N_6712,N_5907,N_5140);
or U6713 (N_6713,N_5348,N_5769);
or U6714 (N_6714,N_5391,N_5619);
and U6715 (N_6715,N_5055,N_5887);
nand U6716 (N_6716,N_5173,N_5526);
nand U6717 (N_6717,N_5841,N_5929);
nand U6718 (N_6718,N_5228,N_5237);
nor U6719 (N_6719,N_5711,N_5981);
or U6720 (N_6720,N_5061,N_5014);
nand U6721 (N_6721,N_5657,N_5069);
nand U6722 (N_6722,N_5170,N_5324);
nand U6723 (N_6723,N_5073,N_5144);
nand U6724 (N_6724,N_5764,N_5722);
nand U6725 (N_6725,N_5456,N_5007);
and U6726 (N_6726,N_5737,N_5087);
or U6727 (N_6727,N_5790,N_5087);
or U6728 (N_6728,N_5498,N_5785);
or U6729 (N_6729,N_5495,N_5401);
and U6730 (N_6730,N_5865,N_5778);
nand U6731 (N_6731,N_5123,N_5638);
or U6732 (N_6732,N_5841,N_5311);
nand U6733 (N_6733,N_5235,N_5052);
and U6734 (N_6734,N_5113,N_5114);
nand U6735 (N_6735,N_5461,N_5740);
or U6736 (N_6736,N_5065,N_5410);
or U6737 (N_6737,N_5027,N_5612);
or U6738 (N_6738,N_5858,N_5367);
nor U6739 (N_6739,N_5617,N_5992);
and U6740 (N_6740,N_5279,N_5488);
or U6741 (N_6741,N_5579,N_5985);
nor U6742 (N_6742,N_5679,N_5392);
and U6743 (N_6743,N_5690,N_5912);
nand U6744 (N_6744,N_5414,N_5480);
or U6745 (N_6745,N_5934,N_5869);
and U6746 (N_6746,N_5381,N_5020);
nor U6747 (N_6747,N_5960,N_5278);
nor U6748 (N_6748,N_5727,N_5090);
or U6749 (N_6749,N_5188,N_5856);
or U6750 (N_6750,N_5039,N_5817);
nand U6751 (N_6751,N_5442,N_5431);
and U6752 (N_6752,N_5794,N_5309);
nand U6753 (N_6753,N_5827,N_5209);
nor U6754 (N_6754,N_5008,N_5402);
nor U6755 (N_6755,N_5555,N_5264);
nor U6756 (N_6756,N_5690,N_5669);
and U6757 (N_6757,N_5727,N_5517);
and U6758 (N_6758,N_5053,N_5095);
and U6759 (N_6759,N_5461,N_5463);
nor U6760 (N_6760,N_5442,N_5793);
or U6761 (N_6761,N_5607,N_5238);
nor U6762 (N_6762,N_5179,N_5239);
or U6763 (N_6763,N_5498,N_5177);
nor U6764 (N_6764,N_5395,N_5003);
and U6765 (N_6765,N_5309,N_5040);
and U6766 (N_6766,N_5798,N_5811);
nand U6767 (N_6767,N_5237,N_5191);
nand U6768 (N_6768,N_5841,N_5026);
or U6769 (N_6769,N_5289,N_5040);
nand U6770 (N_6770,N_5989,N_5140);
or U6771 (N_6771,N_5190,N_5572);
nor U6772 (N_6772,N_5706,N_5079);
nand U6773 (N_6773,N_5328,N_5240);
or U6774 (N_6774,N_5366,N_5582);
or U6775 (N_6775,N_5094,N_5137);
nand U6776 (N_6776,N_5744,N_5259);
nand U6777 (N_6777,N_5150,N_5592);
nand U6778 (N_6778,N_5189,N_5176);
or U6779 (N_6779,N_5150,N_5221);
nor U6780 (N_6780,N_5456,N_5303);
nor U6781 (N_6781,N_5290,N_5124);
or U6782 (N_6782,N_5465,N_5066);
nor U6783 (N_6783,N_5323,N_5360);
and U6784 (N_6784,N_5245,N_5908);
nand U6785 (N_6785,N_5703,N_5649);
or U6786 (N_6786,N_5707,N_5011);
nor U6787 (N_6787,N_5776,N_5241);
nor U6788 (N_6788,N_5157,N_5034);
or U6789 (N_6789,N_5736,N_5022);
nor U6790 (N_6790,N_5659,N_5728);
nand U6791 (N_6791,N_5675,N_5960);
nor U6792 (N_6792,N_5799,N_5208);
nor U6793 (N_6793,N_5874,N_5212);
or U6794 (N_6794,N_5091,N_5249);
nor U6795 (N_6795,N_5216,N_5556);
or U6796 (N_6796,N_5641,N_5591);
nor U6797 (N_6797,N_5494,N_5645);
and U6798 (N_6798,N_5531,N_5869);
nand U6799 (N_6799,N_5481,N_5505);
or U6800 (N_6800,N_5684,N_5987);
nand U6801 (N_6801,N_5293,N_5911);
nand U6802 (N_6802,N_5107,N_5025);
nand U6803 (N_6803,N_5700,N_5400);
and U6804 (N_6804,N_5112,N_5207);
or U6805 (N_6805,N_5568,N_5469);
xor U6806 (N_6806,N_5938,N_5520);
nand U6807 (N_6807,N_5105,N_5754);
nor U6808 (N_6808,N_5725,N_5345);
nand U6809 (N_6809,N_5869,N_5234);
nand U6810 (N_6810,N_5954,N_5661);
and U6811 (N_6811,N_5399,N_5266);
or U6812 (N_6812,N_5904,N_5343);
and U6813 (N_6813,N_5961,N_5559);
and U6814 (N_6814,N_5053,N_5477);
nor U6815 (N_6815,N_5012,N_5359);
nor U6816 (N_6816,N_5738,N_5196);
and U6817 (N_6817,N_5890,N_5407);
and U6818 (N_6818,N_5521,N_5671);
and U6819 (N_6819,N_5025,N_5017);
or U6820 (N_6820,N_5866,N_5898);
and U6821 (N_6821,N_5460,N_5109);
and U6822 (N_6822,N_5278,N_5348);
and U6823 (N_6823,N_5978,N_5366);
or U6824 (N_6824,N_5742,N_5487);
and U6825 (N_6825,N_5146,N_5837);
and U6826 (N_6826,N_5555,N_5810);
nand U6827 (N_6827,N_5270,N_5384);
nand U6828 (N_6828,N_5232,N_5219);
nor U6829 (N_6829,N_5897,N_5178);
nand U6830 (N_6830,N_5911,N_5298);
nand U6831 (N_6831,N_5016,N_5023);
or U6832 (N_6832,N_5341,N_5966);
nand U6833 (N_6833,N_5413,N_5618);
or U6834 (N_6834,N_5366,N_5894);
nor U6835 (N_6835,N_5216,N_5494);
or U6836 (N_6836,N_5384,N_5292);
or U6837 (N_6837,N_5268,N_5206);
or U6838 (N_6838,N_5162,N_5517);
or U6839 (N_6839,N_5701,N_5346);
nand U6840 (N_6840,N_5717,N_5925);
or U6841 (N_6841,N_5478,N_5409);
or U6842 (N_6842,N_5145,N_5356);
nor U6843 (N_6843,N_5221,N_5425);
or U6844 (N_6844,N_5956,N_5797);
and U6845 (N_6845,N_5165,N_5108);
or U6846 (N_6846,N_5727,N_5166);
and U6847 (N_6847,N_5416,N_5550);
or U6848 (N_6848,N_5276,N_5962);
and U6849 (N_6849,N_5524,N_5786);
and U6850 (N_6850,N_5238,N_5299);
nand U6851 (N_6851,N_5539,N_5159);
xnor U6852 (N_6852,N_5363,N_5084);
nand U6853 (N_6853,N_5509,N_5440);
nor U6854 (N_6854,N_5860,N_5950);
or U6855 (N_6855,N_5329,N_5977);
nor U6856 (N_6856,N_5692,N_5502);
or U6857 (N_6857,N_5603,N_5614);
and U6858 (N_6858,N_5061,N_5412);
or U6859 (N_6859,N_5619,N_5740);
nand U6860 (N_6860,N_5182,N_5555);
nand U6861 (N_6861,N_5995,N_5956);
and U6862 (N_6862,N_5085,N_5925);
and U6863 (N_6863,N_5208,N_5816);
or U6864 (N_6864,N_5237,N_5419);
and U6865 (N_6865,N_5980,N_5954);
nand U6866 (N_6866,N_5246,N_5249);
nand U6867 (N_6867,N_5087,N_5520);
nor U6868 (N_6868,N_5303,N_5998);
or U6869 (N_6869,N_5941,N_5770);
and U6870 (N_6870,N_5751,N_5842);
nand U6871 (N_6871,N_5220,N_5866);
or U6872 (N_6872,N_5104,N_5690);
nand U6873 (N_6873,N_5590,N_5662);
and U6874 (N_6874,N_5035,N_5919);
and U6875 (N_6875,N_5285,N_5232);
nor U6876 (N_6876,N_5592,N_5258);
and U6877 (N_6877,N_5518,N_5161);
nand U6878 (N_6878,N_5847,N_5305);
or U6879 (N_6879,N_5311,N_5078);
and U6880 (N_6880,N_5067,N_5954);
or U6881 (N_6881,N_5934,N_5198);
and U6882 (N_6882,N_5122,N_5296);
nor U6883 (N_6883,N_5970,N_5909);
and U6884 (N_6884,N_5148,N_5281);
or U6885 (N_6885,N_5273,N_5252);
or U6886 (N_6886,N_5672,N_5270);
nand U6887 (N_6887,N_5132,N_5069);
nor U6888 (N_6888,N_5455,N_5576);
or U6889 (N_6889,N_5009,N_5185);
nor U6890 (N_6890,N_5085,N_5213);
nor U6891 (N_6891,N_5801,N_5123);
nand U6892 (N_6892,N_5647,N_5877);
and U6893 (N_6893,N_5954,N_5881);
nand U6894 (N_6894,N_5484,N_5321);
nor U6895 (N_6895,N_5030,N_5435);
and U6896 (N_6896,N_5281,N_5925);
nand U6897 (N_6897,N_5964,N_5799);
nand U6898 (N_6898,N_5927,N_5421);
or U6899 (N_6899,N_5909,N_5610);
nand U6900 (N_6900,N_5272,N_5156);
and U6901 (N_6901,N_5120,N_5828);
nand U6902 (N_6902,N_5146,N_5822);
and U6903 (N_6903,N_5240,N_5463);
and U6904 (N_6904,N_5986,N_5604);
nor U6905 (N_6905,N_5921,N_5513);
nand U6906 (N_6906,N_5256,N_5432);
or U6907 (N_6907,N_5713,N_5032);
and U6908 (N_6908,N_5304,N_5455);
nand U6909 (N_6909,N_5699,N_5313);
nor U6910 (N_6910,N_5800,N_5008);
xnor U6911 (N_6911,N_5581,N_5981);
nor U6912 (N_6912,N_5830,N_5841);
or U6913 (N_6913,N_5960,N_5446);
and U6914 (N_6914,N_5679,N_5196);
nand U6915 (N_6915,N_5892,N_5840);
nor U6916 (N_6916,N_5209,N_5557);
and U6917 (N_6917,N_5410,N_5485);
nor U6918 (N_6918,N_5084,N_5185);
xor U6919 (N_6919,N_5933,N_5100);
nand U6920 (N_6920,N_5030,N_5668);
nor U6921 (N_6921,N_5692,N_5446);
nand U6922 (N_6922,N_5229,N_5577);
or U6923 (N_6923,N_5022,N_5797);
nor U6924 (N_6924,N_5736,N_5187);
or U6925 (N_6925,N_5897,N_5140);
nor U6926 (N_6926,N_5965,N_5740);
and U6927 (N_6927,N_5607,N_5283);
and U6928 (N_6928,N_5485,N_5802);
nand U6929 (N_6929,N_5119,N_5895);
or U6930 (N_6930,N_5081,N_5482);
and U6931 (N_6931,N_5961,N_5842);
or U6932 (N_6932,N_5621,N_5009);
or U6933 (N_6933,N_5417,N_5325);
and U6934 (N_6934,N_5788,N_5329);
or U6935 (N_6935,N_5105,N_5135);
nor U6936 (N_6936,N_5376,N_5423);
nand U6937 (N_6937,N_5993,N_5660);
nor U6938 (N_6938,N_5676,N_5105);
nand U6939 (N_6939,N_5407,N_5758);
nand U6940 (N_6940,N_5567,N_5447);
nand U6941 (N_6941,N_5028,N_5414);
or U6942 (N_6942,N_5386,N_5928);
and U6943 (N_6943,N_5892,N_5573);
and U6944 (N_6944,N_5573,N_5521);
or U6945 (N_6945,N_5902,N_5573);
nand U6946 (N_6946,N_5894,N_5342);
or U6947 (N_6947,N_5320,N_5664);
nor U6948 (N_6948,N_5846,N_5603);
or U6949 (N_6949,N_5456,N_5955);
and U6950 (N_6950,N_5605,N_5663);
nor U6951 (N_6951,N_5040,N_5446);
nand U6952 (N_6952,N_5160,N_5451);
or U6953 (N_6953,N_5080,N_5089);
nor U6954 (N_6954,N_5484,N_5047);
nor U6955 (N_6955,N_5387,N_5051);
nor U6956 (N_6956,N_5815,N_5007);
and U6957 (N_6957,N_5868,N_5821);
xnor U6958 (N_6958,N_5913,N_5506);
or U6959 (N_6959,N_5650,N_5664);
xnor U6960 (N_6960,N_5785,N_5667);
nor U6961 (N_6961,N_5740,N_5355);
nand U6962 (N_6962,N_5259,N_5075);
nand U6963 (N_6963,N_5756,N_5187);
nor U6964 (N_6964,N_5626,N_5341);
nand U6965 (N_6965,N_5353,N_5065);
nor U6966 (N_6966,N_5517,N_5396);
nor U6967 (N_6967,N_5089,N_5159);
and U6968 (N_6968,N_5518,N_5800);
nor U6969 (N_6969,N_5680,N_5127);
nor U6970 (N_6970,N_5440,N_5801);
nand U6971 (N_6971,N_5180,N_5868);
nor U6972 (N_6972,N_5679,N_5065);
or U6973 (N_6973,N_5691,N_5167);
or U6974 (N_6974,N_5987,N_5668);
and U6975 (N_6975,N_5997,N_5234);
nand U6976 (N_6976,N_5003,N_5107);
nor U6977 (N_6977,N_5977,N_5137);
nor U6978 (N_6978,N_5144,N_5826);
and U6979 (N_6979,N_5834,N_5261);
or U6980 (N_6980,N_5808,N_5315);
or U6981 (N_6981,N_5426,N_5556);
xor U6982 (N_6982,N_5481,N_5092);
nor U6983 (N_6983,N_5183,N_5379);
and U6984 (N_6984,N_5510,N_5819);
and U6985 (N_6985,N_5610,N_5549);
nor U6986 (N_6986,N_5720,N_5411);
and U6987 (N_6987,N_5137,N_5922);
nor U6988 (N_6988,N_5912,N_5683);
nand U6989 (N_6989,N_5155,N_5737);
and U6990 (N_6990,N_5267,N_5627);
or U6991 (N_6991,N_5606,N_5085);
or U6992 (N_6992,N_5584,N_5421);
or U6993 (N_6993,N_5160,N_5124);
nand U6994 (N_6994,N_5591,N_5949);
or U6995 (N_6995,N_5808,N_5163);
nand U6996 (N_6996,N_5918,N_5972);
nor U6997 (N_6997,N_5706,N_5821);
or U6998 (N_6998,N_5242,N_5930);
or U6999 (N_6999,N_5554,N_5572);
or U7000 (N_7000,N_6730,N_6686);
nor U7001 (N_7001,N_6605,N_6057);
nor U7002 (N_7002,N_6844,N_6722);
nor U7003 (N_7003,N_6525,N_6716);
nand U7004 (N_7004,N_6719,N_6646);
nor U7005 (N_7005,N_6884,N_6704);
nand U7006 (N_7006,N_6827,N_6179);
nor U7007 (N_7007,N_6176,N_6718);
nor U7008 (N_7008,N_6361,N_6239);
or U7009 (N_7009,N_6548,N_6208);
nand U7010 (N_7010,N_6283,N_6602);
nor U7011 (N_7011,N_6786,N_6712);
and U7012 (N_7012,N_6263,N_6741);
nor U7013 (N_7013,N_6643,N_6403);
nor U7014 (N_7014,N_6818,N_6784);
or U7015 (N_7015,N_6628,N_6392);
nand U7016 (N_7016,N_6455,N_6321);
nand U7017 (N_7017,N_6995,N_6408);
nor U7018 (N_7018,N_6214,N_6400);
or U7019 (N_7019,N_6567,N_6039);
or U7020 (N_7020,N_6510,N_6511);
or U7021 (N_7021,N_6865,N_6987);
and U7022 (N_7022,N_6048,N_6217);
nand U7023 (N_7023,N_6087,N_6934);
nor U7024 (N_7024,N_6846,N_6055);
and U7025 (N_7025,N_6919,N_6738);
nor U7026 (N_7026,N_6874,N_6761);
nand U7027 (N_7027,N_6094,N_6853);
and U7028 (N_7028,N_6804,N_6487);
and U7029 (N_7029,N_6880,N_6817);
or U7030 (N_7030,N_6968,N_6090);
nand U7031 (N_7031,N_6886,N_6261);
and U7032 (N_7032,N_6414,N_6042);
nor U7033 (N_7033,N_6689,N_6550);
nand U7034 (N_7034,N_6774,N_6503);
or U7035 (N_7035,N_6514,N_6649);
and U7036 (N_7036,N_6418,N_6611);
and U7037 (N_7037,N_6106,N_6275);
nand U7038 (N_7038,N_6464,N_6703);
and U7039 (N_7039,N_6007,N_6151);
and U7040 (N_7040,N_6492,N_6921);
or U7041 (N_7041,N_6731,N_6759);
and U7042 (N_7042,N_6837,N_6384);
nor U7043 (N_7043,N_6970,N_6972);
and U7044 (N_7044,N_6035,N_6120);
nor U7045 (N_7045,N_6931,N_6808);
nor U7046 (N_7046,N_6389,N_6775);
nand U7047 (N_7047,N_6359,N_6407);
nand U7048 (N_7048,N_6144,N_6073);
nand U7049 (N_7049,N_6269,N_6481);
nand U7050 (N_7050,N_6991,N_6413);
nor U7051 (N_7051,N_6746,N_6566);
and U7052 (N_7052,N_6131,N_6586);
and U7053 (N_7053,N_6427,N_6678);
nor U7054 (N_7054,N_6146,N_6443);
nand U7055 (N_7055,N_6964,N_6847);
or U7056 (N_7056,N_6474,N_6002);
and U7057 (N_7057,N_6982,N_6938);
or U7058 (N_7058,N_6973,N_6658);
nand U7059 (N_7059,N_6875,N_6905);
nand U7060 (N_7060,N_6133,N_6186);
and U7061 (N_7061,N_6171,N_6500);
nor U7062 (N_7062,N_6252,N_6614);
nand U7063 (N_7063,N_6101,N_6249);
or U7064 (N_7064,N_6089,N_6922);
nand U7065 (N_7065,N_6780,N_6218);
nor U7066 (N_7066,N_6635,N_6383);
or U7067 (N_7067,N_6562,N_6612);
nand U7068 (N_7068,N_6054,N_6149);
nand U7069 (N_7069,N_6692,N_6984);
nand U7070 (N_7070,N_6636,N_6810);
or U7071 (N_7071,N_6452,N_6100);
or U7072 (N_7072,N_6713,N_6023);
and U7073 (N_7073,N_6994,N_6422);
and U7074 (N_7074,N_6833,N_6765);
or U7075 (N_7075,N_6341,N_6637);
or U7076 (N_7076,N_6734,N_6793);
or U7077 (N_7077,N_6264,N_6175);
and U7078 (N_7078,N_6822,N_6224);
and U7079 (N_7079,N_6132,N_6721);
and U7080 (N_7080,N_6729,N_6438);
nand U7081 (N_7081,N_6490,N_6673);
and U7082 (N_7082,N_6065,N_6642);
xnor U7083 (N_7083,N_6768,N_6631);
or U7084 (N_7084,N_6084,N_6395);
nor U7085 (N_7085,N_6296,N_6509);
and U7086 (N_7086,N_6109,N_6951);
and U7087 (N_7087,N_6419,N_6573);
and U7088 (N_7088,N_6273,N_6235);
nor U7089 (N_7089,N_6394,N_6346);
and U7090 (N_7090,N_6213,N_6289);
and U7091 (N_7091,N_6410,N_6621);
nor U7092 (N_7092,N_6943,N_6772);
nor U7093 (N_7093,N_6033,N_6879);
nor U7094 (N_7094,N_6486,N_6744);
nor U7095 (N_7095,N_6623,N_6396);
nand U7096 (N_7096,N_6809,N_6032);
or U7097 (N_7097,N_6472,N_6776);
and U7098 (N_7098,N_6368,N_6428);
or U7099 (N_7099,N_6766,N_6197);
nand U7100 (N_7100,N_6430,N_6764);
or U7101 (N_7101,N_6720,N_6163);
or U7102 (N_7102,N_6381,N_6520);
and U7103 (N_7103,N_6652,N_6831);
nand U7104 (N_7104,N_6778,N_6981);
nand U7105 (N_7105,N_6480,N_6282);
and U7106 (N_7106,N_6947,N_6702);
nand U7107 (N_7107,N_6745,N_6290);
nor U7108 (N_7108,N_6390,N_6555);
nor U7109 (N_7109,N_6459,N_6018);
and U7110 (N_7110,N_6295,N_6782);
or U7111 (N_7111,N_6700,N_6022);
and U7112 (N_7112,N_6626,N_6170);
nor U7113 (N_7113,N_6547,N_6963);
nand U7114 (N_7114,N_6536,N_6255);
or U7115 (N_7115,N_6425,N_6851);
nand U7116 (N_7116,N_6328,N_6306);
and U7117 (N_7117,N_6158,N_6749);
or U7118 (N_7118,N_6429,N_6325);
nor U7119 (N_7119,N_6339,N_6103);
nand U7120 (N_7120,N_6667,N_6406);
or U7121 (N_7121,N_6250,N_6788);
nand U7122 (N_7122,N_6156,N_6754);
nand U7123 (N_7123,N_6253,N_6832);
nor U7124 (N_7124,N_6639,N_6236);
nor U7125 (N_7125,N_6501,N_6209);
and U7126 (N_7126,N_6969,N_6811);
or U7127 (N_7127,N_6191,N_6086);
nor U7128 (N_7128,N_6527,N_6949);
or U7129 (N_7129,N_6067,N_6587);
or U7130 (N_7130,N_6929,N_6351);
or U7131 (N_7131,N_6079,N_6228);
nor U7132 (N_7132,N_6551,N_6600);
and U7133 (N_7133,N_6552,N_6796);
nor U7134 (N_7134,N_6985,N_6860);
nand U7135 (N_7135,N_6373,N_6743);
nand U7136 (N_7136,N_6937,N_6902);
and U7137 (N_7137,N_6893,N_6004);
or U7138 (N_7138,N_6823,N_6996);
nand U7139 (N_7139,N_6841,N_6198);
nor U7140 (N_7140,N_6595,N_6767);
and U7141 (N_7141,N_6312,N_6756);
nand U7142 (N_7142,N_6866,N_6983);
nand U7143 (N_7143,N_6226,N_6540);
or U7144 (N_7144,N_6855,N_6141);
and U7145 (N_7145,N_6870,N_6280);
and U7146 (N_7146,N_6961,N_6739);
nand U7147 (N_7147,N_6203,N_6737);
nor U7148 (N_7148,N_6517,N_6225);
xnor U7149 (N_7149,N_6411,N_6461);
and U7150 (N_7150,N_6783,N_6584);
or U7151 (N_7151,N_6518,N_6493);
and U7152 (N_7152,N_6709,N_6498);
nand U7153 (N_7153,N_6303,N_6974);
and U7154 (N_7154,N_6695,N_6155);
nand U7155 (N_7155,N_6168,N_6491);
nand U7156 (N_7156,N_6190,N_6681);
nand U7157 (N_7157,N_6085,N_6593);
and U7158 (N_7158,N_6950,N_6046);
or U7159 (N_7159,N_6183,N_6201);
nand U7160 (N_7160,N_6840,N_6078);
nor U7161 (N_7161,N_6838,N_6558);
and U7162 (N_7162,N_6473,N_6512);
and U7163 (N_7163,N_6115,N_6260);
or U7164 (N_7164,N_6001,N_6535);
nand U7165 (N_7165,N_6244,N_6797);
or U7166 (N_7166,N_6915,N_6672);
nor U7167 (N_7167,N_6760,N_6450);
nor U7168 (N_7168,N_6895,N_6173);
nand U7169 (N_7169,N_6789,N_6670);
nor U7170 (N_7170,N_6869,N_6699);
and U7171 (N_7171,N_6129,N_6080);
and U7172 (N_7172,N_6736,N_6420);
nor U7173 (N_7173,N_6868,N_6959);
nand U7174 (N_7174,N_6458,N_6800);
and U7175 (N_7175,N_6528,N_6694);
or U7176 (N_7176,N_6861,N_6590);
nand U7177 (N_7177,N_6316,N_6139);
nor U7178 (N_7178,N_6640,N_6696);
or U7179 (N_7179,N_6948,N_6653);
or U7180 (N_7180,N_6070,N_6248);
and U7181 (N_7181,N_6380,N_6000);
or U7182 (N_7182,N_6241,N_6708);
nor U7183 (N_7183,N_6656,N_6284);
nand U7184 (N_7184,N_6852,N_6591);
nor U7185 (N_7185,N_6143,N_6082);
and U7186 (N_7186,N_6238,N_6757);
and U7187 (N_7187,N_6638,N_6154);
nor U7188 (N_7188,N_6166,N_6034);
nand U7189 (N_7189,N_6415,N_6469);
nand U7190 (N_7190,N_6231,N_6634);
and U7191 (N_7191,N_6302,N_6012);
or U7192 (N_7192,N_6119,N_6265);
nor U7193 (N_7193,N_6615,N_6051);
or U7194 (N_7194,N_6740,N_6899);
nand U7195 (N_7195,N_6912,N_6799);
nor U7196 (N_7196,N_6401,N_6598);
nand U7197 (N_7197,N_6906,N_6463);
nor U7198 (N_7198,N_6669,N_6690);
or U7199 (N_7199,N_6336,N_6127);
or U7200 (N_7200,N_6954,N_6907);
and U7201 (N_7201,N_6077,N_6358);
or U7202 (N_7202,N_6845,N_6858);
nand U7203 (N_7203,N_6281,N_6113);
and U7204 (N_7204,N_6484,N_6769);
nand U7205 (N_7205,N_6436,N_6362);
nor U7206 (N_7206,N_6539,N_6045);
or U7207 (N_7207,N_6188,N_6409);
or U7208 (N_7208,N_6570,N_6684);
and U7209 (N_7209,N_6385,N_6569);
nand U7210 (N_7210,N_6021,N_6989);
and U7211 (N_7211,N_6076,N_6439);
and U7212 (N_7212,N_6462,N_6148);
nand U7213 (N_7213,N_6763,N_6011);
and U7214 (N_7214,N_6495,N_6262);
nand U7215 (N_7215,N_6522,N_6955);
nor U7216 (N_7216,N_6355,N_6117);
nor U7217 (N_7217,N_6710,N_6583);
or U7218 (N_7218,N_6388,N_6025);
xor U7219 (N_7219,N_6717,N_6125);
and U7220 (N_7220,N_6830,N_6606);
xnor U7221 (N_7221,N_6668,N_6812);
and U7222 (N_7222,N_6999,N_6327);
or U7223 (N_7223,N_6572,N_6102);
or U7224 (N_7224,N_6267,N_6864);
nand U7225 (N_7225,N_6294,N_6299);
or U7226 (N_7226,N_6003,N_6174);
nor U7227 (N_7227,N_6445,N_6180);
nand U7228 (N_7228,N_6935,N_6378);
nor U7229 (N_7229,N_6024,N_6863);
nand U7230 (N_7230,N_6081,N_6580);
nand U7231 (N_7231,N_6805,N_6167);
nand U7232 (N_7232,N_6072,N_6966);
nor U7233 (N_7233,N_6184,N_6609);
or U7234 (N_7234,N_6405,N_6872);
and U7235 (N_7235,N_6071,N_6530);
and U7236 (N_7236,N_6677,N_6816);
or U7237 (N_7237,N_6565,N_6399);
nand U7238 (N_7238,N_6010,N_6885);
nand U7239 (N_7239,N_6376,N_6220);
xnor U7240 (N_7240,N_6978,N_6479);
nor U7241 (N_7241,N_6629,N_6293);
or U7242 (N_7242,N_6502,N_6112);
or U7243 (N_7243,N_6212,N_6013);
and U7244 (N_7244,N_6040,N_6633);
nor U7245 (N_7245,N_6354,N_6664);
or U7246 (N_7246,N_6541,N_6854);
or U7247 (N_7247,N_6930,N_6630);
nor U7248 (N_7248,N_6925,N_6448);
or U7249 (N_7249,N_6862,N_6216);
or U7250 (N_7250,N_6137,N_6140);
nand U7251 (N_7251,N_6457,N_6795);
nand U7252 (N_7252,N_6204,N_6391);
nor U7253 (N_7253,N_6068,N_6271);
and U7254 (N_7254,N_6613,N_6478);
and U7255 (N_7255,N_6733,N_6471);
nor U7256 (N_7256,N_6524,N_6309);
nor U7257 (N_7257,N_6297,N_6229);
nand U7258 (N_7258,N_6485,N_6957);
nor U7259 (N_7259,N_6753,N_6178);
nand U7260 (N_7260,N_6298,N_6971);
nand U7261 (N_7261,N_6210,N_6857);
nand U7262 (N_7262,N_6116,N_6393);
nand U7263 (N_7263,N_6421,N_6932);
nor U7264 (N_7264,N_6849,N_6728);
nand U7265 (N_7265,N_6891,N_6697);
nand U7266 (N_7266,N_6515,N_6601);
or U7267 (N_7267,N_6794,N_6815);
or U7268 (N_7268,N_6751,N_6563);
nand U7269 (N_7269,N_6977,N_6015);
nor U7270 (N_7270,N_6927,N_6211);
or U7271 (N_7271,N_6657,N_6301);
and U7272 (N_7272,N_6432,N_6650);
and U7273 (N_7273,N_6453,N_6227);
or U7274 (N_7274,N_6205,N_6506);
and U7275 (N_7275,N_6560,N_6901);
or U7276 (N_7276,N_6997,N_6993);
and U7277 (N_7277,N_6890,N_6913);
nor U7278 (N_7278,N_6529,N_6582);
nand U7279 (N_7279,N_6813,N_6159);
nor U7280 (N_7280,N_6056,N_6941);
nor U7281 (N_7281,N_6526,N_6437);
nor U7282 (N_7282,N_6988,N_6049);
xnor U7283 (N_7283,N_6898,N_6596);
and U7284 (N_7284,N_6771,N_6758);
nand U7285 (N_7285,N_6559,N_6091);
nor U7286 (N_7286,N_6460,N_6377);
and U7287 (N_7287,N_6122,N_6561);
nor U7288 (N_7288,N_6404,N_6732);
nand U7289 (N_7289,N_6335,N_6641);
nand U7290 (N_7290,N_6504,N_6807);
and U7291 (N_7291,N_6366,N_6234);
nand U7292 (N_7292,N_6918,N_6575);
and U7293 (N_7293,N_6599,N_6288);
nor U7294 (N_7294,N_6343,N_6270);
nand U7295 (N_7295,N_6172,N_6333);
or U7296 (N_7296,N_6417,N_6062);
nor U7297 (N_7297,N_6826,N_6568);
nand U7298 (N_7298,N_6037,N_6016);
xnor U7299 (N_7299,N_6338,N_6747);
nor U7300 (N_7300,N_6367,N_6625);
and U7301 (N_7301,N_6310,N_6546);
or U7302 (N_7302,N_6387,N_6268);
nor U7303 (N_7303,N_6726,N_6342);
and U7304 (N_7304,N_6029,N_6990);
nand U7305 (N_7305,N_6014,N_6256);
or U7306 (N_7306,N_6277,N_6130);
and U7307 (N_7307,N_6074,N_6878);
and U7308 (N_7308,N_6099,N_6892);
nor U7309 (N_7309,N_6451,N_6727);
nor U7310 (N_7310,N_6603,N_6416);
nor U7311 (N_7311,N_6661,N_6352);
nor U7312 (N_7312,N_6701,N_6320);
nor U7313 (N_7313,N_6693,N_6199);
nand U7314 (N_7314,N_6910,N_6365);
nand U7315 (N_7315,N_6126,N_6319);
or U7316 (N_7316,N_6802,N_6223);
nor U7317 (N_7317,N_6556,N_6585);
or U7318 (N_7318,N_6494,N_6960);
nand U7319 (N_7319,N_6324,N_6412);
nand U7320 (N_7320,N_6287,N_6110);
nor U7321 (N_7321,N_6928,N_6476);
or U7322 (N_7322,N_6364,N_6020);
nor U7323 (N_7323,N_6242,N_6781);
nand U7324 (N_7324,N_6124,N_6105);
or U7325 (N_7325,N_6315,N_6247);
xor U7326 (N_7326,N_6647,N_6617);
nand U7327 (N_7327,N_6705,N_6026);
and U7328 (N_7328,N_6592,N_6334);
and U7329 (N_7329,N_6276,N_6069);
and U7330 (N_7330,N_6604,N_6888);
and U7331 (N_7331,N_6006,N_6663);
or U7332 (N_7332,N_6157,N_6724);
and U7333 (N_7333,N_6544,N_6440);
nor U7334 (N_7334,N_6542,N_6979);
and U7335 (N_7335,N_6322,N_6725);
nand U7336 (N_7336,N_6128,N_6152);
nand U7337 (N_7337,N_6571,N_6382);
and U7338 (N_7338,N_6723,N_6791);
or U7339 (N_7339,N_6329,N_6537);
nand U7340 (N_7340,N_6926,N_6292);
or U7341 (N_7341,N_6060,N_6254);
nand U7342 (N_7342,N_6221,N_6347);
nand U7343 (N_7343,N_6353,N_6043);
and U7344 (N_7344,N_6017,N_6967);
and U7345 (N_7345,N_6008,N_6240);
nand U7346 (N_7346,N_6145,N_6616);
nand U7347 (N_7347,N_6521,N_6659);
nor U7348 (N_7348,N_6665,N_6036);
or U7349 (N_7349,N_6588,N_6850);
nor U7350 (N_7350,N_6904,N_6134);
nand U7351 (N_7351,N_6645,N_6750);
and U7352 (N_7352,N_6363,N_6933);
nor U7353 (N_7353,N_6181,N_6532);
nor U7354 (N_7354,N_6369,N_6835);
nor U7355 (N_7355,N_6897,N_6958);
nand U7356 (N_7356,N_6044,N_6516);
and U7357 (N_7357,N_6513,N_6272);
nand U7358 (N_7358,N_6308,N_6924);
and U7359 (N_7359,N_6679,N_6031);
nor U7360 (N_7360,N_6607,N_6192);
and U7361 (N_7361,N_6375,N_6285);
nor U7362 (N_7362,N_6965,N_6956);
or U7363 (N_7363,N_6326,N_6589);
nor U7364 (N_7364,N_6887,N_6028);
xnor U7365 (N_7365,N_6447,N_6944);
and U7366 (N_7366,N_6488,N_6038);
or U7367 (N_7367,N_6859,N_6279);
nand U7368 (N_7368,N_6423,N_6896);
nand U7369 (N_7369,N_6624,N_6196);
or U7370 (N_7370,N_6942,N_6274);
nand U7371 (N_7371,N_6877,N_6632);
and U7372 (N_7372,N_6454,N_6222);
nand U7373 (N_7373,N_6497,N_6666);
and U7374 (N_7374,N_6111,N_6576);
nor U7375 (N_7375,N_6092,N_6803);
nor U7376 (N_7376,N_6779,N_6323);
nand U7377 (N_7377,N_6675,N_6792);
nand U7378 (N_7378,N_6153,N_6998);
or U7379 (N_7379,N_6442,N_6917);
nand U7380 (N_7380,N_6059,N_6194);
or U7381 (N_7381,N_6356,N_6662);
nand U7382 (N_7382,N_6903,N_6259);
nand U7383 (N_7383,N_6441,N_6920);
and U7384 (N_7384,N_6909,N_6519);
and U7385 (N_7385,N_6187,N_6098);
nor U7386 (N_7386,N_6431,N_6135);
or U7387 (N_7387,N_6466,N_6755);
or U7388 (N_7388,N_6711,N_6052);
nor U7389 (N_7389,N_6142,N_6842);
nand U7390 (N_7390,N_6345,N_6574);
nor U7391 (N_7391,N_6762,N_6372);
nand U7392 (N_7392,N_6608,N_6660);
and U7393 (N_7393,N_6348,N_6121);
nor U7394 (N_7394,N_6360,N_6939);
or U7395 (N_7395,N_6064,N_6344);
and U7396 (N_7396,N_6610,N_6233);
nand U7397 (N_7397,N_6900,N_6714);
nor U7398 (N_7398,N_6332,N_6206);
or U7399 (N_7399,N_6300,N_6848);
nor U7400 (N_7400,N_6834,N_6164);
nand U7401 (N_7401,N_6169,N_6165);
or U7402 (N_7402,N_6397,N_6370);
nand U7403 (N_7403,N_6806,N_6200);
or U7404 (N_7404,N_6123,N_6682);
or U7405 (N_7405,N_6337,N_6019);
and U7406 (N_7406,N_6785,N_6053);
or U7407 (N_7407,N_6482,N_6041);
or U7408 (N_7408,N_6821,N_6618);
nand U7409 (N_7409,N_6873,N_6871);
nand U7410 (N_7410,N_6150,N_6108);
or U7411 (N_7411,N_6676,N_6278);
and U7412 (N_7412,N_6202,N_6581);
nor U7413 (N_7413,N_6651,N_6433);
nor U7414 (N_7414,N_6386,N_6047);
and U7415 (N_7415,N_6882,N_6975);
and U7416 (N_7416,N_6554,N_6061);
or U7417 (N_7417,N_6820,N_6507);
nor U7418 (N_7418,N_6465,N_6467);
or U7419 (N_7419,N_6976,N_6477);
and U7420 (N_7420,N_6688,N_6856);
nor U7421 (N_7421,N_6538,N_6883);
nor U7422 (N_7422,N_6685,N_6160);
nand U7423 (N_7423,N_6162,N_6923);
or U7424 (N_7424,N_6083,N_6009);
nor U7425 (N_7425,N_6096,N_6182);
nand U7426 (N_7426,N_6777,N_6379);
and U7427 (N_7427,N_6374,N_6371);
and U7428 (N_7428,N_6946,N_6246);
and U7429 (N_7429,N_6534,N_6398);
nand U7430 (N_7430,N_6671,N_6444);
nor U7431 (N_7431,N_6889,N_6219);
or U7432 (N_7432,N_6350,N_6402);
and U7433 (N_7433,N_6814,N_6237);
nor U7434 (N_7434,N_6908,N_6770);
and U7435 (N_7435,N_6251,N_6523);
nand U7436 (N_7436,N_6449,N_6962);
and U7437 (N_7437,N_6655,N_6489);
or U7438 (N_7438,N_6118,N_6881);
nor U7439 (N_7439,N_6095,N_6185);
or U7440 (N_7440,N_6426,N_6093);
nor U7441 (N_7441,N_6245,N_6620);
nor U7442 (N_7442,N_6557,N_6564);
nand U7443 (N_7443,N_6674,N_6331);
nor U7444 (N_7444,N_6483,N_6136);
and U7445 (N_7445,N_6468,N_6340);
nand U7446 (N_7446,N_6005,N_6195);
nand U7447 (N_7447,N_6953,N_6470);
or U7448 (N_7448,N_6986,N_6742);
and U7449 (N_7449,N_6230,N_6435);
or U7450 (N_7450,N_6258,N_6050);
nand U7451 (N_7451,N_6773,N_6533);
and U7452 (N_7452,N_6475,N_6058);
and U7453 (N_7453,N_6215,N_6286);
or U7454 (N_7454,N_6867,N_6543);
and U7455 (N_7455,N_6828,N_6619);
nor U7456 (N_7456,N_6945,N_6578);
and U7457 (N_7457,N_6314,N_6992);
nand U7458 (N_7458,N_6683,N_6097);
nor U7459 (N_7459,N_6177,N_6232);
nor U7460 (N_7460,N_6207,N_6911);
nor U7461 (N_7461,N_6706,N_6843);
or U7462 (N_7462,N_6138,N_6648);
or U7463 (N_7463,N_6318,N_6107);
and U7464 (N_7464,N_6577,N_6496);
nor U7465 (N_7465,N_6824,N_6499);
or U7466 (N_7466,N_6829,N_6114);
nor U7467 (N_7467,N_6916,N_6066);
nand U7468 (N_7468,N_6549,N_6839);
nor U7469 (N_7469,N_6257,N_6189);
or U7470 (N_7470,N_6307,N_6266);
nand U7471 (N_7471,N_6305,N_6894);
nand U7472 (N_7472,N_6952,N_6752);
and U7473 (N_7473,N_6545,N_6627);
nor U7474 (N_7474,N_6357,N_6707);
and U7475 (N_7475,N_6715,N_6594);
and U7476 (N_7476,N_6748,N_6508);
nor U7477 (N_7477,N_6349,N_6243);
and U7478 (N_7478,N_6456,N_6330);
nor U7479 (N_7479,N_6836,N_6597);
nor U7480 (N_7480,N_6434,N_6825);
and U7481 (N_7481,N_6553,N_6088);
and U7482 (N_7482,N_6063,N_6940);
and U7483 (N_7483,N_6790,N_6193);
nor U7484 (N_7484,N_6313,N_6161);
nor U7485 (N_7485,N_6798,N_6819);
nor U7486 (N_7486,N_6698,N_6075);
xnor U7487 (N_7487,N_6531,N_6687);
and U7488 (N_7488,N_6304,N_6980);
or U7489 (N_7489,N_6680,N_6914);
and U7490 (N_7490,N_6147,N_6104);
or U7491 (N_7491,N_6579,N_6424);
or U7492 (N_7492,N_6027,N_6936);
and U7493 (N_7493,N_6311,N_6622);
xnor U7494 (N_7494,N_6801,N_6291);
and U7495 (N_7495,N_6317,N_6654);
nand U7496 (N_7496,N_6735,N_6030);
and U7497 (N_7497,N_6787,N_6876);
and U7498 (N_7498,N_6644,N_6691);
or U7499 (N_7499,N_6505,N_6446);
nand U7500 (N_7500,N_6905,N_6380);
and U7501 (N_7501,N_6568,N_6467);
or U7502 (N_7502,N_6761,N_6322);
nand U7503 (N_7503,N_6099,N_6554);
and U7504 (N_7504,N_6293,N_6276);
or U7505 (N_7505,N_6611,N_6657);
xor U7506 (N_7506,N_6065,N_6100);
and U7507 (N_7507,N_6947,N_6009);
and U7508 (N_7508,N_6313,N_6461);
nand U7509 (N_7509,N_6335,N_6840);
nand U7510 (N_7510,N_6795,N_6792);
and U7511 (N_7511,N_6800,N_6905);
nand U7512 (N_7512,N_6488,N_6517);
or U7513 (N_7513,N_6027,N_6793);
or U7514 (N_7514,N_6359,N_6659);
nand U7515 (N_7515,N_6536,N_6277);
or U7516 (N_7516,N_6439,N_6697);
and U7517 (N_7517,N_6475,N_6472);
or U7518 (N_7518,N_6503,N_6387);
nand U7519 (N_7519,N_6907,N_6688);
nor U7520 (N_7520,N_6621,N_6023);
nor U7521 (N_7521,N_6062,N_6016);
nor U7522 (N_7522,N_6870,N_6212);
or U7523 (N_7523,N_6240,N_6211);
nand U7524 (N_7524,N_6063,N_6846);
or U7525 (N_7525,N_6671,N_6868);
or U7526 (N_7526,N_6770,N_6081);
or U7527 (N_7527,N_6956,N_6127);
or U7528 (N_7528,N_6659,N_6917);
xnor U7529 (N_7529,N_6420,N_6471);
nor U7530 (N_7530,N_6390,N_6942);
nand U7531 (N_7531,N_6934,N_6323);
nor U7532 (N_7532,N_6790,N_6553);
nor U7533 (N_7533,N_6334,N_6295);
and U7534 (N_7534,N_6835,N_6858);
nand U7535 (N_7535,N_6603,N_6240);
or U7536 (N_7536,N_6331,N_6846);
nor U7537 (N_7537,N_6671,N_6057);
nand U7538 (N_7538,N_6830,N_6003);
and U7539 (N_7539,N_6943,N_6154);
and U7540 (N_7540,N_6953,N_6314);
nor U7541 (N_7541,N_6776,N_6122);
and U7542 (N_7542,N_6877,N_6305);
or U7543 (N_7543,N_6018,N_6475);
or U7544 (N_7544,N_6035,N_6485);
nor U7545 (N_7545,N_6265,N_6504);
and U7546 (N_7546,N_6313,N_6319);
or U7547 (N_7547,N_6542,N_6437);
and U7548 (N_7548,N_6930,N_6601);
nor U7549 (N_7549,N_6989,N_6126);
nand U7550 (N_7550,N_6122,N_6754);
and U7551 (N_7551,N_6091,N_6425);
nand U7552 (N_7552,N_6421,N_6986);
or U7553 (N_7553,N_6803,N_6362);
nor U7554 (N_7554,N_6297,N_6555);
nand U7555 (N_7555,N_6501,N_6393);
and U7556 (N_7556,N_6424,N_6929);
nor U7557 (N_7557,N_6151,N_6602);
or U7558 (N_7558,N_6678,N_6952);
nor U7559 (N_7559,N_6577,N_6231);
or U7560 (N_7560,N_6918,N_6165);
or U7561 (N_7561,N_6489,N_6540);
nand U7562 (N_7562,N_6963,N_6664);
nor U7563 (N_7563,N_6496,N_6034);
nor U7564 (N_7564,N_6605,N_6867);
or U7565 (N_7565,N_6921,N_6442);
nand U7566 (N_7566,N_6192,N_6148);
or U7567 (N_7567,N_6556,N_6795);
nor U7568 (N_7568,N_6765,N_6058);
or U7569 (N_7569,N_6855,N_6815);
and U7570 (N_7570,N_6538,N_6414);
and U7571 (N_7571,N_6805,N_6937);
nor U7572 (N_7572,N_6690,N_6029);
xor U7573 (N_7573,N_6751,N_6958);
nand U7574 (N_7574,N_6054,N_6017);
and U7575 (N_7575,N_6075,N_6914);
and U7576 (N_7576,N_6950,N_6382);
and U7577 (N_7577,N_6341,N_6520);
nand U7578 (N_7578,N_6000,N_6492);
nand U7579 (N_7579,N_6187,N_6327);
nor U7580 (N_7580,N_6483,N_6932);
or U7581 (N_7581,N_6885,N_6986);
nand U7582 (N_7582,N_6895,N_6657);
or U7583 (N_7583,N_6026,N_6773);
nand U7584 (N_7584,N_6103,N_6758);
and U7585 (N_7585,N_6180,N_6458);
or U7586 (N_7586,N_6106,N_6811);
and U7587 (N_7587,N_6302,N_6292);
or U7588 (N_7588,N_6371,N_6798);
xor U7589 (N_7589,N_6583,N_6777);
nand U7590 (N_7590,N_6626,N_6566);
or U7591 (N_7591,N_6779,N_6341);
nor U7592 (N_7592,N_6040,N_6636);
or U7593 (N_7593,N_6325,N_6573);
nand U7594 (N_7594,N_6960,N_6626);
nor U7595 (N_7595,N_6472,N_6910);
nor U7596 (N_7596,N_6444,N_6823);
nor U7597 (N_7597,N_6179,N_6274);
nor U7598 (N_7598,N_6067,N_6702);
and U7599 (N_7599,N_6938,N_6092);
nor U7600 (N_7600,N_6743,N_6189);
nand U7601 (N_7601,N_6351,N_6163);
nand U7602 (N_7602,N_6908,N_6217);
or U7603 (N_7603,N_6856,N_6973);
nor U7604 (N_7604,N_6526,N_6904);
nor U7605 (N_7605,N_6407,N_6793);
and U7606 (N_7606,N_6155,N_6939);
nor U7607 (N_7607,N_6595,N_6449);
nand U7608 (N_7608,N_6057,N_6021);
or U7609 (N_7609,N_6976,N_6015);
nand U7610 (N_7610,N_6725,N_6970);
and U7611 (N_7611,N_6251,N_6324);
nor U7612 (N_7612,N_6119,N_6992);
nand U7613 (N_7613,N_6497,N_6737);
nor U7614 (N_7614,N_6277,N_6994);
or U7615 (N_7615,N_6846,N_6457);
or U7616 (N_7616,N_6340,N_6358);
nand U7617 (N_7617,N_6814,N_6233);
nor U7618 (N_7618,N_6166,N_6433);
or U7619 (N_7619,N_6697,N_6618);
and U7620 (N_7620,N_6246,N_6159);
nor U7621 (N_7621,N_6838,N_6372);
and U7622 (N_7622,N_6813,N_6888);
nand U7623 (N_7623,N_6008,N_6204);
nor U7624 (N_7624,N_6955,N_6214);
or U7625 (N_7625,N_6194,N_6924);
or U7626 (N_7626,N_6963,N_6964);
or U7627 (N_7627,N_6712,N_6515);
or U7628 (N_7628,N_6093,N_6468);
and U7629 (N_7629,N_6181,N_6342);
and U7630 (N_7630,N_6191,N_6357);
xnor U7631 (N_7631,N_6695,N_6086);
and U7632 (N_7632,N_6053,N_6122);
nor U7633 (N_7633,N_6747,N_6609);
and U7634 (N_7634,N_6625,N_6362);
nor U7635 (N_7635,N_6552,N_6914);
nor U7636 (N_7636,N_6102,N_6119);
nor U7637 (N_7637,N_6459,N_6625);
or U7638 (N_7638,N_6998,N_6106);
or U7639 (N_7639,N_6596,N_6128);
xor U7640 (N_7640,N_6545,N_6169);
and U7641 (N_7641,N_6316,N_6602);
or U7642 (N_7642,N_6378,N_6597);
nor U7643 (N_7643,N_6428,N_6991);
and U7644 (N_7644,N_6280,N_6211);
and U7645 (N_7645,N_6234,N_6671);
nand U7646 (N_7646,N_6399,N_6730);
nor U7647 (N_7647,N_6705,N_6976);
or U7648 (N_7648,N_6325,N_6129);
nor U7649 (N_7649,N_6576,N_6912);
nand U7650 (N_7650,N_6574,N_6724);
or U7651 (N_7651,N_6103,N_6879);
nand U7652 (N_7652,N_6855,N_6854);
and U7653 (N_7653,N_6022,N_6764);
nor U7654 (N_7654,N_6348,N_6044);
or U7655 (N_7655,N_6704,N_6297);
nand U7656 (N_7656,N_6368,N_6827);
nor U7657 (N_7657,N_6106,N_6343);
and U7658 (N_7658,N_6088,N_6948);
and U7659 (N_7659,N_6191,N_6133);
and U7660 (N_7660,N_6473,N_6188);
or U7661 (N_7661,N_6277,N_6717);
nand U7662 (N_7662,N_6739,N_6428);
nand U7663 (N_7663,N_6074,N_6023);
nand U7664 (N_7664,N_6614,N_6393);
nand U7665 (N_7665,N_6425,N_6835);
nor U7666 (N_7666,N_6635,N_6430);
and U7667 (N_7667,N_6877,N_6787);
nand U7668 (N_7668,N_6134,N_6401);
nand U7669 (N_7669,N_6795,N_6587);
nand U7670 (N_7670,N_6449,N_6624);
or U7671 (N_7671,N_6783,N_6281);
nor U7672 (N_7672,N_6883,N_6486);
nand U7673 (N_7673,N_6828,N_6444);
or U7674 (N_7674,N_6305,N_6871);
nand U7675 (N_7675,N_6368,N_6077);
nor U7676 (N_7676,N_6894,N_6394);
or U7677 (N_7677,N_6689,N_6248);
nor U7678 (N_7678,N_6382,N_6968);
and U7679 (N_7679,N_6531,N_6497);
or U7680 (N_7680,N_6628,N_6355);
nor U7681 (N_7681,N_6985,N_6089);
nor U7682 (N_7682,N_6251,N_6202);
and U7683 (N_7683,N_6304,N_6212);
and U7684 (N_7684,N_6779,N_6672);
nand U7685 (N_7685,N_6518,N_6990);
nor U7686 (N_7686,N_6534,N_6863);
or U7687 (N_7687,N_6588,N_6561);
nand U7688 (N_7688,N_6810,N_6717);
and U7689 (N_7689,N_6654,N_6591);
and U7690 (N_7690,N_6199,N_6615);
and U7691 (N_7691,N_6829,N_6537);
and U7692 (N_7692,N_6499,N_6080);
or U7693 (N_7693,N_6002,N_6637);
or U7694 (N_7694,N_6501,N_6022);
nor U7695 (N_7695,N_6011,N_6555);
nor U7696 (N_7696,N_6047,N_6093);
nand U7697 (N_7697,N_6032,N_6889);
and U7698 (N_7698,N_6599,N_6087);
and U7699 (N_7699,N_6338,N_6103);
nand U7700 (N_7700,N_6869,N_6851);
and U7701 (N_7701,N_6929,N_6057);
and U7702 (N_7702,N_6007,N_6167);
nor U7703 (N_7703,N_6300,N_6518);
nor U7704 (N_7704,N_6805,N_6282);
or U7705 (N_7705,N_6419,N_6840);
nand U7706 (N_7706,N_6075,N_6393);
nand U7707 (N_7707,N_6112,N_6296);
and U7708 (N_7708,N_6590,N_6878);
nor U7709 (N_7709,N_6643,N_6944);
and U7710 (N_7710,N_6299,N_6635);
and U7711 (N_7711,N_6380,N_6459);
or U7712 (N_7712,N_6919,N_6848);
or U7713 (N_7713,N_6678,N_6003);
nor U7714 (N_7714,N_6905,N_6867);
nor U7715 (N_7715,N_6859,N_6380);
and U7716 (N_7716,N_6697,N_6446);
nor U7717 (N_7717,N_6756,N_6264);
and U7718 (N_7718,N_6674,N_6171);
and U7719 (N_7719,N_6909,N_6971);
nor U7720 (N_7720,N_6645,N_6142);
nor U7721 (N_7721,N_6333,N_6218);
and U7722 (N_7722,N_6175,N_6265);
or U7723 (N_7723,N_6866,N_6359);
nand U7724 (N_7724,N_6780,N_6759);
nand U7725 (N_7725,N_6771,N_6297);
or U7726 (N_7726,N_6410,N_6070);
nor U7727 (N_7727,N_6542,N_6580);
nor U7728 (N_7728,N_6689,N_6962);
and U7729 (N_7729,N_6698,N_6733);
and U7730 (N_7730,N_6838,N_6252);
nor U7731 (N_7731,N_6262,N_6897);
or U7732 (N_7732,N_6937,N_6225);
nand U7733 (N_7733,N_6924,N_6054);
nor U7734 (N_7734,N_6991,N_6455);
nand U7735 (N_7735,N_6081,N_6598);
nor U7736 (N_7736,N_6818,N_6016);
nor U7737 (N_7737,N_6744,N_6784);
nor U7738 (N_7738,N_6469,N_6156);
and U7739 (N_7739,N_6673,N_6844);
and U7740 (N_7740,N_6118,N_6051);
and U7741 (N_7741,N_6634,N_6290);
nor U7742 (N_7742,N_6970,N_6463);
nor U7743 (N_7743,N_6083,N_6775);
nor U7744 (N_7744,N_6925,N_6265);
or U7745 (N_7745,N_6103,N_6925);
nand U7746 (N_7746,N_6897,N_6540);
or U7747 (N_7747,N_6563,N_6880);
or U7748 (N_7748,N_6581,N_6358);
or U7749 (N_7749,N_6901,N_6562);
or U7750 (N_7750,N_6865,N_6726);
nand U7751 (N_7751,N_6802,N_6561);
nand U7752 (N_7752,N_6036,N_6819);
or U7753 (N_7753,N_6859,N_6801);
and U7754 (N_7754,N_6015,N_6953);
and U7755 (N_7755,N_6179,N_6671);
or U7756 (N_7756,N_6595,N_6147);
nor U7757 (N_7757,N_6650,N_6800);
nand U7758 (N_7758,N_6415,N_6891);
nor U7759 (N_7759,N_6145,N_6196);
and U7760 (N_7760,N_6594,N_6907);
and U7761 (N_7761,N_6574,N_6348);
nand U7762 (N_7762,N_6816,N_6106);
nor U7763 (N_7763,N_6530,N_6142);
nand U7764 (N_7764,N_6160,N_6708);
and U7765 (N_7765,N_6434,N_6558);
and U7766 (N_7766,N_6294,N_6184);
and U7767 (N_7767,N_6340,N_6067);
or U7768 (N_7768,N_6072,N_6117);
or U7769 (N_7769,N_6955,N_6212);
or U7770 (N_7770,N_6529,N_6522);
nor U7771 (N_7771,N_6868,N_6993);
and U7772 (N_7772,N_6207,N_6777);
nor U7773 (N_7773,N_6385,N_6192);
xnor U7774 (N_7774,N_6547,N_6341);
and U7775 (N_7775,N_6652,N_6782);
nand U7776 (N_7776,N_6209,N_6901);
nor U7777 (N_7777,N_6935,N_6517);
nand U7778 (N_7778,N_6551,N_6283);
nor U7779 (N_7779,N_6665,N_6327);
nor U7780 (N_7780,N_6616,N_6649);
nor U7781 (N_7781,N_6363,N_6010);
nand U7782 (N_7782,N_6597,N_6382);
nor U7783 (N_7783,N_6899,N_6598);
or U7784 (N_7784,N_6323,N_6549);
and U7785 (N_7785,N_6072,N_6422);
nor U7786 (N_7786,N_6870,N_6675);
and U7787 (N_7787,N_6529,N_6312);
and U7788 (N_7788,N_6433,N_6471);
nor U7789 (N_7789,N_6078,N_6860);
and U7790 (N_7790,N_6149,N_6087);
or U7791 (N_7791,N_6341,N_6809);
nand U7792 (N_7792,N_6603,N_6613);
or U7793 (N_7793,N_6985,N_6895);
nand U7794 (N_7794,N_6795,N_6388);
nor U7795 (N_7795,N_6698,N_6116);
or U7796 (N_7796,N_6664,N_6429);
or U7797 (N_7797,N_6370,N_6203);
nor U7798 (N_7798,N_6556,N_6473);
nand U7799 (N_7799,N_6711,N_6691);
nand U7800 (N_7800,N_6372,N_6045);
and U7801 (N_7801,N_6285,N_6947);
or U7802 (N_7802,N_6963,N_6800);
nand U7803 (N_7803,N_6804,N_6655);
and U7804 (N_7804,N_6849,N_6721);
nand U7805 (N_7805,N_6401,N_6023);
or U7806 (N_7806,N_6905,N_6817);
nand U7807 (N_7807,N_6780,N_6471);
nand U7808 (N_7808,N_6341,N_6094);
nand U7809 (N_7809,N_6158,N_6879);
and U7810 (N_7810,N_6437,N_6013);
xnor U7811 (N_7811,N_6980,N_6233);
nand U7812 (N_7812,N_6777,N_6523);
nor U7813 (N_7813,N_6606,N_6264);
nand U7814 (N_7814,N_6465,N_6781);
or U7815 (N_7815,N_6381,N_6906);
or U7816 (N_7816,N_6393,N_6196);
nand U7817 (N_7817,N_6196,N_6118);
or U7818 (N_7818,N_6689,N_6084);
and U7819 (N_7819,N_6222,N_6649);
nor U7820 (N_7820,N_6739,N_6166);
nor U7821 (N_7821,N_6486,N_6586);
or U7822 (N_7822,N_6431,N_6180);
nand U7823 (N_7823,N_6134,N_6502);
and U7824 (N_7824,N_6388,N_6103);
nor U7825 (N_7825,N_6730,N_6892);
nand U7826 (N_7826,N_6486,N_6024);
nor U7827 (N_7827,N_6169,N_6033);
or U7828 (N_7828,N_6987,N_6758);
nand U7829 (N_7829,N_6869,N_6832);
and U7830 (N_7830,N_6341,N_6209);
nand U7831 (N_7831,N_6928,N_6917);
nand U7832 (N_7832,N_6760,N_6517);
nor U7833 (N_7833,N_6855,N_6402);
nor U7834 (N_7834,N_6706,N_6940);
nor U7835 (N_7835,N_6148,N_6390);
nand U7836 (N_7836,N_6725,N_6889);
nand U7837 (N_7837,N_6299,N_6347);
or U7838 (N_7838,N_6693,N_6726);
or U7839 (N_7839,N_6264,N_6184);
or U7840 (N_7840,N_6588,N_6717);
or U7841 (N_7841,N_6026,N_6464);
and U7842 (N_7842,N_6500,N_6799);
or U7843 (N_7843,N_6984,N_6086);
nor U7844 (N_7844,N_6031,N_6506);
and U7845 (N_7845,N_6106,N_6259);
nor U7846 (N_7846,N_6363,N_6445);
xor U7847 (N_7847,N_6916,N_6879);
and U7848 (N_7848,N_6562,N_6742);
xor U7849 (N_7849,N_6272,N_6297);
and U7850 (N_7850,N_6648,N_6155);
xor U7851 (N_7851,N_6094,N_6427);
nor U7852 (N_7852,N_6331,N_6209);
and U7853 (N_7853,N_6480,N_6891);
or U7854 (N_7854,N_6168,N_6683);
or U7855 (N_7855,N_6275,N_6430);
and U7856 (N_7856,N_6334,N_6074);
nand U7857 (N_7857,N_6862,N_6259);
nor U7858 (N_7858,N_6778,N_6684);
nor U7859 (N_7859,N_6292,N_6243);
nand U7860 (N_7860,N_6246,N_6281);
nand U7861 (N_7861,N_6470,N_6002);
and U7862 (N_7862,N_6654,N_6436);
or U7863 (N_7863,N_6461,N_6043);
nor U7864 (N_7864,N_6536,N_6031);
and U7865 (N_7865,N_6147,N_6620);
nand U7866 (N_7866,N_6910,N_6695);
or U7867 (N_7867,N_6730,N_6046);
nand U7868 (N_7868,N_6872,N_6302);
nand U7869 (N_7869,N_6614,N_6056);
nor U7870 (N_7870,N_6175,N_6159);
and U7871 (N_7871,N_6676,N_6581);
or U7872 (N_7872,N_6452,N_6770);
or U7873 (N_7873,N_6972,N_6577);
nand U7874 (N_7874,N_6168,N_6490);
nand U7875 (N_7875,N_6907,N_6607);
and U7876 (N_7876,N_6870,N_6619);
and U7877 (N_7877,N_6658,N_6872);
and U7878 (N_7878,N_6937,N_6899);
and U7879 (N_7879,N_6506,N_6682);
or U7880 (N_7880,N_6506,N_6640);
nor U7881 (N_7881,N_6039,N_6440);
and U7882 (N_7882,N_6241,N_6311);
and U7883 (N_7883,N_6725,N_6733);
nand U7884 (N_7884,N_6267,N_6709);
nand U7885 (N_7885,N_6305,N_6954);
nor U7886 (N_7886,N_6080,N_6500);
xor U7887 (N_7887,N_6325,N_6025);
or U7888 (N_7888,N_6643,N_6446);
xnor U7889 (N_7889,N_6033,N_6817);
nor U7890 (N_7890,N_6846,N_6393);
nand U7891 (N_7891,N_6430,N_6797);
xnor U7892 (N_7892,N_6251,N_6601);
nor U7893 (N_7893,N_6591,N_6985);
and U7894 (N_7894,N_6141,N_6521);
nand U7895 (N_7895,N_6236,N_6012);
or U7896 (N_7896,N_6700,N_6447);
nor U7897 (N_7897,N_6821,N_6984);
nor U7898 (N_7898,N_6780,N_6370);
and U7899 (N_7899,N_6833,N_6195);
nor U7900 (N_7900,N_6786,N_6844);
and U7901 (N_7901,N_6812,N_6723);
or U7902 (N_7902,N_6607,N_6200);
and U7903 (N_7903,N_6013,N_6277);
or U7904 (N_7904,N_6874,N_6611);
and U7905 (N_7905,N_6369,N_6803);
nand U7906 (N_7906,N_6515,N_6491);
or U7907 (N_7907,N_6868,N_6890);
nor U7908 (N_7908,N_6038,N_6873);
nand U7909 (N_7909,N_6722,N_6186);
nor U7910 (N_7910,N_6754,N_6077);
nand U7911 (N_7911,N_6665,N_6709);
nand U7912 (N_7912,N_6258,N_6949);
nand U7913 (N_7913,N_6968,N_6582);
nand U7914 (N_7914,N_6362,N_6335);
nor U7915 (N_7915,N_6233,N_6656);
nand U7916 (N_7916,N_6615,N_6731);
nor U7917 (N_7917,N_6943,N_6884);
nor U7918 (N_7918,N_6810,N_6406);
or U7919 (N_7919,N_6073,N_6022);
nand U7920 (N_7920,N_6551,N_6705);
or U7921 (N_7921,N_6805,N_6003);
nand U7922 (N_7922,N_6185,N_6017);
or U7923 (N_7923,N_6685,N_6526);
and U7924 (N_7924,N_6507,N_6764);
or U7925 (N_7925,N_6538,N_6212);
or U7926 (N_7926,N_6212,N_6339);
nor U7927 (N_7927,N_6647,N_6893);
and U7928 (N_7928,N_6829,N_6495);
or U7929 (N_7929,N_6520,N_6559);
and U7930 (N_7930,N_6813,N_6944);
nand U7931 (N_7931,N_6847,N_6670);
nor U7932 (N_7932,N_6024,N_6881);
nand U7933 (N_7933,N_6940,N_6392);
nor U7934 (N_7934,N_6953,N_6288);
nand U7935 (N_7935,N_6119,N_6770);
nor U7936 (N_7936,N_6311,N_6724);
nor U7937 (N_7937,N_6294,N_6832);
nor U7938 (N_7938,N_6686,N_6967);
nor U7939 (N_7939,N_6253,N_6323);
nor U7940 (N_7940,N_6684,N_6068);
nor U7941 (N_7941,N_6268,N_6478);
and U7942 (N_7942,N_6330,N_6522);
and U7943 (N_7943,N_6532,N_6815);
and U7944 (N_7944,N_6903,N_6723);
nand U7945 (N_7945,N_6166,N_6870);
and U7946 (N_7946,N_6331,N_6477);
and U7947 (N_7947,N_6202,N_6751);
or U7948 (N_7948,N_6050,N_6972);
nand U7949 (N_7949,N_6703,N_6959);
and U7950 (N_7950,N_6597,N_6093);
or U7951 (N_7951,N_6560,N_6341);
or U7952 (N_7952,N_6987,N_6834);
or U7953 (N_7953,N_6159,N_6692);
nor U7954 (N_7954,N_6929,N_6210);
and U7955 (N_7955,N_6390,N_6772);
and U7956 (N_7956,N_6008,N_6335);
nand U7957 (N_7957,N_6963,N_6763);
nor U7958 (N_7958,N_6562,N_6762);
and U7959 (N_7959,N_6553,N_6908);
and U7960 (N_7960,N_6479,N_6673);
or U7961 (N_7961,N_6941,N_6969);
nor U7962 (N_7962,N_6932,N_6810);
or U7963 (N_7963,N_6201,N_6379);
nor U7964 (N_7964,N_6995,N_6237);
nand U7965 (N_7965,N_6560,N_6230);
or U7966 (N_7966,N_6875,N_6803);
nor U7967 (N_7967,N_6079,N_6769);
nor U7968 (N_7968,N_6735,N_6553);
nand U7969 (N_7969,N_6651,N_6971);
or U7970 (N_7970,N_6197,N_6026);
nand U7971 (N_7971,N_6005,N_6762);
nand U7972 (N_7972,N_6141,N_6933);
nand U7973 (N_7973,N_6313,N_6394);
and U7974 (N_7974,N_6096,N_6310);
and U7975 (N_7975,N_6446,N_6699);
and U7976 (N_7976,N_6229,N_6721);
nor U7977 (N_7977,N_6722,N_6094);
nor U7978 (N_7978,N_6031,N_6097);
nor U7979 (N_7979,N_6247,N_6095);
nand U7980 (N_7980,N_6563,N_6523);
nor U7981 (N_7981,N_6139,N_6936);
nand U7982 (N_7982,N_6107,N_6878);
and U7983 (N_7983,N_6921,N_6329);
and U7984 (N_7984,N_6619,N_6657);
and U7985 (N_7985,N_6205,N_6615);
and U7986 (N_7986,N_6035,N_6281);
nor U7987 (N_7987,N_6529,N_6095);
nand U7988 (N_7988,N_6378,N_6825);
or U7989 (N_7989,N_6800,N_6709);
nand U7990 (N_7990,N_6627,N_6452);
nand U7991 (N_7991,N_6254,N_6668);
or U7992 (N_7992,N_6914,N_6325);
nand U7993 (N_7993,N_6527,N_6578);
nand U7994 (N_7994,N_6942,N_6784);
and U7995 (N_7995,N_6610,N_6850);
or U7996 (N_7996,N_6605,N_6344);
nor U7997 (N_7997,N_6793,N_6673);
and U7998 (N_7998,N_6305,N_6048);
nand U7999 (N_7999,N_6516,N_6665);
nor U8000 (N_8000,N_7942,N_7747);
or U8001 (N_8001,N_7446,N_7201);
and U8002 (N_8002,N_7171,N_7908);
nand U8003 (N_8003,N_7289,N_7903);
and U8004 (N_8004,N_7495,N_7477);
and U8005 (N_8005,N_7025,N_7348);
nor U8006 (N_8006,N_7836,N_7399);
nand U8007 (N_8007,N_7503,N_7368);
or U8008 (N_8008,N_7770,N_7126);
nor U8009 (N_8009,N_7292,N_7657);
or U8010 (N_8010,N_7390,N_7211);
and U8011 (N_8011,N_7443,N_7785);
and U8012 (N_8012,N_7296,N_7595);
or U8013 (N_8013,N_7373,N_7112);
and U8014 (N_8014,N_7269,N_7920);
or U8015 (N_8015,N_7653,N_7267);
nor U8016 (N_8016,N_7034,N_7569);
nand U8017 (N_8017,N_7682,N_7170);
nor U8018 (N_8018,N_7969,N_7887);
and U8019 (N_8019,N_7979,N_7258);
nand U8020 (N_8020,N_7337,N_7691);
or U8021 (N_8021,N_7582,N_7635);
nor U8022 (N_8022,N_7119,N_7820);
nand U8023 (N_8023,N_7197,N_7251);
nand U8024 (N_8024,N_7430,N_7765);
or U8025 (N_8025,N_7159,N_7917);
nor U8026 (N_8026,N_7147,N_7150);
or U8027 (N_8027,N_7875,N_7353);
nor U8028 (N_8028,N_7364,N_7350);
nor U8029 (N_8029,N_7087,N_7900);
or U8030 (N_8030,N_7693,N_7593);
nand U8031 (N_8031,N_7476,N_7506);
nand U8032 (N_8032,N_7907,N_7591);
and U8033 (N_8033,N_7952,N_7273);
and U8034 (N_8034,N_7579,N_7583);
and U8035 (N_8035,N_7946,N_7091);
or U8036 (N_8036,N_7805,N_7723);
or U8037 (N_8037,N_7066,N_7220);
nand U8038 (N_8038,N_7950,N_7982);
nand U8039 (N_8039,N_7391,N_7388);
and U8040 (N_8040,N_7330,N_7431);
or U8041 (N_8041,N_7148,N_7143);
and U8042 (N_8042,N_7849,N_7530);
nor U8043 (N_8043,N_7237,N_7652);
and U8044 (N_8044,N_7687,N_7871);
nor U8045 (N_8045,N_7400,N_7181);
nand U8046 (N_8046,N_7796,N_7169);
nor U8047 (N_8047,N_7560,N_7006);
and U8048 (N_8048,N_7293,N_7363);
or U8049 (N_8049,N_7432,N_7023);
or U8050 (N_8050,N_7800,N_7161);
or U8051 (N_8051,N_7762,N_7242);
or U8052 (N_8052,N_7462,N_7733);
nor U8053 (N_8053,N_7921,N_7288);
nand U8054 (N_8054,N_7297,N_7054);
and U8055 (N_8055,N_7598,N_7532);
nand U8056 (N_8056,N_7214,N_7085);
nand U8057 (N_8057,N_7614,N_7199);
nor U8058 (N_8058,N_7017,N_7885);
or U8059 (N_8059,N_7440,N_7830);
or U8060 (N_8060,N_7478,N_7854);
or U8061 (N_8061,N_7571,N_7387);
or U8062 (N_8062,N_7175,N_7375);
nor U8063 (N_8063,N_7649,N_7114);
and U8064 (N_8064,N_7457,N_7332);
nor U8065 (N_8065,N_7870,N_7265);
nor U8066 (N_8066,N_7922,N_7374);
nand U8067 (N_8067,N_7749,N_7082);
nor U8068 (N_8068,N_7507,N_7782);
nand U8069 (N_8069,N_7702,N_7542);
nand U8070 (N_8070,N_7151,N_7597);
nor U8071 (N_8071,N_7480,N_7426);
and U8072 (N_8072,N_7659,N_7514);
and U8073 (N_8073,N_7642,N_7596);
or U8074 (N_8074,N_7958,N_7323);
nor U8075 (N_8075,N_7102,N_7370);
and U8076 (N_8076,N_7822,N_7898);
or U8077 (N_8077,N_7221,N_7472);
and U8078 (N_8078,N_7680,N_7538);
or U8079 (N_8079,N_7835,N_7972);
and U8080 (N_8080,N_7763,N_7484);
or U8081 (N_8081,N_7573,N_7741);
nor U8082 (N_8082,N_7526,N_7511);
nor U8083 (N_8083,N_7919,N_7909);
nand U8084 (N_8084,N_7306,N_7318);
nand U8085 (N_8085,N_7581,N_7933);
and U8086 (N_8086,N_7456,N_7492);
nor U8087 (N_8087,N_7256,N_7036);
or U8088 (N_8088,N_7302,N_7743);
and U8089 (N_8089,N_7939,N_7962);
nor U8090 (N_8090,N_7473,N_7890);
or U8091 (N_8091,N_7234,N_7717);
nor U8092 (N_8092,N_7157,N_7825);
and U8093 (N_8093,N_7663,N_7522);
or U8094 (N_8094,N_7383,N_7678);
and U8095 (N_8095,N_7137,N_7812);
and U8096 (N_8096,N_7019,N_7216);
nand U8097 (N_8097,N_7708,N_7022);
nand U8098 (N_8098,N_7696,N_7915);
nand U8099 (N_8099,N_7385,N_7524);
nand U8100 (N_8100,N_7018,N_7868);
nor U8101 (N_8101,N_7622,N_7344);
and U8102 (N_8102,N_7677,N_7549);
nand U8103 (N_8103,N_7556,N_7180);
nand U8104 (N_8104,N_7300,N_7746);
xor U8105 (N_8105,N_7978,N_7660);
nor U8106 (N_8106,N_7423,N_7807);
nor U8107 (N_8107,N_7365,N_7925);
and U8108 (N_8108,N_7008,N_7924);
and U8109 (N_8109,N_7224,N_7779);
nor U8110 (N_8110,N_7421,N_7931);
nand U8111 (N_8111,N_7817,N_7059);
or U8112 (N_8112,N_7738,N_7889);
nor U8113 (N_8113,N_7543,N_7517);
nor U8114 (N_8114,N_7638,N_7609);
and U8115 (N_8115,N_7799,N_7294);
nor U8116 (N_8116,N_7343,N_7947);
nor U8117 (N_8117,N_7673,N_7283);
nor U8118 (N_8118,N_7094,N_7389);
or U8119 (N_8119,N_7627,N_7794);
nand U8120 (N_8120,N_7861,N_7498);
or U8121 (N_8121,N_7122,N_7475);
nor U8122 (N_8122,N_7975,N_7155);
or U8123 (N_8123,N_7450,N_7670);
nand U8124 (N_8124,N_7067,N_7239);
nor U8125 (N_8125,N_7781,N_7840);
nor U8126 (N_8126,N_7222,N_7675);
or U8127 (N_8127,N_7434,N_7341);
and U8128 (N_8128,N_7316,N_7177);
or U8129 (N_8129,N_7461,N_7049);
and U8130 (N_8130,N_7883,N_7255);
xor U8131 (N_8131,N_7864,N_7172);
nand U8132 (N_8132,N_7166,N_7356);
nor U8133 (N_8133,N_7880,N_7173);
nand U8134 (N_8134,N_7668,N_7729);
and U8135 (N_8135,N_7482,N_7270);
or U8136 (N_8136,N_7720,N_7879);
and U8137 (N_8137,N_7860,N_7937);
nor U8138 (N_8138,N_7202,N_7757);
and U8139 (N_8139,N_7774,N_7641);
nand U8140 (N_8140,N_7905,N_7715);
nand U8141 (N_8141,N_7756,N_7001);
and U8142 (N_8142,N_7020,N_7710);
nand U8143 (N_8143,N_7415,N_7116);
or U8144 (N_8144,N_7485,N_7096);
nor U8145 (N_8145,N_7966,N_7540);
nand U8146 (N_8146,N_7955,N_7136);
or U8147 (N_8147,N_7661,N_7600);
and U8148 (N_8148,N_7286,N_7531);
nand U8149 (N_8149,N_7088,N_7613);
and U8150 (N_8150,N_7516,N_7384);
nand U8151 (N_8151,N_7829,N_7298);
or U8152 (N_8152,N_7405,N_7455);
nor U8153 (N_8153,N_7030,N_7077);
or U8154 (N_8154,N_7312,N_7204);
nand U8155 (N_8155,N_7011,N_7235);
or U8156 (N_8156,N_7704,N_7973);
and U8157 (N_8157,N_7328,N_7632);
and U8158 (N_8158,N_7865,N_7686);
and U8159 (N_8159,N_7260,N_7699);
and U8160 (N_8160,N_7381,N_7407);
nand U8161 (N_8161,N_7287,N_7402);
nand U8162 (N_8162,N_7414,N_7518);
nand U8163 (N_8163,N_7760,N_7912);
and U8164 (N_8164,N_7099,N_7940);
and U8165 (N_8165,N_7831,N_7301);
and U8166 (N_8166,N_7737,N_7338);
and U8167 (N_8167,N_7427,N_7636);
and U8168 (N_8168,N_7187,N_7508);
and U8169 (N_8169,N_7576,N_7916);
and U8170 (N_8170,N_7182,N_7123);
or U8171 (N_8171,N_7489,N_7113);
nor U8172 (N_8172,N_7333,N_7718);
nor U8173 (N_8173,N_7320,N_7240);
or U8174 (N_8174,N_7953,N_7167);
xor U8175 (N_8175,N_7186,N_7821);
nor U8176 (N_8176,N_7643,N_7156);
and U8177 (N_8177,N_7824,N_7797);
and U8178 (N_8178,N_7499,N_7163);
or U8179 (N_8179,N_7442,N_7042);
nand U8180 (N_8180,N_7910,N_7968);
and U8181 (N_8181,N_7097,N_7366);
or U8182 (N_8182,N_7335,N_7184);
and U8183 (N_8183,N_7090,N_7138);
nand U8184 (N_8184,N_7347,N_7327);
or U8185 (N_8185,N_7873,N_7153);
and U8186 (N_8186,N_7238,N_7935);
or U8187 (N_8187,N_7881,N_7567);
nor U8188 (N_8188,N_7494,N_7559);
and U8189 (N_8189,N_7810,N_7304);
nor U8190 (N_8190,N_7386,N_7192);
or U8191 (N_8191,N_7669,N_7681);
and U8192 (N_8192,N_7447,N_7895);
or U8193 (N_8193,N_7888,N_7439);
nand U8194 (N_8194,N_7002,N_7313);
and U8195 (N_8195,N_7231,N_7533);
nand U8196 (N_8196,N_7321,N_7727);
nand U8197 (N_8197,N_7466,N_7874);
and U8198 (N_8198,N_7984,N_7249);
and U8199 (N_8199,N_7406,N_7869);
nor U8200 (N_8200,N_7392,N_7515);
or U8201 (N_8201,N_7795,N_7108);
or U8202 (N_8202,N_7281,N_7610);
nor U8203 (N_8203,N_7951,N_7878);
nand U8204 (N_8204,N_7588,N_7227);
nor U8205 (N_8205,N_7215,N_7261);
nand U8206 (N_8206,N_7205,N_7026);
nor U8207 (N_8207,N_7814,N_7844);
and U8208 (N_8208,N_7809,N_7314);
and U8209 (N_8209,N_7934,N_7904);
xor U8210 (N_8210,N_7397,N_7587);
or U8211 (N_8211,N_7778,N_7486);
nand U8212 (N_8212,N_7488,N_7007);
nor U8213 (N_8213,N_7118,N_7396);
and U8214 (N_8214,N_7133,N_7010);
nor U8215 (N_8215,N_7291,N_7546);
or U8216 (N_8216,N_7943,N_7505);
and U8217 (N_8217,N_7213,N_7086);
nor U8218 (N_8218,N_7563,N_7395);
or U8219 (N_8219,N_7529,N_7101);
or U8220 (N_8220,N_7124,N_7109);
nor U8221 (N_8221,N_7945,N_7453);
and U8222 (N_8222,N_7590,N_7711);
or U8223 (N_8223,N_7759,N_7063);
nand U8224 (N_8224,N_7057,N_7902);
or U8225 (N_8225,N_7481,N_7911);
and U8226 (N_8226,N_7777,N_7761);
and U8227 (N_8227,N_7217,N_7401);
nor U8228 (N_8228,N_7073,N_7823);
or U8229 (N_8229,N_7557,N_7554);
and U8230 (N_8230,N_7575,N_7896);
or U8231 (N_8231,N_7244,N_7051);
nand U8232 (N_8232,N_7523,N_7120);
and U8233 (N_8233,N_7015,N_7574);
nor U8234 (N_8234,N_7626,N_7944);
nor U8235 (N_8235,N_7142,N_7683);
and U8236 (N_8236,N_7012,N_7206);
nand U8237 (N_8237,N_7245,N_7535);
nor U8238 (N_8238,N_7470,N_7806);
or U8239 (N_8239,N_7319,N_7061);
nand U8240 (N_8240,N_7110,N_7758);
and U8241 (N_8241,N_7928,N_7630);
nor U8242 (N_8242,N_7802,N_7263);
or U8243 (N_8243,N_7801,N_7418);
nand U8244 (N_8244,N_7619,N_7419);
and U8245 (N_8245,N_7991,N_7655);
and U8246 (N_8246,N_7913,N_7158);
or U8247 (N_8247,N_7241,N_7954);
or U8248 (N_8248,N_7404,N_7454);
nand U8249 (N_8249,N_7230,N_7726);
nand U8250 (N_8250,N_7923,N_7268);
or U8251 (N_8251,N_7724,N_7274);
or U8252 (N_8252,N_7060,N_7901);
or U8253 (N_8253,N_7311,N_7621);
or U8254 (N_8254,N_7956,N_7491);
nand U8255 (N_8255,N_7229,N_7735);
and U8256 (N_8256,N_7436,N_7376);
nand U8257 (N_8257,N_7100,N_7845);
nand U8258 (N_8258,N_7617,N_7056);
and U8259 (N_8259,N_7149,N_7891);
or U8260 (N_8260,N_7496,N_7474);
nand U8261 (N_8261,N_7279,N_7985);
and U8262 (N_8262,N_7132,N_7803);
and U8263 (N_8263,N_7135,N_7160);
and U8264 (N_8264,N_7594,N_7633);
and U8265 (N_8265,N_7513,N_7409);
nor U8266 (N_8266,N_7764,N_7618);
xor U8267 (N_8267,N_7317,N_7751);
nor U8268 (N_8268,N_7393,N_7694);
and U8269 (N_8269,N_7716,N_7334);
nand U8270 (N_8270,N_7451,N_7872);
or U8271 (N_8271,N_7045,N_7125);
and U8272 (N_8272,N_7278,N_7188);
and U8273 (N_8273,N_7629,N_7536);
and U8274 (N_8274,N_7558,N_7016);
and U8275 (N_8275,N_7929,N_7534);
nand U8276 (N_8276,N_7483,N_7713);
nor U8277 (N_8277,N_7949,N_7121);
and U8278 (N_8278,N_7562,N_7497);
nand U8279 (N_8279,N_7859,N_7808);
nand U8280 (N_8280,N_7640,N_7083);
and U8281 (N_8281,N_7500,N_7103);
nand U8282 (N_8282,N_7129,N_7326);
and U8283 (N_8283,N_7191,N_7858);
nand U8284 (N_8284,N_7918,N_7468);
and U8285 (N_8285,N_7264,N_7052);
and U8286 (N_8286,N_7307,N_7698);
nor U8287 (N_8287,N_7464,N_7744);
nor U8288 (N_8288,N_7165,N_7745);
and U8289 (N_8289,N_7703,N_7606);
or U8290 (N_8290,N_7882,N_7280);
nor U8291 (N_8291,N_7225,N_7832);
nand U8292 (N_8292,N_7359,N_7413);
nand U8293 (N_8293,N_7420,N_7780);
or U8294 (N_8294,N_7422,N_7974);
nand U8295 (N_8295,N_7322,N_7079);
and U8296 (N_8296,N_7989,N_7380);
or U8297 (N_8297,N_7203,N_7656);
nor U8298 (N_8298,N_7566,N_7959);
and U8299 (N_8299,N_7044,N_7183);
nor U8300 (N_8300,N_7266,N_7117);
nand U8301 (N_8301,N_7843,N_7047);
and U8302 (N_8302,N_7021,N_7324);
and U8303 (N_8303,N_7009,N_7838);
and U8304 (N_8304,N_7226,N_7032);
nor U8305 (N_8305,N_7459,N_7128);
nand U8306 (N_8306,N_7578,N_7601);
nand U8307 (N_8307,N_7866,N_7752);
or U8308 (N_8308,N_7964,N_7075);
nor U8309 (N_8309,N_7185,N_7602);
and U8310 (N_8310,N_7813,N_7971);
nand U8311 (N_8311,N_7377,N_7539);
or U8312 (N_8312,N_7040,N_7349);
and U8313 (N_8313,N_7644,N_7361);
or U8314 (N_8314,N_7469,N_7977);
and U8315 (N_8315,N_7804,N_7193);
nor U8316 (N_8316,N_7379,N_7035);
nand U8317 (N_8317,N_7164,N_7444);
or U8318 (N_8318,N_7519,N_7767);
and U8319 (N_8319,N_7646,N_7707);
nor U8320 (N_8320,N_7709,N_7253);
nor U8321 (N_8321,N_7998,N_7043);
xor U8322 (N_8322,N_7425,N_7967);
and U8323 (N_8323,N_7196,N_7509);
and U8324 (N_8324,N_7254,N_7345);
nor U8325 (N_8325,N_7714,N_7676);
nor U8326 (N_8326,N_7080,N_7788);
nand U8327 (N_8327,N_7223,N_7634);
or U8328 (N_8328,N_7541,N_7104);
or U8329 (N_8329,N_7846,N_7190);
nor U8330 (N_8330,N_7248,N_7605);
nand U8331 (N_8331,N_7862,N_7748);
nand U8332 (N_8332,N_7957,N_7250);
nor U8333 (N_8333,N_7003,N_7892);
nand U8334 (N_8334,N_7354,N_7771);
and U8335 (N_8335,N_7058,N_7271);
nor U8336 (N_8336,N_7564,N_7134);
xor U8337 (N_8337,N_7055,N_7987);
nor U8338 (N_8338,N_7416,N_7815);
or U8339 (N_8339,N_7631,N_7818);
nor U8340 (N_8340,N_7467,N_7315);
nor U8341 (N_8341,N_7679,N_7997);
and U8342 (N_8342,N_7705,N_7072);
nand U8343 (N_8343,N_7435,N_7827);
and U8344 (N_8344,N_7521,N_7154);
or U8345 (N_8345,N_7654,N_7773);
or U8346 (N_8346,N_7510,N_7791);
and U8347 (N_8347,N_7645,N_7615);
nand U8348 (N_8348,N_7233,N_7198);
or U8349 (N_8349,N_7200,N_7792);
nand U8350 (N_8350,N_7550,N_7152);
nor U8351 (N_8351,N_7570,N_7360);
nor U8352 (N_8352,N_7352,N_7284);
nor U8353 (N_8353,N_7127,N_7178);
nor U8354 (N_8354,N_7275,N_7501);
or U8355 (N_8355,N_7078,N_7616);
nand U8356 (N_8356,N_7232,N_7603);
nor U8357 (N_8357,N_7826,N_7168);
nand U8358 (N_8358,N_7029,N_7856);
nand U8359 (N_8359,N_7144,N_7853);
or U8360 (N_8360,N_7033,N_7357);
nand U8361 (N_8361,N_7146,N_7936);
nand U8362 (N_8362,N_7789,N_7775);
or U8363 (N_8363,N_7876,N_7448);
or U8364 (N_8364,N_7076,N_7811);
and U8365 (N_8365,N_7340,N_7276);
nor U8366 (N_8366,N_7068,N_7850);
nand U8367 (N_8367,N_7722,N_7662);
nand U8368 (N_8368,N_7027,N_7624);
and U8369 (N_8369,N_7719,N_7394);
and U8370 (N_8370,N_7189,N_7458);
or U8371 (N_8371,N_7065,N_7048);
and U8372 (N_8372,N_7695,N_7650);
nor U8373 (N_8373,N_7428,N_7069);
nand U8374 (N_8374,N_7179,N_7651);
and U8375 (N_8375,N_7639,N_7512);
and U8376 (N_8376,N_7612,N_7867);
nand U8377 (N_8377,N_7105,N_7408);
or U8378 (N_8378,N_7410,N_7842);
nand U8379 (N_8379,N_7666,N_7339);
nand U8380 (N_8380,N_7684,N_7995);
or U8381 (N_8381,N_7463,N_7648);
or U8382 (N_8382,N_7355,N_7628);
and U8383 (N_8383,N_7926,N_7894);
and U8384 (N_8384,N_7252,N_7433);
nor U8385 (N_8385,N_7692,N_7784);
and U8386 (N_8386,N_7941,N_7766);
and U8387 (N_8387,N_7028,N_7742);
or U8388 (N_8388,N_7981,N_7262);
nand U8389 (N_8389,N_7980,N_7031);
nand U8390 (N_8390,N_7247,N_7604);
nand U8391 (N_8391,N_7671,N_7857);
and U8392 (N_8392,N_7552,N_7378);
nand U8393 (N_8393,N_7664,N_7372);
or U8394 (N_8394,N_7194,N_7310);
nor U8395 (N_8395,N_7014,N_7721);
nor U8396 (N_8396,N_7115,N_7828);
or U8397 (N_8397,N_7607,N_7740);
and U8398 (N_8398,N_7282,N_7371);
or U8399 (N_8399,N_7647,N_7299);
nand U8400 (N_8400,N_7837,N_7728);
nor U8401 (N_8401,N_7927,N_7932);
or U8402 (N_8402,N_7024,N_7062);
and U8403 (N_8403,N_7996,N_7081);
or U8404 (N_8404,N_7712,N_7039);
nor U8405 (N_8405,N_7106,N_7561);
xor U8406 (N_8406,N_7527,N_7986);
nor U8407 (N_8407,N_7819,N_7970);
or U8408 (N_8408,N_7471,N_7685);
nand U8409 (N_8409,N_7930,N_7608);
nand U8410 (N_8410,N_7688,N_7502);
or U8411 (N_8411,N_7309,N_7976);
and U8412 (N_8412,N_7768,N_7212);
nand U8413 (N_8413,N_7382,N_7863);
nor U8414 (N_8414,N_7290,N_7325);
or U8415 (N_8415,N_7487,N_7111);
nor U8416 (N_8416,N_7772,N_7331);
nor U8417 (N_8417,N_7739,N_7877);
and U8418 (N_8418,N_7417,N_7786);
and U8419 (N_8419,N_7336,N_7623);
nand U8420 (N_8420,N_7305,N_7725);
nand U8421 (N_8421,N_7839,N_7246);
or U8422 (N_8422,N_7732,N_7565);
nand U8423 (N_8423,N_7412,N_7460);
and U8424 (N_8424,N_7548,N_7585);
or U8425 (N_8425,N_7914,N_7897);
or U8426 (N_8426,N_7207,N_7537);
and U8427 (N_8427,N_7107,N_7445);
nor U8428 (N_8428,N_7074,N_7665);
nand U8429 (N_8429,N_7787,N_7938);
or U8430 (N_8430,N_7092,N_7611);
nand U8431 (N_8431,N_7769,N_7369);
nand U8432 (N_8432,N_7139,N_7285);
and U8433 (N_8433,N_7449,N_7362);
and U8434 (N_8434,N_7961,N_7783);
nand U8435 (N_8435,N_7790,N_7130);
nand U8436 (N_8436,N_7730,N_7131);
nor U8437 (N_8437,N_7753,N_7899);
and U8438 (N_8438,N_7493,N_7572);
or U8439 (N_8439,N_7544,N_7992);
nand U8440 (N_8440,N_7963,N_7658);
nor U8441 (N_8441,N_7064,N_7555);
and U8442 (N_8442,N_7351,N_7793);
or U8443 (N_8443,N_7236,N_7553);
nand U8444 (N_8444,N_7037,N_7734);
or U8445 (N_8445,N_7990,N_7580);
nand U8446 (N_8446,N_7303,N_7993);
nand U8447 (N_8447,N_7525,N_7438);
or U8448 (N_8448,N_7424,N_7520);
and U8449 (N_8449,N_7545,N_7620);
nor U8450 (N_8450,N_7174,N_7403);
or U8451 (N_8451,N_7209,N_7637);
nor U8452 (N_8452,N_7367,N_7329);
nand U8453 (N_8453,N_7141,N_7568);
or U8454 (N_8454,N_7833,N_7690);
nand U8455 (N_8455,N_7893,N_7441);
nor U8456 (N_8456,N_7437,N_7208);
nand U8457 (N_8457,N_7219,N_7071);
and U8458 (N_8458,N_7776,N_7041);
and U8459 (N_8459,N_7667,N_7672);
nor U8460 (N_8460,N_7697,N_7195);
and U8461 (N_8461,N_7960,N_7346);
nand U8462 (N_8462,N_7834,N_7851);
nand U8463 (N_8463,N_7852,N_7093);
nor U8464 (N_8464,N_7272,N_7140);
nor U8465 (N_8465,N_7295,N_7479);
or U8466 (N_8466,N_7465,N_7855);
nor U8467 (N_8467,N_7398,N_7988);
or U8468 (N_8468,N_7050,N_7625);
nand U8469 (N_8469,N_7218,N_7504);
nand U8470 (N_8470,N_7816,N_7528);
and U8471 (N_8471,N_7089,N_7731);
and U8472 (N_8472,N_7886,N_7070);
nor U8473 (N_8473,N_7259,N_7848);
and U8474 (N_8474,N_7999,N_7906);
and U8475 (N_8475,N_7228,N_7750);
nand U8476 (N_8476,N_7586,N_7095);
and U8477 (N_8477,N_7551,N_7965);
or U8478 (N_8478,N_7162,N_7674);
nand U8479 (N_8479,N_7342,N_7053);
nor U8480 (N_8480,N_7210,N_7592);
nor U8481 (N_8481,N_7046,N_7755);
and U8482 (N_8482,N_7038,N_7706);
nand U8483 (N_8483,N_7994,N_7005);
or U8484 (N_8484,N_7847,N_7013);
nor U8485 (N_8485,N_7701,N_7584);
nand U8486 (N_8486,N_7798,N_7490);
nand U8487 (N_8487,N_7983,N_7841);
nand U8488 (N_8488,N_7145,N_7577);
and U8489 (N_8489,N_7084,N_7736);
or U8490 (N_8490,N_7948,N_7000);
or U8491 (N_8491,N_7176,N_7277);
nor U8492 (N_8492,N_7754,N_7308);
nor U8493 (N_8493,N_7884,N_7429);
and U8494 (N_8494,N_7243,N_7589);
nand U8495 (N_8495,N_7599,N_7547);
nor U8496 (N_8496,N_7358,N_7700);
and U8497 (N_8497,N_7004,N_7452);
nor U8498 (N_8498,N_7411,N_7098);
or U8499 (N_8499,N_7689,N_7257);
nor U8500 (N_8500,N_7184,N_7154);
or U8501 (N_8501,N_7485,N_7314);
nor U8502 (N_8502,N_7493,N_7802);
nor U8503 (N_8503,N_7118,N_7078);
nor U8504 (N_8504,N_7702,N_7796);
or U8505 (N_8505,N_7220,N_7041);
or U8506 (N_8506,N_7627,N_7114);
and U8507 (N_8507,N_7919,N_7585);
or U8508 (N_8508,N_7280,N_7572);
and U8509 (N_8509,N_7326,N_7102);
nor U8510 (N_8510,N_7854,N_7114);
nand U8511 (N_8511,N_7440,N_7221);
and U8512 (N_8512,N_7298,N_7814);
or U8513 (N_8513,N_7440,N_7588);
nand U8514 (N_8514,N_7233,N_7343);
nor U8515 (N_8515,N_7341,N_7679);
nor U8516 (N_8516,N_7872,N_7437);
nand U8517 (N_8517,N_7737,N_7950);
nor U8518 (N_8518,N_7219,N_7337);
nor U8519 (N_8519,N_7685,N_7614);
and U8520 (N_8520,N_7772,N_7348);
nor U8521 (N_8521,N_7387,N_7155);
nand U8522 (N_8522,N_7918,N_7501);
and U8523 (N_8523,N_7785,N_7159);
nor U8524 (N_8524,N_7305,N_7860);
and U8525 (N_8525,N_7999,N_7508);
or U8526 (N_8526,N_7494,N_7349);
nand U8527 (N_8527,N_7390,N_7281);
nand U8528 (N_8528,N_7996,N_7809);
nor U8529 (N_8529,N_7710,N_7708);
nor U8530 (N_8530,N_7487,N_7190);
or U8531 (N_8531,N_7676,N_7464);
nand U8532 (N_8532,N_7055,N_7498);
nand U8533 (N_8533,N_7017,N_7820);
and U8534 (N_8534,N_7820,N_7729);
nor U8535 (N_8535,N_7146,N_7859);
and U8536 (N_8536,N_7707,N_7444);
nand U8537 (N_8537,N_7272,N_7524);
xor U8538 (N_8538,N_7395,N_7941);
or U8539 (N_8539,N_7001,N_7971);
or U8540 (N_8540,N_7296,N_7801);
nor U8541 (N_8541,N_7068,N_7300);
nand U8542 (N_8542,N_7138,N_7589);
or U8543 (N_8543,N_7946,N_7196);
and U8544 (N_8544,N_7486,N_7608);
nand U8545 (N_8545,N_7665,N_7566);
or U8546 (N_8546,N_7955,N_7487);
nor U8547 (N_8547,N_7996,N_7675);
nand U8548 (N_8548,N_7028,N_7483);
nor U8549 (N_8549,N_7961,N_7853);
nand U8550 (N_8550,N_7465,N_7354);
nand U8551 (N_8551,N_7328,N_7146);
nor U8552 (N_8552,N_7272,N_7692);
or U8553 (N_8553,N_7792,N_7915);
and U8554 (N_8554,N_7079,N_7137);
or U8555 (N_8555,N_7975,N_7282);
nand U8556 (N_8556,N_7590,N_7660);
nand U8557 (N_8557,N_7431,N_7233);
or U8558 (N_8558,N_7989,N_7792);
and U8559 (N_8559,N_7645,N_7260);
or U8560 (N_8560,N_7240,N_7420);
and U8561 (N_8561,N_7474,N_7125);
and U8562 (N_8562,N_7604,N_7877);
nor U8563 (N_8563,N_7618,N_7645);
nor U8564 (N_8564,N_7736,N_7874);
nor U8565 (N_8565,N_7055,N_7596);
or U8566 (N_8566,N_7999,N_7919);
nor U8567 (N_8567,N_7509,N_7427);
nand U8568 (N_8568,N_7328,N_7412);
and U8569 (N_8569,N_7628,N_7078);
and U8570 (N_8570,N_7553,N_7444);
or U8571 (N_8571,N_7280,N_7896);
nor U8572 (N_8572,N_7836,N_7969);
or U8573 (N_8573,N_7076,N_7042);
or U8574 (N_8574,N_7826,N_7999);
and U8575 (N_8575,N_7317,N_7353);
nor U8576 (N_8576,N_7882,N_7389);
and U8577 (N_8577,N_7829,N_7324);
nor U8578 (N_8578,N_7617,N_7318);
or U8579 (N_8579,N_7623,N_7790);
or U8580 (N_8580,N_7476,N_7233);
or U8581 (N_8581,N_7230,N_7227);
nand U8582 (N_8582,N_7760,N_7974);
nor U8583 (N_8583,N_7632,N_7075);
nand U8584 (N_8584,N_7858,N_7495);
nor U8585 (N_8585,N_7656,N_7511);
nand U8586 (N_8586,N_7533,N_7862);
nor U8587 (N_8587,N_7801,N_7459);
and U8588 (N_8588,N_7755,N_7924);
nor U8589 (N_8589,N_7105,N_7036);
nor U8590 (N_8590,N_7283,N_7267);
nor U8591 (N_8591,N_7632,N_7040);
nor U8592 (N_8592,N_7536,N_7693);
nor U8593 (N_8593,N_7441,N_7284);
nor U8594 (N_8594,N_7444,N_7380);
nand U8595 (N_8595,N_7046,N_7697);
or U8596 (N_8596,N_7243,N_7876);
nor U8597 (N_8597,N_7862,N_7271);
or U8598 (N_8598,N_7389,N_7664);
or U8599 (N_8599,N_7084,N_7353);
or U8600 (N_8600,N_7978,N_7265);
nor U8601 (N_8601,N_7081,N_7342);
or U8602 (N_8602,N_7263,N_7004);
or U8603 (N_8603,N_7203,N_7323);
and U8604 (N_8604,N_7067,N_7574);
nand U8605 (N_8605,N_7142,N_7931);
nand U8606 (N_8606,N_7188,N_7975);
nand U8607 (N_8607,N_7163,N_7311);
nand U8608 (N_8608,N_7730,N_7667);
and U8609 (N_8609,N_7451,N_7820);
nand U8610 (N_8610,N_7836,N_7651);
or U8611 (N_8611,N_7037,N_7164);
nand U8612 (N_8612,N_7223,N_7872);
and U8613 (N_8613,N_7554,N_7856);
and U8614 (N_8614,N_7286,N_7643);
nor U8615 (N_8615,N_7565,N_7348);
nor U8616 (N_8616,N_7334,N_7812);
nand U8617 (N_8617,N_7760,N_7731);
or U8618 (N_8618,N_7249,N_7781);
nand U8619 (N_8619,N_7630,N_7388);
nand U8620 (N_8620,N_7210,N_7995);
and U8621 (N_8621,N_7674,N_7933);
and U8622 (N_8622,N_7156,N_7108);
or U8623 (N_8623,N_7989,N_7073);
and U8624 (N_8624,N_7665,N_7811);
nor U8625 (N_8625,N_7948,N_7838);
nand U8626 (N_8626,N_7798,N_7966);
or U8627 (N_8627,N_7209,N_7941);
nor U8628 (N_8628,N_7021,N_7564);
nand U8629 (N_8629,N_7117,N_7434);
nand U8630 (N_8630,N_7397,N_7028);
nor U8631 (N_8631,N_7527,N_7692);
or U8632 (N_8632,N_7437,N_7759);
nor U8633 (N_8633,N_7815,N_7494);
and U8634 (N_8634,N_7016,N_7686);
or U8635 (N_8635,N_7964,N_7030);
nor U8636 (N_8636,N_7438,N_7358);
and U8637 (N_8637,N_7270,N_7564);
nor U8638 (N_8638,N_7508,N_7186);
nor U8639 (N_8639,N_7640,N_7768);
or U8640 (N_8640,N_7200,N_7085);
and U8641 (N_8641,N_7062,N_7928);
nor U8642 (N_8642,N_7150,N_7618);
nor U8643 (N_8643,N_7296,N_7584);
nand U8644 (N_8644,N_7054,N_7411);
nand U8645 (N_8645,N_7523,N_7220);
or U8646 (N_8646,N_7030,N_7796);
or U8647 (N_8647,N_7986,N_7293);
nand U8648 (N_8648,N_7450,N_7352);
or U8649 (N_8649,N_7171,N_7045);
nand U8650 (N_8650,N_7724,N_7867);
and U8651 (N_8651,N_7576,N_7585);
and U8652 (N_8652,N_7059,N_7629);
nor U8653 (N_8653,N_7986,N_7691);
and U8654 (N_8654,N_7250,N_7234);
or U8655 (N_8655,N_7950,N_7087);
nand U8656 (N_8656,N_7357,N_7711);
nor U8657 (N_8657,N_7621,N_7438);
or U8658 (N_8658,N_7499,N_7640);
nand U8659 (N_8659,N_7073,N_7884);
nand U8660 (N_8660,N_7079,N_7566);
and U8661 (N_8661,N_7532,N_7497);
nand U8662 (N_8662,N_7722,N_7187);
or U8663 (N_8663,N_7525,N_7096);
and U8664 (N_8664,N_7740,N_7560);
nor U8665 (N_8665,N_7825,N_7849);
nand U8666 (N_8666,N_7842,N_7393);
or U8667 (N_8667,N_7211,N_7106);
and U8668 (N_8668,N_7948,N_7482);
nand U8669 (N_8669,N_7866,N_7475);
nand U8670 (N_8670,N_7705,N_7013);
or U8671 (N_8671,N_7507,N_7625);
and U8672 (N_8672,N_7735,N_7271);
nand U8673 (N_8673,N_7327,N_7391);
nor U8674 (N_8674,N_7136,N_7856);
nor U8675 (N_8675,N_7933,N_7189);
nor U8676 (N_8676,N_7883,N_7684);
nand U8677 (N_8677,N_7328,N_7915);
and U8678 (N_8678,N_7109,N_7073);
or U8679 (N_8679,N_7055,N_7602);
or U8680 (N_8680,N_7794,N_7520);
nand U8681 (N_8681,N_7383,N_7533);
nor U8682 (N_8682,N_7679,N_7690);
or U8683 (N_8683,N_7500,N_7244);
nor U8684 (N_8684,N_7792,N_7014);
nor U8685 (N_8685,N_7251,N_7671);
or U8686 (N_8686,N_7036,N_7187);
nor U8687 (N_8687,N_7642,N_7614);
and U8688 (N_8688,N_7214,N_7883);
or U8689 (N_8689,N_7698,N_7597);
and U8690 (N_8690,N_7582,N_7120);
nor U8691 (N_8691,N_7439,N_7834);
nand U8692 (N_8692,N_7464,N_7359);
nor U8693 (N_8693,N_7280,N_7663);
or U8694 (N_8694,N_7116,N_7902);
and U8695 (N_8695,N_7810,N_7394);
nor U8696 (N_8696,N_7549,N_7645);
and U8697 (N_8697,N_7819,N_7729);
nor U8698 (N_8698,N_7724,N_7829);
nand U8699 (N_8699,N_7016,N_7032);
and U8700 (N_8700,N_7664,N_7857);
nor U8701 (N_8701,N_7650,N_7276);
nor U8702 (N_8702,N_7339,N_7062);
nor U8703 (N_8703,N_7681,N_7258);
nor U8704 (N_8704,N_7557,N_7248);
nor U8705 (N_8705,N_7636,N_7191);
or U8706 (N_8706,N_7494,N_7972);
or U8707 (N_8707,N_7453,N_7776);
and U8708 (N_8708,N_7793,N_7794);
nand U8709 (N_8709,N_7137,N_7548);
or U8710 (N_8710,N_7979,N_7537);
nor U8711 (N_8711,N_7918,N_7758);
or U8712 (N_8712,N_7687,N_7714);
or U8713 (N_8713,N_7746,N_7223);
or U8714 (N_8714,N_7202,N_7994);
or U8715 (N_8715,N_7886,N_7745);
and U8716 (N_8716,N_7731,N_7880);
or U8717 (N_8717,N_7421,N_7362);
and U8718 (N_8718,N_7821,N_7403);
or U8719 (N_8719,N_7371,N_7203);
or U8720 (N_8720,N_7897,N_7105);
or U8721 (N_8721,N_7578,N_7376);
and U8722 (N_8722,N_7404,N_7788);
or U8723 (N_8723,N_7980,N_7101);
nand U8724 (N_8724,N_7339,N_7713);
nor U8725 (N_8725,N_7543,N_7033);
or U8726 (N_8726,N_7774,N_7650);
nand U8727 (N_8727,N_7773,N_7353);
nand U8728 (N_8728,N_7274,N_7473);
nand U8729 (N_8729,N_7909,N_7530);
and U8730 (N_8730,N_7821,N_7536);
and U8731 (N_8731,N_7712,N_7339);
and U8732 (N_8732,N_7140,N_7519);
or U8733 (N_8733,N_7699,N_7868);
nand U8734 (N_8734,N_7432,N_7896);
nor U8735 (N_8735,N_7019,N_7543);
nor U8736 (N_8736,N_7223,N_7660);
and U8737 (N_8737,N_7870,N_7100);
and U8738 (N_8738,N_7309,N_7038);
xor U8739 (N_8739,N_7215,N_7057);
nor U8740 (N_8740,N_7835,N_7794);
nand U8741 (N_8741,N_7753,N_7540);
or U8742 (N_8742,N_7952,N_7231);
and U8743 (N_8743,N_7464,N_7628);
nand U8744 (N_8744,N_7649,N_7490);
and U8745 (N_8745,N_7657,N_7133);
and U8746 (N_8746,N_7630,N_7678);
or U8747 (N_8747,N_7007,N_7509);
or U8748 (N_8748,N_7378,N_7380);
nand U8749 (N_8749,N_7072,N_7310);
nor U8750 (N_8750,N_7012,N_7075);
and U8751 (N_8751,N_7750,N_7820);
and U8752 (N_8752,N_7926,N_7627);
nor U8753 (N_8753,N_7972,N_7636);
or U8754 (N_8754,N_7189,N_7741);
and U8755 (N_8755,N_7340,N_7466);
or U8756 (N_8756,N_7684,N_7129);
nand U8757 (N_8757,N_7378,N_7556);
nand U8758 (N_8758,N_7349,N_7216);
and U8759 (N_8759,N_7232,N_7673);
and U8760 (N_8760,N_7177,N_7962);
or U8761 (N_8761,N_7561,N_7639);
and U8762 (N_8762,N_7797,N_7472);
or U8763 (N_8763,N_7751,N_7358);
and U8764 (N_8764,N_7165,N_7357);
or U8765 (N_8765,N_7939,N_7792);
or U8766 (N_8766,N_7215,N_7044);
or U8767 (N_8767,N_7598,N_7989);
or U8768 (N_8768,N_7345,N_7951);
nand U8769 (N_8769,N_7437,N_7942);
nand U8770 (N_8770,N_7243,N_7783);
nor U8771 (N_8771,N_7796,N_7831);
and U8772 (N_8772,N_7255,N_7903);
or U8773 (N_8773,N_7522,N_7869);
nor U8774 (N_8774,N_7404,N_7384);
nand U8775 (N_8775,N_7186,N_7110);
and U8776 (N_8776,N_7195,N_7660);
nor U8777 (N_8777,N_7359,N_7194);
nand U8778 (N_8778,N_7917,N_7612);
nor U8779 (N_8779,N_7959,N_7392);
nand U8780 (N_8780,N_7897,N_7012);
nor U8781 (N_8781,N_7177,N_7283);
nor U8782 (N_8782,N_7363,N_7417);
and U8783 (N_8783,N_7136,N_7926);
and U8784 (N_8784,N_7010,N_7030);
and U8785 (N_8785,N_7717,N_7866);
nor U8786 (N_8786,N_7636,N_7399);
or U8787 (N_8787,N_7573,N_7152);
nand U8788 (N_8788,N_7791,N_7083);
nor U8789 (N_8789,N_7896,N_7157);
nand U8790 (N_8790,N_7926,N_7660);
and U8791 (N_8791,N_7335,N_7824);
nor U8792 (N_8792,N_7592,N_7925);
or U8793 (N_8793,N_7768,N_7764);
nor U8794 (N_8794,N_7655,N_7163);
nand U8795 (N_8795,N_7932,N_7042);
nor U8796 (N_8796,N_7856,N_7309);
and U8797 (N_8797,N_7733,N_7227);
nor U8798 (N_8798,N_7167,N_7208);
or U8799 (N_8799,N_7780,N_7715);
nor U8800 (N_8800,N_7582,N_7565);
or U8801 (N_8801,N_7382,N_7721);
or U8802 (N_8802,N_7460,N_7028);
nand U8803 (N_8803,N_7432,N_7293);
and U8804 (N_8804,N_7730,N_7036);
nor U8805 (N_8805,N_7817,N_7609);
or U8806 (N_8806,N_7880,N_7783);
or U8807 (N_8807,N_7992,N_7159);
or U8808 (N_8808,N_7492,N_7049);
nor U8809 (N_8809,N_7182,N_7958);
and U8810 (N_8810,N_7997,N_7923);
nor U8811 (N_8811,N_7421,N_7607);
nand U8812 (N_8812,N_7153,N_7133);
or U8813 (N_8813,N_7346,N_7710);
and U8814 (N_8814,N_7603,N_7194);
or U8815 (N_8815,N_7914,N_7448);
or U8816 (N_8816,N_7312,N_7795);
nand U8817 (N_8817,N_7037,N_7940);
nand U8818 (N_8818,N_7541,N_7862);
and U8819 (N_8819,N_7170,N_7823);
and U8820 (N_8820,N_7515,N_7516);
nand U8821 (N_8821,N_7699,N_7051);
nand U8822 (N_8822,N_7871,N_7282);
xnor U8823 (N_8823,N_7860,N_7780);
nor U8824 (N_8824,N_7813,N_7302);
and U8825 (N_8825,N_7353,N_7610);
or U8826 (N_8826,N_7073,N_7596);
and U8827 (N_8827,N_7154,N_7834);
or U8828 (N_8828,N_7266,N_7562);
or U8829 (N_8829,N_7245,N_7024);
nand U8830 (N_8830,N_7857,N_7567);
nor U8831 (N_8831,N_7304,N_7246);
xor U8832 (N_8832,N_7346,N_7736);
nand U8833 (N_8833,N_7565,N_7427);
nand U8834 (N_8834,N_7701,N_7729);
nor U8835 (N_8835,N_7752,N_7262);
and U8836 (N_8836,N_7567,N_7783);
nand U8837 (N_8837,N_7644,N_7579);
or U8838 (N_8838,N_7266,N_7604);
and U8839 (N_8839,N_7333,N_7730);
nor U8840 (N_8840,N_7507,N_7060);
nor U8841 (N_8841,N_7587,N_7836);
nor U8842 (N_8842,N_7345,N_7595);
or U8843 (N_8843,N_7633,N_7404);
nand U8844 (N_8844,N_7130,N_7049);
or U8845 (N_8845,N_7964,N_7043);
and U8846 (N_8846,N_7796,N_7426);
nor U8847 (N_8847,N_7954,N_7531);
or U8848 (N_8848,N_7093,N_7770);
nor U8849 (N_8849,N_7732,N_7255);
or U8850 (N_8850,N_7158,N_7396);
and U8851 (N_8851,N_7493,N_7326);
and U8852 (N_8852,N_7663,N_7391);
nand U8853 (N_8853,N_7683,N_7810);
and U8854 (N_8854,N_7621,N_7870);
and U8855 (N_8855,N_7357,N_7819);
and U8856 (N_8856,N_7987,N_7803);
or U8857 (N_8857,N_7113,N_7891);
nor U8858 (N_8858,N_7124,N_7846);
and U8859 (N_8859,N_7846,N_7152);
or U8860 (N_8860,N_7017,N_7583);
nor U8861 (N_8861,N_7610,N_7333);
and U8862 (N_8862,N_7911,N_7105);
and U8863 (N_8863,N_7709,N_7112);
nor U8864 (N_8864,N_7450,N_7735);
or U8865 (N_8865,N_7312,N_7301);
or U8866 (N_8866,N_7636,N_7873);
or U8867 (N_8867,N_7597,N_7504);
nor U8868 (N_8868,N_7858,N_7460);
nor U8869 (N_8869,N_7329,N_7331);
nand U8870 (N_8870,N_7483,N_7743);
nor U8871 (N_8871,N_7302,N_7405);
nand U8872 (N_8872,N_7152,N_7772);
and U8873 (N_8873,N_7859,N_7506);
nor U8874 (N_8874,N_7040,N_7297);
nand U8875 (N_8875,N_7243,N_7797);
nand U8876 (N_8876,N_7896,N_7811);
or U8877 (N_8877,N_7251,N_7726);
nand U8878 (N_8878,N_7464,N_7555);
nand U8879 (N_8879,N_7270,N_7540);
or U8880 (N_8880,N_7063,N_7267);
nor U8881 (N_8881,N_7517,N_7468);
nand U8882 (N_8882,N_7552,N_7520);
and U8883 (N_8883,N_7937,N_7187);
nor U8884 (N_8884,N_7458,N_7334);
nand U8885 (N_8885,N_7807,N_7110);
and U8886 (N_8886,N_7457,N_7002);
or U8887 (N_8887,N_7433,N_7136);
nor U8888 (N_8888,N_7075,N_7046);
or U8889 (N_8889,N_7157,N_7329);
and U8890 (N_8890,N_7580,N_7299);
and U8891 (N_8891,N_7584,N_7389);
and U8892 (N_8892,N_7036,N_7262);
nand U8893 (N_8893,N_7417,N_7655);
and U8894 (N_8894,N_7346,N_7856);
or U8895 (N_8895,N_7247,N_7446);
and U8896 (N_8896,N_7738,N_7769);
nor U8897 (N_8897,N_7439,N_7058);
nand U8898 (N_8898,N_7103,N_7675);
nand U8899 (N_8899,N_7765,N_7861);
nand U8900 (N_8900,N_7306,N_7977);
and U8901 (N_8901,N_7633,N_7792);
nor U8902 (N_8902,N_7622,N_7188);
nand U8903 (N_8903,N_7924,N_7809);
or U8904 (N_8904,N_7855,N_7443);
or U8905 (N_8905,N_7342,N_7514);
nand U8906 (N_8906,N_7285,N_7100);
nor U8907 (N_8907,N_7470,N_7099);
or U8908 (N_8908,N_7907,N_7602);
and U8909 (N_8909,N_7440,N_7892);
or U8910 (N_8910,N_7324,N_7464);
nor U8911 (N_8911,N_7603,N_7557);
nor U8912 (N_8912,N_7697,N_7225);
nand U8913 (N_8913,N_7510,N_7632);
and U8914 (N_8914,N_7864,N_7025);
nand U8915 (N_8915,N_7843,N_7980);
nor U8916 (N_8916,N_7347,N_7737);
and U8917 (N_8917,N_7313,N_7896);
nor U8918 (N_8918,N_7722,N_7617);
nor U8919 (N_8919,N_7806,N_7801);
and U8920 (N_8920,N_7292,N_7154);
and U8921 (N_8921,N_7760,N_7938);
nor U8922 (N_8922,N_7643,N_7371);
nor U8923 (N_8923,N_7275,N_7420);
nand U8924 (N_8924,N_7574,N_7048);
nand U8925 (N_8925,N_7179,N_7114);
nor U8926 (N_8926,N_7826,N_7446);
nor U8927 (N_8927,N_7780,N_7109);
nand U8928 (N_8928,N_7090,N_7558);
or U8929 (N_8929,N_7255,N_7343);
or U8930 (N_8930,N_7397,N_7222);
or U8931 (N_8931,N_7980,N_7013);
nor U8932 (N_8932,N_7911,N_7983);
xor U8933 (N_8933,N_7876,N_7076);
nand U8934 (N_8934,N_7158,N_7871);
and U8935 (N_8935,N_7032,N_7180);
or U8936 (N_8936,N_7429,N_7810);
nor U8937 (N_8937,N_7264,N_7429);
nor U8938 (N_8938,N_7445,N_7430);
or U8939 (N_8939,N_7262,N_7436);
and U8940 (N_8940,N_7225,N_7005);
nand U8941 (N_8941,N_7302,N_7131);
or U8942 (N_8942,N_7033,N_7503);
nand U8943 (N_8943,N_7431,N_7832);
or U8944 (N_8944,N_7595,N_7694);
nor U8945 (N_8945,N_7256,N_7106);
or U8946 (N_8946,N_7388,N_7851);
nor U8947 (N_8947,N_7745,N_7334);
or U8948 (N_8948,N_7992,N_7658);
and U8949 (N_8949,N_7403,N_7284);
nor U8950 (N_8950,N_7351,N_7624);
nand U8951 (N_8951,N_7558,N_7962);
or U8952 (N_8952,N_7746,N_7518);
and U8953 (N_8953,N_7008,N_7112);
nor U8954 (N_8954,N_7601,N_7036);
nand U8955 (N_8955,N_7377,N_7575);
nand U8956 (N_8956,N_7148,N_7762);
nand U8957 (N_8957,N_7260,N_7104);
nand U8958 (N_8958,N_7177,N_7393);
xnor U8959 (N_8959,N_7151,N_7784);
nor U8960 (N_8960,N_7727,N_7427);
nor U8961 (N_8961,N_7558,N_7569);
nor U8962 (N_8962,N_7584,N_7190);
and U8963 (N_8963,N_7443,N_7127);
nor U8964 (N_8964,N_7369,N_7810);
and U8965 (N_8965,N_7850,N_7032);
nor U8966 (N_8966,N_7874,N_7504);
nor U8967 (N_8967,N_7490,N_7349);
nor U8968 (N_8968,N_7136,N_7067);
nand U8969 (N_8969,N_7716,N_7087);
nor U8970 (N_8970,N_7112,N_7084);
nand U8971 (N_8971,N_7134,N_7146);
nor U8972 (N_8972,N_7752,N_7688);
nor U8973 (N_8973,N_7473,N_7039);
nor U8974 (N_8974,N_7123,N_7752);
nor U8975 (N_8975,N_7930,N_7013);
and U8976 (N_8976,N_7327,N_7757);
nand U8977 (N_8977,N_7884,N_7635);
or U8978 (N_8978,N_7682,N_7677);
and U8979 (N_8979,N_7539,N_7835);
or U8980 (N_8980,N_7128,N_7749);
nand U8981 (N_8981,N_7571,N_7252);
nor U8982 (N_8982,N_7106,N_7660);
nor U8983 (N_8983,N_7807,N_7552);
nand U8984 (N_8984,N_7056,N_7960);
nor U8985 (N_8985,N_7819,N_7756);
nand U8986 (N_8986,N_7802,N_7331);
nand U8987 (N_8987,N_7294,N_7239);
or U8988 (N_8988,N_7820,N_7266);
nand U8989 (N_8989,N_7682,N_7526);
and U8990 (N_8990,N_7306,N_7300);
and U8991 (N_8991,N_7736,N_7148);
and U8992 (N_8992,N_7319,N_7300);
nand U8993 (N_8993,N_7741,N_7644);
nor U8994 (N_8994,N_7712,N_7466);
or U8995 (N_8995,N_7332,N_7956);
nand U8996 (N_8996,N_7354,N_7023);
nor U8997 (N_8997,N_7438,N_7628);
and U8998 (N_8998,N_7243,N_7354);
or U8999 (N_8999,N_7632,N_7462);
and U9000 (N_9000,N_8863,N_8864);
and U9001 (N_9001,N_8611,N_8545);
and U9002 (N_9002,N_8793,N_8956);
nand U9003 (N_9003,N_8785,N_8102);
nor U9004 (N_9004,N_8052,N_8645);
nand U9005 (N_9005,N_8597,N_8766);
and U9006 (N_9006,N_8518,N_8300);
or U9007 (N_9007,N_8696,N_8092);
xnor U9008 (N_9008,N_8192,N_8870);
or U9009 (N_9009,N_8234,N_8682);
nor U9010 (N_9010,N_8888,N_8834);
nor U9011 (N_9011,N_8889,N_8925);
and U9012 (N_9012,N_8561,N_8240);
nand U9013 (N_9013,N_8410,N_8690);
nor U9014 (N_9014,N_8968,N_8097);
and U9015 (N_9015,N_8231,N_8141);
and U9016 (N_9016,N_8995,N_8602);
nor U9017 (N_9017,N_8782,N_8294);
nor U9018 (N_9018,N_8389,N_8124);
nand U9019 (N_9019,N_8081,N_8633);
nor U9020 (N_9020,N_8773,N_8938);
or U9021 (N_9021,N_8164,N_8781);
nor U9022 (N_9022,N_8107,N_8483);
nor U9023 (N_9023,N_8718,N_8387);
and U9024 (N_9024,N_8642,N_8018);
and U9025 (N_9025,N_8087,N_8072);
and U9026 (N_9026,N_8813,N_8810);
or U9027 (N_9027,N_8803,N_8046);
nor U9028 (N_9028,N_8839,N_8400);
or U9029 (N_9029,N_8048,N_8783);
nor U9030 (N_9030,N_8957,N_8599);
and U9031 (N_9031,N_8179,N_8257);
or U9032 (N_9032,N_8574,N_8986);
nand U9033 (N_9033,N_8011,N_8722);
nor U9034 (N_9034,N_8104,N_8233);
and U9035 (N_9035,N_8262,N_8103);
or U9036 (N_9036,N_8306,N_8588);
and U9037 (N_9037,N_8427,N_8249);
nand U9038 (N_9038,N_8003,N_8659);
and U9039 (N_9039,N_8085,N_8002);
or U9040 (N_9040,N_8130,N_8496);
nand U9041 (N_9041,N_8969,N_8648);
and U9042 (N_9042,N_8733,N_8425);
nor U9043 (N_9043,N_8592,N_8279);
and U9044 (N_9044,N_8122,N_8949);
nor U9045 (N_9045,N_8035,N_8355);
nor U9046 (N_9046,N_8579,N_8846);
nand U9047 (N_9047,N_8874,N_8487);
nor U9048 (N_9048,N_8027,N_8896);
nor U9049 (N_9049,N_8150,N_8907);
nand U9050 (N_9050,N_8050,N_8068);
nor U9051 (N_9051,N_8376,N_8833);
and U9052 (N_9052,N_8394,N_8109);
nand U9053 (N_9053,N_8522,N_8503);
nor U9054 (N_9054,N_8190,N_8212);
nand U9055 (N_9055,N_8251,N_8662);
nand U9056 (N_9056,N_8751,N_8587);
or U9057 (N_9057,N_8866,N_8821);
nand U9058 (N_9058,N_8258,N_8537);
and U9059 (N_9059,N_8631,N_8308);
nor U9060 (N_9060,N_8379,N_8559);
nor U9061 (N_9061,N_8033,N_8731);
and U9062 (N_9062,N_8296,N_8643);
or U9063 (N_9063,N_8005,N_8393);
and U9064 (N_9064,N_8418,N_8143);
and U9065 (N_9065,N_8416,N_8026);
or U9066 (N_9066,N_8309,N_8290);
nand U9067 (N_9067,N_8254,N_8570);
nor U9068 (N_9068,N_8719,N_8346);
nand U9069 (N_9069,N_8041,N_8961);
and U9070 (N_9070,N_8182,N_8712);
or U9071 (N_9071,N_8446,N_8276);
or U9072 (N_9072,N_8165,N_8535);
nand U9073 (N_9073,N_8600,N_8827);
nand U9074 (N_9074,N_8553,N_8637);
or U9075 (N_9075,N_8186,N_8057);
and U9076 (N_9076,N_8589,N_8009);
nand U9077 (N_9077,N_8541,N_8621);
and U9078 (N_9078,N_8871,N_8590);
nand U9079 (N_9079,N_8271,N_8530);
nand U9080 (N_9080,N_8170,N_8855);
nor U9081 (N_9081,N_8489,N_8307);
and U9082 (N_9082,N_8322,N_8721);
or U9083 (N_9083,N_8664,N_8460);
nand U9084 (N_9084,N_8241,N_8550);
or U9085 (N_9085,N_8581,N_8204);
nand U9086 (N_9086,N_8449,N_8923);
or U9087 (N_9087,N_8112,N_8804);
nor U9088 (N_9088,N_8649,N_8944);
and U9089 (N_9089,N_8634,N_8504);
nand U9090 (N_9090,N_8922,N_8730);
nand U9091 (N_9091,N_8595,N_8998);
and U9092 (N_9092,N_8129,N_8511);
nand U9093 (N_9093,N_8420,N_8630);
or U9094 (N_9094,N_8685,N_8706);
or U9095 (N_9095,N_8049,N_8434);
and U9096 (N_9096,N_8353,N_8282);
nand U9097 (N_9097,N_8137,N_8554);
nor U9098 (N_9098,N_8572,N_8191);
nor U9099 (N_9099,N_8728,N_8275);
and U9100 (N_9100,N_8937,N_8726);
nand U9101 (N_9101,N_8646,N_8490);
or U9102 (N_9102,N_8264,N_8565);
and U9103 (N_9103,N_8246,N_8983);
or U9104 (N_9104,N_8310,N_8734);
nand U9105 (N_9105,N_8203,N_8914);
and U9106 (N_9106,N_8705,N_8950);
nand U9107 (N_9107,N_8348,N_8845);
or U9108 (N_9108,N_8911,N_8534);
nand U9109 (N_9109,N_8133,N_8209);
and U9110 (N_9110,N_8283,N_8473);
nand U9111 (N_9111,N_8878,N_8096);
or U9112 (N_9112,N_8252,N_8628);
or U9113 (N_9113,N_8178,N_8698);
nor U9114 (N_9114,N_8008,N_8516);
nand U9115 (N_9115,N_8181,N_8876);
nand U9116 (N_9116,N_8510,N_8720);
nor U9117 (N_9117,N_8985,N_8711);
nor U9118 (N_9118,N_8993,N_8082);
nor U9119 (N_9119,N_8683,N_8524);
nor U9120 (N_9120,N_8399,N_8342);
and U9121 (N_9121,N_8612,N_8789);
nand U9122 (N_9122,N_8753,N_8476);
or U9123 (N_9123,N_8029,N_8594);
nand U9124 (N_9124,N_8982,N_8139);
and U9125 (N_9125,N_8532,N_8875);
nand U9126 (N_9126,N_8152,N_8591);
and U9127 (N_9127,N_8681,N_8218);
nand U9128 (N_9128,N_8984,N_8134);
and U9129 (N_9129,N_8397,N_8090);
nand U9130 (N_9130,N_8486,N_8071);
and U9131 (N_9131,N_8975,N_8910);
nand U9132 (N_9132,N_8287,N_8341);
nor U9133 (N_9133,N_8336,N_8172);
or U9134 (N_9134,N_8948,N_8183);
nor U9135 (N_9135,N_8177,N_8135);
nor U9136 (N_9136,N_8635,N_8061);
or U9137 (N_9137,N_8811,N_8759);
and U9138 (N_9138,N_8089,N_8801);
or U9139 (N_9139,N_8185,N_8551);
nand U9140 (N_9140,N_8432,N_8981);
or U9141 (N_9141,N_8429,N_8325);
or U9142 (N_9142,N_8031,N_8247);
nand U9143 (N_9143,N_8277,N_8892);
and U9144 (N_9144,N_8515,N_8442);
nand U9145 (N_9145,N_8064,N_8056);
and U9146 (N_9146,N_8268,N_8661);
nor U9147 (N_9147,N_8067,N_8641);
xor U9148 (N_9148,N_8020,N_8802);
and U9149 (N_9149,N_8672,N_8381);
nand U9150 (N_9150,N_8319,N_8256);
and U9151 (N_9151,N_8676,N_8528);
and U9152 (N_9152,N_8882,N_8780);
or U9153 (N_9153,N_8739,N_8361);
nand U9154 (N_9154,N_8909,N_8059);
and U9155 (N_9155,N_8086,N_8001);
and U9156 (N_9156,N_8737,N_8768);
nor U9157 (N_9157,N_8464,N_8184);
nand U9158 (N_9158,N_8622,N_8229);
and U9159 (N_9159,N_8304,N_8750);
nand U9160 (N_9160,N_8273,N_8312);
nand U9161 (N_9161,N_8408,N_8512);
nand U9162 (N_9162,N_8604,N_8508);
or U9163 (N_9163,N_8941,N_8580);
nor U9164 (N_9164,N_8838,N_8119);
nand U9165 (N_9165,N_8514,N_8270);
and U9166 (N_9166,N_8413,N_8374);
and U9167 (N_9167,N_8208,N_8468);
nand U9168 (N_9168,N_8971,N_8166);
and U9169 (N_9169,N_8852,N_8105);
nor U9170 (N_9170,N_8930,N_8019);
nand U9171 (N_9171,N_8223,N_8378);
and U9172 (N_9172,N_8142,N_8441);
or U9173 (N_9173,N_8349,N_8552);
and U9174 (N_9174,N_8422,N_8851);
nor U9175 (N_9175,N_8558,N_8313);
nand U9176 (N_9176,N_8195,N_8692);
nand U9177 (N_9177,N_8868,N_8638);
nor U9178 (N_9178,N_8673,N_8106);
nor U9179 (N_9179,N_8707,N_8974);
nor U9180 (N_9180,N_8761,N_8154);
nor U9181 (N_9181,N_8458,N_8727);
and U9182 (N_9182,N_8873,N_8776);
nor U9183 (N_9183,N_8653,N_8538);
and U9184 (N_9184,N_8323,N_8363);
or U9185 (N_9185,N_8715,N_8402);
nand U9186 (N_9186,N_8286,N_8808);
nor U9187 (N_9187,N_8474,N_8526);
or U9188 (N_9188,N_8237,N_8140);
or U9189 (N_9189,N_8367,N_8301);
nor U9190 (N_9190,N_8385,N_8610);
and U9191 (N_9191,N_8453,N_8230);
and U9192 (N_9192,N_8853,N_8435);
or U9193 (N_9193,N_8467,N_8132);
nor U9194 (N_9194,N_8384,N_8226);
nor U9195 (N_9195,N_8762,N_8679);
or U9196 (N_9196,N_8797,N_8274);
or U9197 (N_9197,N_8980,N_8639);
nand U9198 (N_9198,N_8831,N_8740);
and U9199 (N_9199,N_8160,N_8098);
nand U9200 (N_9200,N_8702,N_8555);
and U9201 (N_9201,N_8636,N_8828);
nor U9202 (N_9202,N_8830,N_8678);
or U9203 (N_9203,N_8004,N_8284);
or U9204 (N_9204,N_8859,N_8517);
nor U9205 (N_9205,N_8094,N_8560);
nor U9206 (N_9206,N_8025,N_8652);
nor U9207 (N_9207,N_8860,N_8723);
or U9208 (N_9208,N_8916,N_8841);
nor U9209 (N_9209,N_8862,N_8735);
nand U9210 (N_9210,N_8298,N_8812);
nor U9211 (N_9211,N_8593,N_8280);
xor U9212 (N_9212,N_8847,N_8655);
and U9213 (N_9213,N_8421,N_8778);
nor U9214 (N_9214,N_8749,N_8902);
nand U9215 (N_9215,N_8539,N_8585);
nand U9216 (N_9216,N_8239,N_8668);
and U9217 (N_9217,N_8794,N_8343);
or U9218 (N_9218,N_8625,N_8083);
or U9219 (N_9219,N_8644,N_8375);
or U9220 (N_9220,N_8475,N_8962);
nor U9221 (N_9221,N_8564,N_8640);
nand U9222 (N_9222,N_8099,N_8372);
nand U9223 (N_9223,N_8713,N_8525);
nand U9224 (N_9224,N_8777,N_8665);
nand U9225 (N_9225,N_8255,N_8656);
and U9226 (N_9226,N_8278,N_8996);
nand U9227 (N_9227,N_8775,N_8111);
and U9228 (N_9228,N_8055,N_8335);
and U9229 (N_9229,N_8037,N_8651);
or U9230 (N_9230,N_8684,N_8044);
and U9231 (N_9231,N_8695,N_8745);
and U9232 (N_9232,N_8285,N_8471);
or U9233 (N_9233,N_8158,N_8469);
nand U9234 (N_9234,N_8836,N_8125);
or U9235 (N_9235,N_8663,N_8500);
nor U9236 (N_9236,N_8890,N_8670);
nand U9237 (N_9237,N_8350,N_8933);
and U9238 (N_9238,N_8763,N_8114);
or U9239 (N_9239,N_8197,N_8215);
and U9240 (N_9240,N_8791,N_8613);
and U9241 (N_9241,N_8596,N_8459);
nor U9242 (N_9242,N_8603,N_8014);
or U9243 (N_9243,N_8382,N_8054);
nor U9244 (N_9244,N_8314,N_8430);
or U9245 (N_9245,N_8347,N_8201);
and U9246 (N_9246,N_8771,N_8118);
and U9247 (N_9247,N_8932,N_8303);
or U9248 (N_9248,N_8758,N_8492);
nor U9249 (N_9249,N_8607,N_8042);
nand U9250 (N_9250,N_8513,N_8491);
nor U9251 (N_9251,N_8438,N_8199);
or U9252 (N_9252,N_8428,N_8499);
or U9253 (N_9253,N_8955,N_8076);
nand U9254 (N_9254,N_8970,N_8917);
nand U9255 (N_9255,N_8787,N_8481);
and U9256 (N_9256,N_8666,N_8127);
and U9257 (N_9257,N_8318,N_8079);
and U9258 (N_9258,N_8232,N_8360);
nor U9259 (N_9259,N_8686,N_8138);
nor U9260 (N_9260,N_8293,N_8484);
nor U9261 (N_9261,N_8879,N_8764);
xnor U9262 (N_9262,N_8920,N_8894);
and U9263 (N_9263,N_8153,N_8899);
and U9264 (N_9264,N_8624,N_8887);
nand U9265 (N_9265,N_8126,N_8189);
nand U9266 (N_9266,N_8222,N_8359);
nor U9267 (N_9267,N_8886,N_8716);
nand U9268 (N_9268,N_8929,N_8045);
nor U9269 (N_9269,N_8989,N_8131);
nor U9270 (N_9270,N_8462,N_8339);
nand U9271 (N_9271,N_8149,N_8842);
and U9272 (N_9272,N_8835,N_8904);
or U9273 (N_9273,N_8786,N_8582);
nand U9274 (N_9274,N_8034,N_8444);
or U9275 (N_9275,N_8908,N_8893);
or U9276 (N_9276,N_8036,N_8927);
nand U9277 (N_9277,N_8340,N_8704);
nand U9278 (N_9278,N_8945,N_8015);
and U9279 (N_9279,N_8433,N_8479);
and U9280 (N_9280,N_8891,N_8966);
and U9281 (N_9281,N_8242,N_8798);
nand U9282 (N_9282,N_8742,N_8167);
nand U9283 (N_9283,N_8746,N_8939);
nand U9284 (N_9284,N_8465,N_8850);
or U9285 (N_9285,N_8795,N_8299);
nand U9286 (N_9286,N_8338,N_8392);
xnor U9287 (N_9287,N_8368,N_8480);
or U9288 (N_9288,N_8337,N_8669);
or U9289 (N_9289,N_8877,N_8128);
or U9290 (N_9290,N_8988,N_8088);
nand U9291 (N_9291,N_8080,N_8176);
nor U9292 (N_9292,N_8617,N_8245);
and U9293 (N_9293,N_8155,N_8136);
or U9294 (N_9294,N_8997,N_8329);
nor U9295 (N_9295,N_8253,N_8395);
or U9296 (N_9296,N_8028,N_8717);
nor U9297 (N_9297,N_8583,N_8302);
or U9298 (N_9298,N_8063,N_8292);
nand U9299 (N_9299,N_8675,N_8194);
and U9300 (N_9300,N_8832,N_8806);
and U9301 (N_9301,N_8010,N_8440);
nor U9302 (N_9302,N_8963,N_8823);
nand U9303 (N_9303,N_8236,N_8542);
nand U9304 (N_9304,N_8169,N_8324);
or U9305 (N_9305,N_8403,N_8942);
and U9306 (N_9306,N_8447,N_8326);
nor U9307 (N_9307,N_8168,N_8881);
or U9308 (N_9308,N_8770,N_8990);
nand U9309 (N_9309,N_8437,N_8536);
or U9310 (N_9310,N_8405,N_8615);
nor U9311 (N_9311,N_8211,N_8609);
and U9312 (N_9312,N_8305,N_8021);
nand U9313 (N_9313,N_8784,N_8022);
and U9314 (N_9314,N_8912,N_8987);
nor U9315 (N_9315,N_8108,N_8115);
or U9316 (N_9316,N_8216,N_8901);
nand U9317 (N_9317,N_8498,N_8423);
and U9318 (N_9318,N_8573,N_8463);
or U9319 (N_9319,N_8977,N_8461);
nand U9320 (N_9320,N_8123,N_8743);
or U9321 (N_9321,N_8334,N_8578);
xnor U9322 (N_9322,N_8358,N_8819);
nor U9323 (N_9323,N_8225,N_8066);
nand U9324 (N_9324,N_8629,N_8936);
nand U9325 (N_9325,N_8238,N_8947);
nand U9326 (N_9326,N_8872,N_8884);
nor U9327 (N_9327,N_8073,N_8466);
nand U9328 (N_9328,N_8327,N_8865);
and U9329 (N_9329,N_8965,N_8978);
or U9330 (N_9330,N_8404,N_8084);
nand U9331 (N_9331,N_8546,N_8747);
and U9332 (N_9332,N_8171,N_8840);
and U9333 (N_9333,N_8032,N_8352);
nand U9334 (N_9334,N_8576,N_8556);
and U9335 (N_9335,N_8991,N_8390);
nor U9336 (N_9336,N_8210,N_8869);
and U9337 (N_9337,N_8566,N_8012);
or U9338 (N_9338,N_8674,N_8671);
nor U9339 (N_9339,N_8626,N_8934);
and U9340 (N_9340,N_8267,N_8288);
or U9341 (N_9341,N_8219,N_8188);
and U9342 (N_9342,N_8040,N_8657);
nor U9343 (N_9343,N_8605,N_8807);
nor U9344 (N_9344,N_8577,N_8206);
nor U9345 (N_9345,N_8654,N_8744);
and U9346 (N_9346,N_8826,N_8790);
or U9347 (N_9347,N_8456,N_8752);
and U9348 (N_9348,N_8470,N_8356);
or U9349 (N_9349,N_8344,N_8755);
nand U9350 (N_9350,N_8488,N_8448);
or U9351 (N_9351,N_8161,N_8820);
nor U9352 (N_9352,N_8958,N_8151);
nand U9353 (N_9353,N_8482,N_8815);
nor U9354 (N_9354,N_8074,N_8883);
nor U9355 (N_9355,N_8217,N_8691);
and U9356 (N_9356,N_8919,N_8398);
or U9357 (N_9357,N_8162,N_8620);
nor U9358 (N_9358,N_8414,N_8485);
nand U9359 (N_9359,N_8260,N_8412);
or U9360 (N_9360,N_8321,N_8584);
nor U9361 (N_9361,N_8415,N_8024);
or U9362 (N_9362,N_8297,N_8898);
and U9363 (N_9363,N_8994,N_8380);
and U9364 (N_9364,N_8903,N_8954);
nor U9365 (N_9365,N_8051,N_8924);
nor U9366 (N_9366,N_8295,N_8366);
nor U9367 (N_9367,N_8935,N_8885);
nor U9368 (N_9368,N_8992,N_8562);
or U9369 (N_9369,N_8330,N_8450);
nor U9370 (N_9370,N_8494,N_8354);
or U9371 (N_9371,N_8502,N_8601);
nor U9372 (N_9372,N_8013,N_8221);
nand U9373 (N_9373,N_8703,N_8436);
nor U9374 (N_9374,N_8200,N_8159);
nand U9375 (N_9375,N_8999,N_8364);
nor U9376 (N_9376,N_8388,N_8235);
or U9377 (N_9377,N_8523,N_8623);
and U9378 (N_9378,N_8175,N_8953);
or U9379 (N_9379,N_8207,N_8571);
nand U9380 (N_9380,N_8224,N_8091);
nor U9381 (N_9381,N_8362,N_8227);
and U9382 (N_9382,N_8814,N_8976);
nor U9383 (N_9383,N_8757,N_8548);
nand U9384 (N_9384,N_8694,N_8401);
nand U9385 (N_9385,N_8915,N_8660);
or U9386 (N_9386,N_8493,N_8431);
nand U9387 (N_9387,N_8822,N_8895);
xnor U9388 (N_9388,N_8078,N_8047);
or U9389 (N_9389,N_8693,N_8117);
or U9390 (N_9390,N_8861,N_8960);
and U9391 (N_9391,N_8316,N_8365);
nand U9392 (N_9392,N_8809,N_8799);
nor U9393 (N_9393,N_8451,N_8765);
nand U9394 (N_9394,N_8426,N_8101);
or U9395 (N_9395,N_8658,N_8419);
or U9396 (N_9396,N_8501,N_8213);
nor U9397 (N_9397,N_8187,N_8931);
or U9398 (N_9398,N_8913,N_8650);
or U9399 (N_9399,N_8849,N_8272);
xnor U9400 (N_9400,N_8767,N_8598);
nor U9401 (N_9401,N_8825,N_8069);
and U9402 (N_9402,N_8265,N_8320);
or U9403 (N_9403,N_8900,N_8618);
nor U9404 (N_9404,N_8688,N_8824);
or U9405 (N_9405,N_8848,N_8519);
nand U9406 (N_9406,N_8829,N_8311);
nand U9407 (N_9407,N_8406,N_8369);
and U9408 (N_9408,N_8505,N_8699);
nand U9409 (N_9409,N_8529,N_8120);
or U9410 (N_9410,N_8856,N_8043);
or U9411 (N_9411,N_8383,N_8291);
nor U9412 (N_9412,N_8972,N_8805);
nor U9413 (N_9413,N_8928,N_8738);
and U9414 (N_9414,N_8506,N_8144);
or U9415 (N_9415,N_8880,N_8921);
or U9416 (N_9416,N_8053,N_8214);
and U9417 (N_9417,N_8951,N_8926);
nor U9418 (N_9418,N_8077,N_8250);
nor U9419 (N_9419,N_8575,N_8547);
or U9420 (N_9420,N_8754,N_8736);
and U9421 (N_9421,N_8455,N_8608);
or U9422 (N_9422,N_8331,N_8680);
nand U9423 (N_9423,N_8345,N_8544);
nand U9424 (N_9424,N_8193,N_8452);
and U9425 (N_9425,N_8697,N_8454);
and U9426 (N_9426,N_8017,N_8006);
or U9427 (N_9427,N_8220,N_8687);
or U9428 (N_9428,N_8202,N_8606);
nor U9429 (N_9429,N_8248,N_8632);
nor U9430 (N_9430,N_8281,N_8979);
or U9431 (N_9431,N_8586,N_8445);
nand U9432 (N_9432,N_8946,N_8816);
or U9433 (N_9433,N_8509,N_8520);
and U9434 (N_9434,N_8373,N_8093);
or U9435 (N_9435,N_8708,N_8146);
nor U9436 (N_9436,N_8269,N_8351);
nand U9437 (N_9437,N_8614,N_8147);
nor U9438 (N_9438,N_8689,N_8774);
nor U9439 (N_9439,N_8725,N_8243);
or U9440 (N_9440,N_8407,N_8180);
nand U9441 (N_9441,N_8918,N_8837);
or U9442 (N_9442,N_8205,N_8062);
or U9443 (N_9443,N_8732,N_8409);
nand U9444 (N_9444,N_8521,N_8244);
nand U9445 (N_9445,N_8148,N_8779);
or U9446 (N_9446,N_8332,N_8677);
nand U9447 (N_9447,N_8060,N_8800);
nand U9448 (N_9448,N_8616,N_8844);
nand U9449 (N_9449,N_8095,N_8495);
and U9450 (N_9450,N_8391,N_8039);
and U9451 (N_9451,N_8328,N_8943);
nor U9452 (N_9452,N_8163,N_8058);
or U9453 (N_9453,N_8396,N_8619);
and U9454 (N_9454,N_8477,N_8100);
nor U9455 (N_9455,N_8357,N_8075);
and U9456 (N_9456,N_8443,N_8905);
nand U9457 (N_9457,N_8647,N_8457);
nand U9458 (N_9458,N_8370,N_8792);
nor U9459 (N_9459,N_8769,N_8964);
or U9460 (N_9460,N_8424,N_8569);
nor U9461 (N_9461,N_8173,N_8507);
or U9462 (N_9462,N_8315,N_8940);
or U9463 (N_9463,N_8858,N_8741);
or U9464 (N_9464,N_8016,N_8897);
and U9465 (N_9465,N_8709,N_8540);
or U9466 (N_9466,N_8198,N_8817);
and U9467 (N_9467,N_8007,N_8796);
or U9468 (N_9468,N_8377,N_8714);
or U9469 (N_9469,N_8371,N_8478);
nand U9470 (N_9470,N_8317,N_8563);
and U9471 (N_9471,N_8116,N_8857);
nand U9472 (N_9472,N_8070,N_8867);
nand U9473 (N_9473,N_8667,N_8065);
and U9474 (N_9474,N_8568,N_8818);
or U9475 (N_9475,N_8417,N_8110);
nand U9476 (N_9476,N_8266,N_8228);
or U9477 (N_9477,N_8527,N_8531);
and U9478 (N_9478,N_8729,N_8174);
nand U9479 (N_9479,N_8973,N_8121);
and U9480 (N_9480,N_8439,N_8156);
and U9481 (N_9481,N_8038,N_8543);
and U9482 (N_9482,N_8760,N_8567);
nand U9483 (N_9483,N_8756,N_8772);
and U9484 (N_9484,N_8627,N_8557);
nor U9485 (N_9485,N_8710,N_8145);
nand U9486 (N_9486,N_8533,N_8700);
nor U9487 (N_9487,N_8701,N_8959);
nand U9488 (N_9488,N_8549,N_8196);
or U9489 (N_9489,N_8333,N_8000);
and U9490 (N_9490,N_8497,N_8023);
and U9491 (N_9491,N_8748,N_8289);
nor U9492 (N_9492,N_8952,N_8411);
and U9493 (N_9493,N_8854,N_8843);
and U9494 (N_9494,N_8967,N_8263);
nor U9495 (N_9495,N_8906,N_8386);
and U9496 (N_9496,N_8724,N_8259);
and U9497 (N_9497,N_8261,N_8113);
and U9498 (N_9498,N_8157,N_8788);
or U9499 (N_9499,N_8030,N_8472);
xnor U9500 (N_9500,N_8521,N_8079);
and U9501 (N_9501,N_8759,N_8769);
and U9502 (N_9502,N_8866,N_8679);
or U9503 (N_9503,N_8487,N_8744);
nor U9504 (N_9504,N_8358,N_8723);
or U9505 (N_9505,N_8713,N_8371);
nand U9506 (N_9506,N_8186,N_8731);
nand U9507 (N_9507,N_8804,N_8414);
xor U9508 (N_9508,N_8623,N_8541);
or U9509 (N_9509,N_8701,N_8848);
nand U9510 (N_9510,N_8705,N_8936);
and U9511 (N_9511,N_8396,N_8659);
nand U9512 (N_9512,N_8916,N_8135);
nand U9513 (N_9513,N_8486,N_8139);
or U9514 (N_9514,N_8796,N_8560);
nor U9515 (N_9515,N_8748,N_8158);
or U9516 (N_9516,N_8597,N_8979);
nor U9517 (N_9517,N_8766,N_8337);
nand U9518 (N_9518,N_8262,N_8020);
and U9519 (N_9519,N_8885,N_8454);
nand U9520 (N_9520,N_8196,N_8383);
nor U9521 (N_9521,N_8833,N_8727);
nand U9522 (N_9522,N_8312,N_8935);
nor U9523 (N_9523,N_8501,N_8385);
xnor U9524 (N_9524,N_8646,N_8931);
nand U9525 (N_9525,N_8660,N_8633);
nand U9526 (N_9526,N_8758,N_8385);
and U9527 (N_9527,N_8598,N_8947);
nand U9528 (N_9528,N_8188,N_8680);
xor U9529 (N_9529,N_8494,N_8338);
nand U9530 (N_9530,N_8175,N_8499);
nor U9531 (N_9531,N_8567,N_8062);
nand U9532 (N_9532,N_8707,N_8664);
nand U9533 (N_9533,N_8965,N_8283);
nand U9534 (N_9534,N_8294,N_8820);
nor U9535 (N_9535,N_8230,N_8020);
nor U9536 (N_9536,N_8797,N_8195);
or U9537 (N_9537,N_8964,N_8633);
and U9538 (N_9538,N_8770,N_8369);
nor U9539 (N_9539,N_8137,N_8318);
or U9540 (N_9540,N_8113,N_8523);
nor U9541 (N_9541,N_8047,N_8724);
nor U9542 (N_9542,N_8073,N_8165);
nor U9543 (N_9543,N_8282,N_8449);
and U9544 (N_9544,N_8667,N_8835);
nand U9545 (N_9545,N_8563,N_8535);
nor U9546 (N_9546,N_8170,N_8973);
or U9547 (N_9547,N_8619,N_8835);
nor U9548 (N_9548,N_8351,N_8239);
nor U9549 (N_9549,N_8107,N_8578);
and U9550 (N_9550,N_8974,N_8630);
nor U9551 (N_9551,N_8808,N_8974);
nand U9552 (N_9552,N_8977,N_8560);
nor U9553 (N_9553,N_8096,N_8301);
or U9554 (N_9554,N_8359,N_8649);
nand U9555 (N_9555,N_8346,N_8528);
and U9556 (N_9556,N_8755,N_8970);
and U9557 (N_9557,N_8393,N_8866);
nor U9558 (N_9558,N_8511,N_8703);
or U9559 (N_9559,N_8830,N_8810);
nor U9560 (N_9560,N_8821,N_8395);
and U9561 (N_9561,N_8881,N_8677);
nand U9562 (N_9562,N_8643,N_8810);
nor U9563 (N_9563,N_8563,N_8681);
and U9564 (N_9564,N_8118,N_8960);
nand U9565 (N_9565,N_8506,N_8573);
nand U9566 (N_9566,N_8144,N_8626);
and U9567 (N_9567,N_8453,N_8321);
nor U9568 (N_9568,N_8126,N_8375);
and U9569 (N_9569,N_8922,N_8984);
and U9570 (N_9570,N_8786,N_8989);
nor U9571 (N_9571,N_8972,N_8969);
and U9572 (N_9572,N_8346,N_8122);
nand U9573 (N_9573,N_8724,N_8737);
nor U9574 (N_9574,N_8255,N_8115);
nor U9575 (N_9575,N_8530,N_8914);
nor U9576 (N_9576,N_8779,N_8364);
nor U9577 (N_9577,N_8016,N_8420);
or U9578 (N_9578,N_8961,N_8936);
or U9579 (N_9579,N_8040,N_8599);
or U9580 (N_9580,N_8830,N_8051);
nor U9581 (N_9581,N_8023,N_8966);
nand U9582 (N_9582,N_8997,N_8976);
and U9583 (N_9583,N_8609,N_8288);
and U9584 (N_9584,N_8822,N_8220);
and U9585 (N_9585,N_8752,N_8804);
and U9586 (N_9586,N_8400,N_8169);
nor U9587 (N_9587,N_8112,N_8721);
and U9588 (N_9588,N_8935,N_8527);
xnor U9589 (N_9589,N_8644,N_8256);
and U9590 (N_9590,N_8833,N_8730);
nor U9591 (N_9591,N_8268,N_8717);
nand U9592 (N_9592,N_8811,N_8461);
nor U9593 (N_9593,N_8659,N_8789);
or U9594 (N_9594,N_8359,N_8947);
and U9595 (N_9595,N_8241,N_8177);
nand U9596 (N_9596,N_8282,N_8369);
nand U9597 (N_9597,N_8469,N_8838);
and U9598 (N_9598,N_8170,N_8492);
and U9599 (N_9599,N_8559,N_8751);
or U9600 (N_9600,N_8299,N_8098);
nor U9601 (N_9601,N_8401,N_8795);
or U9602 (N_9602,N_8914,N_8820);
or U9603 (N_9603,N_8213,N_8205);
or U9604 (N_9604,N_8608,N_8112);
or U9605 (N_9605,N_8467,N_8901);
nand U9606 (N_9606,N_8538,N_8534);
nor U9607 (N_9607,N_8081,N_8186);
nor U9608 (N_9608,N_8334,N_8248);
nor U9609 (N_9609,N_8353,N_8514);
nor U9610 (N_9610,N_8144,N_8140);
nand U9611 (N_9611,N_8618,N_8300);
and U9612 (N_9612,N_8117,N_8249);
nand U9613 (N_9613,N_8045,N_8104);
or U9614 (N_9614,N_8322,N_8003);
nand U9615 (N_9615,N_8200,N_8465);
or U9616 (N_9616,N_8203,N_8631);
nand U9617 (N_9617,N_8388,N_8765);
and U9618 (N_9618,N_8592,N_8912);
or U9619 (N_9619,N_8888,N_8104);
or U9620 (N_9620,N_8689,N_8060);
or U9621 (N_9621,N_8473,N_8640);
or U9622 (N_9622,N_8136,N_8799);
and U9623 (N_9623,N_8692,N_8904);
or U9624 (N_9624,N_8276,N_8877);
nor U9625 (N_9625,N_8016,N_8769);
nand U9626 (N_9626,N_8336,N_8449);
or U9627 (N_9627,N_8438,N_8880);
or U9628 (N_9628,N_8181,N_8203);
or U9629 (N_9629,N_8307,N_8234);
or U9630 (N_9630,N_8662,N_8750);
and U9631 (N_9631,N_8304,N_8701);
or U9632 (N_9632,N_8802,N_8084);
and U9633 (N_9633,N_8086,N_8790);
and U9634 (N_9634,N_8259,N_8591);
nor U9635 (N_9635,N_8643,N_8699);
nand U9636 (N_9636,N_8686,N_8849);
or U9637 (N_9637,N_8665,N_8080);
and U9638 (N_9638,N_8940,N_8735);
or U9639 (N_9639,N_8135,N_8859);
or U9640 (N_9640,N_8375,N_8215);
or U9641 (N_9641,N_8523,N_8959);
and U9642 (N_9642,N_8210,N_8423);
and U9643 (N_9643,N_8360,N_8660);
or U9644 (N_9644,N_8634,N_8400);
xnor U9645 (N_9645,N_8778,N_8564);
nand U9646 (N_9646,N_8819,N_8575);
and U9647 (N_9647,N_8857,N_8409);
nand U9648 (N_9648,N_8007,N_8287);
nand U9649 (N_9649,N_8975,N_8682);
or U9650 (N_9650,N_8953,N_8990);
nand U9651 (N_9651,N_8362,N_8990);
or U9652 (N_9652,N_8506,N_8454);
and U9653 (N_9653,N_8333,N_8197);
nand U9654 (N_9654,N_8996,N_8301);
nor U9655 (N_9655,N_8309,N_8063);
nand U9656 (N_9656,N_8301,N_8616);
and U9657 (N_9657,N_8516,N_8423);
nor U9658 (N_9658,N_8195,N_8871);
nor U9659 (N_9659,N_8239,N_8770);
or U9660 (N_9660,N_8359,N_8430);
nor U9661 (N_9661,N_8129,N_8812);
and U9662 (N_9662,N_8876,N_8890);
nor U9663 (N_9663,N_8977,N_8216);
nor U9664 (N_9664,N_8564,N_8398);
and U9665 (N_9665,N_8108,N_8684);
nor U9666 (N_9666,N_8566,N_8081);
and U9667 (N_9667,N_8832,N_8236);
and U9668 (N_9668,N_8871,N_8405);
nor U9669 (N_9669,N_8143,N_8318);
or U9670 (N_9670,N_8963,N_8660);
and U9671 (N_9671,N_8178,N_8565);
nor U9672 (N_9672,N_8219,N_8437);
or U9673 (N_9673,N_8304,N_8190);
nand U9674 (N_9674,N_8707,N_8653);
nor U9675 (N_9675,N_8010,N_8907);
and U9676 (N_9676,N_8482,N_8461);
and U9677 (N_9677,N_8768,N_8729);
or U9678 (N_9678,N_8804,N_8820);
nor U9679 (N_9679,N_8754,N_8068);
nor U9680 (N_9680,N_8083,N_8888);
or U9681 (N_9681,N_8498,N_8964);
and U9682 (N_9682,N_8076,N_8452);
nor U9683 (N_9683,N_8591,N_8442);
and U9684 (N_9684,N_8298,N_8543);
nand U9685 (N_9685,N_8648,N_8708);
or U9686 (N_9686,N_8600,N_8436);
or U9687 (N_9687,N_8196,N_8606);
and U9688 (N_9688,N_8417,N_8733);
nor U9689 (N_9689,N_8102,N_8292);
or U9690 (N_9690,N_8723,N_8431);
nand U9691 (N_9691,N_8735,N_8053);
nand U9692 (N_9692,N_8565,N_8872);
nand U9693 (N_9693,N_8344,N_8305);
nand U9694 (N_9694,N_8401,N_8635);
nand U9695 (N_9695,N_8189,N_8650);
or U9696 (N_9696,N_8291,N_8573);
and U9697 (N_9697,N_8468,N_8549);
nand U9698 (N_9698,N_8658,N_8518);
nor U9699 (N_9699,N_8759,N_8362);
nand U9700 (N_9700,N_8056,N_8149);
nor U9701 (N_9701,N_8144,N_8117);
or U9702 (N_9702,N_8674,N_8634);
nor U9703 (N_9703,N_8267,N_8404);
nand U9704 (N_9704,N_8849,N_8711);
or U9705 (N_9705,N_8040,N_8673);
and U9706 (N_9706,N_8354,N_8261);
or U9707 (N_9707,N_8574,N_8469);
nor U9708 (N_9708,N_8137,N_8686);
nand U9709 (N_9709,N_8857,N_8738);
or U9710 (N_9710,N_8218,N_8103);
or U9711 (N_9711,N_8720,N_8979);
nand U9712 (N_9712,N_8076,N_8757);
or U9713 (N_9713,N_8148,N_8427);
nor U9714 (N_9714,N_8166,N_8680);
or U9715 (N_9715,N_8127,N_8939);
or U9716 (N_9716,N_8316,N_8322);
and U9717 (N_9717,N_8457,N_8146);
nor U9718 (N_9718,N_8308,N_8352);
or U9719 (N_9719,N_8088,N_8811);
or U9720 (N_9720,N_8147,N_8670);
and U9721 (N_9721,N_8400,N_8180);
and U9722 (N_9722,N_8028,N_8420);
and U9723 (N_9723,N_8487,N_8466);
nor U9724 (N_9724,N_8925,N_8409);
nor U9725 (N_9725,N_8782,N_8337);
and U9726 (N_9726,N_8968,N_8465);
nor U9727 (N_9727,N_8356,N_8441);
and U9728 (N_9728,N_8790,N_8018);
or U9729 (N_9729,N_8516,N_8784);
or U9730 (N_9730,N_8875,N_8106);
nor U9731 (N_9731,N_8205,N_8031);
or U9732 (N_9732,N_8461,N_8446);
nand U9733 (N_9733,N_8637,N_8168);
nand U9734 (N_9734,N_8563,N_8954);
nor U9735 (N_9735,N_8654,N_8058);
and U9736 (N_9736,N_8255,N_8019);
nand U9737 (N_9737,N_8945,N_8518);
and U9738 (N_9738,N_8838,N_8676);
nand U9739 (N_9739,N_8037,N_8788);
nor U9740 (N_9740,N_8614,N_8128);
and U9741 (N_9741,N_8198,N_8027);
nor U9742 (N_9742,N_8850,N_8067);
or U9743 (N_9743,N_8929,N_8169);
nor U9744 (N_9744,N_8650,N_8141);
xnor U9745 (N_9745,N_8948,N_8579);
or U9746 (N_9746,N_8461,N_8442);
nor U9747 (N_9747,N_8718,N_8269);
and U9748 (N_9748,N_8281,N_8880);
nor U9749 (N_9749,N_8579,N_8909);
nor U9750 (N_9750,N_8509,N_8361);
nand U9751 (N_9751,N_8233,N_8565);
and U9752 (N_9752,N_8584,N_8473);
or U9753 (N_9753,N_8604,N_8715);
nand U9754 (N_9754,N_8541,N_8638);
nand U9755 (N_9755,N_8349,N_8898);
nand U9756 (N_9756,N_8738,N_8329);
and U9757 (N_9757,N_8372,N_8558);
nand U9758 (N_9758,N_8490,N_8038);
nand U9759 (N_9759,N_8917,N_8750);
and U9760 (N_9760,N_8126,N_8022);
nand U9761 (N_9761,N_8435,N_8949);
nor U9762 (N_9762,N_8286,N_8664);
or U9763 (N_9763,N_8973,N_8120);
nand U9764 (N_9764,N_8917,N_8402);
nor U9765 (N_9765,N_8355,N_8826);
or U9766 (N_9766,N_8281,N_8730);
nor U9767 (N_9767,N_8232,N_8991);
nand U9768 (N_9768,N_8323,N_8742);
and U9769 (N_9769,N_8443,N_8456);
and U9770 (N_9770,N_8676,N_8254);
and U9771 (N_9771,N_8627,N_8954);
or U9772 (N_9772,N_8959,N_8389);
or U9773 (N_9773,N_8879,N_8214);
nand U9774 (N_9774,N_8546,N_8750);
nand U9775 (N_9775,N_8325,N_8813);
nor U9776 (N_9776,N_8345,N_8467);
nand U9777 (N_9777,N_8261,N_8300);
nand U9778 (N_9778,N_8600,N_8709);
nand U9779 (N_9779,N_8959,N_8090);
nand U9780 (N_9780,N_8667,N_8629);
and U9781 (N_9781,N_8042,N_8953);
nand U9782 (N_9782,N_8691,N_8754);
nand U9783 (N_9783,N_8277,N_8122);
nand U9784 (N_9784,N_8604,N_8772);
nand U9785 (N_9785,N_8309,N_8432);
nand U9786 (N_9786,N_8662,N_8336);
nand U9787 (N_9787,N_8268,N_8004);
and U9788 (N_9788,N_8258,N_8433);
nor U9789 (N_9789,N_8993,N_8743);
and U9790 (N_9790,N_8890,N_8953);
nor U9791 (N_9791,N_8552,N_8239);
and U9792 (N_9792,N_8520,N_8828);
and U9793 (N_9793,N_8087,N_8117);
or U9794 (N_9794,N_8911,N_8856);
nand U9795 (N_9795,N_8256,N_8488);
and U9796 (N_9796,N_8259,N_8196);
nor U9797 (N_9797,N_8956,N_8763);
and U9798 (N_9798,N_8350,N_8310);
and U9799 (N_9799,N_8280,N_8179);
nor U9800 (N_9800,N_8560,N_8376);
nor U9801 (N_9801,N_8177,N_8429);
and U9802 (N_9802,N_8190,N_8611);
nor U9803 (N_9803,N_8448,N_8167);
nor U9804 (N_9804,N_8141,N_8714);
nor U9805 (N_9805,N_8968,N_8202);
or U9806 (N_9806,N_8358,N_8573);
nand U9807 (N_9807,N_8937,N_8806);
or U9808 (N_9808,N_8367,N_8402);
or U9809 (N_9809,N_8884,N_8041);
nor U9810 (N_9810,N_8884,N_8684);
nand U9811 (N_9811,N_8506,N_8470);
or U9812 (N_9812,N_8339,N_8972);
nor U9813 (N_9813,N_8345,N_8416);
nand U9814 (N_9814,N_8810,N_8570);
nand U9815 (N_9815,N_8008,N_8767);
nand U9816 (N_9816,N_8146,N_8540);
and U9817 (N_9817,N_8234,N_8629);
or U9818 (N_9818,N_8748,N_8654);
and U9819 (N_9819,N_8051,N_8840);
nor U9820 (N_9820,N_8341,N_8926);
and U9821 (N_9821,N_8501,N_8396);
and U9822 (N_9822,N_8532,N_8142);
nand U9823 (N_9823,N_8449,N_8320);
nor U9824 (N_9824,N_8650,N_8194);
nor U9825 (N_9825,N_8071,N_8789);
nor U9826 (N_9826,N_8374,N_8489);
nor U9827 (N_9827,N_8701,N_8651);
and U9828 (N_9828,N_8037,N_8731);
nand U9829 (N_9829,N_8434,N_8118);
nor U9830 (N_9830,N_8724,N_8473);
and U9831 (N_9831,N_8083,N_8803);
and U9832 (N_9832,N_8433,N_8968);
nor U9833 (N_9833,N_8497,N_8453);
nor U9834 (N_9834,N_8230,N_8373);
nor U9835 (N_9835,N_8615,N_8336);
nor U9836 (N_9836,N_8746,N_8952);
or U9837 (N_9837,N_8651,N_8492);
and U9838 (N_9838,N_8797,N_8587);
and U9839 (N_9839,N_8831,N_8513);
or U9840 (N_9840,N_8608,N_8523);
or U9841 (N_9841,N_8420,N_8654);
or U9842 (N_9842,N_8448,N_8512);
xnor U9843 (N_9843,N_8545,N_8383);
and U9844 (N_9844,N_8298,N_8667);
nand U9845 (N_9845,N_8069,N_8796);
nand U9846 (N_9846,N_8046,N_8042);
and U9847 (N_9847,N_8187,N_8351);
or U9848 (N_9848,N_8918,N_8100);
and U9849 (N_9849,N_8247,N_8725);
and U9850 (N_9850,N_8252,N_8821);
and U9851 (N_9851,N_8212,N_8689);
or U9852 (N_9852,N_8578,N_8877);
nor U9853 (N_9853,N_8326,N_8452);
and U9854 (N_9854,N_8861,N_8323);
or U9855 (N_9855,N_8324,N_8958);
nor U9856 (N_9856,N_8038,N_8960);
or U9857 (N_9857,N_8371,N_8065);
nor U9858 (N_9858,N_8269,N_8335);
and U9859 (N_9859,N_8449,N_8425);
nand U9860 (N_9860,N_8333,N_8314);
and U9861 (N_9861,N_8994,N_8894);
nor U9862 (N_9862,N_8987,N_8165);
nor U9863 (N_9863,N_8994,N_8480);
nand U9864 (N_9864,N_8038,N_8081);
nand U9865 (N_9865,N_8356,N_8866);
or U9866 (N_9866,N_8823,N_8611);
or U9867 (N_9867,N_8418,N_8295);
nand U9868 (N_9868,N_8574,N_8414);
or U9869 (N_9869,N_8577,N_8309);
nor U9870 (N_9870,N_8627,N_8456);
and U9871 (N_9871,N_8533,N_8999);
nor U9872 (N_9872,N_8817,N_8617);
and U9873 (N_9873,N_8109,N_8900);
and U9874 (N_9874,N_8819,N_8092);
or U9875 (N_9875,N_8097,N_8448);
and U9876 (N_9876,N_8907,N_8347);
or U9877 (N_9877,N_8560,N_8129);
or U9878 (N_9878,N_8734,N_8295);
nor U9879 (N_9879,N_8316,N_8040);
and U9880 (N_9880,N_8671,N_8230);
nor U9881 (N_9881,N_8449,N_8081);
and U9882 (N_9882,N_8215,N_8607);
or U9883 (N_9883,N_8700,N_8031);
nor U9884 (N_9884,N_8855,N_8783);
nor U9885 (N_9885,N_8831,N_8172);
nor U9886 (N_9886,N_8713,N_8727);
or U9887 (N_9887,N_8595,N_8415);
and U9888 (N_9888,N_8076,N_8841);
nand U9889 (N_9889,N_8097,N_8916);
and U9890 (N_9890,N_8106,N_8599);
and U9891 (N_9891,N_8195,N_8590);
nor U9892 (N_9892,N_8380,N_8514);
or U9893 (N_9893,N_8605,N_8796);
or U9894 (N_9894,N_8327,N_8755);
and U9895 (N_9895,N_8114,N_8022);
nor U9896 (N_9896,N_8416,N_8147);
or U9897 (N_9897,N_8955,N_8159);
or U9898 (N_9898,N_8818,N_8938);
nor U9899 (N_9899,N_8815,N_8228);
nand U9900 (N_9900,N_8084,N_8379);
and U9901 (N_9901,N_8380,N_8443);
nand U9902 (N_9902,N_8507,N_8691);
or U9903 (N_9903,N_8896,N_8852);
nor U9904 (N_9904,N_8463,N_8732);
nor U9905 (N_9905,N_8720,N_8551);
and U9906 (N_9906,N_8312,N_8023);
nor U9907 (N_9907,N_8554,N_8116);
or U9908 (N_9908,N_8563,N_8195);
or U9909 (N_9909,N_8534,N_8252);
nand U9910 (N_9910,N_8613,N_8622);
or U9911 (N_9911,N_8848,N_8477);
and U9912 (N_9912,N_8783,N_8852);
and U9913 (N_9913,N_8876,N_8459);
nand U9914 (N_9914,N_8845,N_8855);
nor U9915 (N_9915,N_8160,N_8001);
or U9916 (N_9916,N_8667,N_8787);
nand U9917 (N_9917,N_8882,N_8536);
nor U9918 (N_9918,N_8242,N_8183);
and U9919 (N_9919,N_8782,N_8131);
or U9920 (N_9920,N_8446,N_8413);
nand U9921 (N_9921,N_8792,N_8061);
nor U9922 (N_9922,N_8088,N_8201);
nor U9923 (N_9923,N_8801,N_8625);
xnor U9924 (N_9924,N_8518,N_8509);
nand U9925 (N_9925,N_8982,N_8230);
and U9926 (N_9926,N_8192,N_8250);
or U9927 (N_9927,N_8930,N_8869);
nand U9928 (N_9928,N_8038,N_8518);
and U9929 (N_9929,N_8545,N_8996);
nor U9930 (N_9930,N_8781,N_8367);
or U9931 (N_9931,N_8666,N_8312);
nand U9932 (N_9932,N_8405,N_8788);
and U9933 (N_9933,N_8829,N_8469);
and U9934 (N_9934,N_8140,N_8351);
nor U9935 (N_9935,N_8094,N_8101);
nand U9936 (N_9936,N_8382,N_8758);
and U9937 (N_9937,N_8819,N_8462);
or U9938 (N_9938,N_8479,N_8025);
or U9939 (N_9939,N_8051,N_8040);
or U9940 (N_9940,N_8940,N_8456);
or U9941 (N_9941,N_8703,N_8015);
and U9942 (N_9942,N_8844,N_8551);
nand U9943 (N_9943,N_8286,N_8688);
nor U9944 (N_9944,N_8024,N_8666);
or U9945 (N_9945,N_8141,N_8682);
nor U9946 (N_9946,N_8092,N_8543);
nor U9947 (N_9947,N_8656,N_8610);
nand U9948 (N_9948,N_8108,N_8672);
and U9949 (N_9949,N_8595,N_8495);
nand U9950 (N_9950,N_8765,N_8230);
and U9951 (N_9951,N_8273,N_8707);
or U9952 (N_9952,N_8440,N_8549);
nand U9953 (N_9953,N_8280,N_8386);
or U9954 (N_9954,N_8479,N_8497);
nand U9955 (N_9955,N_8814,N_8207);
nor U9956 (N_9956,N_8558,N_8862);
nand U9957 (N_9957,N_8974,N_8980);
nor U9958 (N_9958,N_8069,N_8907);
and U9959 (N_9959,N_8931,N_8687);
and U9960 (N_9960,N_8685,N_8375);
and U9961 (N_9961,N_8902,N_8601);
nand U9962 (N_9962,N_8018,N_8940);
nand U9963 (N_9963,N_8475,N_8681);
nor U9964 (N_9964,N_8131,N_8714);
nor U9965 (N_9965,N_8085,N_8206);
and U9966 (N_9966,N_8637,N_8039);
nand U9967 (N_9967,N_8558,N_8811);
and U9968 (N_9968,N_8793,N_8048);
and U9969 (N_9969,N_8078,N_8751);
nand U9970 (N_9970,N_8140,N_8891);
or U9971 (N_9971,N_8311,N_8998);
nor U9972 (N_9972,N_8309,N_8545);
and U9973 (N_9973,N_8332,N_8840);
nand U9974 (N_9974,N_8979,N_8002);
nor U9975 (N_9975,N_8651,N_8675);
and U9976 (N_9976,N_8669,N_8612);
nand U9977 (N_9977,N_8076,N_8332);
and U9978 (N_9978,N_8731,N_8052);
and U9979 (N_9979,N_8963,N_8288);
nand U9980 (N_9980,N_8241,N_8422);
nand U9981 (N_9981,N_8237,N_8906);
nand U9982 (N_9982,N_8208,N_8353);
or U9983 (N_9983,N_8604,N_8482);
nand U9984 (N_9984,N_8290,N_8752);
nor U9985 (N_9985,N_8141,N_8788);
nor U9986 (N_9986,N_8539,N_8733);
nand U9987 (N_9987,N_8544,N_8703);
and U9988 (N_9988,N_8869,N_8112);
or U9989 (N_9989,N_8902,N_8931);
and U9990 (N_9990,N_8660,N_8173);
or U9991 (N_9991,N_8728,N_8290);
or U9992 (N_9992,N_8186,N_8683);
or U9993 (N_9993,N_8465,N_8649);
nand U9994 (N_9994,N_8611,N_8934);
nand U9995 (N_9995,N_8709,N_8794);
nor U9996 (N_9996,N_8710,N_8390);
and U9997 (N_9997,N_8557,N_8720);
and U9998 (N_9998,N_8928,N_8522);
or U9999 (N_9999,N_8758,N_8041);
nand UO_0 (O_0,N_9137,N_9506);
xnor UO_1 (O_1,N_9654,N_9803);
nand UO_2 (O_2,N_9195,N_9483);
nand UO_3 (O_3,N_9982,N_9517);
nand UO_4 (O_4,N_9797,N_9526);
and UO_5 (O_5,N_9757,N_9868);
or UO_6 (O_6,N_9152,N_9773);
and UO_7 (O_7,N_9366,N_9086);
and UO_8 (O_8,N_9055,N_9261);
or UO_9 (O_9,N_9237,N_9186);
and UO_10 (O_10,N_9156,N_9099);
nor UO_11 (O_11,N_9362,N_9096);
or UO_12 (O_12,N_9000,N_9530);
nor UO_13 (O_13,N_9130,N_9464);
or UO_14 (O_14,N_9848,N_9751);
nor UO_15 (O_15,N_9290,N_9238);
and UO_16 (O_16,N_9396,N_9476);
and UO_17 (O_17,N_9593,N_9004);
or UO_18 (O_18,N_9252,N_9762);
or UO_19 (O_19,N_9535,N_9284);
nor UO_20 (O_20,N_9164,N_9932);
and UO_21 (O_21,N_9841,N_9402);
or UO_22 (O_22,N_9381,N_9222);
and UO_23 (O_23,N_9334,N_9107);
or UO_24 (O_24,N_9155,N_9439);
nor UO_25 (O_25,N_9136,N_9918);
nor UO_26 (O_26,N_9983,N_9764);
xnor UO_27 (O_27,N_9980,N_9962);
or UO_28 (O_28,N_9460,N_9853);
and UO_29 (O_29,N_9830,N_9114);
or UO_30 (O_30,N_9511,N_9303);
nor UO_31 (O_31,N_9015,N_9101);
nand UO_32 (O_32,N_9909,N_9429);
nor UO_33 (O_33,N_9394,N_9815);
or UO_34 (O_34,N_9699,N_9822);
nand UO_35 (O_35,N_9628,N_9153);
and UO_36 (O_36,N_9590,N_9564);
or UO_37 (O_37,N_9727,N_9447);
nand UO_38 (O_38,N_9166,N_9554);
nor UO_39 (O_39,N_9617,N_9251);
and UO_40 (O_40,N_9977,N_9837);
and UO_41 (O_41,N_9972,N_9636);
or UO_42 (O_42,N_9360,N_9952);
or UO_43 (O_43,N_9805,N_9187);
nor UO_44 (O_44,N_9927,N_9142);
nand UO_45 (O_45,N_9071,N_9094);
or UO_46 (O_46,N_9311,N_9813);
or UO_47 (O_47,N_9639,N_9631);
xor UO_48 (O_48,N_9789,N_9198);
or UO_49 (O_49,N_9188,N_9646);
xor UO_50 (O_50,N_9782,N_9452);
nor UO_51 (O_51,N_9512,N_9080);
nand UO_52 (O_52,N_9827,N_9338);
nand UO_53 (O_53,N_9772,N_9201);
or UO_54 (O_54,N_9105,N_9790);
nor UO_55 (O_55,N_9598,N_9759);
or UO_56 (O_56,N_9614,N_9191);
nand UO_57 (O_57,N_9482,N_9272);
xor UO_58 (O_58,N_9708,N_9148);
nor UO_59 (O_59,N_9702,N_9093);
and UO_60 (O_60,N_9075,N_9392);
or UO_61 (O_61,N_9776,N_9951);
or UO_62 (O_62,N_9008,N_9994);
or UO_63 (O_63,N_9390,N_9557);
and UO_64 (O_64,N_9486,N_9926);
nand UO_65 (O_65,N_9942,N_9165);
nand UO_66 (O_66,N_9532,N_9622);
and UO_67 (O_67,N_9050,N_9062);
and UO_68 (O_68,N_9289,N_9795);
or UO_69 (O_69,N_9224,N_9042);
nor UO_70 (O_70,N_9601,N_9019);
nand UO_71 (O_71,N_9905,N_9052);
nor UO_72 (O_72,N_9258,N_9022);
and UO_73 (O_73,N_9280,N_9967);
nor UO_74 (O_74,N_9240,N_9007);
or UO_75 (O_75,N_9997,N_9732);
and UO_76 (O_76,N_9014,N_9920);
and UO_77 (O_77,N_9600,N_9016);
nand UO_78 (O_78,N_9663,N_9190);
and UO_79 (O_79,N_9612,N_9767);
or UO_80 (O_80,N_9722,N_9957);
nand UO_81 (O_81,N_9527,N_9226);
or UO_82 (O_82,N_9545,N_9441);
nand UO_83 (O_83,N_9878,N_9494);
nand UO_84 (O_84,N_9978,N_9281);
nand UO_85 (O_85,N_9881,N_9481);
or UO_86 (O_86,N_9265,N_9753);
nand UO_87 (O_87,N_9750,N_9455);
and UO_88 (O_88,N_9876,N_9843);
xor UO_89 (O_89,N_9321,N_9346);
nand UO_90 (O_90,N_9021,N_9863);
or UO_91 (O_91,N_9632,N_9254);
or UO_92 (O_92,N_9048,N_9537);
or UO_93 (O_93,N_9589,N_9037);
nand UO_94 (O_94,N_9500,N_9010);
and UO_95 (O_95,N_9747,N_9673);
nand UO_96 (O_96,N_9451,N_9293);
and UO_97 (O_97,N_9903,N_9309);
xnor UO_98 (O_98,N_9566,N_9703);
nor UO_99 (O_99,N_9748,N_9461);
nand UO_100 (O_100,N_9971,N_9112);
nor UO_101 (O_101,N_9718,N_9051);
nand UO_102 (O_102,N_9276,N_9418);
nor UO_103 (O_103,N_9414,N_9974);
xnor UO_104 (O_104,N_9596,N_9448);
and UO_105 (O_105,N_9259,N_9406);
and UO_106 (O_106,N_9488,N_9074);
and UO_107 (O_107,N_9572,N_9552);
nand UO_108 (O_108,N_9754,N_9315);
nor UO_109 (O_109,N_9111,N_9801);
nor UO_110 (O_110,N_9056,N_9956);
nand UO_111 (O_111,N_9743,N_9161);
xor UO_112 (O_112,N_9025,N_9473);
nor UO_113 (O_113,N_9941,N_9549);
nand UO_114 (O_114,N_9917,N_9219);
and UO_115 (O_115,N_9064,N_9091);
and UO_116 (O_116,N_9648,N_9807);
nand UO_117 (O_117,N_9966,N_9301);
nor UO_118 (O_118,N_9349,N_9756);
or UO_119 (O_119,N_9355,N_9854);
nor UO_120 (O_120,N_9298,N_9277);
nand UO_121 (O_121,N_9594,N_9129);
nor UO_122 (O_122,N_9297,N_9784);
and UO_123 (O_123,N_9291,N_9149);
and UO_124 (O_124,N_9162,N_9913);
nor UO_125 (O_125,N_9811,N_9018);
or UO_126 (O_126,N_9210,N_9735);
nand UO_127 (O_127,N_9002,N_9515);
and UO_128 (O_128,N_9844,N_9432);
nand UO_129 (O_129,N_9307,N_9629);
and UO_130 (O_130,N_9824,N_9911);
or UO_131 (O_131,N_9178,N_9683);
and UO_132 (O_132,N_9860,N_9711);
nand UO_133 (O_133,N_9437,N_9504);
nand UO_134 (O_134,N_9634,N_9568);
or UO_135 (O_135,N_9215,N_9543);
nor UO_136 (O_136,N_9656,N_9832);
nand UO_137 (O_137,N_9184,N_9235);
nor UO_138 (O_138,N_9935,N_9603);
or UO_139 (O_139,N_9279,N_9369);
and UO_140 (O_140,N_9657,N_9700);
or UO_141 (O_141,N_9624,N_9046);
or UO_142 (O_142,N_9724,N_9275);
or UO_143 (O_143,N_9938,N_9078);
and UO_144 (O_144,N_9694,N_9299);
and UO_145 (O_145,N_9828,N_9351);
or UO_146 (O_146,N_9542,N_9412);
and UO_147 (O_147,N_9095,N_9409);
or UO_148 (O_148,N_9523,N_9793);
or UO_149 (O_149,N_9847,N_9550);
or UO_150 (O_150,N_9809,N_9034);
and UO_151 (O_151,N_9682,N_9933);
and UO_152 (O_152,N_9779,N_9092);
nor UO_153 (O_153,N_9625,N_9599);
and UO_154 (O_154,N_9380,N_9892);
and UO_155 (O_155,N_9256,N_9692);
nor UO_156 (O_156,N_9852,N_9395);
nor UO_157 (O_157,N_9497,N_9131);
nor UO_158 (O_158,N_9430,N_9884);
or UO_159 (O_159,N_9348,N_9840);
nor UO_160 (O_160,N_9508,N_9384);
or UO_161 (O_161,N_9431,N_9028);
nor UO_162 (O_162,N_9842,N_9116);
nor UO_163 (O_163,N_9262,N_9559);
or UO_164 (O_164,N_9322,N_9889);
nand UO_165 (O_165,N_9835,N_9049);
nor UO_166 (O_166,N_9317,N_9378);
nor UO_167 (O_167,N_9740,N_9333);
or UO_168 (O_168,N_9861,N_9035);
and UO_169 (O_169,N_9039,N_9465);
or UO_170 (O_170,N_9491,N_9658);
and UO_171 (O_171,N_9709,N_9085);
nand UO_172 (O_172,N_9838,N_9405);
nor UO_173 (O_173,N_9577,N_9819);
nand UO_174 (O_174,N_9791,N_9563);
and UO_175 (O_175,N_9020,N_9653);
and UO_176 (O_176,N_9415,N_9084);
and UO_177 (O_177,N_9584,N_9520);
nor UO_178 (O_178,N_9937,N_9234);
or UO_179 (O_179,N_9597,N_9168);
or UO_180 (O_180,N_9283,N_9505);
nand UO_181 (O_181,N_9312,N_9613);
nor UO_182 (O_182,N_9385,N_9193);
nand UO_183 (O_183,N_9218,N_9744);
and UO_184 (O_184,N_9273,N_9175);
and UO_185 (O_185,N_9445,N_9282);
xor UO_186 (O_186,N_9278,N_9398);
or UO_187 (O_187,N_9522,N_9531);
or UO_188 (O_188,N_9133,N_9534);
nor UO_189 (O_189,N_9851,N_9672);
or UO_190 (O_190,N_9661,N_9245);
and UO_191 (O_191,N_9839,N_9888);
or UO_192 (O_192,N_9898,N_9367);
and UO_193 (O_193,N_9436,N_9516);
nand UO_194 (O_194,N_9825,N_9729);
nor UO_195 (O_195,N_9124,N_9857);
nor UO_196 (O_196,N_9352,N_9691);
nor UO_197 (O_197,N_9061,N_9060);
and UO_198 (O_198,N_9850,N_9407);
and UO_199 (O_199,N_9490,N_9814);
or UO_200 (O_200,N_9045,N_9070);
and UO_201 (O_201,N_9587,N_9944);
nor UO_202 (O_202,N_9003,N_9976);
nor UO_203 (O_203,N_9796,N_9501);
or UO_204 (O_204,N_9287,N_9553);
nor UO_205 (O_205,N_9777,N_9640);
and UO_206 (O_206,N_9033,N_9211);
and UO_207 (O_207,N_9371,N_9263);
and UO_208 (O_208,N_9013,N_9248);
nor UO_209 (O_209,N_9377,N_9698);
nand UO_210 (O_210,N_9975,N_9109);
nor UO_211 (O_211,N_9102,N_9768);
nor UO_212 (O_212,N_9173,N_9474);
nor UO_213 (O_213,N_9221,N_9569);
or UO_214 (O_214,N_9949,N_9931);
and UO_215 (O_215,N_9986,N_9059);
nor UO_216 (O_216,N_9958,N_9073);
or UO_217 (O_217,N_9330,N_9710);
or UO_218 (O_218,N_9410,N_9450);
or UO_219 (O_219,N_9869,N_9134);
and UO_220 (O_220,N_9030,N_9400);
nand UO_221 (O_221,N_9706,N_9484);
nand UO_222 (O_222,N_9328,N_9444);
xor UO_223 (O_223,N_9538,N_9507);
or UO_224 (O_224,N_9110,N_9433);
or UO_225 (O_225,N_9424,N_9582);
or UO_226 (O_226,N_9189,N_9097);
nor UO_227 (O_227,N_9734,N_9741);
nor UO_228 (O_228,N_9585,N_9979);
and UO_229 (O_229,N_9233,N_9896);
and UO_230 (O_230,N_9462,N_9890);
nand UO_231 (O_231,N_9181,N_9364);
nor UO_232 (O_232,N_9468,N_9466);
nor UO_233 (O_233,N_9286,N_9638);
nand UO_234 (O_234,N_9547,N_9054);
or UO_235 (O_235,N_9725,N_9821);
and UO_236 (O_236,N_9574,N_9514);
nor UO_237 (O_237,N_9150,N_9715);
nor UO_238 (O_238,N_9040,N_9082);
and UO_239 (O_239,N_9172,N_9992);
or UO_240 (O_240,N_9655,N_9713);
nor UO_241 (O_241,N_9313,N_9780);
or UO_242 (O_242,N_9183,N_9800);
or UO_243 (O_243,N_9669,N_9339);
or UO_244 (O_244,N_9208,N_9649);
or UO_245 (O_245,N_9470,N_9608);
or UO_246 (O_246,N_9001,N_9088);
and UO_247 (O_247,N_9714,N_9588);
and UO_248 (O_248,N_9945,N_9140);
nand UO_249 (O_249,N_9319,N_9241);
and UO_250 (O_250,N_9122,N_9968);
and UO_251 (O_251,N_9176,N_9539);
nand UO_252 (O_252,N_9242,N_9038);
nor UO_253 (O_253,N_9232,N_9739);
nor UO_254 (O_254,N_9117,N_9266);
nand UO_255 (O_255,N_9645,N_9174);
or UO_256 (O_256,N_9633,N_9372);
or UO_257 (O_257,N_9618,N_9425);
nand UO_258 (O_258,N_9368,N_9864);
nand UO_259 (O_259,N_9318,N_9225);
and UO_260 (O_260,N_9916,N_9914);
or UO_261 (O_261,N_9387,N_9337);
and UO_262 (O_262,N_9434,N_9342);
or UO_263 (O_263,N_9580,N_9223);
and UO_264 (O_264,N_9695,N_9943);
nor UO_265 (O_265,N_9463,N_9145);
nor UO_266 (O_266,N_9244,N_9866);
nor UO_267 (O_267,N_9128,N_9728);
or UO_268 (O_268,N_9677,N_9697);
or UO_269 (O_269,N_9712,N_9806);
or UO_270 (O_270,N_9960,N_9067);
or UO_271 (O_271,N_9573,N_9182);
and UO_272 (O_272,N_9493,N_9820);
or UO_273 (O_273,N_9404,N_9026);
nand UO_274 (O_274,N_9216,N_9373);
and UO_275 (O_275,N_9834,N_9185);
and UO_276 (O_276,N_9637,N_9375);
or UO_277 (O_277,N_9125,N_9421);
and UO_278 (O_278,N_9023,N_9925);
or UO_279 (O_279,N_9964,N_9212);
nand UO_280 (O_280,N_9954,N_9544);
nor UO_281 (O_281,N_9716,N_9749);
nand UO_282 (O_282,N_9541,N_9320);
nand UO_283 (O_283,N_9723,N_9356);
nand UO_284 (O_284,N_9344,N_9867);
nand UO_285 (O_285,N_9341,N_9477);
and UO_286 (O_286,N_9770,N_9882);
nor UO_287 (O_287,N_9704,N_9886);
nand UO_288 (O_288,N_9146,N_9171);
and UO_289 (O_289,N_9157,N_9906);
nand UO_290 (O_290,N_9009,N_9108);
nand UO_291 (O_291,N_9816,N_9332);
and UO_292 (O_292,N_9879,N_9808);
or UO_293 (O_293,N_9257,N_9422);
nand UO_294 (O_294,N_9900,N_9480);
and UO_295 (O_295,N_9467,N_9336);
or UO_296 (O_296,N_9591,N_9119);
nand UO_297 (O_297,N_9662,N_9269);
and UO_298 (O_298,N_9670,N_9382);
or UO_299 (O_299,N_9169,N_9115);
and UO_300 (O_300,N_9685,N_9688);
or UO_301 (O_301,N_9684,N_9681);
nand UO_302 (O_302,N_9781,N_9664);
and UO_303 (O_303,N_9922,N_9737);
nor UO_304 (O_304,N_9546,N_9401);
nand UO_305 (O_305,N_9676,N_9548);
nor UO_306 (O_306,N_9746,N_9154);
and UO_307 (O_307,N_9357,N_9274);
and UO_308 (O_308,N_9250,N_9316);
or UO_309 (O_309,N_9570,N_9817);
or UO_310 (O_310,N_9217,N_9090);
or UO_311 (O_311,N_9874,N_9024);
nand UO_312 (O_312,N_9123,N_9209);
nand UO_313 (O_313,N_9934,N_9571);
nor UO_314 (O_314,N_9620,N_9408);
nor UO_315 (O_315,N_9365,N_9939);
nor UO_316 (O_316,N_9132,N_9243);
or UO_317 (O_317,N_9413,N_9138);
or UO_318 (O_318,N_9619,N_9098);
or UO_319 (O_319,N_9717,N_9229);
nand UO_320 (O_320,N_9032,N_9127);
or UO_321 (O_321,N_9651,N_9513);
nand UO_322 (O_322,N_9205,N_9556);
and UO_323 (O_323,N_9325,N_9794);
nor UO_324 (O_324,N_9005,N_9893);
nand UO_325 (O_325,N_9919,N_9446);
and UO_326 (O_326,N_9475,N_9668);
or UO_327 (O_327,N_9948,N_9247);
nor UO_328 (O_328,N_9731,N_9765);
and UO_329 (O_329,N_9858,N_9973);
nand UO_330 (O_330,N_9044,N_9253);
nand UO_331 (O_331,N_9575,N_9990);
nor UO_332 (O_332,N_9089,N_9562);
and UO_333 (O_333,N_9924,N_9053);
nor UO_334 (O_334,N_9350,N_9179);
and UO_335 (O_335,N_9626,N_9726);
nand UO_336 (O_336,N_9885,N_9420);
nand UO_337 (O_337,N_9862,N_9996);
nand UO_338 (O_338,N_9100,N_9907);
or UO_339 (O_339,N_9989,N_9343);
or UO_340 (O_340,N_9578,N_9659);
and UO_341 (O_341,N_9823,N_9077);
nor UO_342 (O_342,N_9383,N_9592);
or UO_343 (O_343,N_9228,N_9775);
and UO_344 (O_344,N_9160,N_9103);
and UO_345 (O_345,N_9891,N_9623);
nand UO_346 (O_346,N_9999,N_9567);
nor UO_347 (O_347,N_9031,N_9981);
nand UO_348 (O_348,N_9915,N_9170);
or UO_349 (O_349,N_9324,N_9529);
or UO_350 (O_350,N_9167,N_9388);
nor UO_351 (O_351,N_9194,N_9458);
nand UO_352 (O_352,N_9783,N_9533);
nand UO_353 (O_353,N_9985,N_9177);
and UO_354 (O_354,N_9908,N_9605);
nand UO_355 (O_355,N_9586,N_9802);
nand UO_356 (O_356,N_9029,N_9988);
nor UO_357 (O_357,N_9519,N_9921);
nor UO_358 (O_358,N_9652,N_9812);
or UO_359 (O_359,N_9666,N_9068);
or UO_360 (O_360,N_9141,N_9428);
nand UO_361 (O_361,N_9611,N_9471);
nor UO_362 (O_362,N_9701,N_9163);
or UO_363 (O_363,N_9883,N_9399);
nand UO_364 (O_364,N_9158,N_9329);
nor UO_365 (O_365,N_9113,N_9359);
and UO_366 (O_366,N_9180,N_9846);
nor UO_367 (O_367,N_9833,N_9423);
nand UO_368 (O_368,N_9144,N_9302);
nand UO_369 (O_369,N_9327,N_9650);
or UO_370 (O_370,N_9310,N_9370);
or UO_371 (O_371,N_9454,N_9561);
and UO_372 (O_372,N_9788,N_9427);
nand UO_373 (O_373,N_9345,N_9831);
nor UO_374 (O_374,N_9435,N_9300);
nor UO_375 (O_375,N_9079,N_9540);
and UO_376 (O_376,N_9705,N_9785);
nor UO_377 (O_377,N_9621,N_9720);
nand UO_378 (O_378,N_9304,N_9606);
nor UO_379 (O_379,N_9207,N_9761);
or UO_380 (O_380,N_9707,N_9192);
and UO_381 (O_381,N_9680,N_9678);
or UO_382 (O_382,N_9875,N_9950);
or UO_383 (O_383,N_9616,N_9897);
xor UO_384 (O_384,N_9438,N_9871);
nor UO_385 (O_385,N_9442,N_9870);
nand UO_386 (O_386,N_9696,N_9689);
nor UO_387 (O_387,N_9058,N_9353);
or UO_388 (O_388,N_9495,N_9758);
and UO_389 (O_389,N_9912,N_9607);
nor UO_390 (O_390,N_9923,N_9528);
or UO_391 (O_391,N_9928,N_9376);
or UO_392 (O_392,N_9104,N_9693);
nand UO_393 (O_393,N_9766,N_9206);
and UO_394 (O_394,N_9270,N_9118);
nand UO_395 (O_395,N_9011,N_9826);
nor UO_396 (O_396,N_9347,N_9041);
nor UO_397 (O_397,N_9499,N_9798);
and UO_398 (O_398,N_9610,N_9260);
or UO_399 (O_399,N_9296,N_9733);
and UO_400 (O_400,N_9991,N_9403);
or UO_401 (O_401,N_9560,N_9271);
or UO_402 (O_402,N_9873,N_9760);
nand UO_403 (O_403,N_9331,N_9419);
nor UO_404 (O_404,N_9472,N_9081);
nor UO_405 (O_405,N_9391,N_9036);
nand UO_406 (O_406,N_9393,N_9417);
or UO_407 (O_407,N_9609,N_9308);
nand UO_408 (O_408,N_9076,N_9295);
or UO_409 (O_409,N_9083,N_9630);
nor UO_410 (O_410,N_9066,N_9679);
or UO_411 (O_411,N_9660,N_9965);
nand UO_412 (O_412,N_9521,N_9810);
nand UO_413 (O_413,N_9214,N_9121);
nor UO_414 (O_414,N_9249,N_9671);
nand UO_415 (O_415,N_9143,N_9065);
nor UO_416 (O_416,N_9635,N_9665);
nor UO_417 (O_417,N_9456,N_9604);
nor UO_418 (O_418,N_9895,N_9006);
or UO_419 (O_419,N_9440,N_9936);
and UO_420 (O_420,N_9643,N_9910);
nor UO_421 (O_421,N_9998,N_9755);
and UO_422 (O_422,N_9738,N_9363);
nor UO_423 (O_423,N_9930,N_9786);
or UO_424 (O_424,N_9970,N_9953);
nor UO_425 (O_425,N_9929,N_9774);
and UO_426 (O_426,N_9872,N_9220);
and UO_427 (O_427,N_9583,N_9675);
nor UO_428 (O_428,N_9374,N_9294);
and UO_429 (O_429,N_9959,N_9642);
nand UO_430 (O_430,N_9306,N_9993);
or UO_431 (O_431,N_9536,N_9641);
or UO_432 (O_432,N_9027,N_9126);
and UO_433 (O_433,N_9057,N_9203);
nand UO_434 (O_434,N_9961,N_9865);
nand UO_435 (O_435,N_9196,N_9147);
and UO_436 (O_436,N_9855,N_9836);
nor UO_437 (O_437,N_9799,N_9135);
nor UO_438 (O_438,N_9443,N_9627);
and UO_439 (O_439,N_9305,N_9644);
or UO_440 (O_440,N_9719,N_9487);
nand UO_441 (O_441,N_9213,N_9667);
nand UO_442 (O_442,N_9845,N_9752);
nor UO_443 (O_443,N_9969,N_9687);
nand UO_444 (O_444,N_9120,N_9730);
or UO_445 (O_445,N_9106,N_9769);
and UO_446 (O_446,N_9877,N_9524);
and UO_447 (O_447,N_9230,N_9314);
nand UO_448 (O_448,N_9904,N_9047);
nor UO_449 (O_449,N_9901,N_9063);
or UO_450 (O_450,N_9498,N_9416);
nor UO_451 (O_451,N_9647,N_9984);
or UO_452 (O_452,N_9072,N_9457);
or UO_453 (O_453,N_9227,N_9518);
nand UO_454 (O_454,N_9721,N_9255);
or UO_455 (O_455,N_9231,N_9579);
nand UO_456 (O_456,N_9995,N_9340);
or UO_457 (O_457,N_9239,N_9576);
xnor UO_458 (O_458,N_9288,N_9887);
nor UO_459 (O_459,N_9829,N_9818);
nand UO_460 (O_460,N_9742,N_9268);
and UO_461 (O_461,N_9947,N_9354);
or UO_462 (O_462,N_9389,N_9469);
nand UO_463 (O_463,N_9686,N_9489);
or UO_464 (O_464,N_9894,N_9602);
nand UO_465 (O_465,N_9987,N_9449);
nor UO_466 (O_466,N_9386,N_9478);
or UO_467 (O_467,N_9940,N_9361);
nor UO_468 (O_468,N_9763,N_9151);
nor UO_469 (O_469,N_9787,N_9479);
nand UO_470 (O_470,N_9017,N_9012);
xnor UO_471 (O_471,N_9323,N_9555);
xor UO_472 (O_472,N_9411,N_9880);
and UO_473 (O_473,N_9264,N_9856);
and UO_474 (O_474,N_9043,N_9551);
nand UO_475 (O_475,N_9236,N_9335);
nand UO_476 (O_476,N_9963,N_9565);
nor UO_477 (O_477,N_9902,N_9946);
nand UO_478 (O_478,N_9859,N_9492);
nor UO_479 (O_479,N_9139,N_9246);
or UO_480 (O_480,N_9200,N_9379);
or UO_481 (O_481,N_9771,N_9804);
nor UO_482 (O_482,N_9899,N_9087);
nand UO_483 (O_483,N_9690,N_9267);
or UO_484 (O_484,N_9496,N_9581);
nand UO_485 (O_485,N_9502,N_9453);
nand UO_486 (O_486,N_9326,N_9397);
nor UO_487 (O_487,N_9292,N_9674);
or UO_488 (O_488,N_9736,N_9202);
or UO_489 (O_489,N_9778,N_9485);
or UO_490 (O_490,N_9197,N_9510);
nand UO_491 (O_491,N_9525,N_9503);
nor UO_492 (O_492,N_9849,N_9459);
or UO_493 (O_493,N_9509,N_9792);
and UO_494 (O_494,N_9745,N_9204);
nor UO_495 (O_495,N_9285,N_9199);
or UO_496 (O_496,N_9595,N_9069);
nand UO_497 (O_497,N_9426,N_9558);
or UO_498 (O_498,N_9955,N_9615);
or UO_499 (O_499,N_9358,N_9159);
and UO_500 (O_500,N_9650,N_9039);
or UO_501 (O_501,N_9919,N_9769);
or UO_502 (O_502,N_9412,N_9791);
or UO_503 (O_503,N_9872,N_9186);
nand UO_504 (O_504,N_9315,N_9038);
nor UO_505 (O_505,N_9987,N_9782);
nor UO_506 (O_506,N_9993,N_9443);
nand UO_507 (O_507,N_9905,N_9389);
or UO_508 (O_508,N_9809,N_9726);
nand UO_509 (O_509,N_9727,N_9709);
or UO_510 (O_510,N_9610,N_9041);
and UO_511 (O_511,N_9402,N_9423);
and UO_512 (O_512,N_9411,N_9247);
nor UO_513 (O_513,N_9556,N_9417);
nor UO_514 (O_514,N_9449,N_9617);
or UO_515 (O_515,N_9792,N_9973);
or UO_516 (O_516,N_9370,N_9077);
and UO_517 (O_517,N_9829,N_9203);
nand UO_518 (O_518,N_9041,N_9425);
nand UO_519 (O_519,N_9312,N_9060);
nor UO_520 (O_520,N_9723,N_9682);
or UO_521 (O_521,N_9990,N_9386);
or UO_522 (O_522,N_9608,N_9939);
or UO_523 (O_523,N_9510,N_9333);
nor UO_524 (O_524,N_9008,N_9118);
or UO_525 (O_525,N_9566,N_9381);
nor UO_526 (O_526,N_9452,N_9225);
or UO_527 (O_527,N_9844,N_9945);
and UO_528 (O_528,N_9706,N_9991);
nand UO_529 (O_529,N_9379,N_9766);
nand UO_530 (O_530,N_9211,N_9167);
nand UO_531 (O_531,N_9750,N_9768);
nor UO_532 (O_532,N_9569,N_9823);
and UO_533 (O_533,N_9398,N_9284);
or UO_534 (O_534,N_9556,N_9144);
xnor UO_535 (O_535,N_9582,N_9091);
and UO_536 (O_536,N_9092,N_9838);
or UO_537 (O_537,N_9216,N_9387);
nor UO_538 (O_538,N_9138,N_9870);
and UO_539 (O_539,N_9508,N_9847);
nor UO_540 (O_540,N_9799,N_9467);
or UO_541 (O_541,N_9361,N_9014);
or UO_542 (O_542,N_9469,N_9844);
and UO_543 (O_543,N_9965,N_9601);
nor UO_544 (O_544,N_9039,N_9296);
and UO_545 (O_545,N_9829,N_9265);
nor UO_546 (O_546,N_9270,N_9670);
or UO_547 (O_547,N_9937,N_9851);
and UO_548 (O_548,N_9858,N_9648);
nand UO_549 (O_549,N_9450,N_9247);
or UO_550 (O_550,N_9121,N_9748);
nand UO_551 (O_551,N_9236,N_9275);
or UO_552 (O_552,N_9726,N_9831);
and UO_553 (O_553,N_9388,N_9599);
nor UO_554 (O_554,N_9699,N_9823);
nand UO_555 (O_555,N_9976,N_9226);
nor UO_556 (O_556,N_9791,N_9159);
nor UO_557 (O_557,N_9864,N_9601);
nand UO_558 (O_558,N_9492,N_9312);
nor UO_559 (O_559,N_9408,N_9668);
nor UO_560 (O_560,N_9350,N_9537);
and UO_561 (O_561,N_9825,N_9036);
and UO_562 (O_562,N_9587,N_9467);
nand UO_563 (O_563,N_9826,N_9516);
or UO_564 (O_564,N_9430,N_9303);
and UO_565 (O_565,N_9182,N_9658);
nor UO_566 (O_566,N_9243,N_9644);
nor UO_567 (O_567,N_9380,N_9968);
nor UO_568 (O_568,N_9171,N_9084);
nor UO_569 (O_569,N_9024,N_9582);
nor UO_570 (O_570,N_9808,N_9916);
nor UO_571 (O_571,N_9009,N_9912);
nor UO_572 (O_572,N_9604,N_9809);
nand UO_573 (O_573,N_9846,N_9515);
and UO_574 (O_574,N_9379,N_9300);
nor UO_575 (O_575,N_9834,N_9411);
nand UO_576 (O_576,N_9819,N_9013);
nor UO_577 (O_577,N_9889,N_9019);
or UO_578 (O_578,N_9395,N_9682);
or UO_579 (O_579,N_9471,N_9035);
and UO_580 (O_580,N_9681,N_9354);
nand UO_581 (O_581,N_9914,N_9182);
or UO_582 (O_582,N_9557,N_9931);
nand UO_583 (O_583,N_9463,N_9683);
or UO_584 (O_584,N_9236,N_9034);
nand UO_585 (O_585,N_9258,N_9144);
or UO_586 (O_586,N_9022,N_9602);
xnor UO_587 (O_587,N_9194,N_9916);
nor UO_588 (O_588,N_9685,N_9548);
and UO_589 (O_589,N_9666,N_9808);
or UO_590 (O_590,N_9153,N_9194);
or UO_591 (O_591,N_9662,N_9365);
and UO_592 (O_592,N_9616,N_9240);
nor UO_593 (O_593,N_9914,N_9165);
or UO_594 (O_594,N_9427,N_9071);
and UO_595 (O_595,N_9030,N_9159);
and UO_596 (O_596,N_9774,N_9095);
or UO_597 (O_597,N_9126,N_9558);
nand UO_598 (O_598,N_9659,N_9922);
nor UO_599 (O_599,N_9034,N_9950);
nand UO_600 (O_600,N_9998,N_9449);
nand UO_601 (O_601,N_9367,N_9591);
nand UO_602 (O_602,N_9559,N_9355);
nor UO_603 (O_603,N_9427,N_9851);
or UO_604 (O_604,N_9121,N_9681);
nor UO_605 (O_605,N_9344,N_9489);
nand UO_606 (O_606,N_9817,N_9522);
nand UO_607 (O_607,N_9992,N_9455);
nor UO_608 (O_608,N_9127,N_9344);
and UO_609 (O_609,N_9983,N_9517);
nand UO_610 (O_610,N_9756,N_9735);
nand UO_611 (O_611,N_9036,N_9211);
nor UO_612 (O_612,N_9184,N_9649);
nand UO_613 (O_613,N_9066,N_9437);
or UO_614 (O_614,N_9380,N_9782);
nand UO_615 (O_615,N_9128,N_9104);
or UO_616 (O_616,N_9941,N_9674);
nand UO_617 (O_617,N_9215,N_9442);
and UO_618 (O_618,N_9318,N_9003);
or UO_619 (O_619,N_9074,N_9894);
nand UO_620 (O_620,N_9312,N_9218);
nor UO_621 (O_621,N_9630,N_9017);
and UO_622 (O_622,N_9010,N_9355);
and UO_623 (O_623,N_9398,N_9464);
nand UO_624 (O_624,N_9555,N_9520);
nand UO_625 (O_625,N_9937,N_9223);
xor UO_626 (O_626,N_9887,N_9504);
or UO_627 (O_627,N_9230,N_9239);
and UO_628 (O_628,N_9038,N_9693);
and UO_629 (O_629,N_9479,N_9543);
nor UO_630 (O_630,N_9699,N_9878);
nand UO_631 (O_631,N_9239,N_9636);
or UO_632 (O_632,N_9871,N_9275);
nor UO_633 (O_633,N_9635,N_9973);
nor UO_634 (O_634,N_9107,N_9394);
nand UO_635 (O_635,N_9923,N_9207);
or UO_636 (O_636,N_9678,N_9131);
or UO_637 (O_637,N_9125,N_9849);
nand UO_638 (O_638,N_9874,N_9438);
nor UO_639 (O_639,N_9696,N_9244);
and UO_640 (O_640,N_9833,N_9087);
nand UO_641 (O_641,N_9485,N_9355);
nor UO_642 (O_642,N_9248,N_9733);
nor UO_643 (O_643,N_9065,N_9505);
nor UO_644 (O_644,N_9549,N_9761);
or UO_645 (O_645,N_9127,N_9664);
xnor UO_646 (O_646,N_9772,N_9288);
nor UO_647 (O_647,N_9368,N_9923);
xnor UO_648 (O_648,N_9124,N_9146);
and UO_649 (O_649,N_9346,N_9901);
and UO_650 (O_650,N_9241,N_9687);
nor UO_651 (O_651,N_9325,N_9209);
nand UO_652 (O_652,N_9798,N_9548);
nor UO_653 (O_653,N_9775,N_9897);
nand UO_654 (O_654,N_9740,N_9430);
and UO_655 (O_655,N_9469,N_9374);
nor UO_656 (O_656,N_9938,N_9615);
nor UO_657 (O_657,N_9328,N_9514);
and UO_658 (O_658,N_9875,N_9887);
and UO_659 (O_659,N_9829,N_9938);
xnor UO_660 (O_660,N_9149,N_9839);
nand UO_661 (O_661,N_9567,N_9090);
nor UO_662 (O_662,N_9579,N_9239);
nor UO_663 (O_663,N_9756,N_9880);
nor UO_664 (O_664,N_9690,N_9401);
and UO_665 (O_665,N_9803,N_9501);
nor UO_666 (O_666,N_9965,N_9093);
or UO_667 (O_667,N_9730,N_9287);
nor UO_668 (O_668,N_9367,N_9919);
and UO_669 (O_669,N_9620,N_9773);
nand UO_670 (O_670,N_9320,N_9993);
and UO_671 (O_671,N_9123,N_9537);
and UO_672 (O_672,N_9313,N_9103);
nand UO_673 (O_673,N_9462,N_9256);
and UO_674 (O_674,N_9574,N_9195);
or UO_675 (O_675,N_9642,N_9494);
nor UO_676 (O_676,N_9777,N_9228);
or UO_677 (O_677,N_9515,N_9276);
nor UO_678 (O_678,N_9367,N_9490);
nand UO_679 (O_679,N_9686,N_9020);
nand UO_680 (O_680,N_9084,N_9668);
nor UO_681 (O_681,N_9899,N_9656);
and UO_682 (O_682,N_9531,N_9809);
nand UO_683 (O_683,N_9156,N_9608);
or UO_684 (O_684,N_9621,N_9198);
and UO_685 (O_685,N_9542,N_9789);
and UO_686 (O_686,N_9757,N_9706);
or UO_687 (O_687,N_9658,N_9846);
nor UO_688 (O_688,N_9503,N_9963);
or UO_689 (O_689,N_9615,N_9631);
nand UO_690 (O_690,N_9495,N_9795);
nor UO_691 (O_691,N_9707,N_9227);
nor UO_692 (O_692,N_9560,N_9728);
nand UO_693 (O_693,N_9346,N_9532);
nand UO_694 (O_694,N_9377,N_9785);
and UO_695 (O_695,N_9379,N_9227);
or UO_696 (O_696,N_9050,N_9782);
and UO_697 (O_697,N_9774,N_9062);
or UO_698 (O_698,N_9197,N_9962);
nand UO_699 (O_699,N_9880,N_9083);
and UO_700 (O_700,N_9966,N_9981);
or UO_701 (O_701,N_9642,N_9817);
nand UO_702 (O_702,N_9994,N_9758);
nand UO_703 (O_703,N_9024,N_9604);
nand UO_704 (O_704,N_9154,N_9574);
or UO_705 (O_705,N_9687,N_9900);
nor UO_706 (O_706,N_9060,N_9001);
nand UO_707 (O_707,N_9886,N_9640);
nand UO_708 (O_708,N_9309,N_9413);
nor UO_709 (O_709,N_9832,N_9597);
nand UO_710 (O_710,N_9523,N_9931);
or UO_711 (O_711,N_9831,N_9023);
or UO_712 (O_712,N_9741,N_9146);
nand UO_713 (O_713,N_9137,N_9613);
and UO_714 (O_714,N_9049,N_9670);
nand UO_715 (O_715,N_9885,N_9124);
nand UO_716 (O_716,N_9585,N_9311);
nor UO_717 (O_717,N_9161,N_9095);
and UO_718 (O_718,N_9599,N_9778);
nor UO_719 (O_719,N_9621,N_9727);
nand UO_720 (O_720,N_9365,N_9767);
or UO_721 (O_721,N_9231,N_9438);
and UO_722 (O_722,N_9894,N_9325);
or UO_723 (O_723,N_9960,N_9291);
or UO_724 (O_724,N_9288,N_9093);
nand UO_725 (O_725,N_9160,N_9107);
and UO_726 (O_726,N_9048,N_9787);
and UO_727 (O_727,N_9732,N_9525);
nand UO_728 (O_728,N_9601,N_9720);
or UO_729 (O_729,N_9360,N_9094);
and UO_730 (O_730,N_9340,N_9549);
nor UO_731 (O_731,N_9940,N_9098);
nand UO_732 (O_732,N_9784,N_9433);
nor UO_733 (O_733,N_9415,N_9238);
xor UO_734 (O_734,N_9947,N_9952);
or UO_735 (O_735,N_9279,N_9266);
and UO_736 (O_736,N_9370,N_9198);
and UO_737 (O_737,N_9439,N_9773);
nand UO_738 (O_738,N_9233,N_9447);
or UO_739 (O_739,N_9666,N_9315);
or UO_740 (O_740,N_9960,N_9227);
and UO_741 (O_741,N_9062,N_9364);
and UO_742 (O_742,N_9507,N_9396);
and UO_743 (O_743,N_9390,N_9207);
nor UO_744 (O_744,N_9381,N_9922);
or UO_745 (O_745,N_9615,N_9408);
or UO_746 (O_746,N_9717,N_9074);
nor UO_747 (O_747,N_9566,N_9480);
or UO_748 (O_748,N_9273,N_9633);
or UO_749 (O_749,N_9392,N_9208);
xnor UO_750 (O_750,N_9010,N_9596);
or UO_751 (O_751,N_9575,N_9956);
nand UO_752 (O_752,N_9808,N_9705);
or UO_753 (O_753,N_9391,N_9499);
or UO_754 (O_754,N_9986,N_9950);
or UO_755 (O_755,N_9859,N_9860);
or UO_756 (O_756,N_9344,N_9886);
or UO_757 (O_757,N_9040,N_9499);
nor UO_758 (O_758,N_9006,N_9231);
nand UO_759 (O_759,N_9333,N_9112);
nor UO_760 (O_760,N_9612,N_9233);
xnor UO_761 (O_761,N_9401,N_9056);
nand UO_762 (O_762,N_9019,N_9035);
xor UO_763 (O_763,N_9087,N_9572);
and UO_764 (O_764,N_9007,N_9202);
nand UO_765 (O_765,N_9403,N_9932);
and UO_766 (O_766,N_9356,N_9899);
and UO_767 (O_767,N_9179,N_9459);
and UO_768 (O_768,N_9091,N_9415);
or UO_769 (O_769,N_9543,N_9898);
nand UO_770 (O_770,N_9363,N_9754);
nand UO_771 (O_771,N_9059,N_9747);
or UO_772 (O_772,N_9180,N_9877);
nand UO_773 (O_773,N_9211,N_9672);
and UO_774 (O_774,N_9739,N_9137);
and UO_775 (O_775,N_9353,N_9314);
or UO_776 (O_776,N_9923,N_9329);
nand UO_777 (O_777,N_9555,N_9824);
and UO_778 (O_778,N_9279,N_9616);
xor UO_779 (O_779,N_9914,N_9637);
nor UO_780 (O_780,N_9169,N_9217);
nor UO_781 (O_781,N_9084,N_9027);
nor UO_782 (O_782,N_9098,N_9606);
or UO_783 (O_783,N_9085,N_9990);
or UO_784 (O_784,N_9995,N_9852);
or UO_785 (O_785,N_9784,N_9672);
and UO_786 (O_786,N_9184,N_9534);
nor UO_787 (O_787,N_9405,N_9647);
nand UO_788 (O_788,N_9297,N_9372);
nor UO_789 (O_789,N_9994,N_9301);
or UO_790 (O_790,N_9137,N_9650);
and UO_791 (O_791,N_9902,N_9035);
and UO_792 (O_792,N_9393,N_9923);
or UO_793 (O_793,N_9524,N_9609);
and UO_794 (O_794,N_9634,N_9033);
or UO_795 (O_795,N_9755,N_9761);
and UO_796 (O_796,N_9695,N_9917);
or UO_797 (O_797,N_9983,N_9489);
nor UO_798 (O_798,N_9783,N_9606);
nand UO_799 (O_799,N_9868,N_9438);
and UO_800 (O_800,N_9589,N_9246);
nand UO_801 (O_801,N_9529,N_9395);
nand UO_802 (O_802,N_9965,N_9106);
nor UO_803 (O_803,N_9761,N_9117);
xnor UO_804 (O_804,N_9720,N_9699);
nand UO_805 (O_805,N_9915,N_9270);
xor UO_806 (O_806,N_9756,N_9867);
or UO_807 (O_807,N_9511,N_9919);
or UO_808 (O_808,N_9284,N_9504);
nand UO_809 (O_809,N_9609,N_9812);
or UO_810 (O_810,N_9900,N_9850);
or UO_811 (O_811,N_9875,N_9488);
nor UO_812 (O_812,N_9338,N_9886);
nor UO_813 (O_813,N_9946,N_9963);
nor UO_814 (O_814,N_9316,N_9344);
nand UO_815 (O_815,N_9029,N_9047);
or UO_816 (O_816,N_9756,N_9618);
nor UO_817 (O_817,N_9854,N_9746);
and UO_818 (O_818,N_9589,N_9438);
and UO_819 (O_819,N_9233,N_9726);
and UO_820 (O_820,N_9531,N_9404);
or UO_821 (O_821,N_9762,N_9283);
nand UO_822 (O_822,N_9556,N_9409);
or UO_823 (O_823,N_9959,N_9207);
nor UO_824 (O_824,N_9048,N_9019);
or UO_825 (O_825,N_9040,N_9889);
or UO_826 (O_826,N_9872,N_9212);
and UO_827 (O_827,N_9629,N_9276);
nand UO_828 (O_828,N_9020,N_9317);
or UO_829 (O_829,N_9882,N_9923);
or UO_830 (O_830,N_9548,N_9613);
and UO_831 (O_831,N_9418,N_9188);
or UO_832 (O_832,N_9077,N_9741);
nor UO_833 (O_833,N_9750,N_9160);
or UO_834 (O_834,N_9772,N_9712);
nor UO_835 (O_835,N_9531,N_9386);
nand UO_836 (O_836,N_9615,N_9224);
or UO_837 (O_837,N_9175,N_9525);
nand UO_838 (O_838,N_9065,N_9940);
nor UO_839 (O_839,N_9377,N_9869);
nand UO_840 (O_840,N_9955,N_9342);
or UO_841 (O_841,N_9411,N_9224);
or UO_842 (O_842,N_9363,N_9687);
or UO_843 (O_843,N_9472,N_9036);
nor UO_844 (O_844,N_9970,N_9744);
or UO_845 (O_845,N_9651,N_9578);
nor UO_846 (O_846,N_9741,N_9577);
and UO_847 (O_847,N_9115,N_9450);
and UO_848 (O_848,N_9243,N_9131);
nand UO_849 (O_849,N_9247,N_9892);
nand UO_850 (O_850,N_9387,N_9072);
nand UO_851 (O_851,N_9672,N_9964);
nand UO_852 (O_852,N_9054,N_9732);
nor UO_853 (O_853,N_9619,N_9969);
nand UO_854 (O_854,N_9723,N_9443);
and UO_855 (O_855,N_9556,N_9000);
nand UO_856 (O_856,N_9752,N_9717);
nor UO_857 (O_857,N_9798,N_9389);
nor UO_858 (O_858,N_9275,N_9308);
or UO_859 (O_859,N_9914,N_9268);
and UO_860 (O_860,N_9477,N_9570);
or UO_861 (O_861,N_9566,N_9653);
or UO_862 (O_862,N_9201,N_9156);
nand UO_863 (O_863,N_9390,N_9271);
nor UO_864 (O_864,N_9157,N_9323);
or UO_865 (O_865,N_9562,N_9338);
nand UO_866 (O_866,N_9069,N_9146);
nor UO_867 (O_867,N_9272,N_9795);
nor UO_868 (O_868,N_9200,N_9794);
nand UO_869 (O_869,N_9148,N_9989);
nor UO_870 (O_870,N_9631,N_9663);
and UO_871 (O_871,N_9796,N_9839);
and UO_872 (O_872,N_9073,N_9339);
nor UO_873 (O_873,N_9660,N_9746);
nand UO_874 (O_874,N_9602,N_9273);
nor UO_875 (O_875,N_9438,N_9020);
or UO_876 (O_876,N_9199,N_9026);
or UO_877 (O_877,N_9193,N_9967);
nor UO_878 (O_878,N_9608,N_9350);
nand UO_879 (O_879,N_9119,N_9095);
or UO_880 (O_880,N_9781,N_9532);
and UO_881 (O_881,N_9601,N_9868);
nand UO_882 (O_882,N_9349,N_9285);
nor UO_883 (O_883,N_9897,N_9881);
and UO_884 (O_884,N_9760,N_9422);
and UO_885 (O_885,N_9381,N_9608);
nand UO_886 (O_886,N_9213,N_9696);
or UO_887 (O_887,N_9825,N_9678);
nand UO_888 (O_888,N_9472,N_9147);
nand UO_889 (O_889,N_9361,N_9549);
and UO_890 (O_890,N_9155,N_9594);
and UO_891 (O_891,N_9540,N_9223);
nand UO_892 (O_892,N_9716,N_9593);
nand UO_893 (O_893,N_9196,N_9106);
xnor UO_894 (O_894,N_9827,N_9539);
nor UO_895 (O_895,N_9767,N_9226);
or UO_896 (O_896,N_9417,N_9985);
or UO_897 (O_897,N_9790,N_9810);
nand UO_898 (O_898,N_9240,N_9451);
nand UO_899 (O_899,N_9439,N_9548);
nor UO_900 (O_900,N_9204,N_9484);
nand UO_901 (O_901,N_9809,N_9275);
xor UO_902 (O_902,N_9219,N_9734);
and UO_903 (O_903,N_9947,N_9668);
nor UO_904 (O_904,N_9199,N_9537);
and UO_905 (O_905,N_9459,N_9846);
or UO_906 (O_906,N_9232,N_9623);
and UO_907 (O_907,N_9631,N_9304);
and UO_908 (O_908,N_9594,N_9543);
nand UO_909 (O_909,N_9459,N_9659);
or UO_910 (O_910,N_9580,N_9353);
and UO_911 (O_911,N_9230,N_9312);
nor UO_912 (O_912,N_9415,N_9518);
and UO_913 (O_913,N_9901,N_9165);
or UO_914 (O_914,N_9694,N_9967);
nor UO_915 (O_915,N_9300,N_9257);
or UO_916 (O_916,N_9662,N_9240);
or UO_917 (O_917,N_9384,N_9502);
or UO_918 (O_918,N_9554,N_9848);
and UO_919 (O_919,N_9153,N_9429);
nor UO_920 (O_920,N_9146,N_9842);
nor UO_921 (O_921,N_9511,N_9682);
or UO_922 (O_922,N_9501,N_9563);
and UO_923 (O_923,N_9526,N_9029);
or UO_924 (O_924,N_9828,N_9192);
or UO_925 (O_925,N_9301,N_9762);
or UO_926 (O_926,N_9687,N_9909);
nor UO_927 (O_927,N_9209,N_9825);
nand UO_928 (O_928,N_9431,N_9510);
nor UO_929 (O_929,N_9951,N_9674);
nor UO_930 (O_930,N_9836,N_9867);
and UO_931 (O_931,N_9712,N_9509);
and UO_932 (O_932,N_9502,N_9511);
and UO_933 (O_933,N_9416,N_9471);
nand UO_934 (O_934,N_9005,N_9203);
nand UO_935 (O_935,N_9709,N_9975);
nand UO_936 (O_936,N_9341,N_9483);
or UO_937 (O_937,N_9450,N_9405);
nor UO_938 (O_938,N_9584,N_9171);
xor UO_939 (O_939,N_9871,N_9406);
or UO_940 (O_940,N_9814,N_9953);
and UO_941 (O_941,N_9535,N_9015);
or UO_942 (O_942,N_9592,N_9499);
nor UO_943 (O_943,N_9460,N_9562);
or UO_944 (O_944,N_9584,N_9429);
and UO_945 (O_945,N_9848,N_9990);
nor UO_946 (O_946,N_9103,N_9965);
or UO_947 (O_947,N_9275,N_9022);
and UO_948 (O_948,N_9752,N_9155);
and UO_949 (O_949,N_9258,N_9207);
nand UO_950 (O_950,N_9560,N_9688);
and UO_951 (O_951,N_9419,N_9069);
nand UO_952 (O_952,N_9984,N_9335);
nor UO_953 (O_953,N_9296,N_9630);
nor UO_954 (O_954,N_9911,N_9925);
nand UO_955 (O_955,N_9580,N_9257);
nor UO_956 (O_956,N_9118,N_9737);
or UO_957 (O_957,N_9511,N_9982);
or UO_958 (O_958,N_9555,N_9036);
and UO_959 (O_959,N_9499,N_9832);
nand UO_960 (O_960,N_9441,N_9375);
and UO_961 (O_961,N_9738,N_9660);
or UO_962 (O_962,N_9227,N_9159);
nor UO_963 (O_963,N_9193,N_9794);
xnor UO_964 (O_964,N_9652,N_9549);
nor UO_965 (O_965,N_9831,N_9355);
or UO_966 (O_966,N_9082,N_9531);
and UO_967 (O_967,N_9159,N_9924);
nand UO_968 (O_968,N_9801,N_9097);
and UO_969 (O_969,N_9233,N_9362);
nor UO_970 (O_970,N_9313,N_9426);
or UO_971 (O_971,N_9690,N_9996);
or UO_972 (O_972,N_9670,N_9504);
nand UO_973 (O_973,N_9409,N_9113);
and UO_974 (O_974,N_9017,N_9924);
nand UO_975 (O_975,N_9756,N_9295);
and UO_976 (O_976,N_9741,N_9366);
nand UO_977 (O_977,N_9297,N_9627);
or UO_978 (O_978,N_9147,N_9250);
or UO_979 (O_979,N_9885,N_9643);
nand UO_980 (O_980,N_9390,N_9480);
nand UO_981 (O_981,N_9372,N_9724);
nor UO_982 (O_982,N_9065,N_9010);
nand UO_983 (O_983,N_9940,N_9865);
nand UO_984 (O_984,N_9084,N_9022);
nand UO_985 (O_985,N_9109,N_9914);
or UO_986 (O_986,N_9938,N_9487);
and UO_987 (O_987,N_9286,N_9293);
or UO_988 (O_988,N_9546,N_9265);
nor UO_989 (O_989,N_9642,N_9177);
nor UO_990 (O_990,N_9136,N_9242);
or UO_991 (O_991,N_9966,N_9821);
nor UO_992 (O_992,N_9477,N_9109);
nand UO_993 (O_993,N_9409,N_9171);
and UO_994 (O_994,N_9465,N_9640);
nor UO_995 (O_995,N_9436,N_9080);
and UO_996 (O_996,N_9775,N_9217);
or UO_997 (O_997,N_9994,N_9616);
nor UO_998 (O_998,N_9398,N_9437);
nand UO_999 (O_999,N_9706,N_9193);
nor UO_1000 (O_1000,N_9475,N_9801);
or UO_1001 (O_1001,N_9134,N_9984);
nand UO_1002 (O_1002,N_9194,N_9073);
or UO_1003 (O_1003,N_9857,N_9555);
and UO_1004 (O_1004,N_9371,N_9209);
and UO_1005 (O_1005,N_9988,N_9515);
and UO_1006 (O_1006,N_9645,N_9372);
or UO_1007 (O_1007,N_9178,N_9961);
nand UO_1008 (O_1008,N_9842,N_9094);
or UO_1009 (O_1009,N_9610,N_9403);
or UO_1010 (O_1010,N_9465,N_9875);
or UO_1011 (O_1011,N_9730,N_9872);
nor UO_1012 (O_1012,N_9371,N_9549);
nand UO_1013 (O_1013,N_9476,N_9417);
nor UO_1014 (O_1014,N_9249,N_9112);
nand UO_1015 (O_1015,N_9834,N_9213);
nor UO_1016 (O_1016,N_9597,N_9360);
and UO_1017 (O_1017,N_9403,N_9243);
or UO_1018 (O_1018,N_9924,N_9829);
or UO_1019 (O_1019,N_9337,N_9236);
and UO_1020 (O_1020,N_9557,N_9013);
nor UO_1021 (O_1021,N_9353,N_9049);
nand UO_1022 (O_1022,N_9308,N_9891);
nand UO_1023 (O_1023,N_9829,N_9395);
nor UO_1024 (O_1024,N_9334,N_9942);
nand UO_1025 (O_1025,N_9602,N_9471);
and UO_1026 (O_1026,N_9753,N_9108);
nor UO_1027 (O_1027,N_9988,N_9877);
nand UO_1028 (O_1028,N_9423,N_9889);
nor UO_1029 (O_1029,N_9475,N_9366);
or UO_1030 (O_1030,N_9945,N_9653);
nand UO_1031 (O_1031,N_9267,N_9215);
nand UO_1032 (O_1032,N_9516,N_9125);
nor UO_1033 (O_1033,N_9757,N_9745);
or UO_1034 (O_1034,N_9355,N_9209);
nand UO_1035 (O_1035,N_9386,N_9300);
and UO_1036 (O_1036,N_9344,N_9609);
and UO_1037 (O_1037,N_9723,N_9216);
nand UO_1038 (O_1038,N_9190,N_9642);
nor UO_1039 (O_1039,N_9544,N_9699);
nand UO_1040 (O_1040,N_9350,N_9783);
nor UO_1041 (O_1041,N_9017,N_9563);
or UO_1042 (O_1042,N_9308,N_9799);
nand UO_1043 (O_1043,N_9142,N_9899);
or UO_1044 (O_1044,N_9063,N_9508);
nand UO_1045 (O_1045,N_9592,N_9843);
nor UO_1046 (O_1046,N_9027,N_9336);
or UO_1047 (O_1047,N_9700,N_9955);
and UO_1048 (O_1048,N_9977,N_9697);
nand UO_1049 (O_1049,N_9676,N_9140);
nor UO_1050 (O_1050,N_9276,N_9287);
nor UO_1051 (O_1051,N_9491,N_9548);
or UO_1052 (O_1052,N_9176,N_9106);
or UO_1053 (O_1053,N_9996,N_9524);
and UO_1054 (O_1054,N_9512,N_9667);
nand UO_1055 (O_1055,N_9394,N_9173);
nor UO_1056 (O_1056,N_9804,N_9938);
and UO_1057 (O_1057,N_9980,N_9331);
nand UO_1058 (O_1058,N_9688,N_9015);
or UO_1059 (O_1059,N_9713,N_9384);
or UO_1060 (O_1060,N_9162,N_9977);
xor UO_1061 (O_1061,N_9307,N_9244);
or UO_1062 (O_1062,N_9746,N_9032);
nand UO_1063 (O_1063,N_9748,N_9979);
nor UO_1064 (O_1064,N_9187,N_9089);
xor UO_1065 (O_1065,N_9464,N_9731);
or UO_1066 (O_1066,N_9558,N_9596);
nand UO_1067 (O_1067,N_9320,N_9818);
and UO_1068 (O_1068,N_9053,N_9848);
or UO_1069 (O_1069,N_9270,N_9143);
nand UO_1070 (O_1070,N_9714,N_9299);
nand UO_1071 (O_1071,N_9285,N_9840);
nor UO_1072 (O_1072,N_9258,N_9627);
and UO_1073 (O_1073,N_9754,N_9552);
nand UO_1074 (O_1074,N_9655,N_9092);
and UO_1075 (O_1075,N_9199,N_9759);
nor UO_1076 (O_1076,N_9805,N_9823);
nor UO_1077 (O_1077,N_9778,N_9203);
and UO_1078 (O_1078,N_9778,N_9183);
and UO_1079 (O_1079,N_9690,N_9918);
nand UO_1080 (O_1080,N_9817,N_9397);
and UO_1081 (O_1081,N_9574,N_9933);
nor UO_1082 (O_1082,N_9359,N_9955);
nand UO_1083 (O_1083,N_9233,N_9740);
and UO_1084 (O_1084,N_9642,N_9387);
nand UO_1085 (O_1085,N_9650,N_9028);
and UO_1086 (O_1086,N_9454,N_9187);
nor UO_1087 (O_1087,N_9718,N_9667);
and UO_1088 (O_1088,N_9361,N_9019);
or UO_1089 (O_1089,N_9569,N_9944);
or UO_1090 (O_1090,N_9943,N_9478);
nand UO_1091 (O_1091,N_9922,N_9102);
nor UO_1092 (O_1092,N_9584,N_9742);
or UO_1093 (O_1093,N_9074,N_9124);
nand UO_1094 (O_1094,N_9996,N_9372);
and UO_1095 (O_1095,N_9105,N_9135);
or UO_1096 (O_1096,N_9682,N_9915);
or UO_1097 (O_1097,N_9064,N_9081);
nor UO_1098 (O_1098,N_9819,N_9357);
or UO_1099 (O_1099,N_9916,N_9402);
nor UO_1100 (O_1100,N_9635,N_9561);
and UO_1101 (O_1101,N_9386,N_9274);
nor UO_1102 (O_1102,N_9507,N_9998);
or UO_1103 (O_1103,N_9147,N_9675);
nor UO_1104 (O_1104,N_9878,N_9829);
nor UO_1105 (O_1105,N_9966,N_9088);
or UO_1106 (O_1106,N_9692,N_9576);
or UO_1107 (O_1107,N_9553,N_9602);
nand UO_1108 (O_1108,N_9280,N_9169);
and UO_1109 (O_1109,N_9974,N_9545);
or UO_1110 (O_1110,N_9618,N_9912);
and UO_1111 (O_1111,N_9673,N_9846);
nor UO_1112 (O_1112,N_9800,N_9305);
nor UO_1113 (O_1113,N_9901,N_9622);
and UO_1114 (O_1114,N_9439,N_9554);
and UO_1115 (O_1115,N_9450,N_9230);
and UO_1116 (O_1116,N_9445,N_9592);
and UO_1117 (O_1117,N_9932,N_9749);
and UO_1118 (O_1118,N_9915,N_9817);
or UO_1119 (O_1119,N_9521,N_9675);
nand UO_1120 (O_1120,N_9486,N_9968);
or UO_1121 (O_1121,N_9601,N_9240);
or UO_1122 (O_1122,N_9317,N_9989);
nand UO_1123 (O_1123,N_9145,N_9914);
nand UO_1124 (O_1124,N_9024,N_9606);
nor UO_1125 (O_1125,N_9273,N_9578);
or UO_1126 (O_1126,N_9883,N_9784);
and UO_1127 (O_1127,N_9769,N_9103);
and UO_1128 (O_1128,N_9493,N_9917);
nor UO_1129 (O_1129,N_9356,N_9274);
nand UO_1130 (O_1130,N_9663,N_9266);
nor UO_1131 (O_1131,N_9507,N_9196);
and UO_1132 (O_1132,N_9497,N_9694);
nand UO_1133 (O_1133,N_9881,N_9144);
nor UO_1134 (O_1134,N_9386,N_9236);
nor UO_1135 (O_1135,N_9434,N_9372);
nor UO_1136 (O_1136,N_9486,N_9147);
nand UO_1137 (O_1137,N_9436,N_9423);
or UO_1138 (O_1138,N_9716,N_9792);
nor UO_1139 (O_1139,N_9196,N_9740);
and UO_1140 (O_1140,N_9866,N_9078);
and UO_1141 (O_1141,N_9349,N_9977);
nand UO_1142 (O_1142,N_9582,N_9174);
or UO_1143 (O_1143,N_9190,N_9384);
nor UO_1144 (O_1144,N_9628,N_9044);
nand UO_1145 (O_1145,N_9600,N_9781);
xor UO_1146 (O_1146,N_9260,N_9429);
or UO_1147 (O_1147,N_9969,N_9803);
or UO_1148 (O_1148,N_9826,N_9967);
nor UO_1149 (O_1149,N_9859,N_9931);
or UO_1150 (O_1150,N_9628,N_9875);
nand UO_1151 (O_1151,N_9875,N_9246);
nor UO_1152 (O_1152,N_9489,N_9377);
and UO_1153 (O_1153,N_9226,N_9871);
or UO_1154 (O_1154,N_9455,N_9982);
nor UO_1155 (O_1155,N_9188,N_9721);
or UO_1156 (O_1156,N_9509,N_9755);
or UO_1157 (O_1157,N_9773,N_9981);
or UO_1158 (O_1158,N_9604,N_9549);
nor UO_1159 (O_1159,N_9924,N_9428);
or UO_1160 (O_1160,N_9586,N_9122);
xnor UO_1161 (O_1161,N_9769,N_9649);
nor UO_1162 (O_1162,N_9448,N_9126);
nand UO_1163 (O_1163,N_9796,N_9916);
nand UO_1164 (O_1164,N_9542,N_9939);
or UO_1165 (O_1165,N_9534,N_9827);
nor UO_1166 (O_1166,N_9625,N_9588);
and UO_1167 (O_1167,N_9326,N_9930);
nor UO_1168 (O_1168,N_9818,N_9539);
or UO_1169 (O_1169,N_9805,N_9750);
or UO_1170 (O_1170,N_9529,N_9886);
nor UO_1171 (O_1171,N_9849,N_9160);
nand UO_1172 (O_1172,N_9587,N_9939);
nand UO_1173 (O_1173,N_9792,N_9331);
or UO_1174 (O_1174,N_9647,N_9865);
nand UO_1175 (O_1175,N_9205,N_9864);
or UO_1176 (O_1176,N_9053,N_9018);
and UO_1177 (O_1177,N_9733,N_9004);
or UO_1178 (O_1178,N_9588,N_9453);
nand UO_1179 (O_1179,N_9204,N_9093);
nand UO_1180 (O_1180,N_9910,N_9969);
nor UO_1181 (O_1181,N_9549,N_9514);
and UO_1182 (O_1182,N_9337,N_9176);
nand UO_1183 (O_1183,N_9563,N_9150);
xnor UO_1184 (O_1184,N_9805,N_9229);
and UO_1185 (O_1185,N_9524,N_9183);
or UO_1186 (O_1186,N_9086,N_9174);
or UO_1187 (O_1187,N_9010,N_9746);
and UO_1188 (O_1188,N_9685,N_9868);
or UO_1189 (O_1189,N_9406,N_9212);
nor UO_1190 (O_1190,N_9012,N_9025);
or UO_1191 (O_1191,N_9501,N_9633);
and UO_1192 (O_1192,N_9128,N_9361);
or UO_1193 (O_1193,N_9041,N_9623);
nor UO_1194 (O_1194,N_9318,N_9914);
nor UO_1195 (O_1195,N_9868,N_9368);
nand UO_1196 (O_1196,N_9210,N_9757);
nand UO_1197 (O_1197,N_9471,N_9157);
nand UO_1198 (O_1198,N_9863,N_9285);
nand UO_1199 (O_1199,N_9318,N_9817);
nor UO_1200 (O_1200,N_9834,N_9152);
nor UO_1201 (O_1201,N_9847,N_9335);
nand UO_1202 (O_1202,N_9222,N_9241);
or UO_1203 (O_1203,N_9410,N_9201);
nor UO_1204 (O_1204,N_9710,N_9517);
nor UO_1205 (O_1205,N_9084,N_9409);
or UO_1206 (O_1206,N_9407,N_9460);
nor UO_1207 (O_1207,N_9238,N_9659);
and UO_1208 (O_1208,N_9776,N_9387);
or UO_1209 (O_1209,N_9723,N_9622);
nor UO_1210 (O_1210,N_9649,N_9413);
or UO_1211 (O_1211,N_9301,N_9540);
or UO_1212 (O_1212,N_9486,N_9630);
nor UO_1213 (O_1213,N_9433,N_9700);
or UO_1214 (O_1214,N_9196,N_9739);
nor UO_1215 (O_1215,N_9160,N_9755);
or UO_1216 (O_1216,N_9851,N_9095);
nor UO_1217 (O_1217,N_9656,N_9229);
nand UO_1218 (O_1218,N_9935,N_9362);
and UO_1219 (O_1219,N_9685,N_9336);
nor UO_1220 (O_1220,N_9092,N_9813);
and UO_1221 (O_1221,N_9445,N_9596);
and UO_1222 (O_1222,N_9754,N_9291);
and UO_1223 (O_1223,N_9154,N_9534);
or UO_1224 (O_1224,N_9361,N_9313);
nand UO_1225 (O_1225,N_9458,N_9572);
and UO_1226 (O_1226,N_9801,N_9716);
nor UO_1227 (O_1227,N_9308,N_9995);
nand UO_1228 (O_1228,N_9426,N_9348);
and UO_1229 (O_1229,N_9019,N_9066);
nand UO_1230 (O_1230,N_9131,N_9176);
and UO_1231 (O_1231,N_9522,N_9509);
and UO_1232 (O_1232,N_9815,N_9422);
nand UO_1233 (O_1233,N_9602,N_9939);
xnor UO_1234 (O_1234,N_9133,N_9948);
nor UO_1235 (O_1235,N_9004,N_9391);
nand UO_1236 (O_1236,N_9609,N_9293);
and UO_1237 (O_1237,N_9609,N_9186);
or UO_1238 (O_1238,N_9337,N_9276);
nor UO_1239 (O_1239,N_9071,N_9064);
or UO_1240 (O_1240,N_9205,N_9503);
nand UO_1241 (O_1241,N_9707,N_9781);
and UO_1242 (O_1242,N_9636,N_9811);
nand UO_1243 (O_1243,N_9991,N_9152);
nand UO_1244 (O_1244,N_9013,N_9175);
and UO_1245 (O_1245,N_9548,N_9592);
nor UO_1246 (O_1246,N_9131,N_9183);
nor UO_1247 (O_1247,N_9670,N_9004);
xor UO_1248 (O_1248,N_9629,N_9762);
nor UO_1249 (O_1249,N_9285,N_9286);
nand UO_1250 (O_1250,N_9272,N_9587);
nor UO_1251 (O_1251,N_9245,N_9931);
nor UO_1252 (O_1252,N_9709,N_9977);
nand UO_1253 (O_1253,N_9233,N_9570);
nand UO_1254 (O_1254,N_9460,N_9763);
nand UO_1255 (O_1255,N_9201,N_9283);
nand UO_1256 (O_1256,N_9646,N_9642);
and UO_1257 (O_1257,N_9731,N_9846);
nand UO_1258 (O_1258,N_9986,N_9035);
nor UO_1259 (O_1259,N_9089,N_9633);
nor UO_1260 (O_1260,N_9418,N_9266);
nand UO_1261 (O_1261,N_9928,N_9456);
and UO_1262 (O_1262,N_9125,N_9118);
nand UO_1263 (O_1263,N_9032,N_9874);
and UO_1264 (O_1264,N_9593,N_9888);
nand UO_1265 (O_1265,N_9067,N_9037);
xnor UO_1266 (O_1266,N_9308,N_9784);
or UO_1267 (O_1267,N_9100,N_9263);
or UO_1268 (O_1268,N_9087,N_9307);
nand UO_1269 (O_1269,N_9553,N_9102);
or UO_1270 (O_1270,N_9626,N_9243);
or UO_1271 (O_1271,N_9474,N_9557);
and UO_1272 (O_1272,N_9484,N_9548);
or UO_1273 (O_1273,N_9564,N_9902);
and UO_1274 (O_1274,N_9940,N_9633);
and UO_1275 (O_1275,N_9845,N_9791);
and UO_1276 (O_1276,N_9244,N_9976);
and UO_1277 (O_1277,N_9337,N_9537);
and UO_1278 (O_1278,N_9228,N_9917);
nand UO_1279 (O_1279,N_9140,N_9547);
or UO_1280 (O_1280,N_9616,N_9342);
nor UO_1281 (O_1281,N_9579,N_9024);
nor UO_1282 (O_1282,N_9788,N_9345);
nand UO_1283 (O_1283,N_9056,N_9462);
or UO_1284 (O_1284,N_9809,N_9660);
or UO_1285 (O_1285,N_9688,N_9696);
nor UO_1286 (O_1286,N_9776,N_9335);
and UO_1287 (O_1287,N_9626,N_9817);
nand UO_1288 (O_1288,N_9667,N_9928);
nand UO_1289 (O_1289,N_9743,N_9999);
nand UO_1290 (O_1290,N_9401,N_9701);
and UO_1291 (O_1291,N_9889,N_9578);
nor UO_1292 (O_1292,N_9952,N_9285);
nand UO_1293 (O_1293,N_9476,N_9547);
nor UO_1294 (O_1294,N_9652,N_9712);
xnor UO_1295 (O_1295,N_9199,N_9163);
and UO_1296 (O_1296,N_9445,N_9429);
nor UO_1297 (O_1297,N_9959,N_9191);
nor UO_1298 (O_1298,N_9745,N_9151);
nand UO_1299 (O_1299,N_9934,N_9766);
nand UO_1300 (O_1300,N_9192,N_9540);
and UO_1301 (O_1301,N_9131,N_9490);
nor UO_1302 (O_1302,N_9543,N_9829);
or UO_1303 (O_1303,N_9261,N_9402);
and UO_1304 (O_1304,N_9569,N_9987);
and UO_1305 (O_1305,N_9396,N_9418);
nand UO_1306 (O_1306,N_9837,N_9368);
nor UO_1307 (O_1307,N_9974,N_9048);
and UO_1308 (O_1308,N_9331,N_9408);
nor UO_1309 (O_1309,N_9982,N_9621);
nor UO_1310 (O_1310,N_9666,N_9917);
or UO_1311 (O_1311,N_9522,N_9221);
nor UO_1312 (O_1312,N_9320,N_9442);
and UO_1313 (O_1313,N_9247,N_9884);
nor UO_1314 (O_1314,N_9558,N_9326);
and UO_1315 (O_1315,N_9314,N_9155);
nor UO_1316 (O_1316,N_9643,N_9932);
or UO_1317 (O_1317,N_9823,N_9870);
nor UO_1318 (O_1318,N_9759,N_9995);
nand UO_1319 (O_1319,N_9017,N_9167);
and UO_1320 (O_1320,N_9300,N_9618);
nor UO_1321 (O_1321,N_9577,N_9374);
or UO_1322 (O_1322,N_9116,N_9522);
or UO_1323 (O_1323,N_9700,N_9649);
or UO_1324 (O_1324,N_9361,N_9939);
and UO_1325 (O_1325,N_9784,N_9192);
or UO_1326 (O_1326,N_9139,N_9226);
nor UO_1327 (O_1327,N_9946,N_9941);
nand UO_1328 (O_1328,N_9748,N_9355);
nand UO_1329 (O_1329,N_9634,N_9477);
nand UO_1330 (O_1330,N_9522,N_9930);
and UO_1331 (O_1331,N_9776,N_9936);
nor UO_1332 (O_1332,N_9019,N_9421);
and UO_1333 (O_1333,N_9894,N_9189);
nand UO_1334 (O_1334,N_9536,N_9990);
nor UO_1335 (O_1335,N_9337,N_9271);
nor UO_1336 (O_1336,N_9889,N_9223);
nand UO_1337 (O_1337,N_9535,N_9456);
and UO_1338 (O_1338,N_9306,N_9678);
nand UO_1339 (O_1339,N_9096,N_9762);
or UO_1340 (O_1340,N_9829,N_9446);
nand UO_1341 (O_1341,N_9064,N_9478);
nand UO_1342 (O_1342,N_9265,N_9917);
nor UO_1343 (O_1343,N_9254,N_9740);
and UO_1344 (O_1344,N_9646,N_9918);
nor UO_1345 (O_1345,N_9095,N_9300);
or UO_1346 (O_1346,N_9706,N_9041);
nor UO_1347 (O_1347,N_9797,N_9804);
nor UO_1348 (O_1348,N_9957,N_9854);
and UO_1349 (O_1349,N_9167,N_9732);
nor UO_1350 (O_1350,N_9407,N_9258);
nand UO_1351 (O_1351,N_9593,N_9766);
or UO_1352 (O_1352,N_9572,N_9096);
or UO_1353 (O_1353,N_9354,N_9735);
and UO_1354 (O_1354,N_9985,N_9030);
or UO_1355 (O_1355,N_9379,N_9153);
and UO_1356 (O_1356,N_9976,N_9132);
nand UO_1357 (O_1357,N_9770,N_9649);
nor UO_1358 (O_1358,N_9592,N_9988);
and UO_1359 (O_1359,N_9710,N_9944);
nand UO_1360 (O_1360,N_9415,N_9709);
nor UO_1361 (O_1361,N_9605,N_9118);
or UO_1362 (O_1362,N_9455,N_9444);
nand UO_1363 (O_1363,N_9090,N_9695);
or UO_1364 (O_1364,N_9347,N_9099);
or UO_1365 (O_1365,N_9178,N_9018);
nand UO_1366 (O_1366,N_9095,N_9078);
nor UO_1367 (O_1367,N_9438,N_9799);
and UO_1368 (O_1368,N_9736,N_9866);
and UO_1369 (O_1369,N_9813,N_9216);
nor UO_1370 (O_1370,N_9743,N_9608);
nand UO_1371 (O_1371,N_9626,N_9135);
nor UO_1372 (O_1372,N_9006,N_9662);
nand UO_1373 (O_1373,N_9302,N_9666);
or UO_1374 (O_1374,N_9638,N_9226);
nand UO_1375 (O_1375,N_9534,N_9072);
nand UO_1376 (O_1376,N_9952,N_9922);
and UO_1377 (O_1377,N_9221,N_9922);
or UO_1378 (O_1378,N_9805,N_9418);
and UO_1379 (O_1379,N_9821,N_9667);
nand UO_1380 (O_1380,N_9015,N_9052);
nor UO_1381 (O_1381,N_9549,N_9396);
and UO_1382 (O_1382,N_9946,N_9905);
nor UO_1383 (O_1383,N_9216,N_9129);
or UO_1384 (O_1384,N_9941,N_9481);
nor UO_1385 (O_1385,N_9466,N_9891);
or UO_1386 (O_1386,N_9034,N_9116);
or UO_1387 (O_1387,N_9282,N_9537);
nor UO_1388 (O_1388,N_9298,N_9308);
nand UO_1389 (O_1389,N_9486,N_9108);
or UO_1390 (O_1390,N_9534,N_9140);
or UO_1391 (O_1391,N_9521,N_9950);
and UO_1392 (O_1392,N_9121,N_9705);
or UO_1393 (O_1393,N_9191,N_9207);
nor UO_1394 (O_1394,N_9245,N_9545);
or UO_1395 (O_1395,N_9549,N_9550);
nand UO_1396 (O_1396,N_9294,N_9072);
nand UO_1397 (O_1397,N_9530,N_9411);
nand UO_1398 (O_1398,N_9220,N_9531);
or UO_1399 (O_1399,N_9878,N_9676);
nor UO_1400 (O_1400,N_9221,N_9325);
nand UO_1401 (O_1401,N_9922,N_9190);
nor UO_1402 (O_1402,N_9127,N_9601);
nand UO_1403 (O_1403,N_9791,N_9686);
nand UO_1404 (O_1404,N_9194,N_9710);
nor UO_1405 (O_1405,N_9742,N_9904);
or UO_1406 (O_1406,N_9898,N_9622);
nor UO_1407 (O_1407,N_9965,N_9556);
nor UO_1408 (O_1408,N_9656,N_9510);
and UO_1409 (O_1409,N_9811,N_9034);
and UO_1410 (O_1410,N_9604,N_9234);
nor UO_1411 (O_1411,N_9320,N_9326);
and UO_1412 (O_1412,N_9552,N_9821);
or UO_1413 (O_1413,N_9594,N_9957);
or UO_1414 (O_1414,N_9238,N_9457);
nor UO_1415 (O_1415,N_9203,N_9088);
nor UO_1416 (O_1416,N_9390,N_9720);
nand UO_1417 (O_1417,N_9858,N_9192);
or UO_1418 (O_1418,N_9309,N_9934);
nor UO_1419 (O_1419,N_9403,N_9829);
nor UO_1420 (O_1420,N_9005,N_9108);
or UO_1421 (O_1421,N_9383,N_9493);
and UO_1422 (O_1422,N_9271,N_9764);
or UO_1423 (O_1423,N_9786,N_9172);
nand UO_1424 (O_1424,N_9720,N_9920);
nand UO_1425 (O_1425,N_9420,N_9258);
xnor UO_1426 (O_1426,N_9824,N_9982);
nor UO_1427 (O_1427,N_9017,N_9502);
nor UO_1428 (O_1428,N_9269,N_9694);
or UO_1429 (O_1429,N_9657,N_9752);
or UO_1430 (O_1430,N_9469,N_9781);
nand UO_1431 (O_1431,N_9718,N_9948);
and UO_1432 (O_1432,N_9403,N_9393);
and UO_1433 (O_1433,N_9382,N_9663);
nand UO_1434 (O_1434,N_9461,N_9493);
and UO_1435 (O_1435,N_9887,N_9497);
nand UO_1436 (O_1436,N_9266,N_9617);
and UO_1437 (O_1437,N_9366,N_9033);
and UO_1438 (O_1438,N_9315,N_9693);
and UO_1439 (O_1439,N_9238,N_9407);
nor UO_1440 (O_1440,N_9222,N_9463);
and UO_1441 (O_1441,N_9641,N_9459);
nor UO_1442 (O_1442,N_9996,N_9243);
nand UO_1443 (O_1443,N_9158,N_9001);
nand UO_1444 (O_1444,N_9043,N_9654);
nand UO_1445 (O_1445,N_9606,N_9637);
nand UO_1446 (O_1446,N_9783,N_9576);
nand UO_1447 (O_1447,N_9784,N_9725);
xnor UO_1448 (O_1448,N_9345,N_9150);
and UO_1449 (O_1449,N_9354,N_9541);
nor UO_1450 (O_1450,N_9723,N_9844);
nor UO_1451 (O_1451,N_9378,N_9368);
or UO_1452 (O_1452,N_9972,N_9696);
and UO_1453 (O_1453,N_9056,N_9177);
or UO_1454 (O_1454,N_9573,N_9589);
or UO_1455 (O_1455,N_9386,N_9287);
nor UO_1456 (O_1456,N_9335,N_9247);
nand UO_1457 (O_1457,N_9747,N_9840);
nor UO_1458 (O_1458,N_9128,N_9294);
or UO_1459 (O_1459,N_9057,N_9710);
and UO_1460 (O_1460,N_9690,N_9944);
and UO_1461 (O_1461,N_9963,N_9206);
and UO_1462 (O_1462,N_9164,N_9330);
xor UO_1463 (O_1463,N_9749,N_9309);
nor UO_1464 (O_1464,N_9242,N_9072);
and UO_1465 (O_1465,N_9083,N_9690);
nand UO_1466 (O_1466,N_9145,N_9748);
or UO_1467 (O_1467,N_9552,N_9819);
nor UO_1468 (O_1468,N_9465,N_9747);
and UO_1469 (O_1469,N_9240,N_9393);
and UO_1470 (O_1470,N_9908,N_9578);
or UO_1471 (O_1471,N_9083,N_9844);
nand UO_1472 (O_1472,N_9442,N_9640);
or UO_1473 (O_1473,N_9944,N_9275);
and UO_1474 (O_1474,N_9922,N_9993);
nand UO_1475 (O_1475,N_9670,N_9051);
and UO_1476 (O_1476,N_9796,N_9306);
nand UO_1477 (O_1477,N_9334,N_9065);
and UO_1478 (O_1478,N_9550,N_9298);
nor UO_1479 (O_1479,N_9543,N_9998);
nand UO_1480 (O_1480,N_9444,N_9565);
nand UO_1481 (O_1481,N_9557,N_9559);
nand UO_1482 (O_1482,N_9225,N_9285);
or UO_1483 (O_1483,N_9417,N_9251);
and UO_1484 (O_1484,N_9025,N_9656);
or UO_1485 (O_1485,N_9868,N_9717);
nand UO_1486 (O_1486,N_9613,N_9890);
nand UO_1487 (O_1487,N_9962,N_9073);
nand UO_1488 (O_1488,N_9526,N_9276);
xnor UO_1489 (O_1489,N_9993,N_9133);
nand UO_1490 (O_1490,N_9311,N_9746);
or UO_1491 (O_1491,N_9156,N_9173);
or UO_1492 (O_1492,N_9327,N_9576);
and UO_1493 (O_1493,N_9340,N_9354);
nand UO_1494 (O_1494,N_9115,N_9251);
nand UO_1495 (O_1495,N_9333,N_9685);
or UO_1496 (O_1496,N_9212,N_9109);
nor UO_1497 (O_1497,N_9469,N_9731);
or UO_1498 (O_1498,N_9775,N_9171);
nor UO_1499 (O_1499,N_9774,N_9798);
endmodule