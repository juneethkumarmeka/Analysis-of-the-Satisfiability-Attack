module basic_750_5000_1000_5_levels_2xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_26,In_736);
and U1 (N_1,In_401,In_725);
nand U2 (N_2,In_193,In_227);
nand U3 (N_3,In_720,In_36);
or U4 (N_4,In_270,In_595);
or U5 (N_5,In_113,In_32);
nor U6 (N_6,In_271,In_108);
nand U7 (N_7,In_435,In_590);
nand U8 (N_8,In_94,In_541);
or U9 (N_9,In_525,In_417);
or U10 (N_10,In_677,In_218);
and U11 (N_11,In_199,In_705);
and U12 (N_12,In_85,In_150);
and U13 (N_13,In_553,In_33);
nor U14 (N_14,In_416,In_519);
and U15 (N_15,In_578,In_563);
and U16 (N_16,In_548,In_84);
and U17 (N_17,In_302,In_711);
nor U18 (N_18,In_724,In_703);
nand U19 (N_19,In_678,In_247);
nor U20 (N_20,In_122,In_564);
or U21 (N_21,In_687,In_112);
xnor U22 (N_22,In_54,In_344);
or U23 (N_23,In_489,In_430);
or U24 (N_24,In_412,In_371);
and U25 (N_25,In_377,In_597);
nor U26 (N_26,In_614,In_733);
nor U27 (N_27,In_649,In_710);
or U28 (N_28,In_280,In_5);
nand U29 (N_29,In_444,In_305);
nor U30 (N_30,In_605,In_364);
nand U31 (N_31,In_683,In_418);
nor U32 (N_32,In_469,In_49);
nor U33 (N_33,In_447,In_429);
and U34 (N_34,In_507,In_640);
and U35 (N_35,In_537,In_161);
and U36 (N_36,In_496,In_600);
nand U37 (N_37,In_442,In_594);
nand U38 (N_38,In_511,In_482);
and U39 (N_39,In_414,In_410);
nor U40 (N_40,In_27,In_452);
nor U41 (N_41,In_153,In_395);
nand U42 (N_42,In_712,In_249);
or U43 (N_43,In_206,In_77);
and U44 (N_44,In_628,In_319);
nand U45 (N_45,In_251,In_312);
or U46 (N_46,In_556,In_533);
nor U47 (N_47,In_320,In_514);
and U48 (N_48,In_437,In_92);
and U49 (N_49,In_399,In_426);
nand U50 (N_50,In_198,In_722);
and U51 (N_51,In_588,In_627);
and U52 (N_52,In_562,In_528);
or U53 (N_53,In_411,In_635);
or U54 (N_54,In_476,In_680);
and U55 (N_55,In_287,In_236);
nor U56 (N_56,In_689,In_576);
xor U57 (N_57,In_656,In_602);
or U58 (N_58,In_180,In_535);
nand U59 (N_59,In_326,In_532);
or U60 (N_60,In_366,In_168);
or U61 (N_61,In_184,In_645);
or U62 (N_62,In_21,In_70);
or U63 (N_63,In_234,In_453);
nand U64 (N_64,In_598,In_167);
nor U65 (N_65,In_450,In_269);
xnor U66 (N_66,In_531,In_87);
nor U67 (N_67,In_58,In_16);
nand U68 (N_68,In_583,In_373);
or U69 (N_69,In_632,In_730);
and U70 (N_70,In_352,In_672);
and U71 (N_71,In_615,In_299);
and U72 (N_72,In_747,In_455);
and U73 (N_73,In_669,In_370);
and U74 (N_74,In_22,In_498);
nor U75 (N_75,In_291,In_340);
nor U76 (N_76,In_187,In_749);
or U77 (N_77,In_322,In_157);
or U78 (N_78,In_566,In_358);
nand U79 (N_79,In_29,In_580);
nor U80 (N_80,In_443,In_274);
nand U81 (N_81,In_100,In_577);
or U82 (N_82,In_558,In_523);
and U83 (N_83,In_365,In_612);
nor U84 (N_84,In_51,In_59);
nor U85 (N_85,In_509,In_154);
nor U86 (N_86,In_190,In_223);
and U87 (N_87,In_465,In_155);
xor U88 (N_88,In_256,In_132);
nand U89 (N_89,In_698,In_158);
and U90 (N_90,In_494,In_42);
nand U91 (N_91,In_91,In_71);
nand U92 (N_92,In_346,In_50);
nand U93 (N_93,In_125,In_516);
and U94 (N_94,In_93,In_486);
nor U95 (N_95,In_461,In_138);
or U96 (N_96,In_286,In_253);
and U97 (N_97,In_98,In_24);
nand U98 (N_98,In_708,In_679);
or U99 (N_99,In_23,In_436);
nand U100 (N_100,In_502,In_569);
or U101 (N_101,In_464,In_557);
nand U102 (N_102,In_52,In_646);
nand U103 (N_103,In_439,In_409);
and U104 (N_104,In_362,In_263);
xnor U105 (N_105,In_83,In_301);
and U106 (N_106,In_457,In_726);
nand U107 (N_107,In_179,In_428);
nand U108 (N_108,In_636,In_579);
or U109 (N_109,In_473,In_709);
nor U110 (N_110,In_141,In_427);
or U111 (N_111,In_203,In_631);
nand U112 (N_112,In_238,In_6);
and U113 (N_113,In_376,In_232);
nand U114 (N_114,In_729,In_338);
nor U115 (N_115,In_707,In_48);
nor U116 (N_116,In_492,In_652);
and U117 (N_117,In_367,In_647);
nor U118 (N_118,In_466,In_641);
or U119 (N_119,In_369,In_568);
or U120 (N_120,In_723,In_152);
and U121 (N_121,In_147,In_96);
or U122 (N_122,In_262,In_382);
nor U123 (N_123,In_245,In_225);
or U124 (N_124,In_324,In_337);
nand U125 (N_125,In_200,In_34);
or U126 (N_126,In_107,In_611);
nor U127 (N_127,In_480,In_110);
or U128 (N_128,In_695,In_501);
nand U129 (N_129,In_617,In_116);
nor U130 (N_130,In_408,In_420);
nor U131 (N_131,In_375,In_106);
and U132 (N_132,In_446,In_255);
nor U133 (N_133,In_66,In_243);
and U134 (N_134,In_624,In_260);
nor U135 (N_135,In_109,In_570);
and U136 (N_136,In_648,In_214);
or U137 (N_137,In_162,In_146);
or U138 (N_138,In_474,In_304);
nand U139 (N_139,In_294,In_357);
or U140 (N_140,In_172,In_746);
nand U141 (N_141,In_102,In_349);
nor U142 (N_142,In_178,In_35);
nand U143 (N_143,In_675,In_212);
and U144 (N_144,In_37,In_196);
nor U145 (N_145,In_661,In_361);
or U146 (N_146,In_601,In_321);
nand U147 (N_147,In_524,In_385);
and U148 (N_148,In_351,In_504);
nor U149 (N_149,In_117,In_131);
or U150 (N_150,In_651,In_244);
and U151 (N_151,In_252,In_471);
nor U152 (N_152,In_239,In_488);
or U153 (N_153,In_160,In_237);
or U154 (N_154,In_691,In_735);
or U155 (N_155,In_715,In_303);
and U156 (N_156,In_565,In_75);
or U157 (N_157,In_526,In_38);
nand U158 (N_158,In_438,In_462);
nor U159 (N_159,In_663,In_12);
nor U160 (N_160,In_396,In_620);
nand U161 (N_161,In_14,In_622);
nand U162 (N_162,In_194,In_582);
nand U163 (N_163,In_727,In_265);
and U164 (N_164,In_630,In_7);
or U165 (N_165,In_332,In_667);
nor U166 (N_166,In_275,In_419);
xor U167 (N_167,In_470,In_549);
nand U168 (N_168,In_555,In_716);
or U169 (N_169,In_89,In_356);
nor U170 (N_170,In_10,In_266);
and U171 (N_171,In_596,In_387);
or U172 (N_172,In_134,In_475);
or U173 (N_173,In_719,In_374);
and U174 (N_174,In_637,In_378);
and U175 (N_175,In_544,In_19);
nor U176 (N_176,In_115,In_404);
nand U177 (N_177,In_581,In_224);
nor U178 (N_178,In_688,In_664);
nand U179 (N_179,In_561,In_629);
nor U180 (N_180,In_330,In_254);
and U181 (N_181,In_503,In_573);
nor U182 (N_182,In_534,In_159);
or U183 (N_183,In_662,In_542);
nor U184 (N_184,In_120,In_53);
or U185 (N_185,In_311,In_217);
and U186 (N_186,In_642,In_103);
and U187 (N_187,In_88,In_406);
xor U188 (N_188,In_295,In_339);
nand U189 (N_189,In_413,In_522);
and U190 (N_190,In_128,In_621);
nor U191 (N_191,In_717,In_449);
and U192 (N_192,In_171,In_384);
or U193 (N_193,In_500,In_267);
or U194 (N_194,In_659,In_18);
and U195 (N_195,In_101,In_560);
nor U196 (N_196,In_104,In_434);
nor U197 (N_197,In_79,In_281);
and U198 (N_198,In_381,In_572);
or U199 (N_199,In_250,In_741);
or U200 (N_200,In_316,In_634);
nor U201 (N_201,In_676,In_118);
nor U202 (N_202,In_183,In_610);
nor U203 (N_203,In_195,In_421);
nor U204 (N_204,In_424,In_97);
or U205 (N_205,In_201,In_529);
or U206 (N_206,In_415,In_86);
nand U207 (N_207,In_589,In_713);
nand U208 (N_208,In_348,In_30);
or U209 (N_209,In_142,In_379);
and U210 (N_210,In_425,In_701);
and U211 (N_211,In_264,In_55);
or U212 (N_212,In_61,In_3);
and U213 (N_213,In_175,In_586);
or U214 (N_214,In_273,In_306);
or U215 (N_215,In_282,In_56);
or U216 (N_216,In_397,In_28);
and U217 (N_217,In_228,In_111);
or U218 (N_218,In_226,In_495);
and U219 (N_219,In_389,In_78);
or U220 (N_220,In_657,In_403);
nand U221 (N_221,In_137,In_65);
and U222 (N_222,In_284,In_242);
nor U223 (N_223,In_173,In_314);
or U224 (N_224,In_456,In_686);
nor U225 (N_225,In_731,In_259);
nand U226 (N_226,In_213,In_139);
nand U227 (N_227,In_571,In_734);
or U228 (N_228,In_459,In_650);
and U229 (N_229,In_44,In_169);
nor U230 (N_230,In_697,In_329);
nand U231 (N_231,In_547,In_334);
and U232 (N_232,In_441,In_394);
or U233 (N_233,In_230,In_292);
or U234 (N_234,In_665,In_57);
or U235 (N_235,In_174,In_388);
or U236 (N_236,In_658,In_398);
nand U237 (N_237,In_283,In_354);
nor U238 (N_238,In_276,In_221);
nor U239 (N_239,In_95,In_481);
nor U240 (N_240,In_74,In_170);
nor U241 (N_241,In_353,In_467);
or U242 (N_242,In_191,In_550);
or U243 (N_243,In_240,In_743);
and U244 (N_244,In_129,In_740);
nand U245 (N_245,In_81,In_472);
nand U246 (N_246,In_317,In_325);
nor U247 (N_247,In_623,In_653);
nand U248 (N_248,In_114,In_99);
and U249 (N_249,In_335,In_638);
nor U250 (N_250,In_606,In_261);
nand U251 (N_251,In_402,In_197);
nor U252 (N_252,In_391,In_422);
xor U253 (N_253,In_738,In_219);
nand U254 (N_254,In_4,In_593);
and U255 (N_255,In_592,In_136);
or U256 (N_256,In_124,In_510);
nor U257 (N_257,In_490,In_323);
nand U258 (N_258,In_506,In_235);
or U259 (N_259,In_655,In_293);
xor U260 (N_260,In_121,In_135);
nor U261 (N_261,In_505,In_350);
and U262 (N_262,In_15,In_90);
and U263 (N_263,In_17,In_744);
or U264 (N_264,In_468,In_432);
or U265 (N_265,In_60,In_258);
and U266 (N_266,In_204,In_297);
nand U267 (N_267,In_493,In_248);
xor U268 (N_268,In_619,In_508);
nor U269 (N_269,In_451,In_666);
nand U270 (N_270,In_718,In_278);
nand U271 (N_271,In_690,In_298);
nor U272 (N_272,In_372,In_164);
nand U273 (N_273,In_540,In_296);
and U274 (N_274,In_309,In_11);
or U275 (N_275,In_654,In_315);
nand U276 (N_276,In_559,In_272);
and U277 (N_277,In_308,In_599);
nand U278 (N_278,In_290,In_737);
or U279 (N_279,In_328,In_47);
or U280 (N_280,In_554,In_68);
or U281 (N_281,In_8,In_231);
or U282 (N_282,In_608,In_673);
nand U283 (N_283,In_748,In_706);
or U284 (N_284,In_512,In_518);
and U285 (N_285,In_491,In_479);
and U286 (N_286,In_313,In_43);
or U287 (N_287,In_182,In_355);
nand U288 (N_288,In_268,In_538);
nand U289 (N_289,In_127,In_229);
nor U290 (N_290,In_202,In_386);
nand U291 (N_291,In_431,In_714);
nor U292 (N_292,In_625,In_1);
nor U293 (N_293,In_343,In_336);
nand U294 (N_294,In_543,In_407);
nand U295 (N_295,In_591,In_463);
nand U296 (N_296,In_392,In_545);
and U297 (N_297,In_186,In_359);
nand U298 (N_298,In_513,In_9);
or U299 (N_299,In_20,In_674);
nor U300 (N_300,In_307,In_177);
and U301 (N_301,In_575,In_63);
or U302 (N_302,In_693,In_460);
nand U303 (N_303,In_660,In_144);
xnor U304 (N_304,In_520,In_380);
xor U305 (N_305,In_13,In_105);
and U306 (N_306,In_208,In_285);
nor U307 (N_307,In_682,In_433);
nand U308 (N_308,In_210,In_25);
nor U309 (N_309,In_41,In_2);
nand U310 (N_310,In_166,In_0);
or U311 (N_311,In_732,In_458);
or U312 (N_312,In_448,In_644);
or U313 (N_313,In_140,In_216);
nand U314 (N_314,In_477,In_185);
and U315 (N_315,In_64,In_345);
nand U316 (N_316,In_211,In_241);
or U317 (N_317,In_45,In_143);
or U318 (N_318,In_222,In_618);
nand U319 (N_319,In_692,In_668);
and U320 (N_320,In_745,In_574);
nor U321 (N_321,In_205,In_246);
or U322 (N_322,In_633,In_126);
nand U323 (N_323,In_82,In_567);
and U324 (N_324,In_445,In_497);
and U325 (N_325,In_499,In_165);
and U326 (N_326,In_123,In_310);
or U327 (N_327,In_188,In_288);
nor U328 (N_328,In_530,In_699);
nor U329 (N_329,In_220,In_728);
or U330 (N_330,In_584,In_696);
and U331 (N_331,In_721,In_639);
nand U332 (N_332,In_423,In_189);
nor U333 (N_333,In_393,In_149);
and U334 (N_334,In_484,In_76);
nor U335 (N_335,In_483,In_604);
or U336 (N_336,In_626,In_62);
nor U337 (N_337,In_670,In_616);
or U338 (N_338,In_279,In_681);
nor U339 (N_339,In_400,In_609);
nand U340 (N_340,In_342,In_739);
nor U341 (N_341,In_587,In_454);
or U342 (N_342,In_704,In_207);
nand U343 (N_343,In_607,In_39);
nand U344 (N_344,In_192,In_67);
and U345 (N_345,In_390,In_347);
nand U346 (N_346,In_552,In_333);
or U347 (N_347,In_440,In_515);
or U348 (N_348,In_536,In_148);
and U349 (N_349,In_603,In_546);
nor U350 (N_350,In_685,In_702);
or U351 (N_351,In_163,In_80);
nand U352 (N_352,In_383,In_613);
nor U353 (N_353,In_363,In_341);
nand U354 (N_354,In_539,In_327);
nand U355 (N_355,In_300,In_145);
and U356 (N_356,In_72,In_69);
nand U357 (N_357,In_684,In_151);
nor U358 (N_358,In_527,In_31);
or U359 (N_359,In_487,In_73);
and U360 (N_360,In_694,In_478);
nand U361 (N_361,In_643,In_215);
and U362 (N_362,In_585,In_331);
or U363 (N_363,In_289,In_517);
and U364 (N_364,In_257,In_485);
xnor U365 (N_365,In_176,In_521);
nor U366 (N_366,In_233,In_130);
nor U367 (N_367,In_46,In_133);
nor U368 (N_368,In_360,In_318);
nand U369 (N_369,In_181,In_671);
and U370 (N_370,In_277,In_405);
and U371 (N_371,In_368,In_700);
and U372 (N_372,In_156,In_40);
and U373 (N_373,In_551,In_742);
or U374 (N_374,In_209,In_119);
nor U375 (N_375,In_711,In_349);
and U376 (N_376,In_510,In_7);
and U377 (N_377,In_87,In_345);
nand U378 (N_378,In_709,In_541);
xnor U379 (N_379,In_604,In_306);
and U380 (N_380,In_715,In_231);
and U381 (N_381,In_647,In_520);
nand U382 (N_382,In_697,In_493);
nand U383 (N_383,In_142,In_119);
or U384 (N_384,In_7,In_508);
or U385 (N_385,In_240,In_409);
nor U386 (N_386,In_665,In_161);
nand U387 (N_387,In_37,In_485);
or U388 (N_388,In_418,In_214);
nor U389 (N_389,In_597,In_266);
or U390 (N_390,In_74,In_28);
or U391 (N_391,In_519,In_291);
and U392 (N_392,In_575,In_226);
nor U393 (N_393,In_97,In_380);
and U394 (N_394,In_640,In_565);
nand U395 (N_395,In_715,In_682);
or U396 (N_396,In_229,In_466);
nor U397 (N_397,In_397,In_742);
nor U398 (N_398,In_161,In_488);
nand U399 (N_399,In_151,In_304);
or U400 (N_400,In_541,In_95);
nor U401 (N_401,In_526,In_671);
and U402 (N_402,In_522,In_119);
or U403 (N_403,In_412,In_293);
or U404 (N_404,In_160,In_252);
and U405 (N_405,In_73,In_386);
nor U406 (N_406,In_312,In_735);
nand U407 (N_407,In_89,In_488);
and U408 (N_408,In_411,In_284);
nand U409 (N_409,In_286,In_444);
and U410 (N_410,In_202,In_177);
and U411 (N_411,In_252,In_72);
nor U412 (N_412,In_435,In_602);
and U413 (N_413,In_356,In_265);
nor U414 (N_414,In_428,In_626);
nand U415 (N_415,In_182,In_655);
or U416 (N_416,In_362,In_70);
nand U417 (N_417,In_671,In_361);
nand U418 (N_418,In_547,In_379);
or U419 (N_419,In_290,In_623);
and U420 (N_420,In_35,In_404);
and U421 (N_421,In_31,In_328);
or U422 (N_422,In_586,In_554);
or U423 (N_423,In_326,In_738);
nand U424 (N_424,In_434,In_216);
or U425 (N_425,In_643,In_226);
nor U426 (N_426,In_162,In_361);
nand U427 (N_427,In_534,In_218);
nor U428 (N_428,In_484,In_714);
nand U429 (N_429,In_235,In_624);
and U430 (N_430,In_735,In_332);
nor U431 (N_431,In_151,In_626);
and U432 (N_432,In_277,In_749);
nand U433 (N_433,In_441,In_319);
and U434 (N_434,In_580,In_525);
or U435 (N_435,In_177,In_446);
nand U436 (N_436,In_141,In_164);
nand U437 (N_437,In_215,In_8);
and U438 (N_438,In_557,In_544);
nor U439 (N_439,In_223,In_265);
nand U440 (N_440,In_126,In_398);
and U441 (N_441,In_494,In_50);
xnor U442 (N_442,In_392,In_690);
or U443 (N_443,In_709,In_108);
or U444 (N_444,In_7,In_696);
and U445 (N_445,In_148,In_662);
and U446 (N_446,In_19,In_183);
nand U447 (N_447,In_196,In_203);
nand U448 (N_448,In_261,In_25);
and U449 (N_449,In_711,In_215);
and U450 (N_450,In_161,In_706);
or U451 (N_451,In_226,In_119);
nand U452 (N_452,In_543,In_322);
and U453 (N_453,In_619,In_659);
nand U454 (N_454,In_732,In_135);
nor U455 (N_455,In_670,In_509);
and U456 (N_456,In_226,In_162);
nand U457 (N_457,In_463,In_208);
nand U458 (N_458,In_208,In_236);
nand U459 (N_459,In_9,In_157);
nand U460 (N_460,In_1,In_112);
nor U461 (N_461,In_368,In_594);
or U462 (N_462,In_176,In_695);
and U463 (N_463,In_705,In_549);
xor U464 (N_464,In_89,In_678);
nor U465 (N_465,In_21,In_33);
and U466 (N_466,In_175,In_191);
and U467 (N_467,In_36,In_481);
xnor U468 (N_468,In_452,In_210);
nand U469 (N_469,In_15,In_128);
nor U470 (N_470,In_160,In_445);
or U471 (N_471,In_104,In_542);
and U472 (N_472,In_305,In_83);
nor U473 (N_473,In_587,In_445);
or U474 (N_474,In_140,In_411);
nor U475 (N_475,In_630,In_289);
and U476 (N_476,In_707,In_393);
nor U477 (N_477,In_422,In_320);
and U478 (N_478,In_180,In_709);
nor U479 (N_479,In_228,In_460);
and U480 (N_480,In_494,In_211);
nand U481 (N_481,In_552,In_708);
or U482 (N_482,In_258,In_100);
nand U483 (N_483,In_484,In_738);
or U484 (N_484,In_65,In_119);
nor U485 (N_485,In_576,In_575);
nand U486 (N_486,In_740,In_604);
or U487 (N_487,In_576,In_555);
or U488 (N_488,In_344,In_114);
nor U489 (N_489,In_633,In_579);
or U490 (N_490,In_534,In_606);
and U491 (N_491,In_407,In_278);
or U492 (N_492,In_112,In_364);
nand U493 (N_493,In_738,In_510);
nand U494 (N_494,In_34,In_693);
nand U495 (N_495,In_88,In_683);
nor U496 (N_496,In_609,In_366);
nor U497 (N_497,In_672,In_13);
nand U498 (N_498,In_256,In_553);
and U499 (N_499,In_642,In_256);
and U500 (N_500,In_475,In_415);
or U501 (N_501,In_574,In_503);
or U502 (N_502,In_404,In_84);
nor U503 (N_503,In_449,In_194);
nand U504 (N_504,In_742,In_60);
nand U505 (N_505,In_180,In_658);
and U506 (N_506,In_307,In_187);
nor U507 (N_507,In_121,In_197);
or U508 (N_508,In_636,In_164);
nor U509 (N_509,In_659,In_651);
nor U510 (N_510,In_706,In_633);
and U511 (N_511,In_595,In_606);
nor U512 (N_512,In_213,In_566);
xor U513 (N_513,In_117,In_517);
nand U514 (N_514,In_726,In_45);
nor U515 (N_515,In_577,In_203);
nand U516 (N_516,In_399,In_79);
nor U517 (N_517,In_366,In_720);
and U518 (N_518,In_147,In_307);
nor U519 (N_519,In_725,In_535);
and U520 (N_520,In_528,In_288);
nor U521 (N_521,In_187,In_296);
nand U522 (N_522,In_565,In_132);
or U523 (N_523,In_454,In_480);
nor U524 (N_524,In_572,In_301);
nand U525 (N_525,In_464,In_301);
nor U526 (N_526,In_684,In_595);
xnor U527 (N_527,In_405,In_546);
nor U528 (N_528,In_128,In_671);
and U529 (N_529,In_607,In_180);
xnor U530 (N_530,In_271,In_289);
nor U531 (N_531,In_549,In_107);
nor U532 (N_532,In_315,In_457);
nand U533 (N_533,In_388,In_192);
or U534 (N_534,In_399,In_688);
or U535 (N_535,In_613,In_171);
nor U536 (N_536,In_71,In_4);
nor U537 (N_537,In_450,In_10);
nand U538 (N_538,In_439,In_310);
and U539 (N_539,In_631,In_103);
nor U540 (N_540,In_283,In_293);
nor U541 (N_541,In_510,In_435);
and U542 (N_542,In_739,In_12);
or U543 (N_543,In_210,In_81);
nor U544 (N_544,In_615,In_99);
nor U545 (N_545,In_513,In_195);
or U546 (N_546,In_96,In_277);
or U547 (N_547,In_658,In_445);
nor U548 (N_548,In_65,In_650);
nand U549 (N_549,In_657,In_137);
nor U550 (N_550,In_199,In_217);
or U551 (N_551,In_494,In_287);
or U552 (N_552,In_137,In_189);
and U553 (N_553,In_288,In_521);
nor U554 (N_554,In_685,In_179);
nand U555 (N_555,In_537,In_106);
or U556 (N_556,In_549,In_401);
nand U557 (N_557,In_350,In_725);
nand U558 (N_558,In_460,In_644);
or U559 (N_559,In_705,In_374);
nand U560 (N_560,In_314,In_135);
xor U561 (N_561,In_343,In_643);
and U562 (N_562,In_584,In_466);
nand U563 (N_563,In_169,In_573);
nand U564 (N_564,In_708,In_690);
and U565 (N_565,In_477,In_231);
nor U566 (N_566,In_287,In_636);
nand U567 (N_567,In_504,In_630);
nor U568 (N_568,In_654,In_527);
nor U569 (N_569,In_104,In_109);
nor U570 (N_570,In_546,In_254);
nand U571 (N_571,In_575,In_632);
nand U572 (N_572,In_416,In_47);
or U573 (N_573,In_88,In_471);
nor U574 (N_574,In_272,In_41);
nor U575 (N_575,In_157,In_741);
nor U576 (N_576,In_336,In_82);
or U577 (N_577,In_529,In_730);
or U578 (N_578,In_531,In_597);
nor U579 (N_579,In_282,In_124);
nor U580 (N_580,In_309,In_231);
nand U581 (N_581,In_353,In_382);
and U582 (N_582,In_338,In_718);
nor U583 (N_583,In_725,In_603);
nor U584 (N_584,In_59,In_475);
and U585 (N_585,In_407,In_167);
and U586 (N_586,In_460,In_625);
and U587 (N_587,In_296,In_314);
and U588 (N_588,In_467,In_738);
or U589 (N_589,In_63,In_26);
nor U590 (N_590,In_551,In_367);
or U591 (N_591,In_245,In_208);
and U592 (N_592,In_114,In_667);
nor U593 (N_593,In_742,In_400);
nor U594 (N_594,In_223,In_295);
nand U595 (N_595,In_185,In_324);
nand U596 (N_596,In_2,In_405);
or U597 (N_597,In_647,In_229);
nand U598 (N_598,In_578,In_684);
or U599 (N_599,In_517,In_515);
and U600 (N_600,In_429,In_674);
nand U601 (N_601,In_145,In_390);
nor U602 (N_602,In_418,In_386);
nor U603 (N_603,In_405,In_623);
or U604 (N_604,In_175,In_357);
and U605 (N_605,In_483,In_404);
nand U606 (N_606,In_685,In_160);
nand U607 (N_607,In_187,In_124);
or U608 (N_608,In_425,In_616);
and U609 (N_609,In_649,In_439);
or U610 (N_610,In_633,In_242);
nor U611 (N_611,In_700,In_80);
nand U612 (N_612,In_155,In_430);
nand U613 (N_613,In_451,In_372);
and U614 (N_614,In_615,In_376);
nor U615 (N_615,In_58,In_52);
and U616 (N_616,In_327,In_339);
and U617 (N_617,In_605,In_85);
or U618 (N_618,In_33,In_194);
nand U619 (N_619,In_73,In_400);
or U620 (N_620,In_366,In_746);
or U621 (N_621,In_658,In_560);
or U622 (N_622,In_356,In_626);
and U623 (N_623,In_113,In_425);
or U624 (N_624,In_502,In_667);
nor U625 (N_625,In_562,In_32);
and U626 (N_626,In_473,In_2);
nand U627 (N_627,In_152,In_335);
nor U628 (N_628,In_383,In_625);
nor U629 (N_629,In_297,In_329);
nor U630 (N_630,In_495,In_442);
nor U631 (N_631,In_744,In_273);
and U632 (N_632,In_75,In_92);
and U633 (N_633,In_183,In_709);
and U634 (N_634,In_573,In_704);
nand U635 (N_635,In_679,In_403);
nand U636 (N_636,In_689,In_106);
nand U637 (N_637,In_427,In_673);
nand U638 (N_638,In_545,In_300);
and U639 (N_639,In_489,In_410);
nor U640 (N_640,In_166,In_309);
nor U641 (N_641,In_586,In_504);
nor U642 (N_642,In_251,In_599);
or U643 (N_643,In_473,In_98);
or U644 (N_644,In_124,In_266);
and U645 (N_645,In_550,In_649);
or U646 (N_646,In_658,In_417);
nor U647 (N_647,In_513,In_192);
nand U648 (N_648,In_291,In_330);
nand U649 (N_649,In_209,In_478);
or U650 (N_650,In_50,In_748);
nor U651 (N_651,In_544,In_593);
nand U652 (N_652,In_306,In_689);
or U653 (N_653,In_397,In_670);
or U654 (N_654,In_565,In_534);
nor U655 (N_655,In_100,In_39);
and U656 (N_656,In_673,In_726);
nor U657 (N_657,In_386,In_215);
nor U658 (N_658,In_580,In_283);
and U659 (N_659,In_704,In_103);
nor U660 (N_660,In_683,In_500);
nand U661 (N_661,In_110,In_687);
and U662 (N_662,In_355,In_144);
and U663 (N_663,In_61,In_230);
or U664 (N_664,In_515,In_439);
or U665 (N_665,In_113,In_560);
and U666 (N_666,In_616,In_630);
nand U667 (N_667,In_220,In_333);
or U668 (N_668,In_521,In_174);
or U669 (N_669,In_731,In_330);
nor U670 (N_670,In_450,In_108);
or U671 (N_671,In_695,In_598);
nand U672 (N_672,In_215,In_129);
and U673 (N_673,In_346,In_117);
nand U674 (N_674,In_338,In_517);
xor U675 (N_675,In_485,In_695);
and U676 (N_676,In_331,In_569);
nor U677 (N_677,In_82,In_494);
nor U678 (N_678,In_476,In_535);
xor U679 (N_679,In_148,In_139);
or U680 (N_680,In_327,In_211);
nand U681 (N_681,In_484,In_504);
nor U682 (N_682,In_462,In_36);
or U683 (N_683,In_37,In_266);
and U684 (N_684,In_385,In_145);
or U685 (N_685,In_96,In_199);
nor U686 (N_686,In_716,In_522);
nand U687 (N_687,In_668,In_725);
nor U688 (N_688,In_458,In_570);
or U689 (N_689,In_258,In_565);
nor U690 (N_690,In_168,In_35);
nor U691 (N_691,In_640,In_502);
and U692 (N_692,In_608,In_716);
nand U693 (N_693,In_193,In_545);
and U694 (N_694,In_371,In_537);
or U695 (N_695,In_379,In_314);
nor U696 (N_696,In_509,In_59);
nand U697 (N_697,In_101,In_598);
nor U698 (N_698,In_157,In_316);
nand U699 (N_699,In_219,In_305);
nor U700 (N_700,In_281,In_408);
nand U701 (N_701,In_361,In_59);
nor U702 (N_702,In_384,In_373);
nand U703 (N_703,In_166,In_553);
and U704 (N_704,In_409,In_184);
or U705 (N_705,In_584,In_19);
nor U706 (N_706,In_736,In_517);
nand U707 (N_707,In_476,In_358);
nor U708 (N_708,In_121,In_133);
nand U709 (N_709,In_239,In_28);
or U710 (N_710,In_565,In_572);
and U711 (N_711,In_619,In_311);
and U712 (N_712,In_258,In_356);
nor U713 (N_713,In_666,In_610);
and U714 (N_714,In_389,In_377);
and U715 (N_715,In_412,In_288);
or U716 (N_716,In_151,In_682);
and U717 (N_717,In_301,In_447);
nand U718 (N_718,In_23,In_383);
and U719 (N_719,In_415,In_337);
and U720 (N_720,In_476,In_173);
nor U721 (N_721,In_213,In_370);
nor U722 (N_722,In_452,In_636);
nand U723 (N_723,In_131,In_357);
nand U724 (N_724,In_636,In_523);
or U725 (N_725,In_355,In_221);
and U726 (N_726,In_436,In_694);
or U727 (N_727,In_163,In_114);
xor U728 (N_728,In_496,In_219);
or U729 (N_729,In_169,In_471);
nand U730 (N_730,In_114,In_66);
or U731 (N_731,In_649,In_70);
or U732 (N_732,In_351,In_47);
and U733 (N_733,In_642,In_696);
and U734 (N_734,In_94,In_76);
nand U735 (N_735,In_24,In_603);
nor U736 (N_736,In_372,In_63);
and U737 (N_737,In_419,In_207);
xor U738 (N_738,In_619,In_650);
or U739 (N_739,In_344,In_394);
or U740 (N_740,In_693,In_156);
and U741 (N_741,In_627,In_746);
nor U742 (N_742,In_243,In_320);
nand U743 (N_743,In_160,In_482);
xnor U744 (N_744,In_27,In_615);
or U745 (N_745,In_741,In_510);
nor U746 (N_746,In_716,In_51);
or U747 (N_747,In_92,In_736);
or U748 (N_748,In_607,In_19);
nor U749 (N_749,In_74,In_273);
and U750 (N_750,In_376,In_543);
nand U751 (N_751,In_327,In_712);
nor U752 (N_752,In_495,In_366);
and U753 (N_753,In_712,In_155);
xor U754 (N_754,In_746,In_165);
or U755 (N_755,In_88,In_255);
nor U756 (N_756,In_475,In_115);
or U757 (N_757,In_366,In_361);
and U758 (N_758,In_426,In_670);
or U759 (N_759,In_699,In_437);
nor U760 (N_760,In_316,In_222);
and U761 (N_761,In_479,In_405);
nor U762 (N_762,In_169,In_70);
or U763 (N_763,In_1,In_218);
or U764 (N_764,In_234,In_61);
or U765 (N_765,In_252,In_737);
xnor U766 (N_766,In_7,In_315);
and U767 (N_767,In_294,In_98);
nand U768 (N_768,In_196,In_66);
nor U769 (N_769,In_176,In_186);
or U770 (N_770,In_50,In_731);
nor U771 (N_771,In_549,In_301);
and U772 (N_772,In_744,In_435);
nand U773 (N_773,In_319,In_24);
or U774 (N_774,In_204,In_421);
nor U775 (N_775,In_385,In_141);
and U776 (N_776,In_531,In_32);
nor U777 (N_777,In_33,In_452);
nor U778 (N_778,In_170,In_231);
nand U779 (N_779,In_288,In_269);
and U780 (N_780,In_580,In_595);
and U781 (N_781,In_425,In_92);
nor U782 (N_782,In_96,In_478);
and U783 (N_783,In_32,In_141);
or U784 (N_784,In_397,In_274);
and U785 (N_785,In_474,In_135);
and U786 (N_786,In_468,In_91);
nor U787 (N_787,In_308,In_18);
or U788 (N_788,In_356,In_195);
and U789 (N_789,In_633,In_540);
or U790 (N_790,In_73,In_374);
nand U791 (N_791,In_79,In_316);
nor U792 (N_792,In_705,In_262);
nor U793 (N_793,In_173,In_707);
and U794 (N_794,In_227,In_200);
nor U795 (N_795,In_503,In_72);
or U796 (N_796,In_730,In_227);
or U797 (N_797,In_489,In_706);
nand U798 (N_798,In_567,In_615);
nand U799 (N_799,In_577,In_284);
nor U800 (N_800,In_549,In_748);
nor U801 (N_801,In_102,In_175);
or U802 (N_802,In_94,In_508);
nor U803 (N_803,In_678,In_268);
nor U804 (N_804,In_585,In_65);
and U805 (N_805,In_447,In_1);
and U806 (N_806,In_399,In_265);
nor U807 (N_807,In_427,In_527);
and U808 (N_808,In_162,In_458);
or U809 (N_809,In_215,In_693);
nor U810 (N_810,In_296,In_569);
or U811 (N_811,In_112,In_547);
or U812 (N_812,In_24,In_488);
nor U813 (N_813,In_494,In_132);
and U814 (N_814,In_204,In_69);
or U815 (N_815,In_533,In_247);
and U816 (N_816,In_8,In_430);
nor U817 (N_817,In_679,In_49);
nand U818 (N_818,In_418,In_376);
nor U819 (N_819,In_41,In_262);
or U820 (N_820,In_466,In_559);
nor U821 (N_821,In_353,In_527);
or U822 (N_822,In_574,In_409);
and U823 (N_823,In_406,In_182);
xnor U824 (N_824,In_656,In_8);
xnor U825 (N_825,In_500,In_231);
nand U826 (N_826,In_311,In_338);
or U827 (N_827,In_583,In_544);
and U828 (N_828,In_620,In_471);
nand U829 (N_829,In_425,In_335);
nor U830 (N_830,In_368,In_555);
nand U831 (N_831,In_475,In_185);
or U832 (N_832,In_131,In_467);
nor U833 (N_833,In_124,In_634);
nand U834 (N_834,In_7,In_342);
nand U835 (N_835,In_408,In_589);
and U836 (N_836,In_384,In_620);
and U837 (N_837,In_208,In_222);
nand U838 (N_838,In_8,In_164);
nor U839 (N_839,In_147,In_722);
and U840 (N_840,In_5,In_165);
xor U841 (N_841,In_746,In_300);
nand U842 (N_842,In_515,In_194);
or U843 (N_843,In_740,In_361);
or U844 (N_844,In_651,In_338);
and U845 (N_845,In_127,In_643);
or U846 (N_846,In_505,In_219);
or U847 (N_847,In_538,In_340);
nor U848 (N_848,In_206,In_338);
nand U849 (N_849,In_478,In_104);
or U850 (N_850,In_439,In_740);
nor U851 (N_851,In_699,In_700);
and U852 (N_852,In_134,In_143);
or U853 (N_853,In_613,In_706);
nor U854 (N_854,In_646,In_323);
or U855 (N_855,In_108,In_480);
nor U856 (N_856,In_294,In_125);
and U857 (N_857,In_456,In_69);
or U858 (N_858,In_429,In_324);
nand U859 (N_859,In_713,In_210);
nand U860 (N_860,In_230,In_444);
nand U861 (N_861,In_681,In_572);
nand U862 (N_862,In_195,In_567);
nand U863 (N_863,In_14,In_463);
nor U864 (N_864,In_671,In_236);
or U865 (N_865,In_586,In_174);
or U866 (N_866,In_322,In_121);
nor U867 (N_867,In_157,In_87);
nor U868 (N_868,In_384,In_417);
xor U869 (N_869,In_407,In_3);
and U870 (N_870,In_533,In_46);
and U871 (N_871,In_135,In_601);
xnor U872 (N_872,In_169,In_236);
and U873 (N_873,In_24,In_270);
nor U874 (N_874,In_625,In_358);
or U875 (N_875,In_356,In_80);
nor U876 (N_876,In_483,In_202);
and U877 (N_877,In_106,In_225);
nand U878 (N_878,In_441,In_150);
and U879 (N_879,In_200,In_356);
or U880 (N_880,In_54,In_473);
nor U881 (N_881,In_135,In_501);
and U882 (N_882,In_523,In_21);
nor U883 (N_883,In_107,In_748);
nand U884 (N_884,In_730,In_338);
nor U885 (N_885,In_275,In_529);
nand U886 (N_886,In_348,In_631);
nand U887 (N_887,In_321,In_174);
nor U888 (N_888,In_658,In_670);
or U889 (N_889,In_324,In_310);
nand U890 (N_890,In_431,In_223);
nor U891 (N_891,In_180,In_237);
nand U892 (N_892,In_629,In_309);
or U893 (N_893,In_10,In_742);
nor U894 (N_894,In_723,In_164);
nor U895 (N_895,In_739,In_456);
nor U896 (N_896,In_726,In_49);
or U897 (N_897,In_378,In_55);
nor U898 (N_898,In_629,In_436);
nand U899 (N_899,In_149,In_51);
nand U900 (N_900,In_713,In_163);
nor U901 (N_901,In_140,In_291);
and U902 (N_902,In_218,In_191);
nor U903 (N_903,In_414,In_561);
and U904 (N_904,In_243,In_455);
nand U905 (N_905,In_202,In_96);
or U906 (N_906,In_194,In_737);
nand U907 (N_907,In_719,In_352);
and U908 (N_908,In_117,In_147);
nand U909 (N_909,In_730,In_425);
or U910 (N_910,In_714,In_393);
and U911 (N_911,In_725,In_138);
nor U912 (N_912,In_696,In_244);
or U913 (N_913,In_527,In_185);
nor U914 (N_914,In_60,In_262);
nor U915 (N_915,In_499,In_436);
nand U916 (N_916,In_309,In_10);
xor U917 (N_917,In_658,In_711);
or U918 (N_918,In_169,In_709);
xor U919 (N_919,In_169,In_322);
and U920 (N_920,In_47,In_707);
nor U921 (N_921,In_322,In_222);
nor U922 (N_922,In_344,In_170);
and U923 (N_923,In_611,In_507);
nor U924 (N_924,In_271,In_401);
and U925 (N_925,In_497,In_567);
nor U926 (N_926,In_213,In_712);
nand U927 (N_927,In_626,In_217);
and U928 (N_928,In_682,In_285);
or U929 (N_929,In_156,In_580);
nand U930 (N_930,In_439,In_687);
or U931 (N_931,In_591,In_43);
nand U932 (N_932,In_426,In_437);
or U933 (N_933,In_453,In_362);
or U934 (N_934,In_265,In_539);
or U935 (N_935,In_596,In_573);
nand U936 (N_936,In_696,In_280);
nand U937 (N_937,In_502,In_335);
nand U938 (N_938,In_567,In_619);
or U939 (N_939,In_352,In_95);
or U940 (N_940,In_504,In_100);
or U941 (N_941,In_581,In_23);
or U942 (N_942,In_390,In_695);
nand U943 (N_943,In_733,In_282);
and U944 (N_944,In_670,In_225);
nand U945 (N_945,In_143,In_150);
nand U946 (N_946,In_394,In_70);
nor U947 (N_947,In_376,In_364);
nor U948 (N_948,In_669,In_135);
and U949 (N_949,In_266,In_224);
and U950 (N_950,In_633,In_600);
nand U951 (N_951,In_373,In_215);
nand U952 (N_952,In_98,In_618);
xnor U953 (N_953,In_620,In_518);
and U954 (N_954,In_155,In_561);
nor U955 (N_955,In_293,In_1);
or U956 (N_956,In_271,In_747);
nand U957 (N_957,In_483,In_234);
nor U958 (N_958,In_294,In_599);
nand U959 (N_959,In_314,In_414);
nand U960 (N_960,In_133,In_673);
nand U961 (N_961,In_108,In_202);
nor U962 (N_962,In_471,In_677);
and U963 (N_963,In_597,In_288);
nand U964 (N_964,In_217,In_639);
nand U965 (N_965,In_148,In_746);
nand U966 (N_966,In_478,In_133);
nor U967 (N_967,In_184,In_167);
nand U968 (N_968,In_140,In_220);
and U969 (N_969,In_683,In_40);
or U970 (N_970,In_457,In_373);
nand U971 (N_971,In_109,In_126);
or U972 (N_972,In_96,In_78);
nor U973 (N_973,In_488,In_555);
and U974 (N_974,In_31,In_256);
nor U975 (N_975,In_291,In_124);
nand U976 (N_976,In_628,In_239);
or U977 (N_977,In_99,In_553);
and U978 (N_978,In_178,In_611);
and U979 (N_979,In_494,In_285);
and U980 (N_980,In_395,In_630);
nor U981 (N_981,In_414,In_625);
or U982 (N_982,In_491,In_387);
and U983 (N_983,In_609,In_16);
nand U984 (N_984,In_309,In_604);
or U985 (N_985,In_486,In_539);
xor U986 (N_986,In_300,In_249);
and U987 (N_987,In_358,In_458);
or U988 (N_988,In_121,In_497);
or U989 (N_989,In_14,In_134);
nor U990 (N_990,In_393,In_185);
or U991 (N_991,In_11,In_455);
and U992 (N_992,In_321,In_356);
nand U993 (N_993,In_134,In_126);
and U994 (N_994,In_237,In_586);
or U995 (N_995,In_427,In_358);
and U996 (N_996,In_21,In_680);
or U997 (N_997,In_204,In_161);
or U998 (N_998,In_424,In_529);
nor U999 (N_999,In_418,In_356);
or U1000 (N_1000,N_639,N_385);
nor U1001 (N_1001,N_590,N_403);
and U1002 (N_1002,N_553,N_116);
nand U1003 (N_1003,N_79,N_462);
or U1004 (N_1004,N_367,N_978);
or U1005 (N_1005,N_620,N_531);
nor U1006 (N_1006,N_255,N_148);
nor U1007 (N_1007,N_933,N_643);
or U1008 (N_1008,N_88,N_538);
nor U1009 (N_1009,N_912,N_262);
and U1010 (N_1010,N_320,N_684);
and U1011 (N_1011,N_640,N_986);
nor U1012 (N_1012,N_631,N_4);
nand U1013 (N_1013,N_888,N_916);
and U1014 (N_1014,N_605,N_525);
or U1015 (N_1015,N_419,N_586);
nand U1016 (N_1016,N_519,N_170);
nor U1017 (N_1017,N_993,N_144);
and U1018 (N_1018,N_834,N_547);
nor U1019 (N_1019,N_168,N_726);
nor U1020 (N_1020,N_511,N_288);
and U1021 (N_1021,N_767,N_956);
nand U1022 (N_1022,N_158,N_505);
and U1023 (N_1023,N_802,N_446);
and U1024 (N_1024,N_345,N_592);
nor U1025 (N_1025,N_370,N_105);
and U1026 (N_1026,N_881,N_534);
nor U1027 (N_1027,N_233,N_156);
and U1028 (N_1028,N_152,N_861);
nand U1029 (N_1029,N_698,N_151);
nand U1030 (N_1030,N_809,N_472);
and U1031 (N_1031,N_421,N_845);
or U1032 (N_1032,N_545,N_413);
nor U1033 (N_1033,N_527,N_215);
and U1034 (N_1034,N_139,N_234);
and U1035 (N_1035,N_975,N_38);
nand U1036 (N_1036,N_572,N_203);
nor U1037 (N_1037,N_702,N_235);
nand U1038 (N_1038,N_530,N_591);
nand U1039 (N_1039,N_826,N_409);
nor U1040 (N_1040,N_406,N_98);
and U1041 (N_1041,N_117,N_821);
or U1042 (N_1042,N_179,N_688);
or U1043 (N_1043,N_659,N_430);
and U1044 (N_1044,N_914,N_416);
xnor U1045 (N_1045,N_106,N_838);
nand U1046 (N_1046,N_456,N_227);
nor U1047 (N_1047,N_955,N_837);
and U1048 (N_1048,N_526,N_165);
or U1049 (N_1049,N_181,N_954);
or U1050 (N_1050,N_128,N_334);
nand U1051 (N_1051,N_318,N_997);
or U1052 (N_1052,N_849,N_138);
or U1053 (N_1053,N_540,N_625);
or U1054 (N_1054,N_339,N_45);
nand U1055 (N_1055,N_867,N_395);
nand U1056 (N_1056,N_972,N_201);
or U1057 (N_1057,N_321,N_942);
nor U1058 (N_1058,N_304,N_322);
and U1059 (N_1059,N_95,N_828);
nor U1060 (N_1060,N_418,N_184);
or U1061 (N_1061,N_177,N_564);
and U1062 (N_1062,N_758,N_120);
nand U1063 (N_1063,N_11,N_581);
or U1064 (N_1064,N_500,N_617);
or U1065 (N_1065,N_477,N_878);
nor U1066 (N_1066,N_559,N_715);
nand U1067 (N_1067,N_343,N_58);
and U1068 (N_1068,N_424,N_964);
and U1069 (N_1069,N_209,N_101);
nand U1070 (N_1070,N_31,N_238);
nor U1071 (N_1071,N_818,N_727);
or U1072 (N_1072,N_792,N_579);
nand U1073 (N_1073,N_630,N_550);
nand U1074 (N_1074,N_543,N_357);
nor U1075 (N_1075,N_609,N_600);
xnor U1076 (N_1076,N_587,N_100);
and U1077 (N_1077,N_348,N_663);
nand U1078 (N_1078,N_967,N_768);
nand U1079 (N_1079,N_438,N_860);
nand U1080 (N_1080,N_672,N_257);
xor U1081 (N_1081,N_417,N_976);
or U1082 (N_1082,N_515,N_467);
and U1083 (N_1083,N_848,N_296);
nand U1084 (N_1084,N_903,N_72);
or U1085 (N_1085,N_880,N_984);
nand U1086 (N_1086,N_371,N_730);
nor U1087 (N_1087,N_567,N_295);
and U1088 (N_1088,N_466,N_958);
nand U1089 (N_1089,N_745,N_84);
or U1090 (N_1090,N_896,N_610);
or U1091 (N_1091,N_133,N_415);
and U1092 (N_1092,N_405,N_940);
nor U1093 (N_1093,N_351,N_977);
nor U1094 (N_1094,N_762,N_655);
xor U1095 (N_1095,N_223,N_317);
nor U1096 (N_1096,N_966,N_678);
and U1097 (N_1097,N_825,N_626);
nand U1098 (N_1098,N_734,N_426);
or U1099 (N_1099,N_907,N_407);
or U1100 (N_1100,N_573,N_269);
nor U1101 (N_1101,N_192,N_352);
or U1102 (N_1102,N_25,N_769);
and U1103 (N_1103,N_687,N_171);
nor U1104 (N_1104,N_300,N_504);
nand U1105 (N_1105,N_356,N_603);
nand U1106 (N_1106,N_798,N_231);
and U1107 (N_1107,N_16,N_857);
or U1108 (N_1108,N_358,N_824);
and U1109 (N_1109,N_278,N_259);
and U1110 (N_1110,N_281,N_206);
nand U1111 (N_1111,N_930,N_202);
nand U1112 (N_1112,N_902,N_570);
nand U1113 (N_1113,N_740,N_246);
nor U1114 (N_1114,N_196,N_488);
nor U1115 (N_1115,N_782,N_542);
or U1116 (N_1116,N_623,N_283);
nor U1117 (N_1117,N_576,N_991);
and U1118 (N_1118,N_854,N_80);
nor U1119 (N_1119,N_636,N_693);
and U1120 (N_1120,N_868,N_360);
or U1121 (N_1121,N_719,N_90);
nand U1122 (N_1122,N_331,N_219);
and U1123 (N_1123,N_529,N_256);
nor U1124 (N_1124,N_344,N_752);
and U1125 (N_1125,N_901,N_199);
or U1126 (N_1126,N_115,N_354);
nand U1127 (N_1127,N_724,N_260);
nand U1128 (N_1128,N_862,N_756);
nand U1129 (N_1129,N_285,N_738);
or U1130 (N_1130,N_694,N_746);
or U1131 (N_1131,N_588,N_381);
or U1132 (N_1132,N_19,N_271);
nand U1133 (N_1133,N_392,N_582);
nand U1134 (N_1134,N_615,N_654);
and U1135 (N_1135,N_622,N_827);
nor U1136 (N_1136,N_760,N_859);
nand U1137 (N_1137,N_26,N_3);
nor U1138 (N_1138,N_677,N_102);
nand U1139 (N_1139,N_53,N_784);
nor U1140 (N_1140,N_535,N_665);
nand U1141 (N_1141,N_708,N_70);
or U1142 (N_1142,N_228,N_764);
or U1143 (N_1143,N_198,N_110);
and U1144 (N_1144,N_469,N_502);
nand U1145 (N_1145,N_949,N_298);
and U1146 (N_1146,N_983,N_404);
and U1147 (N_1147,N_720,N_8);
and U1148 (N_1148,N_939,N_495);
nor U1149 (N_1149,N_447,N_330);
nand U1150 (N_1150,N_783,N_22);
or U1151 (N_1151,N_69,N_910);
nor U1152 (N_1152,N_869,N_309);
nor U1153 (N_1153,N_660,N_412);
nor U1154 (N_1154,N_887,N_64);
or U1155 (N_1155,N_44,N_160);
nand U1156 (N_1156,N_114,N_539);
or U1157 (N_1157,N_803,N_291);
and U1158 (N_1158,N_815,N_870);
and U1159 (N_1159,N_420,N_479);
and U1160 (N_1160,N_568,N_324);
nand U1161 (N_1161,N_701,N_274);
and U1162 (N_1162,N_154,N_489);
or U1163 (N_1163,N_290,N_453);
and U1164 (N_1164,N_583,N_213);
nand U1165 (N_1165,N_150,N_627);
and U1166 (N_1166,N_61,N_136);
nor U1167 (N_1167,N_207,N_422);
or U1168 (N_1168,N_959,N_458);
nor U1169 (N_1169,N_432,N_463);
nand U1170 (N_1170,N_561,N_808);
or U1171 (N_1171,N_645,N_578);
and U1172 (N_1172,N_516,N_445);
nand U1173 (N_1173,N_178,N_175);
and U1174 (N_1174,N_995,N_691);
nand U1175 (N_1175,N_63,N_261);
nand U1176 (N_1176,N_323,N_491);
xnor U1177 (N_1177,N_624,N_107);
nor U1178 (N_1178,N_990,N_800);
nand U1179 (N_1179,N_315,N_155);
or U1180 (N_1180,N_641,N_565);
and U1181 (N_1181,N_493,N_707);
nor U1182 (N_1182,N_840,N_874);
nor U1183 (N_1183,N_476,N_980);
nand U1184 (N_1184,N_240,N_554);
and U1185 (N_1185,N_595,N_786);
nor U1186 (N_1186,N_87,N_86);
and U1187 (N_1187,N_552,N_364);
nor U1188 (N_1188,N_311,N_931);
nor U1189 (N_1189,N_601,N_706);
or U1190 (N_1190,N_183,N_490);
or U1191 (N_1191,N_936,N_960);
and U1192 (N_1192,N_425,N_174);
and U1193 (N_1193,N_440,N_112);
nand U1194 (N_1194,N_369,N_245);
nand U1195 (N_1195,N_969,N_580);
and U1196 (N_1196,N_408,N_856);
or U1197 (N_1197,N_810,N_366);
and U1198 (N_1198,N_905,N_731);
xnor U1199 (N_1199,N_666,N_17);
nand U1200 (N_1200,N_506,N_119);
nor U1201 (N_1201,N_676,N_523);
nor U1202 (N_1202,N_652,N_51);
nor U1203 (N_1203,N_289,N_944);
nor U1204 (N_1204,N_62,N_671);
nand U1205 (N_1205,N_632,N_108);
nand U1206 (N_1206,N_81,N_236);
or U1207 (N_1207,N_305,N_602);
nor U1208 (N_1208,N_968,N_725);
xor U1209 (N_1209,N_226,N_427);
or U1210 (N_1210,N_680,N_876);
or U1211 (N_1211,N_29,N_950);
nor U1212 (N_1212,N_402,N_889);
nor U1213 (N_1213,N_929,N_471);
nor U1214 (N_1214,N_225,N_464);
nand U1215 (N_1215,N_389,N_753);
or U1216 (N_1216,N_925,N_575);
and U1217 (N_1217,N_723,N_563);
nor U1218 (N_1218,N_548,N_208);
nor U1219 (N_1219,N_536,N_190);
nand U1220 (N_1220,N_21,N_341);
or U1221 (N_1221,N_858,N_66);
and U1222 (N_1222,N_75,N_250);
or U1223 (N_1223,N_822,N_879);
and U1224 (N_1224,N_714,N_717);
or U1225 (N_1225,N_829,N_13);
and U1226 (N_1226,N_328,N_894);
nand U1227 (N_1227,N_584,N_937);
nor U1228 (N_1228,N_599,N_695);
or U1229 (N_1229,N_39,N_164);
and U1230 (N_1230,N_656,N_794);
nand U1231 (N_1231,N_308,N_613);
nor U1232 (N_1232,N_514,N_47);
nand U1233 (N_1233,N_316,N_804);
and U1234 (N_1234,N_770,N_674);
nand U1235 (N_1235,N_823,N_393);
or U1236 (N_1236,N_465,N_350);
or U1237 (N_1237,N_906,N_167);
or U1238 (N_1238,N_843,N_711);
nand U1239 (N_1239,N_985,N_94);
and U1240 (N_1240,N_650,N_23);
nor U1241 (N_1241,N_375,N_598);
nand U1242 (N_1242,N_355,N_710);
nor U1243 (N_1243,N_728,N_833);
and U1244 (N_1244,N_310,N_338);
or U1245 (N_1245,N_91,N_952);
and U1246 (N_1246,N_113,N_638);
nor U1247 (N_1247,N_65,N_55);
or U1248 (N_1248,N_562,N_934);
and U1249 (N_1249,N_195,N_361);
nand U1250 (N_1250,N_492,N_157);
nor U1251 (N_1251,N_411,N_394);
nand U1252 (N_1252,N_461,N_14);
or U1253 (N_1253,N_629,N_470);
or U1254 (N_1254,N_410,N_242);
nor U1255 (N_1255,N_36,N_992);
or U1256 (N_1256,N_455,N_239);
or U1257 (N_1257,N_847,N_382);
nand U1258 (N_1258,N_751,N_301);
and U1259 (N_1259,N_961,N_191);
and U1260 (N_1260,N_846,N_460);
or U1261 (N_1261,N_533,N_941);
or U1262 (N_1262,N_104,N_919);
nor U1263 (N_1263,N_123,N_923);
xor U1264 (N_1264,N_841,N_947);
and U1265 (N_1265,N_89,N_737);
and U1266 (N_1266,N_335,N_507);
nor U1267 (N_1267,N_78,N_92);
nand U1268 (N_1268,N_836,N_673);
nor U1269 (N_1269,N_265,N_48);
xnor U1270 (N_1270,N_789,N_482);
nand U1271 (N_1271,N_313,N_169);
nand U1272 (N_1272,N_635,N_204);
nor U1273 (N_1273,N_377,N_200);
nand U1274 (N_1274,N_773,N_795);
and U1275 (N_1275,N_428,N_544);
or U1276 (N_1276,N_142,N_485);
nand U1277 (N_1277,N_979,N_275);
and U1278 (N_1278,N_917,N_454);
and U1279 (N_1279,N_380,N_899);
and U1280 (N_1280,N_302,N_686);
or U1281 (N_1281,N_153,N_132);
or U1282 (N_1282,N_494,N_400);
nor U1283 (N_1283,N_264,N_263);
and U1284 (N_1284,N_434,N_628);
and U1285 (N_1285,N_657,N_210);
or U1286 (N_1286,N_327,N_67);
nor U1287 (N_1287,N_807,N_34);
nor U1288 (N_1288,N_744,N_337);
nand U1289 (N_1289,N_963,N_46);
xnor U1290 (N_1290,N_741,N_131);
and U1291 (N_1291,N_759,N_254);
xor U1292 (N_1292,N_188,N_682);
nand U1293 (N_1293,N_253,N_386);
nor U1294 (N_1294,N_436,N_697);
and U1295 (N_1295,N_475,N_662);
and U1296 (N_1296,N_222,N_816);
and U1297 (N_1297,N_957,N_921);
nand U1298 (N_1298,N_211,N_266);
nor U1299 (N_1299,N_653,N_374);
and U1300 (N_1300,N_314,N_831);
nor U1301 (N_1301,N_59,N_124);
nand U1302 (N_1302,N_998,N_484);
nand U1303 (N_1303,N_669,N_333);
nor U1304 (N_1304,N_99,N_607);
xnor U1305 (N_1305,N_904,N_109);
or U1306 (N_1306,N_537,N_596);
or U1307 (N_1307,N_483,N_276);
or U1308 (N_1308,N_383,N_9);
or U1309 (N_1309,N_193,N_999);
nand U1310 (N_1310,N_251,N_121);
xor U1311 (N_1311,N_258,N_541);
nor U1312 (N_1312,N_284,N_560);
or U1313 (N_1313,N_633,N_137);
nand U1314 (N_1314,N_487,N_739);
or U1315 (N_1315,N_372,N_486);
or U1316 (N_1316,N_546,N_781);
nand U1317 (N_1317,N_911,N_449);
nor U1318 (N_1318,N_785,N_973);
or U1319 (N_1319,N_329,N_437);
and U1320 (N_1320,N_733,N_229);
nor U1321 (N_1321,N_765,N_649);
or U1322 (N_1322,N_700,N_619);
and U1323 (N_1323,N_474,N_243);
nand U1324 (N_1324,N_7,N_468);
and U1325 (N_1325,N_43,N_683);
and U1326 (N_1326,N_791,N_556);
and U1327 (N_1327,N_608,N_30);
nand U1328 (N_1328,N_448,N_989);
or U1329 (N_1329,N_140,N_129);
and U1330 (N_1330,N_704,N_521);
nand U1331 (N_1331,N_853,N_926);
and U1332 (N_1332,N_42,N_644);
or U1333 (N_1333,N_480,N_951);
and U1334 (N_1334,N_604,N_766);
nor U1335 (N_1335,N_528,N_145);
and U1336 (N_1336,N_52,N_776);
and U1337 (N_1337,N_216,N_557);
nor U1338 (N_1338,N_864,N_166);
and U1339 (N_1339,N_220,N_268);
and U1340 (N_1340,N_722,N_365);
or U1341 (N_1341,N_35,N_850);
nor U1342 (N_1342,N_811,N_873);
nor U1343 (N_1343,N_244,N_287);
and U1344 (N_1344,N_713,N_812);
nor U1345 (N_1345,N_924,N_267);
or U1346 (N_1346,N_496,N_813);
and U1347 (N_1347,N_24,N_230);
nand U1348 (N_1348,N_378,N_801);
nor U1349 (N_1349,N_247,N_908);
or U1350 (N_1350,N_56,N_353);
and U1351 (N_1351,N_597,N_761);
nand U1352 (N_1352,N_326,N_935);
or U1353 (N_1353,N_249,N_306);
and U1354 (N_1354,N_790,N_664);
and U1355 (N_1355,N_60,N_194);
nand U1356 (N_1356,N_126,N_187);
and U1357 (N_1357,N_186,N_146);
nor U1358 (N_1358,N_270,N_135);
and U1359 (N_1359,N_749,N_909);
nand U1360 (N_1360,N_918,N_368);
nor U1361 (N_1361,N_349,N_397);
nand U1362 (N_1362,N_443,N_915);
xnor U1363 (N_1363,N_252,N_705);
nand U1364 (N_1364,N_670,N_224);
or U1365 (N_1365,N_149,N_763);
nand U1366 (N_1366,N_212,N_551);
or U1367 (N_1367,N_780,N_805);
or U1368 (N_1368,N_162,N_787);
and U1369 (N_1369,N_574,N_441);
and U1370 (N_1370,N_297,N_646);
xnor U1371 (N_1371,N_172,N_180);
or U1372 (N_1372,N_913,N_532);
nand U1373 (N_1373,N_71,N_359);
or U1374 (N_1374,N_793,N_32);
and U1375 (N_1375,N_689,N_748);
and U1376 (N_1376,N_130,N_839);
xnor U1377 (N_1377,N_57,N_750);
nor U1378 (N_1378,N_387,N_721);
xnor U1379 (N_1379,N_775,N_76);
nand U1380 (N_1380,N_49,N_920);
nor U1381 (N_1381,N_185,N_895);
nor U1382 (N_1382,N_159,N_272);
nor U1383 (N_1383,N_651,N_696);
and U1384 (N_1384,N_457,N_621);
nand U1385 (N_1385,N_147,N_863);
or U1386 (N_1386,N_981,N_882);
nand U1387 (N_1387,N_886,N_221);
and U1388 (N_1388,N_517,N_732);
or U1389 (N_1389,N_451,N_675);
nor U1390 (N_1390,N_510,N_143);
and U1391 (N_1391,N_423,N_161);
and U1392 (N_1392,N_974,N_742);
or U1393 (N_1393,N_277,N_616);
or U1394 (N_1394,N_612,N_373);
or U1395 (N_1395,N_830,N_499);
or U1396 (N_1396,N_593,N_232);
or U1397 (N_1397,N_82,N_928);
nand U1398 (N_1398,N_141,N_668);
and U1399 (N_1399,N_379,N_932);
and U1400 (N_1400,N_54,N_294);
and U1401 (N_1401,N_340,N_844);
nor U1402 (N_1402,N_391,N_452);
and U1403 (N_1403,N_173,N_15);
nand U1404 (N_1404,N_299,N_96);
nor U1405 (N_1405,N_943,N_197);
or U1406 (N_1406,N_50,N_218);
and U1407 (N_1407,N_661,N_280);
or U1408 (N_1408,N_852,N_512);
and U1409 (N_1409,N_814,N_777);
or U1410 (N_1410,N_842,N_703);
nor U1411 (N_1411,N_658,N_685);
or U1412 (N_1412,N_134,N_97);
nor U1413 (N_1413,N_513,N_214);
nor U1414 (N_1414,N_994,N_241);
nand U1415 (N_1415,N_396,N_37);
nor U1416 (N_1416,N_509,N_735);
or U1417 (N_1417,N_524,N_729);
and U1418 (N_1418,N_819,N_778);
nor U1419 (N_1419,N_127,N_248);
nand U1420 (N_1420,N_293,N_388);
nand U1421 (N_1421,N_459,N_716);
nand U1422 (N_1422,N_571,N_40);
and U1423 (N_1423,N_346,N_384);
or U1424 (N_1424,N_312,N_577);
or U1425 (N_1425,N_5,N_871);
nand U1426 (N_1426,N_755,N_362);
nand U1427 (N_1427,N_401,N_41);
nor U1428 (N_1428,N_893,N_501);
nand U1429 (N_1429,N_788,N_982);
nand U1430 (N_1430,N_1,N_875);
nand U1431 (N_1431,N_962,N_6);
and U1432 (N_1432,N_347,N_892);
and U1433 (N_1433,N_111,N_431);
nor U1434 (N_1434,N_712,N_319);
nand U1435 (N_1435,N_74,N_439);
xnor U1436 (N_1436,N_614,N_332);
nor U1437 (N_1437,N_897,N_429);
or U1438 (N_1438,N_855,N_518);
nor U1439 (N_1439,N_0,N_872);
or U1440 (N_1440,N_779,N_163);
and U1441 (N_1441,N_865,N_2);
nand U1442 (N_1442,N_189,N_558);
nor U1443 (N_1443,N_988,N_28);
and U1444 (N_1444,N_566,N_747);
or U1445 (N_1445,N_637,N_286);
or U1446 (N_1446,N_948,N_503);
or U1447 (N_1447,N_435,N_376);
and U1448 (N_1448,N_699,N_648);
or U1449 (N_1449,N_444,N_877);
nor U1450 (N_1450,N_709,N_594);
or U1451 (N_1451,N_679,N_292);
nor U1452 (N_1452,N_799,N_965);
or U1453 (N_1453,N_103,N_611);
nor U1454 (N_1454,N_692,N_890);
nand U1455 (N_1455,N_806,N_473);
nor U1456 (N_1456,N_498,N_93);
or U1457 (N_1457,N_606,N_549);
or U1458 (N_1458,N_336,N_27);
or U1459 (N_1459,N_497,N_690);
and U1460 (N_1460,N_851,N_885);
nor U1461 (N_1461,N_796,N_883);
or U1462 (N_1462,N_884,N_10);
nand U1463 (N_1463,N_273,N_927);
or U1464 (N_1464,N_971,N_898);
or U1465 (N_1465,N_953,N_478);
and U1466 (N_1466,N_938,N_774);
and U1467 (N_1467,N_832,N_736);
nor U1468 (N_1468,N_866,N_398);
nand U1469 (N_1469,N_891,N_520);
nand U1470 (N_1470,N_771,N_20);
or U1471 (N_1471,N_176,N_797);
and U1472 (N_1472,N_772,N_945);
nand U1473 (N_1473,N_325,N_33);
or U1474 (N_1474,N_522,N_743);
nor U1475 (N_1475,N_122,N_118);
nand U1476 (N_1476,N_481,N_757);
nand U1477 (N_1477,N_681,N_73);
nor U1478 (N_1478,N_237,N_282);
or U1479 (N_1479,N_634,N_508);
nor U1480 (N_1480,N_922,N_642);
nand U1481 (N_1481,N_946,N_205);
xnor U1482 (N_1482,N_835,N_399);
or U1483 (N_1483,N_18,N_85);
nor U1484 (N_1484,N_279,N_125);
nor U1485 (N_1485,N_987,N_647);
nor U1486 (N_1486,N_618,N_900);
nand U1487 (N_1487,N_363,N_718);
or U1488 (N_1488,N_585,N_77);
nor U1489 (N_1489,N_433,N_182);
nor U1490 (N_1490,N_390,N_442);
and U1491 (N_1491,N_996,N_12);
or U1492 (N_1492,N_569,N_83);
or U1493 (N_1493,N_555,N_817);
or U1494 (N_1494,N_303,N_667);
xnor U1495 (N_1495,N_342,N_68);
and U1496 (N_1496,N_414,N_307);
or U1497 (N_1497,N_820,N_217);
and U1498 (N_1498,N_754,N_450);
nand U1499 (N_1499,N_970,N_589);
or U1500 (N_1500,N_644,N_445);
nand U1501 (N_1501,N_676,N_754);
and U1502 (N_1502,N_513,N_979);
nand U1503 (N_1503,N_210,N_494);
nor U1504 (N_1504,N_451,N_46);
or U1505 (N_1505,N_620,N_934);
nor U1506 (N_1506,N_452,N_107);
nor U1507 (N_1507,N_446,N_189);
nor U1508 (N_1508,N_705,N_723);
and U1509 (N_1509,N_842,N_848);
or U1510 (N_1510,N_955,N_142);
or U1511 (N_1511,N_71,N_307);
and U1512 (N_1512,N_302,N_877);
nor U1513 (N_1513,N_847,N_849);
nand U1514 (N_1514,N_271,N_816);
xnor U1515 (N_1515,N_541,N_925);
or U1516 (N_1516,N_469,N_570);
nand U1517 (N_1517,N_255,N_714);
or U1518 (N_1518,N_849,N_881);
nor U1519 (N_1519,N_526,N_300);
nand U1520 (N_1520,N_533,N_66);
nand U1521 (N_1521,N_509,N_385);
nand U1522 (N_1522,N_780,N_599);
or U1523 (N_1523,N_396,N_554);
or U1524 (N_1524,N_991,N_618);
or U1525 (N_1525,N_450,N_676);
nor U1526 (N_1526,N_321,N_207);
nand U1527 (N_1527,N_783,N_46);
nand U1528 (N_1528,N_83,N_300);
or U1529 (N_1529,N_968,N_400);
nand U1530 (N_1530,N_758,N_882);
nor U1531 (N_1531,N_277,N_739);
nand U1532 (N_1532,N_841,N_372);
nand U1533 (N_1533,N_284,N_409);
nor U1534 (N_1534,N_543,N_215);
and U1535 (N_1535,N_919,N_807);
nor U1536 (N_1536,N_288,N_135);
or U1537 (N_1537,N_165,N_427);
or U1538 (N_1538,N_922,N_541);
or U1539 (N_1539,N_678,N_756);
or U1540 (N_1540,N_700,N_570);
and U1541 (N_1541,N_768,N_222);
and U1542 (N_1542,N_577,N_553);
or U1543 (N_1543,N_68,N_24);
nor U1544 (N_1544,N_279,N_747);
nor U1545 (N_1545,N_996,N_907);
and U1546 (N_1546,N_512,N_984);
xor U1547 (N_1547,N_594,N_168);
nand U1548 (N_1548,N_610,N_432);
nor U1549 (N_1549,N_303,N_480);
nand U1550 (N_1550,N_926,N_78);
nor U1551 (N_1551,N_721,N_723);
nor U1552 (N_1552,N_737,N_46);
nor U1553 (N_1553,N_575,N_485);
or U1554 (N_1554,N_447,N_246);
nand U1555 (N_1555,N_429,N_397);
and U1556 (N_1556,N_799,N_6);
nor U1557 (N_1557,N_393,N_477);
xnor U1558 (N_1558,N_3,N_570);
or U1559 (N_1559,N_949,N_700);
nand U1560 (N_1560,N_30,N_733);
nor U1561 (N_1561,N_985,N_532);
or U1562 (N_1562,N_762,N_37);
nor U1563 (N_1563,N_398,N_990);
or U1564 (N_1564,N_658,N_926);
or U1565 (N_1565,N_260,N_42);
nand U1566 (N_1566,N_764,N_22);
nand U1567 (N_1567,N_820,N_390);
nor U1568 (N_1568,N_729,N_293);
or U1569 (N_1569,N_807,N_295);
and U1570 (N_1570,N_593,N_800);
nand U1571 (N_1571,N_203,N_876);
or U1572 (N_1572,N_586,N_817);
nor U1573 (N_1573,N_903,N_703);
nor U1574 (N_1574,N_422,N_967);
nor U1575 (N_1575,N_131,N_829);
nand U1576 (N_1576,N_442,N_508);
or U1577 (N_1577,N_514,N_979);
nand U1578 (N_1578,N_142,N_437);
nand U1579 (N_1579,N_119,N_533);
nand U1580 (N_1580,N_650,N_856);
or U1581 (N_1581,N_30,N_232);
nand U1582 (N_1582,N_860,N_909);
or U1583 (N_1583,N_10,N_982);
xor U1584 (N_1584,N_161,N_441);
and U1585 (N_1585,N_974,N_409);
and U1586 (N_1586,N_257,N_569);
nand U1587 (N_1587,N_345,N_529);
or U1588 (N_1588,N_145,N_938);
nand U1589 (N_1589,N_954,N_475);
or U1590 (N_1590,N_120,N_239);
nor U1591 (N_1591,N_475,N_717);
or U1592 (N_1592,N_21,N_265);
nor U1593 (N_1593,N_203,N_635);
nor U1594 (N_1594,N_549,N_837);
or U1595 (N_1595,N_456,N_714);
nand U1596 (N_1596,N_878,N_115);
or U1597 (N_1597,N_708,N_849);
nand U1598 (N_1598,N_186,N_409);
or U1599 (N_1599,N_69,N_572);
or U1600 (N_1600,N_328,N_110);
nor U1601 (N_1601,N_790,N_237);
nor U1602 (N_1602,N_335,N_431);
nor U1603 (N_1603,N_366,N_945);
and U1604 (N_1604,N_12,N_566);
nor U1605 (N_1605,N_54,N_956);
nand U1606 (N_1606,N_114,N_647);
nor U1607 (N_1607,N_738,N_392);
or U1608 (N_1608,N_234,N_955);
nand U1609 (N_1609,N_945,N_993);
and U1610 (N_1610,N_162,N_295);
nor U1611 (N_1611,N_227,N_325);
nand U1612 (N_1612,N_267,N_542);
nand U1613 (N_1613,N_900,N_305);
and U1614 (N_1614,N_777,N_246);
or U1615 (N_1615,N_860,N_895);
nor U1616 (N_1616,N_968,N_513);
nor U1617 (N_1617,N_26,N_803);
or U1618 (N_1618,N_34,N_376);
nor U1619 (N_1619,N_731,N_503);
or U1620 (N_1620,N_376,N_407);
and U1621 (N_1621,N_771,N_886);
or U1622 (N_1622,N_212,N_162);
nor U1623 (N_1623,N_673,N_776);
or U1624 (N_1624,N_439,N_233);
and U1625 (N_1625,N_821,N_481);
or U1626 (N_1626,N_149,N_941);
and U1627 (N_1627,N_727,N_35);
or U1628 (N_1628,N_271,N_877);
nand U1629 (N_1629,N_596,N_82);
nand U1630 (N_1630,N_705,N_954);
nand U1631 (N_1631,N_565,N_295);
and U1632 (N_1632,N_858,N_277);
nor U1633 (N_1633,N_802,N_63);
and U1634 (N_1634,N_244,N_679);
xor U1635 (N_1635,N_511,N_226);
and U1636 (N_1636,N_792,N_765);
and U1637 (N_1637,N_682,N_831);
nor U1638 (N_1638,N_221,N_364);
or U1639 (N_1639,N_822,N_46);
nor U1640 (N_1640,N_943,N_865);
or U1641 (N_1641,N_660,N_969);
and U1642 (N_1642,N_614,N_240);
nand U1643 (N_1643,N_335,N_865);
nor U1644 (N_1644,N_305,N_213);
nand U1645 (N_1645,N_45,N_180);
or U1646 (N_1646,N_95,N_981);
nand U1647 (N_1647,N_784,N_72);
and U1648 (N_1648,N_159,N_115);
or U1649 (N_1649,N_453,N_689);
nor U1650 (N_1650,N_414,N_270);
nand U1651 (N_1651,N_172,N_535);
nand U1652 (N_1652,N_712,N_809);
or U1653 (N_1653,N_18,N_716);
and U1654 (N_1654,N_997,N_575);
nand U1655 (N_1655,N_247,N_404);
nor U1656 (N_1656,N_31,N_235);
and U1657 (N_1657,N_88,N_398);
nand U1658 (N_1658,N_111,N_469);
nor U1659 (N_1659,N_403,N_692);
and U1660 (N_1660,N_923,N_275);
xor U1661 (N_1661,N_545,N_55);
nand U1662 (N_1662,N_21,N_852);
nand U1663 (N_1663,N_506,N_557);
nand U1664 (N_1664,N_386,N_144);
or U1665 (N_1665,N_691,N_402);
nor U1666 (N_1666,N_333,N_211);
nand U1667 (N_1667,N_961,N_846);
xnor U1668 (N_1668,N_348,N_417);
or U1669 (N_1669,N_429,N_423);
nand U1670 (N_1670,N_839,N_227);
nand U1671 (N_1671,N_727,N_303);
nand U1672 (N_1672,N_34,N_806);
or U1673 (N_1673,N_491,N_67);
xnor U1674 (N_1674,N_108,N_419);
nand U1675 (N_1675,N_622,N_598);
nand U1676 (N_1676,N_571,N_724);
and U1677 (N_1677,N_903,N_847);
nor U1678 (N_1678,N_345,N_322);
nor U1679 (N_1679,N_759,N_118);
nor U1680 (N_1680,N_792,N_538);
nand U1681 (N_1681,N_631,N_746);
or U1682 (N_1682,N_34,N_613);
or U1683 (N_1683,N_435,N_17);
or U1684 (N_1684,N_396,N_864);
nand U1685 (N_1685,N_132,N_480);
and U1686 (N_1686,N_152,N_965);
nand U1687 (N_1687,N_361,N_261);
or U1688 (N_1688,N_345,N_765);
nand U1689 (N_1689,N_410,N_916);
nor U1690 (N_1690,N_898,N_279);
nand U1691 (N_1691,N_579,N_249);
nand U1692 (N_1692,N_296,N_953);
or U1693 (N_1693,N_203,N_438);
nand U1694 (N_1694,N_315,N_152);
or U1695 (N_1695,N_144,N_952);
and U1696 (N_1696,N_471,N_720);
and U1697 (N_1697,N_19,N_252);
or U1698 (N_1698,N_420,N_145);
and U1699 (N_1699,N_823,N_688);
nor U1700 (N_1700,N_278,N_65);
or U1701 (N_1701,N_782,N_491);
nor U1702 (N_1702,N_543,N_725);
and U1703 (N_1703,N_900,N_487);
or U1704 (N_1704,N_117,N_491);
nor U1705 (N_1705,N_194,N_552);
or U1706 (N_1706,N_440,N_992);
nor U1707 (N_1707,N_524,N_585);
and U1708 (N_1708,N_422,N_116);
nor U1709 (N_1709,N_366,N_343);
nor U1710 (N_1710,N_772,N_394);
or U1711 (N_1711,N_330,N_362);
nor U1712 (N_1712,N_62,N_525);
or U1713 (N_1713,N_407,N_938);
or U1714 (N_1714,N_954,N_684);
nor U1715 (N_1715,N_667,N_813);
nor U1716 (N_1716,N_897,N_525);
nor U1717 (N_1717,N_501,N_610);
nand U1718 (N_1718,N_781,N_51);
and U1719 (N_1719,N_904,N_524);
nand U1720 (N_1720,N_903,N_393);
nand U1721 (N_1721,N_453,N_197);
and U1722 (N_1722,N_900,N_233);
or U1723 (N_1723,N_994,N_562);
and U1724 (N_1724,N_464,N_746);
nand U1725 (N_1725,N_247,N_29);
or U1726 (N_1726,N_492,N_763);
and U1727 (N_1727,N_982,N_380);
and U1728 (N_1728,N_265,N_544);
nand U1729 (N_1729,N_331,N_173);
nor U1730 (N_1730,N_187,N_956);
and U1731 (N_1731,N_452,N_292);
or U1732 (N_1732,N_89,N_206);
nand U1733 (N_1733,N_146,N_81);
and U1734 (N_1734,N_301,N_191);
nand U1735 (N_1735,N_489,N_147);
or U1736 (N_1736,N_124,N_480);
xor U1737 (N_1737,N_812,N_360);
xnor U1738 (N_1738,N_854,N_332);
nor U1739 (N_1739,N_831,N_733);
nor U1740 (N_1740,N_780,N_193);
or U1741 (N_1741,N_164,N_714);
and U1742 (N_1742,N_525,N_356);
and U1743 (N_1743,N_297,N_128);
nor U1744 (N_1744,N_741,N_826);
or U1745 (N_1745,N_379,N_938);
or U1746 (N_1746,N_243,N_911);
and U1747 (N_1747,N_732,N_946);
nand U1748 (N_1748,N_269,N_681);
and U1749 (N_1749,N_685,N_916);
and U1750 (N_1750,N_1,N_356);
or U1751 (N_1751,N_305,N_7);
or U1752 (N_1752,N_170,N_361);
or U1753 (N_1753,N_936,N_845);
or U1754 (N_1754,N_316,N_630);
or U1755 (N_1755,N_122,N_348);
nand U1756 (N_1756,N_599,N_749);
or U1757 (N_1757,N_542,N_393);
nand U1758 (N_1758,N_525,N_286);
nand U1759 (N_1759,N_332,N_924);
and U1760 (N_1760,N_738,N_881);
nor U1761 (N_1761,N_349,N_690);
nand U1762 (N_1762,N_193,N_213);
nor U1763 (N_1763,N_844,N_129);
nand U1764 (N_1764,N_421,N_738);
and U1765 (N_1765,N_158,N_471);
or U1766 (N_1766,N_343,N_800);
or U1767 (N_1767,N_64,N_227);
or U1768 (N_1768,N_146,N_769);
and U1769 (N_1769,N_768,N_322);
or U1770 (N_1770,N_267,N_303);
nor U1771 (N_1771,N_678,N_476);
nand U1772 (N_1772,N_881,N_45);
or U1773 (N_1773,N_549,N_839);
and U1774 (N_1774,N_545,N_530);
nor U1775 (N_1775,N_324,N_830);
nor U1776 (N_1776,N_495,N_736);
nand U1777 (N_1777,N_578,N_720);
nand U1778 (N_1778,N_116,N_42);
or U1779 (N_1779,N_870,N_714);
or U1780 (N_1780,N_399,N_596);
nand U1781 (N_1781,N_563,N_184);
nor U1782 (N_1782,N_30,N_751);
nor U1783 (N_1783,N_49,N_763);
or U1784 (N_1784,N_827,N_421);
nand U1785 (N_1785,N_871,N_135);
nor U1786 (N_1786,N_546,N_649);
nor U1787 (N_1787,N_503,N_332);
and U1788 (N_1788,N_622,N_902);
nor U1789 (N_1789,N_885,N_3);
xor U1790 (N_1790,N_391,N_831);
nor U1791 (N_1791,N_531,N_323);
or U1792 (N_1792,N_39,N_140);
and U1793 (N_1793,N_374,N_366);
nand U1794 (N_1794,N_536,N_906);
or U1795 (N_1795,N_943,N_789);
nor U1796 (N_1796,N_325,N_598);
or U1797 (N_1797,N_483,N_817);
nand U1798 (N_1798,N_873,N_105);
nor U1799 (N_1799,N_241,N_406);
and U1800 (N_1800,N_465,N_987);
or U1801 (N_1801,N_435,N_691);
and U1802 (N_1802,N_569,N_712);
nor U1803 (N_1803,N_377,N_66);
nand U1804 (N_1804,N_416,N_531);
nand U1805 (N_1805,N_135,N_271);
or U1806 (N_1806,N_695,N_613);
nand U1807 (N_1807,N_862,N_50);
or U1808 (N_1808,N_452,N_413);
nand U1809 (N_1809,N_315,N_428);
nor U1810 (N_1810,N_295,N_465);
nor U1811 (N_1811,N_352,N_685);
and U1812 (N_1812,N_181,N_492);
or U1813 (N_1813,N_766,N_441);
nor U1814 (N_1814,N_343,N_822);
nor U1815 (N_1815,N_470,N_217);
nor U1816 (N_1816,N_908,N_936);
nor U1817 (N_1817,N_755,N_669);
and U1818 (N_1818,N_987,N_548);
and U1819 (N_1819,N_796,N_84);
and U1820 (N_1820,N_882,N_268);
or U1821 (N_1821,N_589,N_526);
nor U1822 (N_1822,N_778,N_543);
nand U1823 (N_1823,N_34,N_98);
nor U1824 (N_1824,N_645,N_294);
nor U1825 (N_1825,N_945,N_499);
or U1826 (N_1826,N_178,N_177);
or U1827 (N_1827,N_865,N_784);
nor U1828 (N_1828,N_24,N_753);
nand U1829 (N_1829,N_57,N_378);
and U1830 (N_1830,N_58,N_175);
nor U1831 (N_1831,N_549,N_397);
and U1832 (N_1832,N_410,N_974);
nand U1833 (N_1833,N_814,N_45);
and U1834 (N_1834,N_899,N_630);
nand U1835 (N_1835,N_724,N_19);
or U1836 (N_1836,N_323,N_6);
nor U1837 (N_1837,N_296,N_847);
nor U1838 (N_1838,N_35,N_513);
or U1839 (N_1839,N_45,N_763);
nor U1840 (N_1840,N_126,N_260);
nor U1841 (N_1841,N_604,N_125);
or U1842 (N_1842,N_904,N_864);
nand U1843 (N_1843,N_195,N_689);
or U1844 (N_1844,N_174,N_923);
nand U1845 (N_1845,N_557,N_504);
or U1846 (N_1846,N_391,N_155);
or U1847 (N_1847,N_178,N_694);
and U1848 (N_1848,N_23,N_562);
nand U1849 (N_1849,N_725,N_775);
and U1850 (N_1850,N_29,N_910);
and U1851 (N_1851,N_321,N_734);
or U1852 (N_1852,N_734,N_216);
nand U1853 (N_1853,N_635,N_77);
and U1854 (N_1854,N_849,N_144);
and U1855 (N_1855,N_708,N_338);
and U1856 (N_1856,N_352,N_449);
nor U1857 (N_1857,N_721,N_121);
nand U1858 (N_1858,N_856,N_102);
and U1859 (N_1859,N_272,N_301);
nor U1860 (N_1860,N_409,N_95);
or U1861 (N_1861,N_558,N_643);
nor U1862 (N_1862,N_301,N_634);
nand U1863 (N_1863,N_369,N_886);
and U1864 (N_1864,N_961,N_134);
nand U1865 (N_1865,N_203,N_216);
xnor U1866 (N_1866,N_594,N_202);
and U1867 (N_1867,N_608,N_469);
and U1868 (N_1868,N_200,N_611);
and U1869 (N_1869,N_276,N_217);
nand U1870 (N_1870,N_482,N_639);
nand U1871 (N_1871,N_278,N_138);
or U1872 (N_1872,N_870,N_38);
and U1873 (N_1873,N_408,N_568);
and U1874 (N_1874,N_839,N_234);
nor U1875 (N_1875,N_556,N_513);
or U1876 (N_1876,N_363,N_76);
nand U1877 (N_1877,N_359,N_785);
nand U1878 (N_1878,N_123,N_10);
and U1879 (N_1879,N_843,N_271);
and U1880 (N_1880,N_70,N_48);
or U1881 (N_1881,N_763,N_762);
nor U1882 (N_1882,N_805,N_566);
nand U1883 (N_1883,N_36,N_172);
or U1884 (N_1884,N_62,N_570);
or U1885 (N_1885,N_208,N_678);
or U1886 (N_1886,N_753,N_693);
and U1887 (N_1887,N_68,N_854);
nor U1888 (N_1888,N_945,N_130);
and U1889 (N_1889,N_386,N_503);
nor U1890 (N_1890,N_489,N_536);
and U1891 (N_1891,N_240,N_959);
nor U1892 (N_1892,N_457,N_248);
xnor U1893 (N_1893,N_977,N_951);
nand U1894 (N_1894,N_758,N_365);
nand U1895 (N_1895,N_87,N_944);
or U1896 (N_1896,N_823,N_963);
nand U1897 (N_1897,N_447,N_577);
nor U1898 (N_1898,N_857,N_132);
and U1899 (N_1899,N_252,N_21);
nand U1900 (N_1900,N_73,N_308);
nand U1901 (N_1901,N_618,N_212);
or U1902 (N_1902,N_784,N_914);
xor U1903 (N_1903,N_256,N_945);
xnor U1904 (N_1904,N_803,N_597);
nand U1905 (N_1905,N_562,N_494);
nor U1906 (N_1906,N_275,N_985);
nand U1907 (N_1907,N_357,N_734);
or U1908 (N_1908,N_954,N_549);
and U1909 (N_1909,N_556,N_604);
xnor U1910 (N_1910,N_251,N_929);
nor U1911 (N_1911,N_845,N_218);
and U1912 (N_1912,N_23,N_288);
nor U1913 (N_1913,N_872,N_848);
or U1914 (N_1914,N_452,N_235);
and U1915 (N_1915,N_335,N_489);
nand U1916 (N_1916,N_722,N_3);
nand U1917 (N_1917,N_335,N_406);
and U1918 (N_1918,N_334,N_556);
nor U1919 (N_1919,N_996,N_351);
nor U1920 (N_1920,N_880,N_465);
nand U1921 (N_1921,N_561,N_494);
or U1922 (N_1922,N_251,N_828);
nand U1923 (N_1923,N_10,N_198);
and U1924 (N_1924,N_547,N_928);
nor U1925 (N_1925,N_415,N_278);
nand U1926 (N_1926,N_551,N_791);
nor U1927 (N_1927,N_170,N_110);
or U1928 (N_1928,N_811,N_179);
nor U1929 (N_1929,N_249,N_78);
or U1930 (N_1930,N_916,N_154);
nor U1931 (N_1931,N_139,N_964);
or U1932 (N_1932,N_91,N_204);
or U1933 (N_1933,N_54,N_422);
nand U1934 (N_1934,N_536,N_469);
nand U1935 (N_1935,N_582,N_34);
and U1936 (N_1936,N_461,N_897);
and U1937 (N_1937,N_237,N_773);
and U1938 (N_1938,N_704,N_73);
nor U1939 (N_1939,N_438,N_280);
nor U1940 (N_1940,N_559,N_822);
and U1941 (N_1941,N_628,N_682);
nor U1942 (N_1942,N_766,N_675);
nor U1943 (N_1943,N_502,N_68);
or U1944 (N_1944,N_354,N_92);
nor U1945 (N_1945,N_843,N_542);
nor U1946 (N_1946,N_547,N_557);
or U1947 (N_1947,N_909,N_102);
and U1948 (N_1948,N_927,N_697);
nand U1949 (N_1949,N_443,N_277);
nor U1950 (N_1950,N_947,N_665);
or U1951 (N_1951,N_161,N_984);
nand U1952 (N_1952,N_529,N_764);
or U1953 (N_1953,N_50,N_576);
nor U1954 (N_1954,N_933,N_245);
nand U1955 (N_1955,N_448,N_861);
or U1956 (N_1956,N_953,N_315);
nor U1957 (N_1957,N_923,N_789);
or U1958 (N_1958,N_479,N_827);
or U1959 (N_1959,N_691,N_892);
nor U1960 (N_1960,N_324,N_97);
or U1961 (N_1961,N_280,N_653);
nor U1962 (N_1962,N_489,N_852);
and U1963 (N_1963,N_115,N_813);
nor U1964 (N_1964,N_636,N_527);
and U1965 (N_1965,N_113,N_640);
nand U1966 (N_1966,N_89,N_773);
or U1967 (N_1967,N_578,N_867);
or U1968 (N_1968,N_401,N_777);
and U1969 (N_1969,N_239,N_14);
nand U1970 (N_1970,N_651,N_235);
nand U1971 (N_1971,N_901,N_950);
nor U1972 (N_1972,N_105,N_532);
and U1973 (N_1973,N_416,N_946);
or U1974 (N_1974,N_823,N_48);
and U1975 (N_1975,N_283,N_266);
or U1976 (N_1976,N_300,N_698);
nor U1977 (N_1977,N_855,N_596);
or U1978 (N_1978,N_500,N_515);
nor U1979 (N_1979,N_499,N_312);
and U1980 (N_1980,N_630,N_502);
or U1981 (N_1981,N_48,N_108);
nor U1982 (N_1982,N_867,N_383);
nor U1983 (N_1983,N_853,N_514);
nand U1984 (N_1984,N_624,N_564);
and U1985 (N_1985,N_298,N_227);
nand U1986 (N_1986,N_352,N_174);
and U1987 (N_1987,N_483,N_226);
or U1988 (N_1988,N_189,N_147);
nand U1989 (N_1989,N_33,N_457);
nor U1990 (N_1990,N_60,N_746);
nor U1991 (N_1991,N_35,N_688);
or U1992 (N_1992,N_538,N_784);
or U1993 (N_1993,N_943,N_303);
and U1994 (N_1994,N_691,N_663);
and U1995 (N_1995,N_454,N_317);
nand U1996 (N_1996,N_913,N_424);
xnor U1997 (N_1997,N_91,N_972);
nand U1998 (N_1998,N_333,N_851);
nand U1999 (N_1999,N_679,N_104);
or U2000 (N_2000,N_1051,N_1555);
nand U2001 (N_2001,N_1716,N_1312);
or U2002 (N_2002,N_1522,N_1521);
nor U2003 (N_2003,N_1730,N_1021);
nand U2004 (N_2004,N_1872,N_1643);
nand U2005 (N_2005,N_1819,N_1894);
nand U2006 (N_2006,N_1133,N_1975);
nand U2007 (N_2007,N_1771,N_1444);
nor U2008 (N_2008,N_1228,N_1766);
nor U2009 (N_2009,N_1205,N_1029);
nor U2010 (N_2010,N_1800,N_1639);
or U2011 (N_2011,N_1718,N_1092);
and U2012 (N_2012,N_1490,N_1709);
nor U2013 (N_2013,N_1638,N_1456);
and U2014 (N_2014,N_1600,N_1725);
nand U2015 (N_2015,N_1808,N_1791);
nor U2016 (N_2016,N_1708,N_1974);
or U2017 (N_2017,N_1246,N_1668);
xnor U2018 (N_2018,N_1991,N_1353);
nor U2019 (N_2019,N_1785,N_1626);
or U2020 (N_2020,N_1208,N_1996);
nor U2021 (N_2021,N_1673,N_1650);
nor U2022 (N_2022,N_1371,N_1473);
and U2023 (N_2023,N_1729,N_1278);
nor U2024 (N_2024,N_1889,N_1423);
and U2025 (N_2025,N_1903,N_1151);
nand U2026 (N_2026,N_1543,N_1796);
nor U2027 (N_2027,N_1284,N_1052);
or U2028 (N_2028,N_1439,N_1455);
nand U2029 (N_2029,N_1464,N_1534);
and U2030 (N_2030,N_1066,N_1292);
and U2031 (N_2031,N_1050,N_1012);
nand U2032 (N_2032,N_1416,N_1644);
nor U2033 (N_2033,N_1035,N_1765);
or U2034 (N_2034,N_1347,N_1632);
or U2035 (N_2035,N_1101,N_1424);
nand U2036 (N_2036,N_1811,N_1953);
and U2037 (N_2037,N_1307,N_1502);
nor U2038 (N_2038,N_1120,N_1817);
nor U2039 (N_2039,N_1893,N_1550);
nand U2040 (N_2040,N_1601,N_1302);
and U2041 (N_2041,N_1390,N_1666);
xnor U2042 (N_2042,N_1043,N_1062);
or U2043 (N_2043,N_1856,N_1488);
or U2044 (N_2044,N_1373,N_1255);
nand U2045 (N_2045,N_1123,N_1634);
nor U2046 (N_2046,N_1952,N_1535);
xor U2047 (N_2047,N_1265,N_1507);
nor U2048 (N_2048,N_1907,N_1395);
nor U2049 (N_2049,N_1485,N_1129);
and U2050 (N_2050,N_1486,N_1081);
nor U2051 (N_2051,N_1320,N_1781);
nand U2052 (N_2052,N_1589,N_1116);
or U2053 (N_2053,N_1025,N_1004);
nand U2054 (N_2054,N_1619,N_1981);
nand U2055 (N_2055,N_1418,N_1279);
nand U2056 (N_2056,N_1454,N_1868);
nor U2057 (N_2057,N_1193,N_1261);
nor U2058 (N_2058,N_1739,N_1409);
nand U2059 (N_2059,N_1966,N_1482);
and U2060 (N_2060,N_1671,N_1861);
or U2061 (N_2061,N_1176,N_1451);
and U2062 (N_2062,N_1787,N_1111);
nor U2063 (N_2063,N_1512,N_1305);
or U2064 (N_2064,N_1443,N_1252);
or U2065 (N_2065,N_1588,N_1178);
or U2066 (N_2066,N_1828,N_1431);
nor U2067 (N_2067,N_1232,N_1545);
nand U2068 (N_2068,N_1477,N_1175);
or U2069 (N_2069,N_1859,N_1437);
and U2070 (N_2070,N_1096,N_1923);
and U2071 (N_2071,N_1459,N_1964);
and U2072 (N_2072,N_1622,N_1468);
nor U2073 (N_2073,N_1847,N_1959);
nand U2074 (N_2074,N_1264,N_1118);
or U2075 (N_2075,N_1755,N_1023);
nand U2076 (N_2076,N_1380,N_1249);
nand U2077 (N_2077,N_1067,N_1625);
xnor U2078 (N_2078,N_1027,N_1376);
and U2079 (N_2079,N_1406,N_1604);
or U2080 (N_2080,N_1322,N_1807);
nand U2081 (N_2081,N_1105,N_1939);
nor U2082 (N_2082,N_1403,N_1560);
nand U2083 (N_2083,N_1384,N_1737);
and U2084 (N_2084,N_1630,N_1427);
nand U2085 (N_2085,N_1146,N_1690);
nor U2086 (N_2086,N_1815,N_1003);
or U2087 (N_2087,N_1148,N_1707);
and U2088 (N_2088,N_1719,N_1100);
or U2089 (N_2089,N_1792,N_1585);
or U2090 (N_2090,N_1916,N_1372);
or U2091 (N_2091,N_1299,N_1896);
or U2092 (N_2092,N_1359,N_1210);
or U2093 (N_2093,N_1412,N_1654);
nand U2094 (N_2094,N_1017,N_1698);
nand U2095 (N_2095,N_1296,N_1394);
or U2096 (N_2096,N_1421,N_1744);
nor U2097 (N_2097,N_1165,N_1083);
nand U2098 (N_2098,N_1504,N_1295);
nor U2099 (N_2099,N_1759,N_1713);
nand U2100 (N_2100,N_1054,N_1114);
and U2101 (N_2101,N_1263,N_1294);
or U2102 (N_2102,N_1433,N_1014);
or U2103 (N_2103,N_1173,N_1743);
or U2104 (N_2104,N_1607,N_1169);
or U2105 (N_2105,N_1863,N_1987);
and U2106 (N_2106,N_1385,N_1899);
nand U2107 (N_2107,N_1873,N_1233);
nor U2108 (N_2108,N_1321,N_1932);
and U2109 (N_2109,N_1972,N_1084);
or U2110 (N_2110,N_1072,N_1877);
xor U2111 (N_2111,N_1736,N_1876);
and U2112 (N_2112,N_1694,N_1578);
nor U2113 (N_2113,N_1919,N_1881);
or U2114 (N_2114,N_1505,N_1862);
nor U2115 (N_2115,N_1559,N_1442);
or U2116 (N_2116,N_1506,N_1777);
xnor U2117 (N_2117,N_1833,N_1269);
or U2118 (N_2118,N_1287,N_1291);
or U2119 (N_2119,N_1936,N_1885);
or U2120 (N_2120,N_1569,N_1968);
nor U2121 (N_2121,N_1221,N_1662);
and U2122 (N_2122,N_1990,N_1340);
or U2123 (N_2123,N_1127,N_1164);
nand U2124 (N_2124,N_1688,N_1481);
nor U2125 (N_2125,N_1595,N_1115);
nor U2126 (N_2126,N_1989,N_1182);
nor U2127 (N_2127,N_1517,N_1413);
nand U2128 (N_2128,N_1798,N_1648);
nor U2129 (N_2129,N_1710,N_1089);
nand U2130 (N_2130,N_1218,N_1948);
nor U2131 (N_2131,N_1820,N_1323);
and U2132 (N_2132,N_1611,N_1057);
nor U2133 (N_2133,N_1008,N_1620);
and U2134 (N_2134,N_1006,N_1940);
or U2135 (N_2135,N_1194,N_1824);
nor U2136 (N_2136,N_1224,N_1958);
nor U2137 (N_2137,N_1103,N_1928);
and U2138 (N_2138,N_1383,N_1976);
and U2139 (N_2139,N_1326,N_1068);
xor U2140 (N_2140,N_1270,N_1254);
nand U2141 (N_2141,N_1858,N_1695);
nand U2142 (N_2142,N_1276,N_1612);
and U2143 (N_2143,N_1931,N_1259);
xnor U2144 (N_2144,N_1660,N_1495);
and U2145 (N_2145,N_1912,N_1659);
nand U2146 (N_2146,N_1131,N_1309);
and U2147 (N_2147,N_1538,N_1999);
xnor U2148 (N_2148,N_1368,N_1147);
xnor U2149 (N_2149,N_1044,N_1056);
nor U2150 (N_2150,N_1764,N_1592);
nor U2151 (N_2151,N_1187,N_1189);
nand U2152 (N_2152,N_1525,N_1786);
nand U2153 (N_2153,N_1040,N_1922);
nor U2154 (N_2154,N_1703,N_1489);
nand U2155 (N_2155,N_1890,N_1969);
nor U2156 (N_2156,N_1519,N_1962);
or U2157 (N_2157,N_1752,N_1311);
or U2158 (N_2158,N_1298,N_1405);
or U2159 (N_2159,N_1603,N_1658);
or U2160 (N_2160,N_1282,N_1142);
nor U2161 (N_2161,N_1250,N_1908);
nor U2162 (N_2162,N_1854,N_1797);
nor U2163 (N_2163,N_1657,N_1834);
nand U2164 (N_2164,N_1870,N_1157);
nand U2165 (N_2165,N_1945,N_1977);
nor U2166 (N_2166,N_1575,N_1943);
and U2167 (N_2167,N_1801,N_1317);
nand U2168 (N_2168,N_1827,N_1365);
and U2169 (N_2169,N_1190,N_1692);
nand U2170 (N_2170,N_1839,N_1900);
or U2171 (N_2171,N_1720,N_1155);
or U2172 (N_2172,N_1917,N_1678);
nor U2173 (N_2173,N_1714,N_1911);
nor U2174 (N_2174,N_1015,N_1149);
and U2175 (N_2175,N_1060,N_1154);
and U2176 (N_2176,N_1484,N_1310);
nor U2177 (N_2177,N_1196,N_1823);
or U2178 (N_2178,N_1161,N_1135);
or U2179 (N_2179,N_1850,N_1544);
or U2180 (N_2180,N_1393,N_1967);
and U2181 (N_2181,N_1216,N_1767);
nor U2182 (N_2182,N_1857,N_1171);
or U2183 (N_2183,N_1324,N_1774);
nor U2184 (N_2184,N_1582,N_1058);
or U2185 (N_2185,N_1016,N_1509);
and U2186 (N_2186,N_1909,N_1422);
or U2187 (N_2187,N_1350,N_1242);
or U2188 (N_2188,N_1758,N_1770);
nor U2189 (N_2189,N_1346,N_1104);
nand U2190 (N_2190,N_1904,N_1645);
nor U2191 (N_2191,N_1783,N_1110);
xnor U2192 (N_2192,N_1921,N_1816);
xnor U2193 (N_2193,N_1388,N_1426);
nand U2194 (N_2194,N_1170,N_1273);
nor U2195 (N_2195,N_1649,N_1086);
or U2196 (N_2196,N_1590,N_1722);
or U2197 (N_2197,N_1511,N_1831);
nand U2198 (N_2198,N_1458,N_1132);
and U2199 (N_2199,N_1835,N_1957);
or U2200 (N_2200,N_1352,N_1717);
and U2201 (N_2201,N_1887,N_1641);
nand U2202 (N_2202,N_1071,N_1172);
nand U2203 (N_2203,N_1746,N_1567);
nand U2204 (N_2204,N_1059,N_1546);
and U2205 (N_2205,N_1844,N_1961);
or U2206 (N_2206,N_1880,N_1647);
nand U2207 (N_2207,N_1738,N_1530);
and U2208 (N_2208,N_1290,N_1328);
nor U2209 (N_2209,N_1130,N_1865);
nand U2210 (N_2210,N_1204,N_1069);
nand U2211 (N_2211,N_1846,N_1297);
nand U2212 (N_2212,N_1892,N_1950);
nor U2213 (N_2213,N_1217,N_1778);
and U2214 (N_2214,N_1280,N_1000);
or U2215 (N_2215,N_1094,N_1818);
and U2216 (N_2216,N_1386,N_1034);
nand U2217 (N_2217,N_1198,N_1446);
nand U2218 (N_2218,N_1402,N_1301);
nand U2219 (N_2219,N_1669,N_1152);
and U2220 (N_2220,N_1864,N_1753);
and U2221 (N_2221,N_1686,N_1005);
nor U2222 (N_2222,N_1450,N_1757);
or U2223 (N_2223,N_1448,N_1993);
nand U2224 (N_2224,N_1971,N_1822);
nor U2225 (N_2225,N_1536,N_1336);
nor U2226 (N_2226,N_1748,N_1565);
nand U2227 (N_2227,N_1497,N_1126);
and U2228 (N_2228,N_1927,N_1030);
or U2229 (N_2229,N_1606,N_1214);
nand U2230 (N_2230,N_1986,N_1529);
or U2231 (N_2231,N_1853,N_1754);
nand U2232 (N_2232,N_1139,N_1564);
nand U2233 (N_2233,N_1244,N_1556);
and U2234 (N_2234,N_1518,N_1493);
or U2235 (N_2235,N_1011,N_1339);
nor U2236 (N_2236,N_1532,N_1338);
nand U2237 (N_2237,N_1615,N_1061);
nand U2238 (N_2238,N_1226,N_1367);
nand U2239 (N_2239,N_1434,N_1679);
nand U2240 (N_2240,N_1605,N_1240);
or U2241 (N_2241,N_1524,N_1727);
or U2242 (N_2242,N_1197,N_1203);
or U2243 (N_2243,N_1441,N_1732);
nand U2244 (N_2244,N_1082,N_1836);
and U2245 (N_2245,N_1177,N_1274);
and U2246 (N_2246,N_1646,N_1275);
or U2247 (N_2247,N_1624,N_1879);
and U2248 (N_2248,N_1199,N_1676);
or U2249 (N_2249,N_1408,N_1026);
or U2250 (N_2250,N_1851,N_1579);
nand U2251 (N_2251,N_1303,N_1137);
nand U2252 (N_2252,N_1430,N_1075);
nand U2253 (N_2253,N_1803,N_1113);
and U2254 (N_2254,N_1804,N_1185);
and U2255 (N_2255,N_1821,N_1985);
nand U2256 (N_2256,N_1563,N_1665);
nand U2257 (N_2257,N_1573,N_1596);
or U2258 (N_2258,N_1074,N_1202);
nand U2259 (N_2259,N_1209,N_1740);
nor U2260 (N_2260,N_1219,N_1656);
nand U2261 (N_2261,N_1361,N_1784);
nand U2262 (N_2262,N_1001,N_1417);
or U2263 (N_2263,N_1956,N_1915);
nor U2264 (N_2264,N_1306,N_1288);
nor U2265 (N_2265,N_1253,N_1845);
nand U2266 (N_2266,N_1095,N_1188);
or U2267 (N_2267,N_1734,N_1782);
or U2268 (N_2268,N_1195,N_1651);
or U2269 (N_2269,N_1549,N_1156);
or U2270 (N_2270,N_1143,N_1918);
and U2271 (N_2271,N_1160,N_1174);
nor U2272 (N_2272,N_1769,N_1121);
nand U2273 (N_2273,N_1432,N_1772);
xnor U2274 (N_2274,N_1366,N_1047);
and U2275 (N_2275,N_1153,N_1602);
and U2276 (N_2276,N_1539,N_1897);
nor U2277 (N_2277,N_1231,N_1475);
and U2278 (N_2278,N_1663,N_1181);
or U2279 (N_2279,N_1960,N_1982);
nand U2280 (N_2280,N_1735,N_1799);
and U2281 (N_2281,N_1150,N_1077);
nand U2282 (N_2282,N_1938,N_1162);
nor U2283 (N_2283,N_1241,N_1500);
and U2284 (N_2284,N_1461,N_1070);
and U2285 (N_2285,N_1112,N_1723);
or U2286 (N_2286,N_1503,N_1483);
nand U2287 (N_2287,N_1235,N_1984);
or U2288 (N_2288,N_1354,N_1414);
nor U2289 (N_2289,N_1901,N_1080);
or U2290 (N_2290,N_1806,N_1102);
nand U2291 (N_2291,N_1145,N_1552);
or U2292 (N_2292,N_1832,N_1768);
nor U2293 (N_2293,N_1840,N_1262);
nand U2294 (N_2294,N_1705,N_1251);
nor U2295 (N_2295,N_1642,N_1277);
and U2296 (N_2296,N_1934,N_1682);
nand U2297 (N_2297,N_1348,N_1211);
and U2298 (N_2298,N_1470,N_1508);
nor U2299 (N_2299,N_1474,N_1628);
and U2300 (N_2300,N_1223,N_1460);
nor U2301 (N_2301,N_1389,N_1947);
or U2302 (N_2302,N_1236,N_1523);
nand U2303 (N_2303,N_1420,N_1184);
nor U2304 (N_2304,N_1478,N_1627);
or U2305 (N_2305,N_1942,N_1360);
and U2306 (N_2306,N_1558,N_1930);
or U2307 (N_2307,N_1685,N_1449);
and U2308 (N_2308,N_1179,N_1467);
nor U2309 (N_2309,N_1363,N_1019);
nor U2310 (N_2310,N_1515,N_1024);
or U2311 (N_2311,N_1973,N_1410);
and U2312 (N_2312,N_1825,N_1860);
nand U2313 (N_2313,N_1741,N_1526);
nor U2314 (N_2314,N_1598,N_1237);
nand U2315 (N_2315,N_1212,N_1213);
nand U2316 (N_2316,N_1415,N_1581);
nor U2317 (N_2317,N_1227,N_1342);
and U2318 (N_2318,N_1046,N_1843);
nor U2319 (N_2319,N_1941,N_1542);
and U2320 (N_2320,N_1742,N_1002);
nor U2321 (N_2321,N_1479,N_1572);
or U2322 (N_2322,N_1775,N_1436);
or U2323 (N_2323,N_1397,N_1697);
nor U2324 (N_2324,N_1933,N_1548);
nor U2325 (N_2325,N_1480,N_1711);
or U2326 (N_2326,N_1988,N_1547);
and U2327 (N_2327,N_1022,N_1039);
nor U2328 (N_2328,N_1392,N_1239);
nand U2329 (N_2329,N_1954,N_1842);
or U2330 (N_2330,N_1399,N_1268);
and U2331 (N_2331,N_1283,N_1895);
and U2332 (N_2332,N_1810,N_1680);
nor U2333 (N_2333,N_1540,N_1037);
and U2334 (N_2334,N_1913,N_1400);
nand U2335 (N_2335,N_1007,N_1337);
nand U2336 (N_2336,N_1674,N_1963);
and U2337 (N_2337,N_1496,N_1401);
nor U2338 (N_2338,N_1780,N_1566);
nor U2339 (N_2339,N_1379,N_1494);
xor U2340 (N_2340,N_1109,N_1272);
and U2341 (N_2341,N_1574,N_1618);
nor U2342 (N_2342,N_1266,N_1438);
nand U2343 (N_2343,N_1119,N_1498);
and U2344 (N_2344,N_1888,N_1440);
nor U2345 (N_2345,N_1750,N_1762);
nor U2346 (N_2346,N_1107,N_1293);
xnor U2347 (N_2347,N_1093,N_1955);
and U2348 (N_2348,N_1330,N_1374);
nand U2349 (N_2349,N_1979,N_1706);
nor U2350 (N_2350,N_1499,N_1745);
or U2351 (N_2351,N_1681,N_1871);
nor U2352 (N_2352,N_1788,N_1667);
or U2353 (N_2353,N_1878,N_1910);
and U2354 (N_2354,N_1238,N_1476);
nand U2355 (N_2355,N_1537,N_1886);
nand U2356 (N_2356,N_1721,N_1924);
nand U2357 (N_2357,N_1428,N_1661);
nor U2358 (N_2358,N_1701,N_1314);
or U2359 (N_2359,N_1914,N_1382);
nand U2360 (N_2360,N_1733,N_1583);
nand U2361 (N_2361,N_1747,N_1594);
and U2362 (N_2362,N_1884,N_1215);
or U2363 (N_2363,N_1245,N_1304);
and U2364 (N_2364,N_1125,N_1584);
or U2365 (N_2365,N_1159,N_1882);
nor U2366 (N_2366,N_1315,N_1230);
nand U2367 (N_2367,N_1345,N_1576);
nand U2368 (N_2368,N_1141,N_1370);
nand U2369 (N_2369,N_1805,N_1099);
and U2370 (N_2370,N_1124,N_1510);
and U2371 (N_2371,N_1055,N_1180);
nor U2372 (N_2372,N_1281,N_1937);
nor U2373 (N_2373,N_1471,N_1837);
nand U2374 (N_2374,N_1696,N_1183);
or U2375 (N_2375,N_1128,N_1362);
nor U2376 (N_2376,N_1841,N_1201);
nor U2377 (N_2377,N_1629,N_1997);
nand U2378 (N_2378,N_1812,N_1316);
nor U2379 (N_2379,N_1329,N_1411);
and U2380 (N_2380,N_1905,N_1318);
or U2381 (N_2381,N_1983,N_1635);
nand U2382 (N_2382,N_1243,N_1031);
and U2383 (N_2383,N_1849,N_1090);
nor U2384 (N_2384,N_1041,N_1191);
nor U2385 (N_2385,N_1926,N_1613);
or U2386 (N_2386,N_1715,N_1621);
nand U2387 (N_2387,N_1286,N_1728);
nand U2388 (N_2388,N_1063,N_1513);
and U2389 (N_2389,N_1085,N_1462);
nand U2390 (N_2390,N_1088,N_1313);
nor U2391 (N_2391,N_1633,N_1814);
nand U2392 (N_2392,N_1327,N_1013);
and U2393 (N_2393,N_1520,N_1994);
nand U2394 (N_2394,N_1229,N_1852);
and U2395 (N_2395,N_1826,N_1335);
nor U2396 (N_2396,N_1333,N_1790);
and U2397 (N_2397,N_1761,N_1343);
or U2398 (N_2398,N_1465,N_1469);
or U2399 (N_2399,N_1995,N_1396);
or U2400 (N_2400,N_1404,N_1257);
nor U2401 (N_2401,N_1712,N_1271);
xor U2402 (N_2402,N_1756,N_1065);
or U2403 (N_2403,N_1344,N_1992);
or U2404 (N_2404,N_1225,N_1138);
nor U2405 (N_2405,N_1533,N_1935);
nand U2406 (N_2406,N_1200,N_1848);
nand U2407 (N_2407,N_1683,N_1944);
and U2408 (N_2408,N_1491,N_1623);
nand U2409 (N_2409,N_1516,N_1028);
nor U2410 (N_2410,N_1289,N_1136);
and U2411 (N_2411,N_1234,N_1906);
nor U2412 (N_2412,N_1687,N_1435);
nand U2413 (N_2413,N_1773,N_1577);
nand U2414 (N_2414,N_1076,N_1097);
nand U2415 (N_2415,N_1891,N_1453);
or U2416 (N_2416,N_1608,N_1032);
and U2417 (N_2417,N_1541,N_1568);
and U2418 (N_2418,N_1122,N_1098);
or U2419 (N_2419,N_1358,N_1693);
or U2420 (N_2420,N_1751,N_1247);
nor U2421 (N_2421,N_1158,N_1091);
nor U2422 (N_2422,N_1571,N_1898);
nor U2423 (N_2423,N_1970,N_1018);
and U2424 (N_2424,N_1207,N_1531);
nor U2425 (N_2425,N_1597,N_1048);
and U2426 (N_2426,N_1553,N_1675);
or U2427 (N_2427,N_1042,N_1691);
nor U2428 (N_2428,N_1802,N_1463);
nand U2429 (N_2429,N_1073,N_1653);
nor U2430 (N_2430,N_1655,N_1049);
and U2431 (N_2431,N_1168,N_1980);
nor U2432 (N_2432,N_1689,N_1447);
nor U2433 (N_2433,N_1010,N_1920);
nor U2434 (N_2434,N_1355,N_1925);
or U2435 (N_2435,N_1192,N_1670);
and U2436 (N_2436,N_1684,N_1749);
nor U2437 (N_2437,N_1929,N_1779);
nand U2438 (N_2438,N_1949,N_1789);
or U2439 (N_2439,N_1830,N_1036);
and U2440 (N_2440,N_1867,N_1429);
and U2441 (N_2441,N_1457,N_1726);
or U2442 (N_2442,N_1186,N_1672);
nor U2443 (N_2443,N_1855,N_1341);
nand U2444 (N_2444,N_1319,N_1631);
nand U2445 (N_2445,N_1398,N_1637);
xor U2446 (N_2446,N_1978,N_1586);
and U2447 (N_2447,N_1349,N_1357);
nor U2448 (N_2448,N_1760,N_1206);
nor U2449 (N_2449,N_1562,N_1364);
and U2450 (N_2450,N_1325,N_1501);
nor U2451 (N_2451,N_1258,N_1220);
nand U2452 (N_2452,N_1267,N_1425);
nand U2453 (N_2453,N_1492,N_1724);
nand U2454 (N_2454,N_1144,N_1609);
nand U2455 (N_2455,N_1163,N_1664);
and U2456 (N_2456,N_1308,N_1591);
and U2457 (N_2457,N_1407,N_1528);
and U2458 (N_2458,N_1599,N_1763);
nor U2459 (N_2459,N_1079,N_1038);
nor U2460 (N_2460,N_1445,N_1140);
nor U2461 (N_2461,N_1527,N_1776);
and U2462 (N_2462,N_1260,N_1902);
nor U2463 (N_2463,N_1829,N_1285);
and U2464 (N_2464,N_1570,N_1391);
nor U2465 (N_2465,N_1700,N_1838);
or U2466 (N_2466,N_1514,N_1593);
nor U2467 (N_2467,N_1064,N_1452);
nor U2468 (N_2468,N_1378,N_1020);
and U2469 (N_2469,N_1652,N_1375);
nor U2470 (N_2470,N_1248,N_1869);
or U2471 (N_2471,N_1866,N_1332);
and U2472 (N_2472,N_1561,N_1369);
or U2473 (N_2473,N_1166,N_1794);
nand U2474 (N_2474,N_1677,N_1009);
nand U2475 (N_2475,N_1381,N_1636);
nand U2476 (N_2476,N_1809,N_1580);
and U2477 (N_2477,N_1617,N_1731);
or U2478 (N_2478,N_1946,N_1557);
nand U2479 (N_2479,N_1351,N_1965);
and U2480 (N_2480,N_1699,N_1704);
and U2481 (N_2481,N_1883,N_1300);
and U2482 (N_2482,N_1106,N_1222);
nor U2483 (N_2483,N_1033,N_1702);
and U2484 (N_2484,N_1419,N_1387);
nand U2485 (N_2485,N_1998,N_1334);
or U2486 (N_2486,N_1487,N_1874);
nor U2487 (N_2487,N_1587,N_1640);
or U2488 (N_2488,N_1610,N_1377);
and U2489 (N_2489,N_1108,N_1356);
and U2490 (N_2490,N_1134,N_1793);
and U2491 (N_2491,N_1078,N_1554);
nor U2492 (N_2492,N_1875,N_1472);
nor U2493 (N_2493,N_1616,N_1045);
and U2494 (N_2494,N_1951,N_1256);
nand U2495 (N_2495,N_1331,N_1813);
and U2496 (N_2496,N_1117,N_1614);
nand U2497 (N_2497,N_1551,N_1087);
or U2498 (N_2498,N_1167,N_1795);
and U2499 (N_2499,N_1053,N_1466);
or U2500 (N_2500,N_1943,N_1067);
and U2501 (N_2501,N_1416,N_1052);
and U2502 (N_2502,N_1416,N_1139);
and U2503 (N_2503,N_1034,N_1363);
nand U2504 (N_2504,N_1991,N_1627);
and U2505 (N_2505,N_1019,N_1068);
nand U2506 (N_2506,N_1772,N_1195);
nand U2507 (N_2507,N_1503,N_1465);
nor U2508 (N_2508,N_1482,N_1148);
or U2509 (N_2509,N_1875,N_1809);
xor U2510 (N_2510,N_1584,N_1281);
and U2511 (N_2511,N_1405,N_1846);
nand U2512 (N_2512,N_1037,N_1333);
nor U2513 (N_2513,N_1521,N_1149);
or U2514 (N_2514,N_1663,N_1155);
nor U2515 (N_2515,N_1212,N_1670);
and U2516 (N_2516,N_1363,N_1120);
nand U2517 (N_2517,N_1845,N_1602);
or U2518 (N_2518,N_1557,N_1273);
nor U2519 (N_2519,N_1394,N_1061);
and U2520 (N_2520,N_1302,N_1301);
and U2521 (N_2521,N_1615,N_1040);
nor U2522 (N_2522,N_1420,N_1737);
or U2523 (N_2523,N_1136,N_1071);
or U2524 (N_2524,N_1402,N_1243);
xor U2525 (N_2525,N_1500,N_1572);
nor U2526 (N_2526,N_1886,N_1625);
and U2527 (N_2527,N_1074,N_1285);
nor U2528 (N_2528,N_1768,N_1238);
or U2529 (N_2529,N_1288,N_1709);
or U2530 (N_2530,N_1989,N_1197);
xnor U2531 (N_2531,N_1108,N_1530);
or U2532 (N_2532,N_1843,N_1814);
nand U2533 (N_2533,N_1648,N_1484);
nor U2534 (N_2534,N_1710,N_1967);
nand U2535 (N_2535,N_1498,N_1389);
nand U2536 (N_2536,N_1120,N_1194);
nand U2537 (N_2537,N_1726,N_1434);
nand U2538 (N_2538,N_1442,N_1233);
or U2539 (N_2539,N_1024,N_1349);
and U2540 (N_2540,N_1040,N_1855);
or U2541 (N_2541,N_1306,N_1829);
nor U2542 (N_2542,N_1799,N_1456);
or U2543 (N_2543,N_1913,N_1017);
nand U2544 (N_2544,N_1587,N_1405);
nor U2545 (N_2545,N_1884,N_1478);
and U2546 (N_2546,N_1017,N_1640);
nor U2547 (N_2547,N_1077,N_1482);
or U2548 (N_2548,N_1880,N_1892);
nand U2549 (N_2549,N_1065,N_1749);
nor U2550 (N_2550,N_1140,N_1025);
or U2551 (N_2551,N_1054,N_1442);
nand U2552 (N_2552,N_1687,N_1262);
or U2553 (N_2553,N_1345,N_1868);
nand U2554 (N_2554,N_1309,N_1773);
nor U2555 (N_2555,N_1921,N_1066);
and U2556 (N_2556,N_1197,N_1273);
nand U2557 (N_2557,N_1241,N_1065);
nor U2558 (N_2558,N_1072,N_1355);
nor U2559 (N_2559,N_1227,N_1432);
and U2560 (N_2560,N_1865,N_1225);
nor U2561 (N_2561,N_1926,N_1540);
or U2562 (N_2562,N_1066,N_1429);
xor U2563 (N_2563,N_1066,N_1887);
nor U2564 (N_2564,N_1803,N_1911);
or U2565 (N_2565,N_1679,N_1300);
xor U2566 (N_2566,N_1236,N_1741);
nor U2567 (N_2567,N_1486,N_1840);
nor U2568 (N_2568,N_1879,N_1316);
or U2569 (N_2569,N_1094,N_1243);
nand U2570 (N_2570,N_1184,N_1963);
or U2571 (N_2571,N_1763,N_1402);
or U2572 (N_2572,N_1911,N_1167);
nand U2573 (N_2573,N_1261,N_1024);
or U2574 (N_2574,N_1407,N_1772);
or U2575 (N_2575,N_1210,N_1317);
xnor U2576 (N_2576,N_1288,N_1871);
nor U2577 (N_2577,N_1943,N_1715);
nor U2578 (N_2578,N_1780,N_1334);
nand U2579 (N_2579,N_1786,N_1105);
or U2580 (N_2580,N_1513,N_1735);
nor U2581 (N_2581,N_1115,N_1114);
and U2582 (N_2582,N_1765,N_1337);
or U2583 (N_2583,N_1217,N_1664);
nand U2584 (N_2584,N_1622,N_1267);
and U2585 (N_2585,N_1571,N_1041);
nor U2586 (N_2586,N_1305,N_1053);
and U2587 (N_2587,N_1040,N_1242);
and U2588 (N_2588,N_1366,N_1860);
or U2589 (N_2589,N_1861,N_1447);
or U2590 (N_2590,N_1384,N_1469);
nor U2591 (N_2591,N_1059,N_1922);
nand U2592 (N_2592,N_1452,N_1291);
xor U2593 (N_2593,N_1533,N_1664);
or U2594 (N_2594,N_1900,N_1293);
nor U2595 (N_2595,N_1591,N_1127);
or U2596 (N_2596,N_1404,N_1434);
nor U2597 (N_2597,N_1492,N_1639);
and U2598 (N_2598,N_1355,N_1010);
nand U2599 (N_2599,N_1427,N_1560);
nor U2600 (N_2600,N_1437,N_1019);
nor U2601 (N_2601,N_1987,N_1291);
and U2602 (N_2602,N_1333,N_1480);
nor U2603 (N_2603,N_1409,N_1431);
xnor U2604 (N_2604,N_1671,N_1346);
or U2605 (N_2605,N_1895,N_1813);
nand U2606 (N_2606,N_1102,N_1289);
or U2607 (N_2607,N_1961,N_1784);
nand U2608 (N_2608,N_1453,N_1257);
nor U2609 (N_2609,N_1044,N_1046);
or U2610 (N_2610,N_1859,N_1801);
nor U2611 (N_2611,N_1351,N_1957);
and U2612 (N_2612,N_1512,N_1547);
nor U2613 (N_2613,N_1036,N_1591);
and U2614 (N_2614,N_1963,N_1780);
nand U2615 (N_2615,N_1545,N_1999);
or U2616 (N_2616,N_1973,N_1433);
nor U2617 (N_2617,N_1376,N_1279);
and U2618 (N_2618,N_1792,N_1516);
or U2619 (N_2619,N_1932,N_1174);
nor U2620 (N_2620,N_1588,N_1586);
nand U2621 (N_2621,N_1273,N_1766);
nor U2622 (N_2622,N_1378,N_1236);
and U2623 (N_2623,N_1387,N_1151);
nor U2624 (N_2624,N_1574,N_1542);
nand U2625 (N_2625,N_1120,N_1572);
and U2626 (N_2626,N_1177,N_1295);
and U2627 (N_2627,N_1794,N_1208);
nand U2628 (N_2628,N_1664,N_1433);
or U2629 (N_2629,N_1061,N_1030);
nor U2630 (N_2630,N_1572,N_1336);
nand U2631 (N_2631,N_1041,N_1237);
nand U2632 (N_2632,N_1804,N_1897);
nor U2633 (N_2633,N_1211,N_1296);
nor U2634 (N_2634,N_1317,N_1788);
nor U2635 (N_2635,N_1660,N_1063);
nand U2636 (N_2636,N_1073,N_1470);
and U2637 (N_2637,N_1950,N_1371);
and U2638 (N_2638,N_1092,N_1372);
and U2639 (N_2639,N_1345,N_1321);
nand U2640 (N_2640,N_1487,N_1237);
and U2641 (N_2641,N_1822,N_1320);
nor U2642 (N_2642,N_1226,N_1546);
and U2643 (N_2643,N_1853,N_1778);
nand U2644 (N_2644,N_1681,N_1360);
nand U2645 (N_2645,N_1160,N_1882);
nor U2646 (N_2646,N_1693,N_1022);
nand U2647 (N_2647,N_1974,N_1980);
nand U2648 (N_2648,N_1400,N_1060);
nor U2649 (N_2649,N_1919,N_1820);
nor U2650 (N_2650,N_1206,N_1170);
and U2651 (N_2651,N_1039,N_1996);
or U2652 (N_2652,N_1647,N_1891);
and U2653 (N_2653,N_1124,N_1846);
nand U2654 (N_2654,N_1819,N_1901);
and U2655 (N_2655,N_1804,N_1358);
or U2656 (N_2656,N_1731,N_1414);
nand U2657 (N_2657,N_1965,N_1783);
and U2658 (N_2658,N_1253,N_1625);
or U2659 (N_2659,N_1577,N_1505);
nand U2660 (N_2660,N_1164,N_1408);
nor U2661 (N_2661,N_1160,N_1614);
or U2662 (N_2662,N_1368,N_1206);
and U2663 (N_2663,N_1183,N_1161);
nor U2664 (N_2664,N_1649,N_1446);
nor U2665 (N_2665,N_1840,N_1221);
nor U2666 (N_2666,N_1187,N_1862);
nand U2667 (N_2667,N_1169,N_1675);
or U2668 (N_2668,N_1058,N_1306);
and U2669 (N_2669,N_1947,N_1469);
xnor U2670 (N_2670,N_1560,N_1265);
xor U2671 (N_2671,N_1803,N_1849);
nor U2672 (N_2672,N_1405,N_1290);
nor U2673 (N_2673,N_1489,N_1303);
nor U2674 (N_2674,N_1626,N_1999);
or U2675 (N_2675,N_1644,N_1335);
nor U2676 (N_2676,N_1633,N_1121);
nor U2677 (N_2677,N_1378,N_1159);
or U2678 (N_2678,N_1919,N_1917);
or U2679 (N_2679,N_1593,N_1091);
or U2680 (N_2680,N_1223,N_1175);
nor U2681 (N_2681,N_1009,N_1429);
or U2682 (N_2682,N_1384,N_1576);
nor U2683 (N_2683,N_1921,N_1138);
nor U2684 (N_2684,N_1858,N_1089);
nand U2685 (N_2685,N_1992,N_1811);
or U2686 (N_2686,N_1188,N_1153);
nor U2687 (N_2687,N_1826,N_1003);
and U2688 (N_2688,N_1718,N_1548);
and U2689 (N_2689,N_1453,N_1996);
and U2690 (N_2690,N_1749,N_1296);
and U2691 (N_2691,N_1632,N_1332);
or U2692 (N_2692,N_1720,N_1484);
or U2693 (N_2693,N_1218,N_1558);
and U2694 (N_2694,N_1105,N_1126);
or U2695 (N_2695,N_1124,N_1689);
nor U2696 (N_2696,N_1761,N_1071);
nand U2697 (N_2697,N_1149,N_1725);
nor U2698 (N_2698,N_1183,N_1647);
nor U2699 (N_2699,N_1169,N_1447);
nand U2700 (N_2700,N_1008,N_1370);
nor U2701 (N_2701,N_1648,N_1594);
and U2702 (N_2702,N_1681,N_1540);
nand U2703 (N_2703,N_1231,N_1746);
or U2704 (N_2704,N_1504,N_1159);
and U2705 (N_2705,N_1713,N_1704);
nor U2706 (N_2706,N_1529,N_1102);
nand U2707 (N_2707,N_1577,N_1948);
and U2708 (N_2708,N_1962,N_1168);
nor U2709 (N_2709,N_1667,N_1110);
or U2710 (N_2710,N_1434,N_1420);
nor U2711 (N_2711,N_1334,N_1658);
and U2712 (N_2712,N_1809,N_1346);
and U2713 (N_2713,N_1216,N_1668);
and U2714 (N_2714,N_1247,N_1078);
nand U2715 (N_2715,N_1717,N_1254);
nand U2716 (N_2716,N_1812,N_1352);
nand U2717 (N_2717,N_1337,N_1537);
nand U2718 (N_2718,N_1851,N_1513);
or U2719 (N_2719,N_1340,N_1873);
and U2720 (N_2720,N_1040,N_1651);
nand U2721 (N_2721,N_1537,N_1508);
or U2722 (N_2722,N_1540,N_1692);
and U2723 (N_2723,N_1406,N_1787);
and U2724 (N_2724,N_1705,N_1666);
or U2725 (N_2725,N_1707,N_1964);
nand U2726 (N_2726,N_1724,N_1989);
or U2727 (N_2727,N_1599,N_1906);
nand U2728 (N_2728,N_1892,N_1051);
or U2729 (N_2729,N_1789,N_1690);
nand U2730 (N_2730,N_1873,N_1833);
nand U2731 (N_2731,N_1615,N_1029);
nor U2732 (N_2732,N_1126,N_1256);
and U2733 (N_2733,N_1684,N_1079);
xor U2734 (N_2734,N_1693,N_1397);
or U2735 (N_2735,N_1382,N_1801);
and U2736 (N_2736,N_1405,N_1580);
and U2737 (N_2737,N_1067,N_1676);
or U2738 (N_2738,N_1844,N_1108);
nand U2739 (N_2739,N_1846,N_1061);
nand U2740 (N_2740,N_1814,N_1116);
or U2741 (N_2741,N_1410,N_1493);
nor U2742 (N_2742,N_1054,N_1324);
or U2743 (N_2743,N_1116,N_1461);
and U2744 (N_2744,N_1656,N_1002);
nor U2745 (N_2745,N_1763,N_1795);
and U2746 (N_2746,N_1907,N_1817);
or U2747 (N_2747,N_1354,N_1751);
nor U2748 (N_2748,N_1485,N_1476);
nor U2749 (N_2749,N_1818,N_1308);
or U2750 (N_2750,N_1487,N_1717);
nor U2751 (N_2751,N_1306,N_1401);
nand U2752 (N_2752,N_1140,N_1268);
nor U2753 (N_2753,N_1404,N_1955);
xor U2754 (N_2754,N_1188,N_1240);
nor U2755 (N_2755,N_1338,N_1150);
nor U2756 (N_2756,N_1938,N_1986);
and U2757 (N_2757,N_1124,N_1706);
nand U2758 (N_2758,N_1950,N_1959);
nand U2759 (N_2759,N_1172,N_1338);
xnor U2760 (N_2760,N_1970,N_1999);
nor U2761 (N_2761,N_1649,N_1553);
or U2762 (N_2762,N_1496,N_1949);
and U2763 (N_2763,N_1549,N_1650);
or U2764 (N_2764,N_1304,N_1473);
or U2765 (N_2765,N_1256,N_1149);
and U2766 (N_2766,N_1273,N_1889);
nor U2767 (N_2767,N_1835,N_1104);
nand U2768 (N_2768,N_1012,N_1035);
and U2769 (N_2769,N_1441,N_1840);
and U2770 (N_2770,N_1642,N_1129);
and U2771 (N_2771,N_1929,N_1298);
nand U2772 (N_2772,N_1914,N_1273);
and U2773 (N_2773,N_1857,N_1676);
nand U2774 (N_2774,N_1220,N_1396);
or U2775 (N_2775,N_1621,N_1087);
nor U2776 (N_2776,N_1373,N_1032);
nor U2777 (N_2777,N_1956,N_1150);
and U2778 (N_2778,N_1390,N_1447);
or U2779 (N_2779,N_1745,N_1362);
nor U2780 (N_2780,N_1319,N_1935);
nor U2781 (N_2781,N_1262,N_1400);
and U2782 (N_2782,N_1091,N_1499);
nor U2783 (N_2783,N_1982,N_1076);
nor U2784 (N_2784,N_1074,N_1315);
nor U2785 (N_2785,N_1973,N_1006);
nand U2786 (N_2786,N_1837,N_1136);
or U2787 (N_2787,N_1037,N_1095);
nor U2788 (N_2788,N_1311,N_1309);
nand U2789 (N_2789,N_1924,N_1707);
nand U2790 (N_2790,N_1406,N_1694);
or U2791 (N_2791,N_1765,N_1321);
nand U2792 (N_2792,N_1935,N_1435);
and U2793 (N_2793,N_1367,N_1406);
and U2794 (N_2794,N_1340,N_1134);
and U2795 (N_2795,N_1343,N_1243);
and U2796 (N_2796,N_1537,N_1224);
nand U2797 (N_2797,N_1341,N_1701);
nand U2798 (N_2798,N_1190,N_1104);
or U2799 (N_2799,N_1542,N_1624);
and U2800 (N_2800,N_1256,N_1190);
nor U2801 (N_2801,N_1371,N_1910);
nand U2802 (N_2802,N_1835,N_1356);
nor U2803 (N_2803,N_1620,N_1720);
nor U2804 (N_2804,N_1052,N_1879);
xnor U2805 (N_2805,N_1610,N_1155);
nand U2806 (N_2806,N_1750,N_1744);
nand U2807 (N_2807,N_1898,N_1534);
nand U2808 (N_2808,N_1334,N_1971);
nand U2809 (N_2809,N_1587,N_1767);
nand U2810 (N_2810,N_1843,N_1548);
or U2811 (N_2811,N_1197,N_1156);
or U2812 (N_2812,N_1730,N_1808);
and U2813 (N_2813,N_1176,N_1029);
nor U2814 (N_2814,N_1879,N_1120);
and U2815 (N_2815,N_1567,N_1375);
xor U2816 (N_2816,N_1364,N_1113);
and U2817 (N_2817,N_1487,N_1682);
and U2818 (N_2818,N_1755,N_1787);
or U2819 (N_2819,N_1603,N_1749);
nor U2820 (N_2820,N_1440,N_1399);
nand U2821 (N_2821,N_1818,N_1399);
or U2822 (N_2822,N_1692,N_1864);
or U2823 (N_2823,N_1319,N_1261);
or U2824 (N_2824,N_1562,N_1305);
and U2825 (N_2825,N_1407,N_1347);
and U2826 (N_2826,N_1562,N_1623);
nand U2827 (N_2827,N_1291,N_1348);
nand U2828 (N_2828,N_1542,N_1568);
and U2829 (N_2829,N_1132,N_1319);
nand U2830 (N_2830,N_1922,N_1244);
nor U2831 (N_2831,N_1961,N_1041);
and U2832 (N_2832,N_1203,N_1094);
nor U2833 (N_2833,N_1652,N_1115);
nor U2834 (N_2834,N_1841,N_1670);
or U2835 (N_2835,N_1412,N_1703);
nor U2836 (N_2836,N_1827,N_1616);
xnor U2837 (N_2837,N_1560,N_1385);
nand U2838 (N_2838,N_1881,N_1055);
and U2839 (N_2839,N_1335,N_1174);
or U2840 (N_2840,N_1254,N_1358);
or U2841 (N_2841,N_1645,N_1936);
nand U2842 (N_2842,N_1931,N_1362);
nand U2843 (N_2843,N_1661,N_1822);
and U2844 (N_2844,N_1757,N_1083);
or U2845 (N_2845,N_1400,N_1469);
and U2846 (N_2846,N_1914,N_1543);
nor U2847 (N_2847,N_1121,N_1360);
nor U2848 (N_2848,N_1944,N_1659);
nand U2849 (N_2849,N_1904,N_1206);
or U2850 (N_2850,N_1908,N_1995);
nor U2851 (N_2851,N_1887,N_1474);
and U2852 (N_2852,N_1587,N_1875);
nand U2853 (N_2853,N_1567,N_1777);
nor U2854 (N_2854,N_1895,N_1643);
nor U2855 (N_2855,N_1915,N_1432);
nand U2856 (N_2856,N_1619,N_1005);
nor U2857 (N_2857,N_1425,N_1883);
and U2858 (N_2858,N_1864,N_1160);
nor U2859 (N_2859,N_1025,N_1481);
xor U2860 (N_2860,N_1885,N_1077);
and U2861 (N_2861,N_1072,N_1064);
nor U2862 (N_2862,N_1514,N_1432);
nand U2863 (N_2863,N_1727,N_1222);
nand U2864 (N_2864,N_1288,N_1229);
nor U2865 (N_2865,N_1266,N_1743);
and U2866 (N_2866,N_1518,N_1923);
nand U2867 (N_2867,N_1928,N_1253);
nand U2868 (N_2868,N_1886,N_1978);
nand U2869 (N_2869,N_1645,N_1586);
nor U2870 (N_2870,N_1706,N_1200);
or U2871 (N_2871,N_1669,N_1234);
nand U2872 (N_2872,N_1856,N_1738);
nor U2873 (N_2873,N_1349,N_1225);
nand U2874 (N_2874,N_1315,N_1632);
nand U2875 (N_2875,N_1877,N_1325);
or U2876 (N_2876,N_1616,N_1506);
and U2877 (N_2877,N_1476,N_1838);
and U2878 (N_2878,N_1166,N_1721);
and U2879 (N_2879,N_1001,N_1419);
nand U2880 (N_2880,N_1179,N_1822);
nor U2881 (N_2881,N_1608,N_1793);
nand U2882 (N_2882,N_1862,N_1942);
or U2883 (N_2883,N_1717,N_1817);
or U2884 (N_2884,N_1992,N_1579);
nand U2885 (N_2885,N_1591,N_1605);
or U2886 (N_2886,N_1318,N_1641);
and U2887 (N_2887,N_1923,N_1059);
and U2888 (N_2888,N_1834,N_1989);
nor U2889 (N_2889,N_1565,N_1141);
nand U2890 (N_2890,N_1145,N_1338);
nand U2891 (N_2891,N_1017,N_1301);
nand U2892 (N_2892,N_1108,N_1109);
and U2893 (N_2893,N_1808,N_1292);
and U2894 (N_2894,N_1602,N_1998);
and U2895 (N_2895,N_1194,N_1527);
or U2896 (N_2896,N_1057,N_1688);
xnor U2897 (N_2897,N_1174,N_1471);
and U2898 (N_2898,N_1137,N_1960);
nand U2899 (N_2899,N_1833,N_1367);
nor U2900 (N_2900,N_1498,N_1675);
or U2901 (N_2901,N_1279,N_1837);
and U2902 (N_2902,N_1321,N_1359);
nand U2903 (N_2903,N_1608,N_1533);
or U2904 (N_2904,N_1013,N_1579);
and U2905 (N_2905,N_1948,N_1911);
and U2906 (N_2906,N_1414,N_1392);
nor U2907 (N_2907,N_1081,N_1575);
or U2908 (N_2908,N_1725,N_1768);
nand U2909 (N_2909,N_1369,N_1059);
and U2910 (N_2910,N_1166,N_1124);
nand U2911 (N_2911,N_1475,N_1628);
or U2912 (N_2912,N_1507,N_1879);
nand U2913 (N_2913,N_1405,N_1924);
nand U2914 (N_2914,N_1283,N_1004);
or U2915 (N_2915,N_1059,N_1150);
nand U2916 (N_2916,N_1816,N_1451);
xor U2917 (N_2917,N_1720,N_1937);
or U2918 (N_2918,N_1244,N_1281);
nor U2919 (N_2919,N_1449,N_1499);
and U2920 (N_2920,N_1940,N_1692);
and U2921 (N_2921,N_1427,N_1743);
or U2922 (N_2922,N_1236,N_1416);
and U2923 (N_2923,N_1082,N_1987);
nand U2924 (N_2924,N_1439,N_1030);
nor U2925 (N_2925,N_1159,N_1598);
or U2926 (N_2926,N_1939,N_1713);
nor U2927 (N_2927,N_1458,N_1361);
nor U2928 (N_2928,N_1190,N_1450);
or U2929 (N_2929,N_1087,N_1605);
or U2930 (N_2930,N_1658,N_1666);
or U2931 (N_2931,N_1291,N_1265);
nand U2932 (N_2932,N_1726,N_1531);
or U2933 (N_2933,N_1464,N_1278);
or U2934 (N_2934,N_1780,N_1670);
and U2935 (N_2935,N_1168,N_1852);
nand U2936 (N_2936,N_1004,N_1192);
and U2937 (N_2937,N_1732,N_1988);
nor U2938 (N_2938,N_1089,N_1734);
nor U2939 (N_2939,N_1922,N_1431);
nand U2940 (N_2940,N_1613,N_1798);
nor U2941 (N_2941,N_1456,N_1977);
nand U2942 (N_2942,N_1524,N_1910);
nand U2943 (N_2943,N_1439,N_1052);
or U2944 (N_2944,N_1225,N_1064);
nor U2945 (N_2945,N_1725,N_1756);
and U2946 (N_2946,N_1234,N_1031);
nand U2947 (N_2947,N_1868,N_1325);
nand U2948 (N_2948,N_1677,N_1504);
nand U2949 (N_2949,N_1023,N_1506);
and U2950 (N_2950,N_1162,N_1863);
and U2951 (N_2951,N_1755,N_1435);
and U2952 (N_2952,N_1151,N_1910);
or U2953 (N_2953,N_1529,N_1212);
nand U2954 (N_2954,N_1663,N_1048);
nand U2955 (N_2955,N_1839,N_1092);
nand U2956 (N_2956,N_1842,N_1123);
and U2957 (N_2957,N_1840,N_1738);
nor U2958 (N_2958,N_1345,N_1691);
or U2959 (N_2959,N_1169,N_1639);
nand U2960 (N_2960,N_1350,N_1087);
or U2961 (N_2961,N_1568,N_1925);
nor U2962 (N_2962,N_1018,N_1200);
and U2963 (N_2963,N_1544,N_1075);
nor U2964 (N_2964,N_1653,N_1467);
and U2965 (N_2965,N_1176,N_1638);
nand U2966 (N_2966,N_1891,N_1882);
and U2967 (N_2967,N_1397,N_1639);
or U2968 (N_2968,N_1639,N_1926);
or U2969 (N_2969,N_1305,N_1830);
nor U2970 (N_2970,N_1325,N_1330);
nand U2971 (N_2971,N_1335,N_1471);
nor U2972 (N_2972,N_1642,N_1025);
nand U2973 (N_2973,N_1012,N_1794);
or U2974 (N_2974,N_1828,N_1394);
and U2975 (N_2975,N_1485,N_1383);
nand U2976 (N_2976,N_1403,N_1632);
and U2977 (N_2977,N_1036,N_1363);
and U2978 (N_2978,N_1501,N_1899);
or U2979 (N_2979,N_1029,N_1537);
or U2980 (N_2980,N_1788,N_1057);
or U2981 (N_2981,N_1342,N_1963);
nor U2982 (N_2982,N_1545,N_1082);
or U2983 (N_2983,N_1551,N_1841);
nand U2984 (N_2984,N_1115,N_1775);
nand U2985 (N_2985,N_1161,N_1170);
nor U2986 (N_2986,N_1163,N_1690);
and U2987 (N_2987,N_1236,N_1104);
nand U2988 (N_2988,N_1298,N_1476);
and U2989 (N_2989,N_1148,N_1441);
or U2990 (N_2990,N_1370,N_1898);
or U2991 (N_2991,N_1877,N_1426);
and U2992 (N_2992,N_1139,N_1113);
or U2993 (N_2993,N_1205,N_1343);
nand U2994 (N_2994,N_1258,N_1848);
and U2995 (N_2995,N_1105,N_1780);
and U2996 (N_2996,N_1013,N_1207);
nand U2997 (N_2997,N_1439,N_1313);
nand U2998 (N_2998,N_1988,N_1557);
nand U2999 (N_2999,N_1550,N_1306);
nand U3000 (N_3000,N_2904,N_2940);
nand U3001 (N_3001,N_2095,N_2503);
nand U3002 (N_3002,N_2121,N_2052);
nand U3003 (N_3003,N_2082,N_2346);
nor U3004 (N_3004,N_2388,N_2411);
nor U3005 (N_3005,N_2677,N_2282);
nor U3006 (N_3006,N_2421,N_2092);
nand U3007 (N_3007,N_2394,N_2636);
nor U3008 (N_3008,N_2109,N_2047);
or U3009 (N_3009,N_2275,N_2387);
nand U3010 (N_3010,N_2296,N_2350);
xor U3011 (N_3011,N_2139,N_2571);
nand U3012 (N_3012,N_2753,N_2457);
nor U3013 (N_3013,N_2563,N_2236);
and U3014 (N_3014,N_2818,N_2923);
and U3015 (N_3015,N_2698,N_2134);
and U3016 (N_3016,N_2098,N_2631);
or U3017 (N_3017,N_2982,N_2230);
nand U3018 (N_3018,N_2008,N_2269);
and U3019 (N_3019,N_2124,N_2155);
nor U3020 (N_3020,N_2397,N_2413);
or U3021 (N_3021,N_2381,N_2693);
and U3022 (N_3022,N_2347,N_2308);
nor U3023 (N_3023,N_2638,N_2110);
nor U3024 (N_3024,N_2502,N_2432);
and U3025 (N_3025,N_2256,N_2614);
nand U3026 (N_3026,N_2848,N_2748);
nand U3027 (N_3027,N_2015,N_2755);
or U3028 (N_3028,N_2557,N_2500);
or U3029 (N_3029,N_2592,N_2918);
or U3030 (N_3030,N_2512,N_2891);
or U3031 (N_3031,N_2332,N_2646);
nand U3032 (N_3032,N_2882,N_2993);
and U3033 (N_3033,N_2665,N_2348);
nor U3034 (N_3034,N_2170,N_2775);
or U3035 (N_3035,N_2299,N_2661);
and U3036 (N_3036,N_2896,N_2301);
or U3037 (N_3037,N_2611,N_2291);
or U3038 (N_3038,N_2055,N_2228);
nor U3039 (N_3039,N_2612,N_2135);
or U3040 (N_3040,N_2252,N_2177);
and U3041 (N_3041,N_2171,N_2142);
and U3042 (N_3042,N_2566,N_2054);
and U3043 (N_3043,N_2875,N_2710);
and U3044 (N_3044,N_2342,N_2766);
or U3045 (N_3045,N_2009,N_2034);
and U3046 (N_3046,N_2371,N_2527);
and U3047 (N_3047,N_2311,N_2203);
nand U3048 (N_3048,N_2810,N_2328);
and U3049 (N_3049,N_2695,N_2272);
nand U3050 (N_3050,N_2427,N_2556);
and U3051 (N_3051,N_2706,N_2470);
and U3052 (N_3052,N_2339,N_2842);
nor U3053 (N_3053,N_2048,N_2090);
nor U3054 (N_3054,N_2147,N_2788);
nor U3055 (N_3055,N_2243,N_2696);
or U3056 (N_3056,N_2863,N_2830);
nand U3057 (N_3057,N_2231,N_2670);
nand U3058 (N_3058,N_2360,N_2913);
or U3059 (N_3059,N_2319,N_2772);
and U3060 (N_3060,N_2321,N_2042);
nor U3061 (N_3061,N_2154,N_2501);
nor U3062 (N_3062,N_2579,N_2317);
and U3063 (N_3063,N_2545,N_2096);
or U3064 (N_3064,N_2949,N_2261);
nand U3065 (N_3065,N_2425,N_2865);
or U3066 (N_3066,N_2543,N_2149);
nor U3067 (N_3067,N_2552,N_2439);
nand U3068 (N_3068,N_2232,N_2163);
and U3069 (N_3069,N_2524,N_2444);
nor U3070 (N_3070,N_2167,N_2589);
nor U3071 (N_3071,N_2708,N_2724);
xnor U3072 (N_3072,N_2063,N_2590);
nand U3073 (N_3073,N_2811,N_2481);
nor U3074 (N_3074,N_2138,N_2086);
nor U3075 (N_3075,N_2365,N_2870);
nor U3076 (N_3076,N_2518,N_2062);
or U3077 (N_3077,N_2634,N_2085);
or U3078 (N_3078,N_2723,N_2547);
nor U3079 (N_3079,N_2645,N_2560);
or U3080 (N_3080,N_2003,N_2403);
or U3081 (N_3081,N_2655,N_2594);
or U3082 (N_3082,N_2534,N_2866);
nor U3083 (N_3083,N_2292,N_2101);
nor U3084 (N_3084,N_2986,N_2416);
nand U3085 (N_3085,N_2714,N_2654);
nor U3086 (N_3086,N_2314,N_2441);
and U3087 (N_3087,N_2483,N_2424);
nor U3088 (N_3088,N_2701,N_2069);
nor U3089 (N_3089,N_2012,N_2805);
nand U3090 (N_3090,N_2739,N_2129);
or U3091 (N_3091,N_2550,N_2331);
or U3092 (N_3092,N_2697,N_2390);
or U3093 (N_3093,N_2595,N_2694);
nor U3094 (N_3094,N_2798,N_2375);
nor U3095 (N_3095,N_2643,N_2037);
or U3096 (N_3096,N_2983,N_2359);
nand U3097 (N_3097,N_2943,N_2017);
nor U3098 (N_3098,N_2326,N_2757);
nor U3099 (N_3099,N_2843,N_2353);
or U3100 (N_3100,N_2059,N_2599);
nand U3101 (N_3101,N_2660,N_2561);
nor U3102 (N_3102,N_2504,N_2253);
nand U3103 (N_3103,N_2463,N_2459);
nor U3104 (N_3104,N_2649,N_2911);
or U3105 (N_3105,N_2861,N_2893);
nor U3106 (N_3106,N_2068,N_2316);
nand U3107 (N_3107,N_2782,N_2202);
and U3108 (N_3108,N_2945,N_2125);
nor U3109 (N_3109,N_2356,N_2516);
nand U3110 (N_3110,N_2367,N_2482);
and U3111 (N_3111,N_2934,N_2370);
xor U3112 (N_3112,N_2408,N_2309);
or U3113 (N_3113,N_2779,N_2405);
nand U3114 (N_3114,N_2107,N_2574);
or U3115 (N_3115,N_2627,N_2146);
or U3116 (N_3116,N_2270,N_2066);
nor U3117 (N_3117,N_2114,N_2762);
and U3118 (N_3118,N_2450,N_2617);
and U3119 (N_3119,N_2813,N_2192);
nor U3120 (N_3120,N_2156,N_2447);
and U3121 (N_3121,N_2443,N_2931);
nor U3122 (N_3122,N_2219,N_2731);
or U3123 (N_3123,N_2860,N_2173);
and U3124 (N_3124,N_2455,N_2250);
nor U3125 (N_3125,N_2525,N_2473);
nand U3126 (N_3126,N_2554,N_2300);
nor U3127 (N_3127,N_2531,N_2776);
nor U3128 (N_3128,N_2071,N_2277);
nor U3129 (N_3129,N_2548,N_2998);
nand U3130 (N_3130,N_2879,N_2333);
xnor U3131 (N_3131,N_2143,N_2808);
and U3132 (N_3132,N_2832,N_2358);
nor U3133 (N_3133,N_2136,N_2528);
and U3134 (N_3134,N_2814,N_2486);
or U3135 (N_3135,N_2168,N_2799);
or U3136 (N_3136,N_2732,N_2214);
or U3137 (N_3137,N_2248,N_2764);
and U3138 (N_3138,N_2389,N_2623);
and U3139 (N_3139,N_2480,N_2921);
nor U3140 (N_3140,N_2437,N_2064);
or U3141 (N_3141,N_2704,N_2587);
xor U3142 (N_3142,N_2364,N_2099);
or U3143 (N_3143,N_2841,N_2719);
and U3144 (N_3144,N_2188,N_2662);
and U3145 (N_3145,N_2700,N_2488);
and U3146 (N_3146,N_2276,N_2368);
and U3147 (N_3147,N_2576,N_2965);
and U3148 (N_3148,N_2158,N_2336);
and U3149 (N_3149,N_2351,N_2613);
nor U3150 (N_3150,N_2707,N_2602);
nor U3151 (N_3151,N_2692,N_2385);
and U3152 (N_3152,N_2251,N_2958);
nand U3153 (N_3153,N_2744,N_2106);
nand U3154 (N_3154,N_2712,N_2559);
or U3155 (N_3155,N_2991,N_2892);
nand U3156 (N_3156,N_2000,N_2033);
and U3157 (N_3157,N_2874,N_2987);
nor U3158 (N_3158,N_2409,N_2831);
nand U3159 (N_3159,N_2908,N_2324);
or U3160 (N_3160,N_2877,N_2274);
nor U3161 (N_3161,N_2827,N_2304);
nor U3162 (N_3162,N_2323,N_2608);
or U3163 (N_3163,N_2951,N_2476);
nor U3164 (N_3164,N_2784,N_2349);
or U3165 (N_3165,N_2567,N_2377);
and U3166 (N_3166,N_2461,N_2315);
and U3167 (N_3167,N_2889,N_2189);
and U3168 (N_3168,N_2379,N_2615);
xor U3169 (N_3169,N_2376,N_2220);
nor U3170 (N_3170,N_2812,N_2175);
or U3171 (N_3171,N_2577,N_2216);
and U3172 (N_3172,N_2433,N_2094);
nor U3173 (N_3173,N_2920,N_2869);
nand U3174 (N_3174,N_2971,N_2996);
nand U3175 (N_3175,N_2999,N_2051);
and U3176 (N_3176,N_2758,N_2399);
and U3177 (N_3177,N_2873,N_2148);
xnor U3178 (N_3178,N_2065,N_2060);
or U3179 (N_3179,N_2759,N_2464);
or U3180 (N_3180,N_2398,N_2499);
nor U3181 (N_3181,N_2727,N_2484);
nand U3182 (N_3182,N_2607,N_2935);
nor U3183 (N_3183,N_2887,N_2227);
and U3184 (N_3184,N_2910,N_2440);
or U3185 (N_3185,N_2997,N_2372);
and U3186 (N_3186,N_2020,N_2740);
and U3187 (N_3187,N_2043,N_2729);
nand U3188 (N_3188,N_2074,N_2010);
nand U3189 (N_3189,N_2344,N_2329);
nor U3190 (N_3190,N_2485,N_2498);
nand U3191 (N_3191,N_2026,N_2742);
or U3192 (N_3192,N_2838,N_2479);
nand U3193 (N_3193,N_2373,N_2960);
nor U3194 (N_3194,N_2237,N_2294);
nand U3195 (N_3195,N_2036,N_2988);
and U3196 (N_3196,N_2747,N_2083);
or U3197 (N_3197,N_2994,N_2325);
nand U3198 (N_3198,N_2112,N_2180);
and U3199 (N_3199,N_2800,N_2307);
nand U3200 (N_3200,N_2947,N_2787);
and U3201 (N_3201,N_2472,N_2972);
nand U3202 (N_3202,N_2756,N_2950);
or U3203 (N_3203,N_2711,N_2268);
nor U3204 (N_3204,N_2229,N_2050);
and U3205 (N_3205,N_2363,N_2666);
nor U3206 (N_3206,N_2298,N_2293);
or U3207 (N_3207,N_2337,N_2593);
nand U3208 (N_3208,N_2881,N_2953);
and U3209 (N_3209,N_2496,N_2507);
and U3210 (N_3210,N_2070,N_2583);
nor U3211 (N_3211,N_2458,N_2046);
or U3212 (N_3212,N_2538,N_2819);
nor U3213 (N_3213,N_2895,N_2040);
and U3214 (N_3214,N_2233,N_2414);
and U3215 (N_3215,N_2743,N_2391);
nor U3216 (N_3216,N_2213,N_2061);
or U3217 (N_3217,N_2690,N_2658);
and U3218 (N_3218,N_2916,N_2763);
nor U3219 (N_3219,N_2912,N_2151);
nor U3220 (N_3220,N_2285,N_2928);
and U3221 (N_3221,N_2119,N_2508);
nand U3222 (N_3222,N_2572,N_2540);
nand U3223 (N_3223,N_2616,N_2018);
and U3224 (N_3224,N_2944,N_2392);
nor U3225 (N_3225,N_2852,N_2839);
nor U3226 (N_3226,N_2117,N_2312);
or U3227 (N_3227,N_2678,N_2211);
or U3228 (N_3228,N_2871,N_2513);
nor U3229 (N_3229,N_2834,N_2164);
nand U3230 (N_3230,N_2938,N_2279);
nor U3231 (N_3231,N_2878,N_2862);
nand U3232 (N_3232,N_2822,N_2932);
and U3233 (N_3233,N_2954,N_2386);
and U3234 (N_3234,N_2975,N_2976);
or U3235 (N_3235,N_2647,N_2137);
or U3236 (N_3236,N_2773,N_2720);
nor U3237 (N_3237,N_2526,N_2019);
nand U3238 (N_3238,N_2338,N_2990);
nor U3239 (N_3239,N_2777,N_2187);
and U3240 (N_3240,N_2562,N_2930);
xor U3241 (N_3241,N_2880,N_2087);
nor U3242 (N_3242,N_2007,N_2610);
or U3243 (N_3243,N_2014,N_2045);
and U3244 (N_3244,N_2474,N_2900);
nor U3245 (N_3245,N_2400,N_2471);
and U3246 (N_3246,N_2145,N_2283);
xor U3247 (N_3247,N_2166,N_2844);
nor U3248 (N_3248,N_2846,N_2956);
or U3249 (N_3249,N_2401,N_2637);
nor U3250 (N_3250,N_2919,N_2209);
nand U3251 (N_3251,N_2258,N_2505);
nand U3252 (N_3252,N_2084,N_2254);
and U3253 (N_3253,N_2977,N_2395);
nor U3254 (N_3254,N_2575,N_2172);
or U3255 (N_3255,N_2530,N_2366);
nor U3256 (N_3256,N_2717,N_2334);
nand U3257 (N_3257,N_2415,N_2939);
and U3258 (N_3258,N_2741,N_2025);
or U3259 (N_3259,N_2687,N_2453);
nand U3260 (N_3260,N_2907,N_2238);
nor U3261 (N_3261,N_2257,N_2023);
nor U3262 (N_3262,N_2546,N_2406);
nand U3263 (N_3263,N_2454,N_2041);
or U3264 (N_3264,N_2361,N_2186);
and U3265 (N_3265,N_2520,N_2352);
nand U3266 (N_3266,N_2190,N_2621);
and U3267 (N_3267,N_2725,N_2718);
or U3268 (N_3268,N_2224,N_2417);
and U3269 (N_3269,N_2511,N_2709);
nor U3270 (N_3270,N_2162,N_2769);
or U3271 (N_3271,N_2667,N_2259);
nor U3272 (N_3272,N_2533,N_2436);
and U3273 (N_3273,N_2672,N_2849);
nand U3274 (N_3274,N_2628,N_2289);
and U3275 (N_3275,N_2521,N_2952);
nor U3276 (N_3276,N_2449,N_2097);
nand U3277 (N_3277,N_2419,N_2028);
or U3278 (N_3278,N_2102,N_2651);
nand U3279 (N_3279,N_2854,N_2239);
and U3280 (N_3280,N_2885,N_2970);
and U3281 (N_3281,N_2320,N_2768);
and U3282 (N_3282,N_2031,N_2407);
nor U3283 (N_3283,N_2491,N_2100);
and U3284 (N_3284,N_2210,N_2240);
nor U3285 (N_3285,N_2801,N_2824);
or U3286 (N_3286,N_2490,N_2245);
or U3287 (N_3287,N_2797,N_2752);
nor U3288 (N_3288,N_2657,N_2495);
and U3289 (N_3289,N_2206,N_2876);
nand U3290 (N_3290,N_2941,N_2806);
nand U3291 (N_3291,N_2434,N_2013);
xnor U3292 (N_3292,N_2089,N_2199);
or U3293 (N_3293,N_2288,N_2836);
nand U3294 (N_3294,N_2573,N_2194);
nor U3295 (N_3295,N_2789,N_2722);
and U3296 (N_3296,N_2185,N_2430);
nand U3297 (N_3297,N_2738,N_2807);
or U3298 (N_3298,N_2601,N_2073);
nand U3299 (N_3299,N_2635,N_2985);
nor U3300 (N_3300,N_2780,N_2536);
and U3301 (N_3301,N_2157,N_2578);
or U3302 (N_3302,N_2625,N_2835);
or U3303 (N_3303,N_2184,N_2837);
or U3304 (N_3304,N_2855,N_2626);
nand U3305 (N_3305,N_2044,N_2335);
and U3306 (N_3306,N_2297,N_2629);
nand U3307 (N_3307,N_2979,N_2925);
nor U3308 (N_3308,N_2630,N_2584);
nand U3309 (N_3309,N_2933,N_2760);
nor U3310 (N_3310,N_2021,N_2195);
and U3311 (N_3311,N_2541,N_2242);
or U3312 (N_3312,N_2851,N_2144);
and U3313 (N_3313,N_2280,N_2604);
and U3314 (N_3314,N_2682,N_2624);
and U3315 (N_3315,N_2746,N_2641);
or U3316 (N_3316,N_2632,N_2341);
nand U3317 (N_3317,N_2244,N_2153);
nor U3318 (N_3318,N_2537,N_2120);
nand U3319 (N_3319,N_2105,N_2581);
and U3320 (N_3320,N_2897,N_2978);
and U3321 (N_3321,N_2005,N_2123);
nor U3322 (N_3322,N_2803,N_2596);
and U3323 (N_3323,N_2204,N_2703);
nor U3324 (N_3324,N_2428,N_2475);
nand U3325 (N_3325,N_2150,N_2856);
nand U3326 (N_3326,N_2936,N_2633);
nor U3327 (N_3327,N_2659,N_2794);
nor U3328 (N_3328,N_2462,N_2404);
nand U3329 (N_3329,N_2072,N_2116);
nor U3330 (N_3330,N_2809,N_2817);
and U3331 (N_3331,N_2038,N_2795);
and U3332 (N_3332,N_2273,N_2418);
or U3333 (N_3333,N_2039,N_2796);
nand U3334 (N_3334,N_2745,N_2715);
nor U3335 (N_3335,N_2265,N_2858);
nand U3336 (N_3336,N_2681,N_2234);
and U3337 (N_3337,N_2909,N_2489);
or U3338 (N_3338,N_2825,N_2223);
or U3339 (N_3339,N_2529,N_2384);
nand U3340 (N_3340,N_2644,N_2620);
nand U3341 (N_3341,N_2451,N_2362);
nor U3342 (N_3342,N_2679,N_2104);
or U3343 (N_3343,N_2152,N_2791);
and U3344 (N_3344,N_2140,N_2872);
and U3345 (N_3345,N_2606,N_2494);
nor U3346 (N_3346,N_2733,N_2688);
and U3347 (N_3347,N_2542,N_2973);
nor U3348 (N_3348,N_2588,N_2605);
xnor U3349 (N_3349,N_2262,N_2699);
or U3350 (N_3350,N_2968,N_2544);
nor U3351 (N_3351,N_2580,N_2663);
and U3352 (N_3352,N_2517,N_2049);
or U3353 (N_3353,N_2355,N_2751);
and U3354 (N_3354,N_2078,N_2815);
nor U3355 (N_3355,N_2128,N_2108);
nor U3356 (N_3356,N_2278,N_2281);
nor U3357 (N_3357,N_2313,N_2726);
or U3358 (N_3358,N_2438,N_2549);
and U3359 (N_3359,N_2514,N_2989);
nand U3360 (N_3360,N_2035,N_2183);
and U3361 (N_3361,N_2565,N_2422);
and U3362 (N_3362,N_2284,N_2555);
nor U3363 (N_3363,N_2465,N_2761);
nand U3364 (N_3364,N_2380,N_2598);
and U3365 (N_3365,N_2249,N_2922);
and U3366 (N_3366,N_2287,N_2929);
nor U3367 (N_3367,N_2961,N_2027);
and U3368 (N_3368,N_2225,N_2266);
and U3369 (N_3369,N_2196,N_2734);
or U3370 (N_3370,N_2169,N_2469);
and U3371 (N_3371,N_2429,N_2826);
nor U3372 (N_3372,N_2917,N_2016);
nor U3373 (N_3373,N_2067,N_2467);
or U3374 (N_3374,N_2650,N_2222);
nand U3375 (N_3375,N_2212,N_2515);
nor U3376 (N_3376,N_2191,N_2792);
or U3377 (N_3377,N_2648,N_2735);
nand U3378 (N_3378,N_2609,N_2915);
nor U3379 (N_3379,N_2691,N_2081);
and U3380 (N_3380,N_2295,N_2992);
nor U3381 (N_3381,N_2159,N_2619);
or U3382 (N_3382,N_2032,N_2535);
nor U3383 (N_3383,N_2448,N_2318);
nor U3384 (N_3384,N_2378,N_2603);
or U3385 (N_3385,N_2783,N_2959);
or U3386 (N_3386,N_2263,N_2948);
nand U3387 (N_3387,N_2080,N_2200);
nor U3388 (N_3388,N_2509,N_2197);
nor U3389 (N_3389,N_2570,N_2964);
and U3390 (N_3390,N_2410,N_2497);
or U3391 (N_3391,N_2618,N_2771);
nand U3392 (N_3392,N_2804,N_2899);
or U3393 (N_3393,N_2886,N_2460);
nand U3394 (N_3394,N_2456,N_2235);
nor U3395 (N_3395,N_2271,N_2901);
nand U3396 (N_3396,N_2522,N_2664);
and U3397 (N_3397,N_2888,N_2493);
and U3398 (N_3398,N_2053,N_2774);
nor U3399 (N_3399,N_2383,N_2226);
or U3400 (N_3400,N_2656,N_2974);
or U3401 (N_3401,N_2354,N_2426);
nand U3402 (N_3402,N_2510,N_2984);
nor U3403 (N_3403,N_2382,N_2093);
nor U3404 (N_3404,N_2927,N_2668);
nor U3405 (N_3405,N_2115,N_2267);
nor U3406 (N_3406,N_2597,N_2689);
and U3407 (N_3407,N_2770,N_2942);
nand U3408 (N_3408,N_2591,N_2765);
or U3409 (N_3409,N_2906,N_2981);
and U3410 (N_3410,N_2182,N_2305);
and U3411 (N_3411,N_2345,N_2946);
nand U3412 (N_3412,N_2357,N_2058);
nor U3413 (N_3413,N_2290,N_2006);
nor U3414 (N_3414,N_2088,N_2539);
and U3415 (N_3415,N_2452,N_2445);
nor U3416 (N_3416,N_2215,N_2030);
and U3417 (N_3417,N_2178,N_2091);
or U3418 (N_3418,N_2868,N_2523);
nor U3419 (N_3419,N_2310,N_2853);
nor U3420 (N_3420,N_2002,N_2569);
and U3421 (N_3421,N_2676,N_2785);
nor U3422 (N_3422,N_2850,N_2374);
nand U3423 (N_3423,N_2737,N_2011);
and U3424 (N_3424,N_2343,N_2322);
nor U3425 (N_3425,N_2466,N_2793);
xnor U3426 (N_3426,N_2260,N_2716);
or U3427 (N_3427,N_2181,N_2639);
nand U3428 (N_3428,N_2702,N_2412);
and U3429 (N_3429,N_2207,N_2160);
and U3430 (N_3430,N_2963,N_2369);
and U3431 (N_3431,N_2564,N_2840);
and U3432 (N_3432,N_2506,N_2829);
nand U3433 (N_3433,N_2705,N_2478);
nand U3434 (N_3434,N_2179,N_2680);
nor U3435 (N_3435,N_2221,N_2778);
or U3436 (N_3436,N_2898,N_2113);
nor U3437 (N_3437,N_2247,N_2492);
nand U3438 (N_3438,N_2845,N_2029);
nand U3439 (N_3439,N_2859,N_2217);
and U3440 (N_3440,N_2675,N_2781);
nand U3441 (N_3441,N_2582,N_2642);
nor U3442 (N_3442,N_2786,N_2302);
nand U3443 (N_3443,N_2132,N_2057);
and U3444 (N_3444,N_2161,N_2955);
nand U3445 (N_3445,N_2193,N_2914);
and U3446 (N_3446,N_2966,N_2721);
or U3447 (N_3447,N_2468,N_2937);
nor U3448 (N_3448,N_2980,N_2568);
and U3449 (N_3449,N_2133,N_2477);
and U3450 (N_3450,N_2396,N_2327);
and U3451 (N_3451,N_2558,N_2022);
or U3452 (N_3452,N_2201,N_2924);
xor U3453 (N_3453,N_2894,N_2174);
nor U3454 (N_3454,N_2176,N_2131);
nand U3455 (N_3455,N_2111,N_2683);
nor U3456 (N_3456,N_2103,N_2884);
nor U3457 (N_3457,N_2001,N_2754);
and U3458 (N_3458,N_2435,N_2820);
nand U3459 (N_3459,N_2141,N_2246);
nand U3460 (N_3460,N_2004,N_2079);
and U3461 (N_3461,N_2790,N_2995);
or U3462 (N_3462,N_2867,N_2487);
or U3463 (N_3463,N_2431,N_2024);
nor U3464 (N_3464,N_2883,N_2056);
and U3465 (N_3465,N_2864,N_2340);
or U3466 (N_3466,N_2926,N_2306);
and U3467 (N_3467,N_2713,N_2669);
nand U3468 (N_3468,N_2205,N_2640);
nor U3469 (N_3469,N_2905,N_2749);
nor U3470 (N_3470,N_2551,N_2802);
nand U3471 (N_3471,N_2736,N_2728);
nor U3472 (N_3472,N_2816,N_2402);
or U3473 (N_3473,N_2420,N_2730);
or U3474 (N_3474,N_2902,N_2622);
or U3475 (N_3475,N_2586,N_2330);
nor U3476 (N_3476,N_2674,N_2532);
and U3477 (N_3477,N_2821,N_2122);
nor U3478 (N_3478,N_2903,N_2553);
or U3479 (N_3479,N_2165,N_2673);
nor U3480 (N_3480,N_2118,N_2198);
nor U3481 (N_3481,N_2218,N_2303);
and U3482 (N_3482,N_2890,N_2519);
nand U3483 (N_3483,N_2255,N_2833);
or U3484 (N_3484,N_2208,N_2446);
nor U3485 (N_3485,N_2442,N_2967);
and U3486 (N_3486,N_2857,N_2653);
and U3487 (N_3487,N_2685,N_2393);
or U3488 (N_3488,N_2684,N_2962);
nand U3489 (N_3489,N_2127,N_2130);
nor U3490 (N_3490,N_2241,N_2585);
or U3491 (N_3491,N_2671,N_2075);
nor U3492 (N_3492,N_2652,N_2077);
and U3493 (N_3493,N_2076,N_2969);
and U3494 (N_3494,N_2847,N_2600);
or U3495 (N_3495,N_2686,N_2767);
nor U3496 (N_3496,N_2828,N_2126);
or U3497 (N_3497,N_2423,N_2823);
and U3498 (N_3498,N_2264,N_2957);
nand U3499 (N_3499,N_2286,N_2750);
nand U3500 (N_3500,N_2706,N_2644);
and U3501 (N_3501,N_2129,N_2488);
nor U3502 (N_3502,N_2087,N_2610);
or U3503 (N_3503,N_2050,N_2297);
nor U3504 (N_3504,N_2544,N_2242);
or U3505 (N_3505,N_2189,N_2681);
nor U3506 (N_3506,N_2541,N_2503);
nand U3507 (N_3507,N_2932,N_2742);
or U3508 (N_3508,N_2544,N_2737);
nand U3509 (N_3509,N_2006,N_2057);
nor U3510 (N_3510,N_2863,N_2931);
nand U3511 (N_3511,N_2071,N_2466);
nand U3512 (N_3512,N_2275,N_2700);
or U3513 (N_3513,N_2375,N_2810);
and U3514 (N_3514,N_2978,N_2258);
nor U3515 (N_3515,N_2823,N_2903);
nand U3516 (N_3516,N_2980,N_2097);
nor U3517 (N_3517,N_2161,N_2295);
nor U3518 (N_3518,N_2214,N_2465);
or U3519 (N_3519,N_2450,N_2710);
and U3520 (N_3520,N_2956,N_2418);
nor U3521 (N_3521,N_2890,N_2821);
and U3522 (N_3522,N_2096,N_2696);
or U3523 (N_3523,N_2675,N_2125);
nor U3524 (N_3524,N_2198,N_2300);
nand U3525 (N_3525,N_2753,N_2399);
and U3526 (N_3526,N_2049,N_2627);
nand U3527 (N_3527,N_2449,N_2342);
nand U3528 (N_3528,N_2659,N_2382);
or U3529 (N_3529,N_2570,N_2870);
nor U3530 (N_3530,N_2173,N_2413);
and U3531 (N_3531,N_2880,N_2952);
nor U3532 (N_3532,N_2296,N_2683);
and U3533 (N_3533,N_2429,N_2338);
or U3534 (N_3534,N_2689,N_2066);
and U3535 (N_3535,N_2169,N_2050);
nand U3536 (N_3536,N_2416,N_2233);
and U3537 (N_3537,N_2422,N_2988);
nor U3538 (N_3538,N_2159,N_2529);
and U3539 (N_3539,N_2814,N_2454);
or U3540 (N_3540,N_2830,N_2531);
or U3541 (N_3541,N_2794,N_2780);
nand U3542 (N_3542,N_2721,N_2189);
and U3543 (N_3543,N_2852,N_2808);
or U3544 (N_3544,N_2107,N_2953);
or U3545 (N_3545,N_2050,N_2874);
or U3546 (N_3546,N_2568,N_2003);
nand U3547 (N_3547,N_2026,N_2031);
and U3548 (N_3548,N_2094,N_2981);
nor U3549 (N_3549,N_2182,N_2582);
nand U3550 (N_3550,N_2053,N_2766);
or U3551 (N_3551,N_2358,N_2496);
nor U3552 (N_3552,N_2904,N_2261);
and U3553 (N_3553,N_2820,N_2249);
nand U3554 (N_3554,N_2181,N_2224);
nor U3555 (N_3555,N_2867,N_2799);
and U3556 (N_3556,N_2065,N_2607);
nor U3557 (N_3557,N_2954,N_2817);
nand U3558 (N_3558,N_2583,N_2262);
nor U3559 (N_3559,N_2358,N_2236);
or U3560 (N_3560,N_2651,N_2248);
nor U3561 (N_3561,N_2203,N_2297);
nor U3562 (N_3562,N_2651,N_2858);
and U3563 (N_3563,N_2471,N_2859);
nand U3564 (N_3564,N_2374,N_2484);
or U3565 (N_3565,N_2159,N_2616);
xnor U3566 (N_3566,N_2660,N_2664);
nand U3567 (N_3567,N_2381,N_2913);
or U3568 (N_3568,N_2497,N_2191);
and U3569 (N_3569,N_2735,N_2912);
nand U3570 (N_3570,N_2642,N_2058);
nand U3571 (N_3571,N_2248,N_2868);
nor U3572 (N_3572,N_2669,N_2083);
nor U3573 (N_3573,N_2854,N_2866);
or U3574 (N_3574,N_2503,N_2416);
and U3575 (N_3575,N_2173,N_2358);
or U3576 (N_3576,N_2344,N_2245);
nor U3577 (N_3577,N_2632,N_2750);
nand U3578 (N_3578,N_2431,N_2103);
or U3579 (N_3579,N_2871,N_2510);
or U3580 (N_3580,N_2406,N_2563);
nand U3581 (N_3581,N_2916,N_2038);
and U3582 (N_3582,N_2884,N_2343);
or U3583 (N_3583,N_2439,N_2851);
and U3584 (N_3584,N_2574,N_2544);
and U3585 (N_3585,N_2744,N_2559);
or U3586 (N_3586,N_2281,N_2448);
or U3587 (N_3587,N_2225,N_2766);
nand U3588 (N_3588,N_2534,N_2379);
and U3589 (N_3589,N_2794,N_2247);
nand U3590 (N_3590,N_2531,N_2746);
nand U3591 (N_3591,N_2086,N_2889);
nand U3592 (N_3592,N_2645,N_2227);
nor U3593 (N_3593,N_2650,N_2692);
nor U3594 (N_3594,N_2686,N_2604);
and U3595 (N_3595,N_2925,N_2016);
or U3596 (N_3596,N_2655,N_2369);
nand U3597 (N_3597,N_2103,N_2368);
nand U3598 (N_3598,N_2500,N_2492);
or U3599 (N_3599,N_2193,N_2017);
nand U3600 (N_3600,N_2913,N_2395);
nand U3601 (N_3601,N_2631,N_2517);
and U3602 (N_3602,N_2462,N_2626);
nand U3603 (N_3603,N_2590,N_2408);
nand U3604 (N_3604,N_2538,N_2074);
or U3605 (N_3605,N_2194,N_2941);
nand U3606 (N_3606,N_2446,N_2928);
nand U3607 (N_3607,N_2404,N_2203);
xor U3608 (N_3608,N_2515,N_2758);
nor U3609 (N_3609,N_2333,N_2918);
or U3610 (N_3610,N_2630,N_2680);
or U3611 (N_3611,N_2845,N_2054);
or U3612 (N_3612,N_2057,N_2044);
xor U3613 (N_3613,N_2766,N_2612);
nor U3614 (N_3614,N_2590,N_2076);
or U3615 (N_3615,N_2776,N_2208);
nor U3616 (N_3616,N_2089,N_2355);
or U3617 (N_3617,N_2275,N_2670);
or U3618 (N_3618,N_2883,N_2769);
and U3619 (N_3619,N_2330,N_2409);
nor U3620 (N_3620,N_2196,N_2004);
and U3621 (N_3621,N_2176,N_2557);
nand U3622 (N_3622,N_2535,N_2995);
nor U3623 (N_3623,N_2354,N_2841);
or U3624 (N_3624,N_2569,N_2447);
nor U3625 (N_3625,N_2130,N_2013);
nor U3626 (N_3626,N_2254,N_2202);
nor U3627 (N_3627,N_2480,N_2696);
nand U3628 (N_3628,N_2227,N_2046);
and U3629 (N_3629,N_2439,N_2767);
nor U3630 (N_3630,N_2564,N_2422);
and U3631 (N_3631,N_2349,N_2646);
nor U3632 (N_3632,N_2310,N_2037);
and U3633 (N_3633,N_2593,N_2559);
and U3634 (N_3634,N_2634,N_2683);
and U3635 (N_3635,N_2087,N_2881);
and U3636 (N_3636,N_2062,N_2348);
or U3637 (N_3637,N_2225,N_2840);
nand U3638 (N_3638,N_2863,N_2606);
nand U3639 (N_3639,N_2677,N_2735);
or U3640 (N_3640,N_2356,N_2435);
nor U3641 (N_3641,N_2187,N_2472);
nor U3642 (N_3642,N_2587,N_2532);
nor U3643 (N_3643,N_2540,N_2462);
nor U3644 (N_3644,N_2698,N_2843);
and U3645 (N_3645,N_2838,N_2770);
or U3646 (N_3646,N_2161,N_2568);
and U3647 (N_3647,N_2702,N_2700);
nor U3648 (N_3648,N_2550,N_2274);
nor U3649 (N_3649,N_2114,N_2319);
nor U3650 (N_3650,N_2863,N_2416);
nor U3651 (N_3651,N_2962,N_2785);
or U3652 (N_3652,N_2064,N_2119);
nand U3653 (N_3653,N_2546,N_2393);
nor U3654 (N_3654,N_2662,N_2749);
and U3655 (N_3655,N_2816,N_2585);
and U3656 (N_3656,N_2936,N_2705);
or U3657 (N_3657,N_2942,N_2727);
or U3658 (N_3658,N_2673,N_2141);
nor U3659 (N_3659,N_2661,N_2317);
and U3660 (N_3660,N_2508,N_2604);
nor U3661 (N_3661,N_2541,N_2935);
nor U3662 (N_3662,N_2581,N_2418);
and U3663 (N_3663,N_2377,N_2497);
and U3664 (N_3664,N_2467,N_2405);
and U3665 (N_3665,N_2022,N_2625);
nand U3666 (N_3666,N_2961,N_2613);
nand U3667 (N_3667,N_2157,N_2391);
and U3668 (N_3668,N_2773,N_2767);
nand U3669 (N_3669,N_2898,N_2091);
nor U3670 (N_3670,N_2080,N_2166);
nor U3671 (N_3671,N_2307,N_2137);
nand U3672 (N_3672,N_2298,N_2848);
nor U3673 (N_3673,N_2127,N_2050);
or U3674 (N_3674,N_2251,N_2593);
and U3675 (N_3675,N_2298,N_2409);
and U3676 (N_3676,N_2810,N_2312);
or U3677 (N_3677,N_2557,N_2816);
nand U3678 (N_3678,N_2468,N_2601);
or U3679 (N_3679,N_2923,N_2429);
nand U3680 (N_3680,N_2420,N_2131);
and U3681 (N_3681,N_2156,N_2648);
or U3682 (N_3682,N_2568,N_2303);
and U3683 (N_3683,N_2980,N_2386);
or U3684 (N_3684,N_2053,N_2283);
nand U3685 (N_3685,N_2038,N_2970);
nand U3686 (N_3686,N_2542,N_2716);
or U3687 (N_3687,N_2269,N_2398);
and U3688 (N_3688,N_2667,N_2856);
or U3689 (N_3689,N_2337,N_2582);
and U3690 (N_3690,N_2013,N_2034);
nand U3691 (N_3691,N_2178,N_2946);
or U3692 (N_3692,N_2511,N_2440);
nor U3693 (N_3693,N_2538,N_2020);
and U3694 (N_3694,N_2577,N_2866);
or U3695 (N_3695,N_2673,N_2980);
nor U3696 (N_3696,N_2834,N_2410);
xnor U3697 (N_3697,N_2926,N_2153);
or U3698 (N_3698,N_2090,N_2102);
nand U3699 (N_3699,N_2701,N_2182);
or U3700 (N_3700,N_2608,N_2968);
nor U3701 (N_3701,N_2137,N_2474);
or U3702 (N_3702,N_2823,N_2379);
nand U3703 (N_3703,N_2248,N_2015);
and U3704 (N_3704,N_2980,N_2616);
and U3705 (N_3705,N_2655,N_2428);
or U3706 (N_3706,N_2452,N_2970);
and U3707 (N_3707,N_2664,N_2777);
or U3708 (N_3708,N_2265,N_2806);
or U3709 (N_3709,N_2830,N_2698);
nand U3710 (N_3710,N_2103,N_2418);
nor U3711 (N_3711,N_2827,N_2811);
and U3712 (N_3712,N_2803,N_2826);
and U3713 (N_3713,N_2295,N_2431);
nand U3714 (N_3714,N_2701,N_2801);
or U3715 (N_3715,N_2058,N_2112);
nand U3716 (N_3716,N_2953,N_2051);
nor U3717 (N_3717,N_2561,N_2725);
and U3718 (N_3718,N_2317,N_2261);
nor U3719 (N_3719,N_2500,N_2310);
nand U3720 (N_3720,N_2203,N_2195);
xor U3721 (N_3721,N_2386,N_2885);
nand U3722 (N_3722,N_2931,N_2100);
nor U3723 (N_3723,N_2458,N_2989);
and U3724 (N_3724,N_2235,N_2089);
and U3725 (N_3725,N_2368,N_2447);
nor U3726 (N_3726,N_2017,N_2916);
or U3727 (N_3727,N_2351,N_2425);
nand U3728 (N_3728,N_2160,N_2060);
nor U3729 (N_3729,N_2253,N_2319);
and U3730 (N_3730,N_2279,N_2935);
nand U3731 (N_3731,N_2752,N_2443);
and U3732 (N_3732,N_2726,N_2130);
nand U3733 (N_3733,N_2994,N_2004);
nor U3734 (N_3734,N_2015,N_2021);
nand U3735 (N_3735,N_2332,N_2441);
nand U3736 (N_3736,N_2514,N_2427);
nand U3737 (N_3737,N_2899,N_2388);
nor U3738 (N_3738,N_2591,N_2506);
and U3739 (N_3739,N_2768,N_2068);
nor U3740 (N_3740,N_2637,N_2004);
and U3741 (N_3741,N_2667,N_2467);
nor U3742 (N_3742,N_2765,N_2202);
nand U3743 (N_3743,N_2675,N_2250);
and U3744 (N_3744,N_2233,N_2515);
nand U3745 (N_3745,N_2412,N_2627);
and U3746 (N_3746,N_2403,N_2378);
or U3747 (N_3747,N_2971,N_2766);
or U3748 (N_3748,N_2136,N_2441);
nor U3749 (N_3749,N_2872,N_2469);
and U3750 (N_3750,N_2762,N_2812);
or U3751 (N_3751,N_2949,N_2568);
nor U3752 (N_3752,N_2296,N_2413);
nor U3753 (N_3753,N_2046,N_2992);
nand U3754 (N_3754,N_2881,N_2645);
nand U3755 (N_3755,N_2078,N_2296);
and U3756 (N_3756,N_2844,N_2948);
or U3757 (N_3757,N_2400,N_2810);
xor U3758 (N_3758,N_2607,N_2201);
nor U3759 (N_3759,N_2338,N_2445);
and U3760 (N_3760,N_2696,N_2024);
and U3761 (N_3761,N_2573,N_2710);
or U3762 (N_3762,N_2677,N_2800);
and U3763 (N_3763,N_2366,N_2740);
xor U3764 (N_3764,N_2661,N_2581);
or U3765 (N_3765,N_2801,N_2237);
nand U3766 (N_3766,N_2286,N_2740);
or U3767 (N_3767,N_2814,N_2181);
nand U3768 (N_3768,N_2067,N_2105);
and U3769 (N_3769,N_2161,N_2768);
or U3770 (N_3770,N_2972,N_2499);
nand U3771 (N_3771,N_2849,N_2736);
and U3772 (N_3772,N_2662,N_2224);
nor U3773 (N_3773,N_2692,N_2600);
or U3774 (N_3774,N_2144,N_2911);
and U3775 (N_3775,N_2811,N_2105);
nand U3776 (N_3776,N_2662,N_2650);
and U3777 (N_3777,N_2541,N_2211);
nor U3778 (N_3778,N_2248,N_2878);
and U3779 (N_3779,N_2295,N_2163);
nand U3780 (N_3780,N_2926,N_2760);
or U3781 (N_3781,N_2922,N_2311);
and U3782 (N_3782,N_2416,N_2529);
nor U3783 (N_3783,N_2991,N_2791);
and U3784 (N_3784,N_2170,N_2192);
and U3785 (N_3785,N_2428,N_2425);
nand U3786 (N_3786,N_2072,N_2753);
and U3787 (N_3787,N_2349,N_2053);
or U3788 (N_3788,N_2472,N_2777);
nor U3789 (N_3789,N_2164,N_2490);
nand U3790 (N_3790,N_2339,N_2300);
or U3791 (N_3791,N_2294,N_2962);
and U3792 (N_3792,N_2243,N_2559);
xor U3793 (N_3793,N_2184,N_2447);
nand U3794 (N_3794,N_2228,N_2409);
nor U3795 (N_3795,N_2729,N_2666);
nor U3796 (N_3796,N_2649,N_2962);
nor U3797 (N_3797,N_2423,N_2074);
nor U3798 (N_3798,N_2465,N_2525);
nand U3799 (N_3799,N_2953,N_2470);
and U3800 (N_3800,N_2353,N_2721);
and U3801 (N_3801,N_2661,N_2068);
nand U3802 (N_3802,N_2025,N_2095);
or U3803 (N_3803,N_2144,N_2857);
nand U3804 (N_3804,N_2072,N_2866);
and U3805 (N_3805,N_2252,N_2548);
nor U3806 (N_3806,N_2697,N_2543);
or U3807 (N_3807,N_2767,N_2910);
and U3808 (N_3808,N_2474,N_2941);
nor U3809 (N_3809,N_2091,N_2504);
xnor U3810 (N_3810,N_2088,N_2442);
or U3811 (N_3811,N_2171,N_2485);
or U3812 (N_3812,N_2411,N_2929);
nand U3813 (N_3813,N_2268,N_2307);
nand U3814 (N_3814,N_2794,N_2729);
or U3815 (N_3815,N_2144,N_2476);
nand U3816 (N_3816,N_2062,N_2684);
or U3817 (N_3817,N_2564,N_2418);
nand U3818 (N_3818,N_2089,N_2648);
nand U3819 (N_3819,N_2114,N_2204);
nor U3820 (N_3820,N_2894,N_2607);
and U3821 (N_3821,N_2123,N_2815);
and U3822 (N_3822,N_2021,N_2418);
nor U3823 (N_3823,N_2862,N_2678);
and U3824 (N_3824,N_2373,N_2332);
nor U3825 (N_3825,N_2611,N_2589);
nor U3826 (N_3826,N_2962,N_2106);
and U3827 (N_3827,N_2494,N_2678);
nand U3828 (N_3828,N_2482,N_2177);
and U3829 (N_3829,N_2863,N_2471);
or U3830 (N_3830,N_2292,N_2309);
xnor U3831 (N_3831,N_2196,N_2198);
nor U3832 (N_3832,N_2885,N_2843);
nor U3833 (N_3833,N_2205,N_2638);
and U3834 (N_3834,N_2241,N_2464);
and U3835 (N_3835,N_2405,N_2078);
nand U3836 (N_3836,N_2470,N_2443);
and U3837 (N_3837,N_2799,N_2868);
or U3838 (N_3838,N_2427,N_2078);
and U3839 (N_3839,N_2902,N_2834);
or U3840 (N_3840,N_2511,N_2325);
and U3841 (N_3841,N_2235,N_2503);
and U3842 (N_3842,N_2759,N_2242);
and U3843 (N_3843,N_2543,N_2466);
and U3844 (N_3844,N_2990,N_2985);
nand U3845 (N_3845,N_2663,N_2063);
nor U3846 (N_3846,N_2976,N_2378);
or U3847 (N_3847,N_2204,N_2628);
and U3848 (N_3848,N_2073,N_2544);
nor U3849 (N_3849,N_2089,N_2972);
or U3850 (N_3850,N_2126,N_2071);
xnor U3851 (N_3851,N_2611,N_2585);
or U3852 (N_3852,N_2442,N_2926);
or U3853 (N_3853,N_2077,N_2642);
and U3854 (N_3854,N_2173,N_2434);
or U3855 (N_3855,N_2224,N_2635);
nand U3856 (N_3856,N_2829,N_2009);
or U3857 (N_3857,N_2837,N_2805);
nor U3858 (N_3858,N_2169,N_2809);
or U3859 (N_3859,N_2267,N_2451);
xnor U3860 (N_3860,N_2011,N_2613);
nor U3861 (N_3861,N_2355,N_2391);
or U3862 (N_3862,N_2055,N_2337);
or U3863 (N_3863,N_2500,N_2978);
nand U3864 (N_3864,N_2445,N_2770);
nor U3865 (N_3865,N_2481,N_2117);
nand U3866 (N_3866,N_2513,N_2541);
nand U3867 (N_3867,N_2853,N_2441);
and U3868 (N_3868,N_2125,N_2721);
nor U3869 (N_3869,N_2289,N_2784);
and U3870 (N_3870,N_2356,N_2976);
nand U3871 (N_3871,N_2728,N_2059);
nand U3872 (N_3872,N_2138,N_2222);
and U3873 (N_3873,N_2396,N_2902);
nand U3874 (N_3874,N_2461,N_2835);
nor U3875 (N_3875,N_2954,N_2683);
nor U3876 (N_3876,N_2700,N_2467);
or U3877 (N_3877,N_2744,N_2324);
or U3878 (N_3878,N_2047,N_2780);
and U3879 (N_3879,N_2480,N_2769);
or U3880 (N_3880,N_2577,N_2635);
and U3881 (N_3881,N_2267,N_2610);
nand U3882 (N_3882,N_2679,N_2032);
nor U3883 (N_3883,N_2049,N_2850);
and U3884 (N_3884,N_2507,N_2159);
and U3885 (N_3885,N_2896,N_2582);
and U3886 (N_3886,N_2590,N_2759);
and U3887 (N_3887,N_2822,N_2918);
and U3888 (N_3888,N_2164,N_2513);
or U3889 (N_3889,N_2025,N_2708);
nand U3890 (N_3890,N_2065,N_2505);
or U3891 (N_3891,N_2673,N_2221);
or U3892 (N_3892,N_2540,N_2241);
or U3893 (N_3893,N_2719,N_2807);
nor U3894 (N_3894,N_2094,N_2451);
nor U3895 (N_3895,N_2276,N_2369);
nor U3896 (N_3896,N_2894,N_2204);
or U3897 (N_3897,N_2003,N_2013);
and U3898 (N_3898,N_2299,N_2368);
nor U3899 (N_3899,N_2361,N_2613);
or U3900 (N_3900,N_2316,N_2144);
nor U3901 (N_3901,N_2771,N_2946);
nand U3902 (N_3902,N_2598,N_2214);
and U3903 (N_3903,N_2858,N_2595);
and U3904 (N_3904,N_2483,N_2280);
and U3905 (N_3905,N_2973,N_2201);
and U3906 (N_3906,N_2731,N_2361);
and U3907 (N_3907,N_2567,N_2146);
nand U3908 (N_3908,N_2687,N_2156);
nand U3909 (N_3909,N_2691,N_2110);
nand U3910 (N_3910,N_2229,N_2010);
nand U3911 (N_3911,N_2208,N_2371);
or U3912 (N_3912,N_2421,N_2899);
or U3913 (N_3913,N_2319,N_2519);
nor U3914 (N_3914,N_2395,N_2166);
nand U3915 (N_3915,N_2884,N_2095);
and U3916 (N_3916,N_2168,N_2540);
nand U3917 (N_3917,N_2846,N_2555);
and U3918 (N_3918,N_2708,N_2540);
or U3919 (N_3919,N_2688,N_2118);
or U3920 (N_3920,N_2337,N_2139);
or U3921 (N_3921,N_2946,N_2907);
and U3922 (N_3922,N_2492,N_2898);
nand U3923 (N_3923,N_2763,N_2703);
or U3924 (N_3924,N_2626,N_2260);
xnor U3925 (N_3925,N_2995,N_2091);
nor U3926 (N_3926,N_2135,N_2396);
nor U3927 (N_3927,N_2708,N_2790);
and U3928 (N_3928,N_2314,N_2634);
nor U3929 (N_3929,N_2833,N_2783);
or U3930 (N_3930,N_2884,N_2893);
and U3931 (N_3931,N_2884,N_2166);
and U3932 (N_3932,N_2410,N_2516);
nand U3933 (N_3933,N_2367,N_2521);
nand U3934 (N_3934,N_2163,N_2090);
nand U3935 (N_3935,N_2227,N_2677);
and U3936 (N_3936,N_2818,N_2367);
and U3937 (N_3937,N_2921,N_2085);
or U3938 (N_3938,N_2942,N_2878);
and U3939 (N_3939,N_2307,N_2377);
nand U3940 (N_3940,N_2677,N_2220);
nor U3941 (N_3941,N_2677,N_2733);
or U3942 (N_3942,N_2849,N_2857);
and U3943 (N_3943,N_2839,N_2163);
and U3944 (N_3944,N_2686,N_2592);
or U3945 (N_3945,N_2449,N_2849);
nor U3946 (N_3946,N_2572,N_2624);
and U3947 (N_3947,N_2664,N_2610);
and U3948 (N_3948,N_2469,N_2778);
and U3949 (N_3949,N_2665,N_2855);
nor U3950 (N_3950,N_2537,N_2195);
nor U3951 (N_3951,N_2116,N_2154);
or U3952 (N_3952,N_2839,N_2130);
nor U3953 (N_3953,N_2413,N_2419);
and U3954 (N_3954,N_2860,N_2949);
nand U3955 (N_3955,N_2927,N_2149);
and U3956 (N_3956,N_2063,N_2780);
nor U3957 (N_3957,N_2833,N_2234);
nand U3958 (N_3958,N_2781,N_2110);
or U3959 (N_3959,N_2508,N_2399);
nand U3960 (N_3960,N_2742,N_2891);
nand U3961 (N_3961,N_2911,N_2714);
nor U3962 (N_3962,N_2756,N_2333);
xor U3963 (N_3963,N_2400,N_2414);
nor U3964 (N_3964,N_2496,N_2199);
or U3965 (N_3965,N_2940,N_2139);
nor U3966 (N_3966,N_2904,N_2916);
nand U3967 (N_3967,N_2350,N_2054);
or U3968 (N_3968,N_2556,N_2781);
nor U3969 (N_3969,N_2699,N_2000);
nor U3970 (N_3970,N_2728,N_2552);
xor U3971 (N_3971,N_2953,N_2041);
nor U3972 (N_3972,N_2991,N_2554);
nand U3973 (N_3973,N_2453,N_2112);
nor U3974 (N_3974,N_2503,N_2138);
nand U3975 (N_3975,N_2484,N_2850);
and U3976 (N_3976,N_2390,N_2045);
or U3977 (N_3977,N_2373,N_2658);
nand U3978 (N_3978,N_2134,N_2090);
nor U3979 (N_3979,N_2263,N_2772);
nand U3980 (N_3980,N_2270,N_2254);
nand U3981 (N_3981,N_2846,N_2402);
nand U3982 (N_3982,N_2360,N_2171);
nand U3983 (N_3983,N_2613,N_2448);
nor U3984 (N_3984,N_2096,N_2596);
nand U3985 (N_3985,N_2212,N_2265);
nand U3986 (N_3986,N_2664,N_2834);
nand U3987 (N_3987,N_2706,N_2307);
and U3988 (N_3988,N_2977,N_2842);
and U3989 (N_3989,N_2515,N_2274);
nor U3990 (N_3990,N_2962,N_2891);
xor U3991 (N_3991,N_2143,N_2818);
and U3992 (N_3992,N_2876,N_2944);
nand U3993 (N_3993,N_2023,N_2357);
and U3994 (N_3994,N_2619,N_2631);
nor U3995 (N_3995,N_2785,N_2365);
and U3996 (N_3996,N_2512,N_2194);
or U3997 (N_3997,N_2611,N_2938);
and U3998 (N_3998,N_2375,N_2119);
nor U3999 (N_3999,N_2616,N_2042);
and U4000 (N_4000,N_3897,N_3848);
nand U4001 (N_4001,N_3288,N_3998);
nand U4002 (N_4002,N_3626,N_3526);
xor U4003 (N_4003,N_3579,N_3721);
and U4004 (N_4004,N_3282,N_3300);
nor U4005 (N_4005,N_3661,N_3195);
and U4006 (N_4006,N_3126,N_3436);
and U4007 (N_4007,N_3143,N_3454);
and U4008 (N_4008,N_3482,N_3024);
nand U4009 (N_4009,N_3926,N_3017);
or U4010 (N_4010,N_3748,N_3975);
nand U4011 (N_4011,N_3197,N_3620);
nor U4012 (N_4012,N_3874,N_3809);
nor U4013 (N_4013,N_3459,N_3307);
nor U4014 (N_4014,N_3172,N_3398);
and U4015 (N_4015,N_3362,N_3391);
or U4016 (N_4016,N_3909,N_3237);
nand U4017 (N_4017,N_3051,N_3780);
nor U4018 (N_4018,N_3208,N_3228);
or U4019 (N_4019,N_3963,N_3733);
nor U4020 (N_4020,N_3325,N_3373);
or U4021 (N_4021,N_3885,N_3109);
nand U4022 (N_4022,N_3478,N_3512);
nor U4023 (N_4023,N_3054,N_3247);
xnor U4024 (N_4024,N_3778,N_3878);
nand U4025 (N_4025,N_3501,N_3404);
and U4026 (N_4026,N_3789,N_3930);
nor U4027 (N_4027,N_3133,N_3674);
nand U4028 (N_4028,N_3154,N_3792);
and U4029 (N_4029,N_3594,N_3900);
and U4030 (N_4030,N_3921,N_3184);
or U4031 (N_4031,N_3530,N_3424);
nand U4032 (N_4032,N_3899,N_3803);
nand U4033 (N_4033,N_3907,N_3774);
or U4034 (N_4034,N_3074,N_3528);
nor U4035 (N_4035,N_3816,N_3973);
nor U4036 (N_4036,N_3965,N_3444);
and U4037 (N_4037,N_3717,N_3319);
nor U4038 (N_4038,N_3376,N_3922);
or U4039 (N_4039,N_3912,N_3684);
nand U4040 (N_4040,N_3305,N_3953);
or U4041 (N_4041,N_3903,N_3324);
or U4042 (N_4042,N_3120,N_3974);
nor U4043 (N_4043,N_3189,N_3429);
and U4044 (N_4044,N_3776,N_3697);
or U4045 (N_4045,N_3249,N_3954);
nor U4046 (N_4046,N_3915,N_3648);
nand U4047 (N_4047,N_3556,N_3277);
and U4048 (N_4048,N_3862,N_3199);
and U4049 (N_4049,N_3524,N_3531);
nand U4050 (N_4050,N_3418,N_3934);
nor U4051 (N_4051,N_3308,N_3157);
nand U4052 (N_4052,N_3155,N_3700);
nor U4053 (N_4053,N_3236,N_3479);
and U4054 (N_4054,N_3811,N_3132);
or U4055 (N_4055,N_3507,N_3432);
or U4056 (N_4056,N_3165,N_3104);
or U4057 (N_4057,N_3583,N_3160);
nor U4058 (N_4058,N_3884,N_3229);
nor U4059 (N_4059,N_3231,N_3768);
or U4060 (N_4060,N_3353,N_3321);
and U4061 (N_4061,N_3272,N_3093);
nand U4062 (N_4062,N_3895,N_3591);
nand U4063 (N_4063,N_3191,N_3513);
or U4064 (N_4064,N_3536,N_3935);
and U4065 (N_4065,N_3187,N_3474);
nor U4066 (N_4066,N_3727,N_3676);
or U4067 (N_4067,N_3044,N_3703);
nand U4068 (N_4068,N_3629,N_3723);
nand U4069 (N_4069,N_3366,N_3240);
or U4070 (N_4070,N_3538,N_3711);
nand U4071 (N_4071,N_3076,N_3864);
nand U4072 (N_4072,N_3215,N_3204);
xor U4073 (N_4073,N_3053,N_3570);
or U4074 (N_4074,N_3597,N_3254);
or U4075 (N_4075,N_3564,N_3908);
or U4076 (N_4076,N_3483,N_3415);
nand U4077 (N_4077,N_3442,N_3218);
nand U4078 (N_4078,N_3749,N_3781);
or U4079 (N_4079,N_3818,N_3286);
xor U4080 (N_4080,N_3738,N_3535);
nor U4081 (N_4081,N_3057,N_3534);
or U4082 (N_4082,N_3219,N_3639);
nor U4083 (N_4083,N_3421,N_3274);
nor U4084 (N_4084,N_3266,N_3633);
nor U4085 (N_4085,N_3726,N_3735);
nor U4086 (N_4086,N_3110,N_3206);
nor U4087 (N_4087,N_3841,N_3461);
and U4088 (N_4088,N_3549,N_3151);
or U4089 (N_4089,N_3147,N_3081);
or U4090 (N_4090,N_3139,N_3635);
nand U4091 (N_4091,N_3656,N_3599);
and U4092 (N_4092,N_3420,N_3060);
and U4093 (N_4093,N_3007,N_3441);
and U4094 (N_4094,N_3271,N_3381);
or U4095 (N_4095,N_3258,N_3730);
nor U4096 (N_4096,N_3682,N_3622);
and U4097 (N_4097,N_3710,N_3498);
or U4098 (N_4098,N_3281,N_3625);
or U4099 (N_4099,N_3849,N_3980);
nand U4100 (N_4100,N_3539,N_3660);
nand U4101 (N_4101,N_3259,N_3572);
xor U4102 (N_4102,N_3532,N_3744);
or U4103 (N_4103,N_3171,N_3119);
nor U4104 (N_4104,N_3672,N_3425);
xnor U4105 (N_4105,N_3722,N_3244);
or U4106 (N_4106,N_3829,N_3011);
nand U4107 (N_4107,N_3956,N_3791);
or U4108 (N_4108,N_3868,N_3801);
and U4109 (N_4109,N_3890,N_3823);
nor U4110 (N_4110,N_3072,N_3758);
nor U4111 (N_4111,N_3762,N_3417);
xnor U4112 (N_4112,N_3142,N_3018);
nor U4113 (N_4113,N_3031,N_3224);
and U4114 (N_4114,N_3159,N_3509);
nand U4115 (N_4115,N_3357,N_3090);
nor U4116 (N_4116,N_3161,N_3642);
and U4117 (N_4117,N_3506,N_3951);
or U4118 (N_4118,N_3402,N_3222);
and U4119 (N_4119,N_3616,N_3317);
and U4120 (N_4120,N_3323,N_3669);
nor U4121 (N_4121,N_3386,N_3678);
and U4122 (N_4122,N_3784,N_3731);
nand U4123 (N_4123,N_3587,N_3632);
and U4124 (N_4124,N_3799,N_3690);
and U4125 (N_4125,N_3555,N_3872);
nand U4126 (N_4126,N_3099,N_3565);
and U4127 (N_4127,N_3576,N_3964);
xor U4128 (N_4128,N_3743,N_3455);
and U4129 (N_4129,N_3514,N_3059);
and U4130 (N_4130,N_3061,N_3295);
or U4131 (N_4131,N_3527,N_3028);
or U4132 (N_4132,N_3148,N_3447);
and U4133 (N_4133,N_3210,N_3268);
and U4134 (N_4134,N_3405,N_3706);
and U4135 (N_4135,N_3313,N_3430);
and U4136 (N_4136,N_3796,N_3888);
nand U4137 (N_4137,N_3947,N_3794);
nor U4138 (N_4138,N_3709,N_3067);
or U4139 (N_4139,N_3141,N_3001);
nand U4140 (N_4140,N_3752,N_3624);
or U4141 (N_4141,N_3085,N_3611);
and U4142 (N_4142,N_3886,N_3716);
and U4143 (N_4143,N_3248,N_3170);
or U4144 (N_4144,N_3855,N_3857);
and U4145 (N_4145,N_3867,N_3480);
nand U4146 (N_4146,N_3466,N_3440);
nor U4147 (N_4147,N_3005,N_3983);
nand U4148 (N_4148,N_3808,N_3560);
or U4149 (N_4149,N_3894,N_3239);
xor U4150 (N_4150,N_3663,N_3688);
nand U4151 (N_4151,N_3988,N_3203);
or U4152 (N_4152,N_3986,N_3765);
or U4153 (N_4153,N_3056,N_3990);
and U4154 (N_4154,N_3033,N_3102);
and U4155 (N_4155,N_3250,N_3677);
and U4156 (N_4156,N_3994,N_3987);
and U4157 (N_4157,N_3496,N_3377);
nor U4158 (N_4158,N_3100,N_3696);
and U4159 (N_4159,N_3458,N_3837);
xnor U4160 (N_4160,N_3827,N_3223);
nor U4161 (N_4161,N_3438,N_3006);
and U4162 (N_4162,N_3190,N_3860);
nor U4163 (N_4163,N_3844,N_3264);
and U4164 (N_4164,N_3450,N_3260);
or U4165 (N_4165,N_3217,N_3221);
nor U4166 (N_4166,N_3788,N_3253);
or U4167 (N_4167,N_3766,N_3169);
nand U4168 (N_4168,N_3437,N_3227);
nand U4169 (N_4169,N_3123,N_3097);
or U4170 (N_4170,N_3741,N_3972);
and U4171 (N_4171,N_3374,N_3718);
or U4172 (N_4172,N_3449,N_3861);
nor U4173 (N_4173,N_3847,N_3737);
nor U4174 (N_4174,N_3771,N_3675);
nor U4175 (N_4175,N_3544,N_3981);
nor U4176 (N_4176,N_3877,N_3755);
and U4177 (N_4177,N_3692,N_3826);
or U4178 (N_4178,N_3651,N_3108);
nor U4179 (N_4179,N_3403,N_3640);
nand U4180 (N_4180,N_3138,N_3233);
and U4181 (N_4181,N_3529,N_3087);
nand U4182 (N_4182,N_3122,N_3853);
xor U4183 (N_4183,N_3802,N_3783);
nand U4184 (N_4184,N_3773,N_3378);
nor U4185 (N_4185,N_3955,N_3393);
and U4186 (N_4186,N_3601,N_3166);
nor U4187 (N_4187,N_3049,N_3314);
or U4188 (N_4188,N_3959,N_3698);
or U4189 (N_4189,N_3163,N_3763);
nor U4190 (N_4190,N_3623,N_3607);
and U4191 (N_4191,N_3838,N_3186);
nand U4192 (N_4192,N_3495,N_3694);
nand U4193 (N_4193,N_3702,N_3129);
or U4194 (N_4194,N_3604,N_3304);
nand U4195 (N_4195,N_3898,N_3545);
nor U4196 (N_4196,N_3786,N_3106);
or U4197 (N_4197,N_3293,N_3997);
nor U4198 (N_4198,N_3364,N_3645);
nor U4199 (N_4199,N_3380,N_3948);
or U4200 (N_4200,N_3306,N_3043);
and U4201 (N_4201,N_3636,N_3358);
nor U4202 (N_4202,N_3414,N_3365);
nand U4203 (N_4203,N_3095,N_3326);
nand U4204 (N_4204,N_3338,N_3124);
nor U4205 (N_4205,N_3705,N_3606);
or U4206 (N_4206,N_3052,N_3736);
nor U4207 (N_4207,N_3562,N_3029);
nand U4208 (N_4208,N_3416,N_3055);
nand U4209 (N_4209,N_3569,N_3265);
nor U4210 (N_4210,N_3658,N_3379);
nor U4211 (N_4211,N_3234,N_3194);
or U4212 (N_4212,N_3932,N_3654);
nor U4213 (N_4213,N_3671,N_3634);
nand U4214 (N_4214,N_3164,N_3817);
nand U4215 (N_4215,N_3499,N_3284);
or U4216 (N_4216,N_3088,N_3410);
xnor U4217 (N_4217,N_3214,N_3021);
xnor U4218 (N_4218,N_3685,N_3261);
or U4219 (N_4219,N_3232,N_3540);
and U4220 (N_4220,N_3349,N_3002);
nand U4221 (N_4221,N_3027,N_3708);
nand U4222 (N_4222,N_3278,N_3422);
or U4223 (N_4223,N_3940,N_3038);
nor U4224 (N_4224,N_3201,N_3256);
nor U4225 (N_4225,N_3889,N_3828);
and U4226 (N_4226,N_3121,N_3519);
and U4227 (N_4227,N_3263,N_3135);
nor U4228 (N_4228,N_3621,N_3009);
or U4229 (N_4229,N_3946,N_3985);
and U4230 (N_4230,N_3439,N_3875);
nand U4231 (N_4231,N_3580,N_3389);
or U4232 (N_4232,N_3968,N_3650);
and U4233 (N_4233,N_3329,N_3064);
nor U4234 (N_4234,N_3463,N_3746);
nor U4235 (N_4235,N_3020,N_3824);
and U4236 (N_4236,N_3497,N_3352);
nor U4237 (N_4237,N_3891,N_3942);
or U4238 (N_4238,N_3026,N_3967);
nand U4239 (N_4239,N_3595,N_3873);
nand U4240 (N_4240,N_3825,N_3850);
xor U4241 (N_4241,N_3198,N_3945);
and U4242 (N_4242,N_3666,N_3173);
and U4243 (N_4243,N_3557,N_3992);
nor U4244 (N_4244,N_3042,N_3925);
nor U4245 (N_4245,N_3392,N_3941);
and U4246 (N_4246,N_3332,N_3000);
or U4247 (N_4247,N_3558,N_3114);
nand U4248 (N_4248,N_3798,N_3046);
or U4249 (N_4249,N_3168,N_3073);
or U4250 (N_4250,N_3999,N_3918);
or U4251 (N_4251,N_3388,N_3301);
nand U4252 (N_4252,N_3176,N_3759);
and U4253 (N_4253,N_3494,N_3542);
nand U4254 (N_4254,N_3618,N_3695);
or U4255 (N_4255,N_3318,N_3807);
nor U4256 (N_4256,N_3525,N_3851);
nor U4257 (N_4257,N_3916,N_3511);
and U4258 (N_4258,N_3866,N_3036);
or U4259 (N_4259,N_3423,N_3775);
xnor U4260 (N_4260,N_3267,N_3348);
or U4261 (N_4261,N_3728,N_3050);
or U4262 (N_4262,N_3322,N_3615);
and U4263 (N_4263,N_3220,N_3182);
nor U4264 (N_4264,N_3832,N_3516);
nand U4265 (N_4265,N_3019,N_3991);
nand U4266 (N_4266,N_3905,N_3814);
and U4267 (N_4267,N_3846,N_3559);
nor U4268 (N_4268,N_3115,N_3665);
nor U4269 (N_4269,N_3181,N_3071);
and U4270 (N_4270,N_3822,N_3012);
and U4271 (N_4271,N_3150,N_3657);
nor U4272 (N_4272,N_3434,N_3069);
nor U4273 (N_4273,N_3107,N_3724);
nor U4274 (N_4274,N_3729,N_3996);
nor U4275 (N_4275,N_3931,N_3333);
nand U4276 (N_4276,N_3299,N_3681);
nand U4277 (N_4277,N_3294,N_3298);
and U4278 (N_4278,N_3030,N_3966);
nand U4279 (N_4279,N_3128,N_3297);
and U4280 (N_4280,N_3520,N_3476);
nand U4281 (N_4281,N_3910,N_3655);
and U4282 (N_4282,N_3103,N_3679);
nand U4283 (N_4283,N_3091,N_3500);
nand U4284 (N_4284,N_3839,N_3831);
and U4285 (N_4285,N_3785,N_3149);
and U4286 (N_4286,N_3004,N_3035);
nand U4287 (N_4287,N_3982,N_3359);
or U4288 (N_4288,N_3969,N_3670);
or U4289 (N_4289,N_3750,N_3887);
and U4290 (N_4290,N_3384,N_3270);
nand U4291 (N_4291,N_3068,N_3334);
or U4292 (N_4292,N_3772,N_3285);
nor U4293 (N_4293,N_3252,N_3761);
and U4294 (N_4294,N_3486,N_3911);
nor U4295 (N_4295,N_3567,N_3316);
nand U4296 (N_4296,N_3689,N_3659);
nand U4297 (N_4297,N_3287,N_3541);
or U4298 (N_4298,N_3901,N_3086);
and U4299 (N_4299,N_3720,N_3156);
or U4300 (N_4300,N_3105,N_3394);
and U4301 (N_4301,N_3602,N_3586);
nor U4302 (N_4302,N_3464,N_3938);
and U4303 (N_4303,N_3489,N_3976);
nor U4304 (N_4304,N_3754,N_3631);
or U4305 (N_4305,N_3605,N_3638);
and U4306 (N_4306,N_3578,N_3646);
or U4307 (N_4307,N_3315,N_3856);
nor U4308 (N_4308,N_3205,N_3854);
nand U4309 (N_4309,N_3082,N_3577);
nor U4310 (N_4310,N_3207,N_3913);
or U4311 (N_4311,N_3339,N_3243);
nand U4312 (N_4312,N_3815,N_3547);
or U4313 (N_4313,N_3810,N_3008);
nand U4314 (N_4314,N_3238,N_3643);
and U4315 (N_4315,N_3445,N_3821);
or U4316 (N_4316,N_3637,N_3714);
nor U4317 (N_4317,N_3032,N_3504);
nor U4318 (N_4318,N_3034,N_3523);
or U4319 (N_4319,N_3242,N_3834);
or U4320 (N_4320,N_3255,N_3460);
or U4321 (N_4321,N_3769,N_3928);
or U4322 (N_4322,N_3448,N_3715);
nor U4323 (N_4323,N_3995,N_3153);
or U4324 (N_4324,N_3537,N_3667);
nand U4325 (N_4325,N_3058,N_3977);
and U4326 (N_4326,N_3490,N_3593);
or U4327 (N_4327,N_3452,N_3614);
and U4328 (N_4328,N_3943,N_3673);
or U4329 (N_4329,N_3131,N_3734);
or U4330 (N_4330,N_3896,N_3196);
nand U4331 (N_4331,N_3686,N_3664);
or U4332 (N_4332,N_3446,N_3162);
nand U4333 (N_4333,N_3427,N_3978);
nor U4334 (N_4334,N_3211,N_3820);
or U4335 (N_4335,N_3971,N_3309);
nor U4336 (N_4336,N_3335,N_3302);
nor U4337 (N_4337,N_3411,N_3707);
and U4338 (N_4338,N_3573,N_3662);
and U4339 (N_4339,N_3465,N_3041);
nand U4340 (N_4340,N_3096,N_3739);
xor U4341 (N_4341,N_3962,N_3040);
nand U4342 (N_4342,N_3062,N_3701);
and U4343 (N_4343,N_3451,N_3683);
nor U4344 (N_4344,N_3279,N_3371);
or U4345 (N_4345,N_3174,N_3280);
or U4346 (N_4346,N_3883,N_3613);
and U4347 (N_4347,N_3225,N_3797);
and U4348 (N_4348,N_3312,N_3603);
or U4349 (N_4349,N_3691,N_3543);
and U4350 (N_4350,N_3767,N_3732);
nand U4351 (N_4351,N_3551,N_3713);
nor U4352 (N_4352,N_3952,N_3048);
xor U4353 (N_4353,N_3845,N_3399);
nand U4354 (N_4354,N_3443,N_3111);
nor U4355 (N_4355,N_3892,N_3617);
and U4356 (N_4356,N_3342,N_3262);
or U4357 (N_4357,N_3257,N_3116);
nand U4358 (N_4358,N_3876,N_3078);
nor U4359 (N_4359,N_3275,N_3840);
nand U4360 (N_4360,N_3370,N_3283);
or U4361 (N_4361,N_3481,N_3598);
nand U4362 (N_4362,N_3177,N_3241);
and U4363 (N_4363,N_3144,N_3117);
and U4364 (N_4364,N_3047,N_3612);
nand U4365 (N_4365,N_3515,N_3406);
or U4366 (N_4366,N_3508,N_3118);
and U4367 (N_4367,N_3568,N_3193);
nor U4368 (N_4368,N_3098,N_3518);
nand U4369 (N_4369,N_3368,N_3467);
nand U4370 (N_4370,N_3561,N_3344);
nand U4371 (N_4371,N_3488,N_3045);
and U4372 (N_4372,N_3492,N_3209);
nand U4373 (N_4373,N_3296,N_3653);
or U4374 (N_4374,N_3906,N_3320);
nand U4375 (N_4375,N_3944,N_3075);
and U4376 (N_4376,N_3929,N_3014);
nand U4377 (N_4377,N_3600,N_3367);
nand U4378 (N_4378,N_3372,N_3037);
and U4379 (N_4379,N_3079,N_3858);
or U4380 (N_4380,N_3291,N_3533);
and U4381 (N_4381,N_3226,N_3251);
nor U4382 (N_4382,N_3083,N_3395);
xor U4383 (N_4383,N_3125,N_3812);
or U4384 (N_4384,N_3751,N_3958);
and U4385 (N_4385,N_3927,N_3553);
nor U4386 (N_4386,N_3902,N_3369);
or U4387 (N_4387,N_3596,N_3167);
nor U4388 (N_4388,N_3428,N_3094);
or U4389 (N_4389,N_3200,N_3522);
nand U4390 (N_4390,N_3770,N_3584);
nor U4391 (N_4391,N_3077,N_3276);
and U4392 (N_4392,N_3341,N_3409);
nor U4393 (N_4393,N_3022,N_3649);
nand U4394 (N_4394,N_3363,N_3936);
nand U4395 (N_4395,N_3830,N_3468);
nand U4396 (N_4396,N_3039,N_3003);
nor U4397 (N_4397,N_3870,N_3419);
and U4398 (N_4398,N_3782,N_3136);
nor U4399 (N_4399,N_3484,N_3806);
nor U4400 (N_4400,N_3869,N_3188);
and U4401 (N_4401,N_3413,N_3063);
and U4402 (N_4402,N_3340,N_3979);
nand U4403 (N_4403,N_3813,N_3066);
or U4404 (N_4404,N_3949,N_3178);
or U4405 (N_4405,N_3957,N_3647);
and U4406 (N_4406,N_3134,N_3989);
or U4407 (N_4407,N_3375,N_3574);
or U4408 (N_4408,N_3493,N_3882);
or U4409 (N_4409,N_3546,N_3628);
nand U4410 (N_4410,N_3550,N_3548);
or U4411 (N_4411,N_3245,N_3354);
nand U4412 (N_4412,N_3343,N_3871);
and U4413 (N_4413,N_3585,N_3865);
nor U4414 (N_4414,N_3914,N_3347);
nor U4415 (N_4415,N_3015,N_3065);
and U4416 (N_4416,N_3581,N_3092);
and U4417 (N_4417,N_3269,N_3192);
nand U4418 (N_4418,N_3852,N_3202);
or U4419 (N_4419,N_3390,N_3350);
nor U4420 (N_4420,N_3330,N_3470);
nor U4421 (N_4421,N_3216,N_3311);
nor U4422 (N_4422,N_3939,N_3805);
nand U4423 (N_4423,N_3453,N_3431);
and U4424 (N_4424,N_3582,N_3725);
nand U4425 (N_4425,N_3668,N_3753);
and U4426 (N_4426,N_3346,N_3303);
or U4427 (N_4427,N_3327,N_3993);
and U4428 (N_4428,N_3070,N_3385);
nor U4429 (N_4429,N_3158,N_3757);
nand U4430 (N_4430,N_3212,N_3764);
nor U4431 (N_4431,N_3400,N_3641);
or U4432 (N_4432,N_3740,N_3505);
nand U4433 (N_4433,N_3893,N_3472);
nor U4434 (N_4434,N_3292,N_3933);
or U4435 (N_4435,N_3185,N_3473);
or U4436 (N_4436,N_3923,N_3310);
or U4437 (N_4437,N_3704,N_3491);
nor U4438 (N_4438,N_3793,N_3016);
nand U4439 (N_4439,N_3920,N_3880);
and U4440 (N_4440,N_3960,N_3879);
nor U4441 (N_4441,N_3485,N_3747);
nand U4442 (N_4442,N_3331,N_3010);
nor U4443 (N_4443,N_3089,N_3175);
and U4444 (N_4444,N_3502,N_3127);
nor U4445 (N_4445,N_3462,N_3627);
nand U4446 (N_4446,N_3804,N_3588);
or U4447 (N_4447,N_3712,N_3101);
or U4448 (N_4448,N_3795,N_3699);
or U4449 (N_4449,N_3563,N_3836);
nand U4450 (N_4450,N_3859,N_3407);
or U4451 (N_4451,N_3023,N_3113);
or U4452 (N_4452,N_3013,N_3644);
nor U4453 (N_4453,N_3235,N_3457);
or U4454 (N_4454,N_3435,N_3777);
and U4455 (N_4455,N_3383,N_3610);
and U4456 (N_4456,N_3970,N_3652);
nor U4457 (N_4457,N_3609,N_3760);
and U4458 (N_4458,N_3756,N_3779);
or U4459 (N_4459,N_3137,N_3566);
and U4460 (N_4460,N_3590,N_3408);
and U4461 (N_4461,N_3145,N_3503);
and U4462 (N_4462,N_3575,N_3937);
nand U4463 (N_4463,N_3351,N_3904);
nand U4464 (N_4464,N_3843,N_3475);
or U4465 (N_4465,N_3608,N_3140);
nor U4466 (N_4466,N_3881,N_3152);
xnor U4467 (N_4467,N_3517,N_3471);
nor U4468 (N_4468,N_3180,N_3521);
nand U4469 (N_4469,N_3961,N_3924);
or U4470 (N_4470,N_3361,N_3552);
xnor U4471 (N_4471,N_3745,N_3412);
nand U4472 (N_4472,N_3842,N_3917);
nor U4473 (N_4473,N_3337,N_3179);
nand U4474 (N_4474,N_3919,N_3477);
nand U4475 (N_4475,N_3687,N_3130);
or U4476 (N_4476,N_3619,N_3336);
or U4477 (N_4477,N_3833,N_3290);
or U4478 (N_4478,N_3328,N_3356);
and U4479 (N_4479,N_3401,N_3387);
nand U4480 (N_4480,N_3571,N_3719);
and U4481 (N_4481,N_3950,N_3396);
and U4482 (N_4482,N_3456,N_3213);
nand U4483 (N_4483,N_3693,N_3487);
and U4484 (N_4484,N_3589,N_3787);
and U4485 (N_4485,N_3630,N_3084);
or U4486 (N_4486,N_3355,N_3510);
nand U4487 (N_4487,N_3742,N_3146);
nor U4488 (N_4488,N_3230,N_3025);
nand U4489 (N_4489,N_3397,N_3984);
or U4490 (N_4490,N_3835,N_3433);
and U4491 (N_4491,N_3183,N_3382);
and U4492 (N_4492,N_3554,N_3592);
nand U4493 (N_4493,N_3289,N_3680);
or U4494 (N_4494,N_3800,N_3790);
and U4495 (N_4495,N_3080,N_3246);
and U4496 (N_4496,N_3345,N_3273);
and U4497 (N_4497,N_3360,N_3819);
or U4498 (N_4498,N_3426,N_3112);
or U4499 (N_4499,N_3863,N_3469);
or U4500 (N_4500,N_3469,N_3089);
nor U4501 (N_4501,N_3367,N_3075);
nand U4502 (N_4502,N_3299,N_3105);
nand U4503 (N_4503,N_3971,N_3846);
or U4504 (N_4504,N_3131,N_3849);
or U4505 (N_4505,N_3757,N_3144);
and U4506 (N_4506,N_3513,N_3944);
nand U4507 (N_4507,N_3969,N_3804);
or U4508 (N_4508,N_3510,N_3170);
or U4509 (N_4509,N_3917,N_3050);
or U4510 (N_4510,N_3071,N_3024);
nand U4511 (N_4511,N_3832,N_3621);
or U4512 (N_4512,N_3594,N_3714);
and U4513 (N_4513,N_3960,N_3921);
nor U4514 (N_4514,N_3413,N_3982);
nand U4515 (N_4515,N_3791,N_3549);
nand U4516 (N_4516,N_3002,N_3769);
or U4517 (N_4517,N_3793,N_3506);
nand U4518 (N_4518,N_3422,N_3927);
and U4519 (N_4519,N_3595,N_3038);
nor U4520 (N_4520,N_3452,N_3132);
nand U4521 (N_4521,N_3974,N_3321);
nand U4522 (N_4522,N_3885,N_3064);
nor U4523 (N_4523,N_3022,N_3494);
or U4524 (N_4524,N_3777,N_3941);
and U4525 (N_4525,N_3632,N_3499);
nor U4526 (N_4526,N_3621,N_3356);
nand U4527 (N_4527,N_3850,N_3824);
nor U4528 (N_4528,N_3801,N_3648);
nor U4529 (N_4529,N_3026,N_3298);
nor U4530 (N_4530,N_3063,N_3886);
nand U4531 (N_4531,N_3581,N_3998);
and U4532 (N_4532,N_3224,N_3503);
nand U4533 (N_4533,N_3395,N_3355);
and U4534 (N_4534,N_3477,N_3843);
or U4535 (N_4535,N_3986,N_3839);
nor U4536 (N_4536,N_3476,N_3517);
and U4537 (N_4537,N_3351,N_3126);
or U4538 (N_4538,N_3950,N_3738);
and U4539 (N_4539,N_3525,N_3083);
and U4540 (N_4540,N_3115,N_3616);
and U4541 (N_4541,N_3696,N_3527);
or U4542 (N_4542,N_3807,N_3166);
nand U4543 (N_4543,N_3688,N_3206);
or U4544 (N_4544,N_3445,N_3334);
or U4545 (N_4545,N_3168,N_3464);
or U4546 (N_4546,N_3402,N_3467);
and U4547 (N_4547,N_3482,N_3021);
and U4548 (N_4548,N_3576,N_3891);
and U4549 (N_4549,N_3847,N_3360);
xnor U4550 (N_4550,N_3819,N_3672);
nand U4551 (N_4551,N_3357,N_3977);
and U4552 (N_4552,N_3052,N_3770);
nand U4553 (N_4553,N_3669,N_3504);
nor U4554 (N_4554,N_3633,N_3390);
or U4555 (N_4555,N_3540,N_3661);
or U4556 (N_4556,N_3930,N_3298);
nor U4557 (N_4557,N_3863,N_3445);
nand U4558 (N_4558,N_3910,N_3806);
and U4559 (N_4559,N_3632,N_3989);
nand U4560 (N_4560,N_3293,N_3545);
or U4561 (N_4561,N_3681,N_3746);
nor U4562 (N_4562,N_3704,N_3691);
and U4563 (N_4563,N_3740,N_3077);
and U4564 (N_4564,N_3896,N_3937);
or U4565 (N_4565,N_3239,N_3623);
nand U4566 (N_4566,N_3727,N_3355);
nand U4567 (N_4567,N_3136,N_3765);
and U4568 (N_4568,N_3823,N_3508);
and U4569 (N_4569,N_3400,N_3817);
nand U4570 (N_4570,N_3820,N_3382);
or U4571 (N_4571,N_3983,N_3561);
nand U4572 (N_4572,N_3544,N_3069);
nand U4573 (N_4573,N_3525,N_3632);
nand U4574 (N_4574,N_3793,N_3697);
nand U4575 (N_4575,N_3866,N_3685);
and U4576 (N_4576,N_3155,N_3178);
or U4577 (N_4577,N_3603,N_3280);
nand U4578 (N_4578,N_3408,N_3258);
or U4579 (N_4579,N_3514,N_3828);
nor U4580 (N_4580,N_3440,N_3458);
nand U4581 (N_4581,N_3427,N_3260);
and U4582 (N_4582,N_3604,N_3398);
nor U4583 (N_4583,N_3062,N_3866);
nor U4584 (N_4584,N_3195,N_3016);
nand U4585 (N_4585,N_3971,N_3990);
or U4586 (N_4586,N_3292,N_3063);
nand U4587 (N_4587,N_3967,N_3494);
and U4588 (N_4588,N_3188,N_3121);
nor U4589 (N_4589,N_3471,N_3053);
nor U4590 (N_4590,N_3933,N_3957);
or U4591 (N_4591,N_3741,N_3794);
nand U4592 (N_4592,N_3304,N_3102);
nand U4593 (N_4593,N_3591,N_3986);
nand U4594 (N_4594,N_3916,N_3750);
and U4595 (N_4595,N_3510,N_3614);
and U4596 (N_4596,N_3887,N_3989);
nand U4597 (N_4597,N_3125,N_3882);
or U4598 (N_4598,N_3874,N_3691);
nor U4599 (N_4599,N_3505,N_3638);
or U4600 (N_4600,N_3133,N_3507);
or U4601 (N_4601,N_3463,N_3340);
nand U4602 (N_4602,N_3056,N_3623);
or U4603 (N_4603,N_3445,N_3499);
and U4604 (N_4604,N_3484,N_3252);
and U4605 (N_4605,N_3816,N_3932);
nor U4606 (N_4606,N_3384,N_3475);
nor U4607 (N_4607,N_3861,N_3563);
nor U4608 (N_4608,N_3011,N_3804);
or U4609 (N_4609,N_3318,N_3747);
or U4610 (N_4610,N_3752,N_3704);
nor U4611 (N_4611,N_3115,N_3307);
nand U4612 (N_4612,N_3206,N_3150);
nand U4613 (N_4613,N_3666,N_3679);
nand U4614 (N_4614,N_3717,N_3299);
nor U4615 (N_4615,N_3276,N_3709);
nand U4616 (N_4616,N_3858,N_3393);
and U4617 (N_4617,N_3374,N_3981);
or U4618 (N_4618,N_3095,N_3823);
nand U4619 (N_4619,N_3564,N_3152);
and U4620 (N_4620,N_3411,N_3441);
nor U4621 (N_4621,N_3525,N_3840);
or U4622 (N_4622,N_3564,N_3287);
nand U4623 (N_4623,N_3705,N_3136);
or U4624 (N_4624,N_3923,N_3274);
nor U4625 (N_4625,N_3033,N_3231);
or U4626 (N_4626,N_3112,N_3962);
nand U4627 (N_4627,N_3946,N_3515);
nor U4628 (N_4628,N_3507,N_3190);
nor U4629 (N_4629,N_3835,N_3150);
or U4630 (N_4630,N_3410,N_3663);
or U4631 (N_4631,N_3436,N_3591);
or U4632 (N_4632,N_3654,N_3694);
nor U4633 (N_4633,N_3165,N_3217);
and U4634 (N_4634,N_3229,N_3738);
or U4635 (N_4635,N_3526,N_3694);
nand U4636 (N_4636,N_3361,N_3535);
or U4637 (N_4637,N_3157,N_3259);
nand U4638 (N_4638,N_3238,N_3227);
nand U4639 (N_4639,N_3649,N_3967);
nor U4640 (N_4640,N_3489,N_3675);
and U4641 (N_4641,N_3793,N_3817);
xor U4642 (N_4642,N_3895,N_3945);
nor U4643 (N_4643,N_3248,N_3439);
and U4644 (N_4644,N_3985,N_3185);
and U4645 (N_4645,N_3668,N_3107);
nor U4646 (N_4646,N_3472,N_3126);
and U4647 (N_4647,N_3313,N_3419);
nor U4648 (N_4648,N_3133,N_3419);
or U4649 (N_4649,N_3047,N_3532);
nor U4650 (N_4650,N_3574,N_3468);
nand U4651 (N_4651,N_3450,N_3838);
nor U4652 (N_4652,N_3464,N_3321);
and U4653 (N_4653,N_3263,N_3170);
or U4654 (N_4654,N_3357,N_3735);
or U4655 (N_4655,N_3263,N_3650);
or U4656 (N_4656,N_3006,N_3587);
or U4657 (N_4657,N_3405,N_3287);
or U4658 (N_4658,N_3534,N_3401);
nand U4659 (N_4659,N_3097,N_3509);
nor U4660 (N_4660,N_3560,N_3167);
nor U4661 (N_4661,N_3861,N_3151);
or U4662 (N_4662,N_3708,N_3731);
nor U4663 (N_4663,N_3004,N_3786);
nor U4664 (N_4664,N_3645,N_3104);
or U4665 (N_4665,N_3881,N_3275);
nor U4666 (N_4666,N_3987,N_3418);
or U4667 (N_4667,N_3550,N_3400);
nor U4668 (N_4668,N_3023,N_3932);
nor U4669 (N_4669,N_3344,N_3492);
or U4670 (N_4670,N_3669,N_3095);
nand U4671 (N_4671,N_3191,N_3438);
or U4672 (N_4672,N_3154,N_3608);
nand U4673 (N_4673,N_3048,N_3776);
nor U4674 (N_4674,N_3721,N_3779);
nand U4675 (N_4675,N_3067,N_3398);
or U4676 (N_4676,N_3387,N_3724);
or U4677 (N_4677,N_3036,N_3902);
nand U4678 (N_4678,N_3092,N_3388);
nor U4679 (N_4679,N_3388,N_3269);
or U4680 (N_4680,N_3276,N_3780);
nand U4681 (N_4681,N_3530,N_3549);
and U4682 (N_4682,N_3114,N_3115);
and U4683 (N_4683,N_3578,N_3458);
or U4684 (N_4684,N_3935,N_3821);
nor U4685 (N_4685,N_3619,N_3960);
nand U4686 (N_4686,N_3508,N_3871);
or U4687 (N_4687,N_3553,N_3317);
or U4688 (N_4688,N_3724,N_3949);
or U4689 (N_4689,N_3932,N_3160);
and U4690 (N_4690,N_3082,N_3204);
or U4691 (N_4691,N_3160,N_3187);
nand U4692 (N_4692,N_3545,N_3508);
or U4693 (N_4693,N_3936,N_3812);
and U4694 (N_4694,N_3474,N_3410);
nor U4695 (N_4695,N_3129,N_3141);
or U4696 (N_4696,N_3440,N_3557);
nor U4697 (N_4697,N_3930,N_3943);
nand U4698 (N_4698,N_3075,N_3543);
and U4699 (N_4699,N_3921,N_3069);
and U4700 (N_4700,N_3312,N_3549);
and U4701 (N_4701,N_3141,N_3254);
nor U4702 (N_4702,N_3537,N_3396);
nand U4703 (N_4703,N_3038,N_3228);
nand U4704 (N_4704,N_3643,N_3844);
and U4705 (N_4705,N_3418,N_3002);
nor U4706 (N_4706,N_3074,N_3783);
nor U4707 (N_4707,N_3279,N_3996);
nor U4708 (N_4708,N_3468,N_3299);
or U4709 (N_4709,N_3131,N_3371);
and U4710 (N_4710,N_3999,N_3193);
nand U4711 (N_4711,N_3787,N_3753);
nand U4712 (N_4712,N_3457,N_3504);
nand U4713 (N_4713,N_3068,N_3049);
nand U4714 (N_4714,N_3951,N_3767);
or U4715 (N_4715,N_3576,N_3278);
nor U4716 (N_4716,N_3048,N_3499);
nand U4717 (N_4717,N_3176,N_3648);
or U4718 (N_4718,N_3025,N_3358);
and U4719 (N_4719,N_3138,N_3601);
and U4720 (N_4720,N_3568,N_3831);
or U4721 (N_4721,N_3602,N_3088);
and U4722 (N_4722,N_3727,N_3983);
or U4723 (N_4723,N_3583,N_3890);
xor U4724 (N_4724,N_3123,N_3263);
or U4725 (N_4725,N_3180,N_3251);
and U4726 (N_4726,N_3985,N_3123);
and U4727 (N_4727,N_3454,N_3226);
nor U4728 (N_4728,N_3869,N_3595);
nand U4729 (N_4729,N_3073,N_3249);
or U4730 (N_4730,N_3433,N_3370);
and U4731 (N_4731,N_3640,N_3813);
nor U4732 (N_4732,N_3029,N_3548);
or U4733 (N_4733,N_3414,N_3798);
nand U4734 (N_4734,N_3838,N_3713);
or U4735 (N_4735,N_3206,N_3791);
nor U4736 (N_4736,N_3846,N_3793);
xnor U4737 (N_4737,N_3034,N_3610);
or U4738 (N_4738,N_3897,N_3686);
nand U4739 (N_4739,N_3089,N_3405);
nor U4740 (N_4740,N_3770,N_3517);
nand U4741 (N_4741,N_3061,N_3070);
nand U4742 (N_4742,N_3687,N_3364);
and U4743 (N_4743,N_3980,N_3141);
nand U4744 (N_4744,N_3236,N_3873);
nor U4745 (N_4745,N_3788,N_3311);
nand U4746 (N_4746,N_3245,N_3612);
and U4747 (N_4747,N_3302,N_3351);
and U4748 (N_4748,N_3618,N_3084);
nand U4749 (N_4749,N_3305,N_3230);
or U4750 (N_4750,N_3180,N_3955);
nand U4751 (N_4751,N_3451,N_3859);
nand U4752 (N_4752,N_3478,N_3556);
xnor U4753 (N_4753,N_3943,N_3185);
nor U4754 (N_4754,N_3395,N_3729);
nand U4755 (N_4755,N_3370,N_3325);
xnor U4756 (N_4756,N_3286,N_3939);
and U4757 (N_4757,N_3422,N_3817);
nand U4758 (N_4758,N_3561,N_3924);
nor U4759 (N_4759,N_3577,N_3234);
nor U4760 (N_4760,N_3370,N_3165);
nand U4761 (N_4761,N_3435,N_3956);
nor U4762 (N_4762,N_3411,N_3464);
and U4763 (N_4763,N_3008,N_3870);
or U4764 (N_4764,N_3114,N_3614);
nor U4765 (N_4765,N_3913,N_3778);
or U4766 (N_4766,N_3358,N_3253);
and U4767 (N_4767,N_3146,N_3545);
or U4768 (N_4768,N_3649,N_3966);
nand U4769 (N_4769,N_3453,N_3137);
or U4770 (N_4770,N_3624,N_3481);
or U4771 (N_4771,N_3093,N_3392);
or U4772 (N_4772,N_3235,N_3599);
and U4773 (N_4773,N_3398,N_3809);
nand U4774 (N_4774,N_3104,N_3677);
or U4775 (N_4775,N_3327,N_3222);
nand U4776 (N_4776,N_3491,N_3705);
or U4777 (N_4777,N_3700,N_3318);
and U4778 (N_4778,N_3855,N_3879);
nand U4779 (N_4779,N_3979,N_3806);
and U4780 (N_4780,N_3953,N_3417);
nor U4781 (N_4781,N_3317,N_3973);
nand U4782 (N_4782,N_3775,N_3084);
or U4783 (N_4783,N_3055,N_3529);
or U4784 (N_4784,N_3088,N_3404);
or U4785 (N_4785,N_3093,N_3034);
or U4786 (N_4786,N_3855,N_3751);
or U4787 (N_4787,N_3127,N_3921);
or U4788 (N_4788,N_3745,N_3684);
and U4789 (N_4789,N_3971,N_3193);
and U4790 (N_4790,N_3996,N_3376);
or U4791 (N_4791,N_3509,N_3892);
and U4792 (N_4792,N_3253,N_3049);
nand U4793 (N_4793,N_3700,N_3333);
and U4794 (N_4794,N_3647,N_3557);
nand U4795 (N_4795,N_3398,N_3639);
nor U4796 (N_4796,N_3045,N_3477);
or U4797 (N_4797,N_3194,N_3954);
and U4798 (N_4798,N_3781,N_3419);
nand U4799 (N_4799,N_3336,N_3297);
and U4800 (N_4800,N_3850,N_3941);
nor U4801 (N_4801,N_3979,N_3055);
or U4802 (N_4802,N_3217,N_3544);
nor U4803 (N_4803,N_3067,N_3713);
or U4804 (N_4804,N_3525,N_3734);
nor U4805 (N_4805,N_3760,N_3185);
and U4806 (N_4806,N_3856,N_3882);
xnor U4807 (N_4807,N_3676,N_3166);
nor U4808 (N_4808,N_3444,N_3226);
or U4809 (N_4809,N_3992,N_3122);
nor U4810 (N_4810,N_3481,N_3271);
nand U4811 (N_4811,N_3545,N_3521);
nor U4812 (N_4812,N_3747,N_3242);
or U4813 (N_4813,N_3075,N_3707);
nor U4814 (N_4814,N_3338,N_3318);
or U4815 (N_4815,N_3461,N_3371);
or U4816 (N_4816,N_3816,N_3551);
and U4817 (N_4817,N_3092,N_3730);
and U4818 (N_4818,N_3446,N_3868);
or U4819 (N_4819,N_3283,N_3846);
nor U4820 (N_4820,N_3853,N_3228);
or U4821 (N_4821,N_3051,N_3003);
and U4822 (N_4822,N_3758,N_3778);
nand U4823 (N_4823,N_3398,N_3331);
or U4824 (N_4824,N_3202,N_3166);
or U4825 (N_4825,N_3268,N_3400);
nand U4826 (N_4826,N_3767,N_3079);
or U4827 (N_4827,N_3054,N_3561);
nor U4828 (N_4828,N_3028,N_3735);
nor U4829 (N_4829,N_3444,N_3650);
nor U4830 (N_4830,N_3776,N_3465);
and U4831 (N_4831,N_3257,N_3847);
or U4832 (N_4832,N_3036,N_3637);
or U4833 (N_4833,N_3822,N_3415);
nor U4834 (N_4834,N_3977,N_3724);
or U4835 (N_4835,N_3793,N_3176);
xor U4836 (N_4836,N_3146,N_3306);
nor U4837 (N_4837,N_3729,N_3202);
nand U4838 (N_4838,N_3833,N_3192);
nor U4839 (N_4839,N_3747,N_3115);
or U4840 (N_4840,N_3094,N_3929);
nand U4841 (N_4841,N_3219,N_3239);
nor U4842 (N_4842,N_3428,N_3379);
nor U4843 (N_4843,N_3098,N_3418);
or U4844 (N_4844,N_3199,N_3038);
nand U4845 (N_4845,N_3837,N_3459);
or U4846 (N_4846,N_3737,N_3690);
and U4847 (N_4847,N_3179,N_3786);
nand U4848 (N_4848,N_3529,N_3936);
nor U4849 (N_4849,N_3324,N_3702);
or U4850 (N_4850,N_3914,N_3770);
and U4851 (N_4851,N_3763,N_3586);
or U4852 (N_4852,N_3313,N_3492);
and U4853 (N_4853,N_3793,N_3243);
or U4854 (N_4854,N_3648,N_3330);
nor U4855 (N_4855,N_3936,N_3640);
nand U4856 (N_4856,N_3832,N_3934);
and U4857 (N_4857,N_3759,N_3641);
and U4858 (N_4858,N_3079,N_3766);
or U4859 (N_4859,N_3213,N_3290);
or U4860 (N_4860,N_3529,N_3604);
and U4861 (N_4861,N_3358,N_3487);
or U4862 (N_4862,N_3320,N_3851);
and U4863 (N_4863,N_3341,N_3046);
or U4864 (N_4864,N_3351,N_3091);
nand U4865 (N_4865,N_3646,N_3223);
nor U4866 (N_4866,N_3009,N_3764);
and U4867 (N_4867,N_3769,N_3722);
nand U4868 (N_4868,N_3359,N_3564);
nor U4869 (N_4869,N_3503,N_3819);
nand U4870 (N_4870,N_3293,N_3922);
nor U4871 (N_4871,N_3886,N_3191);
and U4872 (N_4872,N_3791,N_3161);
or U4873 (N_4873,N_3712,N_3766);
nor U4874 (N_4874,N_3947,N_3896);
or U4875 (N_4875,N_3926,N_3364);
and U4876 (N_4876,N_3189,N_3019);
nor U4877 (N_4877,N_3992,N_3577);
and U4878 (N_4878,N_3959,N_3536);
or U4879 (N_4879,N_3993,N_3397);
or U4880 (N_4880,N_3128,N_3908);
nand U4881 (N_4881,N_3907,N_3914);
and U4882 (N_4882,N_3093,N_3438);
nor U4883 (N_4883,N_3490,N_3211);
or U4884 (N_4884,N_3684,N_3589);
xnor U4885 (N_4885,N_3260,N_3889);
nand U4886 (N_4886,N_3710,N_3984);
nor U4887 (N_4887,N_3529,N_3486);
and U4888 (N_4888,N_3235,N_3816);
or U4889 (N_4889,N_3032,N_3344);
nor U4890 (N_4890,N_3735,N_3718);
nand U4891 (N_4891,N_3685,N_3469);
and U4892 (N_4892,N_3817,N_3652);
nand U4893 (N_4893,N_3018,N_3314);
or U4894 (N_4894,N_3119,N_3837);
nand U4895 (N_4895,N_3533,N_3640);
nand U4896 (N_4896,N_3019,N_3719);
nor U4897 (N_4897,N_3684,N_3276);
nand U4898 (N_4898,N_3422,N_3472);
or U4899 (N_4899,N_3274,N_3656);
or U4900 (N_4900,N_3727,N_3492);
nor U4901 (N_4901,N_3519,N_3989);
and U4902 (N_4902,N_3318,N_3013);
nand U4903 (N_4903,N_3456,N_3799);
nand U4904 (N_4904,N_3786,N_3597);
and U4905 (N_4905,N_3903,N_3057);
nor U4906 (N_4906,N_3526,N_3076);
nand U4907 (N_4907,N_3184,N_3365);
or U4908 (N_4908,N_3042,N_3800);
and U4909 (N_4909,N_3441,N_3852);
and U4910 (N_4910,N_3502,N_3173);
or U4911 (N_4911,N_3507,N_3554);
or U4912 (N_4912,N_3179,N_3721);
nor U4913 (N_4913,N_3923,N_3574);
nand U4914 (N_4914,N_3589,N_3870);
nand U4915 (N_4915,N_3508,N_3141);
nor U4916 (N_4916,N_3341,N_3265);
or U4917 (N_4917,N_3241,N_3495);
and U4918 (N_4918,N_3568,N_3301);
nor U4919 (N_4919,N_3614,N_3158);
nor U4920 (N_4920,N_3887,N_3162);
and U4921 (N_4921,N_3656,N_3697);
nand U4922 (N_4922,N_3592,N_3359);
nor U4923 (N_4923,N_3255,N_3104);
or U4924 (N_4924,N_3865,N_3821);
xnor U4925 (N_4925,N_3469,N_3998);
or U4926 (N_4926,N_3332,N_3285);
nand U4927 (N_4927,N_3825,N_3195);
xnor U4928 (N_4928,N_3974,N_3775);
nand U4929 (N_4929,N_3280,N_3560);
nor U4930 (N_4930,N_3337,N_3132);
nor U4931 (N_4931,N_3505,N_3108);
nor U4932 (N_4932,N_3312,N_3910);
or U4933 (N_4933,N_3191,N_3505);
nand U4934 (N_4934,N_3543,N_3007);
nand U4935 (N_4935,N_3758,N_3057);
and U4936 (N_4936,N_3437,N_3535);
nor U4937 (N_4937,N_3443,N_3303);
nor U4938 (N_4938,N_3743,N_3083);
nand U4939 (N_4939,N_3783,N_3461);
or U4940 (N_4940,N_3754,N_3103);
or U4941 (N_4941,N_3041,N_3411);
or U4942 (N_4942,N_3420,N_3601);
and U4943 (N_4943,N_3953,N_3577);
nor U4944 (N_4944,N_3760,N_3130);
or U4945 (N_4945,N_3769,N_3625);
nor U4946 (N_4946,N_3977,N_3163);
nor U4947 (N_4947,N_3809,N_3146);
xnor U4948 (N_4948,N_3837,N_3531);
nand U4949 (N_4949,N_3846,N_3369);
nand U4950 (N_4950,N_3654,N_3814);
or U4951 (N_4951,N_3344,N_3176);
xor U4952 (N_4952,N_3682,N_3364);
and U4953 (N_4953,N_3835,N_3598);
nor U4954 (N_4954,N_3355,N_3453);
and U4955 (N_4955,N_3457,N_3547);
nand U4956 (N_4956,N_3472,N_3681);
and U4957 (N_4957,N_3911,N_3614);
nor U4958 (N_4958,N_3720,N_3700);
nand U4959 (N_4959,N_3639,N_3997);
nor U4960 (N_4960,N_3695,N_3476);
nor U4961 (N_4961,N_3921,N_3095);
or U4962 (N_4962,N_3694,N_3773);
nand U4963 (N_4963,N_3345,N_3531);
and U4964 (N_4964,N_3510,N_3938);
and U4965 (N_4965,N_3174,N_3989);
or U4966 (N_4966,N_3054,N_3130);
or U4967 (N_4967,N_3815,N_3000);
nor U4968 (N_4968,N_3515,N_3929);
or U4969 (N_4969,N_3032,N_3578);
nand U4970 (N_4970,N_3771,N_3782);
or U4971 (N_4971,N_3834,N_3496);
and U4972 (N_4972,N_3478,N_3009);
nand U4973 (N_4973,N_3460,N_3111);
nand U4974 (N_4974,N_3270,N_3320);
nand U4975 (N_4975,N_3674,N_3921);
or U4976 (N_4976,N_3572,N_3444);
and U4977 (N_4977,N_3407,N_3624);
and U4978 (N_4978,N_3432,N_3739);
and U4979 (N_4979,N_3849,N_3528);
nor U4980 (N_4980,N_3705,N_3455);
nor U4981 (N_4981,N_3485,N_3824);
and U4982 (N_4982,N_3419,N_3088);
and U4983 (N_4983,N_3804,N_3272);
nor U4984 (N_4984,N_3295,N_3275);
nand U4985 (N_4985,N_3227,N_3198);
nor U4986 (N_4986,N_3906,N_3831);
and U4987 (N_4987,N_3299,N_3227);
or U4988 (N_4988,N_3231,N_3717);
nand U4989 (N_4989,N_3113,N_3951);
and U4990 (N_4990,N_3978,N_3647);
xnor U4991 (N_4991,N_3894,N_3261);
or U4992 (N_4992,N_3075,N_3892);
and U4993 (N_4993,N_3557,N_3913);
nor U4994 (N_4994,N_3690,N_3978);
and U4995 (N_4995,N_3913,N_3733);
nor U4996 (N_4996,N_3999,N_3050);
or U4997 (N_4997,N_3615,N_3825);
nor U4998 (N_4998,N_3590,N_3285);
nand U4999 (N_4999,N_3685,N_3929);
nor UO_0 (O_0,N_4085,N_4437);
or UO_1 (O_1,N_4876,N_4631);
and UO_2 (O_2,N_4970,N_4801);
or UO_3 (O_3,N_4054,N_4786);
or UO_4 (O_4,N_4188,N_4208);
nor UO_5 (O_5,N_4517,N_4798);
and UO_6 (O_6,N_4294,N_4466);
nand UO_7 (O_7,N_4141,N_4377);
or UO_8 (O_8,N_4718,N_4788);
or UO_9 (O_9,N_4057,N_4857);
or UO_10 (O_10,N_4947,N_4866);
nor UO_11 (O_11,N_4845,N_4990);
nor UO_12 (O_12,N_4654,N_4711);
and UO_13 (O_13,N_4261,N_4564);
nand UO_14 (O_14,N_4872,N_4219);
or UO_15 (O_15,N_4722,N_4955);
and UO_16 (O_16,N_4216,N_4996);
nand UO_17 (O_17,N_4033,N_4330);
or UO_18 (O_18,N_4106,N_4563);
or UO_19 (O_19,N_4168,N_4127);
or UO_20 (O_20,N_4257,N_4913);
nand UO_21 (O_21,N_4815,N_4757);
or UO_22 (O_22,N_4074,N_4306);
nor UO_23 (O_23,N_4186,N_4122);
or UO_24 (O_24,N_4272,N_4067);
or UO_25 (O_25,N_4981,N_4781);
and UO_26 (O_26,N_4202,N_4077);
and UO_27 (O_27,N_4602,N_4376);
and UO_28 (O_28,N_4853,N_4280);
or UO_29 (O_29,N_4332,N_4819);
and UO_30 (O_30,N_4748,N_4427);
and UO_31 (O_31,N_4399,N_4941);
nand UO_32 (O_32,N_4824,N_4518);
nor UO_33 (O_33,N_4952,N_4243);
and UO_34 (O_34,N_4509,N_4938);
xor UO_35 (O_35,N_4934,N_4125);
nor UO_36 (O_36,N_4061,N_4855);
nand UO_37 (O_37,N_4449,N_4701);
or UO_38 (O_38,N_4283,N_4587);
nor UO_39 (O_39,N_4615,N_4205);
nor UO_40 (O_40,N_4327,N_4969);
and UO_41 (O_41,N_4155,N_4486);
and UO_42 (O_42,N_4162,N_4575);
or UO_43 (O_43,N_4707,N_4619);
nor UO_44 (O_44,N_4114,N_4369);
and UO_45 (O_45,N_4232,N_4789);
nor UO_46 (O_46,N_4726,N_4265);
or UO_47 (O_47,N_4424,N_4912);
and UO_48 (O_48,N_4165,N_4191);
nor UO_49 (O_49,N_4440,N_4679);
nand UO_50 (O_50,N_4378,N_4173);
nor UO_51 (O_51,N_4764,N_4428);
nand UO_52 (O_52,N_4020,N_4361);
nand UO_53 (O_53,N_4420,N_4292);
nor UO_54 (O_54,N_4861,N_4503);
nor UO_55 (O_55,N_4286,N_4864);
and UO_56 (O_56,N_4348,N_4989);
xor UO_57 (O_57,N_4833,N_4317);
and UO_58 (O_58,N_4953,N_4304);
and UO_59 (O_59,N_4710,N_4945);
nor UO_60 (O_60,N_4003,N_4431);
nor UO_61 (O_61,N_4533,N_4724);
and UO_62 (O_62,N_4562,N_4820);
nor UO_63 (O_63,N_4795,N_4901);
or UO_64 (O_64,N_4779,N_4279);
and UO_65 (O_65,N_4487,N_4406);
nor UO_66 (O_66,N_4800,N_4550);
nand UO_67 (O_67,N_4960,N_4675);
and UO_68 (O_68,N_4195,N_4719);
or UO_69 (O_69,N_4595,N_4805);
or UO_70 (O_70,N_4992,N_4418);
nor UO_71 (O_71,N_4485,N_4210);
nor UO_72 (O_72,N_4190,N_4611);
or UO_73 (O_73,N_4315,N_4612);
and UO_74 (O_74,N_4255,N_4300);
or UO_75 (O_75,N_4390,N_4303);
or UO_76 (O_76,N_4098,N_4018);
or UO_77 (O_77,N_4325,N_4183);
nand UO_78 (O_78,N_4973,N_4007);
and UO_79 (O_79,N_4596,N_4773);
and UO_80 (O_80,N_4759,N_4836);
nand UO_81 (O_81,N_4334,N_4715);
xor UO_82 (O_82,N_4523,N_4357);
xnor UO_83 (O_83,N_4561,N_4600);
nor UO_84 (O_84,N_4551,N_4967);
nor UO_85 (O_85,N_4356,N_4851);
and UO_86 (O_86,N_4481,N_4097);
or UO_87 (O_87,N_4096,N_4763);
or UO_88 (O_88,N_4252,N_4589);
and UO_89 (O_89,N_4863,N_4948);
nand UO_90 (O_90,N_4957,N_4352);
or UO_91 (O_91,N_4343,N_4609);
or UO_92 (O_92,N_4927,N_4438);
nand UO_93 (O_93,N_4075,N_4597);
nor UO_94 (O_94,N_4011,N_4884);
and UO_95 (O_95,N_4796,N_4787);
nor UO_96 (O_96,N_4213,N_4849);
and UO_97 (O_97,N_4289,N_4043);
and UO_98 (O_98,N_4476,N_4408);
xnor UO_99 (O_99,N_4460,N_4966);
or UO_100 (O_100,N_4873,N_4080);
and UO_101 (O_101,N_4834,N_4371);
or UO_102 (O_102,N_4331,N_4887);
and UO_103 (O_103,N_4919,N_4696);
and UO_104 (O_104,N_4549,N_4159);
nand UO_105 (O_105,N_4822,N_4547);
or UO_106 (O_106,N_4359,N_4342);
and UO_107 (O_107,N_4566,N_4986);
nor UO_108 (O_108,N_4178,N_4121);
nor UO_109 (O_109,N_4095,N_4275);
and UO_110 (O_110,N_4883,N_4504);
nor UO_111 (O_111,N_4137,N_4367);
nand UO_112 (O_112,N_4458,N_4678);
nor UO_113 (O_113,N_4015,N_4534);
and UO_114 (O_114,N_4119,N_4682);
and UO_115 (O_115,N_4840,N_4313);
nand UO_116 (O_116,N_4899,N_4312);
or UO_117 (O_117,N_4514,N_4383);
nand UO_118 (O_118,N_4405,N_4917);
or UO_119 (O_119,N_4245,N_4036);
or UO_120 (O_120,N_4598,N_4249);
and UO_121 (O_121,N_4666,N_4142);
nand UO_122 (O_122,N_4439,N_4635);
nand UO_123 (O_123,N_4025,N_4030);
or UO_124 (O_124,N_4374,N_4042);
or UO_125 (O_125,N_4146,N_4531);
nor UO_126 (O_126,N_4687,N_4461);
nor UO_127 (O_127,N_4070,N_4923);
nand UO_128 (O_128,N_4231,N_4634);
nand UO_129 (O_129,N_4591,N_4480);
and UO_130 (O_130,N_4997,N_4850);
nor UO_131 (O_131,N_4005,N_4854);
nand UO_132 (O_132,N_4267,N_4659);
nor UO_133 (O_133,N_4298,N_4637);
or UO_134 (O_134,N_4432,N_4049);
or UO_135 (O_135,N_4740,N_4237);
or UO_136 (O_136,N_4086,N_4254);
and UO_137 (O_137,N_4674,N_4290);
nand UO_138 (O_138,N_4536,N_4078);
nor UO_139 (O_139,N_4001,N_4541);
nand UO_140 (O_140,N_4964,N_4753);
nor UO_141 (O_141,N_4560,N_4818);
and UO_142 (O_142,N_4929,N_4457);
or UO_143 (O_143,N_4484,N_4410);
nand UO_144 (O_144,N_4475,N_4307);
nand UO_145 (O_145,N_4703,N_4738);
nor UO_146 (O_146,N_4120,N_4413);
nand UO_147 (O_147,N_4299,N_4856);
and UO_148 (O_148,N_4991,N_4758);
nand UO_149 (O_149,N_4994,N_4037);
and UO_150 (O_150,N_4502,N_4618);
or UO_151 (O_151,N_4409,N_4230);
and UO_152 (O_152,N_4971,N_4180);
nand UO_153 (O_153,N_4041,N_4101);
nand UO_154 (O_154,N_4130,N_4535);
and UO_155 (O_155,N_4124,N_4278);
or UO_156 (O_156,N_4351,N_4472);
or UO_157 (O_157,N_4895,N_4444);
nand UO_158 (O_158,N_4770,N_4453);
nor UO_159 (O_159,N_4281,N_4847);
and UO_160 (O_160,N_4594,N_4151);
nand UO_161 (O_161,N_4510,N_4639);
or UO_162 (O_162,N_4632,N_4364);
nor UO_163 (O_163,N_4578,N_4143);
and UO_164 (O_164,N_4058,N_4741);
nand UO_165 (O_165,N_4366,N_4823);
and UO_166 (O_166,N_4848,N_4987);
xnor UO_167 (O_167,N_4751,N_4211);
or UO_168 (O_168,N_4791,N_4236);
nand UO_169 (O_169,N_4203,N_4700);
and UO_170 (O_170,N_4749,N_4380);
nor UO_171 (O_171,N_4731,N_4720);
nand UO_172 (O_172,N_4745,N_4468);
and UO_173 (O_173,N_4404,N_4181);
and UO_174 (O_174,N_4209,N_4055);
or UO_175 (O_175,N_4746,N_4337);
and UO_176 (O_176,N_4094,N_4830);
nand UO_177 (O_177,N_4135,N_4580);
xnor UO_178 (O_178,N_4002,N_4425);
nand UO_179 (O_179,N_4527,N_4069);
or UO_180 (O_180,N_4668,N_4985);
xor UO_181 (O_181,N_4782,N_4925);
nor UO_182 (O_182,N_4489,N_4296);
nor UO_183 (O_183,N_4628,N_4047);
nand UO_184 (O_184,N_4318,N_4636);
nor UO_185 (O_185,N_4988,N_4276);
nor UO_186 (O_186,N_4153,N_4998);
nor UO_187 (O_187,N_4645,N_4835);
and UO_188 (O_188,N_4750,N_4525);
or UO_189 (O_189,N_4482,N_4762);
and UO_190 (O_190,N_4241,N_4083);
nor UO_191 (O_191,N_4694,N_4963);
and UO_192 (O_192,N_4262,N_4215);
nor UO_193 (O_193,N_4559,N_4398);
and UO_194 (O_194,N_4869,N_4214);
and UO_195 (O_195,N_4227,N_4508);
nor UO_196 (O_196,N_4898,N_4959);
or UO_197 (O_197,N_4396,N_4302);
or UO_198 (O_198,N_4322,N_4187);
or UO_199 (O_199,N_4630,N_4907);
nand UO_200 (O_200,N_4068,N_4071);
nor UO_201 (O_201,N_4921,N_4123);
and UO_202 (O_202,N_4827,N_4706);
or UO_203 (O_203,N_4138,N_4076);
and UO_204 (O_204,N_4223,N_4056);
or UO_205 (O_205,N_4975,N_4422);
xor UO_206 (O_206,N_4471,N_4900);
nor UO_207 (O_207,N_4350,N_4765);
nor UO_208 (O_208,N_4493,N_4045);
xnor UO_209 (O_209,N_4329,N_4050);
and UO_210 (O_210,N_4933,N_4958);
or UO_211 (O_211,N_4614,N_4004);
nand UO_212 (O_212,N_4584,N_4131);
or UO_213 (O_213,N_4344,N_4980);
nor UO_214 (O_214,N_4776,N_4160);
and UO_215 (O_215,N_4027,N_4282);
nand UO_216 (O_216,N_4736,N_4846);
and UO_217 (O_217,N_4809,N_4426);
nor UO_218 (O_218,N_4251,N_4224);
nand UO_219 (O_219,N_4530,N_4906);
and UO_220 (O_220,N_4553,N_4816);
nand UO_221 (O_221,N_4865,N_4586);
and UO_222 (O_222,N_4051,N_4662);
or UO_223 (O_223,N_4862,N_4113);
nor UO_224 (O_224,N_4295,N_4401);
nand UO_225 (O_225,N_4685,N_4752);
and UO_226 (O_226,N_4538,N_4543);
or UO_227 (O_227,N_4488,N_4200);
nor UO_228 (O_228,N_4347,N_4193);
or UO_229 (O_229,N_4412,N_4868);
nand UO_230 (O_230,N_4653,N_4995);
nand UO_231 (O_231,N_4924,N_4649);
or UO_232 (O_232,N_4260,N_4032);
nor UO_233 (O_233,N_4462,N_4837);
nand UO_234 (O_234,N_4977,N_4397);
nand UO_235 (O_235,N_4081,N_4768);
or UO_236 (O_236,N_4052,N_4402);
nand UO_237 (O_237,N_4381,N_4593);
and UO_238 (O_238,N_4499,N_4291);
nor UO_239 (O_239,N_4506,N_4297);
nor UO_240 (O_240,N_4500,N_4705);
nor UO_241 (O_241,N_4403,N_4017);
nor UO_242 (O_242,N_4680,N_4918);
nor UO_243 (O_243,N_4519,N_4567);
nor UO_244 (O_244,N_4524,N_4128);
or UO_245 (O_245,N_4091,N_4170);
and UO_246 (O_246,N_4035,N_4353);
or UO_247 (O_247,N_4393,N_4144);
and UO_248 (O_248,N_4743,N_4569);
nor UO_249 (O_249,N_4633,N_4175);
nor UO_250 (O_250,N_4698,N_4172);
or UO_251 (O_251,N_4684,N_4807);
and UO_252 (O_252,N_4733,N_4556);
or UO_253 (O_253,N_4670,N_4246);
nand UO_254 (O_254,N_4023,N_4881);
nor UO_255 (O_255,N_4790,N_4182);
nor UO_256 (O_256,N_4258,N_4459);
and UO_257 (O_257,N_4717,N_4365);
nor UO_258 (O_258,N_4326,N_4346);
or UO_259 (O_259,N_4423,N_4250);
and UO_260 (O_260,N_4646,N_4259);
or UO_261 (O_261,N_4844,N_4149);
or UO_262 (O_262,N_4605,N_4039);
nor UO_263 (O_263,N_4780,N_4708);
or UO_264 (O_264,N_4642,N_4742);
nor UO_265 (O_265,N_4529,N_4421);
and UO_266 (O_266,N_4812,N_4092);
nor UO_267 (O_267,N_4665,N_4681);
xor UO_268 (O_268,N_4000,N_4473);
nor UO_269 (O_269,N_4592,N_4648);
or UO_270 (O_270,N_4048,N_4341);
nor UO_271 (O_271,N_4308,N_4450);
and UO_272 (O_272,N_4944,N_4498);
and UO_273 (O_273,N_4414,N_4852);
nor UO_274 (O_274,N_4716,N_4494);
or UO_275 (O_275,N_4099,N_4803);
or UO_276 (O_276,N_4477,N_4419);
nand UO_277 (O_277,N_4238,N_4263);
and UO_278 (O_278,N_4744,N_4916);
nand UO_279 (O_279,N_4574,N_4842);
nor UO_280 (O_280,N_4777,N_4184);
and UO_281 (O_281,N_4915,N_4441);
xor UO_282 (O_282,N_4604,N_4059);
nor UO_283 (O_283,N_4942,N_4910);
nand UO_284 (O_284,N_4363,N_4841);
nand UO_285 (O_285,N_4878,N_4319);
or UO_286 (O_286,N_4288,N_4880);
and UO_287 (O_287,N_4871,N_4735);
or UO_288 (O_288,N_4775,N_4140);
nor UO_289 (O_289,N_4727,N_4368);
and UO_290 (O_290,N_4832,N_4573);
nor UO_291 (O_291,N_4150,N_4558);
nor UO_292 (O_292,N_4570,N_4920);
nand UO_293 (O_293,N_4073,N_4951);
and UO_294 (O_294,N_4676,N_4266);
or UO_295 (O_295,N_4890,N_4394);
xor UO_296 (O_296,N_4522,N_4194);
or UO_297 (O_297,N_4108,N_4174);
or UO_298 (O_298,N_4501,N_4699);
nor UO_299 (O_299,N_4469,N_4658);
nand UO_300 (O_300,N_4747,N_4433);
or UO_301 (O_301,N_4148,N_4470);
nor UO_302 (O_302,N_4009,N_4465);
nand UO_303 (O_303,N_4379,N_4539);
and UO_304 (O_304,N_4582,N_4478);
nand UO_305 (O_305,N_4982,N_4552);
and UO_306 (O_306,N_4640,N_4797);
nor UO_307 (O_307,N_4625,N_4621);
and UO_308 (O_308,N_4169,N_4821);
nand UO_309 (O_309,N_4384,N_4442);
xnor UO_310 (O_310,N_4293,N_4892);
xor UO_311 (O_311,N_4641,N_4277);
nor UO_312 (O_312,N_4652,N_4244);
nand UO_313 (O_313,N_4198,N_4771);
nand UO_314 (O_314,N_4601,N_4521);
and UO_315 (O_315,N_4926,N_4526);
and UO_316 (O_316,N_4495,N_4345);
and UO_317 (O_317,N_4228,N_4756);
or UO_318 (O_318,N_4044,N_4808);
nand UO_319 (O_319,N_4629,N_4152);
or UO_320 (O_320,N_4610,N_4429);
nor UO_321 (O_321,N_4392,N_4022);
xor UO_322 (O_322,N_4134,N_4686);
and UO_323 (O_323,N_4548,N_4732);
and UO_324 (O_324,N_4386,N_4806);
and UO_325 (O_325,N_4937,N_4248);
xor UO_326 (O_326,N_4882,N_4201);
and UO_327 (O_327,N_4360,N_4158);
nor UO_328 (O_328,N_4483,N_4063);
nor UO_329 (O_329,N_4886,N_4507);
or UO_330 (O_330,N_4896,N_4385);
or UO_331 (O_331,N_4217,N_4060);
nand UO_332 (O_332,N_4179,N_4024);
nor UO_333 (O_333,N_4116,N_4794);
nand UO_334 (O_334,N_4111,N_4520);
nand UO_335 (O_335,N_4984,N_4006);
nor UO_336 (O_336,N_4932,N_4839);
xor UO_337 (O_337,N_4166,N_4664);
and UO_338 (O_338,N_4542,N_4774);
and UO_339 (O_339,N_4154,N_4532);
nand UO_340 (O_340,N_4655,N_4673);
nor UO_341 (O_341,N_4199,N_4894);
nand UO_342 (O_342,N_4147,N_4349);
or UO_343 (O_343,N_4761,N_4817);
and UO_344 (O_344,N_4448,N_4336);
nand UO_345 (O_345,N_4133,N_4961);
nor UO_346 (O_346,N_4161,N_4940);
or UO_347 (O_347,N_4065,N_4391);
nor UO_348 (O_348,N_4721,N_4335);
nor UO_349 (O_349,N_4132,N_4739);
and UO_350 (O_350,N_4516,N_4935);
and UO_351 (O_351,N_4657,N_4207);
and UO_352 (O_352,N_4136,N_4965);
nand UO_353 (O_353,N_4546,N_4627);
or UO_354 (O_354,N_4950,N_4983);
nor UO_355 (O_355,N_4922,N_4192);
and UO_356 (O_356,N_4491,N_4447);
and UO_357 (O_357,N_4064,N_4082);
or UO_358 (O_358,N_4577,N_4028);
and UO_359 (O_359,N_4079,N_4324);
or UO_360 (O_360,N_4565,N_4239);
nor UO_361 (O_361,N_4814,N_4226);
nor UO_362 (O_362,N_4118,N_4767);
and UO_363 (O_363,N_4617,N_4772);
xor UO_364 (O_364,N_4626,N_4583);
nor UO_365 (O_365,N_4903,N_4274);
nand UO_366 (O_366,N_4811,N_4220);
nor UO_367 (O_367,N_4599,N_4622);
nor UO_368 (O_368,N_4370,N_4663);
and UO_369 (O_369,N_4309,N_4021);
and UO_370 (O_370,N_4691,N_4513);
or UO_371 (O_371,N_4089,N_4388);
nand UO_372 (O_372,N_4904,N_4338);
nand UO_373 (O_373,N_4242,N_4860);
or UO_374 (O_374,N_4102,N_4831);
and UO_375 (O_375,N_4373,N_4974);
nor UO_376 (O_376,N_4785,N_4088);
or UO_377 (O_377,N_4643,N_4139);
or UO_378 (O_378,N_4197,N_4813);
nor UO_379 (O_379,N_4430,N_4435);
nor UO_380 (O_380,N_4225,N_4375);
nor UO_381 (O_381,N_4683,N_4579);
or UO_382 (O_382,N_4650,N_4874);
and UO_383 (O_383,N_4607,N_4084);
or UO_384 (O_384,N_4072,N_4704);
or UO_385 (O_385,N_4568,N_4667);
or UO_386 (O_386,N_4695,N_4677);
and UO_387 (O_387,N_4613,N_4825);
nor UO_388 (O_388,N_4891,N_4333);
nor UO_389 (O_389,N_4496,N_4647);
and UO_390 (O_390,N_4555,N_4400);
and UO_391 (O_391,N_4688,N_4467);
nor UO_392 (O_392,N_4090,N_4672);
nor UO_393 (O_393,N_4911,N_4693);
nor UO_394 (O_394,N_4490,N_4889);
nand UO_395 (O_395,N_4755,N_4754);
or UO_396 (O_396,N_4620,N_4355);
and UO_397 (O_397,N_4826,N_4407);
or UO_398 (O_398,N_4105,N_4145);
nand UO_399 (O_399,N_4395,N_4544);
and UO_400 (O_400,N_4115,N_4623);
and UO_401 (O_401,N_4117,N_4608);
or UO_402 (O_402,N_4713,N_4712);
nor UO_403 (O_403,N_4010,N_4545);
nand UO_404 (O_404,N_4576,N_4858);
and UO_405 (O_405,N_4233,N_4053);
and UO_406 (O_406,N_4104,N_4867);
and UO_407 (O_407,N_4339,N_4877);
and UO_408 (O_408,N_4040,N_4305);
nor UO_409 (O_409,N_4590,N_4908);
nor UO_410 (O_410,N_4616,N_4737);
nand UO_411 (O_411,N_4661,N_4804);
and UO_412 (O_412,N_4540,N_4492);
nand UO_413 (O_413,N_4870,N_4221);
and UO_414 (O_414,N_4725,N_4799);
nor UO_415 (O_415,N_4455,N_4234);
and UO_416 (O_416,N_4026,N_4167);
and UO_417 (O_417,N_4107,N_4163);
nor UO_418 (O_418,N_4838,N_4164);
xnor UO_419 (O_419,N_4692,N_4511);
nand UO_420 (O_420,N_4434,N_4571);
nor UO_421 (O_421,N_4176,N_4697);
and UO_422 (O_422,N_4949,N_4968);
nand UO_423 (O_423,N_4829,N_4171);
nor UO_424 (O_424,N_4689,N_4316);
nor UO_425 (O_425,N_4656,N_4109);
or UO_426 (O_426,N_4512,N_4936);
nand UO_427 (O_427,N_4766,N_4126);
or UO_428 (O_428,N_4784,N_4212);
and UO_429 (O_429,N_4729,N_4557);
nor UO_430 (O_430,N_4189,N_4783);
nand UO_431 (O_431,N_4387,N_4417);
nor UO_432 (O_432,N_4760,N_4581);
xor UO_433 (O_433,N_4451,N_4793);
nor UO_434 (O_434,N_4879,N_4669);
and UO_435 (O_435,N_4954,N_4885);
or UO_436 (O_436,N_4554,N_4177);
nand UO_437 (O_437,N_4843,N_4382);
and UO_438 (O_438,N_4828,N_4287);
nand UO_439 (O_439,N_4253,N_4928);
or UO_440 (O_440,N_4012,N_4859);
nand UO_441 (O_441,N_4454,N_4702);
nor UO_442 (O_442,N_4247,N_4218);
nor UO_443 (O_443,N_4893,N_4256);
or UO_444 (O_444,N_4320,N_4660);
and UO_445 (O_445,N_4464,N_4270);
or UO_446 (O_446,N_4016,N_4505);
and UO_447 (O_447,N_4285,N_4314);
nand UO_448 (O_448,N_4537,N_4008);
nor UO_449 (O_449,N_4445,N_4588);
and UO_450 (O_450,N_4157,N_4972);
or UO_451 (O_451,N_4962,N_4644);
and UO_452 (O_452,N_4993,N_4235);
nor UO_453 (O_453,N_4671,N_4638);
or UO_454 (O_454,N_4902,N_4651);
and UO_455 (O_455,N_4204,N_4914);
and UO_456 (O_456,N_4606,N_4956);
nor UO_457 (O_457,N_4112,N_4129);
and UO_458 (O_458,N_4269,N_4905);
xnor UO_459 (O_459,N_4976,N_4792);
nand UO_460 (O_460,N_4515,N_4013);
and UO_461 (O_461,N_4019,N_4362);
xnor UO_462 (O_462,N_4875,N_4031);
nand UO_463 (O_463,N_4978,N_4034);
nor UO_464 (O_464,N_4802,N_4301);
and UO_465 (O_465,N_4271,N_4358);
nand UO_466 (O_466,N_4029,N_4268);
and UO_467 (O_467,N_4474,N_4930);
or UO_468 (O_468,N_4196,N_4734);
and UO_469 (O_469,N_4723,N_4415);
or UO_470 (O_470,N_4328,N_4585);
and UO_471 (O_471,N_4284,N_4372);
nor UO_472 (O_472,N_4321,N_4066);
or UO_473 (O_473,N_4810,N_4323);
nand UO_474 (O_474,N_4264,N_4100);
nor UO_475 (O_475,N_4603,N_4103);
and UO_476 (O_476,N_4714,N_4778);
and UO_477 (O_477,N_4479,N_4690);
nand UO_478 (O_478,N_4354,N_4240);
or UO_479 (O_479,N_4273,N_4229);
xor UO_480 (O_480,N_4728,N_4624);
or UO_481 (O_481,N_4456,N_4463);
nand UO_482 (O_482,N_4943,N_4062);
nand UO_483 (O_483,N_4979,N_4730);
or UO_484 (O_484,N_4769,N_4528);
or UO_485 (O_485,N_4156,N_4389);
nor UO_486 (O_486,N_4311,N_4888);
or UO_487 (O_487,N_4452,N_4411);
nor UO_488 (O_488,N_4446,N_4038);
or UO_489 (O_489,N_4897,N_4443);
nand UO_490 (O_490,N_4046,N_4939);
and UO_491 (O_491,N_4340,N_4497);
or UO_492 (O_492,N_4909,N_4436);
nand UO_493 (O_493,N_4185,N_4310);
and UO_494 (O_494,N_4206,N_4709);
nor UO_495 (O_495,N_4931,N_4946);
and UO_496 (O_496,N_4999,N_4572);
or UO_497 (O_497,N_4093,N_4110);
and UO_498 (O_498,N_4087,N_4014);
and UO_499 (O_499,N_4416,N_4222);
or UO_500 (O_500,N_4640,N_4197);
or UO_501 (O_501,N_4825,N_4195);
nor UO_502 (O_502,N_4983,N_4326);
xor UO_503 (O_503,N_4366,N_4279);
nor UO_504 (O_504,N_4612,N_4396);
or UO_505 (O_505,N_4664,N_4926);
or UO_506 (O_506,N_4329,N_4866);
nand UO_507 (O_507,N_4773,N_4126);
and UO_508 (O_508,N_4820,N_4866);
or UO_509 (O_509,N_4333,N_4186);
nor UO_510 (O_510,N_4444,N_4420);
and UO_511 (O_511,N_4461,N_4400);
and UO_512 (O_512,N_4644,N_4376);
nand UO_513 (O_513,N_4359,N_4858);
nand UO_514 (O_514,N_4969,N_4465);
nor UO_515 (O_515,N_4861,N_4308);
nand UO_516 (O_516,N_4343,N_4995);
nand UO_517 (O_517,N_4808,N_4555);
or UO_518 (O_518,N_4390,N_4264);
or UO_519 (O_519,N_4492,N_4476);
nand UO_520 (O_520,N_4155,N_4736);
or UO_521 (O_521,N_4942,N_4523);
nand UO_522 (O_522,N_4553,N_4812);
or UO_523 (O_523,N_4232,N_4076);
xor UO_524 (O_524,N_4701,N_4333);
or UO_525 (O_525,N_4088,N_4525);
nor UO_526 (O_526,N_4788,N_4596);
or UO_527 (O_527,N_4154,N_4605);
and UO_528 (O_528,N_4587,N_4636);
nand UO_529 (O_529,N_4394,N_4101);
nand UO_530 (O_530,N_4223,N_4019);
nand UO_531 (O_531,N_4443,N_4134);
or UO_532 (O_532,N_4532,N_4076);
nand UO_533 (O_533,N_4888,N_4429);
and UO_534 (O_534,N_4205,N_4230);
nor UO_535 (O_535,N_4308,N_4361);
or UO_536 (O_536,N_4253,N_4145);
nor UO_537 (O_537,N_4897,N_4051);
or UO_538 (O_538,N_4873,N_4011);
or UO_539 (O_539,N_4541,N_4677);
nor UO_540 (O_540,N_4556,N_4041);
nand UO_541 (O_541,N_4068,N_4000);
and UO_542 (O_542,N_4922,N_4165);
nor UO_543 (O_543,N_4644,N_4360);
and UO_544 (O_544,N_4535,N_4322);
nor UO_545 (O_545,N_4577,N_4811);
nor UO_546 (O_546,N_4458,N_4176);
nor UO_547 (O_547,N_4454,N_4818);
and UO_548 (O_548,N_4185,N_4120);
or UO_549 (O_549,N_4799,N_4364);
nor UO_550 (O_550,N_4176,N_4478);
and UO_551 (O_551,N_4093,N_4503);
nor UO_552 (O_552,N_4372,N_4691);
nand UO_553 (O_553,N_4426,N_4355);
or UO_554 (O_554,N_4650,N_4019);
or UO_555 (O_555,N_4025,N_4218);
nand UO_556 (O_556,N_4647,N_4401);
nand UO_557 (O_557,N_4041,N_4207);
and UO_558 (O_558,N_4195,N_4337);
nand UO_559 (O_559,N_4873,N_4356);
and UO_560 (O_560,N_4105,N_4535);
or UO_561 (O_561,N_4634,N_4795);
or UO_562 (O_562,N_4161,N_4979);
nand UO_563 (O_563,N_4131,N_4227);
nor UO_564 (O_564,N_4148,N_4962);
nor UO_565 (O_565,N_4174,N_4482);
or UO_566 (O_566,N_4274,N_4888);
or UO_567 (O_567,N_4655,N_4190);
nor UO_568 (O_568,N_4382,N_4011);
or UO_569 (O_569,N_4577,N_4007);
and UO_570 (O_570,N_4170,N_4161);
and UO_571 (O_571,N_4432,N_4846);
nor UO_572 (O_572,N_4789,N_4101);
or UO_573 (O_573,N_4618,N_4744);
nor UO_574 (O_574,N_4899,N_4654);
nor UO_575 (O_575,N_4350,N_4130);
and UO_576 (O_576,N_4114,N_4700);
or UO_577 (O_577,N_4356,N_4096);
and UO_578 (O_578,N_4673,N_4275);
and UO_579 (O_579,N_4272,N_4156);
nand UO_580 (O_580,N_4847,N_4857);
and UO_581 (O_581,N_4168,N_4706);
and UO_582 (O_582,N_4610,N_4528);
and UO_583 (O_583,N_4223,N_4054);
or UO_584 (O_584,N_4419,N_4472);
nand UO_585 (O_585,N_4628,N_4916);
nor UO_586 (O_586,N_4526,N_4728);
nand UO_587 (O_587,N_4375,N_4307);
nand UO_588 (O_588,N_4586,N_4295);
nor UO_589 (O_589,N_4306,N_4727);
or UO_590 (O_590,N_4876,N_4762);
nor UO_591 (O_591,N_4122,N_4802);
nor UO_592 (O_592,N_4958,N_4725);
and UO_593 (O_593,N_4766,N_4031);
nor UO_594 (O_594,N_4716,N_4113);
nand UO_595 (O_595,N_4747,N_4267);
nand UO_596 (O_596,N_4406,N_4887);
nand UO_597 (O_597,N_4981,N_4333);
nor UO_598 (O_598,N_4727,N_4716);
xnor UO_599 (O_599,N_4561,N_4856);
nor UO_600 (O_600,N_4874,N_4351);
or UO_601 (O_601,N_4555,N_4279);
or UO_602 (O_602,N_4648,N_4458);
nand UO_603 (O_603,N_4974,N_4055);
and UO_604 (O_604,N_4299,N_4721);
or UO_605 (O_605,N_4302,N_4965);
nor UO_606 (O_606,N_4484,N_4022);
or UO_607 (O_607,N_4762,N_4779);
nor UO_608 (O_608,N_4386,N_4031);
and UO_609 (O_609,N_4104,N_4998);
nand UO_610 (O_610,N_4347,N_4607);
and UO_611 (O_611,N_4013,N_4387);
nand UO_612 (O_612,N_4911,N_4018);
and UO_613 (O_613,N_4315,N_4934);
and UO_614 (O_614,N_4040,N_4757);
and UO_615 (O_615,N_4916,N_4064);
or UO_616 (O_616,N_4182,N_4605);
or UO_617 (O_617,N_4063,N_4553);
nor UO_618 (O_618,N_4015,N_4037);
nand UO_619 (O_619,N_4859,N_4968);
or UO_620 (O_620,N_4154,N_4798);
and UO_621 (O_621,N_4099,N_4692);
xnor UO_622 (O_622,N_4014,N_4478);
nor UO_623 (O_623,N_4392,N_4376);
nor UO_624 (O_624,N_4900,N_4400);
nand UO_625 (O_625,N_4901,N_4952);
and UO_626 (O_626,N_4557,N_4112);
and UO_627 (O_627,N_4364,N_4070);
nand UO_628 (O_628,N_4184,N_4705);
and UO_629 (O_629,N_4438,N_4381);
nand UO_630 (O_630,N_4960,N_4193);
nand UO_631 (O_631,N_4513,N_4669);
nor UO_632 (O_632,N_4708,N_4339);
and UO_633 (O_633,N_4868,N_4880);
and UO_634 (O_634,N_4561,N_4422);
nor UO_635 (O_635,N_4118,N_4217);
and UO_636 (O_636,N_4479,N_4582);
nand UO_637 (O_637,N_4854,N_4799);
nor UO_638 (O_638,N_4780,N_4385);
nand UO_639 (O_639,N_4612,N_4819);
nor UO_640 (O_640,N_4189,N_4183);
nor UO_641 (O_641,N_4087,N_4747);
or UO_642 (O_642,N_4388,N_4309);
or UO_643 (O_643,N_4547,N_4528);
xor UO_644 (O_644,N_4140,N_4329);
nor UO_645 (O_645,N_4988,N_4317);
or UO_646 (O_646,N_4754,N_4012);
or UO_647 (O_647,N_4823,N_4095);
nand UO_648 (O_648,N_4075,N_4958);
nand UO_649 (O_649,N_4194,N_4251);
or UO_650 (O_650,N_4701,N_4951);
nor UO_651 (O_651,N_4801,N_4815);
nand UO_652 (O_652,N_4708,N_4735);
or UO_653 (O_653,N_4235,N_4876);
and UO_654 (O_654,N_4804,N_4504);
and UO_655 (O_655,N_4846,N_4471);
and UO_656 (O_656,N_4654,N_4017);
and UO_657 (O_657,N_4305,N_4672);
nor UO_658 (O_658,N_4484,N_4226);
and UO_659 (O_659,N_4882,N_4855);
nor UO_660 (O_660,N_4284,N_4831);
or UO_661 (O_661,N_4503,N_4320);
and UO_662 (O_662,N_4265,N_4363);
nand UO_663 (O_663,N_4773,N_4232);
or UO_664 (O_664,N_4233,N_4583);
nor UO_665 (O_665,N_4279,N_4793);
nor UO_666 (O_666,N_4195,N_4937);
nor UO_667 (O_667,N_4099,N_4070);
and UO_668 (O_668,N_4394,N_4161);
nor UO_669 (O_669,N_4597,N_4681);
or UO_670 (O_670,N_4278,N_4287);
xor UO_671 (O_671,N_4932,N_4973);
or UO_672 (O_672,N_4369,N_4836);
nand UO_673 (O_673,N_4201,N_4629);
and UO_674 (O_674,N_4437,N_4255);
and UO_675 (O_675,N_4657,N_4011);
or UO_676 (O_676,N_4963,N_4355);
nand UO_677 (O_677,N_4076,N_4022);
nand UO_678 (O_678,N_4019,N_4003);
and UO_679 (O_679,N_4191,N_4997);
nor UO_680 (O_680,N_4102,N_4714);
xor UO_681 (O_681,N_4154,N_4792);
nor UO_682 (O_682,N_4400,N_4410);
or UO_683 (O_683,N_4923,N_4516);
and UO_684 (O_684,N_4613,N_4373);
and UO_685 (O_685,N_4990,N_4731);
nand UO_686 (O_686,N_4498,N_4002);
or UO_687 (O_687,N_4834,N_4729);
and UO_688 (O_688,N_4200,N_4913);
or UO_689 (O_689,N_4608,N_4018);
or UO_690 (O_690,N_4545,N_4800);
or UO_691 (O_691,N_4301,N_4977);
nand UO_692 (O_692,N_4369,N_4407);
or UO_693 (O_693,N_4518,N_4672);
nand UO_694 (O_694,N_4896,N_4061);
nor UO_695 (O_695,N_4397,N_4586);
or UO_696 (O_696,N_4054,N_4151);
or UO_697 (O_697,N_4471,N_4592);
nand UO_698 (O_698,N_4367,N_4059);
nand UO_699 (O_699,N_4085,N_4365);
xnor UO_700 (O_700,N_4497,N_4085);
and UO_701 (O_701,N_4437,N_4946);
xnor UO_702 (O_702,N_4739,N_4050);
nand UO_703 (O_703,N_4206,N_4912);
and UO_704 (O_704,N_4338,N_4303);
nor UO_705 (O_705,N_4831,N_4072);
nor UO_706 (O_706,N_4538,N_4650);
and UO_707 (O_707,N_4039,N_4240);
nor UO_708 (O_708,N_4472,N_4734);
or UO_709 (O_709,N_4164,N_4576);
nand UO_710 (O_710,N_4094,N_4479);
nand UO_711 (O_711,N_4251,N_4680);
and UO_712 (O_712,N_4536,N_4957);
or UO_713 (O_713,N_4425,N_4644);
nor UO_714 (O_714,N_4587,N_4033);
and UO_715 (O_715,N_4100,N_4075);
nor UO_716 (O_716,N_4707,N_4039);
nand UO_717 (O_717,N_4582,N_4826);
or UO_718 (O_718,N_4759,N_4410);
nand UO_719 (O_719,N_4500,N_4503);
and UO_720 (O_720,N_4520,N_4750);
nand UO_721 (O_721,N_4521,N_4883);
or UO_722 (O_722,N_4643,N_4487);
or UO_723 (O_723,N_4696,N_4934);
nor UO_724 (O_724,N_4405,N_4404);
nor UO_725 (O_725,N_4309,N_4393);
nor UO_726 (O_726,N_4652,N_4503);
nand UO_727 (O_727,N_4615,N_4726);
nand UO_728 (O_728,N_4251,N_4171);
nor UO_729 (O_729,N_4941,N_4746);
nand UO_730 (O_730,N_4188,N_4395);
nor UO_731 (O_731,N_4261,N_4302);
nor UO_732 (O_732,N_4721,N_4439);
nor UO_733 (O_733,N_4764,N_4890);
or UO_734 (O_734,N_4529,N_4369);
nand UO_735 (O_735,N_4665,N_4888);
nor UO_736 (O_736,N_4390,N_4636);
and UO_737 (O_737,N_4115,N_4023);
and UO_738 (O_738,N_4484,N_4209);
and UO_739 (O_739,N_4289,N_4261);
and UO_740 (O_740,N_4680,N_4556);
and UO_741 (O_741,N_4446,N_4319);
xnor UO_742 (O_742,N_4117,N_4887);
or UO_743 (O_743,N_4495,N_4470);
nor UO_744 (O_744,N_4730,N_4415);
nand UO_745 (O_745,N_4501,N_4772);
nand UO_746 (O_746,N_4055,N_4187);
or UO_747 (O_747,N_4936,N_4099);
nand UO_748 (O_748,N_4806,N_4146);
nor UO_749 (O_749,N_4356,N_4016);
or UO_750 (O_750,N_4301,N_4282);
or UO_751 (O_751,N_4908,N_4111);
or UO_752 (O_752,N_4683,N_4820);
and UO_753 (O_753,N_4539,N_4609);
and UO_754 (O_754,N_4580,N_4610);
nand UO_755 (O_755,N_4393,N_4148);
nor UO_756 (O_756,N_4560,N_4327);
nor UO_757 (O_757,N_4122,N_4241);
nor UO_758 (O_758,N_4637,N_4963);
or UO_759 (O_759,N_4396,N_4382);
nor UO_760 (O_760,N_4066,N_4777);
and UO_761 (O_761,N_4601,N_4153);
nand UO_762 (O_762,N_4067,N_4124);
or UO_763 (O_763,N_4442,N_4802);
or UO_764 (O_764,N_4043,N_4533);
and UO_765 (O_765,N_4259,N_4905);
or UO_766 (O_766,N_4354,N_4479);
or UO_767 (O_767,N_4593,N_4619);
nor UO_768 (O_768,N_4695,N_4976);
or UO_769 (O_769,N_4044,N_4380);
nor UO_770 (O_770,N_4691,N_4323);
and UO_771 (O_771,N_4777,N_4766);
nand UO_772 (O_772,N_4735,N_4678);
or UO_773 (O_773,N_4673,N_4331);
and UO_774 (O_774,N_4425,N_4455);
or UO_775 (O_775,N_4429,N_4284);
nor UO_776 (O_776,N_4165,N_4060);
nor UO_777 (O_777,N_4031,N_4451);
xor UO_778 (O_778,N_4735,N_4544);
nor UO_779 (O_779,N_4944,N_4268);
nand UO_780 (O_780,N_4287,N_4130);
and UO_781 (O_781,N_4205,N_4944);
nor UO_782 (O_782,N_4528,N_4126);
nor UO_783 (O_783,N_4420,N_4246);
nand UO_784 (O_784,N_4027,N_4022);
nand UO_785 (O_785,N_4060,N_4018);
nor UO_786 (O_786,N_4846,N_4581);
and UO_787 (O_787,N_4759,N_4564);
or UO_788 (O_788,N_4289,N_4970);
nand UO_789 (O_789,N_4164,N_4917);
and UO_790 (O_790,N_4018,N_4500);
or UO_791 (O_791,N_4529,N_4617);
nor UO_792 (O_792,N_4139,N_4559);
nand UO_793 (O_793,N_4610,N_4849);
nor UO_794 (O_794,N_4442,N_4203);
nand UO_795 (O_795,N_4796,N_4755);
or UO_796 (O_796,N_4957,N_4606);
or UO_797 (O_797,N_4207,N_4539);
or UO_798 (O_798,N_4941,N_4747);
or UO_799 (O_799,N_4185,N_4804);
and UO_800 (O_800,N_4129,N_4167);
nand UO_801 (O_801,N_4162,N_4175);
nand UO_802 (O_802,N_4764,N_4791);
nand UO_803 (O_803,N_4666,N_4952);
and UO_804 (O_804,N_4987,N_4955);
and UO_805 (O_805,N_4771,N_4782);
nor UO_806 (O_806,N_4629,N_4991);
nor UO_807 (O_807,N_4946,N_4132);
and UO_808 (O_808,N_4249,N_4530);
or UO_809 (O_809,N_4487,N_4139);
and UO_810 (O_810,N_4433,N_4812);
xnor UO_811 (O_811,N_4741,N_4507);
nand UO_812 (O_812,N_4064,N_4936);
nor UO_813 (O_813,N_4287,N_4671);
nor UO_814 (O_814,N_4234,N_4616);
and UO_815 (O_815,N_4925,N_4145);
nand UO_816 (O_816,N_4451,N_4267);
nor UO_817 (O_817,N_4182,N_4288);
nor UO_818 (O_818,N_4808,N_4205);
nand UO_819 (O_819,N_4250,N_4645);
and UO_820 (O_820,N_4143,N_4914);
nor UO_821 (O_821,N_4867,N_4311);
xnor UO_822 (O_822,N_4636,N_4622);
and UO_823 (O_823,N_4287,N_4565);
nor UO_824 (O_824,N_4801,N_4495);
and UO_825 (O_825,N_4280,N_4024);
nand UO_826 (O_826,N_4969,N_4614);
or UO_827 (O_827,N_4021,N_4470);
nand UO_828 (O_828,N_4492,N_4287);
nand UO_829 (O_829,N_4993,N_4325);
or UO_830 (O_830,N_4655,N_4170);
xnor UO_831 (O_831,N_4381,N_4495);
or UO_832 (O_832,N_4959,N_4669);
nor UO_833 (O_833,N_4086,N_4570);
nor UO_834 (O_834,N_4847,N_4298);
and UO_835 (O_835,N_4701,N_4051);
or UO_836 (O_836,N_4992,N_4850);
xnor UO_837 (O_837,N_4689,N_4908);
or UO_838 (O_838,N_4903,N_4621);
nor UO_839 (O_839,N_4366,N_4964);
and UO_840 (O_840,N_4966,N_4723);
or UO_841 (O_841,N_4044,N_4326);
nand UO_842 (O_842,N_4734,N_4281);
and UO_843 (O_843,N_4884,N_4655);
nor UO_844 (O_844,N_4625,N_4839);
and UO_845 (O_845,N_4316,N_4695);
nand UO_846 (O_846,N_4386,N_4857);
nand UO_847 (O_847,N_4736,N_4676);
nor UO_848 (O_848,N_4791,N_4188);
nor UO_849 (O_849,N_4825,N_4013);
nand UO_850 (O_850,N_4580,N_4399);
or UO_851 (O_851,N_4443,N_4015);
or UO_852 (O_852,N_4230,N_4525);
and UO_853 (O_853,N_4475,N_4572);
xnor UO_854 (O_854,N_4605,N_4022);
xor UO_855 (O_855,N_4853,N_4582);
or UO_856 (O_856,N_4445,N_4582);
nand UO_857 (O_857,N_4993,N_4122);
nor UO_858 (O_858,N_4353,N_4183);
and UO_859 (O_859,N_4634,N_4326);
nor UO_860 (O_860,N_4227,N_4556);
nor UO_861 (O_861,N_4296,N_4317);
or UO_862 (O_862,N_4389,N_4104);
and UO_863 (O_863,N_4000,N_4608);
and UO_864 (O_864,N_4396,N_4887);
nor UO_865 (O_865,N_4118,N_4988);
and UO_866 (O_866,N_4041,N_4208);
nand UO_867 (O_867,N_4053,N_4773);
and UO_868 (O_868,N_4233,N_4412);
nor UO_869 (O_869,N_4081,N_4565);
and UO_870 (O_870,N_4900,N_4970);
nand UO_871 (O_871,N_4739,N_4269);
nor UO_872 (O_872,N_4136,N_4938);
or UO_873 (O_873,N_4253,N_4871);
or UO_874 (O_874,N_4086,N_4215);
nor UO_875 (O_875,N_4190,N_4199);
or UO_876 (O_876,N_4565,N_4659);
nand UO_877 (O_877,N_4740,N_4701);
or UO_878 (O_878,N_4457,N_4441);
nand UO_879 (O_879,N_4535,N_4670);
nor UO_880 (O_880,N_4562,N_4875);
and UO_881 (O_881,N_4398,N_4051);
nand UO_882 (O_882,N_4911,N_4726);
nor UO_883 (O_883,N_4441,N_4672);
or UO_884 (O_884,N_4449,N_4481);
nand UO_885 (O_885,N_4032,N_4942);
nor UO_886 (O_886,N_4417,N_4811);
and UO_887 (O_887,N_4670,N_4238);
nor UO_888 (O_888,N_4110,N_4161);
nand UO_889 (O_889,N_4903,N_4348);
nor UO_890 (O_890,N_4279,N_4445);
or UO_891 (O_891,N_4092,N_4535);
nor UO_892 (O_892,N_4504,N_4838);
nor UO_893 (O_893,N_4503,N_4532);
nand UO_894 (O_894,N_4657,N_4719);
nand UO_895 (O_895,N_4747,N_4621);
and UO_896 (O_896,N_4109,N_4950);
nor UO_897 (O_897,N_4224,N_4240);
nand UO_898 (O_898,N_4801,N_4898);
and UO_899 (O_899,N_4371,N_4700);
or UO_900 (O_900,N_4403,N_4722);
nor UO_901 (O_901,N_4356,N_4825);
or UO_902 (O_902,N_4806,N_4179);
and UO_903 (O_903,N_4070,N_4058);
or UO_904 (O_904,N_4940,N_4388);
nor UO_905 (O_905,N_4710,N_4265);
and UO_906 (O_906,N_4391,N_4173);
and UO_907 (O_907,N_4918,N_4153);
nor UO_908 (O_908,N_4002,N_4346);
nand UO_909 (O_909,N_4964,N_4515);
and UO_910 (O_910,N_4091,N_4025);
or UO_911 (O_911,N_4323,N_4783);
or UO_912 (O_912,N_4276,N_4731);
nor UO_913 (O_913,N_4244,N_4941);
and UO_914 (O_914,N_4650,N_4469);
nor UO_915 (O_915,N_4726,N_4383);
nor UO_916 (O_916,N_4791,N_4212);
nor UO_917 (O_917,N_4328,N_4304);
nand UO_918 (O_918,N_4348,N_4263);
nor UO_919 (O_919,N_4680,N_4041);
nor UO_920 (O_920,N_4842,N_4257);
nor UO_921 (O_921,N_4992,N_4137);
nor UO_922 (O_922,N_4790,N_4940);
or UO_923 (O_923,N_4972,N_4602);
xnor UO_924 (O_924,N_4360,N_4001);
nor UO_925 (O_925,N_4028,N_4669);
nand UO_926 (O_926,N_4222,N_4642);
nand UO_927 (O_927,N_4622,N_4871);
nand UO_928 (O_928,N_4412,N_4471);
nand UO_929 (O_929,N_4078,N_4370);
nand UO_930 (O_930,N_4723,N_4075);
or UO_931 (O_931,N_4123,N_4144);
and UO_932 (O_932,N_4189,N_4775);
and UO_933 (O_933,N_4335,N_4620);
and UO_934 (O_934,N_4065,N_4658);
nand UO_935 (O_935,N_4252,N_4484);
and UO_936 (O_936,N_4515,N_4454);
and UO_937 (O_937,N_4099,N_4904);
nor UO_938 (O_938,N_4441,N_4269);
nand UO_939 (O_939,N_4787,N_4871);
nor UO_940 (O_940,N_4974,N_4336);
nand UO_941 (O_941,N_4551,N_4745);
and UO_942 (O_942,N_4375,N_4370);
or UO_943 (O_943,N_4261,N_4918);
nor UO_944 (O_944,N_4524,N_4528);
or UO_945 (O_945,N_4021,N_4999);
nand UO_946 (O_946,N_4573,N_4857);
nor UO_947 (O_947,N_4420,N_4800);
nor UO_948 (O_948,N_4413,N_4647);
nor UO_949 (O_949,N_4713,N_4589);
and UO_950 (O_950,N_4287,N_4965);
and UO_951 (O_951,N_4059,N_4490);
nand UO_952 (O_952,N_4046,N_4041);
and UO_953 (O_953,N_4086,N_4468);
and UO_954 (O_954,N_4464,N_4888);
or UO_955 (O_955,N_4650,N_4629);
nor UO_956 (O_956,N_4241,N_4172);
xor UO_957 (O_957,N_4624,N_4956);
nand UO_958 (O_958,N_4082,N_4738);
and UO_959 (O_959,N_4988,N_4357);
nand UO_960 (O_960,N_4414,N_4561);
or UO_961 (O_961,N_4895,N_4687);
and UO_962 (O_962,N_4617,N_4672);
or UO_963 (O_963,N_4484,N_4140);
nor UO_964 (O_964,N_4524,N_4399);
or UO_965 (O_965,N_4672,N_4445);
nand UO_966 (O_966,N_4859,N_4489);
xor UO_967 (O_967,N_4348,N_4106);
nor UO_968 (O_968,N_4347,N_4737);
or UO_969 (O_969,N_4418,N_4239);
nor UO_970 (O_970,N_4874,N_4832);
and UO_971 (O_971,N_4043,N_4685);
nand UO_972 (O_972,N_4470,N_4356);
and UO_973 (O_973,N_4699,N_4320);
or UO_974 (O_974,N_4415,N_4285);
or UO_975 (O_975,N_4740,N_4013);
nand UO_976 (O_976,N_4523,N_4921);
and UO_977 (O_977,N_4113,N_4531);
nand UO_978 (O_978,N_4964,N_4870);
and UO_979 (O_979,N_4348,N_4808);
nand UO_980 (O_980,N_4937,N_4275);
nand UO_981 (O_981,N_4374,N_4940);
or UO_982 (O_982,N_4322,N_4590);
and UO_983 (O_983,N_4115,N_4108);
or UO_984 (O_984,N_4740,N_4167);
or UO_985 (O_985,N_4012,N_4929);
xnor UO_986 (O_986,N_4074,N_4202);
nand UO_987 (O_987,N_4336,N_4996);
and UO_988 (O_988,N_4937,N_4737);
or UO_989 (O_989,N_4442,N_4191);
nor UO_990 (O_990,N_4550,N_4411);
nor UO_991 (O_991,N_4658,N_4756);
nand UO_992 (O_992,N_4080,N_4757);
or UO_993 (O_993,N_4014,N_4032);
or UO_994 (O_994,N_4078,N_4185);
nand UO_995 (O_995,N_4380,N_4245);
and UO_996 (O_996,N_4696,N_4544);
or UO_997 (O_997,N_4056,N_4018);
nand UO_998 (O_998,N_4680,N_4241);
or UO_999 (O_999,N_4776,N_4989);
endmodule