module basic_3000_30000_3500_20_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nand U0 (N_0,In_407,In_1362);
nor U1 (N_1,In_2028,In_1368);
or U2 (N_2,In_746,In_1543);
nand U3 (N_3,In_654,In_2623);
nor U4 (N_4,In_1838,In_2600);
xor U5 (N_5,In_1483,In_667);
nand U6 (N_6,In_688,In_602);
and U7 (N_7,In_1111,In_1952);
and U8 (N_8,In_2892,In_2542);
nand U9 (N_9,In_2449,In_159);
nor U10 (N_10,In_1125,In_981);
nor U11 (N_11,In_2911,In_2766);
nand U12 (N_12,In_2561,In_1786);
xor U13 (N_13,In_1434,In_2876);
or U14 (N_14,In_2953,In_2511);
xor U15 (N_15,In_1373,In_1037);
xor U16 (N_16,In_1470,In_331);
nand U17 (N_17,In_2964,In_709);
xnor U18 (N_18,In_2965,In_2414);
or U19 (N_19,In_2042,In_1767);
and U20 (N_20,In_965,In_2825);
nand U21 (N_21,In_1311,In_1671);
and U22 (N_22,In_2852,In_604);
nand U23 (N_23,In_2612,In_2264);
or U24 (N_24,In_1666,In_1757);
or U25 (N_25,In_176,In_2898);
or U26 (N_26,In_770,In_1741);
nand U27 (N_27,In_1206,In_1508);
and U28 (N_28,In_567,In_2993);
or U29 (N_29,In_628,In_2386);
or U30 (N_30,In_564,In_1637);
and U31 (N_31,In_2118,In_2323);
xnor U32 (N_32,In_2605,In_2249);
or U33 (N_33,In_2236,In_150);
nand U34 (N_34,In_2361,In_361);
xor U35 (N_35,In_608,In_1879);
nand U36 (N_36,In_2270,In_134);
xnor U37 (N_37,In_2975,In_525);
or U38 (N_38,In_2244,In_415);
and U39 (N_39,In_2639,In_1980);
or U40 (N_40,In_98,In_1289);
or U41 (N_41,In_1657,In_863);
nand U42 (N_42,In_199,In_2126);
or U43 (N_43,In_551,In_1673);
and U44 (N_44,In_1572,In_2063);
or U45 (N_45,In_1444,In_218);
or U46 (N_46,In_1376,In_2913);
or U47 (N_47,In_804,In_2266);
or U48 (N_48,In_1151,In_1506);
or U49 (N_49,In_1611,In_231);
and U50 (N_50,In_885,In_2645);
nand U51 (N_51,In_2219,In_546);
or U52 (N_52,In_2690,In_1617);
nand U53 (N_53,In_2676,In_1220);
nor U54 (N_54,In_2874,In_897);
nor U55 (N_55,In_130,In_332);
xnor U56 (N_56,In_1387,In_1453);
nand U57 (N_57,In_2989,In_831);
nand U58 (N_58,In_1643,In_577);
nor U59 (N_59,In_1842,In_1112);
nand U60 (N_60,In_1045,In_2527);
xnor U61 (N_61,In_2159,In_994);
and U62 (N_62,In_521,In_1171);
xor U63 (N_63,In_1312,In_2685);
or U64 (N_64,In_185,In_8);
xor U65 (N_65,In_68,In_275);
nor U66 (N_66,In_341,In_2135);
and U67 (N_67,In_1441,In_623);
and U68 (N_68,In_1272,In_168);
and U69 (N_69,In_1718,In_737);
and U70 (N_70,In_910,In_1050);
or U71 (N_71,In_779,In_2771);
nand U72 (N_72,In_1987,In_1533);
nand U73 (N_73,In_3,In_2954);
xor U74 (N_74,In_310,In_1128);
nand U75 (N_75,In_2785,In_610);
or U76 (N_76,In_146,In_2959);
and U77 (N_77,In_1080,In_2116);
xor U78 (N_78,In_1923,In_2584);
nor U79 (N_79,In_1925,In_2802);
nor U80 (N_80,In_1394,In_834);
nand U81 (N_81,In_1915,In_1325);
and U82 (N_82,In_201,In_340);
and U83 (N_83,In_760,In_1509);
or U84 (N_84,In_780,In_1365);
nand U85 (N_85,In_1450,In_74);
and U86 (N_86,In_1714,In_2501);
and U87 (N_87,In_1680,In_1831);
xor U88 (N_88,In_1343,In_2209);
nor U89 (N_89,In_1263,In_616);
nor U90 (N_90,In_1740,In_225);
or U91 (N_91,In_2640,In_2165);
nor U92 (N_92,In_1809,In_2352);
xnor U93 (N_93,In_2416,In_1224);
nor U94 (N_94,In_850,In_2522);
nand U95 (N_95,In_2288,In_508);
and U96 (N_96,In_1770,In_686);
or U97 (N_97,In_769,In_1722);
and U98 (N_98,In_1492,In_45);
nand U99 (N_99,In_2154,In_2260);
nor U100 (N_100,In_383,In_1735);
nand U101 (N_101,In_2454,In_2458);
and U102 (N_102,In_1203,In_2859);
nor U103 (N_103,In_44,In_43);
nand U104 (N_104,In_1535,In_1101);
nor U105 (N_105,In_1116,In_2908);
and U106 (N_106,In_985,In_999);
nand U107 (N_107,In_1356,In_2936);
xor U108 (N_108,In_1321,In_2553);
nand U109 (N_109,In_2546,In_299);
and U110 (N_110,In_1397,In_1186);
nor U111 (N_111,In_1908,In_2504);
xnor U112 (N_112,In_1213,In_2929);
nor U113 (N_113,In_1609,In_2784);
nand U114 (N_114,In_2935,In_1235);
and U115 (N_115,In_1445,In_2549);
and U116 (N_116,In_1059,In_856);
and U117 (N_117,In_33,In_2298);
nand U118 (N_118,In_2146,In_2337);
or U119 (N_119,In_1984,In_7);
xor U120 (N_120,In_465,In_2143);
or U121 (N_121,In_1703,In_528);
and U122 (N_122,In_24,In_1176);
nor U123 (N_123,In_660,In_783);
and U124 (N_124,In_1456,In_794);
and U125 (N_125,In_148,In_2652);
and U126 (N_126,In_1595,In_466);
xor U127 (N_127,In_2754,In_1791);
and U128 (N_128,In_2314,In_1032);
xnor U129 (N_129,In_1995,In_1184);
nand U130 (N_130,In_224,In_52);
and U131 (N_131,In_392,In_2560);
and U132 (N_132,In_365,In_219);
and U133 (N_133,In_474,In_249);
xnor U134 (N_134,In_427,In_1271);
nor U135 (N_135,In_881,In_1587);
nand U136 (N_136,In_2613,In_1709);
and U137 (N_137,In_2806,In_375);
xor U138 (N_138,In_1839,In_2494);
nor U139 (N_139,In_2174,In_2029);
and U140 (N_140,In_202,In_2114);
nand U141 (N_141,In_2712,In_689);
and U142 (N_142,In_1216,In_252);
or U143 (N_143,In_1275,In_1262);
nand U144 (N_144,In_644,In_2744);
or U145 (N_145,In_478,In_2144);
or U146 (N_146,In_1463,In_2666);
and U147 (N_147,In_2095,In_2719);
nor U148 (N_148,In_82,In_883);
nor U149 (N_149,In_101,In_2944);
xor U150 (N_150,In_898,In_2642);
and U151 (N_151,In_1241,In_380);
nor U152 (N_152,In_1253,In_2073);
nor U153 (N_153,In_1645,In_116);
and U154 (N_154,In_2117,In_2220);
xor U155 (N_155,In_2952,In_510);
xnor U156 (N_156,In_2302,In_2772);
and U157 (N_157,In_1433,In_2464);
nor U158 (N_158,In_1691,In_1968);
nor U159 (N_159,In_270,In_798);
xor U160 (N_160,In_2513,In_1355);
nand U161 (N_161,In_553,In_585);
xor U162 (N_162,In_1665,In_154);
and U163 (N_163,In_1641,In_1288);
xor U164 (N_164,In_2499,In_2239);
or U165 (N_165,In_129,In_1763);
xor U166 (N_166,In_2569,In_1187);
nand U167 (N_167,In_2577,In_1280);
or U168 (N_168,In_204,In_286);
nand U169 (N_169,In_2907,In_890);
or U170 (N_170,In_2216,In_980);
and U171 (N_171,In_1812,In_2069);
or U172 (N_172,In_127,In_1283);
or U173 (N_173,In_2364,In_895);
and U174 (N_174,In_1752,In_1282);
xnor U175 (N_175,In_2039,In_2787);
nor U176 (N_176,In_1008,In_2904);
nand U177 (N_177,In_1326,In_955);
nand U178 (N_178,In_200,In_2141);
nand U179 (N_179,In_2741,In_1823);
and U180 (N_180,In_912,In_1881);
xor U181 (N_181,In_2528,In_1378);
nor U182 (N_182,In_214,In_595);
xnor U183 (N_183,In_953,In_1640);
or U184 (N_184,In_701,In_1423);
nand U185 (N_185,In_2920,In_2503);
xnor U186 (N_186,In_1753,In_489);
or U187 (N_187,In_1999,In_1409);
nor U188 (N_188,In_1619,In_1692);
xor U189 (N_189,In_1464,In_1363);
nand U190 (N_190,In_2038,In_1148);
or U191 (N_191,In_2426,In_2424);
xnor U192 (N_192,In_1883,In_2123);
or U193 (N_193,In_2955,In_385);
nand U194 (N_194,In_2105,In_2196);
or U195 (N_195,In_2997,In_2148);
and U196 (N_196,In_555,In_2207);
xor U197 (N_197,In_77,In_2844);
nand U198 (N_198,In_2113,In_2795);
nand U199 (N_199,In_1511,In_2633);
nor U200 (N_200,In_86,In_533);
nand U201 (N_201,In_2273,In_2714);
nor U202 (N_202,In_964,In_1478);
xnor U203 (N_203,In_2774,In_736);
or U204 (N_204,In_989,In_789);
or U205 (N_205,In_936,In_396);
nand U206 (N_206,In_1079,In_1133);
nor U207 (N_207,In_2064,In_1315);
nand U208 (N_208,In_434,In_2218);
nor U209 (N_209,In_946,In_722);
or U210 (N_210,In_206,In_1331);
nor U211 (N_211,In_1199,In_303);
nand U212 (N_212,In_847,In_922);
nand U213 (N_213,In_1993,In_950);
nand U214 (N_214,In_1399,In_1904);
and U215 (N_215,In_2711,In_1481);
and U216 (N_216,In_824,In_2995);
and U217 (N_217,In_501,In_2444);
xor U218 (N_218,In_2329,In_1070);
nand U219 (N_219,In_1934,In_1574);
and U220 (N_220,In_2743,In_2206);
xnor U221 (N_221,In_70,In_2331);
xor U222 (N_222,In_1856,In_787);
xnor U223 (N_223,In_2791,In_2278);
and U224 (N_224,In_1996,In_2568);
or U225 (N_225,In_2415,In_2851);
nor U226 (N_226,In_2130,In_1559);
xor U227 (N_227,In_2099,In_2023);
or U228 (N_228,In_1690,In_1154);
nor U229 (N_229,In_1290,In_1335);
nor U230 (N_230,In_291,In_2003);
nand U231 (N_231,In_676,In_1351);
or U232 (N_232,In_2841,In_2439);
and U233 (N_233,In_2742,In_1446);
or U234 (N_234,In_1375,In_2518);
nor U235 (N_235,In_1784,In_947);
xor U236 (N_236,In_177,In_1018);
and U237 (N_237,In_1185,In_925);
nor U238 (N_238,In_125,In_2854);
nor U239 (N_239,In_2637,In_1062);
or U240 (N_240,In_2629,In_2779);
and U241 (N_241,In_2410,In_1226);
nor U242 (N_242,In_962,In_1850);
nor U243 (N_243,In_651,In_2375);
and U244 (N_244,In_142,In_638);
or U245 (N_245,In_2438,In_1916);
nor U246 (N_246,In_1575,In_2881);
and U247 (N_247,In_2659,In_2315);
or U248 (N_248,In_1975,In_740);
or U249 (N_249,In_1097,In_2926);
or U250 (N_250,In_468,In_2359);
and U251 (N_251,In_2463,In_2896);
xor U252 (N_252,In_1066,In_1346);
or U253 (N_253,In_2074,In_1500);
nor U254 (N_254,In_842,In_448);
and U255 (N_255,In_2624,In_2864);
nand U256 (N_256,In_1245,In_1659);
nand U257 (N_257,In_2412,In_2491);
and U258 (N_258,In_1540,In_592);
and U259 (N_259,In_1960,In_988);
nor U260 (N_260,In_558,In_290);
or U261 (N_261,In_145,In_1755);
xnor U262 (N_262,In_2047,In_1768);
nand U263 (N_263,In_2265,In_2473);
and U264 (N_264,In_2224,In_869);
and U265 (N_265,In_864,In_2334);
and U266 (N_266,In_2781,In_2340);
nor U267 (N_267,In_581,In_1821);
xor U268 (N_268,In_187,In_149);
and U269 (N_269,In_2222,In_128);
nand U270 (N_270,In_961,In_2902);
xor U271 (N_271,In_1953,In_2548);
nand U272 (N_272,In_2933,In_2187);
nand U273 (N_273,In_2271,In_636);
and U274 (N_274,In_2397,In_1268);
or U275 (N_275,In_1015,In_2835);
or U276 (N_276,In_951,In_2451);
nand U277 (N_277,In_2201,In_2258);
nand U278 (N_278,In_705,In_2713);
or U279 (N_279,In_1589,In_2969);
xnor U280 (N_280,In_1119,In_16);
and U281 (N_281,In_1900,In_265);
nand U282 (N_282,In_2515,In_1238);
nor U283 (N_283,In_1813,In_295);
xor U284 (N_284,In_1708,In_682);
nor U285 (N_285,In_47,In_21);
and U286 (N_286,In_1155,In_1939);
xnor U287 (N_287,In_2013,In_2958);
nand U288 (N_288,In_918,In_2643);
and U289 (N_289,In_1055,In_1026);
nand U290 (N_290,In_1239,In_1254);
xnor U291 (N_291,In_2660,In_900);
and U292 (N_292,In_515,In_2829);
and U293 (N_293,In_1902,In_634);
nor U294 (N_294,In_132,In_313);
xor U295 (N_295,In_1632,In_347);
or U296 (N_296,In_2050,In_1455);
or U297 (N_297,In_475,In_2689);
nor U298 (N_298,In_2554,In_233);
xnor U299 (N_299,In_2108,In_611);
and U300 (N_300,In_2846,In_828);
nand U301 (N_301,In_1158,In_697);
and U302 (N_302,In_2172,In_1568);
nor U303 (N_303,In_2836,In_2801);
and U304 (N_304,In_2371,In_2507);
xnor U305 (N_305,In_738,In_1117);
nand U306 (N_306,In_1894,In_1372);
nor U307 (N_307,In_2671,In_645);
xnor U308 (N_308,In_25,In_1005);
and U309 (N_309,In_2963,In_1033);
xor U310 (N_310,In_2310,In_668);
xnor U311 (N_311,In_580,In_2726);
xor U312 (N_312,In_2004,In_1525);
and U313 (N_313,In_2474,In_1800);
or U314 (N_314,In_2576,In_2931);
or U315 (N_315,In_1056,In_1863);
and U316 (N_316,In_1017,In_2888);
and U317 (N_317,In_2020,In_1488);
nor U318 (N_318,In_1006,In_1109);
nor U319 (N_319,In_986,In_1837);
and U320 (N_320,In_1501,In_405);
nor U321 (N_321,In_1108,In_762);
or U322 (N_322,In_719,In_2725);
nor U323 (N_323,In_2669,In_1638);
and U324 (N_324,In_1635,In_356);
nand U325 (N_325,In_140,In_1287);
and U326 (N_326,In_2609,In_1855);
nand U327 (N_327,In_2872,In_617);
or U328 (N_328,In_1320,In_2098);
xor U329 (N_329,In_839,In_213);
xnor U330 (N_330,In_973,In_1870);
and U331 (N_331,In_714,In_1053);
or U332 (N_332,In_2776,In_124);
nor U333 (N_333,In_1121,In_849);
nor U334 (N_334,In_493,In_472);
nor U335 (N_335,In_2692,In_2535);
nor U336 (N_336,In_2770,In_702);
or U337 (N_337,In_812,In_1776);
nor U338 (N_338,In_1964,In_857);
and U339 (N_339,In_2901,In_2031);
xnor U340 (N_340,In_1065,In_2919);
xor U341 (N_341,In_2565,In_2893);
nand U342 (N_342,In_215,In_180);
or U343 (N_343,In_2205,In_1796);
or U344 (N_344,In_2092,In_92);
and U345 (N_345,In_1240,In_2402);
or U346 (N_346,In_28,In_2573);
and U347 (N_347,In_2005,In_1307);
or U348 (N_348,In_2072,In_255);
and U349 (N_349,In_2909,In_350);
or U350 (N_350,In_2274,In_754);
nor U351 (N_351,In_819,In_30);
xnor U352 (N_352,In_1627,In_1247);
nor U353 (N_353,In_2152,In_613);
xor U354 (N_354,In_1260,In_1382);
nand U355 (N_355,In_1143,In_836);
nand U356 (N_356,In_2747,In_2296);
and U357 (N_357,In_2534,In_2080);
or U358 (N_358,In_244,In_2748);
or U359 (N_359,In_2827,In_748);
or U360 (N_360,In_19,In_2355);
nand U361 (N_361,In_552,In_576);
nor U362 (N_362,In_1270,In_1515);
and U363 (N_363,In_2760,In_1195);
or U364 (N_364,In_1428,In_502);
or U365 (N_365,In_2816,In_2435);
or U366 (N_366,In_438,In_1333);
and U367 (N_367,In_137,In_173);
and U368 (N_368,In_811,In_2523);
and U369 (N_369,In_1947,In_1404);
nand U370 (N_370,In_445,In_1829);
or U371 (N_371,In_1459,In_1771);
nor U372 (N_372,In_488,In_820);
xor U373 (N_373,In_1631,In_2032);
or U374 (N_374,In_2814,In_1107);
nand U375 (N_375,In_2567,In_1712);
xnor U376 (N_376,In_775,In_1798);
nor U377 (N_377,In_460,In_1432);
nand U378 (N_378,In_471,In_2231);
nor U379 (N_379,In_1221,In_85);
nor U380 (N_380,In_2532,In_987);
nand U381 (N_381,In_830,In_1291);
nor U382 (N_382,In_2243,In_578);
nand U383 (N_383,In_1590,In_2188);
nor U384 (N_384,In_2838,In_2650);
nor U385 (N_385,In_84,In_806);
and U386 (N_386,In_549,In_2440);
nor U387 (N_387,In_388,In_2022);
and U388 (N_388,In_2307,In_1664);
or U389 (N_389,In_2670,In_1648);
nand U390 (N_390,In_78,In_938);
and U391 (N_391,In_2750,In_1905);
nand U392 (N_392,In_2267,In_2471);
and U393 (N_393,In_523,In_278);
and U394 (N_394,In_2168,In_2653);
or U395 (N_395,In_1273,In_1988);
nor U396 (N_396,In_1046,In_2376);
xnor U397 (N_397,In_675,In_2984);
or U398 (N_398,In_54,In_2478);
xor U399 (N_399,In_2880,In_2543);
nor U400 (N_400,In_2456,In_2972);
and U401 (N_401,In_2336,In_2313);
nand U402 (N_402,In_1827,In_2661);
nand U403 (N_403,In_2807,In_2540);
nand U404 (N_404,In_2358,In_1435);
or U405 (N_405,In_1930,In_484);
and U406 (N_406,In_1679,In_2133);
nor U407 (N_407,In_657,In_404);
nand U408 (N_408,In_1292,In_2757);
xnor U409 (N_409,In_1913,In_1697);
xor U410 (N_410,In_2780,In_1063);
and U411 (N_411,In_196,In_2163);
and U412 (N_412,In_2192,In_1959);
nor U413 (N_413,In_1678,In_2715);
nand U414 (N_414,In_2385,In_1570);
nor U415 (N_415,In_155,In_1159);
xnor U416 (N_416,In_2716,In_1758);
nor U417 (N_417,In_1380,In_742);
or U418 (N_418,In_2990,In_707);
nand U419 (N_419,In_2813,In_2137);
nor U420 (N_420,In_1388,In_2710);
xor U421 (N_421,In_2539,In_756);
and U422 (N_422,In_309,In_1044);
or U423 (N_423,In_2894,In_2217);
nor U424 (N_424,In_969,In_2380);
xnor U425 (N_425,In_1249,In_1395);
nand U426 (N_426,In_2065,In_1192);
nand U427 (N_427,In_1420,In_242);
and U428 (N_428,In_113,In_2974);
and U429 (N_429,In_685,In_377);
or U430 (N_430,In_1139,In_1424);
and U431 (N_431,In_487,In_1867);
xnor U432 (N_432,In_2508,In_2142);
or U433 (N_433,In_933,In_178);
or U434 (N_434,In_2651,In_1707);
nor U435 (N_435,In_2982,In_635);
xnor U436 (N_436,In_2763,In_937);
xnor U437 (N_437,In_1096,In_1405);
or U438 (N_438,In_1512,In_503);
nand U439 (N_439,In_725,In_391);
or U440 (N_440,In_181,In_2398);
or U441 (N_441,In_1021,In_2976);
or U442 (N_442,In_693,In_855);
and U443 (N_443,In_1354,In_2865);
nor U444 (N_444,In_835,In_2160);
or U445 (N_445,In_626,In_2564);
nor U446 (N_446,In_1076,In_957);
nor U447 (N_447,In_522,In_183);
nand U448 (N_448,In_1799,In_111);
nor U449 (N_449,In_704,In_899);
and U450 (N_450,In_2550,In_2764);
and U451 (N_451,In_1539,In_1701);
or U452 (N_452,In_2899,In_1073);
nand U453 (N_453,In_1898,In_1009);
nand U454 (N_454,In_1985,In_1621);
nand U455 (N_455,In_357,In_2745);
and U456 (N_456,In_2060,In_2998);
nand U457 (N_457,In_2139,In_2405);
and U458 (N_458,In_2203,In_1327);
nor U459 (N_459,In_1149,In_678);
nand U460 (N_460,In_583,In_971);
nor U461 (N_461,In_1193,In_2103);
nand U462 (N_462,In_2996,In_2150);
nor U463 (N_463,In_582,In_1832);
nand U464 (N_464,In_1000,In_476);
xnor U465 (N_465,In_452,In_2756);
xnor U466 (N_466,In_1400,In_248);
and U467 (N_467,In_2082,In_572);
xnor U468 (N_468,In_803,In_1649);
xnor U469 (N_469,In_1379,In_399);
xor U470 (N_470,In_2918,In_2344);
or U471 (N_471,In_2408,In_94);
xor U472 (N_472,In_2610,In_1727);
or U473 (N_473,In_1979,In_858);
and U474 (N_474,In_2429,In_9);
and U475 (N_475,In_2434,In_538);
nor U476 (N_476,In_598,In_1647);
or U477 (N_477,In_417,In_376);
nand U478 (N_478,In_1974,In_6);
and U479 (N_479,In_2585,In_2379);
and U480 (N_480,In_103,In_734);
xor U481 (N_481,In_2370,In_2722);
nor U482 (N_482,In_2979,In_307);
and U483 (N_483,In_2932,In_603);
xnor U484 (N_484,In_1234,In_758);
xor U485 (N_485,In_2736,In_2420);
nand U486 (N_486,In_2285,In_18);
nand U487 (N_487,In_2182,In_2821);
nor U488 (N_488,In_109,In_1808);
xor U489 (N_489,In_2286,In_1804);
nand U490 (N_490,In_1507,In_2592);
nor U491 (N_491,In_1558,In_2240);
nor U492 (N_492,In_2393,In_1945);
nor U493 (N_493,In_490,In_2470);
nand U494 (N_494,In_1991,In_703);
xor U495 (N_495,In_588,In_300);
nand U496 (N_496,In_1505,In_963);
nor U497 (N_497,In_1480,In_845);
xor U498 (N_498,In_324,In_509);
nand U499 (N_499,In_1955,In_500);
xor U500 (N_500,In_1474,In_2915);
nand U501 (N_501,In_1510,In_123);
xnor U502 (N_502,In_954,In_2987);
and U503 (N_503,In_2891,In_526);
nand U504 (N_504,In_1717,In_2981);
nor U505 (N_505,In_669,In_1516);
or U506 (N_506,In_658,In_1495);
nand U507 (N_507,In_464,In_71);
xnor U508 (N_508,In_2247,In_1034);
and U509 (N_509,In_2111,In_2395);
xor U510 (N_510,In_2300,In_164);
or U511 (N_511,In_683,In_942);
or U512 (N_512,In_1135,In_2572);
xnor U513 (N_513,In_832,In_2563);
and U514 (N_514,In_1924,In_69);
nand U515 (N_515,In_1792,In_254);
xnor U516 (N_516,In_135,In_901);
nor U517 (N_517,In_83,In_88);
nor U518 (N_518,In_2696,In_1822);
and U519 (N_519,In_95,In_1725);
and U520 (N_520,In_1940,In_2242);
nor U521 (N_521,In_1316,In_1704);
or U522 (N_522,In_247,In_1921);
nor U523 (N_523,In_2619,In_777);
or U524 (N_524,In_2018,In_1416);
nor U525 (N_525,In_263,In_1145);
xor U526 (N_526,In_2594,In_0);
and U527 (N_527,In_1189,In_1820);
nand U528 (N_528,In_1713,In_1639);
xor U529 (N_529,In_2862,In_2967);
nand U530 (N_530,In_876,In_2903);
xor U531 (N_531,In_1183,In_2102);
nand U532 (N_532,In_1564,In_1897);
nor U533 (N_533,In_782,In_139);
nand U534 (N_534,In_649,In_1744);
or U535 (N_535,In_1676,In_1102);
or U536 (N_536,In_2253,In_1334);
or U537 (N_537,In_1603,In_2171);
or U538 (N_538,In_2204,In_1348);
nor U539 (N_539,In_622,In_198);
or U540 (N_540,In_2490,In_931);
or U541 (N_541,In_1401,In_2052);
or U542 (N_542,In_1598,In_469);
or U543 (N_543,In_1920,In_1297);
xor U544 (N_544,In_991,In_2043);
xor U545 (N_545,In_2962,In_1629);
xnor U546 (N_546,In_245,In_2055);
or U547 (N_547,In_2682,In_2277);
and U548 (N_548,In_393,In_1686);
nor U549 (N_549,In_1688,In_2820);
xnor U550 (N_550,In_413,In_1421);
and U551 (N_551,In_2718,In_1461);
nor U552 (N_552,In_210,In_878);
nor U553 (N_553,In_1557,In_2279);
nand U554 (N_554,In_998,In_720);
xnor U555 (N_555,In_36,In_739);
nor U556 (N_556,In_2447,In_2128);
nor U557 (N_557,In_2980,In_1957);
and U558 (N_558,In_1852,In_2037);
nand U559 (N_559,In_1140,In_1994);
or U560 (N_560,In_308,In_919);
xor U561 (N_561,In_410,In_2430);
and U562 (N_562,In_548,In_2132);
nand U563 (N_563,In_1774,In_1310);
nor U564 (N_564,In_32,In_2497);
nor U565 (N_565,In_1918,In_1522);
and U566 (N_566,In_2890,In_2783);
nand U567 (N_567,In_1257,In_2580);
nand U568 (N_568,In_1103,In_346);
nor U569 (N_569,In_1230,In_1242);
and U570 (N_570,In_1977,In_1653);
nor U571 (N_571,In_455,In_240);
and U572 (N_572,In_949,In_2647);
or U573 (N_573,In_241,In_1358);
and U574 (N_574,In_179,In_2994);
or U575 (N_575,In_2223,In_2949);
xnor U576 (N_576,In_2884,In_2051);
xnor U577 (N_577,In_90,In_436);
xor U578 (N_578,In_2459,In_1422);
and U579 (N_579,In_906,In_1550);
nand U580 (N_580,In_1431,In_1877);
nor U581 (N_581,In_2698,In_1276);
and U582 (N_582,In_11,In_1425);
nor U583 (N_583,In_2134,In_1759);
xor U584 (N_584,In_536,In_1514);
nor U585 (N_585,In_974,In_2401);
xnor U586 (N_586,In_2900,In_1663);
xor U587 (N_587,In_296,In_56);
or U588 (N_588,In_158,In_2895);
nand U589 (N_589,In_1551,In_2365);
nor U590 (N_590,In_1218,In_2593);
nand U591 (N_591,In_2632,In_1534);
nor U592 (N_592,In_710,In_945);
or U593 (N_593,In_2269,In_1085);
xor U594 (N_594,In_1137,In_1231);
xnor U595 (N_595,In_1296,In_236);
and U596 (N_596,In_708,In_2431);
nor U597 (N_597,In_2480,In_766);
nand U598 (N_598,In_2225,In_5);
or U599 (N_599,In_209,In_2200);
and U600 (N_600,In_1584,In_633);
or U601 (N_601,In_1266,In_208);
or U602 (N_602,In_1674,In_2934);
nor U603 (N_603,In_653,In_1857);
nor U604 (N_604,In_2662,In_102);
nand U605 (N_605,In_389,In_627);
or U606 (N_606,In_1178,In_1146);
xnor U607 (N_607,In_1197,In_2831);
or U608 (N_608,In_1020,In_1305);
and U609 (N_609,In_2818,In_1232);
and U610 (N_610,In_2011,In_909);
nand U611 (N_611,In_612,In_2916);
xor U612 (N_612,In_1024,In_799);
and U613 (N_613,In_2552,In_1208);
and U614 (N_614,In_15,In_2178);
xor U615 (N_615,In_2446,In_2012);
xnor U616 (N_616,In_1392,In_1599);
nor U617 (N_617,In_1886,In_2706);
and U618 (N_618,In_2001,In_1951);
nand U619 (N_619,In_1204,In_2484);
nand U620 (N_620,In_1489,In_2603);
nor U621 (N_621,In_1258,In_2487);
nand U622 (N_622,In_338,In_884);
and U623 (N_623,In_506,In_2241);
nand U624 (N_624,In_2252,In_2627);
nor U625 (N_625,In_1202,In_659);
nand U626 (N_626,In_716,In_110);
nand U627 (N_627,In_2985,In_1729);
nand U628 (N_628,In_14,In_1745);
nor U629 (N_629,In_643,In_339);
and U630 (N_630,In_2596,In_1476);
nand U631 (N_631,In_717,In_534);
nand U632 (N_632,In_920,In_2019);
xor U633 (N_633,In_1081,In_2828);
or U634 (N_634,In_2193,In_505);
nor U635 (N_635,In_37,In_1958);
and U636 (N_636,In_1772,In_1911);
xnor U637 (N_637,In_258,In_1858);
nand U638 (N_638,In_1675,In_2819);
and U639 (N_639,In_2280,In_228);
nor U640 (N_640,In_2186,In_430);
nand U641 (N_641,In_1941,In_1656);
nand U642 (N_642,In_172,In_2455);
nor U643 (N_643,In_234,In_2437);
nor U644 (N_644,In_663,In_1328);
nand U645 (N_645,In_458,In_1616);
or U646 (N_646,In_1200,In_1414);
or U647 (N_647,In_2649,In_2589);
and U648 (N_648,In_2833,In_169);
or U649 (N_649,In_1521,In_81);
nor U650 (N_650,In_706,In_1683);
or U651 (N_651,In_2378,In_2655);
or U652 (N_652,In_2161,In_1322);
nor U653 (N_653,In_972,In_418);
nand U654 (N_654,In_752,In_1751);
nand U655 (N_655,In_1219,In_2293);
xnor U656 (N_656,In_1966,In_791);
xor U657 (N_657,In_866,In_397);
xnor U658 (N_658,In_2226,In_382);
nor U659 (N_659,In_1084,In_1191);
and U660 (N_660,In_2992,In_447);
nand U661 (N_661,In_2433,In_1537);
nor U662 (N_662,In_2292,In_1390);
xor U663 (N_663,In_1035,In_1496);
or U664 (N_664,In_282,In_277);
nor U665 (N_665,In_2453,In_923);
nand U666 (N_666,In_280,In_1874);
xor U667 (N_667,In_1699,In_256);
xor U668 (N_668,In_2815,In_46);
nor U669 (N_669,In_1051,In_2396);
xnor U670 (N_670,In_2611,In_2299);
and U671 (N_671,In_99,In_1764);
nand U672 (N_672,In_373,In_1698);
nor U673 (N_673,In_1700,In_2251);
and U674 (N_674,In_1530,In_2654);
or U675 (N_675,In_355,In_1684);
xnor U676 (N_676,In_2425,In_2505);
nand U677 (N_677,In_2921,In_53);
xor U678 (N_678,In_337,In_237);
and U679 (N_679,In_2930,In_2351);
and U680 (N_680,In_939,In_335);
nand U681 (N_681,In_2044,In_1600);
xor U682 (N_682,In_639,In_698);
nor U683 (N_683,In_797,In_1990);
nor U684 (N_684,In_480,In_184);
and U685 (N_685,In_2638,In_854);
and U686 (N_686,In_10,In_976);
and U687 (N_687,In_1869,In_892);
nand U688 (N_688,In_941,In_2185);
and U689 (N_689,In_1485,In_1088);
xor U690 (N_690,In_1164,In_2673);
nand U691 (N_691,In_692,In_940);
nor U692 (N_692,In_2081,In_724);
xnor U693 (N_693,In_378,In_2345);
or U694 (N_694,In_2369,In_2697);
nor U695 (N_695,In_398,In_1526);
nand U696 (N_696,In_956,In_1494);
nor U697 (N_697,In_2794,In_1246);
nor U698 (N_698,In_91,In_1875);
or U699 (N_699,In_2246,In_2804);
or U700 (N_700,In_2792,In_151);
and U701 (N_701,In_1469,In_814);
or U702 (N_702,In_2318,In_2939);
nand U703 (N_703,In_2665,In_1228);
nor U704 (N_704,In_979,In_2153);
nand U705 (N_705,In_1901,In_2628);
xor U706 (N_706,In_12,In_121);
nor U707 (N_707,In_1949,In_1437);
nor U708 (N_708,In_1057,In_2149);
or U709 (N_709,In_191,In_1972);
nand U710 (N_710,In_2656,In_1417);
nor U711 (N_711,In_2467,In_575);
and U712 (N_712,In_259,In_2392);
or U713 (N_713,In_2983,In_2391);
and U714 (N_714,In_344,In_2289);
and U715 (N_715,In_560,In_2068);
nor U716 (N_716,In_605,In_226);
and U717 (N_717,In_370,In_543);
nor U718 (N_718,In_2257,In_1885);
or U719 (N_719,In_1651,In_2418);
nand U720 (N_720,In_2477,In_1519);
xor U721 (N_721,In_182,In_1719);
nand U722 (N_722,In_2399,In_55);
or U723 (N_723,In_419,In_2309);
nand U724 (N_724,In_2704,In_2581);
nor U725 (N_725,In_117,In_1308);
and U726 (N_726,In_1212,In_2341);
nand U727 (N_727,In_700,In_584);
nor U728 (N_728,In_1427,In_1845);
or U729 (N_729,In_2091,In_1083);
nand U730 (N_730,In_1536,In_2007);
and U731 (N_731,In_586,In_1324);
xnor U732 (N_732,In_1969,In_507);
and U733 (N_733,In_1733,In_1591);
nand U734 (N_734,In_2140,In_1352);
or U735 (N_735,In_2536,In_800);
xor U736 (N_736,In_330,In_2834);
or U737 (N_737,In_1787,In_1907);
nand U738 (N_738,In_726,In_2136);
xor U739 (N_739,In_730,In_394);
xnor U740 (N_740,In_594,In_1067);
and U741 (N_741,In_1818,In_414);
and U742 (N_742,In_996,In_796);
nor U743 (N_743,In_369,In_2599);
nand U744 (N_744,In_1252,In_454);
nand U745 (N_745,In_2166,In_761);
and U746 (N_746,In_2701,In_2387);
or U747 (N_747,In_2942,In_1069);
nand U748 (N_748,In_512,In_1805);
and U749 (N_749,In_2797,In_2604);
nand U750 (N_750,In_1491,In_1802);
and U751 (N_751,In_535,In_58);
or U752 (N_752,In_2961,In_1780);
and U753 (N_753,In_1255,In_1095);
or U754 (N_754,In_778,In_810);
nand U755 (N_755,In_2641,In_2107);
nand U756 (N_756,In_934,In_2215);
xor U757 (N_757,In_1314,In_276);
or U758 (N_758,In_34,In_1016);
or U759 (N_759,In_408,In_217);
xor U760 (N_760,In_2860,In_2077);
nor U761 (N_761,In_2502,In_229);
xnor U762 (N_762,In_1410,In_2445);
nand U763 (N_763,In_1398,In_2319);
nand U764 (N_764,In_2769,In_1227);
and U765 (N_765,In_1695,In_1777);
or U766 (N_766,In_1082,In_1769);
or U767 (N_767,In_2110,In_2157);
nand U768 (N_768,In_1594,In_2687);
xor U769 (N_769,In_2033,In_2138);
nand U770 (N_770,In_96,In_227);
or U771 (N_771,In_322,In_916);
nand U772 (N_772,In_2075,In_1369);
or U773 (N_773,In_1750,In_2622);
xor U774 (N_774,In_655,In_2428);
or U775 (N_775,In_1661,In_1906);
xnor U776 (N_776,In_2383,In_1166);
or U777 (N_777,In_597,In_2472);
xnor U778 (N_778,In_648,In_2721);
or U779 (N_779,In_751,In_79);
nand U780 (N_780,In_1801,In_666);
and U781 (N_781,In_2625,In_1910);
nor U782 (N_782,In_2739,In_1458);
xnor U783 (N_783,In_428,In_211);
xnor U784 (N_784,In_1705,In_2729);
or U785 (N_785,In_665,In_1983);
nand U786 (N_786,In_2389,In_1430);
xor U787 (N_787,In_2462,In_2582);
and U788 (N_788,In_409,In_696);
nor U789 (N_789,In_27,In_2620);
nand U790 (N_790,In_1636,In_166);
nand U791 (N_791,In_1634,In_367);
nand U792 (N_792,In_1244,In_2275);
nand U793 (N_793,In_279,In_1814);
or U794 (N_794,In_2000,In_435);
xnor U795 (N_795,In_2839,In_440);
and U796 (N_796,In_2988,In_1721);
nand U797 (N_797,In_1048,In_2571);
xnor U798 (N_798,In_544,In_2311);
nand U799 (N_799,In_2027,In_2030);
xor U800 (N_800,In_790,In_1407);
or U801 (N_801,In_2482,In_20);
and U802 (N_802,In_2817,In_359);
or U803 (N_803,In_2885,In_112);
xnor U804 (N_804,In_1217,In_2956);
or U805 (N_805,In_808,In_333);
or U806 (N_806,In_1694,In_2683);
nor U807 (N_807,In_1672,In_411);
or U808 (N_808,In_2950,In_1871);
xnor U809 (N_809,In_23,In_429);
nor U810 (N_810,In_1563,In_1732);
xor U811 (N_811,In_1278,In_1826);
nand U812 (N_812,In_2343,In_1336);
or U813 (N_813,In_1497,In_2272);
and U814 (N_814,In_1669,In_2853);
nand U815 (N_815,In_165,In_2537);
and U816 (N_816,In_887,In_2120);
nor U817 (N_817,In_763,In_1475);
nand U818 (N_818,In_1477,In_2175);
nor U819 (N_819,In_1794,In_2164);
xnor U820 (N_820,In_1555,In_141);
and U821 (N_821,In_1329,In_2411);
nor U822 (N_822,In_2749,In_2977);
nor U823 (N_823,In_1723,In_1986);
or U824 (N_824,In_600,In_2040);
xor U825 (N_825,In_1788,In_1667);
nand U826 (N_826,In_1350,In_2617);
and U827 (N_827,In_731,In_2256);
or U828 (N_828,In_1565,In_2514);
nor U829 (N_829,In_364,In_2181);
and U830 (N_830,In_2476,In_1819);
and U831 (N_831,In_1361,In_2856);
or U832 (N_832,In_2533,In_467);
or U833 (N_833,In_100,In_325);
nor U834 (N_834,In_747,In_2367);
nor U835 (N_835,In_2948,In_2740);
or U836 (N_836,In_1561,In_1859);
nor U837 (N_837,In_1605,In_1650);
nand U838 (N_838,In_2461,In_195);
xor U839 (N_839,In_400,In_2423);
or U840 (N_840,In_870,In_529);
nor U841 (N_841,In_1295,In_1138);
nor U842 (N_842,In_403,In_2667);
nand U843 (N_843,In_1313,In_2810);
nand U844 (N_844,In_2324,In_2436);
nand U845 (N_845,In_1277,In_1123);
nor U846 (N_846,In_795,In_366);
nor U847 (N_847,In_2422,In_1471);
or U848 (N_848,In_305,In_1060);
nor U849 (N_849,In_59,In_2184);
or U850 (N_850,In_1889,In_1294);
xor U851 (N_851,In_872,In_1223);
and U852 (N_852,In_1579,In_2067);
or U853 (N_853,In_2071,In_959);
and U854 (N_854,In_2541,In_1630);
or U855 (N_855,In_517,In_152);
xor U856 (N_856,In_1895,In_1965);
or U857 (N_857,In_2363,In_2830);
nor U858 (N_858,In_1737,In_2778);
nand U859 (N_859,In_1447,In_1064);
and U860 (N_860,In_877,In_2897);
nand U861 (N_861,In_1765,In_1954);
nor U862 (N_862,In_873,In_1531);
and U863 (N_863,In_2702,In_294);
xnor U864 (N_864,In_1042,In_1157);
and U865 (N_865,In_2158,In_2301);
xnor U866 (N_866,In_1748,In_342);
xor U867 (N_867,In_2583,In_235);
and U868 (N_868,In_1998,In_1677);
nand U869 (N_869,In_2208,In_287);
nand U870 (N_870,In_131,In_514);
nor U871 (N_871,In_630,In_2093);
nor U872 (N_872,In_1013,In_926);
or U873 (N_873,In_2211,In_817);
xor U874 (N_874,In_513,In_713);
and U875 (N_875,In_1860,In_1967);
and U876 (N_876,In_267,In_362);
or U877 (N_877,In_1929,In_1174);
or U878 (N_878,In_2259,In_2886);
nor U879 (N_879,In_1306,In_479);
or U880 (N_880,In_867,In_315);
nand U881 (N_881,In_318,In_1207);
nor U882 (N_882,In_2986,In_2056);
or U883 (N_883,In_784,In_2957);
and U884 (N_884,In_1229,In_1002);
nor U885 (N_885,In_744,In_386);
nor U886 (N_886,In_1383,In_1538);
nand U887 (N_887,In_1518,In_2699);
and U888 (N_888,In_2724,In_119);
nor U889 (N_889,In_1706,In_2538);
nand U890 (N_890,In_2680,In_1546);
xor U891 (N_891,In_571,In_2559);
and U892 (N_892,In_329,In_997);
nor U893 (N_893,In_2937,In_2731);
nand U894 (N_894,In_272,In_968);
nor U895 (N_895,In_2374,In_1731);
and U896 (N_896,In_2684,In_1734);
nand U897 (N_897,In_2053,In_687);
and U898 (N_898,In_2912,In_457);
or U899 (N_899,In_2284,In_1861);
and U900 (N_900,In_2910,In_1882);
xnor U901 (N_901,In_1442,In_2875);
xor U902 (N_902,In_2579,In_2195);
xnor U903 (N_903,In_2283,In_2469);
and U904 (N_904,In_2238,In_671);
or U905 (N_905,In_563,In_161);
nand U906 (N_906,In_1936,In_827);
xor U907 (N_907,In_2131,In_2767);
and U908 (N_908,In_2555,In_992);
and U909 (N_909,In_2421,In_1256);
or U910 (N_910,In_2970,In_860);
and U911 (N_911,In_1236,In_2295);
xnor U912 (N_912,In_2,In_1793);
and U913 (N_913,In_174,In_424);
and U914 (N_914,In_2282,In_545);
and U915 (N_915,In_2214,In_65);
or U916 (N_916,In_2312,In_2151);
and U917 (N_917,In_1092,In_841);
and U918 (N_918,In_1340,In_540);
nand U919 (N_919,In_1188,In_2493);
or U920 (N_920,In_2720,In_1209);
xnor U921 (N_921,In_243,In_2495);
or U922 (N_922,In_1261,In_374);
or U923 (N_923,In_539,In_609);
xor U924 (N_924,In_1806,In_162);
nand U925 (N_925,In_1931,In_2156);
or U926 (N_926,In_774,In_1039);
nor U927 (N_927,In_2250,In_2566);
and U928 (N_928,In_2303,In_1118);
nor U929 (N_929,In_2788,In_792);
nand U930 (N_930,In_1402,In_1330);
nor U931 (N_931,In_632,In_2811);
or U932 (N_932,In_170,In_772);
nor U933 (N_933,In_1556,In_2557);
nor U934 (N_934,In_562,In_2333);
nor U935 (N_935,In_715,In_1467);
nand U936 (N_936,In_2947,In_2703);
nor U937 (N_937,In_1576,In_1341);
nor U938 (N_938,In_1625,In_2973);
or U939 (N_939,In_1696,In_1429);
and U940 (N_940,In_114,In_1816);
xnor U941 (N_941,In_163,In_449);
xnor U942 (N_942,In_1971,In_1120);
nand U943 (N_943,In_1299,In_2232);
xor U944 (N_944,In_422,In_2700);
and U945 (N_945,In_559,In_2101);
nor U946 (N_946,In_1834,In_2227);
xor U947 (N_947,In_2521,In_741);
and U948 (N_948,In_2782,In_1100);
or U949 (N_949,In_2086,In_2737);
nor U950 (N_950,In_2170,In_423);
nor U951 (N_951,In_1866,In_1264);
xor U952 (N_952,In_568,In_2799);
xor U953 (N_953,In_2723,In_776);
nor U954 (N_954,In_1114,In_1332);
xnor U955 (N_955,In_781,In_764);
or U956 (N_956,In_482,In_2826);
xor U957 (N_957,In_2356,In_1233);
and U958 (N_958,In_2866,In_1077);
nor U959 (N_959,In_2212,In_459);
and U960 (N_960,In_354,In_1173);
nand U961 (N_961,In_530,In_2419);
nor U962 (N_962,In_556,In_1385);
and U963 (N_963,In_684,In_1702);
xor U964 (N_964,In_2167,In_2112);
nor U965 (N_965,In_1152,In_2544);
nor U966 (N_966,In_2753,In_1054);
or U967 (N_967,In_1670,In_2648);
or U968 (N_968,In_944,In_2751);
xnor U969 (N_969,In_1618,In_1473);
xor U970 (N_970,In_223,In_1596);
and U971 (N_971,In_1736,In_2530);
nand U972 (N_972,In_908,In_1950);
nor U973 (N_973,In_2443,In_1927);
xor U974 (N_974,In_2317,In_2406);
or U975 (N_975,In_861,In_2366);
nor U976 (N_976,In_2867,In_531);
and U977 (N_977,In_456,In_203);
nor U978 (N_978,In_42,In_1071);
and U979 (N_979,In_390,In_1553);
nor U980 (N_980,In_1302,In_1726);
nor U981 (N_981,In_2591,In_2357);
or U982 (N_982,In_197,In_1090);
nand U983 (N_983,In_193,In_903);
or U984 (N_984,In_1687,In_492);
and U985 (N_985,In_1041,In_2335);
xnor U986 (N_986,In_406,In_1919);
and U987 (N_987,In_75,In_569);
nor U988 (N_988,In_381,In_1147);
or U989 (N_989,In_1614,In_2384);
nand U990 (N_990,In_673,In_2235);
and U991 (N_991,In_2403,In_1795);
or U992 (N_992,In_1865,In_360);
nand U993 (N_993,In_1544,In_574);
nor U994 (N_994,In_1652,In_470);
nor U995 (N_995,In_1309,In_1438);
or U996 (N_996,In_907,In_2923);
xnor U997 (N_997,In_2084,In_765);
nand U998 (N_998,In_721,In_118);
xnor U999 (N_999,In_1668,In_1970);
nor U1000 (N_1000,In_647,In_1577);
or U1001 (N_1001,In_192,In_2306);
nand U1002 (N_1002,In_896,In_22);
and U1003 (N_1003,In_677,In_1624);
xor U1004 (N_1004,In_1439,In_1529);
nor U1005 (N_1005,In_76,In_2162);
nand U1006 (N_1006,In_323,In_1853);
nor U1007 (N_1007,In_1177,In_2180);
nor U1008 (N_1008,In_1824,In_879);
or U1009 (N_1009,In_2083,In_1899);
or U1010 (N_1010,In_1279,In_2109);
nand U1011 (N_1011,In_1010,In_317);
and U1012 (N_1012,In_262,In_2373);
xnor U1013 (N_1013,In_2882,In_160);
xnor U1014 (N_1014,In_439,In_2602);
or U1015 (N_1015,In_1019,In_889);
xor U1016 (N_1016,In_928,In_4);
nor U1017 (N_1017,In_637,In_1811);
nor U1018 (N_1018,In_650,In_1339);
nor U1019 (N_1019,In_2871,In_2849);
nand U1020 (N_1020,In_2837,In_1810);
or U1021 (N_1021,In_587,In_212);
or U1022 (N_1022,In_891,In_2730);
nor U1023 (N_1023,In_1366,In_2348);
nand U1024 (N_1024,In_421,In_1997);
nor U1025 (N_1025,In_1716,In_358);
nor U1026 (N_1026,In_1106,In_809);
and U1027 (N_1027,In_880,In_2524);
nor U1028 (N_1028,In_2350,In_293);
nand U1029 (N_1029,In_554,In_238);
and U1030 (N_1030,In_463,In_1030);
nor U1031 (N_1031,In_2230,In_2388);
or U1032 (N_1032,In_2861,In_2869);
xor U1033 (N_1033,In_1922,In_943);
xnor U1034 (N_1034,In_35,In_284);
and U1035 (N_1035,In_2096,In_2686);
nor U1036 (N_1036,In_2127,In_1403);
xnor U1037 (N_1037,In_1608,In_679);
nor U1038 (N_1038,In_1384,In_1948);
xor U1039 (N_1039,In_297,In_1593);
and U1040 (N_1040,In_1498,In_1344);
or U1041 (N_1041,In_1412,In_2758);
nand U1042 (N_1042,In_126,In_2675);
and U1043 (N_1043,In_579,In_2085);
nor U1044 (N_1044,In_511,In_2058);
and U1045 (N_1045,In_2796,In_825);
or U1046 (N_1046,In_1604,In_2634);
and U1047 (N_1047,In_1523,In_1517);
xnor U1048 (N_1048,In_72,In_292);
xnor U1049 (N_1049,In_1746,In_1783);
and U1050 (N_1050,In_1043,In_750);
and U1051 (N_1051,In_2409,In_983);
nand U1052 (N_1052,In_2960,In_2520);
nor U1053 (N_1053,In_2245,In_2601);
nand U1054 (N_1054,In_1175,In_1779);
xnor U1055 (N_1055,In_1337,In_593);
or U1056 (N_1056,In_2407,In_749);
xnor U1057 (N_1057,In_1047,In_402);
nand U1058 (N_1058,In_156,In_1466);
and U1059 (N_1059,In_1580,In_589);
or U1060 (N_1060,In_882,In_1976);
nor U1061 (N_1061,In_431,In_1773);
or U1062 (N_1062,In_1285,In_793);
nor U1063 (N_1063,In_1377,In_1179);
and U1064 (N_1064,In_2879,In_2574);
and U1065 (N_1065,In_266,In_1396);
and U1066 (N_1066,In_930,In_60);
and U1067 (N_1067,In_1528,In_1374);
and U1068 (N_1068,In_2500,In_888);
xnor U1069 (N_1069,In_2048,In_550);
or U1070 (N_1070,In_1864,In_1583);
and U1071 (N_1071,In_2927,In_1981);
xnor U1072 (N_1072,In_271,In_40);
and U1073 (N_1073,In_520,In_1738);
xor U1074 (N_1074,In_2657,In_2054);
nand U1075 (N_1075,In_2941,In_1942);
nand U1076 (N_1076,In_108,In_1720);
nand U1077 (N_1077,In_1840,In_2873);
nor U1078 (N_1078,In_2848,In_1418);
xor U1079 (N_1079,In_1091,In_2727);
xor U1080 (N_1080,In_2297,In_274);
nand U1081 (N_1081,In_1284,In_2529);
nand U1082 (N_1082,In_2485,In_767);
xnor U1083 (N_1083,In_2076,In_1281);
nand U1084 (N_1084,In_2014,In_1001);
nor U1085 (N_1085,In_1562,In_462);
nand U1086 (N_1086,In_1449,In_2790);
and U1087 (N_1087,In_57,In_1612);
nand U1088 (N_1088,In_1161,In_2705);
or U1089 (N_1089,In_1248,In_1142);
nor U1090 (N_1090,In_1715,In_301);
nor U1091 (N_1091,In_2658,In_2330);
and U1092 (N_1092,In_251,In_1190);
nor U1093 (N_1093,In_1909,In_995);
nor U1094 (N_1094,In_1406,In_1797);
nand U1095 (N_1095,In_735,In_802);
and U1096 (N_1096,In_1785,In_2709);
xor U1097 (N_1097,In_2024,In_1928);
xnor U1098 (N_1098,In_450,In_1803);
or U1099 (N_1099,In_1122,In_2016);
xor U1100 (N_1100,In_64,In_2635);
xor U1101 (N_1101,In_1194,In_1089);
and U1102 (N_1102,In_2382,In_652);
nor U1103 (N_1103,In_753,In_829);
and U1104 (N_1104,In_186,In_1982);
nor U1105 (N_1105,In_2320,In_2229);
xor U1106 (N_1106,In_2618,In_1710);
or U1107 (N_1107,In_353,In_1136);
xor U1108 (N_1108,In_2691,In_207);
or U1109 (N_1109,In_801,In_2598);
and U1110 (N_1110,In_1451,In_273);
and U1111 (N_1111,In_2595,In_2917);
or U1112 (N_1112,In_2481,In_823);
nand U1113 (N_1113,In_2291,In_1022);
or U1114 (N_1114,In_984,In_1760);
nand U1115 (N_1115,In_2304,In_2045);
xor U1116 (N_1116,In_718,In_656);
nand U1117 (N_1117,In_2360,In_461);
and U1118 (N_1118,In_886,In_66);
and U1119 (N_1119,In_1956,In_2255);
xor U1120 (N_1120,In_631,In_1549);
and U1121 (N_1121,In_2349,In_2347);
nor U1122 (N_1122,In_1660,In_788);
nor U1123 (N_1123,In_894,In_838);
or U1124 (N_1124,In_1742,In_2526);
nand U1125 (N_1125,In_599,In_1072);
nor U1126 (N_1126,In_1766,In_519);
and U1127 (N_1127,In_41,In_384);
and U1128 (N_1128,In_2145,In_2194);
xnor U1129 (N_1129,In_2057,In_2570);
or U1130 (N_1130,In_67,In_2644);
or U1131 (N_1131,In_416,In_133);
or U1132 (N_1132,In_1196,In_2586);
nor U1133 (N_1133,In_1415,In_2857);
and U1134 (N_1134,In_851,In_2457);
nor U1135 (N_1135,In_1274,In_2845);
nor U1136 (N_1136,In_1134,In_932);
xor U1137 (N_1137,In_1601,In_2070);
nor U1138 (N_1138,In_993,In_1367);
nand U1139 (N_1139,In_601,In_2732);
xor U1140 (N_1140,In_2786,In_189);
or U1141 (N_1141,In_1884,In_1622);
or U1142 (N_1142,In_2809,In_2631);
and U1143 (N_1143,In_312,In_2450);
and U1144 (N_1144,In_345,In_1040);
and U1145 (N_1145,In_518,In_1620);
nor U1146 (N_1146,In_768,In_2325);
nor U1147 (N_1147,In_1527,In_757);
or U1148 (N_1148,In_2087,In_2294);
and U1149 (N_1149,In_1891,In_147);
and U1150 (N_1150,In_924,In_1393);
nand U1151 (N_1151,In_1762,In_1847);
nand U1152 (N_1152,In_755,In_570);
and U1153 (N_1153,In_2460,In_1003);
nor U1154 (N_1154,In_2590,In_557);
and U1155 (N_1155,In_289,In_2966);
nor U1156 (N_1156,In_2606,In_2868);
nand U1157 (N_1157,In_2210,In_2822);
and U1158 (N_1158,In_1628,In_807);
or U1159 (N_1159,In_542,In_1457);
and U1160 (N_1160,In_1452,In_1267);
xor U1161 (N_1161,In_524,In_1443);
xor U1162 (N_1162,In_948,In_640);
or U1163 (N_1163,In_1181,In_1989);
and U1164 (N_1164,In_2381,In_2290);
xor U1165 (N_1165,In_298,In_1490);
nor U1166 (N_1166,In_1250,In_283);
xor U1167 (N_1167,In_1025,In_2191);
and U1168 (N_1168,In_2506,In_822);
and U1169 (N_1169,In_745,In_1303);
nand U1170 (N_1170,In_2190,In_2305);
nor U1171 (N_1171,In_2938,In_1607);
and U1172 (N_1172,In_106,In_496);
and U1173 (N_1173,In_1479,In_691);
xnor U1174 (N_1174,In_1588,In_1754);
nor U1175 (N_1175,In_2677,In_1058);
nand U1176 (N_1176,In_2688,In_2551);
nor U1177 (N_1177,In_694,In_591);
or U1178 (N_1178,In_253,In_1728);
nand U1179 (N_1179,In_2189,In_1775);
or U1180 (N_1180,In_1552,In_2221);
and U1181 (N_1181,In_759,In_2233);
or U1182 (N_1182,In_670,In_304);
nand U1183 (N_1183,In_2465,In_2800);
or U1184 (N_1184,In_2695,In_2858);
and U1185 (N_1185,In_1569,In_336);
and U1186 (N_1186,In_2510,In_1222);
nand U1187 (N_1187,In_2755,In_2547);
nand U1188 (N_1188,In_2321,In_2621);
nand U1189 (N_1189,In_246,In_2339);
and U1190 (N_1190,In_2432,In_2147);
nor U1191 (N_1191,In_1541,In_2678);
nor U1192 (N_1192,In_2059,In_1426);
nand U1193 (N_1193,In_485,In_136);
nand U1194 (N_1194,In_607,In_1932);
or U1195 (N_1195,In_1386,In_537);
nand U1196 (N_1196,In_2978,In_1162);
nor U1197 (N_1197,In_38,In_1503);
nand U1198 (N_1198,In_1681,In_498);
xor U1199 (N_1199,In_1992,In_349);
or U1200 (N_1200,In_1893,In_311);
nor U1201 (N_1201,In_547,In_1566);
xnor U1202 (N_1202,In_1655,In_590);
nand U1203 (N_1203,In_1011,In_1465);
nand U1204 (N_1204,In_2562,In_268);
xnor U1205 (N_1205,In_1419,In_216);
and U1206 (N_1206,In_2119,In_1567);
nor U1207 (N_1207,In_662,In_1781);
nor U1208 (N_1208,In_2615,In_1520);
nand U1209 (N_1209,In_2261,In_1078);
and U1210 (N_1210,In_2468,In_1251);
or U1211 (N_1211,In_1436,In_2183);
xnor U1212 (N_1212,In_2842,In_1300);
xor U1213 (N_1213,In_541,In_2046);
nand U1214 (N_1214,In_2498,In_2179);
and U1215 (N_1215,In_2199,In_952);
nor U1216 (N_1216,In_917,In_1493);
or U1217 (N_1217,In_2281,In_499);
and U1218 (N_1218,In_1848,In_2354);
and U1219 (N_1219,In_2213,In_2863);
nand U1220 (N_1220,In_143,In_2824);
xnor U1221 (N_1221,In_1061,In_1036);
and U1222 (N_1222,In_1132,In_1571);
xor U1223 (N_1223,In_1210,In_48);
nor U1224 (N_1224,In_2693,In_2525);
nor U1225 (N_1225,In_711,In_813);
and U1226 (N_1226,In_844,In_1144);
or U1227 (N_1227,In_1602,In_302);
nand U1228 (N_1228,In_927,In_1052);
and U1229 (N_1229,In_1318,In_2999);
and U1230 (N_1230,In_2793,In_2263);
or U1231 (N_1231,In_727,In_1872);
nor U1232 (N_1232,In_2448,In_1086);
nand U1233 (N_1233,In_2104,In_2427);
and U1234 (N_1234,In_2017,In_2512);
and U1235 (N_1235,In_2006,In_2049);
nand U1236 (N_1236,In_2877,In_2636);
and U1237 (N_1237,In_220,In_732);
xnor U1238 (N_1238,In_1,In_1319);
or U1239 (N_1239,In_1581,In_646);
xnor U1240 (N_1240,In_805,In_1023);
nor U1241 (N_1241,In_1029,In_1844);
xor U1242 (N_1242,In_2248,In_2708);
xnor U1243 (N_1243,In_1124,In_2177);
xor U1244 (N_1244,In_2088,In_2694);
and U1245 (N_1245,In_2353,In_379);
or U1246 (N_1246,In_1633,In_1215);
or U1247 (N_1247,In_914,In_2173);
and U1248 (N_1248,In_785,In_728);
and U1249 (N_1249,In_681,In_105);
or U1250 (N_1250,In_2663,In_2026);
nor U1251 (N_1251,In_1468,In_1180);
or U1252 (N_1252,In_1074,In_401);
nand U1253 (N_1253,In_1817,In_1917);
xor U1254 (N_1254,In_2089,In_49);
xnor U1255 (N_1255,In_2614,In_2475);
xnor U1256 (N_1256,In_257,In_371);
or U1257 (N_1257,In_1007,In_2197);
xnor U1258 (N_1258,In_2765,In_642);
xnor U1259 (N_1259,In_1127,In_477);
or U1260 (N_1260,In_2556,In_1004);
nor U1261 (N_1261,In_2925,In_1364);
nor U1262 (N_1262,In_960,In_1739);
xnor U1263 (N_1263,In_1961,In_473);
or U1264 (N_1264,In_2588,In_2922);
nor U1265 (N_1265,In_614,In_1014);
xor U1266 (N_1266,In_2400,In_494);
or U1267 (N_1267,In_875,In_1610);
or U1268 (N_1268,In_733,In_786);
or U1269 (N_1269,In_1642,In_395);
and U1270 (N_1270,In_446,In_63);
and U1271 (N_1271,In_2940,In_1682);
nand U1272 (N_1272,In_2870,In_17);
nand U1273 (N_1273,In_368,In_1846);
xnor U1274 (N_1274,In_1830,In_50);
nor U1275 (N_1275,In_1946,In_29);
nor U1276 (N_1276,In_565,In_2681);
xor U1277 (N_1277,In_1347,In_1168);
and U1278 (N_1278,In_1359,In_2728);
or U1279 (N_1279,In_491,In_1110);
xnor U1280 (N_1280,In_232,In_1141);
xor U1281 (N_1281,In_1448,In_2015);
and U1282 (N_1282,In_1615,In_2496);
nor U1283 (N_1283,In_615,In_2517);
xnor U1284 (N_1284,In_840,In_188);
nor U1285 (N_1285,In_443,In_1075);
or U1286 (N_1286,In_387,In_1926);
nand U1287 (N_1287,In_2129,In_1484);
and U1288 (N_1288,In_1685,In_230);
nor U1289 (N_1289,In_532,In_1545);
and U1290 (N_1290,In_1560,In_157);
or U1291 (N_1291,In_2674,In_1104);
nor U1292 (N_1292,In_2121,In_144);
nor U1293 (N_1293,In_1317,In_2228);
nand U1294 (N_1294,In_2777,In_815);
nor U1295 (N_1295,In_1440,In_437);
xnor U1296 (N_1296,In_1890,In_1113);
or U1297 (N_1297,In_31,In_2441);
nand U1298 (N_1298,In_1833,In_314);
xor U1299 (N_1299,In_2578,In_2483);
nor U1300 (N_1300,In_1880,In_352);
xnor U1301 (N_1301,In_1613,In_2452);
nor U1302 (N_1302,In_250,In_2328);
nand U1303 (N_1303,In_2078,In_2575);
xor U1304 (N_1304,In_2733,In_348);
nand U1305 (N_1305,In_2971,In_1851);
nand U1306 (N_1306,In_62,In_39);
xor U1307 (N_1307,In_1878,In_1487);
or U1308 (N_1308,In_967,In_122);
xnor U1309 (N_1309,In_2316,In_61);
and U1310 (N_1310,In_2773,In_343);
or U1311 (N_1311,In_288,In_848);
nand U1312 (N_1312,In_281,In_2021);
nand U1313 (N_1313,In_2106,In_2626);
nand U1314 (N_1314,In_138,In_2466);
and U1315 (N_1315,In_929,In_862);
nand U1316 (N_1316,In_1371,In_306);
nor U1317 (N_1317,In_1782,In_1582);
and U1318 (N_1318,In_2847,In_2010);
xnor U1319 (N_1319,In_2679,In_1349);
and U1320 (N_1320,In_13,In_1662);
or U1321 (N_1321,In_1293,In_451);
nand U1322 (N_1322,In_194,In_2616);
xnor U1323 (N_1323,In_504,In_2812);
or U1324 (N_1324,In_629,In_690);
xnor U1325 (N_1325,In_1843,In_1626);
xor U1326 (N_1326,In_1182,In_2630);
and U1327 (N_1327,In_1342,In_2805);
and U1328 (N_1328,In_2798,In_1962);
and U1329 (N_1329,In_2823,In_2486);
xnor U1330 (N_1330,In_1841,In_1592);
or U1331 (N_1331,In_285,In_2889);
or U1332 (N_1332,In_2707,In_1504);
xnor U1333 (N_1333,In_816,In_566);
and U1334 (N_1334,In_1730,In_833);
or U1335 (N_1335,In_674,In_321);
xnor U1336 (N_1336,In_2587,In_915);
or U1337 (N_1337,In_1873,In_729);
and U1338 (N_1338,In_621,In_661);
xnor U1339 (N_1339,In_1532,In_2034);
nand U1340 (N_1340,In_1165,In_2176);
or U1341 (N_1341,In_966,In_1935);
xor U1342 (N_1342,In_1689,In_1360);
nor U1343 (N_1343,In_1912,In_1606);
or U1344 (N_1344,In_239,In_2646);
nor U1345 (N_1345,In_1623,In_1323);
and U1346 (N_1346,In_93,In_2390);
xor U1347 (N_1347,In_2840,In_2009);
or U1348 (N_1348,In_1513,In_1963);
nor U1349 (N_1349,In_205,In_1585);
xor U1350 (N_1350,In_171,In_1198);
nand U1351 (N_1351,In_1068,In_2545);
nand U1352 (N_1352,In_73,In_260);
or U1353 (N_1353,In_2377,In_2735);
and U1354 (N_1354,In_2945,In_1370);
nor U1355 (N_1355,In_2906,In_852);
nor U1356 (N_1356,In_2803,In_970);
xnor U1357 (N_1357,In_1724,In_1547);
nand U1358 (N_1358,In_26,In_2968);
nor U1359 (N_1359,In_2346,In_1259);
xnor U1360 (N_1360,In_1554,In_2090);
or U1361 (N_1361,In_2752,In_1201);
or U1362 (N_1362,In_902,In_1644);
nand U1363 (N_1363,In_1815,In_1876);
nor U1364 (N_1364,In_1093,In_433);
nor U1365 (N_1365,In_1849,In_625);
or U1366 (N_1366,In_175,In_1130);
nor U1367 (N_1367,In_977,In_1460);
nand U1368 (N_1368,In_2308,In_1131);
nor U1369 (N_1369,In_320,In_868);
xor U1370 (N_1370,In_222,In_1854);
nor U1371 (N_1371,In_1789,In_2850);
and U1372 (N_1372,In_2413,In_2608);
or U1373 (N_1373,In_1150,In_1214);
or U1374 (N_1374,In_2372,In_2155);
nor U1375 (N_1375,In_2332,In_2492);
xor U1376 (N_1376,In_1391,In_1462);
nor U1377 (N_1377,In_2036,In_363);
nand U1378 (N_1378,In_913,In_1486);
nor U1379 (N_1379,In_2672,In_2668);
nand U1380 (N_1380,In_1933,In_2531);
nor U1381 (N_1381,In_846,In_481);
nor U1382 (N_1382,In_2946,In_1499);
xnor U1383 (N_1383,In_2198,In_2322);
xnor U1384 (N_1384,In_1225,In_372);
or U1385 (N_1385,In_2883,In_1892);
or U1386 (N_1386,In_1646,In_2326);
xor U1387 (N_1387,In_1357,In_1031);
xor U1388 (N_1388,In_723,In_1937);
nand U1389 (N_1389,In_2489,In_1269);
nand U1390 (N_1390,In_167,In_2035);
and U1391 (N_1391,In_620,In_1454);
xor U1392 (N_1392,In_664,In_2951);
and U1393 (N_1393,In_1115,In_1153);
or U1394 (N_1394,In_975,In_442);
and U1395 (N_1395,In_2125,In_1482);
nand U1396 (N_1396,In_2062,In_89);
and U1397 (N_1397,In_2237,In_426);
and U1398 (N_1398,In_2276,In_495);
and U1399 (N_1399,In_351,In_2394);
xor U1400 (N_1400,In_1126,In_712);
and U1401 (N_1401,In_441,In_641);
xor U1402 (N_1402,In_2717,In_2789);
xor U1403 (N_1403,In_107,In_483);
nor U1404 (N_1404,In_104,In_516);
and U1405 (N_1405,In_1973,In_1353);
xnor U1406 (N_1406,In_859,In_2509);
nor U1407 (N_1407,In_1747,In_2991);
nand U1408 (N_1408,In_624,In_2855);
or U1409 (N_1409,In_2124,In_821);
and U1410 (N_1410,In_1903,In_2287);
and U1411 (N_1411,In_921,In_905);
nand U1412 (N_1412,In_853,In_874);
or U1413 (N_1413,In_87,In_1524);
nand U1414 (N_1414,In_1807,In_2488);
nor U1415 (N_1415,In_2808,In_420);
and U1416 (N_1416,In_1778,In_1790);
xor U1417 (N_1417,In_2338,In_51);
or U1418 (N_1418,In_1265,In_2519);
or U1419 (N_1419,In_2115,In_2775);
or U1420 (N_1420,In_904,In_1170);
or U1421 (N_1421,In_2025,In_327);
xnor U1422 (N_1422,In_1825,In_1828);
nand U1423 (N_1423,In_2905,In_695);
and U1424 (N_1424,In_2516,In_871);
xor U1425 (N_1425,In_2943,In_221);
and U1426 (N_1426,In_2768,In_1167);
nand U1427 (N_1427,In_771,In_319);
nand U1428 (N_1428,In_2202,In_2262);
xnor U1429 (N_1429,In_497,In_2746);
and U1430 (N_1430,In_1943,In_1896);
nand U1431 (N_1431,In_1012,In_2607);
nor U1432 (N_1432,In_80,In_334);
nand U1433 (N_1433,In_120,In_2417);
and U1434 (N_1434,In_596,In_1887);
nor U1435 (N_1435,In_527,In_1862);
or U1436 (N_1436,In_1389,In_97);
or U1437 (N_1437,In_1978,In_1586);
and U1438 (N_1438,In_2734,In_1542);
xor U1439 (N_1439,In_412,In_425);
nor U1440 (N_1440,In_773,In_1028);
xor U1441 (N_1441,In_1027,In_893);
nand U1442 (N_1442,In_2843,In_1243);
nor U1443 (N_1443,In_1087,In_1338);
or U1444 (N_1444,In_1914,In_1411);
and U1445 (N_1445,In_1835,In_2404);
or U1446 (N_1446,In_1049,In_316);
nor U1447 (N_1447,In_818,In_1038);
or U1448 (N_1448,In_264,In_672);
or U1449 (N_1449,In_1129,In_865);
xor U1450 (N_1450,In_1099,In_326);
nor U1451 (N_1451,In_2234,In_2759);
and U1452 (N_1452,In_606,In_1749);
or U1453 (N_1453,In_2254,In_2442);
nor U1454 (N_1454,In_2342,In_2079);
or U1455 (N_1455,In_2169,In_1756);
xor U1456 (N_1456,In_2066,In_2914);
nor U1457 (N_1457,In_1548,In_2041);
nor U1458 (N_1458,In_486,In_2122);
nor U1459 (N_1459,In_1156,In_153);
nand U1460 (N_1460,In_2762,In_2362);
or U1461 (N_1461,In_1304,In_1237);
nor U1462 (N_1462,In_328,In_699);
and U1463 (N_1463,In_2327,In_1888);
xor U1464 (N_1464,In_2100,In_1160);
nand U1465 (N_1465,In_990,In_261);
and U1466 (N_1466,In_619,In_1693);
or U1467 (N_1467,In_982,In_2664);
nor U1468 (N_1468,In_1743,In_2928);
nor U1469 (N_1469,In_2094,In_2761);
nor U1470 (N_1470,In_2008,In_269);
or U1471 (N_1471,In_573,In_115);
nand U1472 (N_1472,In_190,In_1205);
or U1473 (N_1473,In_1381,In_1711);
or U1474 (N_1474,In_1094,In_958);
and U1475 (N_1475,In_911,In_935);
xnor U1476 (N_1476,In_826,In_2738);
and U1477 (N_1477,In_1938,In_1761);
and U1478 (N_1478,In_978,In_843);
nand U1479 (N_1479,In_1578,In_2268);
and U1480 (N_1480,In_2368,In_1836);
and U1481 (N_1481,In_1944,In_1654);
or U1482 (N_1482,In_1413,In_1868);
or U1483 (N_1483,In_2887,In_1211);
xnor U1484 (N_1484,In_444,In_1169);
and U1485 (N_1485,In_2878,In_1472);
and U1486 (N_1486,In_1658,In_1597);
nor U1487 (N_1487,In_2061,In_1172);
xnor U1488 (N_1488,In_1163,In_2002);
or U1489 (N_1489,In_1502,In_1408);
and U1490 (N_1490,In_837,In_2558);
or U1491 (N_1491,In_2832,In_1098);
nor U1492 (N_1492,In_2924,In_2597);
or U1493 (N_1493,In_743,In_1345);
xor U1494 (N_1494,In_1573,In_1298);
nor U1495 (N_1495,In_2097,In_2479);
and U1496 (N_1496,In_432,In_680);
or U1497 (N_1497,In_1301,In_1105);
or U1498 (N_1498,In_618,In_1286);
nand U1499 (N_1499,In_453,In_561);
or U1500 (N_1500,N_563,N_771);
xnor U1501 (N_1501,N_635,N_311);
xnor U1502 (N_1502,N_268,N_482);
nor U1503 (N_1503,N_853,N_1382);
nand U1504 (N_1504,N_911,N_824);
or U1505 (N_1505,N_219,N_779);
nand U1506 (N_1506,N_1108,N_1230);
nor U1507 (N_1507,N_1426,N_703);
and U1508 (N_1508,N_1104,N_1076);
nand U1509 (N_1509,N_294,N_105);
nand U1510 (N_1510,N_712,N_378);
and U1511 (N_1511,N_478,N_425);
xor U1512 (N_1512,N_422,N_592);
or U1513 (N_1513,N_851,N_1282);
xnor U1514 (N_1514,N_1127,N_816);
or U1515 (N_1515,N_1254,N_708);
nor U1516 (N_1516,N_84,N_1143);
or U1517 (N_1517,N_224,N_947);
xor U1518 (N_1518,N_182,N_313);
or U1519 (N_1519,N_533,N_309);
or U1520 (N_1520,N_1090,N_556);
or U1521 (N_1521,N_354,N_8);
nand U1522 (N_1522,N_432,N_992);
and U1523 (N_1523,N_1101,N_450);
and U1524 (N_1524,N_1201,N_1133);
xnor U1525 (N_1525,N_693,N_167);
xor U1526 (N_1526,N_794,N_350);
xor U1527 (N_1527,N_106,N_162);
and U1528 (N_1528,N_1126,N_178);
and U1529 (N_1529,N_1189,N_652);
nand U1530 (N_1530,N_1263,N_1171);
xor U1531 (N_1531,N_1204,N_869);
or U1532 (N_1532,N_142,N_765);
nand U1533 (N_1533,N_1086,N_341);
and U1534 (N_1534,N_459,N_1052);
and U1535 (N_1535,N_618,N_164);
xnor U1536 (N_1536,N_32,N_250);
nand U1537 (N_1537,N_1423,N_53);
nor U1538 (N_1538,N_1373,N_898);
xor U1539 (N_1539,N_988,N_930);
or U1540 (N_1540,N_395,N_266);
nor U1541 (N_1541,N_1049,N_935);
nand U1542 (N_1542,N_99,N_418);
xnor U1543 (N_1543,N_277,N_1179);
xnor U1544 (N_1544,N_915,N_226);
xor U1545 (N_1545,N_590,N_86);
nand U1546 (N_1546,N_784,N_1285);
xnor U1547 (N_1547,N_1366,N_774);
xor U1548 (N_1548,N_507,N_1464);
nor U1549 (N_1549,N_289,N_767);
xnor U1550 (N_1550,N_279,N_995);
nor U1551 (N_1551,N_545,N_1103);
or U1552 (N_1552,N_104,N_887);
xor U1553 (N_1553,N_1338,N_516);
or U1554 (N_1554,N_241,N_431);
and U1555 (N_1555,N_1190,N_428);
nand U1556 (N_1556,N_134,N_754);
or U1557 (N_1557,N_1438,N_837);
xor U1558 (N_1558,N_486,N_814);
or U1559 (N_1559,N_1094,N_338);
nor U1560 (N_1560,N_717,N_768);
and U1561 (N_1561,N_377,N_1007);
xor U1562 (N_1562,N_473,N_1405);
and U1563 (N_1563,N_144,N_1330);
or U1564 (N_1564,N_382,N_396);
or U1565 (N_1565,N_681,N_657);
and U1566 (N_1566,N_1158,N_136);
and U1567 (N_1567,N_113,N_198);
and U1568 (N_1568,N_1173,N_1401);
nand U1569 (N_1569,N_251,N_588);
and U1570 (N_1570,N_695,N_349);
xor U1571 (N_1571,N_1192,N_892);
nor U1572 (N_1572,N_1390,N_1412);
or U1573 (N_1573,N_153,N_72);
xor U1574 (N_1574,N_936,N_252);
or U1575 (N_1575,N_1031,N_940);
or U1576 (N_1576,N_320,N_442);
and U1577 (N_1577,N_623,N_287);
or U1578 (N_1578,N_1281,N_549);
nor U1579 (N_1579,N_580,N_411);
or U1580 (N_1580,N_616,N_207);
nor U1581 (N_1581,N_729,N_161);
nor U1582 (N_1582,N_743,N_1396);
nor U1583 (N_1583,N_1333,N_1169);
nor U1584 (N_1584,N_686,N_671);
and U1585 (N_1585,N_1456,N_581);
or U1586 (N_1586,N_830,N_68);
and U1587 (N_1587,N_1339,N_974);
nor U1588 (N_1588,N_211,N_228);
nand U1589 (N_1589,N_965,N_1299);
xor U1590 (N_1590,N_557,N_1258);
nand U1591 (N_1591,N_854,N_48);
and U1592 (N_1592,N_66,N_43);
nand U1593 (N_1593,N_352,N_468);
nand U1594 (N_1594,N_1453,N_394);
xor U1595 (N_1595,N_353,N_1208);
nand U1596 (N_1596,N_271,N_532);
or U1597 (N_1597,N_535,N_534);
or U1598 (N_1598,N_945,N_101);
xor U1599 (N_1599,N_400,N_704);
xnor U1600 (N_1600,N_170,N_1089);
xor U1601 (N_1601,N_559,N_1074);
and U1602 (N_1602,N_176,N_679);
or U1603 (N_1603,N_517,N_1278);
nor U1604 (N_1604,N_842,N_610);
nor U1605 (N_1605,N_829,N_682);
or U1606 (N_1606,N_576,N_1245);
nor U1607 (N_1607,N_942,N_777);
nand U1608 (N_1608,N_1165,N_1392);
or U1609 (N_1609,N_985,N_687);
nand U1610 (N_1610,N_436,N_121);
nand U1611 (N_1611,N_430,N_653);
xnor U1612 (N_1612,N_1276,N_10);
nor U1613 (N_1613,N_1153,N_333);
nand U1614 (N_1614,N_269,N_1084);
xor U1615 (N_1615,N_1395,N_487);
nand U1616 (N_1616,N_1020,N_1054);
nand U1617 (N_1617,N_1073,N_462);
or U1618 (N_1618,N_13,N_17);
nand U1619 (N_1619,N_316,N_163);
nor U1620 (N_1620,N_1022,N_1354);
nand U1621 (N_1621,N_319,N_1267);
xor U1622 (N_1622,N_1397,N_359);
nor U1623 (N_1623,N_302,N_326);
nand U1624 (N_1624,N_1082,N_1252);
nor U1625 (N_1625,N_383,N_937);
and U1626 (N_1626,N_221,N_1442);
or U1627 (N_1627,N_553,N_22);
xnor U1628 (N_1628,N_680,N_953);
xnor U1629 (N_1629,N_910,N_877);
nand U1630 (N_1630,N_1273,N_551);
nand U1631 (N_1631,N_978,N_409);
or U1632 (N_1632,N_235,N_550);
nand U1633 (N_1633,N_493,N_280);
nand U1634 (N_1634,N_33,N_1275);
nor U1635 (N_1635,N_47,N_950);
nand U1636 (N_1636,N_1243,N_1055);
or U1637 (N_1637,N_264,N_204);
and U1638 (N_1638,N_1478,N_1280);
nor U1639 (N_1639,N_1212,N_916);
xnor U1640 (N_1640,N_543,N_1160);
nor U1641 (N_1641,N_27,N_329);
and U1642 (N_1642,N_1167,N_640);
xnor U1643 (N_1643,N_360,N_139);
nand U1644 (N_1644,N_1389,N_107);
nand U1645 (N_1645,N_180,N_1130);
nand U1646 (N_1646,N_792,N_1067);
nor U1647 (N_1647,N_633,N_1141);
or U1648 (N_1648,N_1180,N_174);
xnor U1649 (N_1649,N_1145,N_1231);
and U1650 (N_1650,N_701,N_203);
or U1651 (N_1651,N_1213,N_1372);
xor U1652 (N_1652,N_1109,N_843);
nand U1653 (N_1653,N_325,N_299);
or U1654 (N_1654,N_1185,N_683);
or U1655 (N_1655,N_437,N_1378);
xnor U1656 (N_1656,N_725,N_497);
and U1657 (N_1657,N_205,N_598);
nand U1658 (N_1658,N_1293,N_286);
nand U1659 (N_1659,N_1088,N_1044);
xor U1660 (N_1660,N_721,N_647);
nor U1661 (N_1661,N_94,N_278);
and U1662 (N_1662,N_1399,N_702);
nor U1663 (N_1663,N_26,N_751);
and U1664 (N_1664,N_766,N_1488);
and U1665 (N_1665,N_1005,N_539);
or U1666 (N_1666,N_719,N_401);
and U1667 (N_1667,N_1148,N_925);
nor U1668 (N_1668,N_600,N_770);
xnor U1669 (N_1669,N_658,N_14);
nand U1670 (N_1670,N_888,N_1356);
and U1671 (N_1671,N_1321,N_114);
nor U1672 (N_1672,N_1152,N_1159);
xor U1673 (N_1673,N_972,N_4);
and U1674 (N_1674,N_513,N_0);
nand U1675 (N_1675,N_465,N_1410);
nand U1676 (N_1676,N_630,N_1457);
or U1677 (N_1677,N_1241,N_1011);
and U1678 (N_1678,N_710,N_1113);
nand U1679 (N_1679,N_1087,N_1227);
or U1680 (N_1680,N_1146,N_772);
nand U1681 (N_1681,N_1162,N_963);
xnor U1682 (N_1682,N_748,N_674);
and U1683 (N_1683,N_455,N_1223);
or U1684 (N_1684,N_214,N_1199);
nand U1685 (N_1685,N_230,N_255);
or U1686 (N_1686,N_1459,N_272);
and U1687 (N_1687,N_191,N_1398);
and U1688 (N_1688,N_81,N_1137);
or U1689 (N_1689,N_605,N_259);
and U1690 (N_1690,N_195,N_446);
nor U1691 (N_1691,N_620,N_1425);
or U1692 (N_1692,N_1068,N_1250);
or U1693 (N_1693,N_997,N_347);
or U1694 (N_1694,N_926,N_1229);
xor U1695 (N_1695,N_173,N_1347);
nor U1696 (N_1696,N_615,N_909);
and U1697 (N_1697,N_667,N_447);
and U1698 (N_1698,N_1115,N_880);
xor U1699 (N_1699,N_828,N_973);
nand U1700 (N_1700,N_213,N_528);
and U1701 (N_1701,N_65,N_511);
nand U1702 (N_1702,N_518,N_426);
or U1703 (N_1703,N_362,N_836);
and U1704 (N_1704,N_381,N_145);
nor U1705 (N_1705,N_780,N_177);
nand U1706 (N_1706,N_982,N_159);
and U1707 (N_1707,N_498,N_894);
xnor U1708 (N_1708,N_307,N_1370);
nand U1709 (N_1709,N_1487,N_488);
xor U1710 (N_1710,N_626,N_893);
nand U1711 (N_1711,N_1147,N_861);
nand U1712 (N_1712,N_234,N_781);
and U1713 (N_1713,N_983,N_375);
xor U1714 (N_1714,N_21,N_1226);
and U1715 (N_1715,N_438,N_495);
nor U1716 (N_1716,N_496,N_1343);
xnor U1717 (N_1717,N_941,N_569);
and U1718 (N_1718,N_1460,N_645);
nand U1719 (N_1719,N_1219,N_1451);
or U1720 (N_1720,N_202,N_571);
nand U1721 (N_1721,N_1432,N_1262);
and U1722 (N_1722,N_1063,N_1483);
xor U1723 (N_1723,N_698,N_897);
nor U1724 (N_1724,N_1097,N_500);
nor U1725 (N_1725,N_757,N_85);
xnor U1726 (N_1726,N_611,N_1176);
xnor U1727 (N_1727,N_801,N_1375);
nor U1728 (N_1728,N_1448,N_1014);
and U1729 (N_1729,N_262,N_62);
and U1730 (N_1730,N_122,N_1221);
nand U1731 (N_1731,N_1324,N_476);
nand U1732 (N_1732,N_416,N_1393);
nand U1733 (N_1733,N_1239,N_75);
and U1734 (N_1734,N_584,N_736);
and U1735 (N_1735,N_1492,N_1305);
nand U1736 (N_1736,N_1446,N_477);
nand U1737 (N_1737,N_964,N_1462);
or U1738 (N_1738,N_1463,N_89);
and U1739 (N_1739,N_1178,N_1150);
or U1740 (N_1740,N_1482,N_1365);
and U1741 (N_1741,N_1313,N_570);
or U1742 (N_1742,N_283,N_838);
nor U1743 (N_1743,N_256,N_466);
and U1744 (N_1744,N_1186,N_873);
xor U1745 (N_1745,N_954,N_815);
or U1746 (N_1746,N_850,N_28);
or U1747 (N_1747,N_402,N_566);
xor U1748 (N_1748,N_625,N_872);
xor U1749 (N_1749,N_1469,N_1042);
xnor U1750 (N_1750,N_862,N_835);
and U1751 (N_1751,N_1099,N_546);
or U1752 (N_1752,N_419,N_529);
nand U1753 (N_1753,N_454,N_367);
nand U1754 (N_1754,N_300,N_110);
nand U1755 (N_1755,N_527,N_392);
and U1756 (N_1756,N_568,N_445);
nor U1757 (N_1757,N_1182,N_443);
xnor U1758 (N_1758,N_715,N_1009);
or U1759 (N_1759,N_1329,N_323);
nand U1760 (N_1760,N_750,N_397);
nand U1761 (N_1761,N_429,N_714);
nand U1762 (N_1762,N_990,N_902);
or U1763 (N_1763,N_812,N_1363);
and U1764 (N_1764,N_1288,N_998);
and U1765 (N_1765,N_924,N_847);
nor U1766 (N_1766,N_1331,N_220);
nand U1767 (N_1767,N_148,N_515);
nor U1768 (N_1768,N_726,N_467);
or U1769 (N_1769,N_1479,N_669);
xnor U1770 (N_1770,N_1386,N_258);
nand U1771 (N_1771,N_723,N_297);
or U1772 (N_1772,N_1353,N_769);
or U1773 (N_1773,N_1359,N_1349);
and U1774 (N_1774,N_197,N_797);
xnor U1775 (N_1775,N_1207,N_879);
nor U1776 (N_1776,N_175,N_1202);
xor U1777 (N_1777,N_284,N_1081);
xor U1778 (N_1778,N_578,N_222);
nor U1779 (N_1779,N_273,N_510);
and U1780 (N_1780,N_1156,N_629);
nand U1781 (N_1781,N_414,N_1297);
xor U1782 (N_1782,N_91,N_1317);
and U1783 (N_1783,N_210,N_34);
and U1784 (N_1784,N_875,N_749);
and U1785 (N_1785,N_1025,N_1234);
xor U1786 (N_1786,N_811,N_1495);
and U1787 (N_1787,N_1477,N_646);
nor U1788 (N_1788,N_434,N_1345);
and U1789 (N_1789,N_1332,N_718);
and U1790 (N_1790,N_186,N_798);
or U1791 (N_1791,N_544,N_1205);
or U1792 (N_1792,N_1249,N_484);
nor U1793 (N_1793,N_639,N_981);
xor U1794 (N_1794,N_733,N_1421);
nor U1795 (N_1795,N_503,N_263);
xor U1796 (N_1796,N_1322,N_79);
nor U1797 (N_1797,N_330,N_223);
nand U1798 (N_1798,N_596,N_730);
xnor U1799 (N_1799,N_677,N_839);
and U1800 (N_1800,N_1420,N_1406);
nor U1801 (N_1801,N_1140,N_1021);
nand U1802 (N_1802,N_1200,N_166);
xor U1803 (N_1803,N_236,N_469);
nor U1804 (N_1804,N_472,N_308);
xnor U1805 (N_1805,N_490,N_882);
nand U1806 (N_1806,N_934,N_602);
nor U1807 (N_1807,N_1224,N_20);
xor U1808 (N_1808,N_636,N_537);
or U1809 (N_1809,N_460,N_1075);
nor U1810 (N_1810,N_705,N_1050);
xnor U1811 (N_1811,N_825,N_1002);
nand U1812 (N_1812,N_212,N_1255);
xnor U1813 (N_1813,N_831,N_1045);
nor U1814 (N_1814,N_35,N_151);
xnor U1815 (N_1815,N_157,N_318);
nor U1816 (N_1816,N_587,N_356);
and U1817 (N_1817,N_999,N_1222);
or U1818 (N_1818,N_475,N_1105);
nand U1819 (N_1819,N_1489,N_1476);
nand U1820 (N_1820,N_604,N_993);
xnor U1821 (N_1821,N_975,N_1183);
nor U1822 (N_1822,N_334,N_1340);
or U1823 (N_1823,N_12,N_761);
nor U1824 (N_1824,N_337,N_485);
nand U1825 (N_1825,N_1134,N_849);
xor U1826 (N_1826,N_108,N_1010);
xnor U1827 (N_1827,N_470,N_374);
nor U1828 (N_1828,N_822,N_991);
nor U1829 (N_1829,N_508,N_783);
or U1830 (N_1830,N_1121,N_137);
or U1831 (N_1831,N_23,N_100);
or U1832 (N_1832,N_734,N_304);
or U1833 (N_1833,N_1351,N_1290);
or U1834 (N_1834,N_403,N_891);
and U1835 (N_1835,N_711,N_452);
nand U1836 (N_1836,N_1191,N_1220);
xor U1837 (N_1837,N_96,N_83);
or U1838 (N_1838,N_420,N_874);
nand U1839 (N_1839,N_225,N_632);
or U1840 (N_1840,N_1376,N_384);
nand U1841 (N_1841,N_399,N_192);
nor U1842 (N_1842,N_483,N_1077);
nand U1843 (N_1843,N_855,N_716);
nor U1844 (N_1844,N_340,N_685);
nor U1845 (N_1845,N_866,N_1066);
or U1846 (N_1846,N_1362,N_512);
or U1847 (N_1847,N_1428,N_1274);
and U1848 (N_1848,N_1132,N_1166);
or U1849 (N_1849,N_722,N_642);
or U1850 (N_1850,N_1449,N_80);
and U1851 (N_1851,N_1209,N_728);
nor U1852 (N_1852,N_1471,N_50);
xor U1853 (N_1853,N_643,N_987);
nand U1854 (N_1854,N_63,N_1440);
or U1855 (N_1855,N_694,N_135);
nand U1856 (N_1856,N_1327,N_654);
nand U1857 (N_1857,N_773,N_1107);
and U1858 (N_1858,N_379,N_621);
nor U1859 (N_1859,N_624,N_1458);
nand U1860 (N_1860,N_1024,N_668);
nand U1861 (N_1861,N_1323,N_298);
or U1862 (N_1862,N_281,N_1110);
or U1863 (N_1863,N_489,N_826);
xnor U1864 (N_1864,N_1093,N_1315);
nor U1865 (N_1865,N_922,N_1493);
nor U1866 (N_1866,N_1427,N_1026);
and U1867 (N_1867,N_917,N_944);
or U1868 (N_1868,N_720,N_54);
xor U1869 (N_1869,N_457,N_301);
and U1870 (N_1870,N_1265,N_494);
nand U1871 (N_1871,N_1098,N_92);
xnor U1872 (N_1872,N_184,N_984);
and U1873 (N_1873,N_523,N_179);
xnor U1874 (N_1874,N_740,N_724);
nand U1875 (N_1875,N_856,N_276);
xor U1876 (N_1876,N_413,N_38);
or U1877 (N_1877,N_55,N_169);
xnor U1878 (N_1878,N_1218,N_398);
or U1879 (N_1879,N_463,N_29);
or U1880 (N_1880,N_651,N_1038);
and U1881 (N_1881,N_863,N_787);
nor U1882 (N_1882,N_3,N_19);
nor U1883 (N_1883,N_285,N_1102);
or U1884 (N_1884,N_1157,N_933);
nand U1885 (N_1885,N_627,N_1117);
xnor U1886 (N_1886,N_1233,N_295);
nand U1887 (N_1887,N_919,N_1311);
and U1888 (N_1888,N_706,N_143);
xor U1889 (N_1889,N_1187,N_147);
nand U1890 (N_1890,N_42,N_1371);
and U1891 (N_1891,N_1195,N_1289);
xnor U1892 (N_1892,N_775,N_423);
xnor U1893 (N_1893,N_1175,N_742);
xnor U1894 (N_1894,N_1342,N_1337);
or U1895 (N_1895,N_1078,N_129);
and U1896 (N_1896,N_731,N_737);
nand U1897 (N_1897,N_480,N_1346);
or U1898 (N_1898,N_806,N_823);
nand U1899 (N_1899,N_817,N_1374);
xor U1900 (N_1900,N_1416,N_1411);
nand U1901 (N_1901,N_185,N_1296);
nand U1902 (N_1902,N_758,N_479);
or U1903 (N_1903,N_575,N_1308);
xnor U1904 (N_1904,N_1441,N_453);
xor U1905 (N_1905,N_1270,N_120);
nor U1906 (N_1906,N_659,N_907);
nor U1907 (N_1907,N_655,N_1256);
or U1908 (N_1908,N_946,N_116);
nand U1909 (N_1909,N_1260,N_1430);
xnor U1910 (N_1910,N_860,N_1064);
or U1911 (N_1911,N_1053,N_74);
xnor U1912 (N_1912,N_232,N_967);
xor U1913 (N_1913,N_73,N_168);
and U1914 (N_1914,N_1383,N_439);
nor U1915 (N_1915,N_1465,N_763);
nor U1916 (N_1916,N_1072,N_231);
xor U1917 (N_1917,N_421,N_1129);
or U1918 (N_1918,N_593,N_365);
nor U1919 (N_1919,N_601,N_1360);
xnor U1920 (N_1920,N_664,N_1358);
or U1921 (N_1921,N_914,N_638);
xnor U1922 (N_1922,N_1257,N_660);
xnor U1923 (N_1923,N_1325,N_18);
and U1924 (N_1924,N_541,N_391);
nor U1925 (N_1925,N_1272,N_358);
or U1926 (N_1926,N_393,N_547);
and U1927 (N_1927,N_57,N_1193);
nor U1928 (N_1928,N_282,N_526);
or U1929 (N_1929,N_218,N_661);
nor U1930 (N_1930,N_932,N_328);
nor U1931 (N_1931,N_656,N_1112);
or U1932 (N_1932,N_227,N_1404);
nor U1933 (N_1933,N_410,N_118);
or U1934 (N_1934,N_1328,N_1139);
or U1935 (N_1935,N_943,N_745);
xor U1936 (N_1936,N_1135,N_778);
or U1937 (N_1937,N_1000,N_1298);
xor U1938 (N_1938,N_735,N_760);
or U1939 (N_1939,N_867,N_1266);
nand U1940 (N_1940,N_1238,N_433);
nand U1941 (N_1941,N_119,N_1136);
nor U1942 (N_1942,N_474,N_1036);
nor U1943 (N_1943,N_1071,N_574);
nor U1944 (N_1944,N_959,N_614);
nor U1945 (N_1945,N_342,N_2);
nand U1946 (N_1946,N_555,N_270);
xnor U1947 (N_1947,N_155,N_979);
nor U1948 (N_1948,N_267,N_689);
or U1949 (N_1949,N_1170,N_199);
and U1950 (N_1950,N_208,N_805);
xnor U1951 (N_1951,N_1247,N_1164);
nor U1952 (N_1952,N_449,N_77);
and U1953 (N_1953,N_390,N_149);
nor U1954 (N_1954,N_573,N_565);
xor U1955 (N_1955,N_913,N_696);
and U1956 (N_1956,N_804,N_857);
nor U1957 (N_1957,N_803,N_744);
nor U1958 (N_1958,N_216,N_684);
nor U1959 (N_1959,N_809,N_233);
nor U1960 (N_1960,N_1368,N_1450);
and U1961 (N_1961,N_1434,N_904);
or U1962 (N_1962,N_971,N_291);
xnor U1963 (N_1963,N_1481,N_59);
or U1964 (N_1964,N_1118,N_644);
nor U1965 (N_1965,N_790,N_802);
or U1966 (N_1966,N_1437,N_977);
or U1967 (N_1967,N_275,N_1125);
and U1968 (N_1968,N_344,N_1095);
and U1969 (N_1969,N_793,N_789);
or U1970 (N_1970,N_265,N_196);
nor U1971 (N_1971,N_1391,N_921);
and U1972 (N_1972,N_348,N_594);
nand U1973 (N_1973,N_799,N_951);
and U1974 (N_1974,N_562,N_961);
xnor U1975 (N_1975,N_1069,N_868);
xnor U1976 (N_1976,N_165,N_31);
xnor U1977 (N_1977,N_386,N_530);
xnor U1978 (N_1978,N_912,N_818);
xor U1979 (N_1979,N_492,N_955);
or U1980 (N_1980,N_274,N_1413);
or U1981 (N_1981,N_322,N_782);
nor U1982 (N_1982,N_1380,N_1091);
xnor U1983 (N_1983,N_821,N_846);
or U1984 (N_1984,N_692,N_76);
nand U1985 (N_1985,N_899,N_404);
nor U1986 (N_1986,N_435,N_1034);
and U1987 (N_1987,N_1085,N_688);
xnor U1988 (N_1988,N_908,N_1302);
and U1989 (N_1989,N_878,N_548);
nand U1990 (N_1990,N_697,N_1444);
and U1991 (N_1991,N_327,N_69);
xor U1992 (N_1992,N_952,N_1486);
nand U1993 (N_1993,N_244,N_747);
nor U1994 (N_1994,N_1079,N_369);
nor U1995 (N_1995,N_1248,N_732);
or U1996 (N_1996,N_957,N_1122);
xor U1997 (N_1997,N_363,N_1491);
and U1998 (N_1998,N_759,N_583);
nand U1999 (N_1999,N_881,N_331);
nor U2000 (N_2000,N_1138,N_317);
or U2001 (N_2001,N_691,N_1304);
and U2002 (N_2002,N_613,N_949);
nor U2003 (N_2003,N_1083,N_1350);
nor U2004 (N_2004,N_753,N_586);
nor U2005 (N_2005,N_986,N_1361);
nand U2006 (N_2006,N_249,N_380);
and U2007 (N_2007,N_906,N_60);
nor U2008 (N_2008,N_948,N_1381);
xnor U2009 (N_2009,N_927,N_969);
nand U2010 (N_2010,N_852,N_905);
and U2011 (N_2011,N_1377,N_109);
nor U2012 (N_2012,N_125,N_756);
nand U2013 (N_2013,N_585,N_1408);
and U2014 (N_2014,N_310,N_87);
nand U2015 (N_2015,N_785,N_172);
xnor U2016 (N_2016,N_1385,N_1336);
and U2017 (N_2017,N_1008,N_938);
nor U2018 (N_2018,N_597,N_552);
nor U2019 (N_2019,N_1294,N_1387);
and U2020 (N_2020,N_156,N_1027);
nand U2021 (N_2021,N_619,N_190);
nand U2022 (N_2022,N_727,N_538);
nor U2023 (N_2023,N_1418,N_1364);
and U2024 (N_2024,N_321,N_1485);
nor U2025 (N_2025,N_237,N_345);
nor U2026 (N_2026,N_670,N_1033);
and U2027 (N_2027,N_607,N_741);
nor U2028 (N_2028,N_9,N_929);
and U2029 (N_2029,N_412,N_102);
nor U2030 (N_2030,N_524,N_427);
nand U2031 (N_2031,N_366,N_502);
and U2032 (N_2032,N_1177,N_1424);
nor U2033 (N_2033,N_996,N_70);
xor U2034 (N_2034,N_1352,N_464);
xnor U2035 (N_2035,N_800,N_788);
nor U2036 (N_2036,N_1131,N_39);
and U2037 (N_2037,N_889,N_123);
and U2038 (N_2038,N_7,N_1111);
and U2039 (N_2039,N_481,N_305);
nor U2040 (N_2040,N_1384,N_471);
xor U2041 (N_2041,N_200,N_1151);
and U2042 (N_2042,N_456,N_1394);
nand U2043 (N_2043,N_1114,N_388);
or U2044 (N_2044,N_858,N_540);
and U2045 (N_2045,N_608,N_1303);
nand U2046 (N_2046,N_589,N_885);
or U2047 (N_2047,N_11,N_870);
nand U2048 (N_2048,N_980,N_1015);
nand U2049 (N_2049,N_387,N_690);
or U2050 (N_2050,N_776,N_923);
xnor U2051 (N_2051,N_845,N_1096);
nand U2052 (N_2052,N_678,N_1498);
or U2053 (N_2053,N_1174,N_408);
xor U2054 (N_2054,N_1059,N_617);
nor U2055 (N_2055,N_1040,N_520);
and U2056 (N_2056,N_641,N_960);
or U2057 (N_2057,N_1433,N_827);
nand U2058 (N_2058,N_254,N_441);
or U2059 (N_2059,N_368,N_1214);
nor U2060 (N_2060,N_673,N_332);
and U2061 (N_2061,N_1046,N_181);
and U2062 (N_2062,N_890,N_807);
nand U2063 (N_2063,N_525,N_976);
and U2064 (N_2064,N_1123,N_886);
or U2065 (N_2065,N_45,N_127);
nor U2066 (N_2066,N_506,N_713);
nor U2067 (N_2067,N_306,N_44);
xnor U2068 (N_2068,N_82,N_819);
nand U2069 (N_2069,N_339,N_343);
and U2070 (N_2070,N_1215,N_1016);
nand U2071 (N_2071,N_1211,N_813);
nand U2072 (N_2072,N_52,N_1484);
or U2073 (N_2073,N_112,N_1348);
nand U2074 (N_2074,N_1335,N_1369);
or U2075 (N_2075,N_491,N_1070);
or U2076 (N_2076,N_158,N_709);
nor U2077 (N_2077,N_131,N_1017);
and U2078 (N_2078,N_1295,N_595);
xnor U2079 (N_2079,N_962,N_97);
and U2080 (N_2080,N_1242,N_1309);
xor U2081 (N_2081,N_64,N_634);
xnor U2082 (N_2082,N_1436,N_1196);
xnor U2083 (N_2083,N_564,N_290);
or U2084 (N_2084,N_215,N_637);
xnor U2085 (N_2085,N_820,N_504);
xor U2086 (N_2086,N_183,N_373);
xor U2087 (N_2087,N_1210,N_786);
nor U2088 (N_2088,N_1466,N_417);
or U2089 (N_2089,N_1225,N_1168);
and U2090 (N_2090,N_1472,N_1494);
xor U2091 (N_2091,N_61,N_67);
xnor U2092 (N_2092,N_51,N_989);
or U2093 (N_2093,N_1403,N_5);
nand U2094 (N_2094,N_389,N_1473);
and U2095 (N_2095,N_665,N_519);
xor U2096 (N_2096,N_514,N_746);
xor U2097 (N_2097,N_1237,N_146);
and U2098 (N_2098,N_209,N_1048);
xnor U2099 (N_2099,N_124,N_1236);
nor U2100 (N_2100,N_1474,N_1253);
xnor U2101 (N_2101,N_1455,N_40);
nand U2102 (N_2102,N_88,N_649);
and U2103 (N_2103,N_357,N_1019);
xnor U2104 (N_2104,N_834,N_1244);
nor U2105 (N_2105,N_229,N_1161);
xnor U2106 (N_2106,N_15,N_895);
xor U2107 (N_2107,N_1320,N_1443);
nor U2108 (N_2108,N_1047,N_189);
or U2109 (N_2109,N_1480,N_848);
or U2110 (N_2110,N_1119,N_371);
nand U2111 (N_2111,N_1306,N_41);
or U2112 (N_2112,N_840,N_288);
xor U2113 (N_2113,N_1246,N_128);
or U2114 (N_2114,N_1415,N_884);
and U2115 (N_2115,N_1037,N_1181);
nor U2116 (N_2116,N_1409,N_58);
nor U2117 (N_2117,N_1198,N_448);
nor U2118 (N_2118,N_1172,N_346);
and U2119 (N_2119,N_1194,N_542);
and U2120 (N_2120,N_372,N_795);
nand U2121 (N_2121,N_920,N_505);
or U2122 (N_2122,N_1318,N_561);
nor U2123 (N_2123,N_499,N_1407);
and U2124 (N_2124,N_187,N_859);
nor U2125 (N_2125,N_201,N_171);
nand U2126 (N_2126,N_738,N_522);
or U2127 (N_2127,N_1269,N_1240);
nand U2128 (N_2128,N_90,N_188);
or U2129 (N_2129,N_1051,N_1004);
nor U2130 (N_2130,N_833,N_150);
xnor U2131 (N_2131,N_672,N_1326);
nor U2132 (N_2132,N_1334,N_650);
nand U2133 (N_2133,N_599,N_1490);
xnor U2134 (N_2134,N_246,N_662);
and U2135 (N_2135,N_1268,N_152);
and U2136 (N_2136,N_762,N_1467);
xnor U2137 (N_2137,N_903,N_1018);
or U2138 (N_2138,N_579,N_138);
nor U2139 (N_2139,N_16,N_1454);
nand U2140 (N_2140,N_796,N_1216);
and U2141 (N_2141,N_293,N_296);
and U2142 (N_2142,N_253,N_1013);
and U2143 (N_2143,N_1012,N_1310);
nand U2144 (N_2144,N_1287,N_1291);
or U2145 (N_2145,N_1316,N_531);
xor U2146 (N_2146,N_928,N_405);
nand U2147 (N_2147,N_810,N_582);
or U2148 (N_2148,N_1367,N_1154);
nor U2149 (N_2149,N_1475,N_1314);
or U2150 (N_2150,N_56,N_1163);
or U2151 (N_2151,N_126,N_1128);
xor U2152 (N_2152,N_1468,N_1286);
or U2153 (N_2153,N_1001,N_1400);
nor U2154 (N_2154,N_841,N_1422);
nand U2155 (N_2155,N_1203,N_71);
or U2156 (N_2156,N_1235,N_217);
nor U2157 (N_2157,N_1251,N_160);
or U2158 (N_2158,N_572,N_194);
nand U2159 (N_2159,N_1355,N_133);
xor U2160 (N_2160,N_78,N_1061);
or U2161 (N_2161,N_577,N_193);
xnor U2162 (N_2162,N_1312,N_1228);
xor U2163 (N_2163,N_461,N_238);
nand U2164 (N_2164,N_406,N_675);
nor U2165 (N_2165,N_154,N_30);
nor U2166 (N_2166,N_622,N_111);
nor U2167 (N_2167,N_257,N_364);
and U2168 (N_2168,N_1435,N_141);
nand U2169 (N_2169,N_536,N_1058);
nand U2170 (N_2170,N_1496,N_1445);
nor U2171 (N_2171,N_451,N_1144);
and U2172 (N_2172,N_1277,N_1307);
and U2173 (N_2173,N_1461,N_1261);
xnor U2174 (N_2174,N_609,N_591);
xor U2175 (N_2175,N_1217,N_1029);
xor U2176 (N_2176,N_407,N_206);
nand U2177 (N_2177,N_606,N_1116);
nor U2178 (N_2178,N_1344,N_612);
or U2179 (N_2179,N_1057,N_1197);
nor U2180 (N_2180,N_707,N_918);
or U2181 (N_2181,N_1414,N_1056);
nor U2182 (N_2182,N_966,N_631);
nor U2183 (N_2183,N_1499,N_314);
xor U2184 (N_2184,N_351,N_1100);
xor U2185 (N_2185,N_49,N_883);
nor U2186 (N_2186,N_1452,N_239);
xor U2187 (N_2187,N_752,N_1292);
and U2188 (N_2188,N_261,N_1041);
nand U2189 (N_2189,N_1003,N_103);
and U2190 (N_2190,N_968,N_931);
or U2191 (N_2191,N_336,N_663);
or U2192 (N_2192,N_1035,N_292);
nand U2193 (N_2193,N_970,N_1279);
and U2194 (N_2194,N_1497,N_1155);
xor U2195 (N_2195,N_1264,N_130);
nor U2196 (N_2196,N_1284,N_242);
nor U2197 (N_2197,N_24,N_648);
or U2198 (N_2198,N_628,N_755);
xor U2199 (N_2199,N_240,N_958);
nor U2200 (N_2200,N_1188,N_1043);
xor U2201 (N_2201,N_355,N_1092);
nor U2202 (N_2202,N_444,N_1023);
nand U2203 (N_2203,N_603,N_700);
or U2204 (N_2204,N_956,N_376);
or U2205 (N_2205,N_115,N_1300);
and U2206 (N_2206,N_901,N_424);
nor U2207 (N_2207,N_243,N_1431);
xor U2208 (N_2208,N_247,N_25);
xor U2209 (N_2209,N_1120,N_1301);
xnor U2210 (N_2210,N_1080,N_1106);
nand U2211 (N_2211,N_699,N_440);
or U2212 (N_2212,N_509,N_1402);
nor U2213 (N_2213,N_1060,N_303);
nand U2214 (N_2214,N_1470,N_666);
nor U2215 (N_2215,N_245,N_844);
and U2216 (N_2216,N_1149,N_1417);
nand U2217 (N_2217,N_560,N_1184);
xnor U2218 (N_2218,N_739,N_132);
or U2219 (N_2219,N_808,N_37);
nand U2220 (N_2220,N_93,N_1142);
xor U2221 (N_2221,N_896,N_832);
nor U2222 (N_2222,N_315,N_1357);
nand U2223 (N_2223,N_248,N_46);
nand U2224 (N_2224,N_1206,N_1439);
or U2225 (N_2225,N_676,N_370);
nor U2226 (N_2226,N_140,N_385);
and U2227 (N_2227,N_1039,N_994);
or U2228 (N_2228,N_1319,N_521);
nor U2229 (N_2229,N_1419,N_1259);
or U2230 (N_2230,N_415,N_1065);
and U2231 (N_2231,N_95,N_1232);
nand U2232 (N_2232,N_939,N_791);
or U2233 (N_2233,N_554,N_1388);
and U2234 (N_2234,N_1447,N_1341);
and U2235 (N_2235,N_117,N_312);
or U2236 (N_2236,N_871,N_335);
nand U2237 (N_2237,N_1062,N_1028);
nor U2238 (N_2238,N_864,N_1030);
nand U2239 (N_2239,N_876,N_764);
nand U2240 (N_2240,N_1271,N_501);
and U2241 (N_2241,N_865,N_900);
nor U2242 (N_2242,N_1032,N_458);
nor U2243 (N_2243,N_558,N_260);
or U2244 (N_2244,N_361,N_6);
nand U2245 (N_2245,N_1283,N_1);
or U2246 (N_2246,N_1124,N_567);
xor U2247 (N_2247,N_1006,N_324);
and U2248 (N_2248,N_1379,N_1429);
and U2249 (N_2249,N_98,N_36);
xor U2250 (N_2250,N_139,N_1088);
nor U2251 (N_2251,N_174,N_1346);
nor U2252 (N_2252,N_1086,N_1457);
and U2253 (N_2253,N_1043,N_770);
nand U2254 (N_2254,N_153,N_1143);
nor U2255 (N_2255,N_654,N_1421);
or U2256 (N_2256,N_1377,N_1161);
nor U2257 (N_2257,N_1194,N_258);
and U2258 (N_2258,N_588,N_1469);
nand U2259 (N_2259,N_456,N_640);
nor U2260 (N_2260,N_594,N_921);
or U2261 (N_2261,N_1207,N_424);
nand U2262 (N_2262,N_1029,N_846);
nor U2263 (N_2263,N_1370,N_1195);
and U2264 (N_2264,N_1127,N_714);
nand U2265 (N_2265,N_834,N_755);
xnor U2266 (N_2266,N_1404,N_958);
nor U2267 (N_2267,N_533,N_416);
xor U2268 (N_2268,N_27,N_362);
nor U2269 (N_2269,N_1250,N_66);
nand U2270 (N_2270,N_234,N_703);
nand U2271 (N_2271,N_1335,N_442);
or U2272 (N_2272,N_620,N_458);
and U2273 (N_2273,N_110,N_1250);
and U2274 (N_2274,N_1134,N_175);
nor U2275 (N_2275,N_628,N_1352);
and U2276 (N_2276,N_545,N_397);
nor U2277 (N_2277,N_303,N_1253);
or U2278 (N_2278,N_1240,N_1129);
nand U2279 (N_2279,N_1136,N_432);
nand U2280 (N_2280,N_1264,N_1275);
xor U2281 (N_2281,N_413,N_14);
or U2282 (N_2282,N_220,N_445);
and U2283 (N_2283,N_956,N_1138);
or U2284 (N_2284,N_178,N_273);
nand U2285 (N_2285,N_1078,N_28);
or U2286 (N_2286,N_1221,N_278);
nand U2287 (N_2287,N_1346,N_141);
nand U2288 (N_2288,N_580,N_1202);
and U2289 (N_2289,N_1457,N_736);
xor U2290 (N_2290,N_993,N_1041);
nor U2291 (N_2291,N_890,N_290);
nor U2292 (N_2292,N_1214,N_526);
xor U2293 (N_2293,N_48,N_112);
or U2294 (N_2294,N_30,N_1223);
nor U2295 (N_2295,N_917,N_1440);
xor U2296 (N_2296,N_1202,N_265);
or U2297 (N_2297,N_683,N_1402);
and U2298 (N_2298,N_1261,N_1029);
or U2299 (N_2299,N_242,N_783);
and U2300 (N_2300,N_1113,N_149);
xor U2301 (N_2301,N_1232,N_1040);
xnor U2302 (N_2302,N_1250,N_1348);
nand U2303 (N_2303,N_107,N_900);
nand U2304 (N_2304,N_928,N_594);
and U2305 (N_2305,N_293,N_861);
or U2306 (N_2306,N_837,N_368);
nand U2307 (N_2307,N_1270,N_852);
and U2308 (N_2308,N_394,N_1272);
nor U2309 (N_2309,N_230,N_431);
and U2310 (N_2310,N_1112,N_523);
or U2311 (N_2311,N_1489,N_352);
or U2312 (N_2312,N_1473,N_1303);
and U2313 (N_2313,N_1492,N_77);
xor U2314 (N_2314,N_593,N_1150);
xor U2315 (N_2315,N_181,N_944);
or U2316 (N_2316,N_913,N_1375);
nor U2317 (N_2317,N_270,N_92);
xnor U2318 (N_2318,N_1067,N_621);
nor U2319 (N_2319,N_976,N_1223);
and U2320 (N_2320,N_1104,N_737);
xnor U2321 (N_2321,N_459,N_981);
or U2322 (N_2322,N_1143,N_646);
nand U2323 (N_2323,N_274,N_223);
and U2324 (N_2324,N_1379,N_884);
nor U2325 (N_2325,N_725,N_38);
and U2326 (N_2326,N_431,N_100);
or U2327 (N_2327,N_1453,N_585);
or U2328 (N_2328,N_214,N_1374);
xnor U2329 (N_2329,N_21,N_109);
nand U2330 (N_2330,N_275,N_606);
or U2331 (N_2331,N_492,N_1067);
nand U2332 (N_2332,N_1154,N_1067);
xnor U2333 (N_2333,N_1046,N_618);
nor U2334 (N_2334,N_1174,N_1435);
or U2335 (N_2335,N_721,N_188);
xnor U2336 (N_2336,N_571,N_715);
nand U2337 (N_2337,N_1323,N_798);
nor U2338 (N_2338,N_1495,N_40);
xnor U2339 (N_2339,N_104,N_847);
xnor U2340 (N_2340,N_956,N_982);
nor U2341 (N_2341,N_968,N_1331);
nor U2342 (N_2342,N_362,N_1173);
nand U2343 (N_2343,N_633,N_1280);
xnor U2344 (N_2344,N_977,N_83);
xnor U2345 (N_2345,N_1310,N_482);
or U2346 (N_2346,N_1496,N_1009);
and U2347 (N_2347,N_594,N_918);
nor U2348 (N_2348,N_1420,N_575);
xor U2349 (N_2349,N_966,N_793);
and U2350 (N_2350,N_122,N_546);
nor U2351 (N_2351,N_57,N_331);
and U2352 (N_2352,N_77,N_913);
nor U2353 (N_2353,N_431,N_316);
nand U2354 (N_2354,N_1221,N_724);
nor U2355 (N_2355,N_268,N_102);
nand U2356 (N_2356,N_89,N_358);
or U2357 (N_2357,N_472,N_612);
or U2358 (N_2358,N_637,N_707);
xor U2359 (N_2359,N_231,N_1488);
or U2360 (N_2360,N_656,N_317);
xnor U2361 (N_2361,N_1189,N_344);
and U2362 (N_2362,N_506,N_76);
xnor U2363 (N_2363,N_1415,N_119);
nand U2364 (N_2364,N_650,N_877);
or U2365 (N_2365,N_438,N_176);
or U2366 (N_2366,N_742,N_353);
nand U2367 (N_2367,N_131,N_1366);
xor U2368 (N_2368,N_1451,N_919);
xor U2369 (N_2369,N_744,N_118);
nand U2370 (N_2370,N_395,N_25);
nand U2371 (N_2371,N_188,N_1298);
nor U2372 (N_2372,N_233,N_410);
nand U2373 (N_2373,N_393,N_720);
or U2374 (N_2374,N_1003,N_1124);
xnor U2375 (N_2375,N_1236,N_158);
and U2376 (N_2376,N_1279,N_1281);
nor U2377 (N_2377,N_142,N_470);
nor U2378 (N_2378,N_1011,N_469);
or U2379 (N_2379,N_488,N_66);
xnor U2380 (N_2380,N_660,N_111);
nand U2381 (N_2381,N_687,N_1272);
xor U2382 (N_2382,N_346,N_839);
and U2383 (N_2383,N_574,N_1473);
and U2384 (N_2384,N_1048,N_1071);
nor U2385 (N_2385,N_993,N_1406);
and U2386 (N_2386,N_1352,N_1006);
nand U2387 (N_2387,N_1392,N_727);
xnor U2388 (N_2388,N_557,N_1018);
nor U2389 (N_2389,N_955,N_1035);
or U2390 (N_2390,N_1094,N_1363);
and U2391 (N_2391,N_476,N_500);
nand U2392 (N_2392,N_1340,N_1480);
xor U2393 (N_2393,N_1003,N_823);
and U2394 (N_2394,N_438,N_1333);
or U2395 (N_2395,N_1361,N_497);
nor U2396 (N_2396,N_777,N_689);
nand U2397 (N_2397,N_1212,N_1326);
nand U2398 (N_2398,N_863,N_625);
and U2399 (N_2399,N_248,N_1297);
nand U2400 (N_2400,N_1089,N_1210);
xor U2401 (N_2401,N_421,N_403);
or U2402 (N_2402,N_1295,N_924);
nor U2403 (N_2403,N_1339,N_1193);
and U2404 (N_2404,N_438,N_1067);
nor U2405 (N_2405,N_245,N_1002);
and U2406 (N_2406,N_896,N_665);
nand U2407 (N_2407,N_99,N_1071);
xor U2408 (N_2408,N_1242,N_763);
nor U2409 (N_2409,N_914,N_330);
nor U2410 (N_2410,N_892,N_849);
or U2411 (N_2411,N_452,N_1441);
nand U2412 (N_2412,N_1172,N_97);
nand U2413 (N_2413,N_1408,N_102);
nand U2414 (N_2414,N_437,N_528);
and U2415 (N_2415,N_292,N_818);
xor U2416 (N_2416,N_453,N_1282);
and U2417 (N_2417,N_478,N_858);
nand U2418 (N_2418,N_1370,N_36);
nor U2419 (N_2419,N_448,N_1383);
nand U2420 (N_2420,N_95,N_531);
and U2421 (N_2421,N_673,N_856);
nor U2422 (N_2422,N_775,N_1267);
and U2423 (N_2423,N_1128,N_847);
nand U2424 (N_2424,N_71,N_466);
nand U2425 (N_2425,N_1063,N_435);
xor U2426 (N_2426,N_212,N_91);
nand U2427 (N_2427,N_1348,N_357);
nor U2428 (N_2428,N_961,N_1064);
or U2429 (N_2429,N_593,N_864);
nand U2430 (N_2430,N_1402,N_806);
nor U2431 (N_2431,N_1267,N_1005);
and U2432 (N_2432,N_611,N_371);
xor U2433 (N_2433,N_531,N_404);
and U2434 (N_2434,N_457,N_614);
and U2435 (N_2435,N_760,N_1257);
or U2436 (N_2436,N_669,N_1138);
or U2437 (N_2437,N_1224,N_648);
nand U2438 (N_2438,N_857,N_434);
and U2439 (N_2439,N_243,N_1354);
or U2440 (N_2440,N_481,N_1119);
nor U2441 (N_2441,N_187,N_1331);
and U2442 (N_2442,N_1430,N_951);
xor U2443 (N_2443,N_1428,N_1305);
or U2444 (N_2444,N_1321,N_586);
xnor U2445 (N_2445,N_175,N_7);
xor U2446 (N_2446,N_806,N_346);
nor U2447 (N_2447,N_540,N_1093);
nor U2448 (N_2448,N_171,N_454);
or U2449 (N_2449,N_676,N_823);
nand U2450 (N_2450,N_745,N_430);
nor U2451 (N_2451,N_288,N_737);
and U2452 (N_2452,N_751,N_900);
nand U2453 (N_2453,N_16,N_586);
and U2454 (N_2454,N_1083,N_505);
nor U2455 (N_2455,N_1395,N_974);
and U2456 (N_2456,N_1492,N_573);
nor U2457 (N_2457,N_1248,N_939);
or U2458 (N_2458,N_249,N_749);
nand U2459 (N_2459,N_1026,N_1499);
nor U2460 (N_2460,N_199,N_169);
or U2461 (N_2461,N_1097,N_967);
xnor U2462 (N_2462,N_1157,N_1118);
xor U2463 (N_2463,N_725,N_201);
xnor U2464 (N_2464,N_658,N_1320);
nand U2465 (N_2465,N_1203,N_1058);
and U2466 (N_2466,N_530,N_1406);
or U2467 (N_2467,N_301,N_1326);
nand U2468 (N_2468,N_1467,N_259);
and U2469 (N_2469,N_407,N_67);
xor U2470 (N_2470,N_816,N_1173);
xor U2471 (N_2471,N_1322,N_328);
and U2472 (N_2472,N_90,N_569);
and U2473 (N_2473,N_219,N_1107);
xnor U2474 (N_2474,N_291,N_1176);
and U2475 (N_2475,N_1347,N_561);
xnor U2476 (N_2476,N_160,N_1451);
nor U2477 (N_2477,N_1205,N_1225);
xnor U2478 (N_2478,N_472,N_1162);
and U2479 (N_2479,N_260,N_309);
nor U2480 (N_2480,N_745,N_724);
nand U2481 (N_2481,N_799,N_119);
or U2482 (N_2482,N_602,N_191);
xnor U2483 (N_2483,N_1085,N_1474);
nor U2484 (N_2484,N_466,N_342);
and U2485 (N_2485,N_1097,N_1234);
nand U2486 (N_2486,N_1409,N_1266);
nand U2487 (N_2487,N_18,N_1089);
nor U2488 (N_2488,N_752,N_1028);
nor U2489 (N_2489,N_766,N_1413);
or U2490 (N_2490,N_754,N_450);
xnor U2491 (N_2491,N_839,N_1072);
and U2492 (N_2492,N_1309,N_1308);
nand U2493 (N_2493,N_920,N_516);
xnor U2494 (N_2494,N_753,N_293);
nor U2495 (N_2495,N_668,N_819);
and U2496 (N_2496,N_1228,N_298);
and U2497 (N_2497,N_1192,N_1067);
and U2498 (N_2498,N_119,N_996);
and U2499 (N_2499,N_48,N_912);
or U2500 (N_2500,N_71,N_1486);
nor U2501 (N_2501,N_90,N_1205);
nor U2502 (N_2502,N_843,N_1454);
and U2503 (N_2503,N_1329,N_1166);
nor U2504 (N_2504,N_717,N_1313);
xnor U2505 (N_2505,N_1185,N_383);
xnor U2506 (N_2506,N_159,N_908);
nor U2507 (N_2507,N_583,N_666);
nand U2508 (N_2508,N_833,N_1189);
and U2509 (N_2509,N_1175,N_944);
and U2510 (N_2510,N_188,N_922);
xor U2511 (N_2511,N_1251,N_1418);
xnor U2512 (N_2512,N_1315,N_926);
or U2513 (N_2513,N_684,N_179);
and U2514 (N_2514,N_940,N_1043);
or U2515 (N_2515,N_321,N_1195);
or U2516 (N_2516,N_1248,N_51);
and U2517 (N_2517,N_1009,N_986);
nor U2518 (N_2518,N_786,N_1417);
xor U2519 (N_2519,N_1393,N_230);
xnor U2520 (N_2520,N_1168,N_92);
nor U2521 (N_2521,N_326,N_683);
nor U2522 (N_2522,N_1416,N_750);
xnor U2523 (N_2523,N_943,N_982);
xnor U2524 (N_2524,N_169,N_90);
and U2525 (N_2525,N_851,N_803);
nand U2526 (N_2526,N_1406,N_1460);
nor U2527 (N_2527,N_1306,N_177);
nand U2528 (N_2528,N_439,N_372);
xor U2529 (N_2529,N_927,N_722);
and U2530 (N_2530,N_715,N_526);
or U2531 (N_2531,N_330,N_1262);
and U2532 (N_2532,N_457,N_1277);
or U2533 (N_2533,N_1418,N_1039);
xor U2534 (N_2534,N_459,N_808);
nor U2535 (N_2535,N_287,N_263);
nor U2536 (N_2536,N_774,N_938);
nor U2537 (N_2537,N_1033,N_431);
nor U2538 (N_2538,N_691,N_61);
nand U2539 (N_2539,N_1171,N_587);
or U2540 (N_2540,N_168,N_494);
xor U2541 (N_2541,N_1056,N_704);
xnor U2542 (N_2542,N_521,N_1499);
nand U2543 (N_2543,N_1109,N_1298);
and U2544 (N_2544,N_651,N_979);
nor U2545 (N_2545,N_1210,N_609);
or U2546 (N_2546,N_479,N_660);
and U2547 (N_2547,N_1068,N_1178);
nor U2548 (N_2548,N_1382,N_279);
nand U2549 (N_2549,N_941,N_963);
and U2550 (N_2550,N_206,N_128);
xor U2551 (N_2551,N_1165,N_1327);
nand U2552 (N_2552,N_1214,N_370);
and U2553 (N_2553,N_1241,N_154);
nand U2554 (N_2554,N_1064,N_96);
or U2555 (N_2555,N_650,N_1274);
or U2556 (N_2556,N_867,N_883);
nand U2557 (N_2557,N_615,N_24);
and U2558 (N_2558,N_784,N_683);
nor U2559 (N_2559,N_621,N_1253);
xnor U2560 (N_2560,N_1258,N_75);
nand U2561 (N_2561,N_97,N_1019);
nor U2562 (N_2562,N_522,N_911);
and U2563 (N_2563,N_487,N_416);
or U2564 (N_2564,N_577,N_345);
and U2565 (N_2565,N_622,N_1268);
or U2566 (N_2566,N_1185,N_57);
nand U2567 (N_2567,N_1061,N_979);
or U2568 (N_2568,N_148,N_1022);
nand U2569 (N_2569,N_417,N_1073);
xor U2570 (N_2570,N_175,N_1310);
nor U2571 (N_2571,N_50,N_510);
nor U2572 (N_2572,N_1435,N_1002);
nor U2573 (N_2573,N_822,N_1048);
nor U2574 (N_2574,N_771,N_1252);
nand U2575 (N_2575,N_814,N_858);
nand U2576 (N_2576,N_861,N_560);
and U2577 (N_2577,N_1381,N_928);
nand U2578 (N_2578,N_856,N_1368);
and U2579 (N_2579,N_702,N_889);
xor U2580 (N_2580,N_1094,N_1147);
nor U2581 (N_2581,N_1198,N_717);
nor U2582 (N_2582,N_1151,N_831);
nand U2583 (N_2583,N_1355,N_1389);
or U2584 (N_2584,N_642,N_144);
nand U2585 (N_2585,N_514,N_72);
nor U2586 (N_2586,N_967,N_661);
and U2587 (N_2587,N_1293,N_364);
nor U2588 (N_2588,N_580,N_1117);
or U2589 (N_2589,N_1339,N_951);
and U2590 (N_2590,N_442,N_1401);
nand U2591 (N_2591,N_1349,N_1467);
or U2592 (N_2592,N_998,N_304);
nand U2593 (N_2593,N_404,N_346);
nand U2594 (N_2594,N_1192,N_1188);
xor U2595 (N_2595,N_1450,N_408);
xnor U2596 (N_2596,N_1315,N_1239);
or U2597 (N_2597,N_192,N_1089);
or U2598 (N_2598,N_1061,N_92);
or U2599 (N_2599,N_1384,N_222);
or U2600 (N_2600,N_1205,N_792);
xor U2601 (N_2601,N_1141,N_505);
xor U2602 (N_2602,N_171,N_1152);
xnor U2603 (N_2603,N_1393,N_1491);
xor U2604 (N_2604,N_68,N_1459);
nand U2605 (N_2605,N_420,N_854);
or U2606 (N_2606,N_113,N_1053);
nand U2607 (N_2607,N_1255,N_106);
and U2608 (N_2608,N_606,N_1071);
xnor U2609 (N_2609,N_520,N_1084);
and U2610 (N_2610,N_1463,N_1152);
and U2611 (N_2611,N_1206,N_936);
or U2612 (N_2612,N_333,N_354);
nor U2613 (N_2613,N_844,N_1213);
nor U2614 (N_2614,N_297,N_607);
nor U2615 (N_2615,N_598,N_1082);
nand U2616 (N_2616,N_635,N_1209);
nor U2617 (N_2617,N_1288,N_410);
or U2618 (N_2618,N_990,N_29);
or U2619 (N_2619,N_352,N_909);
xor U2620 (N_2620,N_1478,N_1262);
nor U2621 (N_2621,N_420,N_536);
or U2622 (N_2622,N_1264,N_1122);
or U2623 (N_2623,N_889,N_600);
nor U2624 (N_2624,N_70,N_1298);
or U2625 (N_2625,N_1382,N_322);
and U2626 (N_2626,N_1289,N_669);
nand U2627 (N_2627,N_1241,N_486);
and U2628 (N_2628,N_899,N_203);
and U2629 (N_2629,N_978,N_749);
xor U2630 (N_2630,N_1364,N_700);
nand U2631 (N_2631,N_294,N_775);
or U2632 (N_2632,N_1118,N_114);
nor U2633 (N_2633,N_794,N_450);
nor U2634 (N_2634,N_205,N_1026);
xor U2635 (N_2635,N_1256,N_1072);
nor U2636 (N_2636,N_1260,N_464);
or U2637 (N_2637,N_134,N_368);
xnor U2638 (N_2638,N_107,N_892);
xor U2639 (N_2639,N_207,N_1043);
nor U2640 (N_2640,N_1088,N_648);
and U2641 (N_2641,N_619,N_1293);
or U2642 (N_2642,N_188,N_151);
xor U2643 (N_2643,N_1180,N_1327);
or U2644 (N_2644,N_542,N_823);
xor U2645 (N_2645,N_1137,N_373);
nand U2646 (N_2646,N_1432,N_865);
or U2647 (N_2647,N_629,N_689);
or U2648 (N_2648,N_1097,N_975);
or U2649 (N_2649,N_439,N_650);
nand U2650 (N_2650,N_1193,N_742);
xor U2651 (N_2651,N_645,N_1276);
nor U2652 (N_2652,N_379,N_47);
nor U2653 (N_2653,N_1031,N_1345);
and U2654 (N_2654,N_400,N_662);
nor U2655 (N_2655,N_528,N_1424);
nor U2656 (N_2656,N_1485,N_384);
nand U2657 (N_2657,N_29,N_1351);
and U2658 (N_2658,N_890,N_518);
xor U2659 (N_2659,N_237,N_220);
nor U2660 (N_2660,N_1368,N_201);
nand U2661 (N_2661,N_1185,N_214);
and U2662 (N_2662,N_758,N_627);
or U2663 (N_2663,N_1261,N_361);
nand U2664 (N_2664,N_657,N_1307);
nor U2665 (N_2665,N_492,N_840);
and U2666 (N_2666,N_1212,N_546);
and U2667 (N_2667,N_653,N_143);
nand U2668 (N_2668,N_1164,N_192);
nor U2669 (N_2669,N_11,N_1067);
xnor U2670 (N_2670,N_1255,N_1326);
and U2671 (N_2671,N_1290,N_255);
and U2672 (N_2672,N_749,N_188);
and U2673 (N_2673,N_266,N_207);
or U2674 (N_2674,N_1221,N_1141);
and U2675 (N_2675,N_1466,N_242);
or U2676 (N_2676,N_353,N_940);
or U2677 (N_2677,N_1267,N_941);
and U2678 (N_2678,N_378,N_1029);
nor U2679 (N_2679,N_438,N_918);
xnor U2680 (N_2680,N_463,N_122);
xor U2681 (N_2681,N_213,N_1321);
nor U2682 (N_2682,N_461,N_540);
xnor U2683 (N_2683,N_519,N_1173);
nand U2684 (N_2684,N_1219,N_1318);
nand U2685 (N_2685,N_112,N_260);
nand U2686 (N_2686,N_1278,N_1397);
and U2687 (N_2687,N_214,N_756);
and U2688 (N_2688,N_1380,N_1429);
and U2689 (N_2689,N_1419,N_981);
nand U2690 (N_2690,N_1425,N_819);
or U2691 (N_2691,N_1256,N_314);
xnor U2692 (N_2692,N_1303,N_28);
or U2693 (N_2693,N_236,N_472);
nor U2694 (N_2694,N_934,N_547);
xnor U2695 (N_2695,N_405,N_988);
xor U2696 (N_2696,N_36,N_1224);
and U2697 (N_2697,N_861,N_376);
nor U2698 (N_2698,N_883,N_873);
xnor U2699 (N_2699,N_546,N_1055);
or U2700 (N_2700,N_414,N_1301);
nand U2701 (N_2701,N_1220,N_878);
and U2702 (N_2702,N_700,N_1162);
nand U2703 (N_2703,N_443,N_1435);
nor U2704 (N_2704,N_544,N_419);
xor U2705 (N_2705,N_540,N_1065);
xnor U2706 (N_2706,N_1086,N_242);
nand U2707 (N_2707,N_557,N_709);
and U2708 (N_2708,N_297,N_1267);
xnor U2709 (N_2709,N_1105,N_37);
and U2710 (N_2710,N_112,N_447);
nand U2711 (N_2711,N_59,N_355);
nand U2712 (N_2712,N_698,N_603);
xor U2713 (N_2713,N_716,N_1247);
nor U2714 (N_2714,N_498,N_1257);
nand U2715 (N_2715,N_140,N_187);
xnor U2716 (N_2716,N_934,N_82);
or U2717 (N_2717,N_478,N_1373);
nand U2718 (N_2718,N_913,N_1202);
and U2719 (N_2719,N_1355,N_1232);
xor U2720 (N_2720,N_1214,N_347);
nand U2721 (N_2721,N_1219,N_121);
or U2722 (N_2722,N_63,N_684);
xnor U2723 (N_2723,N_542,N_127);
nand U2724 (N_2724,N_66,N_995);
nand U2725 (N_2725,N_356,N_408);
nor U2726 (N_2726,N_1033,N_792);
nand U2727 (N_2727,N_929,N_88);
and U2728 (N_2728,N_728,N_1442);
or U2729 (N_2729,N_1107,N_1408);
xnor U2730 (N_2730,N_362,N_1172);
xnor U2731 (N_2731,N_1080,N_767);
xnor U2732 (N_2732,N_1437,N_1344);
and U2733 (N_2733,N_401,N_1276);
xnor U2734 (N_2734,N_614,N_688);
nand U2735 (N_2735,N_73,N_1123);
or U2736 (N_2736,N_730,N_283);
xnor U2737 (N_2737,N_1029,N_1302);
and U2738 (N_2738,N_790,N_1487);
xnor U2739 (N_2739,N_780,N_276);
nor U2740 (N_2740,N_527,N_338);
or U2741 (N_2741,N_934,N_507);
xor U2742 (N_2742,N_1221,N_627);
or U2743 (N_2743,N_804,N_586);
and U2744 (N_2744,N_379,N_87);
nand U2745 (N_2745,N_1201,N_1169);
nand U2746 (N_2746,N_1442,N_825);
and U2747 (N_2747,N_1444,N_444);
nand U2748 (N_2748,N_1435,N_87);
nand U2749 (N_2749,N_1189,N_555);
nor U2750 (N_2750,N_833,N_413);
and U2751 (N_2751,N_495,N_449);
or U2752 (N_2752,N_105,N_535);
xnor U2753 (N_2753,N_335,N_1433);
and U2754 (N_2754,N_66,N_1108);
nor U2755 (N_2755,N_1224,N_1336);
or U2756 (N_2756,N_637,N_187);
xor U2757 (N_2757,N_297,N_559);
xor U2758 (N_2758,N_93,N_327);
and U2759 (N_2759,N_823,N_1243);
and U2760 (N_2760,N_1318,N_1138);
xnor U2761 (N_2761,N_441,N_256);
xor U2762 (N_2762,N_179,N_974);
or U2763 (N_2763,N_1097,N_1025);
nor U2764 (N_2764,N_3,N_378);
nand U2765 (N_2765,N_641,N_1317);
or U2766 (N_2766,N_150,N_93);
nor U2767 (N_2767,N_982,N_415);
nor U2768 (N_2768,N_334,N_316);
nor U2769 (N_2769,N_392,N_849);
and U2770 (N_2770,N_1159,N_281);
and U2771 (N_2771,N_1063,N_31);
nand U2772 (N_2772,N_419,N_389);
nor U2773 (N_2773,N_514,N_1473);
nor U2774 (N_2774,N_349,N_699);
nor U2775 (N_2775,N_82,N_246);
xor U2776 (N_2776,N_1064,N_181);
xnor U2777 (N_2777,N_397,N_341);
xor U2778 (N_2778,N_797,N_933);
nor U2779 (N_2779,N_1001,N_448);
nor U2780 (N_2780,N_88,N_698);
nand U2781 (N_2781,N_221,N_821);
nor U2782 (N_2782,N_1337,N_667);
nand U2783 (N_2783,N_28,N_82);
nor U2784 (N_2784,N_1498,N_998);
and U2785 (N_2785,N_265,N_1170);
xnor U2786 (N_2786,N_404,N_1187);
nand U2787 (N_2787,N_870,N_941);
nand U2788 (N_2788,N_475,N_368);
or U2789 (N_2789,N_1350,N_1154);
and U2790 (N_2790,N_1056,N_938);
or U2791 (N_2791,N_1038,N_806);
and U2792 (N_2792,N_1244,N_1221);
nand U2793 (N_2793,N_1063,N_505);
or U2794 (N_2794,N_1386,N_892);
or U2795 (N_2795,N_368,N_63);
xnor U2796 (N_2796,N_608,N_322);
or U2797 (N_2797,N_217,N_979);
and U2798 (N_2798,N_894,N_110);
nor U2799 (N_2799,N_312,N_283);
nand U2800 (N_2800,N_1403,N_433);
xor U2801 (N_2801,N_968,N_48);
xor U2802 (N_2802,N_1202,N_1472);
nand U2803 (N_2803,N_868,N_1159);
nand U2804 (N_2804,N_1467,N_1126);
and U2805 (N_2805,N_724,N_492);
and U2806 (N_2806,N_646,N_992);
nor U2807 (N_2807,N_996,N_285);
nor U2808 (N_2808,N_214,N_234);
nor U2809 (N_2809,N_877,N_1037);
and U2810 (N_2810,N_1008,N_1267);
or U2811 (N_2811,N_656,N_434);
and U2812 (N_2812,N_970,N_1035);
or U2813 (N_2813,N_1419,N_308);
xor U2814 (N_2814,N_1046,N_637);
xor U2815 (N_2815,N_709,N_818);
xnor U2816 (N_2816,N_610,N_228);
and U2817 (N_2817,N_363,N_113);
xor U2818 (N_2818,N_244,N_1343);
nor U2819 (N_2819,N_887,N_1320);
nor U2820 (N_2820,N_936,N_1016);
nand U2821 (N_2821,N_395,N_820);
and U2822 (N_2822,N_1124,N_1474);
xor U2823 (N_2823,N_210,N_1307);
nor U2824 (N_2824,N_135,N_1054);
nor U2825 (N_2825,N_244,N_297);
xor U2826 (N_2826,N_1305,N_924);
nor U2827 (N_2827,N_606,N_7);
xnor U2828 (N_2828,N_447,N_934);
nor U2829 (N_2829,N_1266,N_572);
or U2830 (N_2830,N_1395,N_23);
or U2831 (N_2831,N_139,N_1449);
and U2832 (N_2832,N_363,N_1362);
or U2833 (N_2833,N_981,N_123);
and U2834 (N_2834,N_80,N_699);
and U2835 (N_2835,N_360,N_1071);
or U2836 (N_2836,N_383,N_1208);
xor U2837 (N_2837,N_1380,N_507);
and U2838 (N_2838,N_932,N_797);
nor U2839 (N_2839,N_590,N_120);
nor U2840 (N_2840,N_691,N_458);
nand U2841 (N_2841,N_863,N_230);
and U2842 (N_2842,N_932,N_312);
nor U2843 (N_2843,N_480,N_1071);
xnor U2844 (N_2844,N_1437,N_579);
nand U2845 (N_2845,N_827,N_985);
and U2846 (N_2846,N_1337,N_989);
or U2847 (N_2847,N_652,N_896);
nand U2848 (N_2848,N_1440,N_812);
xor U2849 (N_2849,N_1294,N_286);
nand U2850 (N_2850,N_1071,N_125);
xor U2851 (N_2851,N_781,N_519);
xnor U2852 (N_2852,N_948,N_419);
or U2853 (N_2853,N_977,N_1329);
nand U2854 (N_2854,N_626,N_55);
and U2855 (N_2855,N_1320,N_1290);
or U2856 (N_2856,N_1177,N_121);
or U2857 (N_2857,N_583,N_704);
xnor U2858 (N_2858,N_1177,N_325);
nor U2859 (N_2859,N_826,N_429);
and U2860 (N_2860,N_1022,N_330);
or U2861 (N_2861,N_1071,N_603);
xnor U2862 (N_2862,N_352,N_1131);
xnor U2863 (N_2863,N_1381,N_521);
or U2864 (N_2864,N_973,N_809);
nand U2865 (N_2865,N_461,N_903);
nor U2866 (N_2866,N_1056,N_1352);
nand U2867 (N_2867,N_771,N_995);
nor U2868 (N_2868,N_1287,N_351);
xor U2869 (N_2869,N_608,N_347);
nor U2870 (N_2870,N_447,N_418);
nor U2871 (N_2871,N_684,N_1352);
and U2872 (N_2872,N_701,N_678);
xnor U2873 (N_2873,N_1062,N_340);
or U2874 (N_2874,N_515,N_666);
or U2875 (N_2875,N_63,N_411);
and U2876 (N_2876,N_1075,N_853);
nor U2877 (N_2877,N_440,N_1341);
nor U2878 (N_2878,N_1171,N_269);
nand U2879 (N_2879,N_1293,N_134);
xor U2880 (N_2880,N_816,N_603);
or U2881 (N_2881,N_433,N_962);
nand U2882 (N_2882,N_1012,N_219);
and U2883 (N_2883,N_526,N_1083);
and U2884 (N_2884,N_466,N_1271);
nor U2885 (N_2885,N_717,N_662);
xnor U2886 (N_2886,N_703,N_407);
nor U2887 (N_2887,N_774,N_918);
and U2888 (N_2888,N_1437,N_935);
and U2889 (N_2889,N_686,N_167);
nand U2890 (N_2890,N_162,N_15);
or U2891 (N_2891,N_8,N_917);
or U2892 (N_2892,N_229,N_58);
and U2893 (N_2893,N_84,N_1282);
and U2894 (N_2894,N_967,N_1307);
nand U2895 (N_2895,N_1448,N_659);
xnor U2896 (N_2896,N_1095,N_838);
xnor U2897 (N_2897,N_1163,N_1135);
nor U2898 (N_2898,N_1142,N_116);
or U2899 (N_2899,N_369,N_228);
and U2900 (N_2900,N_734,N_746);
or U2901 (N_2901,N_815,N_1284);
nand U2902 (N_2902,N_1445,N_640);
xnor U2903 (N_2903,N_215,N_765);
xnor U2904 (N_2904,N_1390,N_1258);
nand U2905 (N_2905,N_776,N_983);
xnor U2906 (N_2906,N_37,N_1020);
nor U2907 (N_2907,N_1027,N_405);
nor U2908 (N_2908,N_821,N_40);
or U2909 (N_2909,N_205,N_769);
or U2910 (N_2910,N_487,N_1247);
and U2911 (N_2911,N_216,N_387);
nand U2912 (N_2912,N_192,N_1032);
and U2913 (N_2913,N_1127,N_62);
or U2914 (N_2914,N_1365,N_826);
or U2915 (N_2915,N_1468,N_624);
nor U2916 (N_2916,N_574,N_129);
and U2917 (N_2917,N_1208,N_100);
nor U2918 (N_2918,N_1455,N_56);
and U2919 (N_2919,N_92,N_739);
nor U2920 (N_2920,N_1242,N_1305);
xor U2921 (N_2921,N_745,N_993);
xor U2922 (N_2922,N_1426,N_426);
xor U2923 (N_2923,N_1079,N_253);
or U2924 (N_2924,N_859,N_492);
xor U2925 (N_2925,N_851,N_1388);
or U2926 (N_2926,N_264,N_576);
and U2927 (N_2927,N_616,N_840);
or U2928 (N_2928,N_1298,N_925);
nand U2929 (N_2929,N_65,N_1041);
or U2930 (N_2930,N_1210,N_977);
nor U2931 (N_2931,N_256,N_1240);
and U2932 (N_2932,N_338,N_1342);
or U2933 (N_2933,N_923,N_896);
or U2934 (N_2934,N_570,N_1394);
nand U2935 (N_2935,N_85,N_404);
nor U2936 (N_2936,N_979,N_796);
or U2937 (N_2937,N_29,N_391);
nand U2938 (N_2938,N_1436,N_791);
nor U2939 (N_2939,N_292,N_346);
nand U2940 (N_2940,N_1240,N_1354);
or U2941 (N_2941,N_488,N_964);
and U2942 (N_2942,N_525,N_178);
nor U2943 (N_2943,N_974,N_447);
xor U2944 (N_2944,N_271,N_1114);
nor U2945 (N_2945,N_902,N_339);
nand U2946 (N_2946,N_1393,N_702);
and U2947 (N_2947,N_133,N_387);
and U2948 (N_2948,N_1361,N_1409);
nand U2949 (N_2949,N_396,N_257);
or U2950 (N_2950,N_382,N_704);
or U2951 (N_2951,N_83,N_1067);
xnor U2952 (N_2952,N_1266,N_1498);
nand U2953 (N_2953,N_1117,N_1487);
and U2954 (N_2954,N_383,N_1173);
nand U2955 (N_2955,N_1169,N_55);
or U2956 (N_2956,N_586,N_363);
nand U2957 (N_2957,N_81,N_633);
nand U2958 (N_2958,N_1071,N_290);
nand U2959 (N_2959,N_837,N_1203);
or U2960 (N_2960,N_677,N_1438);
nor U2961 (N_2961,N_575,N_595);
nand U2962 (N_2962,N_1419,N_1258);
nand U2963 (N_2963,N_1161,N_155);
or U2964 (N_2964,N_1050,N_993);
nor U2965 (N_2965,N_613,N_1278);
or U2966 (N_2966,N_708,N_637);
or U2967 (N_2967,N_60,N_1450);
nor U2968 (N_2968,N_1041,N_200);
and U2969 (N_2969,N_1498,N_1397);
nor U2970 (N_2970,N_560,N_676);
nand U2971 (N_2971,N_674,N_1096);
and U2972 (N_2972,N_113,N_1484);
xnor U2973 (N_2973,N_27,N_784);
or U2974 (N_2974,N_1094,N_1051);
and U2975 (N_2975,N_1090,N_1363);
or U2976 (N_2976,N_153,N_931);
xnor U2977 (N_2977,N_10,N_837);
or U2978 (N_2978,N_584,N_1480);
nand U2979 (N_2979,N_1027,N_703);
nand U2980 (N_2980,N_988,N_660);
nand U2981 (N_2981,N_1493,N_42);
xor U2982 (N_2982,N_184,N_1427);
and U2983 (N_2983,N_969,N_845);
nor U2984 (N_2984,N_1210,N_566);
nand U2985 (N_2985,N_992,N_277);
xor U2986 (N_2986,N_1323,N_19);
xor U2987 (N_2987,N_13,N_852);
nor U2988 (N_2988,N_686,N_286);
xor U2989 (N_2989,N_110,N_254);
nor U2990 (N_2990,N_872,N_1488);
xnor U2991 (N_2991,N_1108,N_222);
and U2992 (N_2992,N_309,N_1229);
and U2993 (N_2993,N_917,N_47);
nor U2994 (N_2994,N_792,N_1164);
xor U2995 (N_2995,N_1307,N_1148);
xnor U2996 (N_2996,N_50,N_488);
nor U2997 (N_2997,N_1446,N_665);
nand U2998 (N_2998,N_323,N_1093);
and U2999 (N_2999,N_912,N_1311);
and U3000 (N_3000,N_2286,N_2288);
nand U3001 (N_3001,N_1539,N_2574);
nor U3002 (N_3002,N_2987,N_2343);
or U3003 (N_3003,N_1871,N_1838);
and U3004 (N_3004,N_2638,N_1909);
xor U3005 (N_3005,N_1515,N_1517);
nor U3006 (N_3006,N_1701,N_1834);
nand U3007 (N_3007,N_1560,N_2121);
nor U3008 (N_3008,N_1796,N_2631);
nand U3009 (N_3009,N_2065,N_2951);
nand U3010 (N_3010,N_2061,N_1759);
xor U3011 (N_3011,N_1680,N_2986);
xor U3012 (N_3012,N_2613,N_2226);
and U3013 (N_3013,N_1591,N_2349);
xor U3014 (N_3014,N_2992,N_1913);
nand U3015 (N_3015,N_1566,N_2208);
nand U3016 (N_3016,N_1822,N_1824);
nor U3017 (N_3017,N_2344,N_2242);
nand U3018 (N_3018,N_2520,N_1833);
nand U3019 (N_3019,N_2011,N_2253);
nor U3020 (N_3020,N_1638,N_1784);
xor U3021 (N_3021,N_2038,N_2873);
xor U3022 (N_3022,N_2840,N_2458);
and U3023 (N_3023,N_2880,N_1829);
and U3024 (N_3024,N_2018,N_1734);
xor U3025 (N_3025,N_1970,N_1797);
nor U3026 (N_3026,N_2395,N_2280);
and U3027 (N_3027,N_1555,N_2125);
nor U3028 (N_3028,N_2515,N_2417);
nor U3029 (N_3029,N_2846,N_2074);
or U3030 (N_3030,N_2768,N_1595);
nand U3031 (N_3031,N_1685,N_1705);
nand U3032 (N_3032,N_2468,N_2665);
nor U3033 (N_3033,N_1752,N_1804);
or U3034 (N_3034,N_2984,N_2427);
and U3035 (N_3035,N_2776,N_2721);
xor U3036 (N_3036,N_2368,N_1774);
and U3037 (N_3037,N_1636,N_2897);
or U3038 (N_3038,N_1505,N_1847);
or U3039 (N_3039,N_1762,N_2900);
and U3040 (N_3040,N_1621,N_2455);
or U3041 (N_3041,N_2181,N_2975);
and U3042 (N_3042,N_2881,N_2416);
nand U3043 (N_3043,N_2473,N_2157);
and U3044 (N_3044,N_1535,N_2347);
and U3045 (N_3045,N_1894,N_2472);
nand U3046 (N_3046,N_2159,N_2054);
and U3047 (N_3047,N_2488,N_2851);
or U3048 (N_3048,N_1794,N_2722);
xor U3049 (N_3049,N_2719,N_1602);
and U3050 (N_3050,N_2435,N_2034);
nand U3051 (N_3051,N_2747,N_2340);
or U3052 (N_3052,N_2920,N_1520);
nor U3053 (N_3053,N_2329,N_2264);
and U3054 (N_3054,N_2870,N_2444);
or U3055 (N_3055,N_2215,N_1631);
and U3056 (N_3056,N_2799,N_1874);
xor U3057 (N_3057,N_1793,N_2758);
nand U3058 (N_3058,N_1737,N_1519);
or U3059 (N_3059,N_2716,N_2165);
nor U3060 (N_3060,N_2440,N_1528);
nor U3061 (N_3061,N_2677,N_2601);
nand U3062 (N_3062,N_2736,N_2029);
xnor U3063 (N_3063,N_1885,N_1690);
or U3064 (N_3064,N_2112,N_2233);
xnor U3065 (N_3065,N_2672,N_1891);
and U3066 (N_3066,N_1922,N_1882);
nor U3067 (N_3067,N_2718,N_2136);
and U3068 (N_3068,N_1550,N_2192);
nand U3069 (N_3069,N_2466,N_2292);
nand U3070 (N_3070,N_2283,N_1657);
xor U3071 (N_3071,N_2596,N_2558);
nand U3072 (N_3072,N_2265,N_1937);
or U3073 (N_3073,N_1597,N_2807);
xor U3074 (N_3074,N_1574,N_2528);
or U3075 (N_3075,N_2199,N_2757);
or U3076 (N_3076,N_2621,N_2735);
or U3077 (N_3077,N_2274,N_1753);
nor U3078 (N_3078,N_2445,N_2474);
nand U3079 (N_3079,N_2794,N_2801);
nand U3080 (N_3080,N_1647,N_1811);
nand U3081 (N_3081,N_1867,N_1962);
nand U3082 (N_3082,N_1854,N_1691);
xor U3083 (N_3083,N_1604,N_2687);
nand U3084 (N_3084,N_1697,N_2521);
and U3085 (N_3085,N_2235,N_1671);
and U3086 (N_3086,N_2463,N_2365);
xor U3087 (N_3087,N_2971,N_1723);
and U3088 (N_3088,N_2379,N_1892);
nand U3089 (N_3089,N_2839,N_2923);
nor U3090 (N_3090,N_2598,N_1533);
and U3091 (N_3091,N_2066,N_2723);
nor U3092 (N_3092,N_2372,N_2647);
and U3093 (N_3093,N_1659,N_2675);
xor U3094 (N_3094,N_1699,N_2856);
nor U3095 (N_3095,N_2557,N_2308);
xnor U3096 (N_3096,N_1877,N_1567);
xor U3097 (N_3097,N_1789,N_2178);
and U3098 (N_3098,N_2995,N_2590);
or U3099 (N_3099,N_1926,N_2124);
xor U3100 (N_3100,N_2148,N_2693);
or U3101 (N_3101,N_1573,N_2067);
nand U3102 (N_3102,N_2032,N_1989);
or U3103 (N_3103,N_1920,N_2471);
nor U3104 (N_3104,N_1743,N_2163);
and U3105 (N_3105,N_2863,N_2096);
nand U3106 (N_3106,N_2705,N_2015);
and U3107 (N_3107,N_2960,N_1713);
nor U3108 (N_3108,N_2950,N_2707);
nor U3109 (N_3109,N_2778,N_1665);
xnor U3110 (N_3110,N_2775,N_2289);
nand U3111 (N_3111,N_2161,N_2398);
xor U3112 (N_3112,N_2339,N_2037);
nand U3113 (N_3113,N_2115,N_1525);
xnor U3114 (N_3114,N_2016,N_2064);
nor U3115 (N_3115,N_2624,N_2983);
nor U3116 (N_3116,N_2099,N_2554);
or U3117 (N_3117,N_2392,N_2536);
nor U3118 (N_3118,N_2771,N_2421);
or U3119 (N_3119,N_1662,N_1510);
and U3120 (N_3120,N_2966,N_2750);
or U3121 (N_3121,N_2766,N_2056);
nand U3122 (N_3122,N_2953,N_2872);
nor U3123 (N_3123,N_2699,N_1725);
nand U3124 (N_3124,N_2063,N_2105);
xor U3125 (N_3125,N_1571,N_2060);
or U3126 (N_3126,N_2793,N_1582);
xnor U3127 (N_3127,N_2350,N_1850);
nand U3128 (N_3128,N_2439,N_2833);
or U3129 (N_3129,N_2332,N_2564);
nand U3130 (N_3130,N_2715,N_2791);
nor U3131 (N_3131,N_2173,N_1942);
nand U3132 (N_3132,N_2563,N_2709);
nand U3133 (N_3133,N_2451,N_2322);
nor U3134 (N_3134,N_1722,N_2498);
nand U3135 (N_3135,N_2464,N_1741);
nor U3136 (N_3136,N_1546,N_2397);
and U3137 (N_3137,N_2262,N_1982);
xnor U3138 (N_3138,N_2185,N_2772);
xnor U3139 (N_3139,N_1872,N_2737);
and U3140 (N_3140,N_1908,N_2626);
and U3141 (N_3141,N_2519,N_1682);
nor U3142 (N_3142,N_2408,N_2649);
nand U3143 (N_3143,N_1817,N_2634);
and U3144 (N_3144,N_2109,N_2117);
nand U3145 (N_3145,N_2313,N_1740);
and U3146 (N_3146,N_2179,N_2333);
or U3147 (N_3147,N_2635,N_2568);
and U3148 (N_3148,N_2341,N_2250);
or U3149 (N_3149,N_2195,N_1953);
xnor U3150 (N_3150,N_2906,N_2273);
nor U3151 (N_3151,N_1827,N_2695);
nand U3152 (N_3152,N_1767,N_2380);
xor U3153 (N_3153,N_2603,N_2725);
nand U3154 (N_3154,N_2957,N_2166);
nand U3155 (N_3155,N_2353,N_2689);
xor U3156 (N_3156,N_1612,N_2499);
or U3157 (N_3157,N_2360,N_2314);
nor U3158 (N_3158,N_2114,N_2524);
xor U3159 (N_3159,N_1904,N_2324);
or U3160 (N_3160,N_2909,N_2712);
nor U3161 (N_3161,N_1868,N_2935);
or U3162 (N_3162,N_1792,N_1551);
and U3163 (N_3163,N_2714,N_2615);
nand U3164 (N_3164,N_2207,N_1915);
xnor U3165 (N_3165,N_2809,N_1786);
xnor U3166 (N_3166,N_2400,N_2913);
or U3167 (N_3167,N_1531,N_2546);
or U3168 (N_3168,N_1836,N_2550);
xor U3169 (N_3169,N_2278,N_2948);
and U3170 (N_3170,N_1598,N_1512);
xor U3171 (N_3171,N_2113,N_2257);
nand U3172 (N_3172,N_2120,N_2751);
xnor U3173 (N_3173,N_2077,N_1552);
or U3174 (N_3174,N_1732,N_1559);
and U3175 (N_3175,N_2146,N_2510);
nand U3176 (N_3176,N_2625,N_2566);
nor U3177 (N_3177,N_2850,N_2299);
or U3178 (N_3178,N_2248,N_2095);
nand U3179 (N_3179,N_2661,N_2017);
and U3180 (N_3180,N_1637,N_2245);
nand U3181 (N_3181,N_2864,N_1799);
nor U3182 (N_3182,N_2090,N_2260);
nor U3183 (N_3183,N_1808,N_1813);
nand U3184 (N_3184,N_2469,N_2927);
xnor U3185 (N_3185,N_2462,N_2849);
xnor U3186 (N_3186,N_2352,N_2069);
xnor U3187 (N_3187,N_2430,N_2197);
or U3188 (N_3188,N_2938,N_2149);
nor U3189 (N_3189,N_2973,N_2565);
nand U3190 (N_3190,N_2128,N_2654);
or U3191 (N_3191,N_2831,N_2399);
xor U3192 (N_3192,N_2362,N_2355);
nand U3193 (N_3193,N_1695,N_2052);
xor U3194 (N_3194,N_2160,N_2046);
nand U3195 (N_3195,N_2697,N_1603);
xnor U3196 (N_3196,N_2860,N_2652);
xnor U3197 (N_3197,N_2307,N_2828);
xnor U3198 (N_3198,N_1627,N_2806);
and U3199 (N_3199,N_2680,N_2073);
xnor U3200 (N_3200,N_2522,N_2126);
nand U3201 (N_3201,N_1565,N_1619);
nand U3202 (N_3202,N_2559,N_2925);
nand U3203 (N_3203,N_2177,N_2055);
xnor U3204 (N_3204,N_2230,N_2543);
nor U3205 (N_3205,N_1846,N_1773);
nand U3206 (N_3206,N_2949,N_2965);
nor U3207 (N_3207,N_1738,N_1624);
xnor U3208 (N_3208,N_2594,N_1679);
xor U3209 (N_3209,N_1516,N_1879);
nor U3210 (N_3210,N_2062,N_1523);
nand U3211 (N_3211,N_2782,N_2338);
nor U3212 (N_3212,N_1764,N_2614);
or U3213 (N_3213,N_2852,N_2815);
and U3214 (N_3214,N_2764,N_2492);
xnor U3215 (N_3215,N_1934,N_1806);
and U3216 (N_3216,N_1835,N_1664);
nor U3217 (N_3217,N_1852,N_2847);
or U3218 (N_3218,N_1825,N_2495);
xnor U3219 (N_3219,N_2405,N_2502);
nand U3220 (N_3220,N_2182,N_1965);
nand U3221 (N_3221,N_2836,N_2443);
nand U3222 (N_3222,N_1957,N_1581);
nand U3223 (N_3223,N_1666,N_1749);
or U3224 (N_3224,N_2460,N_1949);
and U3225 (N_3225,N_2051,N_2744);
or U3226 (N_3226,N_1991,N_2779);
and U3227 (N_3227,N_2490,N_1675);
or U3228 (N_3228,N_2020,N_1748);
and U3229 (N_3229,N_2952,N_2083);
xnor U3230 (N_3230,N_1720,N_1858);
or U3231 (N_3231,N_2438,N_2739);
and U3232 (N_3232,N_2104,N_2033);
nand U3233 (N_3233,N_1634,N_2317);
and U3234 (N_3234,N_2172,N_2947);
xor U3235 (N_3235,N_1742,N_2921);
xor U3236 (N_3236,N_1673,N_1576);
nand U3237 (N_3237,N_1707,N_2845);
nand U3238 (N_3238,N_1542,N_2236);
nand U3239 (N_3239,N_2529,N_1540);
or U3240 (N_3240,N_1947,N_1783);
nand U3241 (N_3241,N_1974,N_1577);
and U3242 (N_3242,N_2788,N_2537);
xor U3243 (N_3243,N_2143,N_2036);
nand U3244 (N_3244,N_2803,N_2385);
and U3245 (N_3245,N_2817,N_2989);
nand U3246 (N_3246,N_2222,N_2388);
and U3247 (N_3247,N_1980,N_2648);
nand U3248 (N_3248,N_1564,N_1584);
nand U3249 (N_3249,N_2005,N_1655);
xnor U3250 (N_3250,N_2223,N_2664);
and U3251 (N_3251,N_2021,N_1545);
xnor U3252 (N_3252,N_1785,N_2483);
or U3253 (N_3253,N_1534,N_2883);
and U3254 (N_3254,N_2437,N_2926);
xor U3255 (N_3255,N_1860,N_1820);
and U3256 (N_3256,N_2482,N_2760);
and U3257 (N_3257,N_1781,N_1927);
and U3258 (N_3258,N_1661,N_1912);
nand U3259 (N_3259,N_1766,N_1663);
or U3260 (N_3260,N_2560,N_2040);
or U3261 (N_3261,N_1717,N_2454);
and U3262 (N_3262,N_1791,N_2549);
and U3263 (N_3263,N_2946,N_1541);
xnor U3264 (N_3264,N_2701,N_1605);
nand U3265 (N_3265,N_2196,N_1861);
nor U3266 (N_3266,N_1587,N_1807);
or U3267 (N_3267,N_1945,N_2198);
nor U3268 (N_3268,N_2170,N_1809);
nor U3269 (N_3269,N_1626,N_1538);
and U3270 (N_3270,N_2898,N_1964);
or U3271 (N_3271,N_2206,N_2001);
or U3272 (N_3272,N_1630,N_2251);
nor U3273 (N_3273,N_2147,N_1727);
xor U3274 (N_3274,N_1544,N_2452);
and U3275 (N_3275,N_1700,N_2918);
and U3276 (N_3276,N_2369,N_1869);
and U3277 (N_3277,N_2076,N_1961);
and U3278 (N_3278,N_2786,N_2821);
nand U3279 (N_3279,N_2829,N_1589);
nand U3280 (N_3280,N_2057,N_1692);
xor U3281 (N_3281,N_2091,N_2331);
nand U3282 (N_3282,N_2048,N_1898);
and U3283 (N_3283,N_2457,N_2140);
nor U3284 (N_3284,N_1779,N_2282);
nor U3285 (N_3285,N_2303,N_1536);
or U3286 (N_3286,N_2994,N_2361);
xor U3287 (N_3287,N_2434,N_1529);
and U3288 (N_3288,N_2660,N_2577);
xor U3289 (N_3289,N_2587,N_2345);
nand U3290 (N_3290,N_2657,N_2406);
nand U3291 (N_3291,N_2270,N_2356);
xnor U3292 (N_3292,N_1645,N_2008);
or U3293 (N_3293,N_2323,N_1609);
or U3294 (N_3294,N_2859,N_2296);
nor U3295 (N_3295,N_1939,N_1802);
nor U3296 (N_3296,N_2127,N_2942);
and U3297 (N_3297,N_1746,N_2259);
and U3298 (N_3298,N_1640,N_1831);
nand U3299 (N_3299,N_2628,N_2465);
and U3300 (N_3300,N_1928,N_2700);
nor U3301 (N_3301,N_2097,N_2415);
xor U3302 (N_3302,N_2589,N_2713);
and U3303 (N_3303,N_2820,N_2876);
nand U3304 (N_3304,N_2111,N_2669);
nand U3305 (N_3305,N_1726,N_1855);
or U3306 (N_3306,N_2326,N_1986);
nor U3307 (N_3307,N_2619,N_2058);
nor U3308 (N_3308,N_2205,N_2901);
or U3309 (N_3309,N_2028,N_2093);
nand U3310 (N_3310,N_2049,N_2261);
xnor U3311 (N_3311,N_1736,N_2171);
xnor U3312 (N_3312,N_2006,N_1954);
or U3313 (N_3313,N_1890,N_2085);
or U3314 (N_3314,N_1704,N_2375);
and U3315 (N_3315,N_1681,N_2731);
and U3316 (N_3316,N_2742,N_1710);
or U3317 (N_3317,N_2977,N_2879);
nor U3318 (N_3318,N_2783,N_2970);
xor U3319 (N_3319,N_2425,N_2168);
nand U3320 (N_3320,N_1652,N_2878);
xnor U3321 (N_3321,N_1966,N_2228);
or U3322 (N_3322,N_2402,N_2396);
nand U3323 (N_3323,N_1893,N_2305);
nand U3324 (N_3324,N_1578,N_1952);
nor U3325 (N_3325,N_1651,N_1895);
nand U3326 (N_3326,N_2633,N_2275);
nand U3327 (N_3327,N_2348,N_2390);
xnor U3328 (N_3328,N_1521,N_1669);
and U3329 (N_3329,N_2094,N_2886);
and U3330 (N_3330,N_2476,N_2240);
nor U3331 (N_3331,N_2050,N_1696);
xor U3332 (N_3332,N_2187,N_1865);
nand U3333 (N_3333,N_1899,N_2190);
nor U3334 (N_3334,N_2936,N_2941);
xnor U3335 (N_3335,N_1985,N_2180);
and U3336 (N_3336,N_1628,N_1735);
nand U3337 (N_3337,N_2717,N_2745);
or U3338 (N_3338,N_2496,N_2584);
and U3339 (N_3339,N_2756,N_2996);
and U3340 (N_3340,N_2982,N_2221);
xnor U3341 (N_3341,N_2387,N_2068);
and U3342 (N_3342,N_2391,N_2910);
xor U3343 (N_3343,N_2284,N_2746);
and U3344 (N_3344,N_1658,N_2724);
or U3345 (N_3345,N_1563,N_2310);
nand U3346 (N_3346,N_2894,N_1990);
or U3347 (N_3347,N_1729,N_2004);
nand U3348 (N_3348,N_2639,N_2151);
xor U3349 (N_3349,N_2072,N_1756);
or U3350 (N_3350,N_2991,N_2610);
and U3351 (N_3351,N_2403,N_2517);
nand U3352 (N_3352,N_2059,N_2928);
nand U3353 (N_3353,N_2446,N_2548);
nor U3354 (N_3354,N_2583,N_2497);
nand U3355 (N_3355,N_2301,N_2186);
nor U3356 (N_3356,N_2100,N_1754);
xnor U3357 (N_3357,N_2258,N_1818);
or U3358 (N_3358,N_2123,N_2656);
xor U3359 (N_3359,N_2729,N_2754);
nand U3360 (N_3360,N_2899,N_2959);
nor U3361 (N_3361,N_2137,N_1946);
or U3362 (N_3362,N_2777,N_2486);
or U3363 (N_3363,N_2480,N_2075);
or U3364 (N_3364,N_1731,N_2084);
nand U3365 (N_3365,N_2203,N_2263);
xnor U3366 (N_3366,N_2842,N_1914);
or U3367 (N_3367,N_1625,N_2304);
or U3368 (N_3368,N_1608,N_2688);
xor U3369 (N_3369,N_2896,N_1821);
or U3370 (N_3370,N_2968,N_1708);
and U3371 (N_3371,N_1851,N_2903);
or U3372 (N_3372,N_2893,N_2922);
nor U3373 (N_3373,N_2916,N_2044);
or U3374 (N_3374,N_2802,N_2254);
or U3375 (N_3375,N_2007,N_1586);
nor U3376 (N_3376,N_2366,N_1593);
nand U3377 (N_3377,N_2306,N_1557);
and U3378 (N_3378,N_2422,N_2667);
or U3379 (N_3379,N_2853,N_2103);
xor U3380 (N_3380,N_2357,N_2641);
xor U3381 (N_3381,N_2377,N_2266);
and U3382 (N_3382,N_2189,N_1642);
xor U3383 (N_3383,N_2291,N_2122);
nand U3384 (N_3384,N_2431,N_2969);
xnor U3385 (N_3385,N_2389,N_2204);
xnor U3386 (N_3386,N_2071,N_2370);
nand U3387 (N_3387,N_2684,N_2911);
xor U3388 (N_3388,N_2981,N_2875);
or U3389 (N_3389,N_2553,N_1782);
xnor U3390 (N_3390,N_2690,N_2214);
or U3391 (N_3391,N_1606,N_1839);
xor U3392 (N_3392,N_2551,N_2386);
or U3393 (N_3393,N_2080,N_2133);
and U3394 (N_3394,N_1744,N_2600);
nor U3395 (N_3395,N_2604,N_2830);
or U3396 (N_3396,N_1880,N_1810);
or U3397 (N_3397,N_2843,N_2710);
and U3398 (N_3398,N_2732,N_2047);
nand U3399 (N_3399,N_1768,N_2796);
xnor U3400 (N_3400,N_2447,N_2150);
nand U3401 (N_3401,N_2512,N_2741);
nand U3402 (N_3402,N_2383,N_2481);
nand U3403 (N_3403,N_2426,N_2999);
or U3404 (N_3404,N_2030,N_2651);
and U3405 (N_3405,N_2210,N_2116);
xor U3406 (N_3406,N_1568,N_2868);
xor U3407 (N_3407,N_2686,N_2570);
nor U3408 (N_3408,N_1677,N_2153);
and U3409 (N_3409,N_2798,N_2988);
and U3410 (N_3410,N_1569,N_2108);
nor U3411 (N_3411,N_2276,N_2767);
nand U3412 (N_3412,N_1883,N_1607);
xor U3413 (N_3413,N_1644,N_2882);
or U3414 (N_3414,N_1844,N_2407);
nand U3415 (N_3415,N_2837,N_2797);
nor U3416 (N_3416,N_2670,N_2573);
nor U3417 (N_3417,N_2234,N_2618);
xor U3418 (N_3418,N_1522,N_2169);
xnor U3419 (N_3419,N_2671,N_2364);
nand U3420 (N_3420,N_1967,N_1513);
or U3421 (N_3421,N_2698,N_2382);
nor U3422 (N_3422,N_2571,N_1943);
nor U3423 (N_3423,N_2183,N_2131);
xnor U3424 (N_3424,N_1988,N_1968);
xor U3425 (N_3425,N_2142,N_2748);
nor U3426 (N_3426,N_2752,N_2956);
and U3427 (N_3427,N_2325,N_1888);
nand U3428 (N_3428,N_2679,N_2449);
xor U3429 (N_3429,N_2523,N_1973);
nor U3430 (N_3430,N_2293,N_1814);
and U3431 (N_3431,N_2247,N_2394);
and U3432 (N_3432,N_2937,N_2620);
nor U3433 (N_3433,N_1905,N_2964);
nand U3434 (N_3434,N_2201,N_2410);
or U3435 (N_3435,N_1896,N_2184);
nand U3436 (N_3436,N_1635,N_1862);
nand U3437 (N_3437,N_2592,N_2374);
xnor U3438 (N_3438,N_2477,N_2567);
nand U3439 (N_3439,N_2188,N_2838);
nor U3440 (N_3440,N_2042,N_2428);
nor U3441 (N_3441,N_1875,N_2354);
nand U3442 (N_3442,N_2209,N_1757);
or U3443 (N_3443,N_2252,N_2659);
and U3444 (N_3444,N_2743,N_2041);
nand U3445 (N_3445,N_2692,N_1798);
nand U3446 (N_3446,N_2167,N_1676);
or U3447 (N_3447,N_2514,N_1509);
or U3448 (N_3448,N_1715,N_2287);
nand U3449 (N_3449,N_2704,N_2225);
xor U3450 (N_3450,N_1910,N_2871);
and U3451 (N_3451,N_1936,N_2429);
nand U3452 (N_3452,N_2281,N_2993);
xnor U3453 (N_3453,N_2586,N_2552);
nand U3454 (N_3454,N_2022,N_2191);
nor U3455 (N_3455,N_1611,N_2855);
or U3456 (N_3456,N_2433,N_2810);
and U3457 (N_3457,N_1837,N_1866);
nor U3458 (N_3458,N_2834,N_2891);
or U3459 (N_3459,N_1780,N_2424);
and U3460 (N_3460,N_1929,N_2629);
xnor U3461 (N_3461,N_2678,N_2569);
or U3462 (N_3462,N_2367,N_2795);
nand U3463 (N_3463,N_1765,N_2556);
or U3464 (N_3464,N_2762,N_2655);
nor U3465 (N_3465,N_1958,N_2513);
and U3466 (N_3466,N_2441,N_2479);
xor U3467 (N_3467,N_1975,N_2814);
or U3468 (N_3468,N_2418,N_2599);
and U3469 (N_3469,N_2271,N_2193);
and U3470 (N_3470,N_2101,N_2759);
and U3471 (N_3471,N_2774,N_2243);
nand U3472 (N_3472,N_1527,N_2256);
and U3473 (N_3473,N_1594,N_2781);
nand U3474 (N_3474,N_2884,N_2623);
nor U3475 (N_3475,N_1900,N_2773);
nand U3476 (N_3476,N_1590,N_2534);
nor U3477 (N_3477,N_2026,N_2591);
or U3478 (N_3478,N_2087,N_2082);
or U3479 (N_3479,N_2812,N_1500);
or U3480 (N_3480,N_2811,N_2607);
and U3481 (N_3481,N_2738,N_2373);
or U3482 (N_3482,N_2749,N_2681);
and U3483 (N_3483,N_2914,N_1983);
and U3484 (N_3484,N_2475,N_2535);
xor U3485 (N_3485,N_2107,N_1841);
nand U3486 (N_3486,N_1709,N_2943);
xnor U3487 (N_3487,N_2213,N_2990);
and U3488 (N_3488,N_1526,N_2616);
nand U3489 (N_3489,N_1935,N_1897);
nand U3490 (N_3490,N_2593,N_1583);
nand U3491 (N_3491,N_1650,N_1508);
or U3492 (N_3492,N_2024,N_2867);
nor U3493 (N_3493,N_2890,N_2784);
and U3494 (N_3494,N_2432,N_2932);
nand U3495 (N_3495,N_2493,N_1884);
and U3496 (N_3496,N_1554,N_1728);
xnor U3497 (N_3497,N_2409,N_1790);
nand U3498 (N_3498,N_1951,N_1689);
xor U3499 (N_3499,N_2892,N_1623);
nor U3500 (N_3500,N_2816,N_2805);
nor U3501 (N_3501,N_2019,N_2164);
xor U3502 (N_3502,N_2371,N_2027);
or U3503 (N_3503,N_2078,N_2539);
nand U3504 (N_3504,N_2542,N_2877);
xor U3505 (N_3505,N_1805,N_2572);
or U3506 (N_3506,N_1955,N_2889);
nand U3507 (N_3507,N_2682,N_2378);
nand U3508 (N_3508,N_2470,N_1863);
nor U3509 (N_3509,N_2232,N_2268);
and U3510 (N_3510,N_2818,N_1711);
xor U3511 (N_3511,N_2813,N_2787);
and U3512 (N_3512,N_2010,N_2929);
nand U3513 (N_3513,N_2154,N_2980);
and U3514 (N_3514,N_1653,N_2848);
xor U3515 (N_3515,N_2485,N_2316);
and U3516 (N_3516,N_2895,N_2294);
xor U3517 (N_3517,N_1714,N_2606);
nand U3518 (N_3518,N_1543,N_1667);
nor U3519 (N_3519,N_1755,N_2319);
and U3520 (N_3520,N_2401,N_2792);
and U3521 (N_3521,N_2162,N_2645);
xor U3522 (N_3522,N_1549,N_2770);
nand U3523 (N_3523,N_2597,N_2511);
nand U3524 (N_3524,N_2862,N_1801);
and U3525 (N_3525,N_1668,N_1823);
nand U3526 (N_3526,N_1530,N_2376);
nand U3527 (N_3527,N_2217,N_1599);
and U3528 (N_3528,N_1776,N_2555);
xor U3529 (N_3529,N_2320,N_1812);
xnor U3530 (N_3530,N_1948,N_2155);
nand U3531 (N_3531,N_1614,N_1601);
nor U3532 (N_3532,N_1916,N_2249);
or U3533 (N_3533,N_1629,N_1660);
and U3534 (N_3534,N_1887,N_1941);
nor U3535 (N_3535,N_2582,N_2985);
and U3536 (N_3536,N_1562,N_2312);
xor U3537 (N_3537,N_2538,N_2919);
xor U3538 (N_3538,N_2931,N_2532);
nor U3539 (N_3539,N_1683,N_2130);
or U3540 (N_3540,N_2547,N_1706);
xor U3541 (N_3541,N_2753,N_2540);
nor U3542 (N_3542,N_2504,N_2979);
or U3543 (N_3543,N_2808,N_1750);
xor U3544 (N_3544,N_2734,N_2035);
nor U3545 (N_3545,N_2218,N_2579);
or U3546 (N_3546,N_2720,N_2448);
nor U3547 (N_3547,N_2450,N_2643);
xor U3548 (N_3548,N_2861,N_2506);
nand U3549 (N_3549,N_1921,N_2384);
or U3550 (N_3550,N_2826,N_2346);
nand U3551 (N_3551,N_2658,N_1703);
nand U3552 (N_3552,N_1993,N_2436);
nor U3553 (N_3553,N_2733,N_2581);
nand U3554 (N_3554,N_1588,N_2974);
or U3555 (N_3555,N_2944,N_2915);
and U3556 (N_3556,N_1976,N_1940);
nand U3557 (N_3557,N_1881,N_1843);
or U3558 (N_3558,N_1787,N_1532);
nor U3559 (N_3559,N_2650,N_2662);
xnor U3560 (N_3560,N_2216,N_2501);
xor U3561 (N_3561,N_2958,N_1643);
or U3562 (N_3562,N_2381,N_1761);
or U3563 (N_3563,N_1994,N_1501);
or U3564 (N_3564,N_2602,N_2857);
xnor U3565 (N_3565,N_2726,N_2088);
nand U3566 (N_3566,N_2824,N_2622);
nand U3567 (N_3567,N_2089,N_2461);
or U3568 (N_3568,N_2727,N_2706);
or U3569 (N_3569,N_2685,N_1730);
nand U3570 (N_3570,N_1672,N_2315);
and U3571 (N_3571,N_2518,N_1977);
or U3572 (N_3572,N_2819,N_2031);
nand U3573 (N_3573,N_2342,N_2012);
nand U3574 (N_3574,N_1719,N_2269);
xor U3575 (N_3575,N_1944,N_1575);
nand U3576 (N_3576,N_1911,N_2487);
xnor U3577 (N_3577,N_2822,N_2902);
or U3578 (N_3578,N_1777,N_2646);
or U3579 (N_3579,N_1999,N_2702);
or U3580 (N_3580,N_1633,N_1641);
and U3581 (N_3581,N_2972,N_1687);
xor U3582 (N_3582,N_1613,N_1938);
xor U3583 (N_3583,N_1997,N_2013);
and U3584 (N_3584,N_2825,N_1572);
nor U3585 (N_3585,N_2298,N_2930);
nand U3586 (N_3586,N_1721,N_2290);
xor U3587 (N_3587,N_2420,N_2255);
nand U3588 (N_3588,N_1903,N_2780);
xnor U3589 (N_3589,N_1716,N_1684);
xor U3590 (N_3590,N_2351,N_2227);
nor U3591 (N_3591,N_2575,N_2841);
or U3592 (N_3592,N_1960,N_1972);
nor U3593 (N_3593,N_2321,N_2079);
nand U3594 (N_3594,N_1901,N_2674);
and U3595 (N_3595,N_2098,N_2414);
nor U3596 (N_3596,N_1840,N_2605);
xnor U3597 (N_3597,N_2630,N_1561);
or U3598 (N_3598,N_2176,N_2358);
nor U3599 (N_3599,N_2874,N_2404);
and U3600 (N_3600,N_2827,N_1670);
or U3601 (N_3601,N_2561,N_2632);
or U3602 (N_3602,N_2644,N_1886);
or U3603 (N_3603,N_2666,N_1502);
or U3604 (N_3604,N_1503,N_2769);
nand U3605 (N_3605,N_1859,N_2311);
nor U3606 (N_3606,N_2835,N_2334);
nor U3607 (N_3607,N_2609,N_2761);
xnor U3608 (N_3608,N_2102,N_1616);
xnor U3609 (N_3609,N_2231,N_2933);
nor U3610 (N_3610,N_1688,N_1933);
nor U3611 (N_3611,N_1694,N_2070);
and U3612 (N_3612,N_1763,N_2728);
or U3613 (N_3613,N_2145,N_2961);
nand U3614 (N_3614,N_2703,N_1819);
and U3615 (N_3615,N_1579,N_2300);
nor U3616 (N_3616,N_2238,N_2636);
and U3617 (N_3617,N_2765,N_2541);
nor U3618 (N_3618,N_1950,N_1558);
or U3619 (N_3619,N_1504,N_1876);
nand U3620 (N_3620,N_1845,N_1506);
and U3621 (N_3621,N_1646,N_2494);
and U3622 (N_3622,N_2045,N_2611);
nand U3623 (N_3623,N_1615,N_2144);
or U3624 (N_3624,N_2359,N_2442);
or U3625 (N_3625,N_2081,N_1923);
nor U3626 (N_3626,N_2789,N_1733);
xnor U3627 (N_3627,N_1596,N_2413);
nor U3628 (N_3628,N_2092,N_2309);
nand U3629 (N_3629,N_2174,N_2336);
nand U3630 (N_3630,N_2211,N_2976);
nand U3631 (N_3631,N_2907,N_2328);
nand U3632 (N_3632,N_1995,N_2014);
xnor U3633 (N_3633,N_2239,N_2800);
nor U3634 (N_3634,N_1979,N_2673);
nor U3635 (N_3635,N_2578,N_1889);
xnor U3636 (N_3636,N_2866,N_2318);
nand U3637 (N_3637,N_2940,N_2967);
and U3638 (N_3638,N_2954,N_2132);
or U3639 (N_3639,N_1771,N_1984);
nor U3640 (N_3640,N_2585,N_1832);
xnor U3641 (N_3641,N_1878,N_2003);
nor U3642 (N_3642,N_1770,N_1853);
nor U3643 (N_3643,N_2790,N_2194);
nor U3644 (N_3644,N_2484,N_1553);
and U3645 (N_3645,N_2668,N_1992);
nor U3646 (N_3646,N_2478,N_2832);
and U3647 (N_3647,N_2694,N_1981);
nand U3648 (N_3648,N_1873,N_2545);
nor U3649 (N_3649,N_2998,N_2412);
and U3650 (N_3650,N_1849,N_2110);
nor U3651 (N_3651,N_1760,N_1775);
nor U3652 (N_3652,N_1925,N_2588);
and U3653 (N_3653,N_2489,N_1998);
nand U3654 (N_3654,N_1803,N_1856);
and U3655 (N_3655,N_1639,N_2526);
xnor U3656 (N_3656,N_1963,N_2904);
and U3657 (N_3657,N_1864,N_2330);
or U3658 (N_3658,N_2640,N_2934);
nand U3659 (N_3659,N_1919,N_2676);
and U3660 (N_3660,N_1674,N_1622);
or U3661 (N_3661,N_1918,N_2459);
and U3662 (N_3662,N_2978,N_1971);
nand U3663 (N_3663,N_1769,N_1870);
xnor U3664 (N_3664,N_2139,N_2453);
xor U3665 (N_3665,N_1996,N_2267);
xnor U3666 (N_3666,N_1959,N_1751);
or U3667 (N_3667,N_2509,N_2224);
or U3668 (N_3668,N_1698,N_2002);
and U3669 (N_3669,N_1632,N_2887);
or U3670 (N_3670,N_2612,N_2241);
and U3671 (N_3671,N_2000,N_1932);
nand U3672 (N_3672,N_2823,N_1678);
nand U3673 (N_3673,N_2327,N_2804);
nand U3674 (N_3674,N_2627,N_2279);
and U3675 (N_3675,N_2617,N_2295);
nand U3676 (N_3676,N_1648,N_2888);
and U3677 (N_3677,N_2491,N_2663);
xnor U3678 (N_3678,N_2152,N_2963);
xor U3679 (N_3679,N_2562,N_1828);
nor U3680 (N_3680,N_1548,N_2363);
nor U3681 (N_3681,N_2158,N_1848);
xnor U3682 (N_3682,N_1610,N_1524);
xnor U3683 (N_3683,N_1816,N_2229);
nor U3684 (N_3684,N_1969,N_2219);
nand U3685 (N_3685,N_2691,N_2908);
or U3686 (N_3686,N_2302,N_2393);
and U3687 (N_3687,N_1956,N_2955);
or U3688 (N_3688,N_1778,N_2844);
or U3689 (N_3689,N_1842,N_1758);
and U3690 (N_3690,N_2653,N_1772);
nand U3691 (N_3691,N_2530,N_2507);
or U3692 (N_3692,N_2912,N_2595);
xor U3693 (N_3693,N_2730,N_2869);
or U3694 (N_3694,N_2156,N_2106);
nand U3695 (N_3695,N_1815,N_1917);
nor U3696 (N_3696,N_1930,N_1570);
xor U3697 (N_3697,N_2945,N_2212);
or U3698 (N_3698,N_1739,N_1547);
or U3699 (N_3699,N_2335,N_1747);
nor U3700 (N_3700,N_2917,N_1585);
nand U3701 (N_3701,N_2467,N_2763);
nor U3702 (N_3702,N_2858,N_1649);
nor U3703 (N_3703,N_1537,N_2500);
and U3704 (N_3704,N_2865,N_2516);
nand U3705 (N_3705,N_2580,N_2411);
or U3706 (N_3706,N_1702,N_2138);
nand U3707 (N_3707,N_2200,N_1857);
nor U3708 (N_3708,N_2053,N_2272);
nor U3709 (N_3709,N_2285,N_2297);
xor U3710 (N_3710,N_2419,N_1788);
xor U3711 (N_3711,N_1907,N_1693);
or U3712 (N_3712,N_2905,N_1712);
or U3713 (N_3713,N_1511,N_2708);
and U3714 (N_3714,N_1826,N_2637);
or U3715 (N_3715,N_2755,N_1592);
nor U3716 (N_3716,N_1978,N_1507);
xor U3717 (N_3717,N_2962,N_2039);
nor U3718 (N_3718,N_2503,N_1718);
nor U3719 (N_3719,N_1906,N_1987);
nor U3720 (N_3720,N_1795,N_1580);
or U3721 (N_3721,N_2141,N_2525);
or U3722 (N_3722,N_1745,N_2505);
xnor U3723 (N_3723,N_2527,N_1654);
and U3724 (N_3724,N_1656,N_1800);
or U3725 (N_3725,N_2456,N_1518);
nand U3726 (N_3726,N_2043,N_2544);
and U3727 (N_3727,N_1902,N_2997);
and U3728 (N_3728,N_1931,N_2220);
or U3729 (N_3729,N_2118,N_2696);
or U3730 (N_3730,N_2009,N_2129);
and U3731 (N_3731,N_1600,N_2608);
and U3732 (N_3732,N_2337,N_1686);
and U3733 (N_3733,N_2134,N_2785);
nand U3734 (N_3734,N_2576,N_2885);
or U3735 (N_3735,N_1556,N_2711);
or U3736 (N_3736,N_2740,N_1830);
and U3737 (N_3737,N_2023,N_2533);
nor U3738 (N_3738,N_2237,N_1617);
and U3739 (N_3739,N_2531,N_2119);
or U3740 (N_3740,N_2202,N_2086);
nand U3741 (N_3741,N_2508,N_2683);
xnor U3742 (N_3742,N_2423,N_1620);
or U3743 (N_3743,N_1724,N_1618);
nor U3744 (N_3744,N_2246,N_2135);
xnor U3745 (N_3745,N_2854,N_1924);
nor U3746 (N_3746,N_1514,N_2939);
nand U3747 (N_3747,N_2924,N_2175);
nand U3748 (N_3748,N_2244,N_2025);
and U3749 (N_3749,N_2277,N_2642);
nand U3750 (N_3750,N_1788,N_2992);
nand U3751 (N_3751,N_2229,N_1520);
xnor U3752 (N_3752,N_2534,N_1952);
nor U3753 (N_3753,N_1739,N_2778);
xor U3754 (N_3754,N_1812,N_2245);
nor U3755 (N_3755,N_1998,N_1829);
nor U3756 (N_3756,N_1526,N_2687);
nor U3757 (N_3757,N_2182,N_1548);
or U3758 (N_3758,N_1914,N_1762);
and U3759 (N_3759,N_2115,N_1690);
nand U3760 (N_3760,N_1733,N_1515);
nor U3761 (N_3761,N_2695,N_2915);
xnor U3762 (N_3762,N_1855,N_2183);
nand U3763 (N_3763,N_2251,N_1800);
and U3764 (N_3764,N_1825,N_2093);
or U3765 (N_3765,N_2296,N_2984);
nand U3766 (N_3766,N_2673,N_1967);
and U3767 (N_3767,N_2203,N_2221);
nand U3768 (N_3768,N_2408,N_2966);
xor U3769 (N_3769,N_2129,N_2791);
or U3770 (N_3770,N_1798,N_2908);
xnor U3771 (N_3771,N_2530,N_1821);
or U3772 (N_3772,N_2738,N_1734);
nor U3773 (N_3773,N_2815,N_2509);
and U3774 (N_3774,N_2216,N_1967);
xnor U3775 (N_3775,N_2433,N_1689);
xnor U3776 (N_3776,N_2048,N_2956);
xor U3777 (N_3777,N_2545,N_1843);
nand U3778 (N_3778,N_2427,N_2033);
and U3779 (N_3779,N_2803,N_2626);
and U3780 (N_3780,N_2067,N_2309);
nand U3781 (N_3781,N_2923,N_2171);
nor U3782 (N_3782,N_1704,N_1550);
xnor U3783 (N_3783,N_2407,N_1942);
and U3784 (N_3784,N_2886,N_2963);
nand U3785 (N_3785,N_2254,N_2863);
xnor U3786 (N_3786,N_2637,N_2521);
and U3787 (N_3787,N_2104,N_1533);
nor U3788 (N_3788,N_2874,N_2043);
or U3789 (N_3789,N_2139,N_2600);
and U3790 (N_3790,N_2158,N_2346);
and U3791 (N_3791,N_2366,N_1904);
nand U3792 (N_3792,N_1728,N_1683);
nand U3793 (N_3793,N_1595,N_2488);
nor U3794 (N_3794,N_1787,N_1753);
and U3795 (N_3795,N_1729,N_1784);
and U3796 (N_3796,N_1796,N_1735);
xor U3797 (N_3797,N_2628,N_2534);
xnor U3798 (N_3798,N_2965,N_2670);
or U3799 (N_3799,N_2451,N_2986);
and U3800 (N_3800,N_1646,N_1939);
or U3801 (N_3801,N_2839,N_2902);
nor U3802 (N_3802,N_2796,N_2466);
or U3803 (N_3803,N_2137,N_2419);
nand U3804 (N_3804,N_2741,N_1822);
nand U3805 (N_3805,N_1563,N_2756);
and U3806 (N_3806,N_2980,N_1555);
and U3807 (N_3807,N_2998,N_1886);
nor U3808 (N_3808,N_2070,N_1874);
nand U3809 (N_3809,N_1561,N_2801);
xor U3810 (N_3810,N_1999,N_1771);
xnor U3811 (N_3811,N_2260,N_2427);
and U3812 (N_3812,N_2367,N_2245);
nor U3813 (N_3813,N_1731,N_1813);
nand U3814 (N_3814,N_1837,N_2078);
nor U3815 (N_3815,N_2470,N_1563);
nor U3816 (N_3816,N_2529,N_2363);
nand U3817 (N_3817,N_2363,N_2174);
and U3818 (N_3818,N_2506,N_1536);
nand U3819 (N_3819,N_1845,N_2746);
nand U3820 (N_3820,N_2756,N_2084);
nand U3821 (N_3821,N_1835,N_1607);
and U3822 (N_3822,N_2677,N_2984);
or U3823 (N_3823,N_2895,N_1541);
xnor U3824 (N_3824,N_2103,N_2164);
nor U3825 (N_3825,N_2030,N_2201);
and U3826 (N_3826,N_1727,N_1748);
nand U3827 (N_3827,N_1754,N_2622);
or U3828 (N_3828,N_2880,N_1531);
xnor U3829 (N_3829,N_2861,N_1830);
xnor U3830 (N_3830,N_2711,N_1725);
nor U3831 (N_3831,N_2232,N_2040);
nor U3832 (N_3832,N_2418,N_1545);
xor U3833 (N_3833,N_2850,N_2773);
and U3834 (N_3834,N_2105,N_2187);
xor U3835 (N_3835,N_2553,N_2229);
nand U3836 (N_3836,N_2538,N_1887);
xnor U3837 (N_3837,N_1571,N_2906);
nand U3838 (N_3838,N_2500,N_1932);
xnor U3839 (N_3839,N_2478,N_1868);
nor U3840 (N_3840,N_2875,N_1876);
or U3841 (N_3841,N_2329,N_1508);
xor U3842 (N_3842,N_2298,N_1901);
and U3843 (N_3843,N_2706,N_1529);
nand U3844 (N_3844,N_1984,N_2637);
xor U3845 (N_3845,N_2003,N_1827);
nor U3846 (N_3846,N_2642,N_1917);
or U3847 (N_3847,N_1830,N_2134);
nand U3848 (N_3848,N_2846,N_2741);
nor U3849 (N_3849,N_1918,N_1995);
nor U3850 (N_3850,N_2970,N_1603);
and U3851 (N_3851,N_2367,N_1949);
nand U3852 (N_3852,N_1728,N_1732);
nor U3853 (N_3853,N_2997,N_2941);
or U3854 (N_3854,N_1796,N_2783);
or U3855 (N_3855,N_2724,N_2374);
or U3856 (N_3856,N_1608,N_2243);
nor U3857 (N_3857,N_1586,N_1891);
xnor U3858 (N_3858,N_2342,N_2162);
xor U3859 (N_3859,N_2989,N_2643);
xor U3860 (N_3860,N_1568,N_1790);
nand U3861 (N_3861,N_2153,N_1928);
nor U3862 (N_3862,N_2139,N_2734);
nor U3863 (N_3863,N_2356,N_1572);
and U3864 (N_3864,N_2746,N_2441);
and U3865 (N_3865,N_2980,N_1573);
xnor U3866 (N_3866,N_2673,N_2480);
nand U3867 (N_3867,N_2748,N_2746);
xor U3868 (N_3868,N_1786,N_2213);
and U3869 (N_3869,N_2447,N_2698);
xor U3870 (N_3870,N_1601,N_2990);
or U3871 (N_3871,N_1655,N_2935);
nor U3872 (N_3872,N_2445,N_2196);
xnor U3873 (N_3873,N_1825,N_1800);
and U3874 (N_3874,N_2238,N_2769);
or U3875 (N_3875,N_2118,N_1557);
and U3876 (N_3876,N_2615,N_2312);
xnor U3877 (N_3877,N_1506,N_2280);
nand U3878 (N_3878,N_2453,N_2321);
or U3879 (N_3879,N_2347,N_1717);
nor U3880 (N_3880,N_2994,N_1532);
or U3881 (N_3881,N_1568,N_1803);
nor U3882 (N_3882,N_1949,N_2515);
and U3883 (N_3883,N_1735,N_2356);
or U3884 (N_3884,N_2896,N_2636);
or U3885 (N_3885,N_1527,N_1726);
nand U3886 (N_3886,N_1606,N_2602);
or U3887 (N_3887,N_1846,N_2195);
xnor U3888 (N_3888,N_2663,N_2897);
xor U3889 (N_3889,N_1541,N_2369);
and U3890 (N_3890,N_2753,N_1793);
and U3891 (N_3891,N_1992,N_2780);
and U3892 (N_3892,N_2301,N_2710);
nand U3893 (N_3893,N_1507,N_2840);
nor U3894 (N_3894,N_2912,N_2888);
nor U3895 (N_3895,N_1940,N_2448);
and U3896 (N_3896,N_2149,N_1820);
nand U3897 (N_3897,N_2079,N_1526);
xor U3898 (N_3898,N_2638,N_2057);
nand U3899 (N_3899,N_2703,N_2359);
or U3900 (N_3900,N_1801,N_2865);
or U3901 (N_3901,N_2665,N_2367);
xor U3902 (N_3902,N_1958,N_2357);
and U3903 (N_3903,N_2049,N_2561);
nor U3904 (N_3904,N_1501,N_2386);
xnor U3905 (N_3905,N_2310,N_2946);
nand U3906 (N_3906,N_2705,N_2267);
nand U3907 (N_3907,N_2359,N_2820);
nor U3908 (N_3908,N_2623,N_2587);
nor U3909 (N_3909,N_1850,N_2894);
and U3910 (N_3910,N_2773,N_1580);
or U3911 (N_3911,N_2621,N_1998);
and U3912 (N_3912,N_2848,N_1592);
nor U3913 (N_3913,N_2776,N_2580);
xor U3914 (N_3914,N_1526,N_1626);
nand U3915 (N_3915,N_1624,N_1822);
and U3916 (N_3916,N_2216,N_2773);
nor U3917 (N_3917,N_2374,N_1992);
nor U3918 (N_3918,N_2294,N_1819);
nor U3919 (N_3919,N_1958,N_2245);
nor U3920 (N_3920,N_2364,N_2028);
nand U3921 (N_3921,N_2614,N_2336);
xnor U3922 (N_3922,N_1854,N_2216);
nor U3923 (N_3923,N_1804,N_1918);
nand U3924 (N_3924,N_2431,N_2409);
nand U3925 (N_3925,N_1799,N_2499);
or U3926 (N_3926,N_2454,N_2032);
nor U3927 (N_3927,N_2912,N_1866);
nand U3928 (N_3928,N_2560,N_1884);
or U3929 (N_3929,N_1705,N_1743);
and U3930 (N_3930,N_2936,N_2997);
nand U3931 (N_3931,N_2523,N_1636);
and U3932 (N_3932,N_1563,N_2389);
xnor U3933 (N_3933,N_1818,N_1969);
and U3934 (N_3934,N_1965,N_1898);
nor U3935 (N_3935,N_2522,N_2682);
or U3936 (N_3936,N_2839,N_2504);
nor U3937 (N_3937,N_2312,N_1998);
and U3938 (N_3938,N_2053,N_2852);
and U3939 (N_3939,N_2525,N_2446);
and U3940 (N_3940,N_2290,N_1742);
nor U3941 (N_3941,N_1564,N_1979);
nor U3942 (N_3942,N_2294,N_1559);
xor U3943 (N_3943,N_2272,N_2106);
and U3944 (N_3944,N_1505,N_2916);
or U3945 (N_3945,N_2255,N_1821);
and U3946 (N_3946,N_1872,N_1612);
nor U3947 (N_3947,N_2577,N_1760);
or U3948 (N_3948,N_1830,N_2196);
or U3949 (N_3949,N_2845,N_1533);
or U3950 (N_3950,N_1621,N_1599);
nor U3951 (N_3951,N_2985,N_2977);
xnor U3952 (N_3952,N_1601,N_1597);
nor U3953 (N_3953,N_2782,N_2356);
xnor U3954 (N_3954,N_2007,N_1779);
or U3955 (N_3955,N_2869,N_1851);
or U3956 (N_3956,N_2998,N_2123);
or U3957 (N_3957,N_2075,N_1540);
nor U3958 (N_3958,N_1531,N_2011);
nor U3959 (N_3959,N_1976,N_1518);
xnor U3960 (N_3960,N_2062,N_1915);
nor U3961 (N_3961,N_2622,N_1603);
xor U3962 (N_3962,N_2454,N_1583);
or U3963 (N_3963,N_1667,N_2948);
or U3964 (N_3964,N_2101,N_1927);
nor U3965 (N_3965,N_2340,N_2464);
and U3966 (N_3966,N_2559,N_1501);
nor U3967 (N_3967,N_1502,N_1956);
nor U3968 (N_3968,N_2072,N_2322);
nor U3969 (N_3969,N_2644,N_1623);
or U3970 (N_3970,N_2741,N_1642);
nor U3971 (N_3971,N_2225,N_2154);
and U3972 (N_3972,N_1976,N_2193);
and U3973 (N_3973,N_2481,N_1722);
xor U3974 (N_3974,N_2582,N_2056);
nand U3975 (N_3975,N_2568,N_2689);
and U3976 (N_3976,N_2649,N_2197);
or U3977 (N_3977,N_1766,N_1704);
and U3978 (N_3978,N_2188,N_1515);
xor U3979 (N_3979,N_2669,N_2365);
xor U3980 (N_3980,N_1942,N_2483);
nand U3981 (N_3981,N_2230,N_1927);
and U3982 (N_3982,N_2754,N_2968);
xnor U3983 (N_3983,N_2989,N_2574);
nand U3984 (N_3984,N_2939,N_2973);
nand U3985 (N_3985,N_1740,N_2136);
xnor U3986 (N_3986,N_2939,N_2868);
or U3987 (N_3987,N_2769,N_2802);
nand U3988 (N_3988,N_2082,N_2079);
or U3989 (N_3989,N_2545,N_2838);
nand U3990 (N_3990,N_1694,N_2842);
nor U3991 (N_3991,N_2385,N_1912);
nor U3992 (N_3992,N_1519,N_1992);
or U3993 (N_3993,N_1621,N_2709);
or U3994 (N_3994,N_2731,N_2069);
xor U3995 (N_3995,N_1862,N_1503);
or U3996 (N_3996,N_2849,N_1908);
nor U3997 (N_3997,N_2481,N_1711);
or U3998 (N_3998,N_2578,N_2927);
or U3999 (N_3999,N_1560,N_2124);
nand U4000 (N_4000,N_2121,N_2894);
xor U4001 (N_4001,N_2862,N_1705);
nor U4002 (N_4002,N_2730,N_1852);
xor U4003 (N_4003,N_1654,N_2358);
nor U4004 (N_4004,N_2332,N_1679);
nor U4005 (N_4005,N_2499,N_2925);
or U4006 (N_4006,N_1539,N_1974);
nand U4007 (N_4007,N_2356,N_2129);
or U4008 (N_4008,N_2662,N_1560);
and U4009 (N_4009,N_2937,N_2524);
nor U4010 (N_4010,N_2107,N_2155);
and U4011 (N_4011,N_1609,N_2472);
nand U4012 (N_4012,N_2191,N_2821);
nor U4013 (N_4013,N_2036,N_2997);
or U4014 (N_4014,N_2444,N_2121);
and U4015 (N_4015,N_2719,N_2313);
xnor U4016 (N_4016,N_2085,N_1688);
nand U4017 (N_4017,N_1786,N_2331);
xor U4018 (N_4018,N_1550,N_1655);
xor U4019 (N_4019,N_2586,N_2511);
nand U4020 (N_4020,N_1739,N_2917);
nand U4021 (N_4021,N_2059,N_2070);
or U4022 (N_4022,N_2536,N_1724);
xor U4023 (N_4023,N_2217,N_2706);
nor U4024 (N_4024,N_2456,N_1880);
or U4025 (N_4025,N_1700,N_2849);
nor U4026 (N_4026,N_2249,N_1502);
nor U4027 (N_4027,N_2735,N_2603);
xor U4028 (N_4028,N_1780,N_2793);
and U4029 (N_4029,N_1704,N_1883);
nand U4030 (N_4030,N_2673,N_1621);
or U4031 (N_4031,N_2128,N_2805);
nand U4032 (N_4032,N_2116,N_2611);
nor U4033 (N_4033,N_1915,N_2417);
nand U4034 (N_4034,N_2905,N_1590);
or U4035 (N_4035,N_2530,N_1953);
and U4036 (N_4036,N_2125,N_1810);
nand U4037 (N_4037,N_2132,N_2904);
nor U4038 (N_4038,N_1964,N_1639);
nor U4039 (N_4039,N_2292,N_1992);
or U4040 (N_4040,N_1563,N_2631);
and U4041 (N_4041,N_2633,N_1570);
xnor U4042 (N_4042,N_2740,N_2028);
nand U4043 (N_4043,N_2187,N_2796);
or U4044 (N_4044,N_2528,N_1673);
nand U4045 (N_4045,N_2142,N_2323);
nand U4046 (N_4046,N_2751,N_1884);
and U4047 (N_4047,N_2944,N_2184);
xnor U4048 (N_4048,N_2932,N_2286);
nand U4049 (N_4049,N_1838,N_2460);
and U4050 (N_4050,N_2794,N_2687);
nor U4051 (N_4051,N_2510,N_2320);
or U4052 (N_4052,N_2453,N_2730);
nor U4053 (N_4053,N_2240,N_2223);
xnor U4054 (N_4054,N_2993,N_2608);
nand U4055 (N_4055,N_1832,N_2699);
xnor U4056 (N_4056,N_1598,N_2913);
nand U4057 (N_4057,N_2769,N_1871);
nand U4058 (N_4058,N_1745,N_2573);
or U4059 (N_4059,N_2960,N_2093);
and U4060 (N_4060,N_2740,N_2378);
nand U4061 (N_4061,N_2935,N_2478);
xnor U4062 (N_4062,N_2928,N_2847);
xnor U4063 (N_4063,N_2230,N_2491);
and U4064 (N_4064,N_2377,N_1564);
nor U4065 (N_4065,N_2398,N_1669);
xor U4066 (N_4066,N_2220,N_2990);
nand U4067 (N_4067,N_2090,N_1563);
xnor U4068 (N_4068,N_2246,N_2285);
nand U4069 (N_4069,N_1727,N_2470);
and U4070 (N_4070,N_2161,N_2837);
nand U4071 (N_4071,N_2630,N_1749);
nor U4072 (N_4072,N_1914,N_2875);
xor U4073 (N_4073,N_1611,N_1555);
and U4074 (N_4074,N_2679,N_1623);
nor U4075 (N_4075,N_2874,N_2633);
or U4076 (N_4076,N_2837,N_1691);
xor U4077 (N_4077,N_1725,N_2694);
nor U4078 (N_4078,N_2630,N_1637);
nor U4079 (N_4079,N_2175,N_2949);
nand U4080 (N_4080,N_2420,N_1880);
and U4081 (N_4081,N_2718,N_2239);
nand U4082 (N_4082,N_2545,N_1551);
nor U4083 (N_4083,N_1884,N_2154);
xnor U4084 (N_4084,N_1516,N_2422);
and U4085 (N_4085,N_2494,N_2587);
nand U4086 (N_4086,N_2717,N_2262);
nand U4087 (N_4087,N_1737,N_2500);
xor U4088 (N_4088,N_2389,N_1948);
xnor U4089 (N_4089,N_1848,N_2693);
xor U4090 (N_4090,N_1560,N_2066);
or U4091 (N_4091,N_2992,N_1883);
xnor U4092 (N_4092,N_2857,N_2527);
and U4093 (N_4093,N_1917,N_1972);
nand U4094 (N_4094,N_2677,N_1520);
xnor U4095 (N_4095,N_2809,N_2419);
or U4096 (N_4096,N_2143,N_2511);
or U4097 (N_4097,N_2435,N_2397);
nor U4098 (N_4098,N_1569,N_1929);
nor U4099 (N_4099,N_2973,N_2949);
nor U4100 (N_4100,N_1522,N_2473);
nand U4101 (N_4101,N_2286,N_1632);
or U4102 (N_4102,N_2785,N_1691);
and U4103 (N_4103,N_2724,N_1963);
or U4104 (N_4104,N_2140,N_2520);
or U4105 (N_4105,N_1634,N_2941);
xor U4106 (N_4106,N_2883,N_2648);
and U4107 (N_4107,N_2227,N_1950);
and U4108 (N_4108,N_2482,N_2415);
nor U4109 (N_4109,N_2615,N_2448);
nand U4110 (N_4110,N_1695,N_2786);
and U4111 (N_4111,N_2118,N_2204);
xor U4112 (N_4112,N_2141,N_1605);
or U4113 (N_4113,N_1728,N_1747);
or U4114 (N_4114,N_2696,N_2440);
nor U4115 (N_4115,N_2329,N_2858);
nor U4116 (N_4116,N_2459,N_2303);
or U4117 (N_4117,N_2235,N_1747);
nor U4118 (N_4118,N_1652,N_2378);
xor U4119 (N_4119,N_2126,N_2536);
nand U4120 (N_4120,N_1612,N_2484);
xor U4121 (N_4121,N_1908,N_2745);
nand U4122 (N_4122,N_2300,N_2535);
or U4123 (N_4123,N_2735,N_2346);
or U4124 (N_4124,N_1893,N_2799);
nor U4125 (N_4125,N_1666,N_1537);
nand U4126 (N_4126,N_2734,N_2349);
nand U4127 (N_4127,N_2582,N_1564);
or U4128 (N_4128,N_2997,N_1507);
xnor U4129 (N_4129,N_2317,N_1873);
and U4130 (N_4130,N_1949,N_2283);
or U4131 (N_4131,N_2084,N_2167);
nor U4132 (N_4132,N_2747,N_2096);
nor U4133 (N_4133,N_2140,N_2898);
and U4134 (N_4134,N_2985,N_2642);
nand U4135 (N_4135,N_1780,N_1677);
and U4136 (N_4136,N_2905,N_2157);
or U4137 (N_4137,N_2703,N_1575);
xor U4138 (N_4138,N_2073,N_2737);
or U4139 (N_4139,N_1778,N_2946);
and U4140 (N_4140,N_2525,N_2155);
nand U4141 (N_4141,N_2439,N_1591);
xor U4142 (N_4142,N_2261,N_2003);
nand U4143 (N_4143,N_2252,N_2876);
xor U4144 (N_4144,N_2226,N_1607);
nor U4145 (N_4145,N_2791,N_1685);
xnor U4146 (N_4146,N_2168,N_2618);
xnor U4147 (N_4147,N_1502,N_2396);
or U4148 (N_4148,N_2105,N_2934);
nand U4149 (N_4149,N_2792,N_1998);
xor U4150 (N_4150,N_1980,N_2751);
or U4151 (N_4151,N_2105,N_1630);
xnor U4152 (N_4152,N_1806,N_2161);
or U4153 (N_4153,N_1821,N_2945);
nand U4154 (N_4154,N_2639,N_2156);
or U4155 (N_4155,N_2723,N_2469);
nand U4156 (N_4156,N_2249,N_2134);
nand U4157 (N_4157,N_2215,N_1708);
xnor U4158 (N_4158,N_2683,N_2448);
or U4159 (N_4159,N_1983,N_1788);
or U4160 (N_4160,N_1882,N_2312);
xor U4161 (N_4161,N_2235,N_1944);
and U4162 (N_4162,N_2866,N_2613);
or U4163 (N_4163,N_1897,N_2815);
nor U4164 (N_4164,N_2044,N_2215);
xor U4165 (N_4165,N_2737,N_2653);
nand U4166 (N_4166,N_2501,N_1774);
xor U4167 (N_4167,N_2779,N_2325);
and U4168 (N_4168,N_1903,N_2433);
nand U4169 (N_4169,N_2333,N_2665);
or U4170 (N_4170,N_1647,N_2003);
and U4171 (N_4171,N_2834,N_1811);
or U4172 (N_4172,N_1904,N_2064);
or U4173 (N_4173,N_1919,N_2153);
and U4174 (N_4174,N_2650,N_1798);
nand U4175 (N_4175,N_2086,N_1808);
nor U4176 (N_4176,N_2091,N_2970);
and U4177 (N_4177,N_1883,N_2230);
nor U4178 (N_4178,N_2131,N_2217);
nor U4179 (N_4179,N_1737,N_2376);
or U4180 (N_4180,N_1611,N_2317);
xor U4181 (N_4181,N_2784,N_2747);
nor U4182 (N_4182,N_1974,N_2729);
and U4183 (N_4183,N_2007,N_2774);
or U4184 (N_4184,N_2096,N_2367);
or U4185 (N_4185,N_2039,N_2798);
and U4186 (N_4186,N_2620,N_2440);
and U4187 (N_4187,N_1565,N_2900);
or U4188 (N_4188,N_2031,N_1738);
or U4189 (N_4189,N_1901,N_1654);
nand U4190 (N_4190,N_2373,N_2802);
nand U4191 (N_4191,N_2689,N_1836);
xnor U4192 (N_4192,N_2619,N_2296);
or U4193 (N_4193,N_2551,N_1596);
nor U4194 (N_4194,N_2483,N_2911);
nor U4195 (N_4195,N_2707,N_2415);
nand U4196 (N_4196,N_1971,N_2495);
or U4197 (N_4197,N_2723,N_2636);
and U4198 (N_4198,N_2037,N_2710);
nor U4199 (N_4199,N_1847,N_1994);
xnor U4200 (N_4200,N_2018,N_1670);
and U4201 (N_4201,N_2962,N_2475);
nand U4202 (N_4202,N_2533,N_2104);
and U4203 (N_4203,N_2684,N_2801);
nand U4204 (N_4204,N_2327,N_2902);
and U4205 (N_4205,N_2055,N_1957);
or U4206 (N_4206,N_2108,N_1665);
and U4207 (N_4207,N_1660,N_2411);
xor U4208 (N_4208,N_1949,N_1866);
nand U4209 (N_4209,N_1517,N_1825);
and U4210 (N_4210,N_2226,N_2123);
nand U4211 (N_4211,N_2714,N_2424);
or U4212 (N_4212,N_1667,N_2687);
nand U4213 (N_4213,N_2121,N_2050);
nand U4214 (N_4214,N_2325,N_1710);
nor U4215 (N_4215,N_2705,N_1631);
and U4216 (N_4216,N_2266,N_2546);
or U4217 (N_4217,N_2263,N_2186);
or U4218 (N_4218,N_2130,N_2088);
or U4219 (N_4219,N_1725,N_2064);
nand U4220 (N_4220,N_2100,N_2800);
xor U4221 (N_4221,N_2717,N_1957);
or U4222 (N_4222,N_2668,N_1801);
xnor U4223 (N_4223,N_2392,N_2324);
xor U4224 (N_4224,N_1740,N_2297);
xor U4225 (N_4225,N_1507,N_2239);
xor U4226 (N_4226,N_1858,N_1994);
nor U4227 (N_4227,N_1528,N_2931);
nor U4228 (N_4228,N_1957,N_1569);
nand U4229 (N_4229,N_1824,N_1641);
nor U4230 (N_4230,N_2806,N_1574);
nand U4231 (N_4231,N_1617,N_2429);
nor U4232 (N_4232,N_2841,N_2261);
xnor U4233 (N_4233,N_2516,N_2756);
and U4234 (N_4234,N_2233,N_2581);
or U4235 (N_4235,N_2184,N_2834);
nand U4236 (N_4236,N_2206,N_1638);
and U4237 (N_4237,N_2053,N_2313);
nand U4238 (N_4238,N_2710,N_2447);
nor U4239 (N_4239,N_2186,N_2279);
nand U4240 (N_4240,N_2144,N_2192);
and U4241 (N_4241,N_1755,N_1786);
and U4242 (N_4242,N_2072,N_2567);
nor U4243 (N_4243,N_2585,N_1597);
xor U4244 (N_4244,N_1722,N_2082);
xnor U4245 (N_4245,N_1627,N_2890);
nor U4246 (N_4246,N_2725,N_2343);
and U4247 (N_4247,N_2347,N_1986);
nand U4248 (N_4248,N_2596,N_2228);
xor U4249 (N_4249,N_2133,N_2950);
and U4250 (N_4250,N_2937,N_2060);
nand U4251 (N_4251,N_2977,N_2129);
nor U4252 (N_4252,N_1921,N_1806);
and U4253 (N_4253,N_1514,N_2933);
and U4254 (N_4254,N_2953,N_1926);
and U4255 (N_4255,N_2183,N_1656);
nand U4256 (N_4256,N_1564,N_1505);
xor U4257 (N_4257,N_2143,N_2294);
nor U4258 (N_4258,N_2847,N_2372);
or U4259 (N_4259,N_1955,N_1794);
and U4260 (N_4260,N_2541,N_2966);
and U4261 (N_4261,N_1523,N_1750);
nor U4262 (N_4262,N_2496,N_2477);
and U4263 (N_4263,N_1644,N_1792);
and U4264 (N_4264,N_1886,N_1814);
nor U4265 (N_4265,N_2801,N_1536);
and U4266 (N_4266,N_2806,N_1893);
nand U4267 (N_4267,N_2133,N_2961);
or U4268 (N_4268,N_2914,N_1954);
nand U4269 (N_4269,N_2184,N_1585);
nor U4270 (N_4270,N_1809,N_2707);
and U4271 (N_4271,N_2215,N_2979);
nand U4272 (N_4272,N_2175,N_2980);
and U4273 (N_4273,N_2043,N_2957);
nor U4274 (N_4274,N_2363,N_2117);
nand U4275 (N_4275,N_1744,N_2391);
nor U4276 (N_4276,N_2510,N_2841);
and U4277 (N_4277,N_2588,N_1961);
or U4278 (N_4278,N_1757,N_2231);
and U4279 (N_4279,N_2389,N_2681);
nor U4280 (N_4280,N_1887,N_1893);
nand U4281 (N_4281,N_2646,N_2652);
or U4282 (N_4282,N_1707,N_2033);
xor U4283 (N_4283,N_2278,N_2960);
and U4284 (N_4284,N_1785,N_1566);
or U4285 (N_4285,N_2266,N_2610);
or U4286 (N_4286,N_2162,N_2132);
and U4287 (N_4287,N_2037,N_2017);
and U4288 (N_4288,N_1538,N_2737);
nor U4289 (N_4289,N_2911,N_2479);
nor U4290 (N_4290,N_2878,N_1837);
or U4291 (N_4291,N_1732,N_2064);
and U4292 (N_4292,N_2858,N_2007);
or U4293 (N_4293,N_1983,N_1589);
or U4294 (N_4294,N_2561,N_2154);
and U4295 (N_4295,N_1823,N_1814);
or U4296 (N_4296,N_1664,N_2109);
nand U4297 (N_4297,N_2157,N_2787);
nand U4298 (N_4298,N_1559,N_2365);
nand U4299 (N_4299,N_2314,N_2293);
xnor U4300 (N_4300,N_2195,N_2402);
or U4301 (N_4301,N_1746,N_2649);
and U4302 (N_4302,N_1502,N_2870);
nor U4303 (N_4303,N_1786,N_1837);
nor U4304 (N_4304,N_2137,N_2069);
or U4305 (N_4305,N_2198,N_1744);
and U4306 (N_4306,N_2798,N_2475);
or U4307 (N_4307,N_1917,N_2092);
nand U4308 (N_4308,N_2144,N_1880);
and U4309 (N_4309,N_2183,N_1521);
nor U4310 (N_4310,N_2378,N_1741);
nor U4311 (N_4311,N_1856,N_2030);
nand U4312 (N_4312,N_2408,N_2968);
xor U4313 (N_4313,N_2261,N_1965);
and U4314 (N_4314,N_1781,N_1715);
nand U4315 (N_4315,N_1814,N_1882);
and U4316 (N_4316,N_1688,N_1676);
xor U4317 (N_4317,N_2675,N_2295);
nand U4318 (N_4318,N_1755,N_2692);
nor U4319 (N_4319,N_1813,N_2184);
nand U4320 (N_4320,N_1871,N_2463);
nor U4321 (N_4321,N_2521,N_2451);
nand U4322 (N_4322,N_2099,N_1941);
and U4323 (N_4323,N_2908,N_2126);
and U4324 (N_4324,N_2217,N_1630);
nand U4325 (N_4325,N_2067,N_2753);
nor U4326 (N_4326,N_2282,N_2945);
nor U4327 (N_4327,N_2982,N_1607);
xnor U4328 (N_4328,N_1646,N_2316);
nand U4329 (N_4329,N_1852,N_2529);
nand U4330 (N_4330,N_2354,N_1622);
nor U4331 (N_4331,N_1967,N_1509);
and U4332 (N_4332,N_2888,N_2275);
xor U4333 (N_4333,N_2515,N_1853);
xnor U4334 (N_4334,N_2935,N_1770);
xor U4335 (N_4335,N_2076,N_2482);
and U4336 (N_4336,N_2444,N_1578);
and U4337 (N_4337,N_2252,N_2010);
nand U4338 (N_4338,N_2062,N_1538);
nor U4339 (N_4339,N_1865,N_2586);
xor U4340 (N_4340,N_2518,N_2584);
xnor U4341 (N_4341,N_1903,N_2795);
nand U4342 (N_4342,N_2869,N_2293);
or U4343 (N_4343,N_2199,N_2848);
or U4344 (N_4344,N_2131,N_2506);
nor U4345 (N_4345,N_2038,N_2413);
and U4346 (N_4346,N_2074,N_2177);
and U4347 (N_4347,N_2984,N_2673);
or U4348 (N_4348,N_1881,N_2801);
or U4349 (N_4349,N_2981,N_2756);
or U4350 (N_4350,N_2119,N_1668);
and U4351 (N_4351,N_2704,N_1643);
and U4352 (N_4352,N_2823,N_1576);
and U4353 (N_4353,N_1851,N_1779);
nor U4354 (N_4354,N_2854,N_1819);
and U4355 (N_4355,N_2744,N_2851);
or U4356 (N_4356,N_1568,N_1719);
nor U4357 (N_4357,N_2295,N_2664);
nor U4358 (N_4358,N_2265,N_2386);
xnor U4359 (N_4359,N_1931,N_2521);
xor U4360 (N_4360,N_1999,N_2503);
and U4361 (N_4361,N_2897,N_2546);
and U4362 (N_4362,N_2709,N_1720);
xor U4363 (N_4363,N_1818,N_1901);
or U4364 (N_4364,N_2227,N_2694);
or U4365 (N_4365,N_2289,N_2176);
nand U4366 (N_4366,N_2175,N_2896);
and U4367 (N_4367,N_2987,N_2770);
or U4368 (N_4368,N_2171,N_1720);
nor U4369 (N_4369,N_1535,N_2949);
nor U4370 (N_4370,N_2571,N_2572);
and U4371 (N_4371,N_2700,N_2630);
nand U4372 (N_4372,N_2343,N_2727);
nand U4373 (N_4373,N_2712,N_2804);
and U4374 (N_4374,N_1655,N_1671);
xor U4375 (N_4375,N_2730,N_2298);
xor U4376 (N_4376,N_2501,N_2672);
xnor U4377 (N_4377,N_2233,N_2547);
nor U4378 (N_4378,N_2369,N_2791);
nand U4379 (N_4379,N_1729,N_2549);
and U4380 (N_4380,N_2348,N_2082);
or U4381 (N_4381,N_2188,N_1763);
nor U4382 (N_4382,N_2317,N_1638);
nor U4383 (N_4383,N_2642,N_2773);
xor U4384 (N_4384,N_2538,N_2941);
nor U4385 (N_4385,N_2477,N_2423);
nand U4386 (N_4386,N_1660,N_2282);
or U4387 (N_4387,N_2910,N_2328);
and U4388 (N_4388,N_2953,N_2886);
nand U4389 (N_4389,N_2469,N_1600);
nand U4390 (N_4390,N_1866,N_1767);
or U4391 (N_4391,N_2550,N_2209);
and U4392 (N_4392,N_2611,N_2878);
xnor U4393 (N_4393,N_2918,N_2646);
nand U4394 (N_4394,N_1587,N_2044);
and U4395 (N_4395,N_2384,N_1603);
xnor U4396 (N_4396,N_2647,N_2577);
or U4397 (N_4397,N_2464,N_1514);
nor U4398 (N_4398,N_2744,N_2501);
nor U4399 (N_4399,N_2270,N_1717);
xor U4400 (N_4400,N_2538,N_2713);
nand U4401 (N_4401,N_1928,N_2255);
or U4402 (N_4402,N_1666,N_2749);
and U4403 (N_4403,N_2981,N_2986);
xor U4404 (N_4404,N_2603,N_1738);
nand U4405 (N_4405,N_2257,N_1874);
nor U4406 (N_4406,N_2742,N_1882);
nand U4407 (N_4407,N_1797,N_2999);
nand U4408 (N_4408,N_1550,N_1603);
or U4409 (N_4409,N_2310,N_2689);
and U4410 (N_4410,N_1517,N_1780);
and U4411 (N_4411,N_1628,N_2240);
nor U4412 (N_4412,N_2091,N_1892);
and U4413 (N_4413,N_2302,N_1811);
nand U4414 (N_4414,N_2802,N_1628);
and U4415 (N_4415,N_2405,N_2673);
nor U4416 (N_4416,N_1585,N_2527);
or U4417 (N_4417,N_2741,N_2533);
and U4418 (N_4418,N_2545,N_2258);
xor U4419 (N_4419,N_2875,N_1993);
nand U4420 (N_4420,N_2146,N_2326);
xnor U4421 (N_4421,N_2958,N_1561);
nor U4422 (N_4422,N_2953,N_1840);
or U4423 (N_4423,N_2892,N_2958);
nor U4424 (N_4424,N_1950,N_2264);
or U4425 (N_4425,N_1574,N_2379);
or U4426 (N_4426,N_2838,N_1868);
or U4427 (N_4427,N_1865,N_1582);
and U4428 (N_4428,N_2479,N_2790);
xor U4429 (N_4429,N_1998,N_2056);
and U4430 (N_4430,N_1895,N_2740);
xor U4431 (N_4431,N_2917,N_1919);
or U4432 (N_4432,N_2187,N_2837);
and U4433 (N_4433,N_1856,N_1886);
nor U4434 (N_4434,N_1807,N_2412);
nand U4435 (N_4435,N_1870,N_2369);
xnor U4436 (N_4436,N_2970,N_2714);
and U4437 (N_4437,N_2073,N_1979);
and U4438 (N_4438,N_1561,N_2638);
nor U4439 (N_4439,N_2026,N_1655);
or U4440 (N_4440,N_2829,N_2961);
nor U4441 (N_4441,N_1854,N_1820);
nor U4442 (N_4442,N_2048,N_2698);
or U4443 (N_4443,N_1883,N_1723);
nor U4444 (N_4444,N_1901,N_1799);
and U4445 (N_4445,N_1574,N_1513);
nand U4446 (N_4446,N_1713,N_2040);
and U4447 (N_4447,N_2134,N_2847);
or U4448 (N_4448,N_2506,N_2061);
and U4449 (N_4449,N_1734,N_2439);
or U4450 (N_4450,N_2655,N_1578);
and U4451 (N_4451,N_1749,N_2815);
xor U4452 (N_4452,N_1975,N_1544);
nor U4453 (N_4453,N_2871,N_2897);
or U4454 (N_4454,N_2099,N_1578);
nor U4455 (N_4455,N_1509,N_1814);
nor U4456 (N_4456,N_1721,N_2214);
and U4457 (N_4457,N_2870,N_1759);
nand U4458 (N_4458,N_1834,N_1820);
nor U4459 (N_4459,N_2307,N_1803);
or U4460 (N_4460,N_1992,N_2340);
or U4461 (N_4461,N_2659,N_1840);
xnor U4462 (N_4462,N_2651,N_2687);
nor U4463 (N_4463,N_2765,N_2966);
nand U4464 (N_4464,N_2843,N_2816);
xor U4465 (N_4465,N_2708,N_2310);
nand U4466 (N_4466,N_2825,N_1977);
xor U4467 (N_4467,N_2942,N_2341);
xor U4468 (N_4468,N_1665,N_2228);
xor U4469 (N_4469,N_2702,N_2720);
nor U4470 (N_4470,N_2106,N_1775);
xnor U4471 (N_4471,N_1972,N_1583);
or U4472 (N_4472,N_2761,N_2025);
xor U4473 (N_4473,N_1696,N_1611);
and U4474 (N_4474,N_2746,N_1853);
and U4475 (N_4475,N_2774,N_1882);
and U4476 (N_4476,N_2501,N_2642);
nand U4477 (N_4477,N_2407,N_2971);
xor U4478 (N_4478,N_1742,N_1995);
xnor U4479 (N_4479,N_1990,N_2160);
nor U4480 (N_4480,N_2414,N_2390);
xor U4481 (N_4481,N_2437,N_1711);
or U4482 (N_4482,N_2885,N_2311);
or U4483 (N_4483,N_1660,N_2949);
or U4484 (N_4484,N_1513,N_2760);
and U4485 (N_4485,N_1805,N_2210);
nor U4486 (N_4486,N_1763,N_1995);
or U4487 (N_4487,N_2942,N_1610);
nand U4488 (N_4488,N_1883,N_2724);
nor U4489 (N_4489,N_2967,N_2850);
and U4490 (N_4490,N_1757,N_2884);
and U4491 (N_4491,N_2810,N_1724);
or U4492 (N_4492,N_2687,N_2826);
nand U4493 (N_4493,N_2826,N_2823);
xor U4494 (N_4494,N_1936,N_2321);
nor U4495 (N_4495,N_1538,N_2000);
nor U4496 (N_4496,N_2092,N_2267);
nor U4497 (N_4497,N_1711,N_2817);
nand U4498 (N_4498,N_1948,N_1610);
or U4499 (N_4499,N_2282,N_2542);
nor U4500 (N_4500,N_4283,N_3526);
nand U4501 (N_4501,N_4238,N_3270);
or U4502 (N_4502,N_3607,N_4147);
or U4503 (N_4503,N_4004,N_3938);
xnor U4504 (N_4504,N_3757,N_4233);
xnor U4505 (N_4505,N_4080,N_4208);
nand U4506 (N_4506,N_3698,N_3040);
nor U4507 (N_4507,N_3703,N_3684);
xor U4508 (N_4508,N_3795,N_4273);
and U4509 (N_4509,N_4166,N_3858);
and U4510 (N_4510,N_3305,N_4054);
xnor U4511 (N_4511,N_3244,N_3919);
xor U4512 (N_4512,N_4011,N_3697);
nand U4513 (N_4513,N_4258,N_3925);
nand U4514 (N_4514,N_3895,N_3852);
and U4515 (N_4515,N_3171,N_3057);
nor U4516 (N_4516,N_3649,N_4017);
and U4517 (N_4517,N_4456,N_3495);
nand U4518 (N_4518,N_3226,N_3561);
nand U4519 (N_4519,N_3358,N_4149);
nor U4520 (N_4520,N_3438,N_3751);
and U4521 (N_4521,N_3902,N_4463);
xnor U4522 (N_4522,N_4406,N_3179);
nor U4523 (N_4523,N_3664,N_4188);
nor U4524 (N_4524,N_4352,N_3245);
nor U4525 (N_4525,N_3142,N_3110);
or U4526 (N_4526,N_4223,N_3399);
nand U4527 (N_4527,N_3683,N_3378);
and U4528 (N_4528,N_4007,N_3178);
xor U4529 (N_4529,N_3654,N_4246);
nand U4530 (N_4530,N_4105,N_4446);
xnor U4531 (N_4531,N_3322,N_3967);
and U4532 (N_4532,N_3312,N_3289);
or U4533 (N_4533,N_3194,N_3500);
and U4534 (N_4534,N_4315,N_3651);
nand U4535 (N_4535,N_3007,N_3294);
nor U4536 (N_4536,N_3141,N_3523);
nor U4537 (N_4537,N_3944,N_4150);
and U4538 (N_4538,N_3304,N_3137);
nand U4539 (N_4539,N_3782,N_3799);
and U4540 (N_4540,N_3617,N_4178);
or U4541 (N_4541,N_4085,N_3791);
nor U4542 (N_4542,N_4099,N_4399);
or U4543 (N_4543,N_3609,N_3672);
nand U4544 (N_4544,N_3911,N_3994);
nand U4545 (N_4545,N_3143,N_3477);
nand U4546 (N_4546,N_4202,N_3231);
nand U4547 (N_4547,N_4061,N_3360);
nand U4548 (N_4548,N_4047,N_4340);
or U4549 (N_4549,N_4376,N_3107);
xor U4550 (N_4550,N_3824,N_3892);
nor U4551 (N_4551,N_3413,N_3434);
xnor U4552 (N_4552,N_4341,N_3655);
or U4553 (N_4553,N_3104,N_3302);
nand U4554 (N_4554,N_4324,N_3564);
xnor U4555 (N_4555,N_4420,N_3927);
nand U4556 (N_4556,N_3088,N_4243);
nand U4557 (N_4557,N_4318,N_3868);
and U4558 (N_4558,N_3855,N_3769);
nand U4559 (N_4559,N_3587,N_4335);
or U4560 (N_4560,N_3470,N_4450);
or U4561 (N_4561,N_4018,N_3993);
nor U4562 (N_4562,N_4417,N_3329);
xnor U4563 (N_4563,N_3350,N_3199);
or U4564 (N_4564,N_3287,N_3206);
or U4565 (N_4565,N_3550,N_3459);
or U4566 (N_4566,N_3317,N_4141);
and U4567 (N_4567,N_4476,N_3699);
xnor U4568 (N_4568,N_4441,N_3484);
nor U4569 (N_4569,N_3374,N_3532);
and U4570 (N_4570,N_3908,N_4186);
nand U4571 (N_4571,N_3825,N_3747);
xor U4572 (N_4572,N_3991,N_3840);
nor U4573 (N_4573,N_3363,N_3503);
or U4574 (N_4574,N_4302,N_3439);
and U4575 (N_4575,N_4371,N_4355);
and U4576 (N_4576,N_4016,N_4232);
xnor U4577 (N_4577,N_3924,N_4155);
xnor U4578 (N_4578,N_3801,N_4364);
xnor U4579 (N_4579,N_3268,N_3539);
and U4580 (N_4580,N_3036,N_4343);
or U4581 (N_4581,N_3722,N_3075);
nor U4582 (N_4582,N_3514,N_3511);
nand U4583 (N_4583,N_4266,N_3468);
and U4584 (N_4584,N_3936,N_3656);
and U4585 (N_4585,N_3754,N_3896);
or U4586 (N_4586,N_3133,N_3690);
nor U4587 (N_4587,N_3429,N_3175);
and U4588 (N_4588,N_3262,N_4192);
nor U4589 (N_4589,N_3394,N_4091);
xnor U4590 (N_4590,N_3267,N_3610);
and U4591 (N_4591,N_3996,N_3592);
nor U4592 (N_4592,N_3233,N_3605);
nand U4593 (N_4593,N_3202,N_3682);
nand U4594 (N_4594,N_3725,N_4056);
and U4595 (N_4595,N_4485,N_3787);
or U4596 (N_4596,N_3701,N_3939);
nor U4597 (N_4597,N_3685,N_3349);
xor U4598 (N_4598,N_3890,N_3531);
nor U4599 (N_4599,N_3430,N_3147);
nor U4600 (N_4600,N_3023,N_4311);
nor U4601 (N_4601,N_3885,N_3044);
or U4602 (N_4602,N_4455,N_4052);
nor U4603 (N_4603,N_3021,N_3945);
nand U4604 (N_4604,N_3424,N_3116);
nor U4605 (N_4605,N_4127,N_4372);
xor U4606 (N_4606,N_4419,N_3060);
nor U4607 (N_4607,N_3743,N_3876);
xor U4608 (N_4608,N_3686,N_4444);
nor U4609 (N_4609,N_4298,N_4452);
or U4610 (N_4610,N_4221,N_3827);
xor U4611 (N_4611,N_3594,N_3674);
nor U4612 (N_4612,N_4103,N_3185);
and U4613 (N_4613,N_4251,N_3650);
nand U4614 (N_4614,N_3385,N_3337);
and U4615 (N_4615,N_4079,N_4136);
nand U4616 (N_4616,N_4317,N_3067);
xnor U4617 (N_4617,N_4070,N_3572);
or U4618 (N_4618,N_4236,N_4365);
xor U4619 (N_4619,N_3081,N_3553);
nor U4620 (N_4620,N_3933,N_4433);
or U4621 (N_4621,N_4249,N_3502);
xor U4622 (N_4622,N_3538,N_3750);
nand U4623 (N_4623,N_4415,N_4271);
xor U4624 (N_4624,N_4351,N_4021);
xor U4625 (N_4625,N_4043,N_3992);
and U4626 (N_4626,N_3145,N_3386);
and U4627 (N_4627,N_4133,N_3059);
and U4628 (N_4628,N_3762,N_3746);
nand U4629 (N_4629,N_3208,N_4164);
xor U4630 (N_4630,N_4130,N_4175);
or U4631 (N_4631,N_3006,N_3548);
nor U4632 (N_4632,N_4140,N_3634);
xnor U4633 (N_4633,N_3913,N_3794);
xor U4634 (N_4634,N_3547,N_4228);
or U4635 (N_4635,N_4129,N_4459);
and U4636 (N_4636,N_4388,N_3872);
and U4637 (N_4637,N_3718,N_3956);
xor U4638 (N_4638,N_3311,N_3022);
nand U4639 (N_4639,N_3519,N_3481);
and U4640 (N_4640,N_4436,N_4405);
nor U4641 (N_4641,N_3014,N_3125);
or U4642 (N_4642,N_3368,N_3983);
nand U4643 (N_4643,N_3448,N_3971);
xnor U4644 (N_4644,N_3668,N_4172);
and U4645 (N_4645,N_3980,N_3155);
or U4646 (N_4646,N_3087,N_3755);
nand U4647 (N_4647,N_3739,N_4297);
and U4648 (N_4648,N_3917,N_4499);
nor U4649 (N_4649,N_3345,N_4193);
and U4650 (N_4650,N_3623,N_3536);
nand U4651 (N_4651,N_3589,N_3761);
xnor U4652 (N_4652,N_3367,N_4473);
xor U4653 (N_4653,N_3600,N_3570);
nor U4654 (N_4654,N_3568,N_4305);
xnor U4655 (N_4655,N_3065,N_3844);
nor U4656 (N_4656,N_3643,N_4231);
or U4657 (N_4657,N_3581,N_4074);
nand U4658 (N_4658,N_3916,N_3721);
nand U4659 (N_4659,N_3440,N_4209);
nand U4660 (N_4660,N_4346,N_3770);
nand U4661 (N_4661,N_4124,N_3445);
and U4662 (N_4662,N_3841,N_3461);
or U4663 (N_4663,N_3476,N_3740);
nand U4664 (N_4664,N_3928,N_3606);
or U4665 (N_4665,N_3598,N_4089);
nor U4666 (N_4666,N_3615,N_4391);
and U4667 (N_4667,N_4219,N_4057);
xnor U4668 (N_4668,N_3223,N_3574);
or U4669 (N_4669,N_3264,N_4214);
or U4670 (N_4670,N_4122,N_4240);
nor U4671 (N_4671,N_4160,N_3348);
and U4672 (N_4672,N_3914,N_4458);
xnor U4673 (N_4673,N_3156,N_3324);
xnor U4674 (N_4674,N_4098,N_4237);
nand U4675 (N_4675,N_3639,N_3681);
or U4676 (N_4676,N_4220,N_3658);
nand U4677 (N_4677,N_3818,N_3249);
or U4678 (N_4678,N_4059,N_3988);
nand U4679 (N_4679,N_4010,N_4218);
and U4680 (N_4680,N_3077,N_4337);
nand U4681 (N_4681,N_3567,N_3869);
nor U4682 (N_4682,N_3113,N_3693);
nor U4683 (N_4683,N_3237,N_3850);
xor U4684 (N_4684,N_3978,N_4312);
or U4685 (N_4685,N_3504,N_3719);
or U4686 (N_4686,N_3677,N_3976);
xnor U4687 (N_4687,N_3546,N_3282);
xor U4688 (N_4688,N_3704,N_3792);
nand U4689 (N_4689,N_4134,N_3128);
nand U4690 (N_4690,N_3160,N_4264);
or U4691 (N_4691,N_3291,N_4263);
or U4692 (N_4692,N_4148,N_3714);
or U4693 (N_4693,N_4483,N_3744);
or U4694 (N_4694,N_4050,N_4287);
and U4695 (N_4695,N_4395,N_4029);
or U4696 (N_4696,N_3576,N_3695);
nor U4697 (N_4697,N_4006,N_3426);
or U4698 (N_4698,N_3063,N_3715);
nor U4699 (N_4699,N_3454,N_4062);
nor U4700 (N_4700,N_3975,N_3165);
nor U4701 (N_4701,N_4397,N_4204);
and U4702 (N_4702,N_3853,N_3167);
xor U4703 (N_4703,N_4008,N_3357);
xor U4704 (N_4704,N_3987,N_3030);
nand U4705 (N_4705,N_3709,N_3256);
nor U4706 (N_4706,N_3675,N_3497);
nand U4707 (N_4707,N_3344,N_3313);
xor U4708 (N_4708,N_4215,N_4115);
or U4709 (N_4709,N_3730,N_3056);
or U4710 (N_4710,N_4101,N_4300);
and U4711 (N_4711,N_3472,N_4229);
nor U4712 (N_4712,N_4443,N_3408);
or U4713 (N_4713,N_3033,N_4082);
and U4714 (N_4714,N_3877,N_4146);
nand U4715 (N_4715,N_3188,N_3420);
or U4716 (N_4716,N_3402,N_3129);
and U4717 (N_4717,N_3507,N_3665);
nand U4718 (N_4718,N_3947,N_4469);
xnor U4719 (N_4719,N_3802,N_4083);
xnor U4720 (N_4720,N_4400,N_3276);
nand U4721 (N_4721,N_4296,N_3122);
nor U4722 (N_4722,N_4170,N_4189);
and U4723 (N_4723,N_3549,N_3804);
nor U4724 (N_4724,N_4037,N_3283);
nand U4725 (N_4725,N_3124,N_3181);
nor U4726 (N_4726,N_3280,N_3152);
xnor U4727 (N_4727,N_3281,N_4470);
xor U4728 (N_4728,N_3882,N_3227);
xnor U4729 (N_4729,N_3275,N_4191);
nand U4730 (N_4730,N_3812,N_3432);
and U4731 (N_4731,N_3772,N_4289);
and U4732 (N_4732,N_4457,N_3333);
xor U4733 (N_4733,N_3901,N_4200);
nand U4734 (N_4734,N_4131,N_3816);
xnor U4735 (N_4735,N_3528,N_3320);
or U4736 (N_4736,N_3427,N_4269);
nor U4737 (N_4737,N_4109,N_4316);
xor U4738 (N_4738,N_4216,N_3451);
and U4739 (N_4739,N_3222,N_3661);
or U4740 (N_4740,N_3300,N_3692);
xnor U4741 (N_4741,N_4496,N_3881);
and U4742 (N_4742,N_4291,N_3020);
nor U4743 (N_4743,N_4087,N_4253);
or U4744 (N_4744,N_4490,N_3422);
and U4745 (N_4745,N_3829,N_3789);
nand U4746 (N_4746,N_3334,N_4358);
nand U4747 (N_4747,N_4320,N_3177);
or U4748 (N_4748,N_3613,N_3608);
xnor U4749 (N_4749,N_4326,N_3702);
nor U4750 (N_4750,N_4381,N_3308);
nand U4751 (N_4751,N_3105,N_3867);
nand U4752 (N_4752,N_3214,N_3575);
and U4753 (N_4753,N_3204,N_3341);
nor U4754 (N_4754,N_4184,N_3555);
and U4755 (N_4755,N_3323,N_3585);
nand U4756 (N_4756,N_4256,N_3590);
and U4757 (N_4757,N_3455,N_4117);
xnor U4758 (N_4758,N_4396,N_3493);
xnor U4759 (N_4759,N_4331,N_3870);
and U4760 (N_4760,N_3964,N_3370);
xnor U4761 (N_4761,N_3663,N_3298);
nor U4762 (N_4762,N_4033,N_4308);
xnor U4763 (N_4763,N_4234,N_3577);
or U4764 (N_4764,N_3893,N_3954);
and U4765 (N_4765,N_3960,N_3635);
nand U4766 (N_4766,N_3773,N_4063);
or U4767 (N_4767,N_3387,N_4479);
nand U4768 (N_4768,N_4142,N_4494);
and U4769 (N_4769,N_3252,N_3198);
or U4770 (N_4770,N_3392,N_3046);
nand U4771 (N_4771,N_3571,N_4487);
nor U4772 (N_4772,N_3073,N_4427);
and U4773 (N_4773,N_3708,N_4112);
nand U4774 (N_4774,N_4138,N_3779);
nand U4775 (N_4775,N_3900,N_3910);
xnor U4776 (N_4776,N_3723,N_3015);
and U4777 (N_4777,N_4418,N_3002);
nor U4778 (N_4778,N_3330,N_3086);
xor U4779 (N_4779,N_3447,N_3273);
or U4780 (N_4780,N_3494,N_3948);
or U4781 (N_4781,N_3053,N_3822);
and U4782 (N_4782,N_3398,N_4026);
nor U4783 (N_4783,N_4268,N_4244);
xnor U4784 (N_4784,N_3132,N_4199);
nor U4785 (N_4785,N_4387,N_3688);
nor U4786 (N_4786,N_3437,N_4267);
nor U4787 (N_4787,N_3364,N_3071);
nand U4788 (N_4788,N_3638,N_3640);
or U4789 (N_4789,N_3163,N_3080);
nand U4790 (N_4790,N_4116,N_3602);
and U4791 (N_4791,N_3471,N_4293);
and U4792 (N_4792,N_4180,N_4314);
or U4793 (N_4793,N_3213,N_3534);
and U4794 (N_4794,N_3186,N_4414);
nand U4795 (N_4795,N_3556,N_3017);
xor U4796 (N_4796,N_3100,N_4250);
nand U4797 (N_4797,N_3859,N_3771);
xnor U4798 (N_4798,N_3647,N_3235);
nand U4799 (N_4799,N_4161,N_4309);
or U4800 (N_4800,N_3274,N_3756);
or U4801 (N_4801,N_4448,N_3084);
and U4802 (N_4802,N_3079,N_3894);
nor U4803 (N_4803,N_3166,N_3042);
nor U4804 (N_4804,N_4386,N_3940);
and U4805 (N_4805,N_4440,N_3596);
nand U4806 (N_4806,N_3403,N_3072);
xnor U4807 (N_4807,N_3362,N_3431);
xor U4808 (N_4808,N_4349,N_3094);
nor U4809 (N_4809,N_3009,N_3636);
nand U4810 (N_4810,N_3452,N_4282);
and U4811 (N_4811,N_4489,N_3215);
xor U4812 (N_4812,N_4097,N_3808);
xnor U4813 (N_4813,N_3612,N_4128);
and U4814 (N_4814,N_3819,N_3096);
xor U4815 (N_4815,N_3051,N_3909);
xnor U4816 (N_4816,N_4075,N_3485);
and U4817 (N_4817,N_3981,N_3565);
or U4818 (N_4818,N_4212,N_3149);
or U4819 (N_4819,N_4278,N_3435);
xnor U4820 (N_4820,N_4145,N_4373);
nand U4821 (N_4821,N_4435,N_3845);
xnor U4822 (N_4822,N_3527,N_3466);
nand U4823 (N_4823,N_3524,N_4461);
and U4824 (N_4824,N_3669,N_3217);
or U4825 (N_4825,N_3083,N_4077);
nand U4826 (N_4826,N_4286,N_3284);
nor U4827 (N_4827,N_4183,N_3707);
xor U4828 (N_4828,N_3417,N_4424);
or U4829 (N_4829,N_3336,N_3689);
nand U4830 (N_4830,N_3515,N_3098);
nor U4831 (N_4831,N_3182,N_4409);
and U4832 (N_4832,N_3783,N_3861);
xor U4833 (N_4833,N_3114,N_4053);
or U4834 (N_4834,N_3535,N_3196);
nand U4835 (N_4835,N_3776,N_3935);
xnor U4836 (N_4836,N_3260,N_3835);
and U4837 (N_4837,N_4167,N_3295);
or U4838 (N_4838,N_4205,N_3106);
nor U4839 (N_4839,N_4323,N_3250);
xor U4840 (N_4840,N_4000,N_3729);
and U4841 (N_4841,N_4247,N_3279);
nor U4842 (N_4842,N_3011,N_3097);
or U4843 (N_4843,N_3599,N_3013);
or U4844 (N_4844,N_4295,N_4153);
xor U4845 (N_4845,N_3229,N_3923);
and U4846 (N_4846,N_4431,N_4102);
nor U4847 (N_4847,N_3153,N_3319);
or U4848 (N_4848,N_3095,N_3745);
nand U4849 (N_4849,N_3162,N_4347);
and U4850 (N_4850,N_3849,N_3306);
nand U4851 (N_4851,N_4367,N_3483);
and U4852 (N_4852,N_3405,N_3173);
nand U4853 (N_4853,N_3700,N_4094);
and U4854 (N_4854,N_3443,N_4350);
nor U4855 (N_4855,N_3154,N_4190);
or U4856 (N_4856,N_4241,N_4125);
and U4857 (N_4857,N_4447,N_3800);
nand U4858 (N_4858,N_3673,N_3788);
nand U4859 (N_4859,N_3614,N_3506);
or U4860 (N_4860,N_3254,N_4252);
nand U4861 (N_4861,N_3292,N_3404);
nor U4862 (N_4862,N_3343,N_3520);
nor U4863 (N_4863,N_4173,N_4464);
and U4864 (N_4864,N_4438,N_3931);
nand U4865 (N_4865,N_3469,N_3463);
or U4866 (N_4866,N_3865,N_3525);
nor U4867 (N_4867,N_3836,N_3629);
and U4868 (N_4868,N_4211,N_3921);
or U4869 (N_4869,N_3460,N_3748);
nor U4870 (N_4870,N_3889,N_3411);
nand U4871 (N_4871,N_4475,N_4361);
and U4872 (N_4872,N_3860,N_3462);
or U4873 (N_4873,N_3959,N_4303);
or U4874 (N_4874,N_3878,N_3251);
and U4875 (N_4875,N_3726,N_3982);
xor U4876 (N_4876,N_4428,N_4374);
nor U4877 (N_4877,N_3480,N_3657);
and U4878 (N_4878,N_4046,N_3863);
nand U4879 (N_4879,N_4044,N_3724);
and U4880 (N_4880,N_4255,N_4123);
nand U4881 (N_4881,N_3365,N_4009);
nor U4882 (N_4882,N_3028,N_3004);
or U4883 (N_4883,N_3225,N_4156);
nor U4884 (N_4884,N_3645,N_4334);
nand U4885 (N_4885,N_3588,N_3115);
xor U4886 (N_4886,N_3584,N_3929);
nand U4887 (N_4887,N_4113,N_4272);
nand U4888 (N_4888,N_3326,N_3738);
nand U4889 (N_4889,N_3915,N_3180);
or U4890 (N_4890,N_3529,N_4327);
or U4891 (N_4891,N_3218,N_4275);
and U4892 (N_4892,N_4380,N_3321);
xnor U4893 (N_4893,N_3332,N_3784);
and U4894 (N_4894,N_3003,N_3338);
nor U4895 (N_4895,N_3346,N_3421);
nand U4896 (N_4896,N_3966,N_4158);
nand U4897 (N_4897,N_3604,N_3621);
or U4898 (N_4898,N_3101,N_3691);
nand U4899 (N_4899,N_3958,N_3817);
nand U4900 (N_4900,N_3027,N_3126);
or U4901 (N_4901,N_4022,N_3379);
nor U4902 (N_4902,N_3828,N_3170);
or U4903 (N_4903,N_3316,N_4493);
xnor U4904 (N_4904,N_3595,N_3626);
xor U4905 (N_4905,N_3798,N_3766);
nor U4906 (N_4906,N_3029,N_3000);
and U4907 (N_4907,N_4306,N_3382);
xnor U4908 (N_4908,N_4462,N_3951);
or U4909 (N_4909,N_3339,N_3873);
nand U4910 (N_4910,N_3168,N_4423);
or U4911 (N_4911,N_4096,N_4338);
or U4912 (N_4912,N_3157,N_3832);
or U4913 (N_4913,N_3781,N_3545);
nor U4914 (N_4914,N_3957,N_4279);
and U4915 (N_4915,N_3016,N_3705);
xor U4916 (N_4916,N_3353,N_4333);
and U4917 (N_4917,N_4430,N_3834);
nor U4918 (N_4918,N_4321,N_3962);
or U4919 (N_4919,N_4472,N_3209);
nor U4920 (N_4920,N_3409,N_3941);
nand U4921 (N_4921,N_3039,N_3973);
nor U4922 (N_4922,N_3487,N_4362);
or U4923 (N_4923,N_3236,N_3591);
nor U4924 (N_4924,N_3395,N_3499);
and U4925 (N_4925,N_3191,N_4495);
and U4926 (N_4926,N_3415,N_4329);
nor U4927 (N_4927,N_4261,N_3898);
nor U4928 (N_4928,N_3542,N_4084);
nor U4929 (N_4929,N_4114,N_3920);
nor U4930 (N_4930,N_4280,N_3883);
and U4931 (N_4931,N_3340,N_3012);
nor U4932 (N_4932,N_3752,N_3266);
nor U4933 (N_4933,N_4014,N_4195);
xnor U4934 (N_4934,N_3479,N_3049);
or U4935 (N_4935,N_3625,N_3174);
or U4936 (N_4936,N_3243,N_3307);
xor U4937 (N_4937,N_4345,N_3052);
nand U4938 (N_4938,N_3880,N_4210);
or U4939 (N_4939,N_3995,N_3735);
nor U4940 (N_4940,N_3820,N_4379);
and U4941 (N_4941,N_3833,N_3904);
or U4942 (N_4942,N_4181,N_4377);
or U4943 (N_4943,N_3372,N_3031);
xnor U4944 (N_4944,N_4299,N_4072);
xor U4945 (N_4945,N_3774,N_3058);
xnor U4946 (N_4946,N_3790,N_3169);
xnor U4947 (N_4947,N_4437,N_3257);
and U4948 (N_4948,N_3670,N_3884);
xor U4949 (N_4949,N_3297,N_4393);
or U4950 (N_4950,N_3847,N_4151);
xor U4951 (N_4951,N_3303,N_3117);
nor U4952 (N_4952,N_3239,N_3024);
nor U4953 (N_4953,N_4310,N_3158);
and U4954 (N_4954,N_4325,N_4132);
or U4955 (N_4955,N_4226,N_3391);
nor U4956 (N_4956,N_3373,N_3619);
xor U4957 (N_4957,N_4254,N_3963);
nor U4958 (N_4958,N_4168,N_3741);
nor U4959 (N_4959,N_3777,N_4005);
nor U4960 (N_4960,N_3134,N_3473);
nand U4961 (N_4961,N_3176,N_3008);
or U4962 (N_4962,N_3823,N_3102);
or U4963 (N_4963,N_3522,N_3821);
nor U4964 (N_4964,N_3566,N_3839);
nand U4965 (N_4965,N_3069,N_3666);
nor U4966 (N_4966,N_3355,N_4019);
and U4967 (N_4967,N_3573,N_4265);
nand U4968 (N_4968,N_4319,N_4404);
nand U4969 (N_4969,N_3293,N_4126);
nor U4970 (N_4970,N_4139,N_3785);
nor U4971 (N_4971,N_3247,N_3159);
xor U4972 (N_4972,N_4093,N_4179);
and U4973 (N_4973,N_4067,N_4432);
nand U4974 (N_4974,N_3441,N_3197);
xnor U4975 (N_4975,N_3488,N_3758);
nor U4976 (N_4976,N_3035,N_3383);
and U4977 (N_4977,N_4027,N_4344);
nand U4978 (N_4978,N_3622,N_3230);
nor U4979 (N_4979,N_3616,N_4051);
nor U4980 (N_4980,N_3109,N_3457);
or U4981 (N_4981,N_4292,N_3050);
and U4982 (N_4982,N_3809,N_3136);
nand U4983 (N_4983,N_3261,N_3559);
nand U4984 (N_4984,N_4086,N_3676);
and U4985 (N_4985,N_4230,N_3127);
and U4986 (N_4986,N_3864,N_4012);
or U4987 (N_4987,N_3371,N_3263);
nor U4988 (N_4988,N_3121,N_3637);
or U4989 (N_4989,N_3899,N_4259);
nor U4990 (N_4990,N_3135,N_3793);
nand U4991 (N_4991,N_3361,N_4045);
nor U4992 (N_4992,N_4366,N_3150);
nor U4993 (N_4993,N_3203,N_4270);
xor U4994 (N_4994,N_4330,N_4294);
or U4995 (N_4995,N_4171,N_3767);
nor U4996 (N_4996,N_3120,N_4454);
nand U4997 (N_4997,N_3043,N_3089);
and U4998 (N_4998,N_3811,N_3854);
and U4999 (N_4999,N_3148,N_4492);
xnor U5000 (N_5000,N_3711,N_3753);
or U5001 (N_5001,N_3093,N_3512);
or U5002 (N_5002,N_3659,N_3146);
and U5003 (N_5003,N_3796,N_3418);
nor U5004 (N_5004,N_4137,N_4385);
or U5005 (N_5005,N_3765,N_3414);
nor U5006 (N_5006,N_4023,N_4328);
nor U5007 (N_5007,N_3848,N_4357);
xnor U5008 (N_5008,N_3189,N_4071);
xor U5009 (N_5009,N_3221,N_3513);
nor U5010 (N_5010,N_3815,N_3489);
and U5011 (N_5011,N_4144,N_4110);
nor U5012 (N_5012,N_3554,N_3200);
nand U5013 (N_5013,N_3974,N_3026);
or U5014 (N_5014,N_4486,N_4066);
xor U5015 (N_5015,N_3130,N_3641);
nor U5016 (N_5016,N_3201,N_4488);
or U5017 (N_5017,N_3055,N_3271);
or U5018 (N_5018,N_3038,N_3047);
xnor U5019 (N_5019,N_3578,N_3749);
nor U5020 (N_5020,N_3648,N_4162);
nor U5021 (N_5021,N_3679,N_3558);
and U5022 (N_5022,N_4368,N_4135);
nand U5023 (N_5023,N_3579,N_3453);
xnor U5024 (N_5024,N_3351,N_3240);
xnor U5025 (N_5025,N_3342,N_4453);
or U5026 (N_5026,N_4092,N_3140);
nor U5027 (N_5027,N_3569,N_3627);
and U5028 (N_5028,N_3464,N_3837);
nand U5029 (N_5029,N_3248,N_3482);
or U5030 (N_5030,N_3064,N_3517);
nor U5031 (N_5031,N_3210,N_3205);
nand U5032 (N_5032,N_3376,N_3212);
nand U5033 (N_5033,N_4058,N_3803);
or U5034 (N_5034,N_4100,N_3986);
nand U5035 (N_5035,N_4106,N_3667);
or U5036 (N_5036,N_3710,N_4354);
and U5037 (N_5037,N_3025,N_3259);
xnor U5038 (N_5038,N_3897,N_3680);
xnor U5039 (N_5039,N_3032,N_3846);
or U5040 (N_5040,N_3074,N_4198);
nor U5041 (N_5041,N_3377,N_3492);
nand U5042 (N_5042,N_3934,N_3242);
nor U5043 (N_5043,N_3359,N_3888);
nand U5044 (N_5044,N_4451,N_4078);
nand U5045 (N_5045,N_4336,N_3078);
xor U5046 (N_5046,N_4260,N_3131);
xor U5047 (N_5047,N_4410,N_4426);
and U5048 (N_5048,N_4143,N_4108);
or U5049 (N_5049,N_3068,N_4095);
and U5050 (N_5050,N_3301,N_3428);
and U5051 (N_5051,N_3632,N_3874);
xor U5052 (N_5052,N_3552,N_3253);
nand U5053 (N_5053,N_4040,N_3932);
and U5054 (N_5054,N_3092,N_3216);
and U5055 (N_5055,N_4090,N_3611);
or U5056 (N_5056,N_4356,N_3269);
and U5057 (N_5057,N_4384,N_3325);
and U5058 (N_5058,N_3760,N_3597);
or U5059 (N_5059,N_4425,N_3108);
nand U5060 (N_5060,N_3396,N_3763);
nor U5061 (N_5061,N_4201,N_3694);
nor U5062 (N_5062,N_3423,N_4163);
or U5063 (N_5063,N_3985,N_4088);
nor U5064 (N_5064,N_3436,N_4304);
nor U5065 (N_5065,N_3583,N_3943);
nor U5066 (N_5066,N_3618,N_4360);
xnor U5067 (N_5067,N_3458,N_3331);
nor U5068 (N_5068,N_4025,N_4482);
xnor U5069 (N_5069,N_3090,N_3593);
nand U5070 (N_5070,N_3544,N_3857);
xor U5071 (N_5071,N_3687,N_3949);
nor U5072 (N_5072,N_4392,N_3410);
nor U5073 (N_5073,N_3970,N_3805);
xor U5074 (N_5074,N_4342,N_3989);
or U5075 (N_5075,N_4001,N_4245);
xor U5076 (N_5076,N_4307,N_3838);
and U5077 (N_5077,N_3258,N_3123);
or U5078 (N_5078,N_3562,N_3728);
nor U5079 (N_5079,N_3384,N_4119);
and U5080 (N_5080,N_3318,N_4407);
and U5081 (N_5081,N_4111,N_4081);
xnor U5082 (N_5082,N_4322,N_3509);
xor U5083 (N_5083,N_3151,N_3732);
nand U5084 (N_5084,N_3419,N_3891);
xor U5085 (N_5085,N_3620,N_3630);
nand U5086 (N_5086,N_3219,N_3112);
and U5087 (N_5087,N_4032,N_3644);
nor U5088 (N_5088,N_3082,N_4107);
or U5089 (N_5089,N_4174,N_3510);
or U5090 (N_5090,N_3918,N_3875);
nor U5091 (N_5091,N_3490,N_4348);
and U5092 (N_5092,N_3813,N_3521);
and U5093 (N_5093,N_3830,N_3193);
and U5094 (N_5094,N_3653,N_3907);
xnor U5095 (N_5095,N_3786,N_4020);
xor U5096 (N_5096,N_4498,N_3955);
nand U5097 (N_5097,N_3491,N_3518);
nand U5098 (N_5098,N_4313,N_3062);
or U5099 (N_5099,N_3190,N_3232);
nand U5100 (N_5100,N_4442,N_4466);
nor U5101 (N_5101,N_4378,N_4068);
nand U5102 (N_5102,N_3652,N_3449);
and U5103 (N_5103,N_3633,N_3843);
nand U5104 (N_5104,N_3990,N_3400);
and U5105 (N_5105,N_3646,N_3731);
nand U5106 (N_5106,N_3508,N_3501);
nand U5107 (N_5107,N_3290,N_3224);
and U5108 (N_5108,N_3034,N_4382);
xor U5109 (N_5109,N_3906,N_3706);
or U5110 (N_5110,N_3866,N_3851);
and U5111 (N_5111,N_3352,N_3972);
xnor U5112 (N_5112,N_3717,N_4480);
nand U5113 (N_5113,N_3187,N_4104);
nor U5114 (N_5114,N_4467,N_4030);
nor U5115 (N_5115,N_4227,N_4239);
and U5116 (N_5116,N_3733,N_4034);
or U5117 (N_5117,N_4398,N_4169);
or U5118 (N_5118,N_4481,N_3272);
and U5119 (N_5119,N_4048,N_3207);
and U5120 (N_5120,N_3968,N_3328);
nand U5121 (N_5121,N_3950,N_3161);
nor U5122 (N_5122,N_4439,N_3807);
nor U5123 (N_5123,N_3085,N_4217);
or U5124 (N_5124,N_4235,N_3862);
nand U5125 (N_5125,N_4497,N_3366);
xor U5126 (N_5126,N_3465,N_3712);
nand U5127 (N_5127,N_3347,N_3335);
nor U5128 (N_5128,N_4434,N_3952);
xnor U5129 (N_5129,N_3797,N_4197);
and U5130 (N_5130,N_4274,N_3211);
xnor U5131 (N_5131,N_3642,N_3380);
nor U5132 (N_5132,N_4038,N_3977);
nand U5133 (N_5133,N_3091,N_3433);
nand U5134 (N_5134,N_4154,N_3879);
and U5135 (N_5135,N_4383,N_3425);
nor U5136 (N_5136,N_4049,N_3887);
or U5137 (N_5137,N_3192,N_3238);
and U5138 (N_5138,N_3164,N_3456);
and U5139 (N_5139,N_4301,N_3118);
and U5140 (N_5140,N_4035,N_4262);
nor U5141 (N_5141,N_3814,N_3764);
nor U5142 (N_5142,N_3624,N_4339);
and U5143 (N_5143,N_4449,N_4353);
xor U5144 (N_5144,N_3716,N_4248);
nand U5145 (N_5145,N_3582,N_3327);
nor U5146 (N_5146,N_3314,N_3099);
or U5147 (N_5147,N_3184,N_4390);
nand U5148 (N_5148,N_3389,N_3942);
and U5149 (N_5149,N_4242,N_4389);
nand U5150 (N_5150,N_4196,N_4468);
nor U5151 (N_5151,N_3228,N_4363);
or U5152 (N_5152,N_3183,N_3671);
and U5153 (N_5153,N_3005,N_3139);
xnor U5154 (N_5154,N_4402,N_4478);
nor U5155 (N_5155,N_4036,N_3780);
nand U5156 (N_5156,N_3019,N_3277);
or U5157 (N_5157,N_4064,N_3937);
xnor U5158 (N_5158,N_3903,N_3416);
and U5159 (N_5159,N_3001,N_3530);
nor U5160 (N_5160,N_3969,N_3580);
nand U5161 (N_5161,N_3486,N_4411);
nor U5162 (N_5162,N_4073,N_3631);
xnor U5163 (N_5163,N_3768,N_4491);
xor U5164 (N_5164,N_3999,N_3720);
xnor U5165 (N_5165,N_4288,N_3048);
nand U5166 (N_5166,N_3543,N_4277);
xor U5167 (N_5167,N_3241,N_3930);
and U5168 (N_5168,N_4055,N_3286);
or U5169 (N_5169,N_3288,N_3478);
or U5170 (N_5170,N_4065,N_4421);
nand U5171 (N_5171,N_3010,N_3467);
xnor U5172 (N_5172,N_3998,N_3778);
xor U5173 (N_5173,N_4465,N_3736);
nor U5174 (N_5174,N_3138,N_3397);
nor U5175 (N_5175,N_4165,N_4224);
nand U5176 (N_5176,N_4477,N_4460);
xnor U5177 (N_5177,N_3742,N_3054);
or U5178 (N_5178,N_3111,N_3381);
or U5179 (N_5179,N_3965,N_4015);
and U5180 (N_5180,N_4285,N_3922);
xor U5181 (N_5181,N_3541,N_3540);
nand U5182 (N_5182,N_3401,N_3912);
or U5183 (N_5183,N_3871,N_3563);
xor U5184 (N_5184,N_3103,N_4187);
nor U5185 (N_5185,N_4118,N_4069);
or U5186 (N_5186,N_3406,N_3810);
or U5187 (N_5187,N_3551,N_4222);
nor U5188 (N_5188,N_3678,N_3195);
nor U5189 (N_5189,N_3037,N_3660);
nand U5190 (N_5190,N_4028,N_4159);
and U5191 (N_5191,N_4207,N_3450);
xnor U5192 (N_5192,N_4401,N_3713);
and U5193 (N_5193,N_4002,N_4121);
nand U5194 (N_5194,N_3953,N_4290);
and U5195 (N_5195,N_3375,N_3560);
xnor U5196 (N_5196,N_4120,N_3388);
nor U5197 (N_5197,N_3533,N_4257);
nand U5198 (N_5198,N_4213,N_3979);
and U5199 (N_5199,N_3356,N_4369);
and U5200 (N_5200,N_3390,N_3309);
nand U5201 (N_5201,N_3842,N_3172);
or U5202 (N_5202,N_3265,N_4408);
nor U5203 (N_5203,N_3061,N_4474);
nand U5204 (N_5204,N_4276,N_4484);
xor U5205 (N_5205,N_4422,N_3537);
nor U5206 (N_5206,N_4375,N_3255);
and U5207 (N_5207,N_4157,N_4152);
or U5208 (N_5208,N_3557,N_3299);
nor U5209 (N_5209,N_3727,N_3601);
xnor U5210 (N_5210,N_4041,N_4031);
xnor U5211 (N_5211,N_4024,N_4039);
nor U5212 (N_5212,N_3412,N_3474);
nor U5213 (N_5213,N_3734,N_3070);
and U5214 (N_5214,N_3278,N_3926);
and U5215 (N_5215,N_3119,N_3628);
nand U5216 (N_5216,N_3826,N_3446);
and U5217 (N_5217,N_4359,N_4225);
xnor U5218 (N_5218,N_3354,N_3505);
xnor U5219 (N_5219,N_4182,N_3407);
nand U5220 (N_5220,N_4445,N_3234);
nand U5221 (N_5221,N_4176,N_4413);
or U5222 (N_5222,N_4281,N_3516);
xor U5223 (N_5223,N_3696,N_3806);
nand U5224 (N_5224,N_3315,N_3961);
and U5225 (N_5225,N_4003,N_3759);
and U5226 (N_5226,N_4013,N_3997);
nand U5227 (N_5227,N_4416,N_4042);
and U5228 (N_5228,N_3285,N_3737);
nand U5229 (N_5229,N_3444,N_4284);
nand U5230 (N_5230,N_3775,N_3886);
and U5231 (N_5231,N_3018,N_3045);
and U5232 (N_5232,N_3369,N_4177);
and U5233 (N_5233,N_4403,N_3041);
nor U5234 (N_5234,N_4206,N_3393);
nor U5235 (N_5235,N_4076,N_3984);
nand U5236 (N_5236,N_3066,N_3442);
xnor U5237 (N_5237,N_3310,N_3662);
or U5238 (N_5238,N_3076,N_4194);
nand U5239 (N_5239,N_4060,N_4185);
or U5240 (N_5240,N_4394,N_3946);
nand U5241 (N_5241,N_3475,N_3496);
xnor U5242 (N_5242,N_3498,N_4203);
nand U5243 (N_5243,N_4471,N_4332);
nand U5244 (N_5244,N_4370,N_4412);
or U5245 (N_5245,N_3586,N_3905);
or U5246 (N_5246,N_3603,N_3144);
nand U5247 (N_5247,N_3246,N_3856);
nand U5248 (N_5248,N_3831,N_4429);
and U5249 (N_5249,N_3220,N_3296);
and U5250 (N_5250,N_3698,N_4254);
and U5251 (N_5251,N_3799,N_3043);
nand U5252 (N_5252,N_4400,N_3364);
or U5253 (N_5253,N_3521,N_3528);
xnor U5254 (N_5254,N_4300,N_4301);
and U5255 (N_5255,N_4366,N_3658);
and U5256 (N_5256,N_3895,N_3478);
and U5257 (N_5257,N_3410,N_4235);
nand U5258 (N_5258,N_4004,N_4170);
and U5259 (N_5259,N_4229,N_4346);
or U5260 (N_5260,N_3070,N_4161);
and U5261 (N_5261,N_4124,N_3687);
and U5262 (N_5262,N_3692,N_3989);
and U5263 (N_5263,N_4461,N_3328);
and U5264 (N_5264,N_3752,N_3134);
nand U5265 (N_5265,N_3086,N_3970);
nand U5266 (N_5266,N_3970,N_4054);
or U5267 (N_5267,N_3368,N_3177);
xor U5268 (N_5268,N_3810,N_4153);
nor U5269 (N_5269,N_4147,N_4483);
xnor U5270 (N_5270,N_4484,N_3519);
nand U5271 (N_5271,N_3957,N_4307);
and U5272 (N_5272,N_4133,N_3375);
nor U5273 (N_5273,N_4147,N_4284);
xor U5274 (N_5274,N_4378,N_3670);
nand U5275 (N_5275,N_3745,N_4313);
xor U5276 (N_5276,N_3449,N_3424);
or U5277 (N_5277,N_3987,N_3756);
nor U5278 (N_5278,N_3664,N_3697);
xor U5279 (N_5279,N_3728,N_3805);
nor U5280 (N_5280,N_3930,N_3242);
nand U5281 (N_5281,N_3112,N_3073);
xnor U5282 (N_5282,N_4181,N_3055);
or U5283 (N_5283,N_3718,N_4115);
nand U5284 (N_5284,N_3802,N_3535);
nand U5285 (N_5285,N_3347,N_3528);
xnor U5286 (N_5286,N_4344,N_3597);
nor U5287 (N_5287,N_3482,N_4363);
xnor U5288 (N_5288,N_3621,N_4219);
and U5289 (N_5289,N_4059,N_3702);
or U5290 (N_5290,N_3361,N_4433);
xnor U5291 (N_5291,N_3621,N_3400);
nor U5292 (N_5292,N_3909,N_4289);
nor U5293 (N_5293,N_3867,N_4035);
xor U5294 (N_5294,N_4304,N_3978);
or U5295 (N_5295,N_3007,N_3580);
nor U5296 (N_5296,N_3000,N_4307);
and U5297 (N_5297,N_3496,N_3869);
or U5298 (N_5298,N_3312,N_3296);
or U5299 (N_5299,N_3970,N_3675);
or U5300 (N_5300,N_4457,N_3630);
and U5301 (N_5301,N_3100,N_4227);
nor U5302 (N_5302,N_3161,N_3025);
and U5303 (N_5303,N_4232,N_4172);
nand U5304 (N_5304,N_3524,N_3460);
and U5305 (N_5305,N_3284,N_4347);
nor U5306 (N_5306,N_3851,N_3795);
nor U5307 (N_5307,N_4399,N_3075);
and U5308 (N_5308,N_3217,N_4236);
nor U5309 (N_5309,N_3369,N_3113);
xnor U5310 (N_5310,N_4490,N_3675);
nand U5311 (N_5311,N_4022,N_4338);
nor U5312 (N_5312,N_3862,N_3425);
and U5313 (N_5313,N_3637,N_3011);
nand U5314 (N_5314,N_3776,N_3010);
xor U5315 (N_5315,N_4306,N_4203);
nor U5316 (N_5316,N_3223,N_3178);
nor U5317 (N_5317,N_3892,N_3232);
nor U5318 (N_5318,N_3710,N_3610);
or U5319 (N_5319,N_3495,N_3424);
and U5320 (N_5320,N_3166,N_4242);
nand U5321 (N_5321,N_4095,N_4081);
nand U5322 (N_5322,N_3221,N_3467);
nand U5323 (N_5323,N_4122,N_4008);
nand U5324 (N_5324,N_3346,N_3341);
nor U5325 (N_5325,N_3057,N_3748);
xor U5326 (N_5326,N_3903,N_3486);
and U5327 (N_5327,N_4258,N_4068);
and U5328 (N_5328,N_4293,N_3325);
or U5329 (N_5329,N_4099,N_4035);
nor U5330 (N_5330,N_4479,N_4293);
xor U5331 (N_5331,N_3629,N_3731);
or U5332 (N_5332,N_3278,N_4015);
xnor U5333 (N_5333,N_3203,N_3749);
and U5334 (N_5334,N_4161,N_4392);
nand U5335 (N_5335,N_3407,N_3257);
nor U5336 (N_5336,N_4188,N_3027);
or U5337 (N_5337,N_3536,N_4289);
or U5338 (N_5338,N_3813,N_4131);
nand U5339 (N_5339,N_3131,N_3023);
nor U5340 (N_5340,N_3104,N_4245);
xnor U5341 (N_5341,N_3324,N_3761);
xor U5342 (N_5342,N_3149,N_3724);
nand U5343 (N_5343,N_4325,N_3376);
xor U5344 (N_5344,N_4480,N_4307);
nand U5345 (N_5345,N_3572,N_4463);
xnor U5346 (N_5346,N_3920,N_4048);
or U5347 (N_5347,N_3040,N_3964);
nor U5348 (N_5348,N_3611,N_4292);
xor U5349 (N_5349,N_4135,N_4429);
and U5350 (N_5350,N_4357,N_3798);
xnor U5351 (N_5351,N_4186,N_3282);
xor U5352 (N_5352,N_3951,N_3551);
and U5353 (N_5353,N_3100,N_3003);
nor U5354 (N_5354,N_3967,N_4012);
xnor U5355 (N_5355,N_3392,N_4303);
nor U5356 (N_5356,N_3938,N_4281);
nor U5357 (N_5357,N_3861,N_3100);
xnor U5358 (N_5358,N_4289,N_4032);
xnor U5359 (N_5359,N_3902,N_3605);
and U5360 (N_5360,N_3197,N_3690);
nor U5361 (N_5361,N_4173,N_3837);
xnor U5362 (N_5362,N_4201,N_4164);
or U5363 (N_5363,N_3923,N_4461);
or U5364 (N_5364,N_3456,N_3775);
or U5365 (N_5365,N_3727,N_3481);
nand U5366 (N_5366,N_3649,N_4459);
nor U5367 (N_5367,N_3207,N_3940);
xnor U5368 (N_5368,N_4486,N_3106);
xor U5369 (N_5369,N_4165,N_3619);
or U5370 (N_5370,N_4338,N_4105);
nor U5371 (N_5371,N_4345,N_3322);
nor U5372 (N_5372,N_4355,N_3620);
nand U5373 (N_5373,N_4423,N_3454);
or U5374 (N_5374,N_4471,N_4054);
and U5375 (N_5375,N_3333,N_4217);
or U5376 (N_5376,N_3519,N_3490);
and U5377 (N_5377,N_3222,N_3224);
or U5378 (N_5378,N_3007,N_4365);
nor U5379 (N_5379,N_3907,N_3033);
nor U5380 (N_5380,N_3474,N_3190);
or U5381 (N_5381,N_3327,N_4291);
nand U5382 (N_5382,N_3687,N_3858);
and U5383 (N_5383,N_3455,N_3245);
xnor U5384 (N_5384,N_4196,N_4421);
or U5385 (N_5385,N_3005,N_3871);
and U5386 (N_5386,N_4398,N_3994);
xnor U5387 (N_5387,N_3174,N_3994);
or U5388 (N_5388,N_3780,N_3079);
and U5389 (N_5389,N_3978,N_3225);
and U5390 (N_5390,N_3285,N_4083);
and U5391 (N_5391,N_4029,N_3521);
and U5392 (N_5392,N_3191,N_4280);
and U5393 (N_5393,N_4178,N_4275);
nand U5394 (N_5394,N_3292,N_4128);
xor U5395 (N_5395,N_3586,N_4467);
and U5396 (N_5396,N_3362,N_3964);
and U5397 (N_5397,N_3680,N_3876);
or U5398 (N_5398,N_3189,N_4323);
nor U5399 (N_5399,N_4074,N_3249);
nor U5400 (N_5400,N_3668,N_3212);
nand U5401 (N_5401,N_3548,N_3944);
xor U5402 (N_5402,N_4344,N_4422);
nor U5403 (N_5403,N_4058,N_3389);
xor U5404 (N_5404,N_3823,N_3931);
xor U5405 (N_5405,N_3193,N_3286);
and U5406 (N_5406,N_4174,N_3254);
nor U5407 (N_5407,N_4110,N_4183);
nand U5408 (N_5408,N_3738,N_4362);
xor U5409 (N_5409,N_4052,N_4171);
nand U5410 (N_5410,N_4458,N_3203);
and U5411 (N_5411,N_3370,N_3451);
nand U5412 (N_5412,N_3658,N_3428);
and U5413 (N_5413,N_3686,N_4087);
nand U5414 (N_5414,N_3072,N_3849);
or U5415 (N_5415,N_4242,N_3237);
xor U5416 (N_5416,N_3442,N_4483);
nor U5417 (N_5417,N_3464,N_4268);
nor U5418 (N_5418,N_3053,N_4326);
nand U5419 (N_5419,N_3951,N_3369);
xor U5420 (N_5420,N_3187,N_3815);
nor U5421 (N_5421,N_3189,N_4270);
and U5422 (N_5422,N_3389,N_3124);
nor U5423 (N_5423,N_4145,N_4429);
nand U5424 (N_5424,N_3455,N_3466);
nand U5425 (N_5425,N_3922,N_3100);
xor U5426 (N_5426,N_4167,N_4158);
and U5427 (N_5427,N_4092,N_3193);
nor U5428 (N_5428,N_3956,N_4352);
nor U5429 (N_5429,N_3743,N_4377);
nand U5430 (N_5430,N_3758,N_3237);
xor U5431 (N_5431,N_3029,N_3344);
and U5432 (N_5432,N_3359,N_3033);
nor U5433 (N_5433,N_4069,N_3058);
nor U5434 (N_5434,N_4337,N_3941);
or U5435 (N_5435,N_3689,N_4204);
xnor U5436 (N_5436,N_3476,N_4381);
nand U5437 (N_5437,N_3169,N_3453);
and U5438 (N_5438,N_3332,N_3302);
nand U5439 (N_5439,N_3504,N_4021);
and U5440 (N_5440,N_3565,N_3783);
and U5441 (N_5441,N_4179,N_4290);
and U5442 (N_5442,N_3409,N_3098);
xor U5443 (N_5443,N_3814,N_3171);
and U5444 (N_5444,N_4081,N_3619);
and U5445 (N_5445,N_4388,N_4409);
or U5446 (N_5446,N_3751,N_3367);
or U5447 (N_5447,N_3565,N_3947);
xor U5448 (N_5448,N_3744,N_3065);
nand U5449 (N_5449,N_4210,N_3138);
xor U5450 (N_5450,N_3526,N_4021);
nor U5451 (N_5451,N_3909,N_3523);
or U5452 (N_5452,N_3011,N_3423);
xor U5453 (N_5453,N_3510,N_4489);
nand U5454 (N_5454,N_3343,N_3460);
nor U5455 (N_5455,N_3328,N_4255);
and U5456 (N_5456,N_4463,N_3057);
or U5457 (N_5457,N_4340,N_4115);
or U5458 (N_5458,N_4101,N_4118);
nor U5459 (N_5459,N_3389,N_3556);
or U5460 (N_5460,N_3419,N_3533);
or U5461 (N_5461,N_3747,N_3229);
nand U5462 (N_5462,N_3013,N_4042);
xor U5463 (N_5463,N_3774,N_3591);
nand U5464 (N_5464,N_4364,N_3775);
xnor U5465 (N_5465,N_4190,N_3356);
and U5466 (N_5466,N_4078,N_4222);
or U5467 (N_5467,N_3900,N_4473);
or U5468 (N_5468,N_4281,N_4121);
xnor U5469 (N_5469,N_3191,N_4439);
nand U5470 (N_5470,N_3780,N_3472);
and U5471 (N_5471,N_4299,N_4368);
nor U5472 (N_5472,N_3873,N_4204);
and U5473 (N_5473,N_3710,N_4425);
nand U5474 (N_5474,N_3722,N_3595);
xor U5475 (N_5475,N_4305,N_3214);
or U5476 (N_5476,N_3112,N_3768);
xor U5477 (N_5477,N_3823,N_4175);
nor U5478 (N_5478,N_3211,N_3712);
nor U5479 (N_5479,N_4267,N_3500);
and U5480 (N_5480,N_3098,N_3646);
xnor U5481 (N_5481,N_3993,N_3337);
or U5482 (N_5482,N_4270,N_3527);
or U5483 (N_5483,N_3445,N_3706);
and U5484 (N_5484,N_3225,N_3783);
nand U5485 (N_5485,N_3757,N_4440);
and U5486 (N_5486,N_4337,N_3205);
or U5487 (N_5487,N_4375,N_3637);
nand U5488 (N_5488,N_3325,N_4015);
or U5489 (N_5489,N_4256,N_3125);
nor U5490 (N_5490,N_4338,N_3683);
xnor U5491 (N_5491,N_3707,N_4112);
nor U5492 (N_5492,N_3122,N_3746);
xor U5493 (N_5493,N_4172,N_3591);
nand U5494 (N_5494,N_3581,N_3059);
and U5495 (N_5495,N_4371,N_3091);
nor U5496 (N_5496,N_3322,N_3870);
nor U5497 (N_5497,N_3128,N_3658);
xor U5498 (N_5498,N_3134,N_3632);
and U5499 (N_5499,N_3131,N_4420);
or U5500 (N_5500,N_3423,N_3242);
and U5501 (N_5501,N_4467,N_3998);
xnor U5502 (N_5502,N_4204,N_3289);
xnor U5503 (N_5503,N_3638,N_3580);
xnor U5504 (N_5504,N_3516,N_3425);
nor U5505 (N_5505,N_3464,N_4230);
or U5506 (N_5506,N_4407,N_3416);
xor U5507 (N_5507,N_3536,N_4181);
xnor U5508 (N_5508,N_4476,N_3289);
or U5509 (N_5509,N_4192,N_3426);
or U5510 (N_5510,N_3077,N_4361);
nand U5511 (N_5511,N_4175,N_4323);
nor U5512 (N_5512,N_4428,N_3093);
nor U5513 (N_5513,N_3391,N_3153);
nand U5514 (N_5514,N_4045,N_4080);
and U5515 (N_5515,N_4067,N_3606);
xor U5516 (N_5516,N_3995,N_3094);
xor U5517 (N_5517,N_4393,N_3766);
nand U5518 (N_5518,N_3498,N_3536);
nor U5519 (N_5519,N_4161,N_4001);
nand U5520 (N_5520,N_4488,N_4353);
or U5521 (N_5521,N_3595,N_4005);
nor U5522 (N_5522,N_4088,N_4087);
xnor U5523 (N_5523,N_3249,N_3433);
and U5524 (N_5524,N_3936,N_4161);
or U5525 (N_5525,N_3693,N_3915);
nor U5526 (N_5526,N_3734,N_4339);
nand U5527 (N_5527,N_4018,N_3122);
nand U5528 (N_5528,N_4117,N_3419);
or U5529 (N_5529,N_3840,N_3676);
and U5530 (N_5530,N_3274,N_4415);
xnor U5531 (N_5531,N_4186,N_3818);
or U5532 (N_5532,N_3623,N_3424);
xnor U5533 (N_5533,N_4240,N_3765);
nand U5534 (N_5534,N_3338,N_3290);
nand U5535 (N_5535,N_3890,N_3982);
nor U5536 (N_5536,N_3678,N_3006);
or U5537 (N_5537,N_3893,N_3409);
or U5538 (N_5538,N_3209,N_3867);
and U5539 (N_5539,N_3357,N_4122);
xor U5540 (N_5540,N_3183,N_3017);
nand U5541 (N_5541,N_4189,N_3520);
nand U5542 (N_5542,N_3198,N_3216);
xor U5543 (N_5543,N_4143,N_3427);
or U5544 (N_5544,N_3187,N_3605);
and U5545 (N_5545,N_3648,N_3026);
or U5546 (N_5546,N_3468,N_3060);
xnor U5547 (N_5547,N_3748,N_4189);
nor U5548 (N_5548,N_4146,N_4124);
and U5549 (N_5549,N_3403,N_3268);
and U5550 (N_5550,N_3558,N_3977);
and U5551 (N_5551,N_3010,N_3558);
nor U5552 (N_5552,N_4403,N_4291);
and U5553 (N_5553,N_3890,N_3231);
nand U5554 (N_5554,N_3961,N_3050);
xnor U5555 (N_5555,N_3593,N_3917);
or U5556 (N_5556,N_3173,N_4356);
and U5557 (N_5557,N_4079,N_4328);
nor U5558 (N_5558,N_3651,N_4494);
nor U5559 (N_5559,N_4194,N_3370);
and U5560 (N_5560,N_3717,N_3812);
nand U5561 (N_5561,N_4402,N_3500);
or U5562 (N_5562,N_3491,N_4229);
or U5563 (N_5563,N_4278,N_3520);
nor U5564 (N_5564,N_3443,N_4287);
and U5565 (N_5565,N_3620,N_3538);
nor U5566 (N_5566,N_3336,N_3508);
and U5567 (N_5567,N_3829,N_3510);
and U5568 (N_5568,N_3399,N_3007);
nand U5569 (N_5569,N_4244,N_3798);
nor U5570 (N_5570,N_4172,N_3688);
nor U5571 (N_5571,N_3447,N_3863);
xor U5572 (N_5572,N_3029,N_3041);
and U5573 (N_5573,N_3503,N_3257);
xor U5574 (N_5574,N_4414,N_3601);
and U5575 (N_5575,N_3932,N_3654);
or U5576 (N_5576,N_3461,N_3738);
nand U5577 (N_5577,N_3149,N_4361);
nor U5578 (N_5578,N_4172,N_4434);
or U5579 (N_5579,N_3269,N_3919);
nand U5580 (N_5580,N_3243,N_3397);
nand U5581 (N_5581,N_3276,N_4308);
or U5582 (N_5582,N_3126,N_4412);
nor U5583 (N_5583,N_4014,N_3905);
nor U5584 (N_5584,N_3840,N_3596);
nand U5585 (N_5585,N_3546,N_3884);
nand U5586 (N_5586,N_3444,N_3083);
or U5587 (N_5587,N_4497,N_4195);
or U5588 (N_5588,N_3843,N_4031);
or U5589 (N_5589,N_4045,N_4282);
nor U5590 (N_5590,N_3713,N_3382);
nand U5591 (N_5591,N_4089,N_3211);
nor U5592 (N_5592,N_3163,N_3159);
and U5593 (N_5593,N_3862,N_3269);
nor U5594 (N_5594,N_3452,N_4357);
nand U5595 (N_5595,N_3601,N_4244);
and U5596 (N_5596,N_3546,N_3780);
and U5597 (N_5597,N_4296,N_3257);
and U5598 (N_5598,N_3092,N_4251);
and U5599 (N_5599,N_4473,N_4482);
or U5600 (N_5600,N_3908,N_4269);
and U5601 (N_5601,N_4499,N_4416);
xnor U5602 (N_5602,N_3017,N_4235);
xor U5603 (N_5603,N_4141,N_4216);
xnor U5604 (N_5604,N_3984,N_3621);
or U5605 (N_5605,N_3928,N_4486);
nor U5606 (N_5606,N_3505,N_3449);
and U5607 (N_5607,N_4394,N_3163);
xor U5608 (N_5608,N_3748,N_3397);
xor U5609 (N_5609,N_4479,N_3092);
and U5610 (N_5610,N_4044,N_3502);
nand U5611 (N_5611,N_3969,N_3917);
nor U5612 (N_5612,N_3514,N_3172);
nand U5613 (N_5613,N_3985,N_3133);
and U5614 (N_5614,N_4091,N_3696);
xnor U5615 (N_5615,N_3595,N_4121);
nand U5616 (N_5616,N_4117,N_3698);
xnor U5617 (N_5617,N_3249,N_4141);
and U5618 (N_5618,N_4370,N_4402);
nor U5619 (N_5619,N_3952,N_4156);
or U5620 (N_5620,N_4102,N_3306);
nand U5621 (N_5621,N_4443,N_3998);
and U5622 (N_5622,N_3109,N_3191);
xnor U5623 (N_5623,N_3523,N_3276);
and U5624 (N_5624,N_3147,N_4386);
and U5625 (N_5625,N_3986,N_3159);
nand U5626 (N_5626,N_4499,N_4342);
nand U5627 (N_5627,N_4452,N_3472);
nor U5628 (N_5628,N_4025,N_3951);
or U5629 (N_5629,N_3465,N_3808);
xnor U5630 (N_5630,N_3237,N_3886);
nand U5631 (N_5631,N_4348,N_3311);
nand U5632 (N_5632,N_3329,N_3803);
nor U5633 (N_5633,N_3816,N_4466);
and U5634 (N_5634,N_3079,N_3750);
or U5635 (N_5635,N_3492,N_3763);
nor U5636 (N_5636,N_3597,N_3500);
or U5637 (N_5637,N_4098,N_4305);
and U5638 (N_5638,N_3476,N_4075);
nor U5639 (N_5639,N_4102,N_3040);
nor U5640 (N_5640,N_3794,N_3399);
or U5641 (N_5641,N_3435,N_4301);
or U5642 (N_5642,N_3954,N_3068);
xnor U5643 (N_5643,N_3646,N_3835);
xnor U5644 (N_5644,N_3346,N_3042);
and U5645 (N_5645,N_3578,N_3570);
and U5646 (N_5646,N_3870,N_3081);
xnor U5647 (N_5647,N_4130,N_3129);
nor U5648 (N_5648,N_3371,N_4363);
or U5649 (N_5649,N_3581,N_3719);
xor U5650 (N_5650,N_4328,N_4280);
and U5651 (N_5651,N_3299,N_3065);
nand U5652 (N_5652,N_3494,N_4460);
or U5653 (N_5653,N_3994,N_4060);
xor U5654 (N_5654,N_3388,N_3651);
nor U5655 (N_5655,N_4215,N_3372);
and U5656 (N_5656,N_4013,N_4186);
or U5657 (N_5657,N_3720,N_3411);
nand U5658 (N_5658,N_3240,N_3795);
xor U5659 (N_5659,N_4470,N_3875);
nor U5660 (N_5660,N_3544,N_3334);
nor U5661 (N_5661,N_3555,N_3286);
nor U5662 (N_5662,N_4014,N_3085);
and U5663 (N_5663,N_3330,N_4267);
nor U5664 (N_5664,N_3861,N_3106);
nand U5665 (N_5665,N_4480,N_3644);
or U5666 (N_5666,N_3074,N_3159);
and U5667 (N_5667,N_3185,N_4067);
or U5668 (N_5668,N_4422,N_4456);
xnor U5669 (N_5669,N_4378,N_3189);
nor U5670 (N_5670,N_3620,N_3925);
and U5671 (N_5671,N_4282,N_3772);
xor U5672 (N_5672,N_3053,N_3788);
nor U5673 (N_5673,N_4396,N_4294);
nor U5674 (N_5674,N_3158,N_4149);
nor U5675 (N_5675,N_4411,N_3409);
and U5676 (N_5676,N_3681,N_4415);
nand U5677 (N_5677,N_3183,N_3844);
or U5678 (N_5678,N_3301,N_3267);
xnor U5679 (N_5679,N_3693,N_3869);
or U5680 (N_5680,N_3856,N_3077);
and U5681 (N_5681,N_4382,N_4420);
and U5682 (N_5682,N_4146,N_4173);
nand U5683 (N_5683,N_4103,N_3342);
and U5684 (N_5684,N_3143,N_4061);
xnor U5685 (N_5685,N_3975,N_4311);
nor U5686 (N_5686,N_3227,N_4113);
and U5687 (N_5687,N_4387,N_4052);
nor U5688 (N_5688,N_3308,N_3859);
or U5689 (N_5689,N_3574,N_4471);
xnor U5690 (N_5690,N_3888,N_3686);
and U5691 (N_5691,N_4287,N_3142);
nor U5692 (N_5692,N_3560,N_3943);
nand U5693 (N_5693,N_3869,N_3569);
xor U5694 (N_5694,N_3204,N_3603);
or U5695 (N_5695,N_3187,N_4440);
nand U5696 (N_5696,N_3563,N_3660);
nand U5697 (N_5697,N_4104,N_3489);
xor U5698 (N_5698,N_3951,N_3138);
and U5699 (N_5699,N_3202,N_3639);
or U5700 (N_5700,N_3066,N_3918);
xor U5701 (N_5701,N_4244,N_3817);
nor U5702 (N_5702,N_4110,N_4280);
xor U5703 (N_5703,N_3391,N_3767);
xor U5704 (N_5704,N_4081,N_3495);
nor U5705 (N_5705,N_3385,N_4466);
nand U5706 (N_5706,N_3390,N_3978);
and U5707 (N_5707,N_3576,N_4424);
nand U5708 (N_5708,N_4022,N_3466);
or U5709 (N_5709,N_4296,N_3708);
or U5710 (N_5710,N_3409,N_4156);
and U5711 (N_5711,N_3444,N_3165);
or U5712 (N_5712,N_3849,N_4295);
or U5713 (N_5713,N_3335,N_3356);
nor U5714 (N_5714,N_3759,N_4350);
or U5715 (N_5715,N_4254,N_3532);
and U5716 (N_5716,N_3812,N_3572);
or U5717 (N_5717,N_4030,N_4294);
or U5718 (N_5718,N_3151,N_4404);
and U5719 (N_5719,N_3534,N_4073);
nor U5720 (N_5720,N_3126,N_3018);
and U5721 (N_5721,N_3724,N_4260);
nand U5722 (N_5722,N_4093,N_3301);
xnor U5723 (N_5723,N_3479,N_4045);
and U5724 (N_5724,N_3597,N_4229);
xnor U5725 (N_5725,N_3338,N_4162);
or U5726 (N_5726,N_3013,N_4068);
nand U5727 (N_5727,N_4342,N_4495);
or U5728 (N_5728,N_3386,N_3941);
xor U5729 (N_5729,N_3578,N_3364);
xnor U5730 (N_5730,N_4224,N_3927);
or U5731 (N_5731,N_4251,N_3743);
nand U5732 (N_5732,N_3904,N_4049);
xnor U5733 (N_5733,N_4380,N_3025);
xnor U5734 (N_5734,N_3616,N_3110);
or U5735 (N_5735,N_3032,N_3905);
or U5736 (N_5736,N_3837,N_3090);
and U5737 (N_5737,N_4315,N_3750);
nand U5738 (N_5738,N_3466,N_3098);
or U5739 (N_5739,N_3868,N_3702);
or U5740 (N_5740,N_4248,N_4320);
nor U5741 (N_5741,N_3491,N_3015);
and U5742 (N_5742,N_4227,N_3132);
or U5743 (N_5743,N_3062,N_3639);
xor U5744 (N_5744,N_4192,N_4367);
or U5745 (N_5745,N_3455,N_3951);
xnor U5746 (N_5746,N_3222,N_3355);
or U5747 (N_5747,N_3496,N_4311);
or U5748 (N_5748,N_4346,N_3082);
xor U5749 (N_5749,N_3369,N_3997);
xnor U5750 (N_5750,N_3976,N_3492);
xor U5751 (N_5751,N_4381,N_3894);
nand U5752 (N_5752,N_4360,N_3510);
xnor U5753 (N_5753,N_3467,N_3910);
nand U5754 (N_5754,N_4401,N_3927);
or U5755 (N_5755,N_4381,N_3895);
xnor U5756 (N_5756,N_3758,N_3922);
and U5757 (N_5757,N_4038,N_3893);
nand U5758 (N_5758,N_4176,N_4182);
nand U5759 (N_5759,N_4381,N_3101);
and U5760 (N_5760,N_4427,N_3063);
nor U5761 (N_5761,N_3097,N_3587);
or U5762 (N_5762,N_3769,N_4331);
and U5763 (N_5763,N_3300,N_3413);
nor U5764 (N_5764,N_4346,N_3524);
nor U5765 (N_5765,N_4436,N_3377);
and U5766 (N_5766,N_3028,N_3236);
nor U5767 (N_5767,N_4296,N_4166);
nor U5768 (N_5768,N_4059,N_3557);
and U5769 (N_5769,N_3203,N_4462);
xnor U5770 (N_5770,N_4112,N_3793);
nor U5771 (N_5771,N_4339,N_3957);
and U5772 (N_5772,N_3945,N_4172);
and U5773 (N_5773,N_4054,N_4179);
and U5774 (N_5774,N_4333,N_3993);
nand U5775 (N_5775,N_3203,N_3467);
xnor U5776 (N_5776,N_3095,N_3384);
and U5777 (N_5777,N_3264,N_3400);
and U5778 (N_5778,N_3386,N_4438);
xor U5779 (N_5779,N_4481,N_3262);
nor U5780 (N_5780,N_4213,N_3819);
nand U5781 (N_5781,N_3534,N_4473);
nor U5782 (N_5782,N_3193,N_3025);
xnor U5783 (N_5783,N_3614,N_3541);
and U5784 (N_5784,N_4339,N_3764);
nand U5785 (N_5785,N_4038,N_4189);
or U5786 (N_5786,N_4466,N_4371);
xor U5787 (N_5787,N_3780,N_3882);
or U5788 (N_5788,N_3256,N_4188);
nor U5789 (N_5789,N_3203,N_3825);
and U5790 (N_5790,N_3781,N_3639);
or U5791 (N_5791,N_3690,N_4484);
nor U5792 (N_5792,N_4251,N_3649);
and U5793 (N_5793,N_3385,N_3615);
nand U5794 (N_5794,N_3771,N_3110);
and U5795 (N_5795,N_3448,N_3965);
or U5796 (N_5796,N_4245,N_3599);
and U5797 (N_5797,N_4445,N_3531);
xnor U5798 (N_5798,N_3996,N_4184);
xnor U5799 (N_5799,N_4400,N_3958);
or U5800 (N_5800,N_3471,N_3653);
or U5801 (N_5801,N_3441,N_3778);
or U5802 (N_5802,N_4227,N_3365);
or U5803 (N_5803,N_4289,N_4449);
or U5804 (N_5804,N_4437,N_4132);
and U5805 (N_5805,N_3677,N_3809);
xnor U5806 (N_5806,N_3834,N_3607);
xor U5807 (N_5807,N_4184,N_3601);
nor U5808 (N_5808,N_4097,N_4067);
xnor U5809 (N_5809,N_4433,N_3047);
xnor U5810 (N_5810,N_4387,N_3963);
nor U5811 (N_5811,N_3719,N_3600);
or U5812 (N_5812,N_3936,N_3556);
or U5813 (N_5813,N_3790,N_3436);
nor U5814 (N_5814,N_3335,N_4198);
xnor U5815 (N_5815,N_3450,N_3561);
and U5816 (N_5816,N_3952,N_3762);
nand U5817 (N_5817,N_3893,N_3883);
and U5818 (N_5818,N_4148,N_3413);
nor U5819 (N_5819,N_3833,N_3765);
nor U5820 (N_5820,N_3496,N_3688);
nor U5821 (N_5821,N_4220,N_3259);
nor U5822 (N_5822,N_3213,N_3053);
and U5823 (N_5823,N_4149,N_4295);
nor U5824 (N_5824,N_4112,N_3613);
and U5825 (N_5825,N_4121,N_3524);
nor U5826 (N_5826,N_4438,N_3234);
nand U5827 (N_5827,N_4235,N_4111);
nand U5828 (N_5828,N_4129,N_3036);
nand U5829 (N_5829,N_3189,N_4289);
nand U5830 (N_5830,N_3676,N_3013);
and U5831 (N_5831,N_3428,N_4002);
and U5832 (N_5832,N_3481,N_4408);
or U5833 (N_5833,N_3947,N_3172);
or U5834 (N_5834,N_3219,N_3461);
and U5835 (N_5835,N_3927,N_3788);
and U5836 (N_5836,N_3508,N_4085);
xnor U5837 (N_5837,N_3217,N_3849);
and U5838 (N_5838,N_3832,N_4495);
nand U5839 (N_5839,N_3518,N_3379);
or U5840 (N_5840,N_3777,N_3655);
nand U5841 (N_5841,N_4060,N_4129);
nand U5842 (N_5842,N_4362,N_3075);
nand U5843 (N_5843,N_3501,N_3184);
xor U5844 (N_5844,N_4153,N_3625);
nor U5845 (N_5845,N_4135,N_3603);
xnor U5846 (N_5846,N_3213,N_4137);
nor U5847 (N_5847,N_4344,N_4010);
and U5848 (N_5848,N_3967,N_4061);
or U5849 (N_5849,N_3446,N_3696);
nor U5850 (N_5850,N_3008,N_4322);
xnor U5851 (N_5851,N_4213,N_4205);
or U5852 (N_5852,N_4036,N_4000);
and U5853 (N_5853,N_4477,N_3109);
nor U5854 (N_5854,N_3621,N_3472);
nor U5855 (N_5855,N_4424,N_3651);
nor U5856 (N_5856,N_4261,N_3931);
xnor U5857 (N_5857,N_3924,N_4443);
or U5858 (N_5858,N_4050,N_3884);
nor U5859 (N_5859,N_4327,N_3402);
or U5860 (N_5860,N_4003,N_4208);
nand U5861 (N_5861,N_3346,N_4470);
nor U5862 (N_5862,N_4253,N_3377);
or U5863 (N_5863,N_4045,N_4445);
nand U5864 (N_5864,N_3222,N_3337);
nor U5865 (N_5865,N_3165,N_4246);
and U5866 (N_5866,N_3156,N_3883);
and U5867 (N_5867,N_4350,N_3785);
xnor U5868 (N_5868,N_3842,N_3861);
and U5869 (N_5869,N_4282,N_4492);
nand U5870 (N_5870,N_4149,N_3310);
nand U5871 (N_5871,N_4230,N_3309);
nor U5872 (N_5872,N_3334,N_3149);
xnor U5873 (N_5873,N_3294,N_3564);
nand U5874 (N_5874,N_4281,N_4149);
nand U5875 (N_5875,N_3339,N_4003);
or U5876 (N_5876,N_3222,N_3500);
nand U5877 (N_5877,N_3273,N_3071);
nand U5878 (N_5878,N_4372,N_3898);
nand U5879 (N_5879,N_3091,N_3042);
or U5880 (N_5880,N_3998,N_3616);
nor U5881 (N_5881,N_3684,N_3798);
and U5882 (N_5882,N_4270,N_3106);
or U5883 (N_5883,N_3704,N_4367);
or U5884 (N_5884,N_3073,N_3187);
and U5885 (N_5885,N_4368,N_3884);
and U5886 (N_5886,N_3205,N_4192);
or U5887 (N_5887,N_3484,N_3490);
nor U5888 (N_5888,N_3795,N_3102);
nor U5889 (N_5889,N_4176,N_4064);
nor U5890 (N_5890,N_4130,N_3118);
nor U5891 (N_5891,N_4317,N_3511);
and U5892 (N_5892,N_3288,N_3628);
and U5893 (N_5893,N_3311,N_3818);
nand U5894 (N_5894,N_4217,N_4021);
or U5895 (N_5895,N_4124,N_3678);
and U5896 (N_5896,N_4255,N_4417);
or U5897 (N_5897,N_4102,N_3103);
and U5898 (N_5898,N_3322,N_4382);
or U5899 (N_5899,N_3053,N_4140);
and U5900 (N_5900,N_3851,N_3779);
xor U5901 (N_5901,N_3323,N_3957);
and U5902 (N_5902,N_4468,N_3990);
nand U5903 (N_5903,N_4026,N_3884);
and U5904 (N_5904,N_3529,N_3834);
or U5905 (N_5905,N_4481,N_3560);
nand U5906 (N_5906,N_4312,N_3650);
or U5907 (N_5907,N_3607,N_4068);
xnor U5908 (N_5908,N_3237,N_4168);
or U5909 (N_5909,N_3038,N_3349);
nor U5910 (N_5910,N_3684,N_3140);
nor U5911 (N_5911,N_3236,N_4251);
or U5912 (N_5912,N_3394,N_4378);
or U5913 (N_5913,N_3217,N_4314);
xnor U5914 (N_5914,N_3433,N_3722);
nand U5915 (N_5915,N_3807,N_4243);
xor U5916 (N_5916,N_4262,N_3175);
nor U5917 (N_5917,N_3808,N_3569);
and U5918 (N_5918,N_3186,N_3406);
or U5919 (N_5919,N_3197,N_3250);
and U5920 (N_5920,N_4087,N_4058);
nand U5921 (N_5921,N_4342,N_3735);
xnor U5922 (N_5922,N_4260,N_3836);
or U5923 (N_5923,N_3801,N_3411);
and U5924 (N_5924,N_3381,N_3343);
xnor U5925 (N_5925,N_4015,N_3266);
and U5926 (N_5926,N_4181,N_4240);
and U5927 (N_5927,N_4069,N_3182);
nand U5928 (N_5928,N_4498,N_4270);
or U5929 (N_5929,N_4492,N_4173);
nand U5930 (N_5930,N_3389,N_3246);
nand U5931 (N_5931,N_3990,N_3577);
nor U5932 (N_5932,N_3522,N_3487);
nor U5933 (N_5933,N_3327,N_4029);
or U5934 (N_5934,N_3721,N_3787);
and U5935 (N_5935,N_3925,N_4306);
nor U5936 (N_5936,N_4353,N_3080);
nor U5937 (N_5937,N_3282,N_3587);
nand U5938 (N_5938,N_3442,N_4231);
nand U5939 (N_5939,N_3877,N_4485);
and U5940 (N_5940,N_3677,N_3747);
nor U5941 (N_5941,N_3763,N_4163);
xor U5942 (N_5942,N_4363,N_4146);
xnor U5943 (N_5943,N_3024,N_3308);
and U5944 (N_5944,N_3883,N_4186);
xor U5945 (N_5945,N_3902,N_3704);
or U5946 (N_5946,N_3297,N_3126);
nor U5947 (N_5947,N_3488,N_4351);
or U5948 (N_5948,N_4266,N_4417);
and U5949 (N_5949,N_3150,N_3861);
xor U5950 (N_5950,N_4164,N_4172);
nand U5951 (N_5951,N_4383,N_3509);
and U5952 (N_5952,N_3638,N_4270);
or U5953 (N_5953,N_3647,N_3471);
nor U5954 (N_5954,N_3317,N_4206);
nand U5955 (N_5955,N_3886,N_3240);
nor U5956 (N_5956,N_3994,N_3604);
nand U5957 (N_5957,N_3456,N_3129);
or U5958 (N_5958,N_3639,N_3743);
and U5959 (N_5959,N_4289,N_4242);
and U5960 (N_5960,N_3271,N_3977);
nand U5961 (N_5961,N_3281,N_3613);
nand U5962 (N_5962,N_3955,N_4470);
and U5963 (N_5963,N_3241,N_3802);
nand U5964 (N_5964,N_3099,N_3873);
nor U5965 (N_5965,N_3513,N_4409);
xor U5966 (N_5966,N_4337,N_3459);
and U5967 (N_5967,N_3887,N_4451);
and U5968 (N_5968,N_3521,N_4188);
nor U5969 (N_5969,N_3515,N_3207);
and U5970 (N_5970,N_3102,N_3535);
xor U5971 (N_5971,N_4213,N_3681);
nor U5972 (N_5972,N_3544,N_4034);
or U5973 (N_5973,N_4011,N_4495);
nand U5974 (N_5974,N_3612,N_3164);
nand U5975 (N_5975,N_3682,N_3880);
xor U5976 (N_5976,N_3621,N_3161);
xnor U5977 (N_5977,N_3226,N_3646);
nand U5978 (N_5978,N_4107,N_3885);
nand U5979 (N_5979,N_4484,N_3389);
or U5980 (N_5980,N_4377,N_3874);
and U5981 (N_5981,N_3137,N_3496);
or U5982 (N_5982,N_3100,N_4035);
xnor U5983 (N_5983,N_3996,N_3310);
and U5984 (N_5984,N_3613,N_4249);
and U5985 (N_5985,N_3580,N_3611);
xnor U5986 (N_5986,N_4075,N_3528);
nand U5987 (N_5987,N_3687,N_3805);
or U5988 (N_5988,N_4274,N_3472);
and U5989 (N_5989,N_4478,N_4100);
and U5990 (N_5990,N_3018,N_3053);
xor U5991 (N_5991,N_4321,N_3396);
nand U5992 (N_5992,N_3572,N_3039);
nand U5993 (N_5993,N_3890,N_4367);
nand U5994 (N_5994,N_3963,N_3294);
and U5995 (N_5995,N_4034,N_4292);
and U5996 (N_5996,N_3733,N_3725);
xor U5997 (N_5997,N_3147,N_3810);
or U5998 (N_5998,N_3376,N_3374);
or U5999 (N_5999,N_4481,N_3996);
nor U6000 (N_6000,N_4688,N_5644);
nand U6001 (N_6001,N_5938,N_5518);
or U6002 (N_6002,N_5930,N_5413);
and U6003 (N_6003,N_4660,N_4837);
or U6004 (N_6004,N_4831,N_4643);
nor U6005 (N_6005,N_4830,N_4926);
xor U6006 (N_6006,N_5609,N_4707);
and U6007 (N_6007,N_5582,N_5179);
xor U6008 (N_6008,N_4961,N_5757);
or U6009 (N_6009,N_5293,N_5982);
nor U6010 (N_6010,N_5633,N_5491);
nor U6011 (N_6011,N_5987,N_4963);
xor U6012 (N_6012,N_4645,N_5035);
and U6013 (N_6013,N_5911,N_5925);
or U6014 (N_6014,N_4572,N_4813);
and U6015 (N_6015,N_5124,N_5102);
xor U6016 (N_6016,N_5089,N_4674);
and U6017 (N_6017,N_5349,N_5027);
xnor U6018 (N_6018,N_5555,N_5683);
nand U6019 (N_6019,N_5343,N_4905);
xor U6020 (N_6020,N_5876,N_5507);
nand U6021 (N_6021,N_5794,N_4852);
and U6022 (N_6022,N_4578,N_5081);
nand U6023 (N_6023,N_4916,N_4618);
nand U6024 (N_6024,N_4894,N_4784);
nor U6025 (N_6025,N_4612,N_5273);
nand U6026 (N_6026,N_5473,N_4842);
nor U6027 (N_6027,N_4622,N_5997);
xnor U6028 (N_6028,N_4540,N_5074);
nand U6029 (N_6029,N_5064,N_4577);
nand U6030 (N_6030,N_4717,N_5317);
xnor U6031 (N_6031,N_4644,N_5178);
and U6032 (N_6032,N_4599,N_4689);
nand U6033 (N_6033,N_5039,N_5013);
or U6034 (N_6034,N_5126,N_5798);
nand U6035 (N_6035,N_4914,N_5923);
nor U6036 (N_6036,N_4747,N_5976);
nor U6037 (N_6037,N_4507,N_5914);
nor U6038 (N_6038,N_4770,N_5988);
or U6039 (N_6039,N_5482,N_4972);
xnor U6040 (N_6040,N_4721,N_5575);
and U6041 (N_6041,N_4866,N_4874);
xor U6042 (N_6042,N_5447,N_5493);
and U6043 (N_6043,N_4878,N_5568);
and U6044 (N_6044,N_4939,N_5395);
nand U6045 (N_6045,N_5990,N_5773);
nor U6046 (N_6046,N_5044,N_5279);
and U6047 (N_6047,N_5772,N_5951);
and U6048 (N_6048,N_5655,N_5407);
nand U6049 (N_6049,N_4898,N_5600);
or U6050 (N_6050,N_5420,N_5656);
nor U6051 (N_6051,N_5402,N_5077);
or U6052 (N_6052,N_4956,N_4918);
and U6053 (N_6053,N_5776,N_4606);
nor U6054 (N_6054,N_4930,N_5836);
or U6055 (N_6055,N_4710,N_5409);
or U6056 (N_6056,N_5549,N_5672);
nor U6057 (N_6057,N_4724,N_5980);
or U6058 (N_6058,N_4949,N_4818);
or U6059 (N_6059,N_4508,N_4774);
and U6060 (N_6060,N_5245,N_5623);
and U6061 (N_6061,N_5536,N_5675);
and U6062 (N_6062,N_5226,N_5524);
nor U6063 (N_6063,N_5437,N_4803);
nor U6064 (N_6064,N_4735,N_5635);
or U6065 (N_6065,N_5770,N_4969);
nor U6066 (N_6066,N_5585,N_5153);
xnor U6067 (N_6067,N_5134,N_5452);
xor U6068 (N_6068,N_5466,N_5517);
or U6069 (N_6069,N_5330,N_5065);
and U6070 (N_6070,N_5168,N_5338);
nor U6071 (N_6071,N_5543,N_4880);
xor U6072 (N_6072,N_4532,N_4863);
or U6073 (N_6073,N_4545,N_5985);
and U6074 (N_6074,N_4822,N_4590);
xor U6075 (N_6075,N_5691,N_5658);
and U6076 (N_6076,N_4619,N_4664);
nand U6077 (N_6077,N_4746,N_4865);
nor U6078 (N_6078,N_5239,N_5526);
xnor U6079 (N_6079,N_4760,N_4742);
nand U6080 (N_6080,N_5753,N_5870);
nand U6081 (N_6081,N_4738,N_5268);
nor U6082 (N_6082,N_5712,N_5458);
xor U6083 (N_6083,N_5598,N_5442);
xor U6084 (N_6084,N_4904,N_5778);
nor U6085 (N_6085,N_5121,N_4889);
or U6086 (N_6086,N_5266,N_5786);
xor U6087 (N_6087,N_5047,N_4858);
and U6088 (N_6088,N_4758,N_4517);
xnor U6089 (N_6089,N_5744,N_5165);
and U6090 (N_6090,N_5640,N_4811);
xor U6091 (N_6091,N_5570,N_5132);
nand U6092 (N_6092,N_4713,N_5058);
or U6093 (N_6093,N_5768,N_4712);
nand U6094 (N_6094,N_5596,N_5328);
nor U6095 (N_6095,N_5784,N_4684);
and U6096 (N_6096,N_5544,N_4555);
and U6097 (N_6097,N_5201,N_5857);
nor U6098 (N_6098,N_5036,N_5125);
or U6099 (N_6099,N_5935,N_5189);
and U6100 (N_6100,N_5759,N_4665);
xnor U6101 (N_6101,N_5022,N_5117);
xnor U6102 (N_6102,N_4902,N_5119);
nand U6103 (N_6103,N_5638,N_5352);
or U6104 (N_6104,N_4616,N_5780);
nor U6105 (N_6105,N_5244,N_5831);
xor U6106 (N_6106,N_4593,N_5503);
nand U6107 (N_6107,N_5200,N_4654);
or U6108 (N_6108,N_4629,N_5823);
xor U6109 (N_6109,N_4698,N_4994);
xnor U6110 (N_6110,N_5916,N_5922);
nand U6111 (N_6111,N_4675,N_5112);
or U6112 (N_6112,N_5385,N_5894);
and U6113 (N_6113,N_5900,N_4788);
or U6114 (N_6114,N_4873,N_4705);
and U6115 (N_6115,N_5885,N_4936);
or U6116 (N_6116,N_5711,N_5299);
nand U6117 (N_6117,N_5969,N_4562);
nor U6118 (N_6118,N_5586,N_5954);
nor U6119 (N_6119,N_4792,N_5705);
xor U6120 (N_6120,N_5869,N_5896);
or U6121 (N_6121,N_4657,N_5043);
xor U6122 (N_6122,N_5158,N_4838);
nand U6123 (N_6123,N_5008,N_4623);
and U6124 (N_6124,N_4631,N_5681);
nor U6125 (N_6125,N_5505,N_4809);
nor U6126 (N_6126,N_5028,N_5700);
xor U6127 (N_6127,N_4607,N_5878);
and U6128 (N_6128,N_5872,N_4666);
nor U6129 (N_6129,N_5030,N_5372);
nor U6130 (N_6130,N_5811,N_5687);
and U6131 (N_6131,N_5141,N_5080);
nand U6132 (N_6132,N_5525,N_4557);
or U6133 (N_6133,N_5004,N_5217);
xor U6134 (N_6134,N_5653,N_5240);
and U6135 (N_6135,N_4649,N_4828);
nor U6136 (N_6136,N_5924,N_5172);
nor U6137 (N_6137,N_5664,N_5157);
nor U6138 (N_6138,N_4598,N_4762);
nand U6139 (N_6139,N_5706,N_5356);
and U6140 (N_6140,N_5803,N_5694);
nand U6141 (N_6141,N_4626,N_5436);
xnor U6142 (N_6142,N_4810,N_4663);
xor U6143 (N_6143,N_5187,N_5715);
and U6144 (N_6144,N_5406,N_5629);
nor U6145 (N_6145,N_4843,N_5854);
nor U6146 (N_6146,N_5079,N_4530);
xnor U6147 (N_6147,N_5825,N_5581);
xnor U6148 (N_6148,N_4648,N_4563);
nor U6149 (N_6149,N_5461,N_5634);
nand U6150 (N_6150,N_4756,N_5136);
nand U6151 (N_6151,N_4832,N_4857);
and U6152 (N_6152,N_5070,N_5417);
and U6153 (N_6153,N_4833,N_4642);
nand U6154 (N_6154,N_5860,N_4806);
nor U6155 (N_6155,N_4846,N_5438);
nor U6156 (N_6156,N_5267,N_4521);
nand U6157 (N_6157,N_4933,N_5408);
nand U6158 (N_6158,N_5843,N_5531);
nor U6159 (N_6159,N_4789,N_4708);
nor U6160 (N_6160,N_5781,N_5054);
nand U6161 (N_6161,N_5650,N_5090);
or U6162 (N_6162,N_4864,N_5465);
xor U6163 (N_6163,N_5326,N_5766);
and U6164 (N_6164,N_4932,N_5237);
or U6165 (N_6165,N_5783,N_5589);
xor U6166 (N_6166,N_4510,N_5289);
xnor U6167 (N_6167,N_5865,N_5208);
or U6168 (N_6168,N_5177,N_5147);
nand U6169 (N_6169,N_4680,N_4552);
or U6170 (N_6170,N_5485,N_5073);
or U6171 (N_6171,N_5820,N_5418);
xnor U6172 (N_6172,N_5845,N_4501);
or U6173 (N_6173,N_4585,N_5416);
xnor U6174 (N_6174,N_4977,N_5796);
xnor U6175 (N_6175,N_5154,N_5419);
nand U6176 (N_6176,N_5309,N_5410);
nand U6177 (N_6177,N_5169,N_4716);
nor U6178 (N_6178,N_5040,N_5238);
xnor U6179 (N_6179,N_5354,N_5731);
nand U6180 (N_6180,N_5383,N_4888);
nor U6181 (N_6181,N_4693,N_4714);
and U6182 (N_6182,N_5921,N_5001);
xnor U6183 (N_6183,N_5632,N_5898);
nor U6184 (N_6184,N_5999,N_5193);
and U6185 (N_6185,N_5445,N_5232);
nor U6186 (N_6186,N_5254,N_4901);
nand U6187 (N_6187,N_5327,N_5184);
xor U6188 (N_6188,N_4951,N_5311);
xor U6189 (N_6189,N_4962,N_5470);
and U6190 (N_6190,N_5053,N_4906);
xnor U6191 (N_6191,N_4536,N_5535);
and U6192 (N_6192,N_4887,N_5649);
nor U6193 (N_6193,N_4668,N_4825);
and U6194 (N_6194,N_5403,N_5093);
xnor U6195 (N_6195,N_5926,N_4610);
nor U6196 (N_6196,N_5790,N_5981);
nor U6197 (N_6197,N_5862,N_4817);
nor U6198 (N_6198,N_5944,N_4958);
xor U6199 (N_6199,N_5821,N_5498);
nand U6200 (N_6200,N_4935,N_5906);
nor U6201 (N_6201,N_5630,N_5603);
or U6202 (N_6202,N_4669,N_4815);
or U6203 (N_6203,N_4730,N_5584);
or U6204 (N_6204,N_5713,N_4537);
xnor U6205 (N_6205,N_4591,N_4635);
and U6206 (N_6206,N_4512,N_4928);
or U6207 (N_6207,N_4927,N_4709);
nand U6208 (N_6208,N_5241,N_5539);
or U6209 (N_6209,N_4736,N_4613);
nand U6210 (N_6210,N_5859,N_5646);
or U6211 (N_6211,N_5204,N_4686);
xor U6212 (N_6212,N_5155,N_5218);
and U6213 (N_6213,N_5903,N_5056);
nand U6214 (N_6214,N_5280,N_5880);
and U6215 (N_6215,N_5974,N_5032);
nor U6216 (N_6216,N_4764,N_5929);
nand U6217 (N_6217,N_5983,N_4611);
or U6218 (N_6218,N_4952,N_4869);
and U6219 (N_6219,N_5627,N_4702);
and U6220 (N_6220,N_4777,N_4920);
and U6221 (N_6221,N_5099,N_4615);
or U6222 (N_6222,N_5977,N_4547);
nor U6223 (N_6223,N_5550,N_4690);
nor U6224 (N_6224,N_5523,N_5449);
nand U6225 (N_6225,N_4847,N_5353);
nor U6226 (N_6226,N_5942,N_4526);
xor U6227 (N_6227,N_4614,N_5451);
xor U6228 (N_6228,N_5874,N_4794);
nand U6229 (N_6229,N_4573,N_5488);
or U6230 (N_6230,N_5384,N_5487);
and U6231 (N_6231,N_4979,N_4795);
nor U6232 (N_6232,N_5486,N_5197);
or U6233 (N_6233,N_5888,N_4890);
or U6234 (N_6234,N_5152,N_5135);
or U6235 (N_6235,N_4621,N_5378);
or U6236 (N_6236,N_4658,N_5243);
nor U6237 (N_6237,N_4672,N_5703);
xor U6238 (N_6238,N_5897,N_5370);
nand U6239 (N_6239,N_5167,N_4995);
nor U6240 (N_6240,N_4604,N_5529);
nand U6241 (N_6241,N_5214,N_4625);
xnor U6242 (N_6242,N_5733,N_5839);
nor U6243 (N_6243,N_4681,N_4543);
xor U6244 (N_6244,N_4551,N_5499);
and U6245 (N_6245,N_4715,N_4500);
nor U6246 (N_6246,N_4694,N_5918);
nand U6247 (N_6247,N_4872,N_5717);
xor U6248 (N_6248,N_5986,N_4923);
and U6249 (N_6249,N_5213,N_4749);
and U6250 (N_6250,N_4778,N_5611);
xor U6251 (N_6251,N_5024,N_5509);
and U6252 (N_6252,N_5334,N_5957);
xnor U6253 (N_6253,N_5714,N_5963);
or U6254 (N_6254,N_5615,N_5034);
nand U6255 (N_6255,N_4983,N_5490);
or U6256 (N_6256,N_4656,N_4617);
nor U6257 (N_6257,N_5263,N_4785);
or U6258 (N_6258,N_5676,N_5910);
or U6259 (N_6259,N_4542,N_5802);
or U6260 (N_6260,N_4691,N_5062);
xor U6261 (N_6261,N_4791,N_4881);
and U6262 (N_6262,N_5367,N_5984);
and U6263 (N_6263,N_5745,N_4876);
nor U6264 (N_6264,N_5399,N_5212);
nand U6265 (N_6265,N_5883,N_4950);
nor U6266 (N_6266,N_5852,N_5091);
or U6267 (N_6267,N_5005,N_4516);
nor U6268 (N_6268,N_5521,N_5247);
nand U6269 (N_6269,N_4525,N_5002);
nand U6270 (N_6270,N_5194,N_5667);
nand U6271 (N_6271,N_5592,N_5527);
nand U6272 (N_6272,N_4883,N_5350);
or U6273 (N_6273,N_5561,N_5173);
xnor U6274 (N_6274,N_5665,N_5608);
xnor U6275 (N_6275,N_5978,N_5789);
nand U6276 (N_6276,N_4862,N_5949);
nor U6277 (N_6277,N_5631,N_5701);
xnor U6278 (N_6278,N_5313,N_4720);
or U6279 (N_6279,N_4560,N_4588);
xor U6280 (N_6280,N_4974,N_5068);
or U6281 (N_6281,N_4759,N_5552);
xnor U6282 (N_6282,N_4761,N_5729);
nor U6283 (N_6283,N_5782,N_5434);
and U6284 (N_6284,N_5994,N_5995);
nand U6285 (N_6285,N_5260,N_4799);
or U6286 (N_6286,N_4984,N_5016);
nor U6287 (N_6287,N_5373,N_5542);
nand U6288 (N_6288,N_4841,N_5248);
nor U6289 (N_6289,N_5702,N_5257);
or U6290 (N_6290,N_5743,N_5967);
and U6291 (N_6291,N_5899,N_4955);
xor U6292 (N_6292,N_4741,N_4909);
and U6293 (N_6293,N_5730,N_5159);
and U6294 (N_6294,N_5433,N_5962);
nand U6295 (N_6295,N_5432,N_4780);
and U6296 (N_6296,N_5021,N_5606);
nor U6297 (N_6297,N_5306,N_5310);
nor U6298 (N_6298,N_5139,N_5365);
or U6299 (N_6299,N_5774,N_5775);
or U6300 (N_6300,N_4937,N_5483);
nand U6301 (N_6301,N_5685,N_5075);
nand U6302 (N_6302,N_4524,N_4587);
nor U6303 (N_6303,N_4548,N_5826);
nor U6304 (N_6304,N_5163,N_5689);
or U6305 (N_6305,N_5915,N_5278);
nand U6306 (N_6306,N_5363,N_5613);
nor U6307 (N_6307,N_4790,N_5619);
nand U6308 (N_6308,N_4699,N_5140);
or U6309 (N_6309,N_5858,N_5863);
nand U6310 (N_6310,N_5097,N_5810);
xor U6311 (N_6311,N_5332,N_5873);
and U6312 (N_6312,N_5292,N_5610);
nand U6313 (N_6313,N_5959,N_4752);
nand U6314 (N_6314,N_5738,N_5283);
xor U6315 (N_6315,N_4734,N_5264);
nor U6316 (N_6316,N_5941,N_4965);
or U6317 (N_6317,N_5128,N_5249);
or U6318 (N_6318,N_5726,N_5622);
xor U6319 (N_6319,N_5103,N_5000);
xor U6320 (N_6320,N_4827,N_5377);
nand U6321 (N_6321,N_4739,N_4620);
nand U6322 (N_6322,N_5566,N_5513);
nand U6323 (N_6323,N_5386,N_5428);
xnor U6324 (N_6324,N_4719,N_5031);
and U6325 (N_6325,N_5955,N_5236);
nor U6326 (N_6326,N_4533,N_4772);
and U6327 (N_6327,N_5892,N_5844);
nand U6328 (N_6328,N_5666,N_5797);
or U6329 (N_6329,N_5697,N_5092);
and U6330 (N_6330,N_5932,N_5651);
and U6331 (N_6331,N_4670,N_4849);
or U6332 (N_6332,N_4556,N_5115);
xor U6333 (N_6333,N_5716,N_4594);
nor U6334 (N_6334,N_5720,N_5206);
nor U6335 (N_6335,N_5602,N_5749);
or U6336 (N_6336,N_5252,N_5939);
or U6337 (N_6337,N_4892,N_4966);
nor U6338 (N_6338,N_5752,N_5459);
xor U6339 (N_6339,N_5818,N_5756);
and U6340 (N_6340,N_5851,N_5884);
nand U6341 (N_6341,N_5946,N_4743);
nand U6342 (N_6342,N_5286,N_4934);
xnor U6343 (N_6343,N_4677,N_5992);
nand U6344 (N_6344,N_4605,N_5813);
xnor U6345 (N_6345,N_5095,N_5788);
xnor U6346 (N_6346,N_4652,N_4659);
xor U6347 (N_6347,N_5078,N_4988);
or U6348 (N_6348,N_4704,N_5736);
and U6349 (N_6349,N_5430,N_5072);
and U6350 (N_6350,N_5828,N_5979);
and U6351 (N_6351,N_4655,N_5989);
nor U6352 (N_6352,N_5412,N_4978);
or U6353 (N_6353,N_5175,N_5253);
nand U6354 (N_6354,N_5284,N_4509);
or U6355 (N_6355,N_5440,N_5366);
or U6356 (N_6356,N_5323,N_4519);
nor U6357 (N_6357,N_4816,N_5038);
nor U6358 (N_6358,N_5389,N_5699);
and U6359 (N_6359,N_5719,N_5545);
and U6360 (N_6360,N_5934,N_5133);
or U6361 (N_6361,N_4506,N_4859);
nand U6362 (N_6362,N_4941,N_5364);
and U6363 (N_6363,N_5255,N_5494);
and U6364 (N_6364,N_4513,N_4630);
and U6365 (N_6365,N_5497,N_4824);
and U6366 (N_6366,N_5500,N_5960);
xor U6367 (N_6367,N_5620,N_4581);
and U6368 (N_6368,N_5741,N_5710);
nor U6369 (N_6369,N_5554,N_5421);
nand U6370 (N_6370,N_5607,N_4940);
xnor U6371 (N_6371,N_5708,N_5496);
nand U6372 (N_6372,N_4718,N_5120);
nand U6373 (N_6373,N_5131,N_4678);
xor U6374 (N_6374,N_4993,N_5342);
nand U6375 (N_6375,N_4679,N_5693);
nor U6376 (N_6376,N_4997,N_5130);
and U6377 (N_6377,N_5742,N_5006);
nand U6378 (N_6378,N_4751,N_4579);
nand U6379 (N_6379,N_5576,N_5562);
nand U6380 (N_6380,N_5269,N_5740);
or U6381 (N_6381,N_5947,N_4753);
xnor U6382 (N_6382,N_5076,N_5164);
nand U6383 (N_6383,N_5577,N_4600);
xnor U6384 (N_6384,N_5871,N_4685);
nand U6385 (N_6385,N_4797,N_5297);
nand U6386 (N_6386,N_5265,N_5840);
or U6387 (N_6387,N_5642,N_4755);
and U6388 (N_6388,N_5591,N_4885);
or U6389 (N_6389,N_5762,N_5456);
or U6390 (N_6390,N_5795,N_4697);
nor U6391 (N_6391,N_5645,N_5750);
xnor U6392 (N_6392,N_5282,N_5014);
xnor U6393 (N_6393,N_5541,N_5042);
or U6394 (N_6394,N_4504,N_5231);
nand U6395 (N_6395,N_5015,N_5948);
xor U6396 (N_6396,N_5382,N_5515);
or U6397 (N_6397,N_5037,N_4948);
or U6398 (N_6398,N_5170,N_5067);
nor U6399 (N_6399,N_5537,N_5732);
or U6400 (N_6400,N_5877,N_5060);
nand U6401 (N_6401,N_5300,N_4529);
and U6402 (N_6402,N_5387,N_5495);
nand U6403 (N_6403,N_5636,N_5288);
or U6404 (N_6404,N_5106,N_5492);
and U6405 (N_6405,N_5104,N_5302);
nor U6406 (N_6406,N_4583,N_4706);
nor U6407 (N_6407,N_5808,N_5684);
and U6408 (N_6408,N_4938,N_4973);
and U6409 (N_6409,N_5052,N_5142);
nand U6410 (N_6410,N_4682,N_5023);
and U6411 (N_6411,N_4919,N_5472);
or U6412 (N_6412,N_5180,N_5936);
nand U6413 (N_6413,N_5891,N_4999);
xnor U6414 (N_6414,N_5435,N_5734);
or U6415 (N_6415,N_4535,N_5567);
and U6416 (N_6416,N_5850,N_4725);
and U6417 (N_6417,N_5540,N_5837);
and U6418 (N_6418,N_5025,N_5118);
or U6419 (N_6419,N_5320,N_4609);
or U6420 (N_6420,N_4737,N_4592);
nand U6421 (N_6421,N_4515,N_5322);
nand U6422 (N_6422,N_5340,N_5071);
xor U6423 (N_6423,N_5970,N_5307);
nor U6424 (N_6424,N_5392,N_4754);
nor U6425 (N_6425,N_4886,N_5626);
nor U6426 (N_6426,N_4564,N_5325);
and U6427 (N_6427,N_5422,N_5534);
and U6428 (N_6428,N_4954,N_5904);
xnor U6429 (N_6429,N_5361,N_5893);
nor U6430 (N_6430,N_5057,N_5186);
or U6431 (N_6431,N_5595,N_4653);
nor U6432 (N_6432,N_5415,N_4602);
xor U6433 (N_6433,N_4893,N_5725);
xnor U6434 (N_6434,N_4757,N_4808);
and U6435 (N_6435,N_5460,N_4823);
nand U6436 (N_6436,N_5920,N_4836);
and U6437 (N_6437,N_5376,N_5573);
or U6438 (N_6438,N_5151,N_4854);
nand U6439 (N_6439,N_5108,N_5815);
xnor U6440 (N_6440,N_4596,N_5824);
or U6441 (N_6441,N_5051,N_5546);
xor U6442 (N_6442,N_5565,N_5202);
nor U6443 (N_6443,N_5329,N_5116);
nand U6444 (N_6444,N_5617,N_5448);
or U6445 (N_6445,N_5569,N_4646);
nor U6446 (N_6446,N_4917,N_5879);
or U6447 (N_6447,N_5431,N_4981);
nor U6448 (N_6448,N_5258,N_5398);
nand U6449 (N_6449,N_5659,N_5150);
or U6450 (N_6450,N_5271,N_5479);
nand U6451 (N_6451,N_5624,N_5114);
nand U6452 (N_6452,N_5477,N_4687);
xor U6453 (N_6453,N_4899,N_4576);
nor U6454 (N_6454,N_4727,N_5933);
nand U6455 (N_6455,N_5522,N_4821);
nor U6456 (N_6456,N_5246,N_4511);
nand U6457 (N_6457,N_5662,N_5059);
xnor U6458 (N_6458,N_4527,N_5557);
nand U6459 (N_6459,N_4913,N_5663);
nor U6460 (N_6460,N_5512,N_5274);
nor U6461 (N_6461,N_5272,N_5853);
xor U6462 (N_6462,N_5604,N_4539);
xnor U6463 (N_6463,N_4903,N_5145);
or U6464 (N_6464,N_5511,N_4990);
xor U6465 (N_6465,N_5501,N_5599);
xor U6466 (N_6466,N_5358,N_5087);
xnor U6467 (N_6467,N_4518,N_5270);
or U6468 (N_6468,N_4647,N_5069);
nand U6469 (N_6469,N_5760,N_5261);
or U6470 (N_6470,N_5553,N_5318);
nor U6471 (N_6471,N_5704,N_4884);
and U6472 (N_6472,N_4701,N_5380);
nand U6473 (N_6473,N_4769,N_4840);
or U6474 (N_6474,N_4776,N_4733);
or U6475 (N_6475,N_5209,N_5185);
and U6476 (N_6476,N_4731,N_5160);
and U6477 (N_6477,N_5799,N_4975);
xnor U6478 (N_6478,N_5901,N_5441);
xor U6479 (N_6479,N_5026,N_5695);
and U6480 (N_6480,N_4553,N_5673);
and U6481 (N_6481,N_4546,N_5429);
or U6482 (N_6482,N_5597,N_5199);
and U6483 (N_6483,N_5680,N_4798);
xor U6484 (N_6484,N_4877,N_4566);
nor U6485 (N_6485,N_5453,N_5203);
or U6486 (N_6486,N_5425,N_4985);
and U6487 (N_6487,N_5314,N_4744);
nand U6488 (N_6488,N_5834,N_4853);
or U6489 (N_6489,N_4986,N_5003);
nor U6490 (N_6490,N_5688,N_5785);
xor U6491 (N_6491,N_5198,N_5801);
nor U6492 (N_6492,N_5777,N_5110);
nor U6493 (N_6493,N_5192,N_4711);
xnor U6494 (N_6494,N_5285,N_5812);
or U6495 (N_6495,N_5393,N_5183);
nand U6496 (N_6496,N_5471,N_4775);
nor U6497 (N_6497,N_5887,N_5748);
xor U6498 (N_6498,N_5296,N_4700);
and U6499 (N_6499,N_5864,N_4584);
xnor U6500 (N_6500,N_5331,N_5519);
nand U6501 (N_6501,N_5643,N_5414);
or U6502 (N_6502,N_4971,N_5912);
nand U6503 (N_6503,N_4912,N_5207);
xor U6504 (N_6504,N_5833,N_4550);
nand U6505 (N_6505,N_4559,N_5648);
nand U6506 (N_6506,N_5463,N_5682);
xor U6507 (N_6507,N_5009,N_5560);
or U6508 (N_6508,N_4860,N_4871);
nor U6509 (N_6509,N_5335,N_4554);
nand U6510 (N_6510,N_4748,N_5138);
nand U6511 (N_6511,N_5469,N_5669);
nor U6512 (N_6512,N_5765,N_4793);
nand U6513 (N_6513,N_5590,N_5661);
and U6514 (N_6514,N_5162,N_5621);
xnor U6515 (N_6515,N_5275,N_5109);
and U6516 (N_6516,N_5055,N_5333);
xnor U6517 (N_6517,N_4632,N_4915);
nor U6518 (N_6518,N_5234,N_5787);
and U6519 (N_6519,N_5290,N_5146);
nand U6520 (N_6520,N_5294,N_5861);
nor U6521 (N_6521,N_5909,N_4947);
or U6522 (N_6522,N_4967,N_5446);
xnor U6523 (N_6523,N_4503,N_5084);
or U6524 (N_6524,N_5305,N_5769);
or U6525 (N_6525,N_5019,N_5895);
nand U6526 (N_6526,N_5122,N_4633);
xor U6527 (N_6527,N_5250,N_4726);
nor U6528 (N_6528,N_5262,N_5029);
nand U6529 (N_6529,N_5144,N_5698);
xnor U6530 (N_6530,N_5228,N_5578);
nand U6531 (N_6531,N_5639,N_4851);
nand U6532 (N_6532,N_4641,N_4570);
nand U6533 (N_6533,N_5601,N_5652);
and U6534 (N_6534,N_5816,N_4834);
nand U6535 (N_6535,N_4544,N_5875);
nor U6536 (N_6536,N_4960,N_4597);
nor U6537 (N_6537,N_4637,N_5847);
and U6538 (N_6538,N_5913,N_5316);
nor U6539 (N_6539,N_5945,N_4944);
or U6540 (N_6540,N_4931,N_5657);
or U6541 (N_6541,N_4505,N_5975);
and U6542 (N_6542,N_4812,N_5242);
nand U6543 (N_6543,N_5641,N_5276);
or U6544 (N_6544,N_5190,N_5829);
and U6545 (N_6545,N_5754,N_4768);
nor U6546 (N_6546,N_4745,N_5443);
nor U6547 (N_6547,N_5722,N_5502);
or U6548 (N_6548,N_5007,N_4541);
xnor U6549 (N_6549,N_5220,N_5692);
and U6550 (N_6550,N_4534,N_5618);
and U6551 (N_6551,N_5830,N_4856);
xor U6552 (N_6552,N_5908,N_5508);
nor U6553 (N_6553,N_4946,N_4959);
and U6554 (N_6554,N_5961,N_5807);
or U6555 (N_6555,N_4844,N_5547);
or U6556 (N_6556,N_5956,N_5312);
nand U6557 (N_6557,N_5571,N_5761);
and U6558 (N_6558,N_4839,N_5674);
nand U6559 (N_6559,N_5747,N_5971);
and U6560 (N_6560,N_5222,N_4636);
and U6561 (N_6561,N_4805,N_5806);
or U6562 (N_6562,N_4703,N_4662);
or U6563 (N_6563,N_4855,N_5308);
and U6564 (N_6564,N_5690,N_5696);
and U6565 (N_6565,N_5149,N_4814);
nor U6566 (N_6566,N_5235,N_4565);
or U6567 (N_6567,N_5574,N_5324);
and U6568 (N_6568,N_5259,N_5181);
and U6569 (N_6569,N_5045,N_5551);
nor U6570 (N_6570,N_5127,N_4502);
or U6571 (N_6571,N_4942,N_5588);
xnor U6572 (N_6572,N_5346,N_5856);
nor U6573 (N_6573,N_5905,N_5176);
xnor U6574 (N_6574,N_5475,N_4921);
and U6575 (N_6575,N_5396,N_5593);
nor U6576 (N_6576,N_4729,N_5968);
or U6577 (N_6577,N_4875,N_5137);
nand U6578 (N_6578,N_5063,N_5902);
nand U6579 (N_6579,N_5506,N_5998);
nor U6580 (N_6580,N_4651,N_5866);
and U6581 (N_6581,N_4867,N_4771);
nand U6582 (N_6582,N_5937,N_5041);
nand U6583 (N_6583,N_4671,N_4987);
nand U6584 (N_6584,N_5129,N_5504);
or U6585 (N_6585,N_5457,N_4523);
xnor U6586 (N_6586,N_5362,N_5085);
or U6587 (N_6587,N_4896,N_5791);
xor U6588 (N_6588,N_4826,N_5670);
and U6589 (N_6589,N_4695,N_5048);
xnor U6590 (N_6590,N_4861,N_4807);
or U6591 (N_6591,N_5819,N_5476);
and U6592 (N_6592,N_5855,N_5654);
xor U6593 (N_6593,N_4845,N_4582);
xnor U6594 (N_6594,N_5890,N_5625);
nor U6595 (N_6595,N_5427,N_5345);
nor U6596 (N_6596,N_4879,N_4786);
xnor U6597 (N_6597,N_4945,N_4908);
xor U6598 (N_6598,N_4802,N_5718);
nand U6599 (N_6599,N_5277,N_5224);
or U6600 (N_6600,N_4829,N_5677);
and U6601 (N_6601,N_5668,N_5298);
and U6602 (N_6602,N_5919,N_5215);
or U6603 (N_6603,N_5728,N_5143);
or U6604 (N_6604,N_5304,N_5375);
nand U6605 (N_6605,N_5814,N_5156);
nor U6606 (N_6606,N_4531,N_5287);
nand U6607 (N_6607,N_4634,N_4589);
nand U6608 (N_6608,N_5341,N_5724);
nor U6609 (N_6609,N_4766,N_5404);
nor U6610 (N_6610,N_5931,N_5763);
nor U6611 (N_6611,N_4989,N_5755);
or U6612 (N_6612,N_5017,N_5779);
or U6613 (N_6613,N_5940,N_5827);
or U6614 (N_6614,N_4891,N_4801);
and U6615 (N_6615,N_5405,N_4796);
and U6616 (N_6616,N_4895,N_5559);
nand U6617 (N_6617,N_5484,N_5671);
nand U6618 (N_6618,N_5281,N_4996);
nor U6619 (N_6619,N_4650,N_4957);
or U6620 (N_6620,N_5478,N_4640);
xnor U6621 (N_6621,N_4992,N_5583);
xor U6622 (N_6622,N_5454,N_5809);
and U6623 (N_6623,N_5793,N_5612);
nor U6624 (N_6624,N_5301,N_5587);
nand U6625 (N_6625,N_5223,N_5804);
xor U6626 (N_6626,N_5368,N_5303);
nor U6627 (N_6627,N_5556,N_4568);
xnor U6628 (N_6628,N_5792,N_4538);
nand U6629 (N_6629,N_5061,N_4558);
xor U6630 (N_6630,N_4820,N_4740);
xor U6631 (N_6631,N_5737,N_5291);
nand U6632 (N_6632,N_4953,N_4767);
and U6633 (N_6633,N_5450,N_4522);
xor U6634 (N_6634,N_4528,N_5917);
and U6635 (N_6635,N_5161,N_4980);
and U6636 (N_6636,N_5123,N_5391);
or U6637 (N_6637,N_4929,N_4897);
nor U6638 (N_6638,N_5211,N_5082);
xnor U6639 (N_6639,N_5889,N_5735);
nand U6640 (N_6640,N_4514,N_4787);
nand U6641 (N_6641,N_5538,N_4603);
xnor U6642 (N_6642,N_5171,N_5191);
xor U6643 (N_6643,N_5390,N_5467);
nand U6644 (N_6644,N_5174,N_4943);
and U6645 (N_6645,N_5727,N_5229);
xnor U6646 (N_6646,N_5105,N_5489);
or U6647 (N_6647,N_5835,N_5401);
xnor U6648 (N_6648,N_5397,N_5336);
or U6649 (N_6649,N_4569,N_5337);
xnor U6650 (N_6650,N_4661,N_4922);
and U6651 (N_6651,N_5528,N_5532);
and U6652 (N_6652,N_4765,N_4924);
nand U6653 (N_6653,N_4763,N_5344);
or U6654 (N_6654,N_5033,N_4870);
and U6655 (N_6655,N_5679,N_5010);
nand U6656 (N_6656,N_4722,N_4673);
nand U6657 (N_6657,N_5066,N_5950);
nor U6658 (N_6658,N_4571,N_5548);
nand U6659 (N_6659,N_5958,N_5339);
xor U6660 (N_6660,N_4750,N_5094);
and U6661 (N_6661,N_5832,N_4964);
xnor U6662 (N_6662,N_5012,N_5849);
xor U6663 (N_6663,N_5817,N_5295);
nand U6664 (N_6664,N_4998,N_5096);
and U6665 (N_6665,N_4835,N_5928);
or U6666 (N_6666,N_5707,N_5357);
xnor U6667 (N_6667,N_5347,N_5468);
nor U6668 (N_6668,N_5227,N_5379);
nand U6669 (N_6669,N_4628,N_5088);
nor U6670 (N_6670,N_5927,N_4638);
or U6671 (N_6671,N_4732,N_5886);
nand U6672 (N_6672,N_5480,N_4800);
nor U6673 (N_6673,N_5965,N_4925);
and U6674 (N_6674,N_5216,N_5319);
xor U6675 (N_6675,N_5558,N_5083);
and U6676 (N_6676,N_5315,N_5256);
xnor U6677 (N_6677,N_4520,N_5423);
or U6678 (N_6678,N_5846,N_5520);
and U6679 (N_6679,N_5050,N_5374);
xnor U6680 (N_6680,N_5359,N_5182);
nand U6681 (N_6681,N_4911,N_5481);
and U6682 (N_6682,N_5907,N_5210);
and U6683 (N_6683,N_4848,N_5251);
nor U6684 (N_6684,N_5221,N_4601);
and U6685 (N_6685,N_4882,N_5101);
or U6686 (N_6686,N_5767,N_5952);
or U6687 (N_6687,N_5046,N_4608);
nor U6688 (N_6688,N_4549,N_5205);
and U6689 (N_6689,N_5868,N_5426);
xnor U6690 (N_6690,N_5972,N_5321);
nand U6691 (N_6691,N_5219,N_4595);
nor U6692 (N_6692,N_5424,N_4676);
and U6693 (N_6693,N_5616,N_4779);
xnor U6694 (N_6694,N_5230,N_5739);
nor U6695 (N_6695,N_4819,N_4868);
or U6696 (N_6696,N_5758,N_4683);
xor U6697 (N_6697,N_5351,N_4627);
or U6698 (N_6698,N_5464,N_5533);
or U6699 (N_6699,N_5993,N_5678);
and U6700 (N_6700,N_4982,N_5381);
xor U6701 (N_6701,N_5966,N_5225);
xnor U6702 (N_6702,N_5563,N_5660);
nand U6703 (N_6703,N_5822,N_4907);
or U6704 (N_6704,N_4804,N_4728);
xor U6705 (N_6705,N_4580,N_5751);
nor U6706 (N_6706,N_4781,N_5113);
and U6707 (N_6707,N_5510,N_5020);
and U6708 (N_6708,N_5746,N_4976);
or U6709 (N_6709,N_5514,N_5516);
nand U6710 (N_6710,N_4574,N_5018);
or U6711 (N_6711,N_5098,N_4567);
xor U6712 (N_6712,N_5107,N_5086);
xnor U6713 (N_6713,N_5195,N_5444);
xnor U6714 (N_6714,N_5647,N_5388);
nand U6715 (N_6715,N_4667,N_4639);
or U6716 (N_6716,N_5842,N_5964);
nand U6717 (N_6717,N_5764,N_4561);
nor U6718 (N_6718,N_5530,N_5572);
and U6719 (N_6719,N_5881,N_5411);
nand U6720 (N_6720,N_5369,N_5233);
nor U6721 (N_6721,N_5841,N_5867);
nand U6722 (N_6722,N_5943,N_5614);
nand U6723 (N_6723,N_4900,N_4696);
nor U6724 (N_6724,N_4723,N_4586);
and U6725 (N_6725,N_5100,N_4991);
nand U6726 (N_6726,N_4575,N_4692);
and U6727 (N_6727,N_5049,N_5011);
xnor U6728 (N_6728,N_5709,N_5474);
nand U6729 (N_6729,N_5594,N_4968);
nand U6730 (N_6730,N_4624,N_4773);
and U6731 (N_6731,N_4782,N_5188);
xor U6732 (N_6732,N_5721,N_5148);
nand U6733 (N_6733,N_5991,N_5196);
nor U6734 (N_6734,N_5371,N_4850);
or U6735 (N_6735,N_5723,N_5360);
xor U6736 (N_6736,N_5637,N_5605);
nor U6737 (N_6737,N_4970,N_5686);
xnor U6738 (N_6738,N_5771,N_5580);
nand U6739 (N_6739,N_5348,N_5628);
nor U6740 (N_6740,N_5996,N_5455);
nand U6741 (N_6741,N_5805,N_5953);
or U6742 (N_6742,N_5579,N_5400);
or U6743 (N_6743,N_5838,N_4910);
nor U6744 (N_6744,N_5848,N_5800);
xnor U6745 (N_6745,N_5355,N_4783);
nor U6746 (N_6746,N_5439,N_5564);
nand U6747 (N_6747,N_5394,N_5111);
or U6748 (N_6748,N_5166,N_5462);
or U6749 (N_6749,N_5882,N_5973);
or U6750 (N_6750,N_5497,N_5492);
nor U6751 (N_6751,N_5821,N_5017);
nor U6752 (N_6752,N_4961,N_5013);
nor U6753 (N_6753,N_5611,N_4856);
nor U6754 (N_6754,N_5604,N_5961);
or U6755 (N_6755,N_5843,N_4882);
xor U6756 (N_6756,N_5073,N_5759);
nand U6757 (N_6757,N_5387,N_5793);
nor U6758 (N_6758,N_5736,N_5442);
and U6759 (N_6759,N_5259,N_5228);
nor U6760 (N_6760,N_5136,N_5788);
or U6761 (N_6761,N_5290,N_4695);
nand U6762 (N_6762,N_5188,N_4756);
or U6763 (N_6763,N_5844,N_5504);
xnor U6764 (N_6764,N_4579,N_4629);
xor U6765 (N_6765,N_5467,N_4642);
nand U6766 (N_6766,N_5880,N_5024);
xnor U6767 (N_6767,N_5581,N_4588);
and U6768 (N_6768,N_4995,N_4944);
xor U6769 (N_6769,N_5460,N_5937);
xnor U6770 (N_6770,N_5774,N_5503);
or U6771 (N_6771,N_5314,N_4534);
nor U6772 (N_6772,N_5886,N_4786);
xor U6773 (N_6773,N_5632,N_4962);
and U6774 (N_6774,N_4630,N_5781);
xor U6775 (N_6775,N_5982,N_5064);
or U6776 (N_6776,N_4656,N_5749);
or U6777 (N_6777,N_5434,N_4644);
or U6778 (N_6778,N_5803,N_5588);
nor U6779 (N_6779,N_5895,N_5213);
and U6780 (N_6780,N_5977,N_4891);
or U6781 (N_6781,N_4832,N_5961);
or U6782 (N_6782,N_5468,N_5939);
or U6783 (N_6783,N_4529,N_4725);
xor U6784 (N_6784,N_5942,N_5671);
xnor U6785 (N_6785,N_4917,N_4972);
nand U6786 (N_6786,N_5074,N_5694);
and U6787 (N_6787,N_4976,N_4555);
xor U6788 (N_6788,N_5430,N_5664);
and U6789 (N_6789,N_5335,N_5691);
xnor U6790 (N_6790,N_5492,N_5817);
xor U6791 (N_6791,N_5623,N_5880);
or U6792 (N_6792,N_4583,N_5822);
nor U6793 (N_6793,N_5905,N_4647);
nor U6794 (N_6794,N_4623,N_5846);
or U6795 (N_6795,N_5910,N_5050);
nor U6796 (N_6796,N_5152,N_5966);
nor U6797 (N_6797,N_5494,N_4701);
nand U6798 (N_6798,N_5367,N_5799);
nor U6799 (N_6799,N_5049,N_4965);
or U6800 (N_6800,N_5911,N_5000);
and U6801 (N_6801,N_5322,N_4616);
or U6802 (N_6802,N_4881,N_5009);
or U6803 (N_6803,N_5322,N_4830);
or U6804 (N_6804,N_5619,N_5455);
and U6805 (N_6805,N_5480,N_5401);
and U6806 (N_6806,N_5488,N_4608);
and U6807 (N_6807,N_5989,N_4932);
and U6808 (N_6808,N_5890,N_5756);
and U6809 (N_6809,N_5528,N_5123);
or U6810 (N_6810,N_4771,N_5653);
or U6811 (N_6811,N_5990,N_5784);
or U6812 (N_6812,N_4684,N_5356);
or U6813 (N_6813,N_5250,N_5331);
nand U6814 (N_6814,N_5413,N_5693);
nand U6815 (N_6815,N_4569,N_4513);
or U6816 (N_6816,N_5256,N_5262);
or U6817 (N_6817,N_4622,N_5134);
nand U6818 (N_6818,N_5840,N_4827);
nand U6819 (N_6819,N_5770,N_5420);
and U6820 (N_6820,N_5094,N_5432);
nand U6821 (N_6821,N_5238,N_4861);
nand U6822 (N_6822,N_5633,N_4739);
nand U6823 (N_6823,N_4626,N_5467);
nand U6824 (N_6824,N_5734,N_5155);
and U6825 (N_6825,N_5039,N_4855);
or U6826 (N_6826,N_4640,N_5122);
nor U6827 (N_6827,N_5000,N_4707);
nand U6828 (N_6828,N_5436,N_5615);
nor U6829 (N_6829,N_5666,N_4793);
nand U6830 (N_6830,N_5928,N_4581);
or U6831 (N_6831,N_5348,N_5723);
nand U6832 (N_6832,N_5338,N_4636);
and U6833 (N_6833,N_5794,N_5839);
nand U6834 (N_6834,N_5457,N_4650);
or U6835 (N_6835,N_5835,N_5048);
and U6836 (N_6836,N_5993,N_5588);
xor U6837 (N_6837,N_5096,N_4982);
nor U6838 (N_6838,N_4679,N_5510);
xor U6839 (N_6839,N_5392,N_5264);
and U6840 (N_6840,N_5672,N_4517);
or U6841 (N_6841,N_5988,N_4568);
or U6842 (N_6842,N_5650,N_4562);
xnor U6843 (N_6843,N_5593,N_4735);
and U6844 (N_6844,N_4880,N_5076);
nand U6845 (N_6845,N_5127,N_5938);
nand U6846 (N_6846,N_4613,N_5086);
or U6847 (N_6847,N_4590,N_4974);
nand U6848 (N_6848,N_4939,N_4521);
and U6849 (N_6849,N_5918,N_5997);
or U6850 (N_6850,N_5056,N_4556);
nor U6851 (N_6851,N_5396,N_4520);
xor U6852 (N_6852,N_4998,N_5134);
and U6853 (N_6853,N_4616,N_5306);
xnor U6854 (N_6854,N_5574,N_5025);
xor U6855 (N_6855,N_5426,N_4532);
or U6856 (N_6856,N_5043,N_5028);
nor U6857 (N_6857,N_5222,N_4971);
nand U6858 (N_6858,N_4964,N_4878);
nor U6859 (N_6859,N_5887,N_4619);
and U6860 (N_6860,N_5810,N_5866);
nor U6861 (N_6861,N_5254,N_5349);
and U6862 (N_6862,N_5710,N_4543);
xor U6863 (N_6863,N_5274,N_5417);
nor U6864 (N_6864,N_5964,N_5004);
and U6865 (N_6865,N_5036,N_4706);
nand U6866 (N_6866,N_5255,N_4678);
nor U6867 (N_6867,N_5869,N_5078);
nor U6868 (N_6868,N_5520,N_5468);
nor U6869 (N_6869,N_5987,N_5332);
or U6870 (N_6870,N_4771,N_5440);
or U6871 (N_6871,N_5438,N_5130);
nand U6872 (N_6872,N_5258,N_4765);
and U6873 (N_6873,N_5339,N_5073);
or U6874 (N_6874,N_5502,N_4576);
and U6875 (N_6875,N_5892,N_5692);
nor U6876 (N_6876,N_5140,N_5370);
and U6877 (N_6877,N_4652,N_5414);
nor U6878 (N_6878,N_5730,N_4524);
nand U6879 (N_6879,N_5469,N_5419);
or U6880 (N_6880,N_5339,N_4787);
nor U6881 (N_6881,N_4955,N_5022);
or U6882 (N_6882,N_5644,N_5243);
nor U6883 (N_6883,N_5980,N_5384);
or U6884 (N_6884,N_5258,N_5794);
and U6885 (N_6885,N_5100,N_4628);
or U6886 (N_6886,N_5063,N_5552);
nor U6887 (N_6887,N_4717,N_5671);
and U6888 (N_6888,N_5674,N_5361);
or U6889 (N_6889,N_5068,N_5449);
and U6890 (N_6890,N_5811,N_5502);
xor U6891 (N_6891,N_5423,N_5630);
xor U6892 (N_6892,N_4992,N_5886);
and U6893 (N_6893,N_4624,N_4707);
and U6894 (N_6894,N_5495,N_5046);
nor U6895 (N_6895,N_5291,N_4703);
and U6896 (N_6896,N_4562,N_5626);
nand U6897 (N_6897,N_5779,N_5061);
nand U6898 (N_6898,N_5351,N_5794);
nor U6899 (N_6899,N_4909,N_5091);
and U6900 (N_6900,N_5708,N_5885);
xor U6901 (N_6901,N_4553,N_5627);
nand U6902 (N_6902,N_5371,N_5598);
xor U6903 (N_6903,N_4739,N_4847);
xnor U6904 (N_6904,N_5056,N_4700);
or U6905 (N_6905,N_5643,N_5408);
nand U6906 (N_6906,N_5068,N_5703);
or U6907 (N_6907,N_5900,N_5011);
nor U6908 (N_6908,N_5048,N_5527);
xnor U6909 (N_6909,N_5006,N_5933);
xor U6910 (N_6910,N_5584,N_5767);
or U6911 (N_6911,N_4573,N_5084);
xnor U6912 (N_6912,N_5480,N_5813);
nand U6913 (N_6913,N_5026,N_4808);
and U6914 (N_6914,N_5631,N_5970);
nor U6915 (N_6915,N_5901,N_5455);
and U6916 (N_6916,N_5920,N_5333);
and U6917 (N_6917,N_5880,N_4822);
nand U6918 (N_6918,N_5450,N_4909);
nand U6919 (N_6919,N_5097,N_4642);
xnor U6920 (N_6920,N_5043,N_5806);
xor U6921 (N_6921,N_5470,N_5166);
or U6922 (N_6922,N_5760,N_5439);
and U6923 (N_6923,N_4519,N_4562);
or U6924 (N_6924,N_5520,N_5222);
or U6925 (N_6925,N_5161,N_5363);
xnor U6926 (N_6926,N_4887,N_4581);
xnor U6927 (N_6927,N_4815,N_5756);
and U6928 (N_6928,N_5015,N_5878);
xnor U6929 (N_6929,N_5994,N_4508);
or U6930 (N_6930,N_5223,N_4713);
nor U6931 (N_6931,N_4759,N_5674);
and U6932 (N_6932,N_4910,N_4766);
nand U6933 (N_6933,N_5699,N_5494);
xor U6934 (N_6934,N_5545,N_4897);
or U6935 (N_6935,N_5852,N_5394);
nand U6936 (N_6936,N_5210,N_5376);
xnor U6937 (N_6937,N_4625,N_4610);
nand U6938 (N_6938,N_5779,N_5954);
xor U6939 (N_6939,N_4806,N_4509);
nor U6940 (N_6940,N_5528,N_4755);
or U6941 (N_6941,N_5149,N_5791);
xnor U6942 (N_6942,N_5206,N_4509);
nand U6943 (N_6943,N_4597,N_5316);
and U6944 (N_6944,N_5814,N_5382);
xnor U6945 (N_6945,N_5823,N_5433);
nor U6946 (N_6946,N_4912,N_4554);
nand U6947 (N_6947,N_5705,N_5623);
nor U6948 (N_6948,N_4568,N_5314);
nor U6949 (N_6949,N_5000,N_5734);
nand U6950 (N_6950,N_5999,N_5642);
or U6951 (N_6951,N_5022,N_5945);
nor U6952 (N_6952,N_5577,N_4662);
nand U6953 (N_6953,N_5981,N_4576);
and U6954 (N_6954,N_4740,N_5953);
or U6955 (N_6955,N_4967,N_5934);
nand U6956 (N_6956,N_4802,N_5587);
nor U6957 (N_6957,N_5235,N_5700);
nor U6958 (N_6958,N_5185,N_5647);
or U6959 (N_6959,N_4690,N_5228);
nor U6960 (N_6960,N_5625,N_5394);
xnor U6961 (N_6961,N_5152,N_4939);
nor U6962 (N_6962,N_4958,N_5963);
and U6963 (N_6963,N_4608,N_5707);
or U6964 (N_6964,N_5650,N_4950);
nand U6965 (N_6965,N_5995,N_4850);
or U6966 (N_6966,N_4621,N_5420);
nor U6967 (N_6967,N_5843,N_5642);
xnor U6968 (N_6968,N_5981,N_5192);
xnor U6969 (N_6969,N_5078,N_4743);
nand U6970 (N_6970,N_5396,N_4543);
xnor U6971 (N_6971,N_4552,N_5156);
nor U6972 (N_6972,N_5516,N_5400);
or U6973 (N_6973,N_5235,N_5025);
xor U6974 (N_6974,N_4578,N_5821);
xnor U6975 (N_6975,N_5840,N_4698);
xnor U6976 (N_6976,N_5873,N_5051);
or U6977 (N_6977,N_5917,N_5942);
or U6978 (N_6978,N_4704,N_5083);
or U6979 (N_6979,N_4808,N_4892);
xor U6980 (N_6980,N_5707,N_5572);
xor U6981 (N_6981,N_5604,N_5046);
nand U6982 (N_6982,N_4929,N_5449);
xor U6983 (N_6983,N_4841,N_5715);
and U6984 (N_6984,N_5452,N_5048);
or U6985 (N_6985,N_4849,N_5863);
or U6986 (N_6986,N_5989,N_4518);
and U6987 (N_6987,N_4742,N_4615);
xnor U6988 (N_6988,N_5949,N_5555);
nor U6989 (N_6989,N_5560,N_5026);
and U6990 (N_6990,N_5893,N_5856);
xnor U6991 (N_6991,N_4637,N_4593);
and U6992 (N_6992,N_5788,N_5766);
nor U6993 (N_6993,N_5870,N_4625);
and U6994 (N_6994,N_5360,N_4911);
or U6995 (N_6995,N_5706,N_5695);
xnor U6996 (N_6996,N_5615,N_4928);
nand U6997 (N_6997,N_5869,N_5962);
xor U6998 (N_6998,N_5204,N_4758);
nand U6999 (N_6999,N_5966,N_5600);
nand U7000 (N_7000,N_5098,N_5029);
or U7001 (N_7001,N_5021,N_4738);
nor U7002 (N_7002,N_5487,N_5062);
and U7003 (N_7003,N_5002,N_4684);
and U7004 (N_7004,N_5768,N_5134);
xnor U7005 (N_7005,N_4874,N_5856);
nor U7006 (N_7006,N_5754,N_5285);
or U7007 (N_7007,N_5705,N_5561);
and U7008 (N_7008,N_4849,N_5134);
nor U7009 (N_7009,N_4863,N_5878);
or U7010 (N_7010,N_5047,N_4834);
or U7011 (N_7011,N_5282,N_4503);
or U7012 (N_7012,N_4721,N_4659);
and U7013 (N_7013,N_5215,N_5764);
nand U7014 (N_7014,N_5167,N_5572);
and U7015 (N_7015,N_5344,N_5746);
and U7016 (N_7016,N_4869,N_5527);
and U7017 (N_7017,N_4919,N_5721);
or U7018 (N_7018,N_5711,N_5289);
or U7019 (N_7019,N_5356,N_5463);
xnor U7020 (N_7020,N_4632,N_5273);
nand U7021 (N_7021,N_5030,N_5812);
and U7022 (N_7022,N_5258,N_4625);
and U7023 (N_7023,N_5831,N_5366);
and U7024 (N_7024,N_5163,N_5747);
xor U7025 (N_7025,N_5470,N_5818);
or U7026 (N_7026,N_5000,N_5616);
and U7027 (N_7027,N_4574,N_4931);
and U7028 (N_7028,N_5892,N_4844);
nand U7029 (N_7029,N_5030,N_5452);
or U7030 (N_7030,N_5154,N_5145);
nor U7031 (N_7031,N_5176,N_5269);
xor U7032 (N_7032,N_4874,N_5873);
nand U7033 (N_7033,N_5105,N_5051);
and U7034 (N_7034,N_5925,N_4699);
nand U7035 (N_7035,N_4864,N_5018);
xnor U7036 (N_7036,N_5114,N_5561);
nor U7037 (N_7037,N_5335,N_4573);
xor U7038 (N_7038,N_5760,N_5804);
nand U7039 (N_7039,N_5869,N_5060);
xnor U7040 (N_7040,N_5476,N_4691);
nand U7041 (N_7041,N_5698,N_5718);
nand U7042 (N_7042,N_4807,N_4984);
nor U7043 (N_7043,N_5575,N_4506);
and U7044 (N_7044,N_4953,N_5592);
or U7045 (N_7045,N_5873,N_5126);
nand U7046 (N_7046,N_5031,N_4752);
or U7047 (N_7047,N_5040,N_4753);
xnor U7048 (N_7048,N_4854,N_4527);
nand U7049 (N_7049,N_4627,N_4722);
and U7050 (N_7050,N_5732,N_5197);
xor U7051 (N_7051,N_4554,N_5287);
nand U7052 (N_7052,N_5675,N_5601);
xnor U7053 (N_7053,N_5618,N_4818);
or U7054 (N_7054,N_5283,N_4932);
nor U7055 (N_7055,N_5862,N_4776);
or U7056 (N_7056,N_5148,N_5633);
or U7057 (N_7057,N_5347,N_5595);
xnor U7058 (N_7058,N_4563,N_4601);
nor U7059 (N_7059,N_5274,N_4936);
and U7060 (N_7060,N_5619,N_5342);
xor U7061 (N_7061,N_5811,N_5284);
or U7062 (N_7062,N_5983,N_4557);
or U7063 (N_7063,N_5832,N_5764);
nand U7064 (N_7064,N_5568,N_4869);
nand U7065 (N_7065,N_5623,N_4680);
xor U7066 (N_7066,N_5376,N_5702);
and U7067 (N_7067,N_5058,N_5253);
nand U7068 (N_7068,N_5443,N_5100);
nor U7069 (N_7069,N_4889,N_5714);
nand U7070 (N_7070,N_5721,N_5662);
or U7071 (N_7071,N_5816,N_5308);
and U7072 (N_7072,N_5527,N_5595);
and U7073 (N_7073,N_5539,N_5027);
xor U7074 (N_7074,N_5217,N_5549);
nor U7075 (N_7075,N_5802,N_4923);
nor U7076 (N_7076,N_5323,N_5899);
or U7077 (N_7077,N_5644,N_5307);
xor U7078 (N_7078,N_5594,N_5486);
and U7079 (N_7079,N_5712,N_5809);
and U7080 (N_7080,N_5937,N_5927);
nand U7081 (N_7081,N_5943,N_5414);
nand U7082 (N_7082,N_5976,N_5673);
nor U7083 (N_7083,N_4609,N_5851);
or U7084 (N_7084,N_5935,N_5788);
nor U7085 (N_7085,N_5155,N_5174);
nand U7086 (N_7086,N_4980,N_4745);
nand U7087 (N_7087,N_4506,N_5707);
and U7088 (N_7088,N_5361,N_5592);
and U7089 (N_7089,N_4601,N_5108);
or U7090 (N_7090,N_4611,N_5279);
nand U7091 (N_7091,N_5482,N_4909);
nand U7092 (N_7092,N_5948,N_4775);
and U7093 (N_7093,N_5426,N_5449);
or U7094 (N_7094,N_5939,N_5667);
nand U7095 (N_7095,N_5749,N_5386);
or U7096 (N_7096,N_5136,N_5025);
nand U7097 (N_7097,N_4844,N_5787);
nand U7098 (N_7098,N_5564,N_5303);
and U7099 (N_7099,N_4918,N_4694);
nand U7100 (N_7100,N_5442,N_5558);
nand U7101 (N_7101,N_5046,N_4794);
xnor U7102 (N_7102,N_5922,N_5519);
xor U7103 (N_7103,N_5219,N_5641);
and U7104 (N_7104,N_5693,N_5955);
xnor U7105 (N_7105,N_5244,N_5427);
or U7106 (N_7106,N_5490,N_4765);
and U7107 (N_7107,N_5495,N_5621);
nand U7108 (N_7108,N_5254,N_5824);
or U7109 (N_7109,N_5664,N_4522);
or U7110 (N_7110,N_5252,N_4663);
and U7111 (N_7111,N_5070,N_5999);
xor U7112 (N_7112,N_5481,N_4507);
xnor U7113 (N_7113,N_4956,N_5108);
nor U7114 (N_7114,N_5123,N_4743);
and U7115 (N_7115,N_5221,N_5929);
and U7116 (N_7116,N_5383,N_5315);
and U7117 (N_7117,N_5797,N_4663);
nor U7118 (N_7118,N_4913,N_5546);
xnor U7119 (N_7119,N_4898,N_5665);
nand U7120 (N_7120,N_4630,N_4637);
and U7121 (N_7121,N_5932,N_5727);
nand U7122 (N_7122,N_5168,N_5357);
or U7123 (N_7123,N_4729,N_5647);
and U7124 (N_7124,N_4893,N_4794);
and U7125 (N_7125,N_4567,N_5804);
nand U7126 (N_7126,N_5472,N_5920);
xor U7127 (N_7127,N_4999,N_4507);
xor U7128 (N_7128,N_5436,N_4830);
nand U7129 (N_7129,N_5879,N_4567);
xnor U7130 (N_7130,N_5809,N_5796);
nor U7131 (N_7131,N_4626,N_5504);
and U7132 (N_7132,N_5088,N_5494);
nand U7133 (N_7133,N_5839,N_5185);
xor U7134 (N_7134,N_5753,N_5927);
nor U7135 (N_7135,N_4603,N_5104);
nor U7136 (N_7136,N_5018,N_5233);
and U7137 (N_7137,N_5664,N_5711);
nor U7138 (N_7138,N_5456,N_4699);
or U7139 (N_7139,N_5088,N_5877);
nor U7140 (N_7140,N_5180,N_5139);
xor U7141 (N_7141,N_5554,N_5817);
xnor U7142 (N_7142,N_4810,N_4728);
or U7143 (N_7143,N_5093,N_5943);
and U7144 (N_7144,N_5183,N_4503);
and U7145 (N_7145,N_4939,N_5236);
nor U7146 (N_7146,N_4736,N_5786);
nor U7147 (N_7147,N_5755,N_4798);
or U7148 (N_7148,N_5957,N_5715);
nor U7149 (N_7149,N_5132,N_5504);
and U7150 (N_7150,N_4905,N_4813);
and U7151 (N_7151,N_4822,N_4850);
and U7152 (N_7152,N_5155,N_4810);
or U7153 (N_7153,N_4645,N_4822);
or U7154 (N_7154,N_5590,N_4786);
nor U7155 (N_7155,N_5846,N_4730);
and U7156 (N_7156,N_4898,N_5744);
nand U7157 (N_7157,N_5268,N_5355);
xor U7158 (N_7158,N_5915,N_5390);
nand U7159 (N_7159,N_5797,N_5690);
xnor U7160 (N_7160,N_4633,N_4785);
nor U7161 (N_7161,N_4783,N_5864);
xnor U7162 (N_7162,N_5824,N_4687);
xor U7163 (N_7163,N_5465,N_4642);
or U7164 (N_7164,N_4771,N_5256);
nor U7165 (N_7165,N_5209,N_4582);
or U7166 (N_7166,N_5164,N_5402);
nor U7167 (N_7167,N_4520,N_5205);
nand U7168 (N_7168,N_5324,N_5567);
and U7169 (N_7169,N_4644,N_5545);
xor U7170 (N_7170,N_4717,N_4524);
nand U7171 (N_7171,N_5693,N_4961);
and U7172 (N_7172,N_5196,N_5608);
nand U7173 (N_7173,N_5124,N_5697);
nand U7174 (N_7174,N_4834,N_4863);
and U7175 (N_7175,N_5058,N_5962);
and U7176 (N_7176,N_5699,N_5833);
and U7177 (N_7177,N_5503,N_5004);
nand U7178 (N_7178,N_4727,N_5279);
nand U7179 (N_7179,N_4896,N_5045);
or U7180 (N_7180,N_5312,N_5301);
and U7181 (N_7181,N_4746,N_5702);
nand U7182 (N_7182,N_5219,N_5146);
nand U7183 (N_7183,N_5516,N_4866);
nor U7184 (N_7184,N_5762,N_4837);
nand U7185 (N_7185,N_5071,N_5105);
xnor U7186 (N_7186,N_5673,N_4983);
and U7187 (N_7187,N_5437,N_4685);
xor U7188 (N_7188,N_5723,N_5231);
and U7189 (N_7189,N_5933,N_5552);
nor U7190 (N_7190,N_5288,N_4891);
nand U7191 (N_7191,N_5908,N_4565);
and U7192 (N_7192,N_5283,N_5641);
nand U7193 (N_7193,N_5981,N_5414);
nand U7194 (N_7194,N_5277,N_4677);
or U7195 (N_7195,N_5911,N_4638);
or U7196 (N_7196,N_4665,N_4935);
or U7197 (N_7197,N_4891,N_5721);
and U7198 (N_7198,N_5293,N_5843);
nor U7199 (N_7199,N_4870,N_5803);
or U7200 (N_7200,N_4834,N_5138);
and U7201 (N_7201,N_4792,N_4793);
nand U7202 (N_7202,N_5571,N_5019);
xor U7203 (N_7203,N_5033,N_4960);
xnor U7204 (N_7204,N_4939,N_4672);
nor U7205 (N_7205,N_4674,N_4987);
nand U7206 (N_7206,N_5910,N_5168);
nand U7207 (N_7207,N_5595,N_4860);
or U7208 (N_7208,N_4680,N_5972);
or U7209 (N_7209,N_5654,N_5736);
or U7210 (N_7210,N_5057,N_5769);
and U7211 (N_7211,N_5458,N_5150);
and U7212 (N_7212,N_5151,N_4715);
nand U7213 (N_7213,N_4559,N_5356);
nor U7214 (N_7214,N_4864,N_5762);
nor U7215 (N_7215,N_5028,N_4973);
or U7216 (N_7216,N_5118,N_5087);
xor U7217 (N_7217,N_4907,N_5647);
and U7218 (N_7218,N_4795,N_4567);
xnor U7219 (N_7219,N_4816,N_4698);
nor U7220 (N_7220,N_4648,N_4731);
or U7221 (N_7221,N_5706,N_4702);
or U7222 (N_7222,N_5733,N_4824);
nor U7223 (N_7223,N_5172,N_5442);
and U7224 (N_7224,N_4782,N_5488);
or U7225 (N_7225,N_5787,N_4685);
nand U7226 (N_7226,N_5614,N_4992);
nor U7227 (N_7227,N_4664,N_4761);
nand U7228 (N_7228,N_5140,N_4757);
xnor U7229 (N_7229,N_5512,N_5090);
nor U7230 (N_7230,N_5168,N_5123);
nand U7231 (N_7231,N_4522,N_4737);
and U7232 (N_7232,N_5994,N_5706);
nor U7233 (N_7233,N_5236,N_5500);
nor U7234 (N_7234,N_5501,N_4877);
xor U7235 (N_7235,N_5349,N_4745);
and U7236 (N_7236,N_5494,N_5039);
and U7237 (N_7237,N_5778,N_4742);
or U7238 (N_7238,N_4977,N_4809);
nor U7239 (N_7239,N_5615,N_5164);
or U7240 (N_7240,N_5922,N_5092);
nand U7241 (N_7241,N_5420,N_4806);
or U7242 (N_7242,N_5336,N_5907);
nand U7243 (N_7243,N_4665,N_5605);
nor U7244 (N_7244,N_5245,N_5965);
nand U7245 (N_7245,N_4746,N_4662);
or U7246 (N_7246,N_4536,N_4874);
or U7247 (N_7247,N_5284,N_5880);
or U7248 (N_7248,N_5536,N_5526);
nor U7249 (N_7249,N_5947,N_5262);
xor U7250 (N_7250,N_5910,N_4863);
nor U7251 (N_7251,N_5894,N_5376);
nor U7252 (N_7252,N_5283,N_5424);
nor U7253 (N_7253,N_4630,N_5560);
xnor U7254 (N_7254,N_5079,N_5797);
nand U7255 (N_7255,N_5315,N_5039);
and U7256 (N_7256,N_5438,N_5190);
or U7257 (N_7257,N_4834,N_4566);
nor U7258 (N_7258,N_5673,N_5878);
and U7259 (N_7259,N_4596,N_5918);
and U7260 (N_7260,N_5926,N_5224);
xnor U7261 (N_7261,N_5671,N_4627);
xnor U7262 (N_7262,N_4814,N_5791);
and U7263 (N_7263,N_5319,N_4713);
xor U7264 (N_7264,N_5046,N_4702);
and U7265 (N_7265,N_4801,N_5862);
nor U7266 (N_7266,N_4858,N_5277);
xor U7267 (N_7267,N_5196,N_4926);
nor U7268 (N_7268,N_5670,N_5701);
nor U7269 (N_7269,N_5895,N_5180);
or U7270 (N_7270,N_4561,N_5884);
nand U7271 (N_7271,N_5053,N_5286);
nor U7272 (N_7272,N_5380,N_4894);
or U7273 (N_7273,N_4977,N_5863);
xor U7274 (N_7274,N_5039,N_5964);
xnor U7275 (N_7275,N_5041,N_5566);
xnor U7276 (N_7276,N_5566,N_5934);
or U7277 (N_7277,N_5520,N_5054);
nand U7278 (N_7278,N_5545,N_4937);
xnor U7279 (N_7279,N_5972,N_4702);
or U7280 (N_7280,N_5025,N_4694);
nor U7281 (N_7281,N_4630,N_5227);
and U7282 (N_7282,N_5505,N_5033);
nor U7283 (N_7283,N_5923,N_4517);
or U7284 (N_7284,N_5868,N_4593);
nand U7285 (N_7285,N_5505,N_5623);
nor U7286 (N_7286,N_4528,N_4924);
and U7287 (N_7287,N_4585,N_4607);
nor U7288 (N_7288,N_5200,N_5060);
nand U7289 (N_7289,N_4802,N_5324);
xnor U7290 (N_7290,N_4982,N_5919);
or U7291 (N_7291,N_4820,N_4764);
nand U7292 (N_7292,N_5915,N_4796);
nand U7293 (N_7293,N_4955,N_5512);
nor U7294 (N_7294,N_4826,N_4759);
nand U7295 (N_7295,N_5740,N_5179);
or U7296 (N_7296,N_4876,N_5058);
or U7297 (N_7297,N_5534,N_4537);
nand U7298 (N_7298,N_5026,N_5035);
nor U7299 (N_7299,N_5496,N_5209);
nand U7300 (N_7300,N_5409,N_4932);
and U7301 (N_7301,N_5381,N_5911);
nor U7302 (N_7302,N_4588,N_5892);
nand U7303 (N_7303,N_4541,N_4962);
nor U7304 (N_7304,N_4674,N_4979);
xnor U7305 (N_7305,N_5285,N_4713);
xnor U7306 (N_7306,N_5130,N_5004);
xnor U7307 (N_7307,N_5511,N_5021);
xnor U7308 (N_7308,N_5776,N_4554);
nand U7309 (N_7309,N_5781,N_5859);
xor U7310 (N_7310,N_4666,N_5722);
nor U7311 (N_7311,N_5336,N_5459);
and U7312 (N_7312,N_5992,N_5109);
or U7313 (N_7313,N_5505,N_5660);
xor U7314 (N_7314,N_5398,N_5893);
nand U7315 (N_7315,N_4760,N_4853);
nand U7316 (N_7316,N_5542,N_4640);
nor U7317 (N_7317,N_5783,N_5618);
xnor U7318 (N_7318,N_4988,N_5958);
nor U7319 (N_7319,N_5618,N_5091);
nand U7320 (N_7320,N_5507,N_5019);
xnor U7321 (N_7321,N_5140,N_4501);
nor U7322 (N_7322,N_4773,N_5350);
and U7323 (N_7323,N_5965,N_5197);
and U7324 (N_7324,N_5854,N_5181);
nor U7325 (N_7325,N_5955,N_4888);
nand U7326 (N_7326,N_5623,N_5307);
xor U7327 (N_7327,N_4939,N_5041);
nand U7328 (N_7328,N_5666,N_5845);
xor U7329 (N_7329,N_4895,N_5817);
nor U7330 (N_7330,N_5133,N_5620);
and U7331 (N_7331,N_5622,N_5244);
nor U7332 (N_7332,N_5800,N_4930);
xor U7333 (N_7333,N_5303,N_5750);
or U7334 (N_7334,N_5216,N_4656);
nand U7335 (N_7335,N_5270,N_5369);
or U7336 (N_7336,N_5089,N_5752);
xnor U7337 (N_7337,N_5822,N_5806);
and U7338 (N_7338,N_5517,N_5771);
nand U7339 (N_7339,N_5157,N_5444);
nand U7340 (N_7340,N_5905,N_5886);
xor U7341 (N_7341,N_4541,N_5624);
nor U7342 (N_7342,N_4716,N_4756);
nand U7343 (N_7343,N_5862,N_5148);
or U7344 (N_7344,N_4604,N_5029);
nand U7345 (N_7345,N_5441,N_5445);
nor U7346 (N_7346,N_5673,N_4870);
and U7347 (N_7347,N_5580,N_5026);
nand U7348 (N_7348,N_4966,N_5880);
nor U7349 (N_7349,N_5514,N_4800);
and U7350 (N_7350,N_4839,N_4810);
nand U7351 (N_7351,N_5945,N_4636);
and U7352 (N_7352,N_4767,N_5434);
or U7353 (N_7353,N_4924,N_4711);
or U7354 (N_7354,N_4658,N_5008);
and U7355 (N_7355,N_5325,N_5202);
or U7356 (N_7356,N_4816,N_5044);
nand U7357 (N_7357,N_5957,N_5467);
nand U7358 (N_7358,N_4769,N_5034);
nand U7359 (N_7359,N_5392,N_4921);
nand U7360 (N_7360,N_5430,N_5056);
or U7361 (N_7361,N_5322,N_5791);
nand U7362 (N_7362,N_5368,N_4968);
nand U7363 (N_7363,N_5891,N_5671);
and U7364 (N_7364,N_4746,N_5555);
or U7365 (N_7365,N_4506,N_5882);
xor U7366 (N_7366,N_5377,N_5029);
and U7367 (N_7367,N_5697,N_4643);
nand U7368 (N_7368,N_5480,N_4518);
or U7369 (N_7369,N_5391,N_5155);
nand U7370 (N_7370,N_4569,N_4639);
and U7371 (N_7371,N_5636,N_5861);
or U7372 (N_7372,N_5139,N_5650);
or U7373 (N_7373,N_5414,N_4580);
and U7374 (N_7374,N_5449,N_5032);
nor U7375 (N_7375,N_5308,N_4568);
or U7376 (N_7376,N_5355,N_4825);
xor U7377 (N_7377,N_4735,N_5644);
xnor U7378 (N_7378,N_5819,N_5607);
nor U7379 (N_7379,N_5110,N_4725);
nor U7380 (N_7380,N_5124,N_5836);
or U7381 (N_7381,N_5998,N_5377);
nand U7382 (N_7382,N_5587,N_5813);
nand U7383 (N_7383,N_4699,N_5813);
nor U7384 (N_7384,N_5361,N_5108);
and U7385 (N_7385,N_5397,N_4910);
nor U7386 (N_7386,N_5480,N_5797);
xor U7387 (N_7387,N_5453,N_4701);
xor U7388 (N_7388,N_5625,N_5168);
nor U7389 (N_7389,N_5511,N_5715);
or U7390 (N_7390,N_5133,N_5330);
xor U7391 (N_7391,N_5815,N_5891);
nand U7392 (N_7392,N_5824,N_4944);
or U7393 (N_7393,N_5778,N_5362);
nand U7394 (N_7394,N_5841,N_4791);
or U7395 (N_7395,N_5156,N_5993);
nor U7396 (N_7396,N_5547,N_5584);
nand U7397 (N_7397,N_5837,N_5143);
nor U7398 (N_7398,N_5380,N_4853);
nand U7399 (N_7399,N_5921,N_5222);
xor U7400 (N_7400,N_5985,N_5645);
xor U7401 (N_7401,N_5621,N_5672);
and U7402 (N_7402,N_4519,N_4616);
or U7403 (N_7403,N_5474,N_5272);
and U7404 (N_7404,N_5845,N_4594);
nor U7405 (N_7405,N_4916,N_5773);
xor U7406 (N_7406,N_5167,N_5864);
nor U7407 (N_7407,N_5435,N_5271);
and U7408 (N_7408,N_5228,N_4604);
nor U7409 (N_7409,N_4646,N_4988);
xor U7410 (N_7410,N_5616,N_5523);
nor U7411 (N_7411,N_5986,N_4548);
or U7412 (N_7412,N_5842,N_4840);
and U7413 (N_7413,N_5371,N_5660);
nand U7414 (N_7414,N_5223,N_4593);
nand U7415 (N_7415,N_5368,N_5636);
or U7416 (N_7416,N_5778,N_5257);
or U7417 (N_7417,N_4764,N_4605);
xor U7418 (N_7418,N_5859,N_4610);
xnor U7419 (N_7419,N_4619,N_5822);
or U7420 (N_7420,N_5794,N_4558);
and U7421 (N_7421,N_4546,N_5344);
xor U7422 (N_7422,N_5290,N_4884);
and U7423 (N_7423,N_5757,N_4893);
xor U7424 (N_7424,N_4970,N_5468);
or U7425 (N_7425,N_5814,N_5886);
or U7426 (N_7426,N_5997,N_5158);
nor U7427 (N_7427,N_5660,N_5441);
xor U7428 (N_7428,N_5093,N_4787);
nor U7429 (N_7429,N_4603,N_5162);
nor U7430 (N_7430,N_5937,N_4814);
nor U7431 (N_7431,N_4840,N_4829);
nor U7432 (N_7432,N_5031,N_5018);
nand U7433 (N_7433,N_4526,N_4885);
or U7434 (N_7434,N_5010,N_5485);
or U7435 (N_7435,N_5028,N_4854);
nor U7436 (N_7436,N_4725,N_4560);
xor U7437 (N_7437,N_5423,N_5805);
xor U7438 (N_7438,N_5179,N_5928);
or U7439 (N_7439,N_4699,N_5003);
and U7440 (N_7440,N_5600,N_5754);
and U7441 (N_7441,N_4566,N_5573);
xnor U7442 (N_7442,N_5324,N_5374);
and U7443 (N_7443,N_5064,N_5804);
nand U7444 (N_7444,N_5563,N_5737);
and U7445 (N_7445,N_4702,N_5553);
nor U7446 (N_7446,N_4780,N_5651);
nor U7447 (N_7447,N_5113,N_5032);
nor U7448 (N_7448,N_5068,N_5234);
nor U7449 (N_7449,N_4894,N_4895);
and U7450 (N_7450,N_4606,N_5556);
xnor U7451 (N_7451,N_5118,N_5664);
nand U7452 (N_7452,N_5722,N_5078);
nor U7453 (N_7453,N_4904,N_5962);
nand U7454 (N_7454,N_5262,N_5837);
xnor U7455 (N_7455,N_4559,N_4503);
xnor U7456 (N_7456,N_5299,N_4548);
or U7457 (N_7457,N_5436,N_5480);
xnor U7458 (N_7458,N_5245,N_4543);
xor U7459 (N_7459,N_4645,N_5419);
xnor U7460 (N_7460,N_5212,N_5236);
nand U7461 (N_7461,N_4763,N_5483);
nor U7462 (N_7462,N_5268,N_5545);
and U7463 (N_7463,N_5430,N_5090);
or U7464 (N_7464,N_5458,N_4741);
and U7465 (N_7465,N_5230,N_5414);
or U7466 (N_7466,N_4705,N_5508);
or U7467 (N_7467,N_5184,N_4761);
and U7468 (N_7468,N_5330,N_5287);
or U7469 (N_7469,N_5143,N_5874);
xor U7470 (N_7470,N_5336,N_5232);
or U7471 (N_7471,N_4901,N_5853);
nand U7472 (N_7472,N_4759,N_5749);
and U7473 (N_7473,N_5438,N_5775);
nand U7474 (N_7474,N_4537,N_4626);
or U7475 (N_7475,N_5092,N_5719);
or U7476 (N_7476,N_5623,N_5862);
and U7477 (N_7477,N_5512,N_5876);
and U7478 (N_7478,N_5232,N_4650);
nand U7479 (N_7479,N_5285,N_5247);
xnor U7480 (N_7480,N_5175,N_4853);
and U7481 (N_7481,N_5044,N_5170);
and U7482 (N_7482,N_5461,N_5589);
xor U7483 (N_7483,N_5700,N_5822);
xnor U7484 (N_7484,N_4847,N_4621);
xor U7485 (N_7485,N_5724,N_5649);
and U7486 (N_7486,N_4703,N_5161);
nand U7487 (N_7487,N_5477,N_4686);
xnor U7488 (N_7488,N_5348,N_5171);
or U7489 (N_7489,N_5639,N_5524);
nand U7490 (N_7490,N_5328,N_4748);
nand U7491 (N_7491,N_5120,N_5918);
and U7492 (N_7492,N_4985,N_4648);
nand U7493 (N_7493,N_4905,N_4750);
or U7494 (N_7494,N_5637,N_4688);
or U7495 (N_7495,N_4724,N_5560);
xor U7496 (N_7496,N_5403,N_5040);
nor U7497 (N_7497,N_5922,N_4642);
or U7498 (N_7498,N_5113,N_5630);
or U7499 (N_7499,N_4839,N_4992);
xnor U7500 (N_7500,N_7148,N_6367);
and U7501 (N_7501,N_6852,N_7015);
and U7502 (N_7502,N_7251,N_6180);
xor U7503 (N_7503,N_7175,N_6307);
or U7504 (N_7504,N_7159,N_6335);
nor U7505 (N_7505,N_6044,N_7256);
nand U7506 (N_7506,N_6060,N_6828);
or U7507 (N_7507,N_7496,N_6276);
or U7508 (N_7508,N_7086,N_6043);
or U7509 (N_7509,N_7187,N_6315);
and U7510 (N_7510,N_6354,N_7419);
xor U7511 (N_7511,N_6869,N_6213);
and U7512 (N_7512,N_6314,N_7336);
nor U7513 (N_7513,N_6322,N_6170);
nor U7514 (N_7514,N_6110,N_6544);
nor U7515 (N_7515,N_6208,N_6706);
or U7516 (N_7516,N_6453,N_6870);
and U7517 (N_7517,N_6616,N_6358);
and U7518 (N_7518,N_7166,N_7369);
or U7519 (N_7519,N_7316,N_6030);
nor U7520 (N_7520,N_6301,N_7169);
and U7521 (N_7521,N_7351,N_6565);
xor U7522 (N_7522,N_7042,N_6466);
nor U7523 (N_7523,N_7073,N_7285);
nand U7524 (N_7524,N_7374,N_6951);
nand U7525 (N_7525,N_6617,N_7453);
and U7526 (N_7526,N_6000,N_7286);
nand U7527 (N_7527,N_6943,N_6730);
nor U7528 (N_7528,N_7459,N_6272);
nor U7529 (N_7529,N_6778,N_7079);
and U7530 (N_7530,N_6142,N_6561);
nor U7531 (N_7531,N_7326,N_7139);
nor U7532 (N_7532,N_6871,N_7360);
nor U7533 (N_7533,N_6411,N_6250);
or U7534 (N_7534,N_6189,N_6143);
and U7535 (N_7535,N_7051,N_6967);
nand U7536 (N_7536,N_7184,N_7147);
xor U7537 (N_7537,N_7120,N_7119);
or U7538 (N_7538,N_6837,N_7335);
xor U7539 (N_7539,N_7047,N_6663);
and U7540 (N_7540,N_6239,N_6868);
xor U7541 (N_7541,N_7392,N_6963);
nand U7542 (N_7542,N_7080,N_6686);
or U7543 (N_7543,N_7477,N_6102);
and U7544 (N_7544,N_7221,N_6097);
or U7545 (N_7545,N_6210,N_6111);
xor U7546 (N_7546,N_7087,N_7261);
xor U7547 (N_7547,N_6710,N_6693);
and U7548 (N_7548,N_6678,N_6506);
nor U7549 (N_7549,N_6292,N_7058);
nor U7550 (N_7550,N_7274,N_6540);
or U7551 (N_7551,N_6896,N_6287);
nor U7552 (N_7552,N_6149,N_7240);
or U7553 (N_7553,N_7259,N_6619);
nand U7554 (N_7554,N_6045,N_7010);
nand U7555 (N_7555,N_6578,N_7269);
nand U7556 (N_7556,N_6118,N_7299);
nor U7557 (N_7557,N_6222,N_6817);
nand U7558 (N_7558,N_6878,N_7262);
nand U7559 (N_7559,N_6254,N_7408);
nand U7560 (N_7560,N_6542,N_7065);
xor U7561 (N_7561,N_6692,N_6586);
nand U7562 (N_7562,N_6297,N_7355);
nor U7563 (N_7563,N_6327,N_6843);
xor U7564 (N_7564,N_6526,N_7099);
nand U7565 (N_7565,N_6701,N_6401);
or U7566 (N_7566,N_6700,N_6038);
xor U7567 (N_7567,N_6621,N_6995);
or U7568 (N_7568,N_6822,N_7331);
nand U7569 (N_7569,N_6650,N_7263);
nor U7570 (N_7570,N_6491,N_6167);
xor U7571 (N_7571,N_7378,N_6086);
and U7572 (N_7572,N_7228,N_7224);
nor U7573 (N_7573,N_6488,N_6691);
nor U7574 (N_7574,N_6976,N_6465);
and U7575 (N_7575,N_7070,N_7029);
nor U7576 (N_7576,N_6410,N_6115);
and U7577 (N_7577,N_6009,N_6187);
or U7578 (N_7578,N_6298,N_7445);
nand U7579 (N_7579,N_6742,N_6428);
nand U7580 (N_7580,N_7101,N_7050);
and U7581 (N_7581,N_7179,N_6626);
nand U7582 (N_7582,N_6894,N_6863);
or U7583 (N_7583,N_6198,N_6237);
and U7584 (N_7584,N_7386,N_6027);
and U7585 (N_7585,N_6763,N_6734);
nand U7586 (N_7586,N_6741,N_7370);
nand U7587 (N_7587,N_7442,N_6932);
and U7588 (N_7588,N_6338,N_7132);
nor U7589 (N_7589,N_6560,N_6429);
nand U7590 (N_7590,N_7188,N_6849);
nand U7591 (N_7591,N_6886,N_7491);
nand U7592 (N_7592,N_6439,N_6685);
nand U7593 (N_7593,N_6786,N_6673);
xnor U7594 (N_7594,N_6842,N_6585);
and U7595 (N_7595,N_7232,N_6061);
and U7596 (N_7596,N_6773,N_6620);
or U7597 (N_7597,N_7174,N_6015);
xor U7598 (N_7598,N_7458,N_7154);
nand U7599 (N_7599,N_7110,N_6305);
nor U7600 (N_7600,N_6472,N_6670);
xnor U7601 (N_7601,N_6225,N_7094);
nand U7602 (N_7602,N_7034,N_7171);
and U7603 (N_7603,N_7217,N_6860);
nor U7604 (N_7604,N_6994,N_7338);
and U7605 (N_7605,N_6675,N_7095);
xnor U7606 (N_7606,N_6241,N_7401);
nor U7607 (N_7607,N_6395,N_6722);
or U7608 (N_7608,N_6820,N_7332);
nand U7609 (N_7609,N_6386,N_6368);
or U7610 (N_7610,N_7462,N_6028);
xor U7611 (N_7611,N_6193,N_6515);
xnor U7612 (N_7612,N_6255,N_6851);
xor U7613 (N_7613,N_7267,N_7125);
and U7614 (N_7614,N_7093,N_7032);
nor U7615 (N_7615,N_6037,N_7384);
nand U7616 (N_7616,N_6486,N_6014);
or U7617 (N_7617,N_6764,N_6853);
nand U7618 (N_7618,N_7046,N_7487);
or U7619 (N_7619,N_6775,N_6771);
or U7620 (N_7620,N_6668,N_6478);
and U7621 (N_7621,N_6952,N_6231);
or U7622 (N_7622,N_6072,N_6376);
xnor U7623 (N_7623,N_7353,N_7287);
and U7624 (N_7624,N_6985,N_6532);
and U7625 (N_7625,N_6294,N_6036);
and U7626 (N_7626,N_6873,N_6503);
or U7627 (N_7627,N_6484,N_6343);
xor U7628 (N_7628,N_6081,N_7216);
and U7629 (N_7629,N_6854,N_6330);
or U7630 (N_7630,N_6965,N_6993);
or U7631 (N_7631,N_6059,N_6520);
and U7632 (N_7632,N_6823,N_7118);
nand U7633 (N_7633,N_6024,N_7172);
nand U7634 (N_7634,N_6169,N_6404);
xor U7635 (N_7635,N_7466,N_6676);
xor U7636 (N_7636,N_7035,N_6933);
nand U7637 (N_7637,N_6783,N_6726);
xnor U7638 (N_7638,N_6594,N_6725);
nand U7639 (N_7639,N_7354,N_6275);
nor U7640 (N_7640,N_6375,N_7135);
nand U7641 (N_7641,N_6648,N_6988);
nor U7642 (N_7642,N_7303,N_6555);
and U7643 (N_7643,N_7106,N_7003);
nand U7644 (N_7644,N_6447,N_6895);
xor U7645 (N_7645,N_7253,N_6291);
and U7646 (N_7646,N_7182,N_6321);
and U7647 (N_7647,N_6805,N_6328);
nor U7648 (N_7648,N_6940,N_6482);
or U7649 (N_7649,N_6107,N_6039);
xnor U7650 (N_7650,N_7218,N_7385);
or U7651 (N_7651,N_6845,N_6891);
or U7652 (N_7652,N_6247,N_7464);
or U7653 (N_7653,N_6510,N_6002);
nor U7654 (N_7654,N_6899,N_7140);
nor U7655 (N_7655,N_7243,N_6598);
and U7656 (N_7656,N_6025,N_6062);
nand U7657 (N_7657,N_7468,N_7470);
nor U7658 (N_7658,N_6419,N_6076);
nand U7659 (N_7659,N_6541,N_6504);
or U7660 (N_7660,N_6113,N_6904);
and U7661 (N_7661,N_6847,N_6052);
nand U7662 (N_7662,N_6957,N_6412);
nor U7663 (N_7663,N_6796,N_7318);
or U7664 (N_7664,N_6385,N_6906);
nand U7665 (N_7665,N_7089,N_6887);
and U7666 (N_7666,N_6144,N_7198);
nand U7667 (N_7667,N_6454,N_7455);
or U7668 (N_7668,N_6013,N_6529);
xor U7669 (N_7669,N_6205,N_6604);
nor U7670 (N_7670,N_7022,N_6268);
or U7671 (N_7671,N_6825,N_6001);
and U7672 (N_7672,N_6393,N_6492);
or U7673 (N_7673,N_7072,N_7078);
nor U7674 (N_7674,N_6166,N_6217);
or U7675 (N_7675,N_7381,N_6662);
nor U7676 (N_7676,N_6093,N_7438);
nor U7677 (N_7677,N_6681,N_7031);
nor U7678 (N_7678,N_7199,N_6318);
nand U7679 (N_7679,N_6339,N_7001);
and U7680 (N_7680,N_7157,N_7241);
and U7681 (N_7681,N_6117,N_6575);
and U7682 (N_7682,N_7129,N_7498);
and U7683 (N_7683,N_7479,N_7493);
nor U7684 (N_7684,N_7478,N_7225);
nand U7685 (N_7685,N_7446,N_6151);
nand U7686 (N_7686,N_7163,N_6426);
xnor U7687 (N_7687,N_7201,N_6416);
or U7688 (N_7688,N_6096,N_6876);
nand U7689 (N_7689,N_6483,N_7002);
nor U7690 (N_7690,N_6928,N_6751);
xnor U7691 (N_7691,N_6601,N_6260);
nor U7692 (N_7692,N_7048,N_6020);
xor U7693 (N_7693,N_6070,N_7363);
xnor U7694 (N_7694,N_6754,N_6194);
or U7695 (N_7695,N_6802,N_6377);
nand U7696 (N_7696,N_6090,N_7437);
nand U7697 (N_7697,N_6396,N_6089);
nand U7698 (N_7698,N_7308,N_7111);
nand U7699 (N_7699,N_6155,N_6135);
or U7700 (N_7700,N_6229,N_6538);
nor U7701 (N_7701,N_6912,N_6644);
nand U7702 (N_7702,N_6122,N_6073);
and U7703 (N_7703,N_6104,N_6183);
nor U7704 (N_7704,N_7113,N_6640);
xnor U7705 (N_7705,N_7314,N_7309);
or U7706 (N_7706,N_7451,N_7289);
nor U7707 (N_7707,N_6859,N_7114);
and U7708 (N_7708,N_7481,N_6679);
or U7709 (N_7709,N_7246,N_6402);
and U7710 (N_7710,N_7030,N_6266);
xnor U7711 (N_7711,N_6890,N_7038);
or U7712 (N_7712,N_6168,N_6069);
or U7713 (N_7713,N_6862,N_6991);
nor U7714 (N_7714,N_6079,N_7238);
and U7715 (N_7715,N_6924,N_6739);
nand U7716 (N_7716,N_6903,N_6035);
nand U7717 (N_7717,N_7415,N_7327);
nor U7718 (N_7718,N_7317,N_6827);
xor U7719 (N_7719,N_6065,N_6005);
nor U7720 (N_7720,N_6197,N_6989);
or U7721 (N_7721,N_7143,N_6085);
xor U7722 (N_7722,N_7069,N_6078);
xor U7723 (N_7723,N_6969,N_7206);
nor U7724 (N_7724,N_6190,N_6782);
nor U7725 (N_7725,N_6109,N_6941);
and U7726 (N_7726,N_6579,N_6092);
xnor U7727 (N_7727,N_6527,N_7420);
and U7728 (N_7728,N_6926,N_7024);
and U7729 (N_7729,N_6975,N_6731);
nor U7730 (N_7730,N_6793,N_6622);
nand U7731 (N_7731,N_6577,N_6974);
xor U7732 (N_7732,N_6175,N_7176);
nand U7733 (N_7733,N_6206,N_6557);
xnor U7734 (N_7734,N_6407,N_6505);
or U7735 (N_7735,N_6211,N_6087);
and U7736 (N_7736,N_7480,N_6753);
or U7737 (N_7737,N_6497,N_6106);
nand U7738 (N_7738,N_6935,N_7431);
and U7739 (N_7739,N_7016,N_6592);
and U7740 (N_7740,N_7472,N_7195);
xor U7741 (N_7741,N_6264,N_6769);
nand U7742 (N_7742,N_6902,N_6792);
and U7743 (N_7743,N_6784,N_6067);
and U7744 (N_7744,N_6664,N_6865);
and U7745 (N_7745,N_6137,N_6643);
nand U7746 (N_7746,N_6958,N_6955);
nand U7747 (N_7747,N_7227,N_6979);
nand U7748 (N_7748,N_6549,N_7011);
or U7749 (N_7749,N_6745,N_6159);
nand U7750 (N_7750,N_6336,N_6129);
or U7751 (N_7751,N_7194,N_6815);
and U7752 (N_7752,N_7068,N_6750);
nand U7753 (N_7753,N_6382,N_6641);
nor U7754 (N_7754,N_6178,N_6179);
or U7755 (N_7755,N_6232,N_7250);
or U7756 (N_7756,N_6489,N_6204);
xor U7757 (N_7757,N_7325,N_7337);
nand U7758 (N_7758,N_6942,N_6639);
or U7759 (N_7759,N_7105,N_7142);
or U7760 (N_7760,N_7364,N_6939);
nand U7761 (N_7761,N_6344,N_6680);
nor U7762 (N_7762,N_6591,N_6729);
nor U7763 (N_7763,N_6576,N_7208);
xor U7764 (N_7764,N_7060,N_6425);
nand U7765 (N_7765,N_6732,N_6398);
nor U7766 (N_7766,N_6451,N_6334);
xnor U7767 (N_7767,N_6273,N_6471);
xor U7768 (N_7768,N_7304,N_6571);
or U7769 (N_7769,N_7434,N_6308);
nand U7770 (N_7770,N_6761,N_6160);
nor U7771 (N_7771,N_6997,N_7495);
nor U7772 (N_7772,N_6953,N_6238);
xor U7773 (N_7773,N_7151,N_6657);
nor U7774 (N_7774,N_6552,N_7145);
and U7775 (N_7775,N_6534,N_7026);
or U7776 (N_7776,N_6123,N_7074);
nor U7777 (N_7777,N_7405,N_6223);
nand U7778 (N_7778,N_6171,N_7191);
or U7779 (N_7779,N_6911,N_6120);
xor U7780 (N_7780,N_6119,N_7380);
nor U7781 (N_7781,N_6281,N_6219);
nor U7782 (N_7782,N_6262,N_6400);
nand U7783 (N_7783,N_6518,N_7203);
or U7784 (N_7784,N_7357,N_6799);
or U7785 (N_7785,N_6444,N_6116);
and U7786 (N_7786,N_7350,N_6636);
nand U7787 (N_7787,N_6360,N_7411);
and U7788 (N_7788,N_6186,N_7117);
nand U7789 (N_7789,N_6893,N_7280);
nor U7790 (N_7790,N_7102,N_6790);
nand U7791 (N_7791,N_7367,N_6258);
and U7792 (N_7792,N_7229,N_6177);
nor U7793 (N_7793,N_6509,N_6480);
nand U7794 (N_7794,N_6188,N_6574);
nor U7795 (N_7795,N_6346,N_6968);
or U7796 (N_7796,N_7312,N_7168);
and U7797 (N_7797,N_6758,N_6733);
or U7798 (N_7798,N_6776,N_7282);
xnor U7799 (N_7799,N_7435,N_6253);
or U7800 (N_7800,N_7319,N_7213);
nor U7801 (N_7801,N_6708,N_6345);
or U7802 (N_7802,N_6645,N_6176);
or U7803 (N_7803,N_6284,N_7160);
or U7804 (N_7804,N_6448,N_7009);
nand U7805 (N_7805,N_6618,N_6514);
nand U7806 (N_7806,N_6788,N_6033);
nand U7807 (N_7807,N_6835,N_7084);
or U7808 (N_7808,N_6533,N_7348);
and U7809 (N_7809,N_6913,N_6295);
xor U7810 (N_7810,N_7146,N_7413);
nor U7811 (N_7811,N_6537,N_7247);
nand U7812 (N_7812,N_6257,N_6218);
nand U7813 (N_7813,N_6779,N_7271);
xor U7814 (N_7814,N_6858,N_7448);
nor U7815 (N_7815,N_7340,N_7368);
xor U7816 (N_7816,N_6744,N_7008);
or U7817 (N_7817,N_6512,N_6789);
nor U7818 (N_7818,N_7422,N_7379);
xor U7819 (N_7819,N_6811,N_6406);
or U7820 (N_7820,N_7085,N_6612);
xnor U7821 (N_7821,N_6587,N_6422);
nor U7822 (N_7822,N_7347,N_6813);
or U7823 (N_7823,N_6804,N_6332);
nor U7824 (N_7824,N_7215,N_6918);
and U7825 (N_7825,N_6234,N_7233);
or U7826 (N_7826,N_6630,N_6140);
nor U7827 (N_7827,N_7257,N_6839);
nor U7828 (N_7828,N_6589,N_6163);
xor U7829 (N_7829,N_6103,N_6524);
or U7830 (N_7830,N_7020,N_6256);
nor U7831 (N_7831,N_7124,N_6606);
nor U7832 (N_7832,N_6495,N_6535);
nand U7833 (N_7833,N_6289,N_6554);
nor U7834 (N_7834,N_6249,N_7063);
nand U7835 (N_7835,N_6007,N_6814);
nor U7836 (N_7836,N_7320,N_6145);
or U7837 (N_7837,N_7334,N_7185);
nor U7838 (N_7838,N_6525,N_6199);
xnor U7839 (N_7839,N_6808,N_6596);
nand U7840 (N_7840,N_7417,N_6930);
nand U7841 (N_7841,N_7043,N_6909);
nor U7842 (N_7842,N_6702,N_6908);
nor U7843 (N_7843,N_7362,N_7018);
and U7844 (N_7844,N_6768,N_6203);
nand U7845 (N_7845,N_6767,N_7397);
and U7846 (N_7846,N_7281,N_7219);
xnor U7847 (N_7847,N_6174,N_6597);
nor U7848 (N_7848,N_6371,N_6202);
or U7849 (N_7849,N_7077,N_6456);
nor U7850 (N_7850,N_7393,N_7366);
nor U7851 (N_7851,N_6818,N_6660);
nor U7852 (N_7852,N_6323,N_6875);
xor U7853 (N_7853,N_7329,N_6154);
and U7854 (N_7854,N_7301,N_6785);
nor U7855 (N_7855,N_7040,N_6653);
or U7856 (N_7856,N_6624,N_6511);
and U7857 (N_7857,N_7483,N_6987);
xor U7858 (N_7858,N_7284,N_6271);
or U7859 (N_7859,N_6165,N_6468);
nand U7860 (N_7860,N_6138,N_6695);
or U7861 (N_7861,N_6564,N_6424);
or U7862 (N_7862,N_6800,N_7115);
nor U7863 (N_7863,N_7400,N_7014);
or U7864 (N_7864,N_7447,N_6770);
and U7865 (N_7865,N_6302,N_7323);
and U7866 (N_7866,N_7432,N_6359);
nor U7867 (N_7867,N_6777,N_7162);
nand U7868 (N_7868,N_7499,N_7190);
nor U7869 (N_7869,N_6267,N_6493);
xnor U7870 (N_7870,N_6714,N_7398);
nand U7871 (N_7871,N_6522,N_7409);
nor U7872 (N_7872,N_6973,N_7096);
xnor U7873 (N_7873,N_7012,N_6916);
nor U7874 (N_7874,N_6834,N_7399);
and U7875 (N_7875,N_6282,N_7053);
and U7876 (N_7876,N_7028,N_7097);
xnor U7877 (N_7877,N_7359,N_7144);
and U7878 (N_7878,N_7244,N_6934);
xor U7879 (N_7879,N_6801,N_6944);
xnor U7880 (N_7880,N_6915,N_6403);
nor U7881 (N_7881,N_6684,N_6373);
nand U7882 (N_7882,N_6050,N_6531);
xnor U7883 (N_7883,N_6759,N_7231);
and U7884 (N_7884,N_6659,N_6080);
nand U7885 (N_7885,N_6667,N_7473);
and U7886 (N_7886,N_6048,N_6476);
nor U7887 (N_7887,N_6477,N_7311);
xor U7888 (N_7888,N_6195,N_6420);
xor U7889 (N_7889,N_6463,N_6927);
or U7890 (N_7890,N_6711,N_7361);
and U7891 (N_7891,N_6341,N_6569);
nand U7892 (N_7892,N_7330,N_6088);
and U7893 (N_7893,N_7277,N_7436);
nor U7894 (N_7894,N_6724,N_7450);
nor U7895 (N_7895,N_6885,N_7297);
or U7896 (N_7896,N_6185,N_6459);
and U7897 (N_7897,N_7109,N_6923);
nor U7898 (N_7898,N_6889,N_7457);
xnor U7899 (N_7899,N_6409,N_7088);
or U7900 (N_7900,N_7180,N_6765);
xnor U7901 (N_7901,N_6917,N_6992);
nand U7902 (N_7902,N_7222,N_6721);
or U7903 (N_7903,N_7039,N_7130);
xnor U7904 (N_7904,N_6948,N_6689);
and U7905 (N_7905,N_7212,N_7258);
xnor U7906 (N_7906,N_7486,N_6583);
xnor U7907 (N_7907,N_7234,N_6674);
or U7908 (N_7908,N_7476,N_6697);
or U7909 (N_7909,N_6687,N_6966);
nand U7910 (N_7910,N_7196,N_7025);
or U7911 (N_7911,N_6436,N_6856);
xor U7912 (N_7912,N_7375,N_6156);
and U7913 (N_7913,N_6746,N_6405);
nor U7914 (N_7914,N_6300,N_7428);
xor U7915 (N_7915,N_6055,N_7383);
xnor U7916 (N_7916,N_7441,N_6325);
or U7917 (N_7917,N_6430,N_6164);
nand U7918 (N_7918,N_6629,N_6513);
nor U7919 (N_7919,N_6632,N_6372);
nor U7920 (N_7920,N_6666,N_7341);
and U7921 (N_7921,N_7279,N_6011);
nand U7922 (N_7922,N_6830,N_6914);
and U7923 (N_7923,N_6573,N_7298);
nand U7924 (N_7924,N_7183,N_6872);
nand U7925 (N_7925,N_6348,N_6091);
xor U7926 (N_7926,N_7292,N_6831);
nor U7927 (N_7927,N_7211,N_7021);
and U7928 (N_7928,N_6920,N_6907);
nand U7929 (N_7929,N_7425,N_7346);
xor U7930 (N_7930,N_7342,N_6200);
nor U7931 (N_7931,N_7235,N_6631);
nand U7932 (N_7932,N_7153,N_6718);
nor U7933 (N_7933,N_6922,N_7005);
xor U7934 (N_7934,N_7414,N_6867);
and U7935 (N_7935,N_6628,N_6688);
xnor U7936 (N_7936,N_6153,N_7107);
nand U7937 (N_7937,N_7141,N_6350);
and U7938 (N_7938,N_7427,N_6329);
nor U7939 (N_7939,N_6124,N_6846);
xnor U7940 (N_7940,N_6387,N_7165);
nor U7941 (N_7941,N_6351,N_6665);
or U7942 (N_7942,N_6998,N_6568);
nand U7943 (N_7943,N_7291,N_6251);
or U7944 (N_7944,N_7252,N_7387);
or U7945 (N_7945,N_7158,N_6543);
xor U7946 (N_7946,N_7463,N_6242);
xnor U7947 (N_7947,N_6442,N_6600);
and U7948 (N_7948,N_7410,N_6240);
nor U7949 (N_7949,N_6614,N_7091);
or U7950 (N_7950,N_6530,N_6954);
xor U7951 (N_7951,N_7193,N_7137);
and U7952 (N_7952,N_6704,N_6071);
nand U7953 (N_7953,N_6607,N_6184);
nor U7954 (N_7954,N_6647,N_6824);
xnor U7955 (N_7955,N_6464,N_6879);
nand U7956 (N_7956,N_6357,N_7465);
and U7957 (N_7957,N_6634,N_6550);
and U7958 (N_7958,N_6971,N_7352);
nand U7959 (N_7959,N_7333,N_6635);
xor U7960 (N_7960,N_6905,N_7245);
xor U7961 (N_7961,N_6580,N_7150);
nor U7962 (N_7962,N_6806,N_7000);
and U7963 (N_7963,N_6029,N_7161);
nand U7964 (N_7964,N_6602,N_6937);
or U7965 (N_7965,N_6836,N_6130);
nor U7966 (N_7966,N_6669,N_7443);
or U7967 (N_7967,N_6945,N_7192);
nand U7968 (N_7968,N_7306,N_6245);
xnor U7969 (N_7969,N_7412,N_6233);
or U7970 (N_7970,N_6016,N_6326);
or U7971 (N_7971,N_7181,N_6649);
xnor U7972 (N_7972,N_6982,N_6599);
and U7973 (N_7973,N_7220,N_6460);
nor U7974 (N_7974,N_7239,N_7469);
nand U7975 (N_7975,N_6787,N_7156);
or U7976 (N_7976,N_6546,N_7372);
and U7977 (N_7977,N_7076,N_6008);
nor U7978 (N_7978,N_7230,N_6394);
nand U7979 (N_7979,N_6479,N_6136);
and U7980 (N_7980,N_6749,N_7310);
and U7981 (N_7981,N_6427,N_6850);
and U7982 (N_7982,N_7373,N_6049);
xnor U7983 (N_7983,N_6516,N_7126);
nand U7984 (N_7984,N_7083,N_6553);
or U7985 (N_7985,N_7467,N_7056);
or U7986 (N_7986,N_7064,N_6625);
xnor U7987 (N_7987,N_6990,N_7452);
nor U7988 (N_7988,N_6608,N_6074);
xor U7989 (N_7989,N_6735,N_7433);
xor U7990 (N_7990,N_6057,N_6068);
nand U7991 (N_7991,N_7062,N_7345);
nand U7992 (N_7992,N_7210,N_7055);
nand U7993 (N_7993,N_6572,N_7484);
nor U7994 (N_7994,N_6157,N_7237);
or U7995 (N_7995,N_6959,N_6435);
nor U7996 (N_7996,N_7315,N_6004);
or U7997 (N_7997,N_6084,N_6774);
and U7998 (N_7998,N_7307,N_6125);
or U7999 (N_7999,N_7272,N_6502);
nand U8000 (N_8000,N_6235,N_7328);
nor U8001 (N_8001,N_6539,N_7100);
nand U8002 (N_8002,N_6970,N_6369);
xor U8003 (N_8003,N_6054,N_6418);
and U8004 (N_8004,N_7189,N_7236);
nor U8005 (N_8005,N_6288,N_6244);
xor U8006 (N_8006,N_6481,N_7418);
or U8007 (N_8007,N_7059,N_6449);
or U8008 (N_8008,N_6999,N_6717);
nor U8009 (N_8009,N_7489,N_6795);
and U8010 (N_8010,N_6517,N_6652);
nand U8011 (N_8011,N_6848,N_7390);
or U8012 (N_8012,N_6757,N_7164);
nor U8013 (N_8013,N_6521,N_6391);
nand U8014 (N_8014,N_7178,N_7045);
and U8015 (N_8015,N_7391,N_6523);
nor U8016 (N_8016,N_6821,N_6457);
and U8017 (N_8017,N_7322,N_6415);
nor U8018 (N_8018,N_6173,N_6042);
and U8019 (N_8019,N_7313,N_6723);
and U8020 (N_8020,N_6582,N_6365);
nor U8021 (N_8021,N_6021,N_7121);
and U8022 (N_8022,N_6715,N_7249);
xor U8023 (N_8023,N_6545,N_6293);
and U8024 (N_8024,N_6651,N_6040);
nand U8025 (N_8025,N_6603,N_6392);
xor U8026 (N_8026,N_6212,N_6022);
xor U8027 (N_8027,N_6812,N_7057);
nor U8028 (N_8028,N_6310,N_6181);
xor U8029 (N_8029,N_6347,N_6342);
nor U8030 (N_8030,N_7377,N_6559);
nor U8031 (N_8031,N_6637,N_6320);
and U8032 (N_8032,N_7293,N_7296);
nor U8033 (N_8033,N_6034,N_7497);
nor U8034 (N_8034,N_7023,N_7294);
nand U8035 (N_8035,N_6984,N_6519);
xnor U8036 (N_8036,N_6063,N_7344);
or U8037 (N_8037,N_6230,N_6311);
and U8038 (N_8038,N_6064,N_6780);
nand U8039 (N_8039,N_6752,N_6977);
and U8040 (N_8040,N_6026,N_7116);
xnor U8041 (N_8041,N_7134,N_6209);
or U8042 (N_8042,N_7104,N_6041);
nor U8043 (N_8043,N_6593,N_7358);
and U8044 (N_8044,N_6551,N_6162);
xnor U8045 (N_8045,N_6032,N_6433);
nor U8046 (N_8046,N_6423,N_6370);
or U8047 (N_8047,N_6844,N_6114);
and U8048 (N_8048,N_7482,N_6743);
or U8049 (N_8049,N_7264,N_7167);
xor U8050 (N_8050,N_7122,N_7090);
xnor U8051 (N_8051,N_6707,N_6450);
nor U8052 (N_8052,N_7128,N_6962);
and U8053 (N_8053,N_6019,N_7017);
xor U8054 (N_8054,N_6224,N_6611);
xnor U8055 (N_8055,N_7223,N_6956);
or U8056 (N_8056,N_7424,N_6132);
or U8057 (N_8057,N_7302,N_6263);
or U8058 (N_8058,N_6921,N_7349);
nand U8059 (N_8059,N_7123,N_6158);
nor U8060 (N_8060,N_7067,N_6470);
and U8061 (N_8061,N_7204,N_6296);
xnor U8062 (N_8062,N_6980,N_6978);
xor U8063 (N_8063,N_6877,N_6270);
or U8064 (N_8064,N_7066,N_6996);
and U8065 (N_8065,N_6981,N_6898);
or U8066 (N_8066,N_6452,N_7019);
or U8067 (N_8067,N_7108,N_7092);
xnor U8068 (N_8068,N_6888,N_6748);
xnor U8069 (N_8069,N_6131,N_6201);
or U8070 (N_8070,N_6265,N_6498);
xor U8071 (N_8071,N_6766,N_6866);
nand U8072 (N_8072,N_6494,N_6443);
or U8073 (N_8073,N_6243,N_7376);
and U8074 (N_8074,N_7037,N_6128);
nor U8075 (N_8075,N_7305,N_7265);
xnor U8076 (N_8076,N_6023,N_7131);
nand U8077 (N_8077,N_6075,N_6384);
or U8078 (N_8078,N_6857,N_6499);
nor U8079 (N_8079,N_7214,N_6082);
nor U8080 (N_8080,N_6324,N_6855);
or U8081 (N_8081,N_6964,N_6152);
nand U8082 (N_8082,N_6936,N_7395);
nor U8083 (N_8083,N_7049,N_7013);
xor U8084 (N_8084,N_6646,N_6414);
and U8085 (N_8085,N_7275,N_6192);
or U8086 (N_8086,N_6058,N_7044);
or U8087 (N_8087,N_6389,N_6832);
and U8088 (N_8088,N_6947,N_7209);
and U8089 (N_8089,N_6547,N_6901);
nor U8090 (N_8090,N_7343,N_6248);
and U8091 (N_8091,N_6261,N_6283);
xor U8092 (N_8092,N_7098,N_6672);
or U8093 (N_8093,N_7276,N_6133);
xor U8094 (N_8094,N_6148,N_6809);
and U8095 (N_8095,N_7295,N_6826);
nor U8096 (N_8096,N_6883,N_6473);
xnor U8097 (N_8097,N_6897,N_7324);
and U8098 (N_8098,N_7389,N_6077);
and U8099 (N_8099,N_6127,N_6829);
and U8100 (N_8100,N_6010,N_6018);
or U8101 (N_8101,N_6556,N_6438);
and U8102 (N_8102,N_7081,N_6950);
xnor U8103 (N_8103,N_6196,N_7288);
and U8104 (N_8104,N_7403,N_6794);
nor U8105 (N_8105,N_6349,N_7426);
or U8106 (N_8106,N_7027,N_6705);
nand U8107 (N_8107,N_6810,N_7075);
or U8108 (N_8108,N_7254,N_6613);
nand U8109 (N_8109,N_6485,N_6563);
xnor U8110 (N_8110,N_6738,N_6755);
nor U8111 (N_8111,N_7365,N_7149);
nor U8112 (N_8112,N_7430,N_6946);
or U8113 (N_8113,N_6474,N_6226);
xor U8114 (N_8114,N_6280,N_6207);
and U8115 (N_8115,N_6737,N_6441);
and U8116 (N_8116,N_6446,N_7006);
and U8117 (N_8117,N_6861,N_7273);
and U8118 (N_8118,N_6432,N_6709);
xnor U8119 (N_8119,N_6841,N_6126);
nand U8120 (N_8120,N_6929,N_6252);
nand U8121 (N_8121,N_6772,N_7173);
or U8122 (N_8122,N_6797,N_6274);
nor U8123 (N_8123,N_6609,N_7444);
nand U8124 (N_8124,N_6736,N_6756);
nor U8125 (N_8125,N_6864,N_6101);
nand U8126 (N_8126,N_7429,N_6807);
xor U8127 (N_8127,N_6501,N_6655);
xnor U8128 (N_8128,N_7449,N_7460);
and U8129 (N_8129,N_6031,N_6658);
xnor U8130 (N_8130,N_6819,N_6172);
xor U8131 (N_8131,N_7268,N_7471);
and U8132 (N_8132,N_7082,N_6259);
or U8133 (N_8133,N_6654,N_7242);
or U8134 (N_8134,N_7494,N_6319);
and U8135 (N_8135,N_6610,N_6399);
and U8136 (N_8136,N_6374,N_7170);
and U8137 (N_8137,N_7255,N_6703);
nor U8138 (N_8138,N_6228,N_6445);
nor U8139 (N_8139,N_6884,N_6661);
or U8140 (N_8140,N_7177,N_6378);
and U8141 (N_8141,N_7207,N_6380);
or U8142 (N_8142,N_6100,N_7202);
xor U8143 (N_8143,N_6053,N_7488);
nand U8144 (N_8144,N_7356,N_6803);
nor U8145 (N_8145,N_6458,N_7396);
and U8146 (N_8146,N_6548,N_6627);
nor U8147 (N_8147,N_7402,N_6983);
nor U8148 (N_8148,N_6408,N_6046);
xnor U8149 (N_8149,N_7474,N_6269);
nor U8150 (N_8150,N_6146,N_7071);
xnor U8151 (N_8151,N_6006,N_6562);
and U8152 (N_8152,N_7388,N_6938);
xnor U8153 (N_8153,N_7321,N_7004);
nor U8154 (N_8154,N_6833,N_7394);
nor U8155 (N_8155,N_6816,N_6881);
xor U8156 (N_8156,N_7278,N_6919);
xor U8157 (N_8157,N_6366,N_7440);
xnor U8158 (N_8158,N_6353,N_6355);
and U8159 (N_8159,N_6727,N_6469);
xor U8160 (N_8160,N_6719,N_6961);
nor U8161 (N_8161,N_7200,N_7423);
nand U8162 (N_8162,N_6051,N_6246);
and U8163 (N_8163,N_6720,N_7283);
nand U8164 (N_8164,N_6216,N_6615);
or U8165 (N_8165,N_6671,N_6098);
nand U8166 (N_8166,N_6134,N_6417);
or U8167 (N_8167,N_6012,N_6121);
or U8168 (N_8168,N_6397,N_7382);
and U8169 (N_8169,N_6567,N_7155);
and U8170 (N_8170,N_7152,N_6716);
nand U8171 (N_8171,N_6352,N_6303);
xnor U8172 (N_8172,N_7127,N_6633);
or U8173 (N_8173,N_6747,N_6900);
xnor U8174 (N_8174,N_7033,N_6623);
nor U8175 (N_8175,N_6638,N_6017);
nand U8176 (N_8176,N_6570,N_6434);
and U8177 (N_8177,N_7112,N_7490);
xnor U8178 (N_8178,N_6379,N_6437);
or U8179 (N_8179,N_6312,N_7300);
nand U8180 (N_8180,N_6220,N_7186);
nand U8181 (N_8181,N_6713,N_6316);
xor U8182 (N_8182,N_7407,N_6083);
xor U8183 (N_8183,N_6690,N_6362);
xnor U8184 (N_8184,N_6487,N_6390);
nor U8185 (N_8185,N_6840,N_6781);
nor U8186 (N_8186,N_6528,N_6642);
or U8187 (N_8187,N_6698,N_6388);
nand U8188 (N_8188,N_6356,N_6696);
xor U8189 (N_8189,N_7421,N_6139);
nor U8190 (N_8190,N_6299,N_6413);
nand U8191 (N_8191,N_6910,N_6095);
nand U8192 (N_8192,N_7492,N_6304);
and U8193 (N_8193,N_6340,N_7054);
xnor U8194 (N_8194,N_6683,N_6337);
xor U8195 (N_8195,N_6986,N_7406);
and U8196 (N_8196,N_6191,N_6581);
nand U8197 (N_8197,N_6108,N_6236);
nand U8198 (N_8198,N_6141,N_6105);
nor U8199 (N_8199,N_6383,N_6892);
xor U8200 (N_8200,N_6762,N_6925);
nand U8201 (N_8201,N_6094,N_7416);
xnor U8202 (N_8202,N_6182,N_6455);
nand U8203 (N_8203,N_6496,N_6331);
and U8204 (N_8204,N_6507,N_6791);
nor U8205 (N_8205,N_7136,N_6590);
nand U8206 (N_8206,N_6215,N_6047);
nand U8207 (N_8207,N_6313,N_6798);
and U8208 (N_8208,N_6286,N_6363);
nand U8209 (N_8209,N_7371,N_6694);
nand U8210 (N_8210,N_6099,N_6467);
and U8211 (N_8211,N_7052,N_6285);
xnor U8212 (N_8212,N_7041,N_6147);
and U8213 (N_8213,N_6361,N_6278);
and U8214 (N_8214,N_6462,N_7205);
or U8215 (N_8215,N_6508,N_7226);
xor U8216 (N_8216,N_6566,N_7461);
nand U8217 (N_8217,N_6656,N_6056);
nand U8218 (N_8218,N_6728,N_6221);
nor U8219 (N_8219,N_6536,N_7290);
nor U8220 (N_8220,N_7339,N_7036);
xnor U8221 (N_8221,N_6712,N_7266);
nand U8222 (N_8222,N_6874,N_7061);
xnor U8223 (N_8223,N_7133,N_6290);
and U8224 (N_8224,N_7260,N_6500);
nor U8225 (N_8225,N_6949,N_7138);
nor U8226 (N_8226,N_7454,N_6972);
nand U8227 (N_8227,N_6333,N_6740);
or U8228 (N_8228,N_6112,N_6475);
nor U8229 (N_8229,N_6306,N_7475);
nand U8230 (N_8230,N_7456,N_6558);
or U8231 (N_8231,N_6461,N_6699);
nor U8232 (N_8232,N_6440,N_6381);
and U8233 (N_8233,N_6490,N_7197);
xor U8234 (N_8234,N_7270,N_6277);
nand U8235 (N_8235,N_6677,N_6960);
nor U8236 (N_8236,N_6838,N_6317);
and U8237 (N_8237,N_7248,N_6309);
nor U8238 (N_8238,N_6605,N_7007);
nor U8239 (N_8239,N_6214,N_7439);
and U8240 (N_8240,N_6364,N_6760);
or U8241 (N_8241,N_6227,N_6003);
and U8242 (N_8242,N_6066,N_6431);
nor U8243 (N_8243,N_7103,N_6161);
or U8244 (N_8244,N_6882,N_6584);
xor U8245 (N_8245,N_6880,N_6595);
xor U8246 (N_8246,N_6931,N_7404);
and U8247 (N_8247,N_6279,N_6682);
xnor U8248 (N_8248,N_6421,N_6588);
nand U8249 (N_8249,N_6150,N_7485);
xnor U8250 (N_8250,N_7307,N_6502);
xor U8251 (N_8251,N_6502,N_6569);
nand U8252 (N_8252,N_6780,N_6856);
or U8253 (N_8253,N_6553,N_6419);
nand U8254 (N_8254,N_6078,N_6120);
or U8255 (N_8255,N_6767,N_6732);
or U8256 (N_8256,N_7453,N_6526);
nand U8257 (N_8257,N_6061,N_7303);
and U8258 (N_8258,N_6057,N_6148);
nand U8259 (N_8259,N_6587,N_6090);
or U8260 (N_8260,N_7259,N_7492);
nor U8261 (N_8261,N_6259,N_6821);
or U8262 (N_8262,N_7314,N_6708);
and U8263 (N_8263,N_6986,N_6911);
xnor U8264 (N_8264,N_6839,N_7139);
and U8265 (N_8265,N_7129,N_6752);
xnor U8266 (N_8266,N_6091,N_7417);
and U8267 (N_8267,N_6155,N_6203);
nand U8268 (N_8268,N_6606,N_6597);
xnor U8269 (N_8269,N_6478,N_7094);
nand U8270 (N_8270,N_7251,N_6548);
nand U8271 (N_8271,N_6792,N_7056);
nand U8272 (N_8272,N_7373,N_7113);
or U8273 (N_8273,N_6801,N_6236);
nor U8274 (N_8274,N_7100,N_6336);
and U8275 (N_8275,N_7101,N_7468);
and U8276 (N_8276,N_6182,N_7409);
nand U8277 (N_8277,N_6823,N_7050);
or U8278 (N_8278,N_6487,N_7006);
nor U8279 (N_8279,N_6532,N_7465);
nand U8280 (N_8280,N_6869,N_7438);
nand U8281 (N_8281,N_7165,N_6366);
nand U8282 (N_8282,N_7102,N_7307);
xnor U8283 (N_8283,N_6570,N_6580);
xnor U8284 (N_8284,N_6860,N_6974);
nor U8285 (N_8285,N_6819,N_6121);
and U8286 (N_8286,N_7047,N_6260);
or U8287 (N_8287,N_6018,N_6254);
xnor U8288 (N_8288,N_7011,N_6864);
nor U8289 (N_8289,N_6318,N_6047);
nand U8290 (N_8290,N_6263,N_6732);
nand U8291 (N_8291,N_6598,N_7022);
or U8292 (N_8292,N_7367,N_6004);
nand U8293 (N_8293,N_6832,N_6012);
xnor U8294 (N_8294,N_7292,N_6849);
xor U8295 (N_8295,N_6859,N_7020);
nand U8296 (N_8296,N_6133,N_6844);
and U8297 (N_8297,N_6247,N_6026);
and U8298 (N_8298,N_6517,N_6740);
or U8299 (N_8299,N_6767,N_6200);
xor U8300 (N_8300,N_6400,N_7246);
or U8301 (N_8301,N_7415,N_6122);
or U8302 (N_8302,N_6524,N_6319);
nor U8303 (N_8303,N_6127,N_6482);
nor U8304 (N_8304,N_7486,N_6103);
nor U8305 (N_8305,N_7399,N_6186);
nor U8306 (N_8306,N_7125,N_7438);
nand U8307 (N_8307,N_6466,N_6662);
nand U8308 (N_8308,N_6925,N_6291);
nand U8309 (N_8309,N_7073,N_7381);
nor U8310 (N_8310,N_6997,N_7474);
xor U8311 (N_8311,N_7301,N_7477);
xor U8312 (N_8312,N_6541,N_7363);
and U8313 (N_8313,N_7493,N_6918);
nor U8314 (N_8314,N_6426,N_6676);
nor U8315 (N_8315,N_6032,N_7173);
or U8316 (N_8316,N_6250,N_7182);
or U8317 (N_8317,N_6129,N_6056);
nand U8318 (N_8318,N_6153,N_6114);
xnor U8319 (N_8319,N_7114,N_7077);
nor U8320 (N_8320,N_7351,N_6711);
or U8321 (N_8321,N_7237,N_7124);
and U8322 (N_8322,N_6230,N_6468);
nand U8323 (N_8323,N_6714,N_6657);
or U8324 (N_8324,N_7387,N_6081);
nand U8325 (N_8325,N_6917,N_7262);
xnor U8326 (N_8326,N_6794,N_6714);
and U8327 (N_8327,N_7206,N_6562);
xnor U8328 (N_8328,N_6387,N_6505);
and U8329 (N_8329,N_6938,N_6468);
nand U8330 (N_8330,N_6913,N_6546);
and U8331 (N_8331,N_7086,N_6473);
nand U8332 (N_8332,N_6425,N_6182);
or U8333 (N_8333,N_6818,N_6133);
xor U8334 (N_8334,N_7413,N_6703);
and U8335 (N_8335,N_6989,N_6355);
xnor U8336 (N_8336,N_6251,N_6313);
nand U8337 (N_8337,N_6583,N_6525);
nand U8338 (N_8338,N_6494,N_7092);
nand U8339 (N_8339,N_7282,N_6223);
nor U8340 (N_8340,N_6581,N_6585);
nand U8341 (N_8341,N_7372,N_6051);
xnor U8342 (N_8342,N_6417,N_6196);
nor U8343 (N_8343,N_7228,N_6771);
xor U8344 (N_8344,N_6145,N_6293);
nand U8345 (N_8345,N_6267,N_6125);
nor U8346 (N_8346,N_6249,N_7112);
xnor U8347 (N_8347,N_6585,N_7135);
or U8348 (N_8348,N_6223,N_7071);
nand U8349 (N_8349,N_6416,N_7018);
nor U8350 (N_8350,N_6531,N_7309);
nand U8351 (N_8351,N_6915,N_6436);
nand U8352 (N_8352,N_6845,N_6952);
nand U8353 (N_8353,N_7133,N_6585);
nor U8354 (N_8354,N_7356,N_6762);
xor U8355 (N_8355,N_6587,N_7099);
and U8356 (N_8356,N_6280,N_6122);
nor U8357 (N_8357,N_7433,N_6148);
and U8358 (N_8358,N_7472,N_6139);
nor U8359 (N_8359,N_7139,N_6453);
xnor U8360 (N_8360,N_6251,N_6787);
xnor U8361 (N_8361,N_6071,N_7201);
and U8362 (N_8362,N_6743,N_6220);
and U8363 (N_8363,N_6484,N_6490);
nand U8364 (N_8364,N_6673,N_7166);
nand U8365 (N_8365,N_7145,N_6068);
nand U8366 (N_8366,N_7139,N_7370);
nor U8367 (N_8367,N_6225,N_6055);
nand U8368 (N_8368,N_6331,N_7300);
and U8369 (N_8369,N_7494,N_7413);
nor U8370 (N_8370,N_6145,N_6398);
or U8371 (N_8371,N_7345,N_6316);
nand U8372 (N_8372,N_6005,N_6453);
or U8373 (N_8373,N_6175,N_6993);
and U8374 (N_8374,N_7156,N_6700);
nor U8375 (N_8375,N_7291,N_6315);
xor U8376 (N_8376,N_7434,N_6057);
or U8377 (N_8377,N_7375,N_6547);
or U8378 (N_8378,N_7026,N_6532);
and U8379 (N_8379,N_6039,N_6584);
or U8380 (N_8380,N_6165,N_7180);
and U8381 (N_8381,N_7234,N_6551);
nor U8382 (N_8382,N_7448,N_6937);
and U8383 (N_8383,N_7193,N_6601);
nand U8384 (N_8384,N_6048,N_6101);
or U8385 (N_8385,N_6979,N_6573);
and U8386 (N_8386,N_7071,N_7401);
nor U8387 (N_8387,N_7492,N_6257);
nor U8388 (N_8388,N_7169,N_6124);
nand U8389 (N_8389,N_6727,N_6872);
nand U8390 (N_8390,N_6442,N_6559);
or U8391 (N_8391,N_7069,N_6422);
and U8392 (N_8392,N_6149,N_6122);
and U8393 (N_8393,N_6473,N_7167);
or U8394 (N_8394,N_7346,N_6382);
xnor U8395 (N_8395,N_7295,N_6768);
nand U8396 (N_8396,N_7494,N_6998);
or U8397 (N_8397,N_6171,N_7241);
and U8398 (N_8398,N_7470,N_6327);
nor U8399 (N_8399,N_6471,N_6650);
or U8400 (N_8400,N_6213,N_7183);
nor U8401 (N_8401,N_6304,N_7208);
and U8402 (N_8402,N_6649,N_7249);
xor U8403 (N_8403,N_7323,N_6027);
or U8404 (N_8404,N_6507,N_6018);
or U8405 (N_8405,N_6486,N_6675);
nor U8406 (N_8406,N_7365,N_7162);
and U8407 (N_8407,N_6259,N_6075);
nand U8408 (N_8408,N_6751,N_6259);
nor U8409 (N_8409,N_7070,N_6850);
xnor U8410 (N_8410,N_7325,N_6853);
and U8411 (N_8411,N_6175,N_6482);
xor U8412 (N_8412,N_6601,N_6490);
xnor U8413 (N_8413,N_6227,N_6428);
nor U8414 (N_8414,N_6889,N_6386);
nand U8415 (N_8415,N_6870,N_6069);
xnor U8416 (N_8416,N_6898,N_6042);
nor U8417 (N_8417,N_6757,N_6242);
nor U8418 (N_8418,N_6042,N_6940);
xor U8419 (N_8419,N_6957,N_6613);
and U8420 (N_8420,N_6779,N_6143);
and U8421 (N_8421,N_6407,N_6420);
and U8422 (N_8422,N_6656,N_6904);
xor U8423 (N_8423,N_6439,N_7311);
xor U8424 (N_8424,N_6154,N_6099);
nand U8425 (N_8425,N_6046,N_6933);
nand U8426 (N_8426,N_6390,N_6526);
nand U8427 (N_8427,N_6232,N_7208);
xor U8428 (N_8428,N_6819,N_6663);
nand U8429 (N_8429,N_7382,N_6477);
nand U8430 (N_8430,N_6074,N_6639);
nor U8431 (N_8431,N_6747,N_7131);
xnor U8432 (N_8432,N_6170,N_7452);
or U8433 (N_8433,N_6212,N_6335);
xor U8434 (N_8434,N_6962,N_6907);
or U8435 (N_8435,N_7411,N_7195);
nand U8436 (N_8436,N_6866,N_7131);
nor U8437 (N_8437,N_7056,N_7211);
nand U8438 (N_8438,N_6298,N_6626);
and U8439 (N_8439,N_7201,N_6104);
xor U8440 (N_8440,N_7294,N_6658);
xor U8441 (N_8441,N_6009,N_7328);
nand U8442 (N_8442,N_7259,N_7019);
or U8443 (N_8443,N_6047,N_6688);
xor U8444 (N_8444,N_7009,N_6009);
nor U8445 (N_8445,N_7478,N_7327);
nor U8446 (N_8446,N_6280,N_6431);
xnor U8447 (N_8447,N_6591,N_6233);
and U8448 (N_8448,N_6870,N_6841);
nand U8449 (N_8449,N_7122,N_7284);
xnor U8450 (N_8450,N_6431,N_6864);
or U8451 (N_8451,N_7201,N_7360);
nor U8452 (N_8452,N_6591,N_7077);
nor U8453 (N_8453,N_6643,N_6384);
and U8454 (N_8454,N_6062,N_6348);
and U8455 (N_8455,N_7392,N_6586);
nand U8456 (N_8456,N_6701,N_6950);
nand U8457 (N_8457,N_6251,N_6200);
xnor U8458 (N_8458,N_7488,N_7453);
nor U8459 (N_8459,N_7044,N_6077);
or U8460 (N_8460,N_6177,N_7122);
nor U8461 (N_8461,N_6339,N_6736);
nor U8462 (N_8462,N_7157,N_7479);
nand U8463 (N_8463,N_7042,N_7122);
nand U8464 (N_8464,N_6850,N_6202);
nor U8465 (N_8465,N_6574,N_7025);
and U8466 (N_8466,N_6326,N_7458);
and U8467 (N_8467,N_7025,N_6577);
nor U8468 (N_8468,N_6443,N_6041);
nand U8469 (N_8469,N_6528,N_6178);
or U8470 (N_8470,N_6802,N_6707);
nand U8471 (N_8471,N_6461,N_7029);
nand U8472 (N_8472,N_6756,N_6459);
xnor U8473 (N_8473,N_7006,N_7174);
nand U8474 (N_8474,N_6272,N_6750);
or U8475 (N_8475,N_6205,N_7364);
xnor U8476 (N_8476,N_7113,N_7201);
nor U8477 (N_8477,N_6448,N_6021);
and U8478 (N_8478,N_6490,N_6858);
or U8479 (N_8479,N_6531,N_6479);
nand U8480 (N_8480,N_7274,N_6753);
or U8481 (N_8481,N_7425,N_6447);
and U8482 (N_8482,N_7250,N_7004);
nor U8483 (N_8483,N_6044,N_7416);
or U8484 (N_8484,N_6586,N_7121);
or U8485 (N_8485,N_6220,N_6978);
xnor U8486 (N_8486,N_6450,N_6115);
nand U8487 (N_8487,N_7245,N_6770);
and U8488 (N_8488,N_6634,N_6256);
nor U8489 (N_8489,N_6387,N_6668);
and U8490 (N_8490,N_6998,N_6925);
and U8491 (N_8491,N_6882,N_7165);
xnor U8492 (N_8492,N_6924,N_6516);
or U8493 (N_8493,N_7495,N_6668);
and U8494 (N_8494,N_6768,N_7100);
nor U8495 (N_8495,N_7027,N_7099);
or U8496 (N_8496,N_6341,N_6786);
nor U8497 (N_8497,N_7464,N_7471);
nand U8498 (N_8498,N_6879,N_6674);
or U8499 (N_8499,N_6695,N_6429);
nor U8500 (N_8500,N_6588,N_7334);
or U8501 (N_8501,N_7493,N_6356);
xnor U8502 (N_8502,N_7110,N_6155);
or U8503 (N_8503,N_6397,N_7409);
or U8504 (N_8504,N_6304,N_6646);
nor U8505 (N_8505,N_6964,N_6802);
and U8506 (N_8506,N_6960,N_6066);
nand U8507 (N_8507,N_6300,N_6273);
nor U8508 (N_8508,N_7069,N_6523);
or U8509 (N_8509,N_6273,N_6680);
nand U8510 (N_8510,N_6308,N_6078);
nand U8511 (N_8511,N_6153,N_7407);
or U8512 (N_8512,N_6305,N_6724);
nor U8513 (N_8513,N_7291,N_7090);
nand U8514 (N_8514,N_7299,N_7355);
nand U8515 (N_8515,N_6987,N_7162);
and U8516 (N_8516,N_6299,N_6755);
and U8517 (N_8517,N_6537,N_6004);
or U8518 (N_8518,N_7217,N_7249);
nand U8519 (N_8519,N_7300,N_6063);
nor U8520 (N_8520,N_7139,N_6405);
and U8521 (N_8521,N_7139,N_6257);
nor U8522 (N_8522,N_7350,N_7154);
or U8523 (N_8523,N_6707,N_6071);
xnor U8524 (N_8524,N_6468,N_6113);
nand U8525 (N_8525,N_7198,N_7113);
nand U8526 (N_8526,N_7063,N_6657);
or U8527 (N_8527,N_6355,N_6348);
xor U8528 (N_8528,N_7430,N_6327);
or U8529 (N_8529,N_6963,N_7294);
and U8530 (N_8530,N_7442,N_6190);
or U8531 (N_8531,N_6159,N_7202);
xnor U8532 (N_8532,N_7224,N_6037);
or U8533 (N_8533,N_6570,N_7034);
and U8534 (N_8534,N_6996,N_7478);
or U8535 (N_8535,N_7337,N_7414);
nand U8536 (N_8536,N_6324,N_7185);
xor U8537 (N_8537,N_6175,N_7149);
nor U8538 (N_8538,N_6037,N_6675);
nand U8539 (N_8539,N_6489,N_6799);
xnor U8540 (N_8540,N_7465,N_6855);
nor U8541 (N_8541,N_6505,N_6961);
or U8542 (N_8542,N_6261,N_7074);
nand U8543 (N_8543,N_6752,N_6571);
nor U8544 (N_8544,N_6093,N_6779);
or U8545 (N_8545,N_7170,N_7273);
nor U8546 (N_8546,N_6195,N_6103);
xnor U8547 (N_8547,N_7135,N_6943);
or U8548 (N_8548,N_6453,N_6578);
nor U8549 (N_8549,N_6438,N_6344);
nand U8550 (N_8550,N_6291,N_6897);
nand U8551 (N_8551,N_6989,N_6814);
nand U8552 (N_8552,N_7243,N_7372);
or U8553 (N_8553,N_6778,N_6024);
nand U8554 (N_8554,N_6970,N_7123);
nand U8555 (N_8555,N_6176,N_6914);
nor U8556 (N_8556,N_6059,N_7048);
xnor U8557 (N_8557,N_7275,N_6561);
or U8558 (N_8558,N_6025,N_6934);
nor U8559 (N_8559,N_6506,N_6844);
and U8560 (N_8560,N_6797,N_6612);
and U8561 (N_8561,N_6110,N_7436);
xnor U8562 (N_8562,N_7400,N_7114);
and U8563 (N_8563,N_6910,N_6584);
or U8564 (N_8564,N_6777,N_6643);
nor U8565 (N_8565,N_6462,N_6496);
and U8566 (N_8566,N_6242,N_6150);
nand U8567 (N_8567,N_7098,N_6448);
nand U8568 (N_8568,N_7258,N_7421);
xor U8569 (N_8569,N_6956,N_6734);
or U8570 (N_8570,N_6957,N_6886);
xnor U8571 (N_8571,N_6120,N_6880);
nand U8572 (N_8572,N_6074,N_6317);
xnor U8573 (N_8573,N_6088,N_6595);
and U8574 (N_8574,N_6407,N_6156);
and U8575 (N_8575,N_6066,N_7149);
and U8576 (N_8576,N_6381,N_6375);
and U8577 (N_8577,N_7193,N_6370);
nand U8578 (N_8578,N_6044,N_6460);
or U8579 (N_8579,N_6900,N_6037);
and U8580 (N_8580,N_6794,N_6207);
nor U8581 (N_8581,N_6960,N_7345);
and U8582 (N_8582,N_6078,N_6977);
nand U8583 (N_8583,N_6178,N_7407);
and U8584 (N_8584,N_6169,N_6447);
or U8585 (N_8585,N_7309,N_7371);
xnor U8586 (N_8586,N_6102,N_6909);
nand U8587 (N_8587,N_6175,N_6846);
and U8588 (N_8588,N_7457,N_6132);
and U8589 (N_8589,N_6151,N_6725);
nand U8590 (N_8590,N_7131,N_7493);
and U8591 (N_8591,N_6418,N_6715);
or U8592 (N_8592,N_6646,N_6645);
and U8593 (N_8593,N_6810,N_7213);
nor U8594 (N_8594,N_7197,N_7188);
or U8595 (N_8595,N_6161,N_7071);
or U8596 (N_8596,N_6116,N_7220);
nor U8597 (N_8597,N_6941,N_6475);
nor U8598 (N_8598,N_6802,N_6539);
nor U8599 (N_8599,N_6062,N_6360);
nor U8600 (N_8600,N_7344,N_7198);
xor U8601 (N_8601,N_7370,N_7400);
and U8602 (N_8602,N_6970,N_6338);
nand U8603 (N_8603,N_7457,N_6377);
nand U8604 (N_8604,N_6243,N_7420);
or U8605 (N_8605,N_6635,N_7377);
nor U8606 (N_8606,N_6822,N_7195);
or U8607 (N_8607,N_6167,N_6232);
and U8608 (N_8608,N_6072,N_7002);
and U8609 (N_8609,N_6738,N_6490);
nand U8610 (N_8610,N_6375,N_7003);
or U8611 (N_8611,N_7242,N_6506);
nand U8612 (N_8612,N_6766,N_6030);
or U8613 (N_8613,N_6878,N_7098);
nand U8614 (N_8614,N_7406,N_7296);
and U8615 (N_8615,N_6929,N_7221);
xnor U8616 (N_8616,N_6207,N_6896);
xnor U8617 (N_8617,N_6845,N_6442);
and U8618 (N_8618,N_7160,N_6648);
nand U8619 (N_8619,N_6416,N_6141);
or U8620 (N_8620,N_7211,N_6024);
or U8621 (N_8621,N_7141,N_6616);
nand U8622 (N_8622,N_6312,N_6958);
nor U8623 (N_8623,N_6248,N_6110);
or U8624 (N_8624,N_6830,N_7125);
xor U8625 (N_8625,N_6526,N_6373);
xor U8626 (N_8626,N_7234,N_6460);
or U8627 (N_8627,N_7469,N_7236);
xor U8628 (N_8628,N_7463,N_7115);
and U8629 (N_8629,N_6978,N_6519);
or U8630 (N_8630,N_6383,N_7259);
nor U8631 (N_8631,N_7250,N_7434);
and U8632 (N_8632,N_7430,N_6398);
nor U8633 (N_8633,N_6019,N_7183);
and U8634 (N_8634,N_7322,N_7284);
and U8635 (N_8635,N_6055,N_6703);
nand U8636 (N_8636,N_6749,N_6569);
nor U8637 (N_8637,N_6740,N_6099);
and U8638 (N_8638,N_6645,N_7257);
xnor U8639 (N_8639,N_6454,N_7225);
and U8640 (N_8640,N_6249,N_6575);
and U8641 (N_8641,N_7097,N_6771);
xor U8642 (N_8642,N_6638,N_6548);
or U8643 (N_8643,N_6066,N_6894);
xnor U8644 (N_8644,N_7280,N_6896);
or U8645 (N_8645,N_6910,N_7313);
and U8646 (N_8646,N_7379,N_6751);
and U8647 (N_8647,N_6010,N_7452);
nand U8648 (N_8648,N_6966,N_6610);
xor U8649 (N_8649,N_6014,N_6800);
nor U8650 (N_8650,N_6205,N_6400);
or U8651 (N_8651,N_6391,N_6166);
xor U8652 (N_8652,N_6889,N_6939);
and U8653 (N_8653,N_7358,N_6007);
or U8654 (N_8654,N_6135,N_6264);
or U8655 (N_8655,N_6738,N_7089);
nand U8656 (N_8656,N_6485,N_6408);
nor U8657 (N_8657,N_6712,N_6874);
xor U8658 (N_8658,N_7192,N_7459);
and U8659 (N_8659,N_7143,N_7294);
or U8660 (N_8660,N_7325,N_6522);
and U8661 (N_8661,N_6764,N_7104);
or U8662 (N_8662,N_7162,N_6593);
nor U8663 (N_8663,N_6974,N_6640);
xor U8664 (N_8664,N_6953,N_6011);
and U8665 (N_8665,N_7411,N_7491);
nand U8666 (N_8666,N_6146,N_6827);
and U8667 (N_8667,N_7040,N_7411);
xnor U8668 (N_8668,N_6578,N_7023);
nor U8669 (N_8669,N_7119,N_6344);
and U8670 (N_8670,N_6162,N_7224);
and U8671 (N_8671,N_6339,N_7449);
nand U8672 (N_8672,N_6666,N_6413);
and U8673 (N_8673,N_7272,N_6404);
nor U8674 (N_8674,N_6105,N_7209);
xnor U8675 (N_8675,N_7130,N_6024);
xnor U8676 (N_8676,N_7395,N_6356);
nor U8677 (N_8677,N_6511,N_6144);
or U8678 (N_8678,N_6954,N_6302);
or U8679 (N_8679,N_7349,N_6965);
nand U8680 (N_8680,N_6452,N_6710);
xor U8681 (N_8681,N_6501,N_6596);
and U8682 (N_8682,N_6396,N_7344);
or U8683 (N_8683,N_6237,N_6469);
or U8684 (N_8684,N_6326,N_7058);
or U8685 (N_8685,N_6600,N_6225);
xnor U8686 (N_8686,N_7442,N_7036);
nor U8687 (N_8687,N_6570,N_6210);
nor U8688 (N_8688,N_6818,N_6838);
or U8689 (N_8689,N_6947,N_7159);
xor U8690 (N_8690,N_6026,N_6542);
or U8691 (N_8691,N_7454,N_6450);
xor U8692 (N_8692,N_7448,N_6112);
or U8693 (N_8693,N_7417,N_6687);
nor U8694 (N_8694,N_7357,N_6888);
or U8695 (N_8695,N_6333,N_6279);
nor U8696 (N_8696,N_6596,N_6927);
nor U8697 (N_8697,N_6716,N_6384);
xnor U8698 (N_8698,N_7464,N_6252);
nand U8699 (N_8699,N_7469,N_7308);
nor U8700 (N_8700,N_7108,N_6607);
or U8701 (N_8701,N_7453,N_6910);
or U8702 (N_8702,N_6058,N_7012);
nand U8703 (N_8703,N_7200,N_6143);
nor U8704 (N_8704,N_6184,N_6145);
xnor U8705 (N_8705,N_7459,N_7219);
or U8706 (N_8706,N_7078,N_7228);
or U8707 (N_8707,N_6071,N_6246);
or U8708 (N_8708,N_7474,N_6927);
nand U8709 (N_8709,N_6107,N_6484);
xor U8710 (N_8710,N_7456,N_6451);
or U8711 (N_8711,N_7048,N_6536);
xnor U8712 (N_8712,N_6922,N_7031);
nor U8713 (N_8713,N_6039,N_6838);
xor U8714 (N_8714,N_6121,N_6417);
nor U8715 (N_8715,N_7455,N_6457);
and U8716 (N_8716,N_6213,N_6827);
xor U8717 (N_8717,N_6960,N_7464);
xnor U8718 (N_8718,N_7350,N_6660);
nand U8719 (N_8719,N_7155,N_7051);
nor U8720 (N_8720,N_6227,N_7110);
nand U8721 (N_8721,N_6161,N_6921);
nand U8722 (N_8722,N_7145,N_6407);
nor U8723 (N_8723,N_7300,N_6240);
nand U8724 (N_8724,N_6329,N_6768);
and U8725 (N_8725,N_7155,N_6315);
xnor U8726 (N_8726,N_6781,N_6902);
or U8727 (N_8727,N_6204,N_6449);
and U8728 (N_8728,N_6413,N_6460);
and U8729 (N_8729,N_7144,N_6193);
xor U8730 (N_8730,N_7026,N_7126);
xnor U8731 (N_8731,N_7333,N_6940);
or U8732 (N_8732,N_6150,N_7492);
or U8733 (N_8733,N_6482,N_6274);
nand U8734 (N_8734,N_7101,N_6928);
and U8735 (N_8735,N_6298,N_6313);
nand U8736 (N_8736,N_6650,N_6998);
nor U8737 (N_8737,N_6474,N_6572);
xor U8738 (N_8738,N_7008,N_6806);
xor U8739 (N_8739,N_7372,N_6657);
or U8740 (N_8740,N_6282,N_7013);
or U8741 (N_8741,N_6694,N_6380);
xnor U8742 (N_8742,N_6010,N_6852);
nor U8743 (N_8743,N_6707,N_6634);
nor U8744 (N_8744,N_6219,N_7129);
xor U8745 (N_8745,N_6462,N_7301);
nand U8746 (N_8746,N_6331,N_6420);
or U8747 (N_8747,N_6380,N_6967);
or U8748 (N_8748,N_6068,N_7000);
and U8749 (N_8749,N_7360,N_7291);
nor U8750 (N_8750,N_7117,N_6859);
xnor U8751 (N_8751,N_7201,N_6470);
nor U8752 (N_8752,N_7122,N_6644);
xnor U8753 (N_8753,N_6300,N_7272);
nand U8754 (N_8754,N_7320,N_6091);
nor U8755 (N_8755,N_6241,N_6949);
xor U8756 (N_8756,N_6274,N_6430);
nand U8757 (N_8757,N_6529,N_6080);
nor U8758 (N_8758,N_6113,N_6675);
or U8759 (N_8759,N_6379,N_6002);
xnor U8760 (N_8760,N_7437,N_6687);
xor U8761 (N_8761,N_6497,N_6978);
nor U8762 (N_8762,N_6764,N_7179);
and U8763 (N_8763,N_6767,N_6786);
nand U8764 (N_8764,N_6659,N_6389);
and U8765 (N_8765,N_6281,N_6975);
xor U8766 (N_8766,N_6880,N_6969);
nor U8767 (N_8767,N_7112,N_6964);
and U8768 (N_8768,N_7429,N_6489);
and U8769 (N_8769,N_6442,N_7280);
nor U8770 (N_8770,N_6385,N_6870);
or U8771 (N_8771,N_7469,N_6616);
or U8772 (N_8772,N_6196,N_6623);
nor U8773 (N_8773,N_6122,N_6068);
xnor U8774 (N_8774,N_7236,N_6382);
nor U8775 (N_8775,N_6970,N_6528);
and U8776 (N_8776,N_6736,N_7447);
nor U8777 (N_8777,N_7193,N_6691);
xnor U8778 (N_8778,N_6080,N_6629);
and U8779 (N_8779,N_7185,N_6959);
nand U8780 (N_8780,N_7327,N_6133);
xnor U8781 (N_8781,N_6714,N_6973);
nand U8782 (N_8782,N_6755,N_6133);
nor U8783 (N_8783,N_6643,N_6337);
xor U8784 (N_8784,N_7403,N_6361);
xor U8785 (N_8785,N_6963,N_6734);
nand U8786 (N_8786,N_6882,N_7181);
and U8787 (N_8787,N_6960,N_6742);
and U8788 (N_8788,N_6317,N_7009);
and U8789 (N_8789,N_6214,N_6125);
nor U8790 (N_8790,N_7240,N_7351);
and U8791 (N_8791,N_7149,N_6872);
xnor U8792 (N_8792,N_7385,N_7065);
nand U8793 (N_8793,N_6531,N_6776);
and U8794 (N_8794,N_6964,N_6015);
and U8795 (N_8795,N_6344,N_7019);
xor U8796 (N_8796,N_6883,N_7143);
or U8797 (N_8797,N_7143,N_6380);
nand U8798 (N_8798,N_6795,N_7186);
or U8799 (N_8799,N_6811,N_7280);
nor U8800 (N_8800,N_6830,N_6548);
or U8801 (N_8801,N_6114,N_6115);
xor U8802 (N_8802,N_6500,N_6865);
xnor U8803 (N_8803,N_6507,N_6735);
nand U8804 (N_8804,N_7024,N_7217);
nor U8805 (N_8805,N_6571,N_6490);
and U8806 (N_8806,N_6334,N_6594);
and U8807 (N_8807,N_6586,N_6688);
and U8808 (N_8808,N_6774,N_6479);
xor U8809 (N_8809,N_6956,N_6478);
or U8810 (N_8810,N_7386,N_6117);
nor U8811 (N_8811,N_6381,N_6115);
nand U8812 (N_8812,N_6379,N_6131);
nor U8813 (N_8813,N_6324,N_7014);
xnor U8814 (N_8814,N_6112,N_7011);
nor U8815 (N_8815,N_7161,N_6331);
nand U8816 (N_8816,N_6442,N_7295);
nand U8817 (N_8817,N_6110,N_6538);
nand U8818 (N_8818,N_6042,N_6787);
or U8819 (N_8819,N_7027,N_6689);
or U8820 (N_8820,N_7405,N_7281);
and U8821 (N_8821,N_6172,N_6749);
and U8822 (N_8822,N_6073,N_7237);
or U8823 (N_8823,N_6057,N_6522);
nand U8824 (N_8824,N_7446,N_7113);
or U8825 (N_8825,N_6493,N_6882);
or U8826 (N_8826,N_6081,N_7405);
nand U8827 (N_8827,N_6007,N_7454);
and U8828 (N_8828,N_6632,N_6169);
nand U8829 (N_8829,N_6695,N_6702);
nand U8830 (N_8830,N_6556,N_6663);
and U8831 (N_8831,N_6756,N_6581);
nor U8832 (N_8832,N_7497,N_7152);
nor U8833 (N_8833,N_6426,N_6459);
and U8834 (N_8834,N_6818,N_6758);
nand U8835 (N_8835,N_6573,N_6146);
nand U8836 (N_8836,N_7496,N_7471);
nand U8837 (N_8837,N_6417,N_6394);
xor U8838 (N_8838,N_7240,N_7480);
xnor U8839 (N_8839,N_6926,N_7121);
nand U8840 (N_8840,N_7025,N_6007);
and U8841 (N_8841,N_7339,N_7464);
or U8842 (N_8842,N_6224,N_6577);
and U8843 (N_8843,N_7031,N_6141);
nor U8844 (N_8844,N_6065,N_6932);
nor U8845 (N_8845,N_7308,N_7288);
nor U8846 (N_8846,N_7171,N_7008);
nor U8847 (N_8847,N_6930,N_7367);
and U8848 (N_8848,N_6597,N_6210);
xor U8849 (N_8849,N_6198,N_6704);
nor U8850 (N_8850,N_6023,N_7111);
xor U8851 (N_8851,N_6465,N_6690);
nand U8852 (N_8852,N_6204,N_7197);
nand U8853 (N_8853,N_7370,N_6507);
xnor U8854 (N_8854,N_6389,N_6342);
xor U8855 (N_8855,N_6280,N_6521);
nor U8856 (N_8856,N_6099,N_7070);
or U8857 (N_8857,N_6406,N_6824);
nor U8858 (N_8858,N_6760,N_6319);
nor U8859 (N_8859,N_7415,N_6397);
nor U8860 (N_8860,N_7376,N_7098);
nand U8861 (N_8861,N_6022,N_6786);
nor U8862 (N_8862,N_6033,N_6693);
and U8863 (N_8863,N_7031,N_7262);
and U8864 (N_8864,N_6759,N_6888);
nor U8865 (N_8865,N_7412,N_6380);
xnor U8866 (N_8866,N_6427,N_6846);
or U8867 (N_8867,N_6760,N_6990);
nor U8868 (N_8868,N_7383,N_6271);
nand U8869 (N_8869,N_6234,N_6013);
nand U8870 (N_8870,N_6242,N_7475);
xor U8871 (N_8871,N_6774,N_6504);
nor U8872 (N_8872,N_6556,N_6109);
and U8873 (N_8873,N_6479,N_6655);
nand U8874 (N_8874,N_7004,N_7177);
or U8875 (N_8875,N_6011,N_7211);
and U8876 (N_8876,N_6965,N_6099);
nand U8877 (N_8877,N_6723,N_6289);
and U8878 (N_8878,N_7431,N_6550);
nor U8879 (N_8879,N_7282,N_6760);
nand U8880 (N_8880,N_7255,N_6492);
xor U8881 (N_8881,N_6951,N_6026);
nor U8882 (N_8882,N_7036,N_7457);
xor U8883 (N_8883,N_6359,N_6775);
or U8884 (N_8884,N_7471,N_6546);
nand U8885 (N_8885,N_6054,N_7294);
xnor U8886 (N_8886,N_7449,N_6495);
nor U8887 (N_8887,N_6240,N_6719);
and U8888 (N_8888,N_6910,N_6173);
and U8889 (N_8889,N_7022,N_7366);
nand U8890 (N_8890,N_7445,N_7379);
or U8891 (N_8891,N_7136,N_6011);
or U8892 (N_8892,N_6393,N_6742);
nor U8893 (N_8893,N_7448,N_7068);
or U8894 (N_8894,N_7141,N_6973);
nand U8895 (N_8895,N_6646,N_7001);
nand U8896 (N_8896,N_6634,N_6483);
xnor U8897 (N_8897,N_7387,N_6742);
or U8898 (N_8898,N_6812,N_7191);
nor U8899 (N_8899,N_6110,N_6397);
nor U8900 (N_8900,N_7174,N_6599);
xnor U8901 (N_8901,N_6872,N_7257);
or U8902 (N_8902,N_6812,N_6340);
or U8903 (N_8903,N_6423,N_6105);
nand U8904 (N_8904,N_6777,N_6518);
nand U8905 (N_8905,N_6425,N_6360);
or U8906 (N_8906,N_6356,N_7223);
nand U8907 (N_8907,N_6808,N_7374);
and U8908 (N_8908,N_7127,N_6401);
nand U8909 (N_8909,N_6347,N_6674);
xor U8910 (N_8910,N_6553,N_7495);
and U8911 (N_8911,N_6532,N_7144);
nand U8912 (N_8912,N_6632,N_6012);
and U8913 (N_8913,N_7092,N_6756);
xnor U8914 (N_8914,N_6463,N_7299);
and U8915 (N_8915,N_6130,N_7172);
and U8916 (N_8916,N_6698,N_6923);
or U8917 (N_8917,N_7044,N_6638);
and U8918 (N_8918,N_6570,N_6578);
and U8919 (N_8919,N_6736,N_7277);
xnor U8920 (N_8920,N_7476,N_6409);
xor U8921 (N_8921,N_6450,N_6212);
and U8922 (N_8922,N_7258,N_6506);
nor U8923 (N_8923,N_6485,N_6591);
and U8924 (N_8924,N_7030,N_7009);
nor U8925 (N_8925,N_6769,N_6360);
xor U8926 (N_8926,N_6790,N_6566);
nor U8927 (N_8927,N_7407,N_6366);
xnor U8928 (N_8928,N_6493,N_6153);
and U8929 (N_8929,N_7197,N_6054);
xnor U8930 (N_8930,N_6042,N_6204);
or U8931 (N_8931,N_6833,N_6752);
nor U8932 (N_8932,N_6299,N_7128);
nor U8933 (N_8933,N_7474,N_6137);
nor U8934 (N_8934,N_6715,N_6324);
or U8935 (N_8935,N_6566,N_7371);
nor U8936 (N_8936,N_6052,N_7138);
or U8937 (N_8937,N_6645,N_7132);
or U8938 (N_8938,N_7367,N_7250);
nor U8939 (N_8939,N_7301,N_6537);
and U8940 (N_8940,N_7074,N_6700);
or U8941 (N_8941,N_6601,N_7026);
or U8942 (N_8942,N_6650,N_6468);
nor U8943 (N_8943,N_7198,N_7379);
nor U8944 (N_8944,N_7208,N_7470);
or U8945 (N_8945,N_6736,N_6885);
nor U8946 (N_8946,N_6684,N_7200);
xnor U8947 (N_8947,N_7060,N_6349);
nor U8948 (N_8948,N_7287,N_6239);
nor U8949 (N_8949,N_6070,N_7052);
and U8950 (N_8950,N_7480,N_6952);
nand U8951 (N_8951,N_6833,N_6016);
or U8952 (N_8952,N_6102,N_6805);
and U8953 (N_8953,N_6811,N_6424);
nand U8954 (N_8954,N_7453,N_6740);
and U8955 (N_8955,N_7115,N_6877);
or U8956 (N_8956,N_6737,N_6034);
nand U8957 (N_8957,N_6599,N_6841);
and U8958 (N_8958,N_6883,N_7472);
nor U8959 (N_8959,N_6720,N_7477);
nor U8960 (N_8960,N_7411,N_6614);
or U8961 (N_8961,N_6256,N_6628);
nor U8962 (N_8962,N_7452,N_6073);
or U8963 (N_8963,N_6199,N_7217);
xor U8964 (N_8964,N_7294,N_6291);
nor U8965 (N_8965,N_6457,N_7262);
and U8966 (N_8966,N_6731,N_6519);
nor U8967 (N_8967,N_7242,N_6340);
nand U8968 (N_8968,N_6613,N_6008);
xor U8969 (N_8969,N_6502,N_7317);
nor U8970 (N_8970,N_6206,N_7242);
and U8971 (N_8971,N_6394,N_6605);
nor U8972 (N_8972,N_6687,N_6260);
and U8973 (N_8973,N_7233,N_7010);
xor U8974 (N_8974,N_7110,N_6949);
and U8975 (N_8975,N_6778,N_6153);
or U8976 (N_8976,N_6742,N_6555);
nor U8977 (N_8977,N_6559,N_7208);
and U8978 (N_8978,N_7236,N_6242);
nand U8979 (N_8979,N_6518,N_6249);
nand U8980 (N_8980,N_7341,N_7468);
nor U8981 (N_8981,N_7132,N_6367);
nand U8982 (N_8982,N_6036,N_6416);
xnor U8983 (N_8983,N_6883,N_7103);
or U8984 (N_8984,N_7474,N_6194);
xor U8985 (N_8985,N_6217,N_6872);
or U8986 (N_8986,N_6968,N_6635);
or U8987 (N_8987,N_6348,N_6551);
nor U8988 (N_8988,N_6278,N_7475);
nor U8989 (N_8989,N_6961,N_6640);
xor U8990 (N_8990,N_6627,N_7045);
and U8991 (N_8991,N_6876,N_6030);
nand U8992 (N_8992,N_6753,N_6447);
nand U8993 (N_8993,N_6718,N_6715);
or U8994 (N_8994,N_6867,N_6674);
nor U8995 (N_8995,N_7259,N_7338);
nor U8996 (N_8996,N_7099,N_6119);
xor U8997 (N_8997,N_6861,N_6196);
xor U8998 (N_8998,N_6690,N_6217);
nand U8999 (N_8999,N_6173,N_7489);
nor U9000 (N_9000,N_8177,N_8697);
nand U9001 (N_9001,N_8566,N_8771);
and U9002 (N_9002,N_7928,N_8818);
and U9003 (N_9003,N_7953,N_8823);
xnor U9004 (N_9004,N_7693,N_7547);
nor U9005 (N_9005,N_8123,N_8762);
xnor U9006 (N_9006,N_8600,N_8283);
nand U9007 (N_9007,N_8825,N_8513);
and U9008 (N_9008,N_7633,N_8396);
and U9009 (N_9009,N_7513,N_8217);
nor U9010 (N_9010,N_8258,N_8474);
or U9011 (N_9011,N_7692,N_8964);
or U9012 (N_9012,N_8419,N_8336);
nand U9013 (N_9013,N_7872,N_8004);
nor U9014 (N_9014,N_8181,N_8564);
or U9015 (N_9015,N_8398,N_7667);
or U9016 (N_9016,N_8851,N_8480);
xnor U9017 (N_9017,N_8200,N_8218);
and U9018 (N_9018,N_8432,N_8351);
or U9019 (N_9019,N_8394,N_8953);
nor U9020 (N_9020,N_7676,N_8751);
or U9021 (N_9021,N_8210,N_8760);
or U9022 (N_9022,N_8881,N_8977);
nand U9023 (N_9023,N_8379,N_8111);
and U9024 (N_9024,N_8548,N_8867);
or U9025 (N_9025,N_8046,N_8254);
nor U9026 (N_9026,N_8520,N_8877);
nand U9027 (N_9027,N_7833,N_8387);
nand U9028 (N_9028,N_8051,N_7531);
xnor U9029 (N_9029,N_7587,N_7836);
and U9030 (N_9030,N_8289,N_8882);
and U9031 (N_9031,N_8524,N_8541);
nor U9032 (N_9032,N_7689,N_8163);
and U9033 (N_9033,N_7727,N_8276);
xor U9034 (N_9034,N_7996,N_8244);
nor U9035 (N_9035,N_8984,N_8641);
or U9036 (N_9036,N_7550,N_8993);
nor U9037 (N_9037,N_8628,N_8786);
and U9038 (N_9038,N_8106,N_7604);
nand U9039 (N_9039,N_8365,N_7565);
nor U9040 (N_9040,N_7556,N_7519);
nor U9041 (N_9041,N_8059,N_8206);
nor U9042 (N_9042,N_8457,N_7680);
nor U9043 (N_9043,N_8793,N_8311);
nand U9044 (N_9044,N_8060,N_7706);
xor U9045 (N_9045,N_8640,N_8648);
xor U9046 (N_9046,N_8515,N_8452);
and U9047 (N_9047,N_8035,N_8001);
or U9048 (N_9048,N_8341,N_8089);
nor U9049 (N_9049,N_8159,N_8145);
nand U9050 (N_9050,N_7823,N_7535);
and U9051 (N_9051,N_7522,N_7523);
nor U9052 (N_9052,N_7528,N_8944);
nand U9053 (N_9053,N_7895,N_8691);
nand U9054 (N_9054,N_8601,N_8523);
nand U9055 (N_9055,N_8027,N_8553);
nand U9056 (N_9056,N_7591,N_7827);
or U9057 (N_9057,N_8837,N_8402);
and U9058 (N_9058,N_8608,N_7934);
or U9059 (N_9059,N_8647,N_8579);
xnor U9060 (N_9060,N_7721,N_7758);
nand U9061 (N_9061,N_8033,N_8602);
nand U9062 (N_9062,N_7866,N_8550);
and U9063 (N_9063,N_8589,N_7725);
or U9064 (N_9064,N_8836,N_7746);
nand U9065 (N_9065,N_8805,N_7908);
or U9066 (N_9066,N_7506,N_7651);
nand U9067 (N_9067,N_8479,N_7977);
and U9068 (N_9068,N_7784,N_7955);
nor U9069 (N_9069,N_8108,N_8727);
or U9070 (N_9070,N_8265,N_8312);
or U9071 (N_9071,N_7923,N_8334);
nor U9072 (N_9072,N_8963,N_8031);
or U9073 (N_9073,N_8887,N_8140);
or U9074 (N_9074,N_7790,N_8325);
xor U9075 (N_9075,N_7674,N_8686);
nand U9076 (N_9076,N_8531,N_8885);
and U9077 (N_9077,N_8496,N_8086);
nand U9078 (N_9078,N_8139,N_8293);
nand U9079 (N_9079,N_8758,N_8649);
and U9080 (N_9080,N_8448,N_8291);
nor U9081 (N_9081,N_7780,N_8676);
nor U9082 (N_9082,N_8779,N_8362);
or U9083 (N_9083,N_7538,N_7954);
xor U9084 (N_9084,N_7601,N_8143);
nor U9085 (N_9085,N_8006,N_8785);
and U9086 (N_9086,N_8892,N_8503);
nor U9087 (N_9087,N_8739,N_8831);
and U9088 (N_9088,N_7792,N_8835);
nor U9089 (N_9089,N_7643,N_8395);
xnor U9090 (N_9090,N_8976,N_8471);
xor U9091 (N_9091,N_8516,N_8838);
and U9092 (N_9092,N_8767,N_8952);
xor U9093 (N_9093,N_8209,N_8078);
nor U9094 (N_9094,N_8850,N_8847);
nor U9095 (N_9095,N_7553,N_8631);
nand U9096 (N_9096,N_8295,N_7558);
nor U9097 (N_9097,N_8302,N_7828);
xor U9098 (N_9098,N_8439,N_8546);
nor U9099 (N_9099,N_8603,N_8588);
or U9100 (N_9100,N_8067,N_8063);
nand U9101 (N_9101,N_8083,N_8715);
xor U9102 (N_9102,N_8991,N_7933);
or U9103 (N_9103,N_7940,N_8382);
nand U9104 (N_9104,N_8383,N_8700);
and U9105 (N_9105,N_8079,N_8274);
nand U9106 (N_9106,N_7505,N_7576);
nand U9107 (N_9107,N_8207,N_8346);
and U9108 (N_9108,N_8458,N_8912);
or U9109 (N_9109,N_8569,N_8766);
nand U9110 (N_9110,N_7814,N_8107);
and U9111 (N_9111,N_7831,N_8205);
xnor U9112 (N_9112,N_7798,N_8983);
or U9113 (N_9113,N_8121,N_7672);
or U9114 (N_9114,N_8790,N_7838);
nand U9115 (N_9115,N_7670,N_8570);
and U9116 (N_9116,N_8330,N_7647);
xor U9117 (N_9117,N_8247,N_8152);
nor U9118 (N_9118,N_8454,N_7624);
or U9119 (N_9119,N_8252,N_8655);
xnor U9120 (N_9120,N_7902,N_8975);
nand U9121 (N_9121,N_8896,N_8598);
and U9122 (N_9122,N_8948,N_7991);
xnor U9123 (N_9123,N_8696,N_8685);
or U9124 (N_9124,N_8642,N_7857);
or U9125 (N_9125,N_7888,N_8164);
nor U9126 (N_9126,N_7976,N_7541);
nor U9127 (N_9127,N_8626,N_8441);
nand U9128 (N_9128,N_8465,N_7919);
nand U9129 (N_9129,N_8088,N_7883);
or U9130 (N_9130,N_8702,N_8359);
nor U9131 (N_9131,N_7545,N_7776);
or U9132 (N_9132,N_7697,N_7865);
xor U9133 (N_9133,N_8194,N_8817);
and U9134 (N_9134,N_8022,N_8014);
or U9135 (N_9135,N_8663,N_7551);
nor U9136 (N_9136,N_8591,N_8476);
nand U9137 (N_9137,N_8373,N_7809);
nor U9138 (N_9138,N_7966,N_7724);
or U9139 (N_9139,N_7921,N_8486);
or U9140 (N_9140,N_8040,N_7943);
nand U9141 (N_9141,N_8661,N_8216);
or U9142 (N_9142,N_8594,N_8352);
xor U9143 (N_9143,N_8775,N_7543);
nor U9144 (N_9144,N_7677,N_7532);
nand U9145 (N_9145,N_8129,N_8269);
nor U9146 (N_9146,N_7770,N_7573);
nand U9147 (N_9147,N_7589,N_8543);
and U9148 (N_9148,N_8861,N_8041);
xor U9149 (N_9149,N_8604,N_8888);
nand U9150 (N_9150,N_8481,N_8618);
nor U9151 (N_9151,N_8856,N_8183);
or U9152 (N_9152,N_7615,N_7621);
or U9153 (N_9153,N_8552,N_7652);
nor U9154 (N_9154,N_7690,N_7962);
xor U9155 (N_9155,N_7822,N_8554);
nor U9156 (N_9156,N_7552,N_8556);
and U9157 (N_9157,N_8392,N_7518);
or U9158 (N_9158,N_8609,N_7859);
or U9159 (N_9159,N_8148,N_7851);
and U9160 (N_9160,N_8803,N_8495);
or U9161 (N_9161,N_8461,N_8363);
xor U9162 (N_9162,N_8386,N_7956);
nand U9163 (N_9163,N_8561,N_8037);
xor U9164 (N_9164,N_8555,N_8860);
and U9165 (N_9165,N_7634,N_8468);
and U9166 (N_9166,N_7585,N_8298);
xnor U9167 (N_9167,N_7679,N_7625);
nor U9168 (N_9168,N_7942,N_8931);
xor U9169 (N_9169,N_8630,N_8572);
and U9170 (N_9170,N_7975,N_8511);
nand U9171 (N_9171,N_8199,N_7970);
or U9172 (N_9172,N_8299,N_7862);
and U9173 (N_9173,N_7892,N_8248);
xor U9174 (N_9174,N_8968,N_8733);
nor U9175 (N_9175,N_8822,N_7834);
nand U9176 (N_9176,N_8021,N_8162);
and U9177 (N_9177,N_8095,N_8845);
nor U9178 (N_9178,N_8144,N_7779);
nor U9179 (N_9179,N_8300,N_8911);
or U9180 (N_9180,N_8469,N_7918);
and U9181 (N_9181,N_7596,N_8728);
and U9182 (N_9182,N_8693,N_8287);
nor U9183 (N_9183,N_8273,N_8239);
or U9184 (N_9184,N_8320,N_8377);
and U9185 (N_9185,N_8673,N_8493);
nor U9186 (N_9186,N_7569,N_7570);
xnor U9187 (N_9187,N_8403,N_8622);
nor U9188 (N_9188,N_7613,N_8488);
xor U9189 (N_9189,N_8571,N_8985);
nand U9190 (N_9190,N_7717,N_8434);
nand U9191 (N_9191,N_7752,N_8366);
or U9192 (N_9192,N_7765,N_7713);
xnor U9193 (N_9193,N_7906,N_7959);
or U9194 (N_9194,N_8406,N_8651);
and U9195 (N_9195,N_7747,N_8455);
or U9196 (N_9196,N_8369,N_7716);
nand U9197 (N_9197,N_8783,N_7797);
nand U9198 (N_9198,N_7743,N_8189);
xnor U9199 (N_9199,N_8407,N_8639);
and U9200 (N_9200,N_8580,N_8337);
nand U9201 (N_9201,N_8150,N_7623);
nor U9202 (N_9202,N_8220,N_7517);
or U9203 (N_9203,N_8101,N_7782);
xnor U9204 (N_9204,N_8750,N_8871);
nand U9205 (N_9205,N_8716,N_8195);
or U9206 (N_9206,N_8869,N_8381);
nor U9207 (N_9207,N_8710,N_8744);
nand U9208 (N_9208,N_7773,N_8819);
nand U9209 (N_9209,N_7914,N_7537);
or U9210 (N_9210,N_7696,N_8583);
nand U9211 (N_9211,N_7876,N_7728);
nand U9212 (N_9212,N_7577,N_8732);
nor U9213 (N_9213,N_8076,N_8081);
or U9214 (N_9214,N_7867,N_7911);
nor U9215 (N_9215,N_8978,N_7571);
nor U9216 (N_9216,N_8376,N_8947);
or U9217 (N_9217,N_8301,N_8521);
xnor U9218 (N_9218,N_8400,N_8657);
nand U9219 (N_9219,N_8412,N_8918);
nor U9220 (N_9220,N_7656,N_8806);
nor U9221 (N_9221,N_8592,N_8862);
nand U9222 (N_9222,N_7994,N_8234);
nand U9223 (N_9223,N_8534,N_7771);
or U9224 (N_9224,N_7967,N_8763);
xnor U9225 (N_9225,N_8935,N_7903);
nand U9226 (N_9226,N_8322,N_7945);
and U9227 (N_9227,N_7764,N_8131);
nor U9228 (N_9228,N_8080,N_7864);
or U9229 (N_9229,N_8946,N_8921);
nand U9230 (N_9230,N_8201,N_7600);
and U9231 (N_9231,N_8443,N_8354);
and U9232 (N_9232,N_8280,N_7607);
nand U9233 (N_9233,N_8753,N_8587);
and U9234 (N_9234,N_8232,N_8011);
nand U9235 (N_9235,N_8192,N_7761);
xnor U9236 (N_9236,N_8128,N_7971);
nor U9237 (N_9237,N_7999,N_8787);
or U9238 (N_9238,N_8768,N_7626);
xnor U9239 (N_9239,N_7586,N_8389);
and U9240 (N_9240,N_8824,N_7694);
nor U9241 (N_9241,N_8137,N_8241);
nand U9242 (N_9242,N_7731,N_7509);
or U9243 (N_9243,N_8310,N_8429);
xor U9244 (N_9244,N_7960,N_8242);
nand U9245 (N_9245,N_8627,N_7636);
nor U9246 (N_9246,N_8979,N_8605);
xnor U9247 (N_9247,N_8082,N_8615);
or U9248 (N_9248,N_8582,N_8380);
nand U9249 (N_9249,N_8416,N_8499);
nand U9250 (N_9250,N_7830,N_8694);
or U9251 (N_9251,N_8789,N_8709);
nand U9252 (N_9252,N_7546,N_7846);
nor U9253 (N_9253,N_8134,N_7969);
xor U9254 (N_9254,N_8110,N_8026);
xnor U9255 (N_9255,N_7875,N_8084);
xor U9256 (N_9256,N_7981,N_8249);
or U9257 (N_9257,N_7756,N_8595);
nor U9258 (N_9258,N_8318,N_8430);
xor U9259 (N_9259,N_8634,N_7567);
nand U9260 (N_9260,N_7768,N_8436);
nand U9261 (N_9261,N_7755,N_8726);
or U9262 (N_9262,N_8472,N_7597);
nand U9263 (N_9263,N_8250,N_8510);
and U9264 (N_9264,N_8119,N_7654);
xor U9265 (N_9265,N_8538,N_8054);
nor U9266 (N_9266,N_7946,N_7794);
xnor U9267 (N_9267,N_7803,N_8245);
or U9268 (N_9268,N_8251,N_8857);
xnor U9269 (N_9269,N_8502,N_8662);
nand U9270 (N_9270,N_8208,N_7642);
and U9271 (N_9271,N_8928,N_8230);
nor U9272 (N_9272,N_7832,N_7578);
nand U9273 (N_9273,N_7631,N_7843);
or U9274 (N_9274,N_8506,N_7548);
nor U9275 (N_9275,N_8808,N_7901);
xor U9276 (N_9276,N_8155,N_8166);
or U9277 (N_9277,N_8883,N_7845);
and U9278 (N_9278,N_8064,N_7741);
or U9279 (N_9279,N_8122,N_8719);
nand U9280 (N_9280,N_7791,N_8563);
or U9281 (N_9281,N_7516,N_8738);
and U9282 (N_9282,N_7849,N_8872);
and U9283 (N_9283,N_8275,N_8184);
or U9284 (N_9284,N_8874,N_8530);
and U9285 (N_9285,N_8675,N_8174);
or U9286 (N_9286,N_7612,N_8623);
or U9287 (N_9287,N_8408,N_8186);
nor U9288 (N_9288,N_7575,N_7881);
or U9289 (N_9289,N_7869,N_8423);
and U9290 (N_9290,N_8752,N_7639);
or U9291 (N_9291,N_8316,N_8927);
and U9292 (N_9292,N_8741,N_8816);
nor U9293 (N_9293,N_8171,N_8364);
or U9294 (N_9294,N_8492,N_7512);
and U9295 (N_9295,N_8453,N_8629);
or U9296 (N_9296,N_8990,N_8425);
nand U9297 (N_9297,N_8942,N_8168);
nor U9298 (N_9298,N_7563,N_7748);
or U9299 (N_9299,N_8297,N_8656);
xnor U9300 (N_9300,N_8029,N_8904);
nand U9301 (N_9301,N_8489,N_7941);
or U9302 (N_9302,N_8449,N_8795);
nor U9303 (N_9303,N_7718,N_7742);
nand U9304 (N_9304,N_8136,N_8853);
nand U9305 (N_9305,N_8072,N_8539);
and U9306 (N_9306,N_7950,N_8482);
xnor U9307 (N_9307,N_8706,N_8329);
nand U9308 (N_9308,N_8483,N_8682);
and U9309 (N_9309,N_8126,N_7530);
nor U9310 (N_9310,N_8043,N_8923);
nor U9311 (N_9311,N_8670,N_7990);
xor U9312 (N_9312,N_7719,N_8939);
nor U9313 (N_9313,N_8257,N_8090);
xor U9314 (N_9314,N_7944,N_8282);
nand U9315 (N_9315,N_8562,N_8669);
nor U9316 (N_9316,N_8999,N_7584);
nand U9317 (N_9317,N_7712,N_8243);
nor U9318 (N_9318,N_8420,N_7844);
nor U9319 (N_9319,N_8460,N_7520);
or U9320 (N_9320,N_8982,N_7769);
or U9321 (N_9321,N_7760,N_8328);
nand U9322 (N_9322,N_8485,N_7819);
and U9323 (N_9323,N_8922,N_8533);
nor U9324 (N_9324,N_7661,N_8307);
and U9325 (N_9325,N_8668,N_8438);
nor U9326 (N_9326,N_8950,N_7708);
and U9327 (N_9327,N_7858,N_8813);
and U9328 (N_9328,N_8104,N_8165);
nand U9329 (N_9329,N_7778,N_7599);
and U9330 (N_9330,N_8478,N_7504);
nor U9331 (N_9331,N_8529,N_7985);
xor U9332 (N_9332,N_8451,N_8970);
and U9333 (N_9333,N_8607,N_8013);
and U9334 (N_9334,N_8925,N_7815);
nand U9335 (N_9335,N_8091,N_7659);
or U9336 (N_9336,N_8459,N_8288);
xor U9337 (N_9337,N_8353,N_8005);
nand U9338 (N_9338,N_8278,N_8214);
and U9339 (N_9339,N_7666,N_8565);
or U9340 (N_9340,N_8677,N_8370);
nand U9341 (N_9341,N_7957,N_8262);
xnor U9342 (N_9342,N_7663,N_7890);
or U9343 (N_9343,N_7852,N_7861);
nor U9344 (N_9344,N_7754,N_7655);
nand U9345 (N_9345,N_8358,N_8672);
and U9346 (N_9346,N_8343,N_8305);
nand U9347 (N_9347,N_8893,N_8321);
and U9348 (N_9348,N_7637,N_7525);
nand U9349 (N_9349,N_7650,N_8309);
and U9350 (N_9350,N_8418,N_8294);
xnor U9351 (N_9351,N_8431,N_8135);
nand U9352 (N_9352,N_8030,N_7734);
nand U9353 (N_9353,N_8812,N_7789);
and U9354 (N_9354,N_8507,N_7885);
nand U9355 (N_9355,N_8854,N_8794);
xor U9356 (N_9356,N_8225,N_8116);
or U9357 (N_9357,N_8052,N_8666);
and U9358 (N_9358,N_8138,N_8367);
xor U9359 (N_9359,N_8723,N_7648);
nor U9360 (N_9360,N_8018,N_8017);
nor U9361 (N_9361,N_8391,N_8926);
nand U9362 (N_9362,N_7978,N_7590);
and U9363 (N_9363,N_8019,N_8518);
and U9364 (N_9364,N_7606,N_8315);
xnor U9365 (N_9365,N_8246,N_8167);
nand U9366 (N_9366,N_7687,N_7658);
nand U9367 (N_9367,N_8842,N_8338);
and U9368 (N_9368,N_8442,N_7653);
or U9369 (N_9369,N_8832,N_8105);
nand U9370 (N_9370,N_8290,N_8074);
and U9371 (N_9371,N_8497,N_7753);
nand U9372 (N_9372,N_7929,N_8378);
and U9373 (N_9373,N_7703,N_8114);
xnor U9374 (N_9374,N_8036,N_8858);
or U9375 (N_9375,N_8444,N_7580);
nor U9376 (N_9376,N_8196,N_8992);
and U9377 (N_9377,N_8271,N_8292);
nor U9378 (N_9378,N_7524,N_8303);
nor U9379 (N_9379,N_8075,N_8742);
nor U9380 (N_9380,N_8774,N_8528);
nor U9381 (N_9381,N_8178,N_7704);
and U9382 (N_9382,N_7774,N_8141);
and U9383 (N_9383,N_7788,N_7909);
xor U9384 (N_9384,N_8833,N_7856);
nor U9385 (N_9385,N_8317,N_8193);
nor U9386 (N_9386,N_8734,N_7926);
and U9387 (N_9387,N_7763,N_8901);
nor U9388 (N_9388,N_8834,N_8617);
nor U9389 (N_9389,N_7560,N_8097);
or U9390 (N_9390,N_8221,N_8938);
and U9391 (N_9391,N_8718,N_8955);
and U9392 (N_9392,N_8259,N_7877);
nand U9393 (N_9393,N_8304,N_7947);
nor U9394 (N_9394,N_7611,N_8801);
nor U9395 (N_9395,N_8575,N_8536);
nor U9396 (N_9396,N_8843,N_8578);
xor U9397 (N_9397,N_8849,N_7891);
or U9398 (N_9398,N_8053,N_8047);
and U9399 (N_9399,N_7841,N_8223);
and U9400 (N_9400,N_8224,N_7638);
nor U9401 (N_9401,N_8056,N_7913);
or U9402 (N_9402,N_8695,N_7796);
or U9403 (N_9403,N_7886,N_7810);
or U9404 (N_9404,N_8997,N_8707);
xor U9405 (N_9405,N_8490,N_8113);
and U9406 (N_9406,N_8898,N_8340);
and U9407 (N_9407,N_7900,N_8087);
and U9408 (N_9408,N_7958,N_8308);
or U9409 (N_9409,N_8314,N_7618);
and U9410 (N_9410,N_7562,N_8109);
or U9411 (N_9411,N_7740,N_8125);
xor U9412 (N_9412,N_8974,N_8680);
or U9413 (N_9413,N_8477,N_8807);
and U9414 (N_9414,N_8830,N_7539);
nor U9415 (N_9415,N_7529,N_8498);
xor U9416 (N_9416,N_7668,N_7781);
nor U9417 (N_9417,N_8045,N_8919);
nor U9418 (N_9418,N_8172,N_7566);
nand U9419 (N_9419,N_8235,N_8721);
or U9420 (N_9420,N_7894,N_7644);
nor U9421 (N_9421,N_8450,N_8773);
and U9422 (N_9422,N_8401,N_8897);
nand U9423 (N_9423,N_8375,N_8180);
xor U9424 (N_9424,N_8537,N_7738);
or U9425 (N_9425,N_8714,N_8098);
nand U9426 (N_9426,N_8701,N_8704);
nand U9427 (N_9427,N_8558,N_7993);
or U9428 (N_9428,N_8809,N_8447);
or U9429 (N_9429,N_8428,N_7632);
xor U9430 (N_9430,N_7549,N_7873);
and U9431 (N_9431,N_8446,N_8093);
xor U9432 (N_9432,N_7835,N_8038);
or U9433 (N_9433,N_8745,N_8149);
nor U9434 (N_9434,N_8722,N_8679);
nand U9435 (N_9435,N_7987,N_8612);
xnor U9436 (N_9436,N_7922,N_7848);
and U9437 (N_9437,N_8777,N_8909);
nand U9438 (N_9438,N_8638,N_7744);
and U9439 (N_9439,N_8961,N_8240);
xnor U9440 (N_9440,N_7777,N_8917);
or U9441 (N_9441,N_8724,N_8509);
or U9442 (N_9442,N_7581,N_8466);
nor U9443 (N_9443,N_8757,N_8988);
and U9444 (N_9444,N_7709,N_7605);
nor U9445 (N_9445,N_7868,N_7917);
xor U9446 (N_9446,N_8559,N_7963);
and U9447 (N_9447,N_7602,N_8255);
or U9448 (N_9448,N_7630,N_8573);
nor U9449 (N_9449,N_7593,N_8156);
and U9450 (N_9450,N_7893,N_7715);
xor U9451 (N_9451,N_8981,N_8190);
and U9452 (N_9452,N_8296,N_8659);
nor U9453 (N_9453,N_8410,N_7598);
and U9454 (N_9454,N_7804,N_8348);
nand U9455 (N_9455,N_8426,N_7592);
or U9456 (N_9456,N_8435,N_8527);
or U9457 (N_9457,N_7766,N_8263);
nor U9458 (N_9458,N_8039,N_8417);
nand U9459 (N_9459,N_8705,N_8219);
and U9460 (N_9460,N_7688,N_8414);
xnor U9461 (N_9461,N_7629,N_7821);
xor U9462 (N_9462,N_8099,N_8157);
or U9463 (N_9463,N_8796,N_8028);
xor U9464 (N_9464,N_8233,N_8687);
nand U9465 (N_9465,N_8913,N_8547);
and U9466 (N_9466,N_8781,N_7732);
nor U9467 (N_9467,N_8971,N_8023);
and U9468 (N_9468,N_8103,N_7646);
xnor U9469 (N_9469,N_8962,N_7603);
or U9470 (N_9470,N_8003,N_8132);
xnor U9471 (N_9471,N_8683,N_7785);
nand U9472 (N_9472,N_8737,N_8799);
xor U9473 (N_9473,N_7899,N_7916);
nor U9474 (N_9474,N_7555,N_7588);
nor U9475 (N_9475,N_8972,N_8226);
nor U9476 (N_9476,N_7811,N_8042);
nand U9477 (N_9477,N_8829,N_8908);
nand U9478 (N_9478,N_8256,N_8933);
nor U9479 (N_9479,N_8397,N_8130);
xor U9480 (N_9480,N_8065,N_7887);
nor U9481 (N_9481,N_8285,N_8187);
and U9482 (N_9482,N_8995,N_7511);
xor U9483 (N_9483,N_8413,N_7735);
or U9484 (N_9484,N_8660,N_7952);
nor U9485 (N_9485,N_8540,N_7840);
and U9486 (N_9486,N_8788,N_8611);
or U9487 (N_9487,N_8671,N_8957);
or U9488 (N_9488,N_8462,N_8525);
xor U9489 (N_9489,N_8996,N_8585);
xnor U9490 (N_9490,N_7898,N_8385);
or U9491 (N_9491,N_8526,N_8755);
xnor U9492 (N_9492,N_8712,N_8501);
nand U9493 (N_9493,N_8231,N_8868);
nand U9494 (N_9494,N_7701,N_7561);
and U9495 (N_9495,N_8484,N_8009);
and U9496 (N_9496,N_8765,N_7787);
nand U9497 (N_9497,N_8650,N_7729);
and U9498 (N_9498,N_8117,N_8058);
xnor U9499 (N_9499,N_7767,N_8127);
and U9500 (N_9500,N_7979,N_8024);
nor U9501 (N_9501,N_7514,N_8986);
nand U9502 (N_9502,N_8327,N_7808);
nand U9503 (N_9503,N_8949,N_8720);
nand U9504 (N_9504,N_8266,N_8586);
xnor U9505 (N_9505,N_7502,N_7510);
nand U9506 (N_9506,N_7896,N_8260);
or U9507 (N_9507,N_8681,N_7806);
and U9508 (N_9508,N_8204,N_7574);
xnor U9509 (N_9509,N_8690,N_7932);
nor U9510 (N_9510,N_8185,N_7820);
nand U9511 (N_9511,N_8512,N_7964);
nand U9512 (N_9512,N_8319,N_8487);
and U9513 (N_9513,N_8658,N_8272);
xnor U9514 (N_9514,N_8020,N_7860);
xor U9515 (N_9515,N_7965,N_7936);
xor U9516 (N_9516,N_8597,N_8331);
xor U9517 (N_9517,N_7730,N_8549);
xnor U9518 (N_9518,N_8202,N_8071);
or U9519 (N_9519,N_7825,N_7912);
and U9520 (N_9520,N_7837,N_8153);
or U9521 (N_9521,N_7905,N_8574);
nor U9522 (N_9522,N_8494,N_8906);
and U9523 (N_9523,N_8945,N_8596);
and U9524 (N_9524,N_8717,N_8748);
and U9525 (N_9525,N_7707,N_8930);
and U9526 (N_9526,N_7608,N_8731);
nand U9527 (N_9527,N_8368,N_8173);
and U9528 (N_9528,N_8576,N_8371);
nor U9529 (N_9529,N_7714,N_8878);
xnor U9530 (N_9530,N_8440,N_7995);
or U9531 (N_9531,N_8198,N_8621);
or U9532 (N_9532,N_7772,N_8176);
nor U9533 (N_9533,N_8902,N_8708);
or U9534 (N_9534,N_8624,N_8772);
xnor U9535 (N_9535,N_8112,N_8924);
xor U9536 (N_9536,N_8907,N_8170);
nor U9537 (N_9537,N_8855,N_8593);
nand U9538 (N_9538,N_7839,N_8711);
or U9539 (N_9539,N_8844,N_8409);
and U9540 (N_9540,N_8270,N_8865);
xor U9541 (N_9541,N_8665,N_7984);
nand U9542 (N_9542,N_7847,N_8620);
xnor U9543 (N_9543,N_8848,N_8517);
nor U9544 (N_9544,N_7526,N_8966);
or U9545 (N_9545,N_7948,N_8880);
or U9546 (N_9546,N_7974,N_7521);
nor U9547 (N_9547,N_8929,N_8333);
or U9548 (N_9548,N_8875,N_7980);
nand U9549 (N_9549,N_8960,N_7816);
nand U9550 (N_9550,N_7671,N_8619);
xnor U9551 (N_9551,N_7720,N_7920);
nand U9552 (N_9552,N_8798,N_8994);
nand U9553 (N_9553,N_8780,N_8505);
nand U9554 (N_9554,N_8475,N_8286);
or U9555 (N_9555,N_8264,N_8032);
nor U9556 (N_9556,N_8188,N_7824);
nor U9557 (N_9557,N_8535,N_8749);
or U9558 (N_9558,N_7705,N_8954);
and U9559 (N_9559,N_8070,N_7540);
or U9560 (N_9560,N_8903,N_8890);
or U9561 (N_9561,N_8782,N_7759);
and U9562 (N_9562,N_8584,N_8910);
nand U9563 (N_9563,N_7826,N_8581);
and U9564 (N_9564,N_8491,N_7863);
and U9565 (N_9565,N_8916,N_8002);
and U9566 (N_9566,N_8522,N_7685);
nand U9567 (N_9567,N_8764,N_8743);
nor U9568 (N_9568,N_8519,N_8077);
or U9569 (N_9569,N_8729,N_7675);
or U9570 (N_9570,N_7817,N_7681);
or U9571 (N_9571,N_8182,N_7750);
xor U9572 (N_9572,N_7925,N_8100);
nor U9573 (N_9573,N_8866,N_8102);
or U9574 (N_9574,N_8827,N_8313);
or U9575 (N_9575,N_8007,N_7924);
or U9576 (N_9576,N_8012,N_7927);
nor U9577 (N_9577,N_7842,N_7813);
nand U9578 (N_9578,N_8147,N_8895);
or U9579 (N_9579,N_8160,N_7582);
and U9580 (N_9580,N_8770,N_7628);
or U9581 (N_9581,N_8544,N_7878);
nor U9582 (N_9582,N_7915,N_8055);
or U9583 (N_9583,N_7931,N_7951);
nor U9584 (N_9584,N_8820,N_7880);
nand U9585 (N_9585,N_7879,N_8900);
xnor U9586 (N_9586,N_8551,N_8213);
and U9587 (N_9587,N_8802,N_8094);
and U9588 (N_9588,N_8645,N_8388);
nor U9589 (N_9589,N_8987,N_7657);
and U9590 (N_9590,N_8654,N_7882);
nand U9591 (N_9591,N_8215,N_7800);
or U9592 (N_9592,N_7662,N_8158);
nand U9593 (N_9593,N_7988,N_7594);
and U9594 (N_9594,N_7855,N_8884);
xnor U9595 (N_9595,N_8821,N_8937);
or U9596 (N_9596,N_8010,N_8169);
nor U9597 (N_9597,N_7939,N_8967);
nor U9598 (N_9598,N_7664,N_8306);
xnor U9599 (N_9599,N_8852,N_7961);
and U9600 (N_9600,N_8415,N_7610);
or U9601 (N_9601,N_8048,N_7897);
nand U9602 (N_9602,N_7749,N_8560);
xor U9603 (N_9603,N_8124,N_8889);
nor U9604 (N_9604,N_8936,N_8644);
nor U9605 (N_9605,N_8814,N_7500);
xor U9606 (N_9606,N_8355,N_8016);
and U9607 (N_9607,N_7627,N_8633);
and U9608 (N_9608,N_8236,N_8899);
nand U9609 (N_9609,N_7938,N_8227);
or U9610 (N_9610,N_8356,N_8073);
nand U9611 (N_9611,N_7660,N_8161);
nor U9612 (N_9612,N_8360,N_7542);
or U9613 (N_9613,N_8653,N_7673);
xor U9614 (N_9614,N_8980,N_7572);
and U9615 (N_9615,N_8674,N_8500);
or U9616 (N_9616,N_7684,N_8068);
or U9617 (N_9617,N_7686,N_7733);
and U9618 (N_9618,N_7983,N_8118);
nor U9619 (N_9619,N_8590,N_8464);
or U9620 (N_9620,N_7699,N_8228);
or U9621 (N_9621,N_8151,N_8635);
and U9622 (N_9622,N_8859,N_7982);
or U9623 (N_9623,N_8614,N_7739);
or U9624 (N_9624,N_8735,N_8034);
nor U9625 (N_9625,N_8632,N_8736);
nand U9626 (N_9626,N_8678,N_8754);
nand U9627 (N_9627,N_8342,N_7937);
nand U9628 (N_9628,N_8345,N_8277);
xnor U9629 (N_9629,N_7829,N_7620);
xor U9630 (N_9630,N_7807,N_7870);
xnor U9631 (N_9631,N_8361,N_8756);
and U9632 (N_9632,N_8725,N_7854);
and U9633 (N_9633,N_7850,N_8335);
nand U9634 (N_9634,N_8514,N_8253);
xor U9635 (N_9635,N_8092,N_7564);
nand U9636 (N_9636,N_8421,N_7795);
nand U9637 (N_9637,N_8914,N_7536);
nor U9638 (N_9638,N_8864,N_8399);
nand U9639 (N_9639,N_8828,N_8905);
or U9640 (N_9640,N_8958,N_8085);
or U9641 (N_9641,N_8577,N_7640);
or U9642 (N_9642,N_7695,N_7723);
nand U9643 (N_9643,N_8332,N_8393);
nand U9644 (N_9644,N_8689,N_7989);
xor U9645 (N_9645,N_8713,N_8606);
xor U9646 (N_9646,N_8840,N_7641);
nor U9647 (N_9647,N_7998,N_8846);
nor U9648 (N_9648,N_8470,N_7871);
and U9649 (N_9649,N_7874,N_8636);
or U9650 (N_9650,N_8969,N_8326);
or U9651 (N_9651,N_8212,N_8324);
or U9652 (N_9652,N_7544,N_8769);
nor U9653 (N_9653,N_8810,N_8179);
and U9654 (N_9654,N_8467,N_8504);
xor U9655 (N_9655,N_8115,N_8545);
xnor U9656 (N_9656,N_8175,N_8357);
or U9657 (N_9657,N_8956,N_7557);
or U9658 (N_9658,N_8066,N_8154);
nor U9659 (N_9659,N_7757,N_8684);
or U9660 (N_9660,N_8229,N_8238);
nor U9661 (N_9661,N_7669,N_7997);
nand U9662 (N_9662,N_8870,N_7889);
xnor U9663 (N_9663,N_8008,N_7904);
nor U9664 (N_9664,N_8759,N_8384);
or U9665 (N_9665,N_8989,N_8934);
xor U9666 (N_9666,N_7884,N_7907);
or U9667 (N_9667,N_7745,N_7930);
nor U9668 (N_9668,N_8211,N_8433);
xnor U9669 (N_9669,N_8998,N_8374);
or U9670 (N_9670,N_7614,N_8797);
or U9671 (N_9671,N_8049,N_8941);
and U9672 (N_9672,N_8652,N_8692);
and U9673 (N_9673,N_7935,N_7711);
nor U9674 (N_9674,N_8405,N_8268);
xor U9675 (N_9675,N_8339,N_8776);
and U9676 (N_9676,N_8625,N_8932);
nor U9677 (N_9677,N_8698,N_8940);
xnor U9678 (N_9678,N_7775,N_7554);
and U9679 (N_9679,N_7786,N_8133);
or U9680 (N_9680,N_7683,N_8050);
nand U9681 (N_9681,N_8791,N_7710);
or U9682 (N_9682,N_8761,N_7802);
nand U9683 (N_9683,N_8778,N_7793);
nor U9684 (N_9684,N_8667,N_8699);
and U9685 (N_9685,N_8841,N_7910);
or U9686 (N_9686,N_8800,N_8747);
xnor U9687 (N_9687,N_7619,N_8920);
xor U9688 (N_9688,N_8203,N_8730);
nor U9689 (N_9689,N_7736,N_8025);
xnor U9690 (N_9690,N_8427,N_7722);
nor U9691 (N_9691,N_7665,N_8456);
xnor U9692 (N_9692,N_8891,N_8411);
and U9693 (N_9693,N_7698,N_7783);
xor U9694 (N_9694,N_8894,N_7682);
or U9695 (N_9695,N_7583,N_7818);
or U9696 (N_9696,N_8965,N_8873);
and U9697 (N_9697,N_7949,N_7678);
or U9698 (N_9698,N_8959,N_8267);
nand U9699 (N_9699,N_8532,N_8703);
nor U9700 (N_9700,N_7616,N_8044);
nor U9701 (N_9701,N_7986,N_7515);
and U9702 (N_9702,N_7737,N_8281);
xnor U9703 (N_9703,N_8879,N_8222);
nor U9704 (N_9704,N_8804,N_8863);
and U9705 (N_9705,N_8284,N_7503);
xnor U9706 (N_9706,N_8120,N_8826);
nand U9707 (N_9707,N_8323,N_8951);
and U9708 (N_9708,N_7533,N_8191);
nand U9709 (N_9709,N_8062,N_8613);
or U9710 (N_9710,N_8915,N_7559);
nor U9711 (N_9711,N_7799,N_8557);
or U9712 (N_9712,N_8664,N_7691);
nand U9713 (N_9713,N_7527,N_8061);
nor U9714 (N_9714,N_7853,N_8508);
and U9715 (N_9715,N_8422,N_8599);
nand U9716 (N_9716,N_8740,N_7534);
and U9717 (N_9717,N_8096,N_7617);
nand U9718 (N_9718,N_7751,N_7968);
xor U9719 (N_9719,N_7762,N_8643);
xnor U9720 (N_9720,N_8746,N_8815);
nand U9721 (N_9721,N_8616,N_7501);
or U9722 (N_9722,N_7645,N_8839);
or U9723 (N_9723,N_7568,N_7992);
or U9724 (N_9724,N_8146,N_7649);
nand U9725 (N_9725,N_8943,N_7508);
nor U9726 (N_9726,N_7595,N_8973);
xnor U9727 (N_9727,N_7805,N_7579);
nand U9728 (N_9728,N_8142,N_8567);
or U9729 (N_9729,N_8811,N_8347);
or U9730 (N_9730,N_8237,N_8688);
and U9731 (N_9731,N_7702,N_8069);
nor U9732 (N_9732,N_7972,N_7801);
and U9733 (N_9733,N_7726,N_8792);
and U9734 (N_9734,N_8404,N_8372);
nand U9735 (N_9735,N_8424,N_8344);
or U9736 (N_9736,N_8646,N_8057);
and U9737 (N_9737,N_8610,N_8876);
and U9738 (N_9738,N_8568,N_8350);
or U9739 (N_9739,N_8445,N_8197);
nor U9740 (N_9740,N_7635,N_7609);
xor U9741 (N_9741,N_8015,N_8886);
nand U9742 (N_9742,N_8261,N_8349);
and U9743 (N_9743,N_8784,N_8637);
nor U9744 (N_9744,N_8000,N_8279);
nor U9745 (N_9745,N_8437,N_7812);
xnor U9746 (N_9746,N_8473,N_8463);
or U9747 (N_9747,N_7700,N_7507);
or U9748 (N_9748,N_8542,N_7622);
nor U9749 (N_9749,N_8390,N_7973);
nor U9750 (N_9750,N_7672,N_7711);
xnor U9751 (N_9751,N_8048,N_7792);
nor U9752 (N_9752,N_8187,N_7956);
or U9753 (N_9753,N_8055,N_8228);
nand U9754 (N_9754,N_7849,N_8474);
or U9755 (N_9755,N_7558,N_8005);
or U9756 (N_9756,N_7803,N_8957);
and U9757 (N_9757,N_8534,N_7844);
or U9758 (N_9758,N_7570,N_7645);
or U9759 (N_9759,N_8148,N_7556);
and U9760 (N_9760,N_8426,N_7510);
nand U9761 (N_9761,N_7967,N_8916);
nor U9762 (N_9762,N_7879,N_8172);
and U9763 (N_9763,N_8468,N_7500);
nand U9764 (N_9764,N_8766,N_8326);
and U9765 (N_9765,N_8410,N_8741);
nor U9766 (N_9766,N_8849,N_7960);
nor U9767 (N_9767,N_8997,N_8217);
nand U9768 (N_9768,N_8459,N_8434);
xor U9769 (N_9769,N_8191,N_8119);
nand U9770 (N_9770,N_8886,N_8967);
and U9771 (N_9771,N_8071,N_7711);
nor U9772 (N_9772,N_7605,N_8024);
xor U9773 (N_9773,N_8456,N_8596);
nand U9774 (N_9774,N_7536,N_8806);
nand U9775 (N_9775,N_7916,N_7995);
or U9776 (N_9776,N_8111,N_8166);
nor U9777 (N_9777,N_7995,N_7989);
xor U9778 (N_9778,N_8647,N_7508);
xnor U9779 (N_9779,N_8991,N_8703);
nor U9780 (N_9780,N_8138,N_7560);
or U9781 (N_9781,N_8249,N_8256);
nor U9782 (N_9782,N_8999,N_7888);
or U9783 (N_9783,N_7644,N_8904);
and U9784 (N_9784,N_8124,N_8405);
xor U9785 (N_9785,N_8244,N_7823);
nor U9786 (N_9786,N_8051,N_8489);
and U9787 (N_9787,N_7857,N_8162);
nor U9788 (N_9788,N_8893,N_7976);
xor U9789 (N_9789,N_7617,N_8682);
or U9790 (N_9790,N_7737,N_7792);
nor U9791 (N_9791,N_7676,N_8687);
nor U9792 (N_9792,N_7772,N_8968);
and U9793 (N_9793,N_8411,N_8976);
or U9794 (N_9794,N_7988,N_7918);
or U9795 (N_9795,N_8206,N_8116);
xnor U9796 (N_9796,N_7533,N_8127);
or U9797 (N_9797,N_7523,N_7929);
and U9798 (N_9798,N_7616,N_8319);
or U9799 (N_9799,N_8798,N_7954);
nand U9800 (N_9800,N_8064,N_8364);
and U9801 (N_9801,N_8428,N_7570);
and U9802 (N_9802,N_8060,N_8456);
xnor U9803 (N_9803,N_7896,N_8280);
nor U9804 (N_9804,N_8948,N_8275);
and U9805 (N_9805,N_8642,N_7809);
nand U9806 (N_9806,N_7904,N_8638);
nand U9807 (N_9807,N_8409,N_7508);
or U9808 (N_9808,N_8285,N_8390);
xor U9809 (N_9809,N_7934,N_8619);
or U9810 (N_9810,N_8317,N_7870);
nand U9811 (N_9811,N_8840,N_8131);
nand U9812 (N_9812,N_7734,N_7620);
or U9813 (N_9813,N_8470,N_7947);
nand U9814 (N_9814,N_8823,N_8723);
or U9815 (N_9815,N_7918,N_8182);
xor U9816 (N_9816,N_8833,N_8291);
nor U9817 (N_9817,N_7977,N_7775);
or U9818 (N_9818,N_8025,N_8894);
or U9819 (N_9819,N_8394,N_8500);
or U9820 (N_9820,N_8039,N_8696);
or U9821 (N_9821,N_8748,N_8460);
nand U9822 (N_9822,N_7822,N_8299);
xnor U9823 (N_9823,N_8222,N_7873);
nor U9824 (N_9824,N_8260,N_8710);
nor U9825 (N_9825,N_8154,N_8865);
nand U9826 (N_9826,N_7656,N_7653);
nor U9827 (N_9827,N_8641,N_8202);
and U9828 (N_9828,N_7929,N_7963);
nand U9829 (N_9829,N_7557,N_7680);
and U9830 (N_9830,N_8038,N_8428);
and U9831 (N_9831,N_7554,N_8062);
or U9832 (N_9832,N_8855,N_7617);
and U9833 (N_9833,N_8590,N_8867);
and U9834 (N_9834,N_8517,N_7742);
and U9835 (N_9835,N_7690,N_7623);
xor U9836 (N_9836,N_8246,N_8212);
and U9837 (N_9837,N_8644,N_8816);
nand U9838 (N_9838,N_8137,N_7577);
xor U9839 (N_9839,N_8672,N_7603);
nor U9840 (N_9840,N_8532,N_8187);
or U9841 (N_9841,N_8776,N_8233);
nor U9842 (N_9842,N_7680,N_7856);
nor U9843 (N_9843,N_7968,N_7957);
and U9844 (N_9844,N_8583,N_7751);
nand U9845 (N_9845,N_8756,N_8910);
xnor U9846 (N_9846,N_7548,N_8098);
xor U9847 (N_9847,N_8029,N_8501);
nand U9848 (N_9848,N_8844,N_8179);
and U9849 (N_9849,N_8759,N_8600);
and U9850 (N_9850,N_8466,N_7994);
or U9851 (N_9851,N_7561,N_8200);
xor U9852 (N_9852,N_8283,N_8080);
xor U9853 (N_9853,N_8331,N_7986);
or U9854 (N_9854,N_7679,N_7983);
nor U9855 (N_9855,N_7824,N_7979);
nor U9856 (N_9856,N_8854,N_8124);
nor U9857 (N_9857,N_8443,N_8226);
and U9858 (N_9858,N_7804,N_8845);
xor U9859 (N_9859,N_7892,N_7729);
nand U9860 (N_9860,N_8026,N_7561);
or U9861 (N_9861,N_8543,N_8284);
and U9862 (N_9862,N_8759,N_8772);
nand U9863 (N_9863,N_7808,N_8920);
or U9864 (N_9864,N_8177,N_8252);
nor U9865 (N_9865,N_8554,N_7655);
nor U9866 (N_9866,N_8176,N_8474);
and U9867 (N_9867,N_8723,N_8953);
nor U9868 (N_9868,N_7556,N_8425);
xnor U9869 (N_9869,N_8030,N_8871);
nor U9870 (N_9870,N_7779,N_8859);
nand U9871 (N_9871,N_8018,N_8663);
nor U9872 (N_9872,N_8980,N_7524);
nand U9873 (N_9873,N_7876,N_8044);
xnor U9874 (N_9874,N_8745,N_8338);
xor U9875 (N_9875,N_8009,N_8918);
nand U9876 (N_9876,N_8474,N_8224);
and U9877 (N_9877,N_8209,N_8520);
xnor U9878 (N_9878,N_8636,N_8825);
nor U9879 (N_9879,N_8796,N_7796);
and U9880 (N_9880,N_8918,N_8384);
or U9881 (N_9881,N_8650,N_8334);
nor U9882 (N_9882,N_7640,N_8846);
xor U9883 (N_9883,N_8945,N_8919);
nand U9884 (N_9884,N_8495,N_7709);
nand U9885 (N_9885,N_8134,N_8958);
and U9886 (N_9886,N_8408,N_8321);
or U9887 (N_9887,N_7512,N_8385);
xnor U9888 (N_9888,N_7547,N_7823);
or U9889 (N_9889,N_7935,N_7998);
or U9890 (N_9890,N_7929,N_8694);
and U9891 (N_9891,N_8999,N_8707);
or U9892 (N_9892,N_7746,N_7719);
or U9893 (N_9893,N_8853,N_7535);
xnor U9894 (N_9894,N_7764,N_7866);
or U9895 (N_9895,N_8166,N_7644);
or U9896 (N_9896,N_8558,N_8537);
nor U9897 (N_9897,N_8229,N_7735);
xor U9898 (N_9898,N_8683,N_8902);
or U9899 (N_9899,N_8056,N_8557);
or U9900 (N_9900,N_8046,N_8427);
nor U9901 (N_9901,N_8159,N_8928);
and U9902 (N_9902,N_8580,N_8321);
and U9903 (N_9903,N_7693,N_8618);
xnor U9904 (N_9904,N_7637,N_7973);
nor U9905 (N_9905,N_8756,N_7816);
and U9906 (N_9906,N_8590,N_8451);
or U9907 (N_9907,N_7707,N_7500);
and U9908 (N_9908,N_8756,N_8837);
or U9909 (N_9909,N_7559,N_8750);
xnor U9910 (N_9910,N_7783,N_8553);
nor U9911 (N_9911,N_7586,N_7670);
nand U9912 (N_9912,N_8585,N_7682);
xnor U9913 (N_9913,N_7721,N_8837);
nor U9914 (N_9914,N_8437,N_8691);
nand U9915 (N_9915,N_8457,N_8781);
nand U9916 (N_9916,N_8431,N_8409);
nand U9917 (N_9917,N_8341,N_7969);
nand U9918 (N_9918,N_8165,N_8781);
or U9919 (N_9919,N_8914,N_8719);
xor U9920 (N_9920,N_8697,N_7504);
xnor U9921 (N_9921,N_7540,N_8495);
nor U9922 (N_9922,N_8261,N_8221);
and U9923 (N_9923,N_8750,N_8661);
and U9924 (N_9924,N_8048,N_8617);
or U9925 (N_9925,N_8609,N_8080);
nor U9926 (N_9926,N_8281,N_8463);
xor U9927 (N_9927,N_8486,N_8626);
nand U9928 (N_9928,N_8292,N_8461);
xnor U9929 (N_9929,N_7577,N_7665);
xor U9930 (N_9930,N_7977,N_8582);
or U9931 (N_9931,N_8155,N_8932);
nor U9932 (N_9932,N_8447,N_8108);
nor U9933 (N_9933,N_7857,N_7516);
and U9934 (N_9934,N_7518,N_8559);
and U9935 (N_9935,N_8104,N_7657);
or U9936 (N_9936,N_8296,N_8272);
nor U9937 (N_9937,N_7560,N_8696);
and U9938 (N_9938,N_8980,N_8796);
and U9939 (N_9939,N_7992,N_7953);
nor U9940 (N_9940,N_8743,N_8766);
nand U9941 (N_9941,N_8397,N_8073);
xor U9942 (N_9942,N_8424,N_8512);
nor U9943 (N_9943,N_8744,N_7789);
xnor U9944 (N_9944,N_8438,N_8967);
or U9945 (N_9945,N_7791,N_8369);
or U9946 (N_9946,N_8958,N_8362);
or U9947 (N_9947,N_8882,N_7606);
nand U9948 (N_9948,N_8601,N_8768);
or U9949 (N_9949,N_8759,N_8821);
xnor U9950 (N_9950,N_8771,N_8546);
and U9951 (N_9951,N_8530,N_8479);
nand U9952 (N_9952,N_8932,N_8989);
nand U9953 (N_9953,N_8740,N_7734);
or U9954 (N_9954,N_7826,N_7909);
nor U9955 (N_9955,N_8763,N_7883);
and U9956 (N_9956,N_8776,N_8902);
or U9957 (N_9957,N_7501,N_7762);
or U9958 (N_9958,N_8704,N_7795);
nand U9959 (N_9959,N_8595,N_8686);
xnor U9960 (N_9960,N_8462,N_8842);
xor U9961 (N_9961,N_8542,N_7763);
and U9962 (N_9962,N_7595,N_8365);
nand U9963 (N_9963,N_8009,N_8519);
nor U9964 (N_9964,N_8194,N_8889);
nand U9965 (N_9965,N_8296,N_7520);
or U9966 (N_9966,N_8607,N_7882);
or U9967 (N_9967,N_7590,N_8855);
and U9968 (N_9968,N_8718,N_8020);
nor U9969 (N_9969,N_8258,N_8146);
and U9970 (N_9970,N_8501,N_8424);
nand U9971 (N_9971,N_7749,N_8278);
and U9972 (N_9972,N_8166,N_8696);
and U9973 (N_9973,N_8050,N_8448);
xor U9974 (N_9974,N_8558,N_8081);
and U9975 (N_9975,N_8002,N_7655);
nand U9976 (N_9976,N_8060,N_8515);
xor U9977 (N_9977,N_7968,N_8431);
xnor U9978 (N_9978,N_8543,N_8393);
nand U9979 (N_9979,N_8543,N_8655);
or U9980 (N_9980,N_8098,N_7581);
nor U9981 (N_9981,N_8625,N_7735);
nor U9982 (N_9982,N_8620,N_7635);
nand U9983 (N_9983,N_8137,N_8356);
and U9984 (N_9984,N_7757,N_8991);
nand U9985 (N_9985,N_8626,N_8162);
and U9986 (N_9986,N_7561,N_8127);
nor U9987 (N_9987,N_8245,N_8442);
nor U9988 (N_9988,N_7795,N_8775);
nor U9989 (N_9989,N_8418,N_7827);
xnor U9990 (N_9990,N_7780,N_8917);
xnor U9991 (N_9991,N_7634,N_8735);
and U9992 (N_9992,N_8498,N_8191);
and U9993 (N_9993,N_8740,N_8323);
or U9994 (N_9994,N_8972,N_8524);
nand U9995 (N_9995,N_7630,N_8162);
nand U9996 (N_9996,N_8632,N_7881);
xor U9997 (N_9997,N_8000,N_7647);
or U9998 (N_9998,N_8637,N_8130);
xnor U9999 (N_9999,N_8483,N_8940);
nor U10000 (N_10000,N_8100,N_8959);
nor U10001 (N_10001,N_8482,N_8197);
nor U10002 (N_10002,N_7798,N_8412);
or U10003 (N_10003,N_7768,N_8813);
or U10004 (N_10004,N_8692,N_8783);
nor U10005 (N_10005,N_8185,N_8336);
nor U10006 (N_10006,N_7607,N_8262);
nand U10007 (N_10007,N_7663,N_8683);
nand U10008 (N_10008,N_8059,N_8885);
xnor U10009 (N_10009,N_8563,N_8308);
and U10010 (N_10010,N_8841,N_8719);
xnor U10011 (N_10011,N_8392,N_7675);
nand U10012 (N_10012,N_8872,N_8201);
nand U10013 (N_10013,N_7930,N_8657);
nand U10014 (N_10014,N_7899,N_8413);
or U10015 (N_10015,N_7778,N_7890);
and U10016 (N_10016,N_8483,N_8493);
xor U10017 (N_10017,N_7748,N_8074);
nor U10018 (N_10018,N_7541,N_8040);
nor U10019 (N_10019,N_8507,N_8925);
nor U10020 (N_10020,N_7907,N_8100);
or U10021 (N_10021,N_7524,N_7963);
nor U10022 (N_10022,N_7625,N_8334);
or U10023 (N_10023,N_8339,N_8316);
xor U10024 (N_10024,N_7794,N_8508);
nor U10025 (N_10025,N_8377,N_8090);
and U10026 (N_10026,N_8276,N_8385);
nand U10027 (N_10027,N_8803,N_8206);
nor U10028 (N_10028,N_8017,N_8845);
and U10029 (N_10029,N_8817,N_8781);
or U10030 (N_10030,N_8848,N_7893);
nor U10031 (N_10031,N_8643,N_8674);
or U10032 (N_10032,N_7636,N_8261);
and U10033 (N_10033,N_7531,N_8357);
or U10034 (N_10034,N_8618,N_8332);
xnor U10035 (N_10035,N_8143,N_8862);
and U10036 (N_10036,N_8540,N_8627);
and U10037 (N_10037,N_8355,N_8395);
and U10038 (N_10038,N_8662,N_7690);
or U10039 (N_10039,N_8331,N_8703);
and U10040 (N_10040,N_8873,N_8692);
nor U10041 (N_10041,N_8999,N_8070);
and U10042 (N_10042,N_8327,N_8760);
or U10043 (N_10043,N_7552,N_7513);
nor U10044 (N_10044,N_8237,N_7975);
xnor U10045 (N_10045,N_8919,N_8761);
and U10046 (N_10046,N_7780,N_8221);
and U10047 (N_10047,N_8140,N_7810);
nand U10048 (N_10048,N_8249,N_8281);
nor U10049 (N_10049,N_8400,N_8717);
xnor U10050 (N_10050,N_8115,N_8658);
or U10051 (N_10051,N_8786,N_8606);
and U10052 (N_10052,N_8280,N_8211);
nor U10053 (N_10053,N_8637,N_8062);
or U10054 (N_10054,N_7891,N_8871);
xnor U10055 (N_10055,N_8664,N_8011);
nor U10056 (N_10056,N_7555,N_8982);
and U10057 (N_10057,N_8054,N_8848);
nand U10058 (N_10058,N_7811,N_7936);
or U10059 (N_10059,N_8462,N_8583);
nand U10060 (N_10060,N_8745,N_8612);
nor U10061 (N_10061,N_8444,N_8265);
nor U10062 (N_10062,N_7535,N_7936);
xnor U10063 (N_10063,N_8038,N_7856);
and U10064 (N_10064,N_7951,N_7691);
nand U10065 (N_10065,N_7799,N_8014);
xor U10066 (N_10066,N_7808,N_8588);
xnor U10067 (N_10067,N_8428,N_8563);
or U10068 (N_10068,N_7931,N_8686);
nor U10069 (N_10069,N_8372,N_8340);
or U10070 (N_10070,N_7520,N_8361);
nor U10071 (N_10071,N_8121,N_7805);
nor U10072 (N_10072,N_8182,N_7914);
nand U10073 (N_10073,N_8132,N_8346);
nand U10074 (N_10074,N_8200,N_7914);
nor U10075 (N_10075,N_7773,N_8249);
nor U10076 (N_10076,N_8251,N_8303);
nor U10077 (N_10077,N_8116,N_7788);
nor U10078 (N_10078,N_8621,N_8149);
or U10079 (N_10079,N_8048,N_7793);
nand U10080 (N_10080,N_7769,N_7679);
nor U10081 (N_10081,N_7649,N_8111);
xnor U10082 (N_10082,N_7783,N_8537);
nor U10083 (N_10083,N_7871,N_8717);
or U10084 (N_10084,N_7545,N_7956);
or U10085 (N_10085,N_7527,N_7731);
and U10086 (N_10086,N_7777,N_8819);
nand U10087 (N_10087,N_8727,N_7959);
or U10088 (N_10088,N_8999,N_8995);
nand U10089 (N_10089,N_8968,N_8259);
nor U10090 (N_10090,N_8867,N_8263);
nor U10091 (N_10091,N_8508,N_8235);
nor U10092 (N_10092,N_8099,N_8986);
and U10093 (N_10093,N_8818,N_8209);
xor U10094 (N_10094,N_7972,N_8505);
nand U10095 (N_10095,N_7714,N_7667);
nand U10096 (N_10096,N_8154,N_8509);
nor U10097 (N_10097,N_7549,N_7623);
xnor U10098 (N_10098,N_8909,N_8770);
nand U10099 (N_10099,N_7937,N_7786);
nand U10100 (N_10100,N_8755,N_8622);
nand U10101 (N_10101,N_8085,N_8071);
xor U10102 (N_10102,N_8956,N_8485);
and U10103 (N_10103,N_7973,N_8631);
or U10104 (N_10104,N_7986,N_8818);
or U10105 (N_10105,N_7978,N_8280);
nor U10106 (N_10106,N_8144,N_8483);
nand U10107 (N_10107,N_8096,N_7831);
or U10108 (N_10108,N_7638,N_8234);
xor U10109 (N_10109,N_8234,N_8256);
and U10110 (N_10110,N_8186,N_7791);
or U10111 (N_10111,N_8736,N_8347);
or U10112 (N_10112,N_8417,N_7929);
and U10113 (N_10113,N_8616,N_8214);
nand U10114 (N_10114,N_8412,N_8457);
nor U10115 (N_10115,N_8394,N_8385);
xnor U10116 (N_10116,N_7757,N_8106);
or U10117 (N_10117,N_8091,N_8672);
and U10118 (N_10118,N_7602,N_8776);
or U10119 (N_10119,N_8809,N_7999);
or U10120 (N_10120,N_7991,N_7899);
xor U10121 (N_10121,N_8085,N_8721);
nor U10122 (N_10122,N_8048,N_7854);
nand U10123 (N_10123,N_8595,N_7783);
and U10124 (N_10124,N_8684,N_8357);
and U10125 (N_10125,N_7707,N_8764);
nor U10126 (N_10126,N_8011,N_7704);
or U10127 (N_10127,N_8695,N_8350);
or U10128 (N_10128,N_8083,N_8852);
nand U10129 (N_10129,N_7798,N_7666);
nand U10130 (N_10130,N_8480,N_8995);
nand U10131 (N_10131,N_8023,N_7567);
nand U10132 (N_10132,N_8649,N_8341);
or U10133 (N_10133,N_8683,N_7610);
nor U10134 (N_10134,N_8373,N_8225);
or U10135 (N_10135,N_8176,N_8456);
xnor U10136 (N_10136,N_8820,N_8315);
nor U10137 (N_10137,N_8697,N_8438);
xnor U10138 (N_10138,N_8950,N_8320);
and U10139 (N_10139,N_7927,N_8815);
nand U10140 (N_10140,N_7807,N_7665);
and U10141 (N_10141,N_8088,N_8972);
or U10142 (N_10142,N_7903,N_7971);
xnor U10143 (N_10143,N_8189,N_7774);
and U10144 (N_10144,N_8898,N_7832);
nor U10145 (N_10145,N_7652,N_7653);
nand U10146 (N_10146,N_8319,N_7627);
or U10147 (N_10147,N_8082,N_8878);
nand U10148 (N_10148,N_8418,N_8883);
and U10149 (N_10149,N_8647,N_7989);
xnor U10150 (N_10150,N_7616,N_8958);
and U10151 (N_10151,N_8071,N_7959);
or U10152 (N_10152,N_8037,N_7759);
and U10153 (N_10153,N_8183,N_8440);
nor U10154 (N_10154,N_8140,N_7934);
nor U10155 (N_10155,N_7702,N_8119);
nor U10156 (N_10156,N_8390,N_7953);
nand U10157 (N_10157,N_8682,N_8605);
xor U10158 (N_10158,N_8905,N_8542);
nand U10159 (N_10159,N_8348,N_8039);
nor U10160 (N_10160,N_8843,N_7916);
and U10161 (N_10161,N_7993,N_8169);
or U10162 (N_10162,N_8319,N_8581);
xnor U10163 (N_10163,N_8337,N_8903);
nand U10164 (N_10164,N_7718,N_8414);
or U10165 (N_10165,N_8475,N_7782);
nor U10166 (N_10166,N_8033,N_8081);
and U10167 (N_10167,N_8557,N_8297);
nand U10168 (N_10168,N_8563,N_8273);
xor U10169 (N_10169,N_8429,N_8246);
xnor U10170 (N_10170,N_8566,N_8049);
and U10171 (N_10171,N_7928,N_8429);
or U10172 (N_10172,N_8884,N_8273);
nor U10173 (N_10173,N_8191,N_8894);
nand U10174 (N_10174,N_8146,N_7573);
nor U10175 (N_10175,N_8702,N_8712);
or U10176 (N_10176,N_7710,N_8697);
and U10177 (N_10177,N_8561,N_7952);
nor U10178 (N_10178,N_7595,N_7922);
nand U10179 (N_10179,N_8507,N_8308);
nand U10180 (N_10180,N_7534,N_8612);
xnor U10181 (N_10181,N_8235,N_7631);
xor U10182 (N_10182,N_8216,N_8726);
or U10183 (N_10183,N_8098,N_8793);
xnor U10184 (N_10184,N_8236,N_8016);
and U10185 (N_10185,N_8430,N_8473);
nor U10186 (N_10186,N_8018,N_7979);
or U10187 (N_10187,N_7834,N_8109);
nor U10188 (N_10188,N_8295,N_8626);
or U10189 (N_10189,N_8180,N_7682);
xnor U10190 (N_10190,N_8239,N_7608);
nor U10191 (N_10191,N_8558,N_8997);
nand U10192 (N_10192,N_8769,N_7874);
and U10193 (N_10193,N_8618,N_8520);
and U10194 (N_10194,N_7951,N_7948);
nor U10195 (N_10195,N_8195,N_8573);
xnor U10196 (N_10196,N_8759,N_8588);
nand U10197 (N_10197,N_7750,N_8642);
nand U10198 (N_10198,N_7726,N_8622);
nand U10199 (N_10199,N_8794,N_8467);
nor U10200 (N_10200,N_8829,N_8934);
or U10201 (N_10201,N_7827,N_7753);
or U10202 (N_10202,N_8275,N_8965);
and U10203 (N_10203,N_8376,N_7857);
xnor U10204 (N_10204,N_8759,N_8325);
and U10205 (N_10205,N_7981,N_8599);
xnor U10206 (N_10206,N_8671,N_7646);
nor U10207 (N_10207,N_8762,N_7708);
nor U10208 (N_10208,N_7616,N_7518);
nand U10209 (N_10209,N_8597,N_8514);
nand U10210 (N_10210,N_8191,N_7551);
and U10211 (N_10211,N_8278,N_8978);
or U10212 (N_10212,N_7789,N_8397);
or U10213 (N_10213,N_8942,N_8287);
xor U10214 (N_10214,N_7749,N_8662);
xnor U10215 (N_10215,N_7750,N_8167);
nor U10216 (N_10216,N_7911,N_7909);
nand U10217 (N_10217,N_7837,N_8459);
xnor U10218 (N_10218,N_8175,N_8585);
xnor U10219 (N_10219,N_7988,N_8762);
nand U10220 (N_10220,N_8825,N_8188);
nand U10221 (N_10221,N_8233,N_8226);
and U10222 (N_10222,N_7586,N_8502);
nor U10223 (N_10223,N_8709,N_8578);
and U10224 (N_10224,N_7724,N_7506);
or U10225 (N_10225,N_7978,N_7990);
xor U10226 (N_10226,N_8411,N_8254);
nand U10227 (N_10227,N_8967,N_7564);
nand U10228 (N_10228,N_7558,N_7637);
or U10229 (N_10229,N_7508,N_7608);
nor U10230 (N_10230,N_7691,N_8161);
xnor U10231 (N_10231,N_7617,N_8302);
and U10232 (N_10232,N_8359,N_8567);
xnor U10233 (N_10233,N_7943,N_7906);
nand U10234 (N_10234,N_8603,N_7724);
and U10235 (N_10235,N_8475,N_7501);
or U10236 (N_10236,N_7725,N_8224);
and U10237 (N_10237,N_8994,N_8850);
xnor U10238 (N_10238,N_7663,N_7631);
nor U10239 (N_10239,N_8509,N_8002);
nor U10240 (N_10240,N_8428,N_8333);
xnor U10241 (N_10241,N_8178,N_8236);
nor U10242 (N_10242,N_8865,N_8732);
xnor U10243 (N_10243,N_8982,N_7552);
or U10244 (N_10244,N_8837,N_8773);
nor U10245 (N_10245,N_8191,N_8919);
or U10246 (N_10246,N_8366,N_8926);
and U10247 (N_10247,N_8757,N_8232);
xor U10248 (N_10248,N_7943,N_8552);
or U10249 (N_10249,N_8849,N_7886);
nor U10250 (N_10250,N_7950,N_8396);
or U10251 (N_10251,N_8272,N_8980);
xnor U10252 (N_10252,N_8058,N_8510);
xor U10253 (N_10253,N_8897,N_8334);
xnor U10254 (N_10254,N_8525,N_8754);
and U10255 (N_10255,N_7835,N_8450);
and U10256 (N_10256,N_8292,N_8449);
nor U10257 (N_10257,N_8150,N_7946);
or U10258 (N_10258,N_8575,N_7732);
nand U10259 (N_10259,N_8108,N_8827);
and U10260 (N_10260,N_8222,N_8862);
nand U10261 (N_10261,N_7597,N_8724);
nor U10262 (N_10262,N_7787,N_8537);
or U10263 (N_10263,N_8649,N_8793);
nand U10264 (N_10264,N_8465,N_8017);
and U10265 (N_10265,N_8550,N_8172);
or U10266 (N_10266,N_8800,N_7610);
nand U10267 (N_10267,N_8577,N_8459);
and U10268 (N_10268,N_8834,N_7963);
xor U10269 (N_10269,N_8725,N_7543);
and U10270 (N_10270,N_7787,N_8199);
xnor U10271 (N_10271,N_8966,N_7866);
nand U10272 (N_10272,N_7574,N_8518);
nor U10273 (N_10273,N_8440,N_8637);
xnor U10274 (N_10274,N_7609,N_7629);
and U10275 (N_10275,N_8916,N_8243);
nor U10276 (N_10276,N_8485,N_8940);
nand U10277 (N_10277,N_8179,N_7715);
and U10278 (N_10278,N_8121,N_8587);
and U10279 (N_10279,N_7640,N_7770);
and U10280 (N_10280,N_8659,N_8137);
and U10281 (N_10281,N_8259,N_8910);
nor U10282 (N_10282,N_8822,N_8680);
or U10283 (N_10283,N_8533,N_8044);
nand U10284 (N_10284,N_8261,N_8248);
nand U10285 (N_10285,N_8547,N_8817);
xnor U10286 (N_10286,N_8050,N_8354);
and U10287 (N_10287,N_8621,N_7707);
xor U10288 (N_10288,N_8054,N_8147);
nor U10289 (N_10289,N_8631,N_8743);
nand U10290 (N_10290,N_8757,N_8576);
xnor U10291 (N_10291,N_7869,N_7571);
nand U10292 (N_10292,N_8067,N_8263);
and U10293 (N_10293,N_8428,N_8473);
or U10294 (N_10294,N_8087,N_8949);
nor U10295 (N_10295,N_8137,N_8016);
or U10296 (N_10296,N_7764,N_7661);
nand U10297 (N_10297,N_7791,N_8442);
or U10298 (N_10298,N_8345,N_7962);
xor U10299 (N_10299,N_8181,N_8130);
nor U10300 (N_10300,N_8321,N_7740);
xor U10301 (N_10301,N_8378,N_7930);
nand U10302 (N_10302,N_8849,N_7751);
nand U10303 (N_10303,N_8498,N_7689);
and U10304 (N_10304,N_8888,N_8227);
xnor U10305 (N_10305,N_8301,N_7985);
and U10306 (N_10306,N_7848,N_8195);
and U10307 (N_10307,N_8823,N_8857);
nand U10308 (N_10308,N_8890,N_7599);
and U10309 (N_10309,N_8874,N_7737);
nand U10310 (N_10310,N_8796,N_8194);
nand U10311 (N_10311,N_8121,N_7829);
and U10312 (N_10312,N_8973,N_7830);
or U10313 (N_10313,N_8130,N_8389);
nor U10314 (N_10314,N_7782,N_8233);
or U10315 (N_10315,N_7947,N_8264);
nand U10316 (N_10316,N_8865,N_8158);
nor U10317 (N_10317,N_7687,N_7939);
nor U10318 (N_10318,N_8368,N_8019);
and U10319 (N_10319,N_8694,N_8887);
nor U10320 (N_10320,N_8928,N_8851);
or U10321 (N_10321,N_8169,N_8315);
or U10322 (N_10322,N_7803,N_7859);
or U10323 (N_10323,N_8578,N_8860);
xnor U10324 (N_10324,N_8624,N_7909);
and U10325 (N_10325,N_7571,N_8692);
nand U10326 (N_10326,N_8014,N_7889);
and U10327 (N_10327,N_7976,N_8037);
nor U10328 (N_10328,N_8940,N_8605);
and U10329 (N_10329,N_7830,N_8968);
nor U10330 (N_10330,N_8069,N_8952);
or U10331 (N_10331,N_8998,N_8190);
nor U10332 (N_10332,N_8141,N_8570);
or U10333 (N_10333,N_8633,N_8630);
nand U10334 (N_10334,N_7562,N_8121);
nand U10335 (N_10335,N_8096,N_8225);
nand U10336 (N_10336,N_7940,N_7585);
and U10337 (N_10337,N_7733,N_8243);
nor U10338 (N_10338,N_8121,N_8383);
or U10339 (N_10339,N_8885,N_8837);
xor U10340 (N_10340,N_8104,N_8285);
or U10341 (N_10341,N_8905,N_8869);
or U10342 (N_10342,N_8368,N_8234);
nor U10343 (N_10343,N_8950,N_8173);
nor U10344 (N_10344,N_8222,N_8894);
nor U10345 (N_10345,N_8323,N_8889);
nor U10346 (N_10346,N_7797,N_8629);
nor U10347 (N_10347,N_8047,N_7809);
nor U10348 (N_10348,N_8811,N_7968);
nand U10349 (N_10349,N_7639,N_7835);
or U10350 (N_10350,N_8604,N_7605);
nand U10351 (N_10351,N_8169,N_8652);
nand U10352 (N_10352,N_8433,N_8101);
xor U10353 (N_10353,N_7891,N_7624);
xor U10354 (N_10354,N_8656,N_8105);
xnor U10355 (N_10355,N_8164,N_7914);
nor U10356 (N_10356,N_8679,N_7843);
nand U10357 (N_10357,N_7685,N_8511);
nor U10358 (N_10358,N_8841,N_8840);
nor U10359 (N_10359,N_7880,N_7905);
nor U10360 (N_10360,N_8989,N_8245);
nand U10361 (N_10361,N_7592,N_8625);
and U10362 (N_10362,N_8395,N_8573);
and U10363 (N_10363,N_8525,N_7795);
xnor U10364 (N_10364,N_8689,N_7788);
xnor U10365 (N_10365,N_8660,N_8454);
xor U10366 (N_10366,N_7788,N_7663);
nand U10367 (N_10367,N_8054,N_7734);
and U10368 (N_10368,N_8062,N_8267);
nand U10369 (N_10369,N_8292,N_8602);
nand U10370 (N_10370,N_8078,N_8906);
xor U10371 (N_10371,N_8642,N_7906);
xor U10372 (N_10372,N_8446,N_8777);
or U10373 (N_10373,N_8359,N_8022);
xor U10374 (N_10374,N_8106,N_8990);
nand U10375 (N_10375,N_8467,N_8462);
nor U10376 (N_10376,N_8454,N_7601);
nor U10377 (N_10377,N_8656,N_7989);
nand U10378 (N_10378,N_7643,N_8072);
xnor U10379 (N_10379,N_7746,N_8935);
and U10380 (N_10380,N_7930,N_8694);
xor U10381 (N_10381,N_7744,N_7734);
nor U10382 (N_10382,N_7838,N_8796);
nand U10383 (N_10383,N_7599,N_8503);
or U10384 (N_10384,N_8463,N_7534);
and U10385 (N_10385,N_7517,N_8724);
nand U10386 (N_10386,N_8068,N_8315);
nor U10387 (N_10387,N_7697,N_8694);
and U10388 (N_10388,N_8930,N_8498);
and U10389 (N_10389,N_7695,N_8279);
or U10390 (N_10390,N_8261,N_7849);
nand U10391 (N_10391,N_8488,N_8598);
nor U10392 (N_10392,N_8935,N_8652);
xnor U10393 (N_10393,N_8588,N_8141);
and U10394 (N_10394,N_8922,N_8039);
xnor U10395 (N_10395,N_8480,N_7725);
and U10396 (N_10396,N_8781,N_7638);
or U10397 (N_10397,N_7633,N_8403);
nand U10398 (N_10398,N_8065,N_8508);
or U10399 (N_10399,N_7525,N_7846);
nor U10400 (N_10400,N_8274,N_7548);
or U10401 (N_10401,N_7611,N_8254);
or U10402 (N_10402,N_8349,N_8671);
and U10403 (N_10403,N_8239,N_8618);
xor U10404 (N_10404,N_7826,N_7513);
nor U10405 (N_10405,N_7694,N_8840);
or U10406 (N_10406,N_7990,N_8063);
or U10407 (N_10407,N_8287,N_8118);
nor U10408 (N_10408,N_8801,N_8292);
and U10409 (N_10409,N_8748,N_8645);
nor U10410 (N_10410,N_8060,N_7834);
nor U10411 (N_10411,N_8348,N_8055);
and U10412 (N_10412,N_8262,N_7579);
or U10413 (N_10413,N_8769,N_8951);
xnor U10414 (N_10414,N_7923,N_7647);
xor U10415 (N_10415,N_7894,N_8673);
and U10416 (N_10416,N_7960,N_7614);
xnor U10417 (N_10417,N_7831,N_7776);
and U10418 (N_10418,N_7528,N_8412);
and U10419 (N_10419,N_7893,N_8834);
and U10420 (N_10420,N_8035,N_7822);
nand U10421 (N_10421,N_8858,N_8790);
or U10422 (N_10422,N_7816,N_8449);
or U10423 (N_10423,N_7839,N_7803);
and U10424 (N_10424,N_8335,N_7693);
and U10425 (N_10425,N_8399,N_7665);
and U10426 (N_10426,N_8034,N_8831);
xnor U10427 (N_10427,N_7602,N_8818);
or U10428 (N_10428,N_8046,N_8460);
or U10429 (N_10429,N_7543,N_7989);
nor U10430 (N_10430,N_8299,N_8677);
nand U10431 (N_10431,N_8225,N_8132);
and U10432 (N_10432,N_8263,N_7881);
xor U10433 (N_10433,N_8295,N_8565);
nor U10434 (N_10434,N_8938,N_8240);
and U10435 (N_10435,N_7910,N_7513);
xnor U10436 (N_10436,N_7548,N_8633);
nand U10437 (N_10437,N_8606,N_7731);
or U10438 (N_10438,N_8437,N_8284);
nor U10439 (N_10439,N_8754,N_8524);
nor U10440 (N_10440,N_7972,N_7657);
nand U10441 (N_10441,N_7937,N_7922);
or U10442 (N_10442,N_8348,N_7902);
xnor U10443 (N_10443,N_8182,N_8951);
nor U10444 (N_10444,N_7555,N_8335);
xnor U10445 (N_10445,N_8611,N_8700);
nor U10446 (N_10446,N_8750,N_7627);
and U10447 (N_10447,N_8182,N_8359);
nand U10448 (N_10448,N_7802,N_8886);
and U10449 (N_10449,N_8458,N_8361);
or U10450 (N_10450,N_8271,N_8107);
and U10451 (N_10451,N_8846,N_8396);
nor U10452 (N_10452,N_8997,N_7838);
xnor U10453 (N_10453,N_8497,N_8173);
or U10454 (N_10454,N_8902,N_8113);
or U10455 (N_10455,N_8737,N_8051);
or U10456 (N_10456,N_7630,N_8353);
xnor U10457 (N_10457,N_7563,N_8079);
and U10458 (N_10458,N_7646,N_8486);
nor U10459 (N_10459,N_8069,N_8438);
nor U10460 (N_10460,N_8685,N_8627);
nand U10461 (N_10461,N_8910,N_7749);
xnor U10462 (N_10462,N_8258,N_8534);
and U10463 (N_10463,N_7859,N_8906);
nor U10464 (N_10464,N_7604,N_8034);
or U10465 (N_10465,N_8435,N_8638);
and U10466 (N_10466,N_7627,N_7751);
and U10467 (N_10467,N_8324,N_7625);
nor U10468 (N_10468,N_8686,N_7999);
xor U10469 (N_10469,N_7768,N_8618);
and U10470 (N_10470,N_8108,N_7603);
nand U10471 (N_10471,N_8585,N_8431);
xnor U10472 (N_10472,N_8484,N_8138);
and U10473 (N_10473,N_8929,N_8776);
or U10474 (N_10474,N_7857,N_7518);
xor U10475 (N_10475,N_8952,N_8896);
nand U10476 (N_10476,N_8743,N_7908);
nand U10477 (N_10477,N_8894,N_7994);
and U10478 (N_10478,N_7813,N_8349);
or U10479 (N_10479,N_8190,N_8321);
nor U10480 (N_10480,N_8700,N_8929);
nor U10481 (N_10481,N_7892,N_8779);
xor U10482 (N_10482,N_7752,N_8285);
nand U10483 (N_10483,N_7597,N_8902);
nand U10484 (N_10484,N_8155,N_8243);
nand U10485 (N_10485,N_8856,N_7626);
or U10486 (N_10486,N_7722,N_8718);
and U10487 (N_10487,N_8051,N_7933);
nand U10488 (N_10488,N_7600,N_7912);
xor U10489 (N_10489,N_7923,N_8241);
nand U10490 (N_10490,N_7708,N_7789);
or U10491 (N_10491,N_8168,N_8583);
xor U10492 (N_10492,N_7559,N_8230);
nor U10493 (N_10493,N_8472,N_8485);
nor U10494 (N_10494,N_7522,N_8308);
nor U10495 (N_10495,N_8209,N_8504);
nand U10496 (N_10496,N_7976,N_8327);
and U10497 (N_10497,N_7523,N_8438);
or U10498 (N_10498,N_7556,N_8767);
or U10499 (N_10499,N_8323,N_8555);
xnor U10500 (N_10500,N_9339,N_9265);
and U10501 (N_10501,N_9830,N_10286);
or U10502 (N_10502,N_10159,N_10361);
xor U10503 (N_10503,N_10385,N_9142);
nor U10504 (N_10504,N_10331,N_10447);
nor U10505 (N_10505,N_10197,N_9132);
xor U10506 (N_10506,N_9783,N_10469);
xnor U10507 (N_10507,N_10373,N_10493);
xnor U10508 (N_10508,N_10342,N_10364);
and U10509 (N_10509,N_9283,N_10076);
and U10510 (N_10510,N_9719,N_9342);
or U10511 (N_10511,N_9129,N_9742);
or U10512 (N_10512,N_9947,N_10104);
and U10513 (N_10513,N_9954,N_10395);
xnor U10514 (N_10514,N_9413,N_9236);
nand U10515 (N_10515,N_9647,N_10036);
nand U10516 (N_10516,N_9455,N_9688);
and U10517 (N_10517,N_9471,N_9516);
and U10518 (N_10518,N_9047,N_10021);
or U10519 (N_10519,N_9800,N_10055);
nor U10520 (N_10520,N_10437,N_10013);
nand U10521 (N_10521,N_9023,N_9210);
and U10522 (N_10522,N_10056,N_9391);
nand U10523 (N_10523,N_9670,N_10350);
nor U10524 (N_10524,N_9257,N_9224);
nor U10525 (N_10525,N_10397,N_9259);
nand U10526 (N_10526,N_9502,N_9765);
and U10527 (N_10527,N_9357,N_9535);
nand U10528 (N_10528,N_10495,N_10306);
or U10529 (N_10529,N_9086,N_9794);
nor U10530 (N_10530,N_9465,N_10169);
and U10531 (N_10531,N_10067,N_10434);
nor U10532 (N_10532,N_9809,N_10232);
nor U10533 (N_10533,N_10253,N_10173);
or U10534 (N_10534,N_9043,N_9513);
or U10535 (N_10535,N_9228,N_9204);
xnor U10536 (N_10536,N_10356,N_9088);
nor U10537 (N_10537,N_10498,N_9634);
and U10538 (N_10538,N_9948,N_10047);
or U10539 (N_10539,N_9031,N_10236);
xor U10540 (N_10540,N_9763,N_10140);
and U10541 (N_10541,N_9810,N_9450);
nor U10542 (N_10542,N_9355,N_9917);
nor U10543 (N_10543,N_9706,N_10488);
and U10544 (N_10544,N_10222,N_10320);
nand U10545 (N_10545,N_9686,N_9926);
nor U10546 (N_10546,N_9790,N_9896);
xnor U10547 (N_10547,N_9496,N_9118);
and U10548 (N_10548,N_9856,N_9667);
xor U10549 (N_10549,N_9508,N_9576);
or U10550 (N_10550,N_9051,N_9982);
nor U10551 (N_10551,N_9337,N_9099);
or U10552 (N_10552,N_9890,N_10422);
and U10553 (N_10553,N_9072,N_9317);
nor U10554 (N_10554,N_10280,N_9264);
nand U10555 (N_10555,N_9212,N_9389);
nand U10556 (N_10556,N_9082,N_9555);
or U10557 (N_10557,N_9924,N_10151);
nand U10558 (N_10558,N_9594,N_9770);
or U10559 (N_10559,N_9928,N_9638);
xor U10560 (N_10560,N_10287,N_9219);
and U10561 (N_10561,N_9749,N_10157);
xor U10562 (N_10562,N_9536,N_9093);
nand U10563 (N_10563,N_9444,N_9320);
and U10564 (N_10564,N_9373,N_9834);
or U10565 (N_10565,N_9523,N_10072);
nand U10566 (N_10566,N_10112,N_9044);
nand U10567 (N_10567,N_10419,N_9167);
xnor U10568 (N_10568,N_9549,N_9939);
nor U10569 (N_10569,N_9714,N_10088);
and U10570 (N_10570,N_10011,N_9838);
xnor U10571 (N_10571,N_10249,N_9522);
nor U10572 (N_10572,N_9187,N_9836);
xnor U10573 (N_10573,N_9806,N_9194);
nor U10574 (N_10574,N_9661,N_9307);
or U10575 (N_10575,N_9933,N_9478);
and U10576 (N_10576,N_10353,N_10409);
and U10577 (N_10577,N_9642,N_10439);
xnor U10578 (N_10578,N_9814,N_9037);
xnor U10579 (N_10579,N_9873,N_10051);
or U10580 (N_10580,N_9530,N_10476);
or U10581 (N_10581,N_9493,N_10024);
and U10582 (N_10582,N_9973,N_9696);
or U10583 (N_10583,N_10129,N_10089);
nor U10584 (N_10584,N_9211,N_10374);
nand U10585 (N_10585,N_10283,N_10475);
nand U10586 (N_10586,N_9060,N_9936);
xnor U10587 (N_10587,N_9610,N_10341);
nand U10588 (N_10588,N_9728,N_10180);
or U10589 (N_10589,N_9408,N_9930);
nor U10590 (N_10590,N_9664,N_10177);
nor U10591 (N_10591,N_10053,N_10445);
or U10592 (N_10592,N_9967,N_9232);
nor U10593 (N_10593,N_10212,N_10202);
nand U10594 (N_10594,N_9779,N_9857);
xnor U10595 (N_10595,N_9281,N_9677);
or U10596 (N_10596,N_10473,N_10048);
nor U10597 (N_10597,N_10334,N_10225);
nor U10598 (N_10598,N_10243,N_10292);
nor U10599 (N_10599,N_9533,N_9921);
nor U10600 (N_10600,N_9461,N_9018);
nand U10601 (N_10601,N_9835,N_10126);
nand U10602 (N_10602,N_9633,N_9216);
nand U10603 (N_10603,N_9899,N_9468);
and U10604 (N_10604,N_9971,N_9720);
nand U10605 (N_10605,N_9148,N_9700);
nand U10606 (N_10606,N_9286,N_10430);
nand U10607 (N_10607,N_9263,N_10268);
and U10608 (N_10608,N_9520,N_9575);
xor U10609 (N_10609,N_10207,N_10137);
nand U10610 (N_10610,N_10153,N_10150);
nand U10611 (N_10611,N_9149,N_9112);
or U10612 (N_10612,N_9472,N_9510);
and U10613 (N_10613,N_9115,N_9230);
or U10614 (N_10614,N_10124,N_9207);
and U10615 (N_10615,N_9808,N_10368);
or U10616 (N_10616,N_9394,N_9662);
or U10617 (N_10617,N_9152,N_9143);
and U10618 (N_10618,N_9126,N_10110);
or U10619 (N_10619,N_10022,N_9891);
or U10620 (N_10620,N_9858,N_10133);
nand U10621 (N_10621,N_9932,N_9803);
nand U10622 (N_10622,N_9985,N_9287);
and U10623 (N_10623,N_9256,N_9826);
and U10624 (N_10624,N_9441,N_9267);
or U10625 (N_10625,N_9305,N_10261);
or U10626 (N_10626,N_10101,N_10044);
xnor U10627 (N_10627,N_10269,N_9027);
nand U10628 (N_10628,N_9903,N_9386);
or U10629 (N_10629,N_9711,N_9692);
xnor U10630 (N_10630,N_10081,N_9900);
nand U10631 (N_10631,N_9600,N_9285);
nand U10632 (N_10632,N_9713,N_9909);
and U10633 (N_10633,N_9901,N_10233);
or U10634 (N_10634,N_9447,N_9937);
and U10635 (N_10635,N_10192,N_9704);
and U10636 (N_10636,N_9325,N_9291);
or U10637 (N_10637,N_9761,N_9300);
nor U10638 (N_10638,N_10193,N_10194);
and U10639 (N_10639,N_10317,N_9243);
xor U10640 (N_10640,N_10310,N_9295);
xnor U10641 (N_10641,N_9382,N_9871);
or U10642 (N_10642,N_9592,N_9403);
and U10643 (N_10643,N_9079,N_10058);
nand U10644 (N_10644,N_9990,N_10172);
and U10645 (N_10645,N_10214,N_10463);
nand U10646 (N_10646,N_9608,N_10230);
nor U10647 (N_10647,N_9248,N_9850);
and U10648 (N_10648,N_9613,N_9153);
xor U10649 (N_10649,N_9306,N_9262);
xnor U10650 (N_10650,N_10034,N_9843);
xor U10651 (N_10651,N_10102,N_9246);
xor U10652 (N_10652,N_9254,N_10348);
and U10653 (N_10653,N_9802,N_10064);
nor U10654 (N_10654,N_10464,N_9318);
xor U10655 (N_10655,N_9495,N_9528);
and U10656 (N_10656,N_10059,N_9828);
and U10657 (N_10657,N_9147,N_9116);
nor U10658 (N_10658,N_10494,N_9334);
nor U10659 (N_10659,N_9723,N_10443);
or U10660 (N_10660,N_9620,N_9807);
nor U10661 (N_10661,N_10438,N_10378);
or U10662 (N_10662,N_9229,N_9327);
nor U10663 (N_10663,N_9073,N_9326);
nor U10664 (N_10664,N_9344,N_9128);
xor U10665 (N_10665,N_9547,N_10389);
nor U10666 (N_10666,N_9546,N_9832);
or U10667 (N_10667,N_10267,N_9021);
nand U10668 (N_10668,N_10497,N_9619);
and U10669 (N_10669,N_10198,N_9294);
and U10670 (N_10670,N_9226,N_9369);
nor U10671 (N_10671,N_9273,N_9693);
nor U10672 (N_10672,N_10060,N_9577);
xor U10673 (N_10673,N_9847,N_9867);
nand U10674 (N_10674,N_9599,N_9505);
xnor U10675 (N_10675,N_10403,N_9239);
xor U10676 (N_10676,N_10315,N_9451);
and U10677 (N_10677,N_10357,N_10027);
xnor U10678 (N_10678,N_10239,N_9905);
and U10679 (N_10679,N_10390,N_9422);
xor U10680 (N_10680,N_9480,N_9584);
and U10681 (N_10681,N_9851,N_9712);
nor U10682 (N_10682,N_10467,N_9078);
xor U10683 (N_10683,N_10296,N_10041);
nand U10684 (N_10684,N_9952,N_10431);
or U10685 (N_10685,N_9484,N_9590);
xor U10686 (N_10686,N_9296,N_9103);
nand U10687 (N_10687,N_10483,N_10136);
nand U10688 (N_10688,N_9379,N_9362);
xor U10689 (N_10689,N_9883,N_9722);
and U10690 (N_10690,N_9241,N_10131);
or U10691 (N_10691,N_10371,N_9639);
and U10692 (N_10692,N_10108,N_10100);
xor U10693 (N_10693,N_10185,N_9504);
xor U10694 (N_10694,N_9804,N_9597);
nor U10695 (N_10695,N_9427,N_9151);
xor U10696 (N_10696,N_10250,N_9063);
xor U10697 (N_10697,N_10039,N_9815);
nor U10698 (N_10698,N_9687,N_9902);
or U10699 (N_10699,N_10470,N_10127);
or U10700 (N_10700,N_10226,N_9573);
xnor U10701 (N_10701,N_9423,N_10071);
and U10702 (N_10702,N_9282,N_9587);
xor U10703 (N_10703,N_9284,N_10105);
nand U10704 (N_10704,N_9345,N_9034);
nor U10705 (N_10705,N_10481,N_9785);
nor U10706 (N_10706,N_9012,N_9956);
xor U10707 (N_10707,N_10466,N_9481);
nor U10708 (N_10708,N_9271,N_9884);
xor U10709 (N_10709,N_10444,N_10307);
nand U10710 (N_10710,N_10279,N_9026);
nand U10711 (N_10711,N_9359,N_9668);
xor U10712 (N_10712,N_10082,N_10418);
and U10713 (N_10713,N_9048,N_9155);
nand U10714 (N_10714,N_9940,N_9812);
nand U10715 (N_10715,N_10454,N_9964);
and U10716 (N_10716,N_9065,N_10183);
and U10717 (N_10717,N_10156,N_9154);
nor U10718 (N_10718,N_9558,N_9058);
nand U10719 (N_10719,N_9864,N_9893);
and U10720 (N_10720,N_9245,N_10401);
and U10721 (N_10721,N_9949,N_9439);
xnor U10722 (N_10722,N_9097,N_9341);
or U10723 (N_10723,N_9085,N_9368);
nor U10724 (N_10724,N_9612,N_9643);
nand U10725 (N_10725,N_9489,N_9768);
or U10726 (N_10726,N_10456,N_10363);
and U10727 (N_10727,N_9776,N_10125);
and U10728 (N_10728,N_9360,N_10284);
and U10729 (N_10729,N_9069,N_9446);
nand U10730 (N_10730,N_10008,N_9727);
nor U10731 (N_10731,N_9518,N_9565);
or U10732 (N_10732,N_9583,N_9562);
or U10733 (N_10733,N_9708,N_10042);
or U10734 (N_10734,N_9467,N_9240);
xor U10735 (N_10735,N_9974,N_9372);
or U10736 (N_10736,N_9080,N_9158);
or U10737 (N_10737,N_10103,N_10309);
xor U10738 (N_10738,N_10369,N_9557);
nor U10739 (N_10739,N_9186,N_10235);
or U10740 (N_10740,N_10297,N_9560);
and U10741 (N_10741,N_9421,N_9426);
or U10742 (N_10742,N_10086,N_10229);
or U10743 (N_10743,N_9998,N_9797);
and U10744 (N_10744,N_10449,N_9448);
nand U10745 (N_10745,N_10410,N_10303);
or U10746 (N_10746,N_10486,N_10366);
xor U10747 (N_10747,N_10333,N_10360);
nor U10748 (N_10748,N_9636,N_10455);
nor U10749 (N_10749,N_9313,N_9580);
nor U10750 (N_10750,N_10408,N_9874);
and U10751 (N_10751,N_9989,N_10245);
nand U10752 (N_10752,N_9007,N_9578);
and U10753 (N_10753,N_9199,N_10121);
nor U10754 (N_10754,N_9113,N_9569);
or U10755 (N_10755,N_10291,N_9679);
or U10756 (N_10756,N_9473,N_10045);
or U10757 (N_10757,N_9895,N_9981);
xor U10758 (N_10758,N_9880,N_10035);
or U10759 (N_10759,N_9004,N_10391);
or U10760 (N_10760,N_9579,N_9920);
nand U10761 (N_10761,N_9778,N_9258);
nor U10762 (N_10762,N_10223,N_9059);
or U10763 (N_10763,N_9744,N_10147);
and U10764 (N_10764,N_9321,N_9602);
nand U10765 (N_10765,N_9328,N_10294);
nor U10766 (N_10766,N_10149,N_9529);
nor U10767 (N_10767,N_9332,N_10012);
or U10768 (N_10768,N_10255,N_9675);
and U10769 (N_10769,N_10271,N_9564);
nor U10770 (N_10770,N_9651,N_9351);
and U10771 (N_10771,N_9125,N_9338);
xnor U10772 (N_10772,N_9010,N_10425);
and U10773 (N_10773,N_10171,N_10043);
nand U10774 (N_10774,N_10407,N_9221);
nand U10775 (N_10775,N_9792,N_10116);
xnor U10776 (N_10776,N_9630,N_9469);
nand U10777 (N_10777,N_9526,N_9650);
or U10778 (N_10778,N_10347,N_9092);
nand U10779 (N_10779,N_9617,N_10465);
or U10780 (N_10780,N_9738,N_10380);
xnor U10781 (N_10781,N_10282,N_9213);
or U10782 (N_10782,N_9683,N_10029);
nand U10783 (N_10783,N_9003,N_10352);
or U10784 (N_10784,N_9865,N_9214);
xnor U10785 (N_10785,N_9984,N_10162);
nand U10786 (N_10786,N_9657,N_10336);
and U10787 (N_10787,N_9537,N_9497);
xor U10788 (N_10788,N_10033,N_10312);
or U10789 (N_10789,N_9754,N_9209);
or U10790 (N_10790,N_9791,N_9784);
nor U10791 (N_10791,N_9729,N_9519);
and U10792 (N_10792,N_10077,N_9656);
xnor U10793 (N_10793,N_9242,N_9799);
and U10794 (N_10794,N_9595,N_9877);
xnor U10795 (N_10795,N_9420,N_10379);
or U10796 (N_10796,N_10016,N_10479);
xor U10797 (N_10797,N_9474,N_9388);
or U10798 (N_10798,N_9999,N_9127);
or U10799 (N_10799,N_10050,N_10384);
or U10800 (N_10800,N_10079,N_10091);
and U10801 (N_10801,N_10109,N_9994);
xnor U10802 (N_10802,N_9237,N_10161);
or U10803 (N_10803,N_9629,N_9795);
xnor U10804 (N_10804,N_9868,N_9255);
or U10805 (N_10805,N_10281,N_9816);
and U10806 (N_10806,N_9514,N_9008);
or U10807 (N_10807,N_9190,N_9916);
nor U10808 (N_10808,N_9424,N_9491);
nand U10809 (N_10809,N_9411,N_9684);
and U10810 (N_10810,N_9995,N_9965);
xnor U10811 (N_10811,N_10452,N_9943);
and U10812 (N_10812,N_9122,N_10095);
and U10813 (N_10813,N_10323,N_9637);
nor U10814 (N_10814,N_9030,N_9013);
xnor U10815 (N_10815,N_10240,N_10117);
or U10816 (N_10816,N_9615,N_9658);
xor U10817 (N_10817,N_10383,N_9346);
or U10818 (N_10818,N_10200,N_10424);
nand U10819 (N_10819,N_10251,N_9171);
nor U10820 (N_10820,N_9582,N_9139);
nor U10821 (N_10821,N_10038,N_10491);
xor U10822 (N_10822,N_9494,N_9596);
and U10823 (N_10823,N_10453,N_10062);
or U10824 (N_10824,N_10311,N_10019);
or U10825 (N_10825,N_9840,N_9377);
and U10826 (N_10826,N_9333,N_9436);
nand U10827 (N_10827,N_10496,N_10417);
xnor U10828 (N_10828,N_9781,N_9591);
or U10829 (N_10829,N_9855,N_9534);
nor U10830 (N_10830,N_10004,N_9299);
or U10831 (N_10831,N_9066,N_9951);
or U10832 (N_10832,N_9039,N_9598);
or U10833 (N_10833,N_9046,N_9813);
and U10834 (N_10834,N_9882,N_10241);
xnor U10835 (N_10835,N_9009,N_9314);
or U10836 (N_10836,N_9527,N_9160);
nor U10837 (N_10837,N_9750,N_9911);
xnor U10838 (N_10838,N_9801,N_10365);
nand U10839 (N_10839,N_10477,N_10111);
xnor U10840 (N_10840,N_9348,N_10040);
xor U10841 (N_10841,N_9798,N_9201);
and U10842 (N_10842,N_9133,N_9681);
or U10843 (N_10843,N_10487,N_10474);
nand U10844 (N_10844,N_9550,N_9014);
xnor U10845 (N_10845,N_9041,N_10330);
and U10846 (N_10846,N_9780,N_9177);
nor U10847 (N_10847,N_10097,N_9866);
nor U10848 (N_10848,N_9067,N_9347);
or U10849 (N_10849,N_9992,N_9938);
or U10850 (N_10850,N_9746,N_9825);
nor U10851 (N_10851,N_10204,N_9217);
nand U10852 (N_10852,N_10227,N_9870);
nor U10853 (N_10853,N_9084,N_10399);
and U10854 (N_10854,N_10351,N_10168);
and U10855 (N_10855,N_9957,N_9611);
nand U10856 (N_10856,N_9297,N_9517);
xor U10857 (N_10857,N_9454,N_10224);
or U10858 (N_10858,N_9969,N_9676);
nand U10859 (N_10859,N_9350,N_9701);
xnor U10860 (N_10860,N_9897,N_10370);
xnor U10861 (N_10861,N_9769,N_9384);
nand U10862 (N_10862,N_9352,N_9401);
nor U10863 (N_10863,N_9741,N_10414);
or U10864 (N_10864,N_10023,N_10460);
nand U10865 (N_10865,N_9365,N_9691);
and U10866 (N_10866,N_9498,N_9507);
and U10867 (N_10867,N_9886,N_10244);
nand U10868 (N_10868,N_9782,N_9852);
and U10869 (N_10869,N_10388,N_9089);
nand U10870 (N_10870,N_9609,N_9324);
and U10871 (N_10871,N_9753,N_9961);
xnor U10872 (N_10872,N_9404,N_9280);
or U10873 (N_10873,N_10381,N_9453);
nand U10874 (N_10874,N_10237,N_9845);
or U10875 (N_10875,N_9913,N_9251);
and U10876 (N_10876,N_10482,N_9788);
nand U10877 (N_10877,N_9077,N_10302);
and U10878 (N_10878,N_10134,N_9980);
nand U10879 (N_10879,N_10295,N_9195);
or U10880 (N_10880,N_9572,N_9771);
or U10881 (N_10881,N_9433,N_9872);
nand U10882 (N_10882,N_9690,N_10258);
nor U10883 (N_10883,N_9793,N_9552);
xor U10884 (N_10884,N_9730,N_9945);
or U10885 (N_10885,N_9682,N_9392);
xnor U10886 (N_10886,N_9482,N_10318);
and U10887 (N_10887,N_9457,N_10484);
or U10888 (N_10888,N_10265,N_10423);
xnor U10889 (N_10889,N_9340,N_10325);
nand U10890 (N_10890,N_9588,N_9381);
xnor U10891 (N_10891,N_9185,N_9755);
nor U10892 (N_10892,N_9174,N_9414);
or U10893 (N_10893,N_9509,N_9912);
or U10894 (N_10894,N_9095,N_10078);
nand U10895 (N_10895,N_9958,N_9925);
xnor U10896 (N_10896,N_9006,N_9292);
xor U10897 (N_10897,N_10049,N_9894);
nor U10898 (N_10898,N_9492,N_10376);
nand U10899 (N_10899,N_9290,N_9163);
or U10900 (N_10900,N_9545,N_10090);
xnor U10901 (N_10901,N_9197,N_9252);
xor U10902 (N_10902,N_10184,N_9206);
or U10903 (N_10903,N_10328,N_9997);
nand U10904 (N_10904,N_9398,N_9172);
xor U10905 (N_10905,N_10106,N_9053);
xor U10906 (N_10906,N_9070,N_9499);
nand U10907 (N_10907,N_9036,N_9136);
nand U10908 (N_10908,N_9309,N_9218);
and U10909 (N_10909,N_9929,N_9275);
and U10910 (N_10910,N_9966,N_9068);
nand U10911 (N_10911,N_9694,N_9748);
or U10912 (N_10912,N_10057,N_10206);
xnor U10913 (N_10913,N_10305,N_9378);
nor U10914 (N_10914,N_10068,N_9861);
nor U10915 (N_10915,N_9370,N_9293);
nor U10916 (N_10916,N_9503,N_10063);
xnor U10917 (N_10917,N_9119,N_9543);
nor U10918 (N_10918,N_9652,N_9308);
and U10919 (N_10919,N_10002,N_9574);
xor U10920 (N_10920,N_9076,N_9906);
and U10921 (N_10921,N_9017,N_9644);
nor U10922 (N_10922,N_10329,N_10094);
nor U10923 (N_10923,N_9490,N_9963);
and U10924 (N_10924,N_9544,N_9789);
nand U10925 (N_10925,N_9390,N_9848);
nand U10926 (N_10926,N_9824,N_10429);
xnor U10927 (N_10927,N_9500,N_10179);
nand U10928 (N_10928,N_10070,N_9083);
or U10929 (N_10929,N_9184,N_9200);
or U10930 (N_10930,N_10396,N_10248);
or U10931 (N_10931,N_9972,N_10152);
or U10932 (N_10932,N_9343,N_9434);
xor U10933 (N_10933,N_10472,N_9709);
nand U10934 (N_10934,N_9751,N_9626);
nand U10935 (N_10935,N_9170,N_9567);
and U10936 (N_10936,N_10324,N_9501);
nor U10937 (N_10937,N_9653,N_10181);
or U10938 (N_10938,N_10398,N_9570);
or U10939 (N_10939,N_9485,N_10362);
nor U10940 (N_10940,N_9918,N_10132);
nand U10941 (N_10941,N_9739,N_9539);
nand U10942 (N_10942,N_9055,N_10413);
nand U10943 (N_10943,N_9968,N_9669);
xor U10944 (N_10944,N_10092,N_9205);
and U10945 (N_10945,N_9358,N_9025);
nand U10946 (N_10946,N_9960,N_9462);
xnor U10947 (N_10947,N_9024,N_9946);
and U10948 (N_10948,N_9898,N_9878);
and U10949 (N_10949,N_9437,N_9697);
nand U10950 (N_10950,N_10107,N_9397);
or U10951 (N_10951,N_9459,N_9604);
nand U10952 (N_10952,N_9117,N_10099);
or U10953 (N_10953,N_9585,N_9137);
nand U10954 (N_10954,N_9942,N_9193);
nand U10955 (N_10955,N_9235,N_10231);
xnor U10956 (N_10956,N_9758,N_9707);
or U10957 (N_10957,N_9409,N_9336);
nand U10958 (N_10958,N_9640,N_9892);
nand U10959 (N_10959,N_9762,N_9622);
xor U10960 (N_10960,N_9202,N_9361);
xnor U10961 (N_10961,N_10014,N_10468);
nor U10962 (N_10962,N_10450,N_9772);
or U10963 (N_10963,N_9168,N_10075);
nor U10964 (N_10964,N_9548,N_9056);
xor U10965 (N_10965,N_9144,N_10167);
nand U10966 (N_10966,N_9512,N_10478);
and U10967 (N_10967,N_10451,N_9660);
xor U10968 (N_10968,N_9996,N_10319);
nor U10969 (N_10969,N_9987,N_9915);
nand U10970 (N_10970,N_9179,N_9515);
nand U10971 (N_10971,N_9736,N_10080);
nand U10972 (N_10972,N_9425,N_9104);
nor U10973 (N_10973,N_9935,N_9551);
nand U10974 (N_10974,N_9673,N_9203);
and U10975 (N_10975,N_9475,N_9910);
or U10976 (N_10976,N_9532,N_9822);
xnor U10977 (N_10977,N_10499,N_9849);
xnor U10978 (N_10978,N_9166,N_9674);
nand U10979 (N_10979,N_9111,N_9191);
nor U10980 (N_10980,N_10120,N_9860);
xor U10981 (N_10981,N_9173,N_9466);
xor U10982 (N_10982,N_9098,N_10354);
nor U10983 (N_10983,N_10337,N_9182);
xnor U10984 (N_10984,N_10026,N_9220);
xor U10985 (N_10985,N_10440,N_10344);
nor U10986 (N_10986,N_10358,N_10030);
or U10987 (N_10987,N_10135,N_9247);
and U10988 (N_10988,N_9011,N_9571);
and U10989 (N_10989,N_9443,N_9542);
nor U10990 (N_10990,N_9703,N_9463);
xor U10991 (N_10991,N_10301,N_9888);
xnor U10992 (N_10992,N_9854,N_9716);
and U10993 (N_10993,N_10073,N_9429);
nand U10994 (N_10994,N_9774,N_10145);
nor U10995 (N_10995,N_9641,N_9623);
xnor U10996 (N_10996,N_10142,N_10187);
and U10997 (N_10997,N_10196,N_9022);
nor U10998 (N_10998,N_9135,N_10393);
nand U10999 (N_10999,N_10448,N_9385);
nand U11000 (N_11000,N_9724,N_9811);
xnor U11001 (N_11001,N_10195,N_9511);
nand U11002 (N_11002,N_9624,N_9887);
xor U11003 (N_11003,N_9045,N_9715);
and U11004 (N_11004,N_10158,N_10266);
xor U11005 (N_11005,N_9628,N_10174);
xor U11006 (N_11006,N_9908,N_9107);
nor U11007 (N_11007,N_10205,N_10377);
xnor U11008 (N_11008,N_9371,N_10216);
nor U11009 (N_11009,N_9879,N_10367);
nor U11010 (N_11010,N_9123,N_10001);
and U11011 (N_11011,N_9432,N_9015);
xnor U11012 (N_11012,N_9563,N_9016);
and U11013 (N_11013,N_9827,N_10432);
nand U11014 (N_11014,N_9914,N_9074);
and U11015 (N_11015,N_9227,N_9405);
nand U11016 (N_11016,N_9181,N_9274);
nand U11017 (N_11017,N_9839,N_9438);
xor U11018 (N_11018,N_9354,N_9101);
nand U11019 (N_11019,N_9665,N_9818);
nor U11020 (N_11020,N_10199,N_9464);
nand U11021 (N_11021,N_9417,N_9428);
nor U11022 (N_11022,N_9955,N_9020);
nor U11023 (N_11023,N_9141,N_9764);
and U11024 (N_11024,N_10405,N_10154);
xnor U11025 (N_11025,N_9521,N_9796);
xnor U11026 (N_11026,N_9331,N_10359);
and U11027 (N_11027,N_10052,N_9767);
xor U11028 (N_11028,N_9625,N_9725);
nor U11029 (N_11029,N_10128,N_10256);
and U11030 (N_11030,N_9418,N_10304);
and U11031 (N_11031,N_9396,N_10093);
xnor U11032 (N_11032,N_9435,N_9487);
or U11033 (N_11033,N_10340,N_9071);
nor U11034 (N_11034,N_9260,N_9178);
xnor U11035 (N_11035,N_9869,N_9506);
nor U11036 (N_11036,N_9541,N_10221);
xor U11037 (N_11037,N_9261,N_10201);
xnor U11038 (N_11038,N_10262,N_9150);
or U11039 (N_11039,N_10163,N_9192);
nand U11040 (N_11040,N_9033,N_9310);
and U11041 (N_11041,N_9698,N_10113);
xor U11042 (N_11042,N_9540,N_9164);
xor U11043 (N_11043,N_9322,N_9556);
and U11044 (N_11044,N_9366,N_10436);
nor U11045 (N_11045,N_10300,N_9648);
nor U11046 (N_11046,N_9479,N_9950);
xor U11047 (N_11047,N_10404,N_9988);
or U11048 (N_11048,N_9747,N_10186);
and U11049 (N_11049,N_9430,N_10246);
and U11050 (N_11050,N_10308,N_10355);
or U11051 (N_11051,N_9635,N_10375);
or U11052 (N_11052,N_10416,N_10122);
nor U11053 (N_11053,N_10228,N_9740);
nor U11054 (N_11054,N_9934,N_9941);
nand U11055 (N_11055,N_9986,N_9919);
xor U11056 (N_11056,N_9001,N_9175);
nor U11057 (N_11057,N_9817,N_9614);
or U11058 (N_11058,N_9993,N_9607);
or U11059 (N_11059,N_9064,N_9586);
xnor U11060 (N_11060,N_10166,N_10066);
nor U11061 (N_11061,N_9904,N_9554);
or U11062 (N_11062,N_10332,N_10459);
nor U11063 (N_11063,N_10433,N_9442);
or U11064 (N_11064,N_9659,N_9831);
nor U11065 (N_11065,N_9419,N_10278);
nand U11066 (N_11066,N_10260,N_9655);
and U11067 (N_11067,N_10406,N_9645);
and U11068 (N_11068,N_10096,N_9075);
or U11069 (N_11069,N_10234,N_9250);
nor U11070 (N_11070,N_10217,N_9568);
and U11071 (N_11071,N_9488,N_9244);
and U11072 (N_11072,N_9249,N_10435);
and U11073 (N_11073,N_9605,N_10165);
nor U11074 (N_11074,N_9829,N_9819);
xor U11075 (N_11075,N_9367,N_10471);
or U11076 (N_11076,N_9091,N_9962);
xnor U11077 (N_11077,N_10031,N_9215);
or U11078 (N_11078,N_9276,N_9140);
xnor U11079 (N_11079,N_9124,N_9049);
xor U11080 (N_11080,N_10338,N_10046);
nor U11081 (N_11081,N_10005,N_10028);
or U11082 (N_11082,N_9975,N_9298);
nor U11083 (N_11083,N_9159,N_10208);
or U11084 (N_11084,N_9416,N_9054);
and U11085 (N_11085,N_10346,N_10146);
xor U11086 (N_11086,N_10400,N_9663);
or U11087 (N_11087,N_10492,N_10321);
nand U11088 (N_11088,N_9524,N_10191);
nor U11089 (N_11089,N_10277,N_10190);
or U11090 (N_11090,N_9272,N_9102);
and U11091 (N_11091,N_9105,N_10037);
and U11092 (N_11092,N_9198,N_9477);
and U11093 (N_11093,N_10421,N_10242);
nor U11094 (N_11094,N_10148,N_10020);
or U11095 (N_11095,N_9689,N_9616);
xor U11096 (N_11096,N_10220,N_9889);
and U11097 (N_11097,N_9038,N_9120);
nor U11098 (N_11098,N_9162,N_9702);
nand U11099 (N_11099,N_10327,N_10442);
nand U11100 (N_11100,N_9138,N_9695);
or U11101 (N_11101,N_10461,N_9876);
xnor U11102 (N_11102,N_10018,N_10273);
xnor U11103 (N_11103,N_10219,N_9743);
and U11104 (N_11104,N_9759,N_9062);
nand U11105 (N_11105,N_9970,N_10010);
nor U11106 (N_11106,N_9374,N_9363);
nor U11107 (N_11107,N_10210,N_9319);
and U11108 (N_11108,N_9090,N_10316);
nor U11109 (N_11109,N_9983,N_9050);
nand U11110 (N_11110,N_9991,N_10458);
and U11111 (N_11111,N_9268,N_9821);
and U11112 (N_11112,N_9029,N_9631);
and U11113 (N_11113,N_10335,N_9589);
nor U11114 (N_11114,N_10025,N_9094);
or U11115 (N_11115,N_9846,N_9161);
and U11116 (N_11116,N_10144,N_9412);
xor U11117 (N_11117,N_9735,N_9165);
xnor U11118 (N_11118,N_9380,N_9183);
or U11119 (N_11119,N_10061,N_9823);
xor U11120 (N_11120,N_10189,N_10130);
nor U11121 (N_11121,N_9927,N_10009);
nand U11122 (N_11122,N_10382,N_9766);
xnor U11123 (N_11123,N_10209,N_10485);
nand U11124 (N_11124,N_9431,N_9531);
and U11125 (N_11125,N_9238,N_10290);
or U11126 (N_11126,N_9944,N_9820);
nor U11127 (N_11127,N_9134,N_10293);
nand U11128 (N_11128,N_9837,N_10087);
nand U11129 (N_11129,N_10114,N_9907);
nand U11130 (N_11130,N_9859,N_9277);
or U11131 (N_11131,N_9678,N_9052);
xor U11132 (N_11132,N_9559,N_9335);
xnor U11133 (N_11133,N_9005,N_9393);
nand U11134 (N_11134,N_9188,N_9976);
xnor U11135 (N_11135,N_10138,N_10402);
nor U11136 (N_11136,N_9862,N_9316);
or U11137 (N_11137,N_9476,N_9196);
or U11138 (N_11138,N_9844,N_10238);
or U11139 (N_11139,N_9145,N_9169);
nor U11140 (N_11140,N_9035,N_9156);
nand U11141 (N_11141,N_9233,N_9106);
or U11142 (N_11142,N_9731,N_10415);
or U11143 (N_11143,N_9114,N_9376);
and U11144 (N_11144,N_10420,N_9110);
xnor U11145 (N_11145,N_10314,N_10392);
or U11146 (N_11146,N_9649,N_9737);
or U11147 (N_11147,N_10480,N_10457);
and U11148 (N_11148,N_9978,N_9402);
and U11149 (N_11149,N_9279,N_9019);
xor U11150 (N_11150,N_9486,N_9225);
xnor U11151 (N_11151,N_9288,N_9756);
nand U11152 (N_11152,N_10462,N_9449);
or U11153 (N_11153,N_10247,N_9407);
or U11154 (N_11154,N_10322,N_10175);
nor U11155 (N_11155,N_9356,N_10000);
nand U11156 (N_11156,N_9666,N_10254);
nand U11157 (N_11157,N_9959,N_10188);
nor U11158 (N_11158,N_9881,N_9603);
or U11159 (N_11159,N_9842,N_10182);
xnor U11160 (N_11160,N_10313,N_9400);
nand U11161 (N_11161,N_9253,N_9760);
xnor U11162 (N_11162,N_10387,N_10115);
nand U11163 (N_11163,N_9452,N_9705);
and U11164 (N_11164,N_9087,N_10326);
or U11165 (N_11165,N_9953,N_10032);
xor U11166 (N_11166,N_9726,N_10289);
xor U11167 (N_11167,N_9266,N_9538);
or U11168 (N_11168,N_10288,N_9329);
and U11169 (N_11169,N_9234,N_9734);
and U11170 (N_11170,N_9718,N_9180);
nand U11171 (N_11171,N_9627,N_9301);
and U11172 (N_11172,N_9732,N_10003);
nand U11173 (N_11173,N_10394,N_9108);
nor U11174 (N_11174,N_9146,N_9786);
xor U11175 (N_11175,N_10065,N_10215);
nor U11176 (N_11176,N_9289,N_9470);
nor U11177 (N_11177,N_10446,N_9863);
and U11178 (N_11178,N_9757,N_9922);
and U11179 (N_11179,N_9395,N_9923);
or U11180 (N_11180,N_10349,N_9566);
nand U11181 (N_11181,N_9121,N_9853);
nor U11182 (N_11182,N_10264,N_10274);
and U11183 (N_11183,N_10141,N_10178);
nand U11184 (N_11184,N_10119,N_10083);
and U11185 (N_11185,N_10218,N_9733);
nor U11186 (N_11186,N_10155,N_10343);
nor U11187 (N_11187,N_10007,N_10170);
nor U11188 (N_11188,N_10203,N_9773);
and U11189 (N_11189,N_10263,N_9375);
or U11190 (N_11190,N_9311,N_9081);
or U11191 (N_11191,N_10285,N_9330);
xor U11192 (N_11192,N_9302,N_9787);
nor U11193 (N_11193,N_9745,N_10372);
xnor U11194 (N_11194,N_9977,N_9752);
and U11195 (N_11195,N_10143,N_9040);
or U11196 (N_11196,N_9654,N_10441);
xor U11197 (N_11197,N_9445,N_9775);
xnor U11198 (N_11198,N_9777,N_9672);
nand U11199 (N_11199,N_9130,N_10074);
xor U11200 (N_11200,N_10069,N_9315);
or U11201 (N_11201,N_10345,N_10386);
xor U11202 (N_11202,N_9671,N_9456);
nor U11203 (N_11203,N_10259,N_9028);
nor U11204 (N_11204,N_9157,N_9269);
nor U11205 (N_11205,N_9000,N_9223);
or U11206 (N_11206,N_9581,N_9410);
nor U11207 (N_11207,N_10085,N_10299);
or U11208 (N_11208,N_10257,N_10252);
or U11209 (N_11209,N_10426,N_9349);
or U11210 (N_11210,N_9440,N_9231);
and U11211 (N_11211,N_10015,N_9270);
nor U11212 (N_11212,N_9979,N_10017);
nor U11213 (N_11213,N_10276,N_9383);
xnor U11214 (N_11214,N_9312,N_10211);
or U11215 (N_11215,N_10411,N_10176);
and U11216 (N_11216,N_10118,N_10164);
nor U11217 (N_11217,N_9553,N_9032);
nor U11218 (N_11218,N_9189,N_9606);
and U11219 (N_11219,N_10084,N_10428);
nor U11220 (N_11220,N_10490,N_9303);
and U11221 (N_11221,N_10427,N_10054);
nand U11222 (N_11222,N_9176,N_9222);
or U11223 (N_11223,N_10160,N_10006);
nand U11224 (N_11224,N_9323,N_10272);
nand U11225 (N_11225,N_10339,N_10098);
and U11226 (N_11226,N_9061,N_9885);
xor U11227 (N_11227,N_9680,N_9399);
and U11228 (N_11228,N_9621,N_9304);
xnor U11229 (N_11229,N_9710,N_9685);
nand U11230 (N_11230,N_9525,N_9593);
nor U11231 (N_11231,N_10270,N_9717);
or U11232 (N_11232,N_9131,N_9100);
xnor U11233 (N_11233,N_9931,N_9387);
nor U11234 (N_11234,N_9646,N_9875);
or U11235 (N_11235,N_9805,N_10123);
nand U11236 (N_11236,N_10489,N_9415);
xnor U11237 (N_11237,N_10275,N_9601);
nand U11238 (N_11238,N_10298,N_9632);
and U11239 (N_11239,N_10139,N_9460);
and U11240 (N_11240,N_10412,N_9109);
nand U11241 (N_11241,N_9278,N_9406);
nor U11242 (N_11242,N_9699,N_9618);
nor U11243 (N_11243,N_9458,N_9721);
or U11244 (N_11244,N_9057,N_9353);
or U11245 (N_11245,N_9096,N_9841);
nand U11246 (N_11246,N_9208,N_9002);
nand U11247 (N_11247,N_9833,N_9042);
nand U11248 (N_11248,N_9561,N_10213);
nor U11249 (N_11249,N_9483,N_9364);
nand U11250 (N_11250,N_9949,N_10126);
nor U11251 (N_11251,N_9419,N_9837);
nor U11252 (N_11252,N_10227,N_9303);
or U11253 (N_11253,N_9342,N_9950);
nor U11254 (N_11254,N_10061,N_10244);
xor U11255 (N_11255,N_9613,N_9591);
and U11256 (N_11256,N_9965,N_9941);
or U11257 (N_11257,N_9963,N_9045);
nor U11258 (N_11258,N_9746,N_9834);
nor U11259 (N_11259,N_9147,N_10497);
or U11260 (N_11260,N_9709,N_9067);
nor U11261 (N_11261,N_9540,N_9672);
nor U11262 (N_11262,N_9906,N_9516);
xor U11263 (N_11263,N_10226,N_9354);
nand U11264 (N_11264,N_10275,N_10150);
or U11265 (N_11265,N_10221,N_9529);
nand U11266 (N_11266,N_9161,N_10161);
xor U11267 (N_11267,N_9204,N_9425);
and U11268 (N_11268,N_9094,N_10395);
and U11269 (N_11269,N_9039,N_10428);
xnor U11270 (N_11270,N_9043,N_10078);
and U11271 (N_11271,N_10301,N_9471);
or U11272 (N_11272,N_9013,N_10040);
nor U11273 (N_11273,N_9669,N_9135);
and U11274 (N_11274,N_9908,N_9964);
nor U11275 (N_11275,N_10475,N_9649);
nand U11276 (N_11276,N_9968,N_9711);
nand U11277 (N_11277,N_9463,N_9179);
nand U11278 (N_11278,N_9067,N_10383);
nand U11279 (N_11279,N_9137,N_10416);
nor U11280 (N_11280,N_9069,N_10159);
nor U11281 (N_11281,N_9993,N_10126);
nand U11282 (N_11282,N_9597,N_10064);
nor U11283 (N_11283,N_9817,N_9043);
nor U11284 (N_11284,N_10165,N_9925);
or U11285 (N_11285,N_10172,N_10076);
xnor U11286 (N_11286,N_9242,N_9142);
xnor U11287 (N_11287,N_10230,N_10172);
and U11288 (N_11288,N_10102,N_10153);
or U11289 (N_11289,N_9594,N_9504);
or U11290 (N_11290,N_9004,N_9730);
or U11291 (N_11291,N_9093,N_9046);
xor U11292 (N_11292,N_9955,N_9645);
xor U11293 (N_11293,N_10303,N_10228);
nor U11294 (N_11294,N_10333,N_9411);
and U11295 (N_11295,N_9269,N_10145);
xnor U11296 (N_11296,N_9082,N_9649);
xnor U11297 (N_11297,N_9063,N_9320);
or U11298 (N_11298,N_10482,N_9433);
nor U11299 (N_11299,N_9082,N_9732);
and U11300 (N_11300,N_9734,N_9845);
or U11301 (N_11301,N_10393,N_9535);
or U11302 (N_11302,N_10292,N_9203);
nor U11303 (N_11303,N_9748,N_10377);
nand U11304 (N_11304,N_10186,N_9069);
nor U11305 (N_11305,N_9432,N_9508);
nor U11306 (N_11306,N_10303,N_10386);
nor U11307 (N_11307,N_9424,N_9191);
or U11308 (N_11308,N_9385,N_10391);
or U11309 (N_11309,N_9293,N_10040);
nor U11310 (N_11310,N_9519,N_9832);
nand U11311 (N_11311,N_9733,N_10219);
nand U11312 (N_11312,N_9245,N_9578);
or U11313 (N_11313,N_9619,N_10285);
xor U11314 (N_11314,N_10434,N_9737);
and U11315 (N_11315,N_9614,N_10399);
xnor U11316 (N_11316,N_9208,N_9957);
or U11317 (N_11317,N_9253,N_9176);
or U11318 (N_11318,N_10288,N_9806);
xnor U11319 (N_11319,N_9859,N_9106);
xnor U11320 (N_11320,N_10230,N_9359);
nand U11321 (N_11321,N_9089,N_9106);
and U11322 (N_11322,N_9389,N_9093);
and U11323 (N_11323,N_9443,N_10343);
xnor U11324 (N_11324,N_9838,N_10223);
xnor U11325 (N_11325,N_9487,N_9273);
and U11326 (N_11326,N_9149,N_9953);
or U11327 (N_11327,N_9833,N_10422);
nand U11328 (N_11328,N_10009,N_9410);
and U11329 (N_11329,N_10307,N_9762);
nor U11330 (N_11330,N_10384,N_9995);
nor U11331 (N_11331,N_9288,N_9968);
or U11332 (N_11332,N_10309,N_9754);
xor U11333 (N_11333,N_10138,N_10245);
nand U11334 (N_11334,N_9440,N_9371);
and U11335 (N_11335,N_10139,N_9731);
and U11336 (N_11336,N_10199,N_9869);
or U11337 (N_11337,N_9249,N_10296);
or U11338 (N_11338,N_9038,N_10364);
xor U11339 (N_11339,N_9223,N_10046);
and U11340 (N_11340,N_9446,N_10157);
and U11341 (N_11341,N_10294,N_10150);
nand U11342 (N_11342,N_9378,N_10214);
or U11343 (N_11343,N_10473,N_10097);
nand U11344 (N_11344,N_10323,N_9663);
xor U11345 (N_11345,N_9942,N_10480);
xnor U11346 (N_11346,N_9676,N_9576);
and U11347 (N_11347,N_9475,N_9887);
and U11348 (N_11348,N_10465,N_10250);
and U11349 (N_11349,N_9935,N_10430);
and U11350 (N_11350,N_9669,N_10134);
xor U11351 (N_11351,N_9850,N_10435);
xor U11352 (N_11352,N_9768,N_9910);
xnor U11353 (N_11353,N_9731,N_9571);
and U11354 (N_11354,N_10049,N_9007);
nor U11355 (N_11355,N_9869,N_10212);
and U11356 (N_11356,N_9703,N_10393);
and U11357 (N_11357,N_9892,N_9981);
xor U11358 (N_11358,N_10399,N_10380);
nor U11359 (N_11359,N_10213,N_9710);
and U11360 (N_11360,N_10231,N_9002);
or U11361 (N_11361,N_9936,N_9795);
or U11362 (N_11362,N_10191,N_9872);
or U11363 (N_11363,N_10173,N_9530);
and U11364 (N_11364,N_9463,N_10027);
xor U11365 (N_11365,N_10148,N_10263);
or U11366 (N_11366,N_9697,N_10068);
nand U11367 (N_11367,N_9453,N_9919);
xor U11368 (N_11368,N_10145,N_10409);
or U11369 (N_11369,N_9771,N_9343);
and U11370 (N_11370,N_9074,N_9270);
xor U11371 (N_11371,N_10178,N_9153);
nor U11372 (N_11372,N_9673,N_9125);
and U11373 (N_11373,N_9060,N_9771);
xnor U11374 (N_11374,N_9963,N_10179);
and U11375 (N_11375,N_10098,N_9961);
or U11376 (N_11376,N_10122,N_10222);
or U11377 (N_11377,N_9390,N_9962);
nor U11378 (N_11378,N_10290,N_9062);
nand U11379 (N_11379,N_9215,N_9135);
nand U11380 (N_11380,N_9036,N_9571);
and U11381 (N_11381,N_9649,N_9967);
xor U11382 (N_11382,N_10054,N_10458);
and U11383 (N_11383,N_10368,N_9167);
nand U11384 (N_11384,N_10031,N_9986);
or U11385 (N_11385,N_9224,N_9913);
nor U11386 (N_11386,N_10228,N_10199);
nor U11387 (N_11387,N_10399,N_10029);
and U11388 (N_11388,N_9684,N_9176);
nand U11389 (N_11389,N_9204,N_9402);
and U11390 (N_11390,N_9194,N_9463);
xor U11391 (N_11391,N_9956,N_9809);
and U11392 (N_11392,N_9480,N_9692);
or U11393 (N_11393,N_9713,N_10374);
nand U11394 (N_11394,N_9228,N_9563);
nand U11395 (N_11395,N_9598,N_9764);
nand U11396 (N_11396,N_9796,N_9506);
or U11397 (N_11397,N_9376,N_9426);
nor U11398 (N_11398,N_9758,N_9024);
and U11399 (N_11399,N_10227,N_9119);
or U11400 (N_11400,N_9334,N_9318);
and U11401 (N_11401,N_9427,N_9206);
xnor U11402 (N_11402,N_9504,N_10380);
nand U11403 (N_11403,N_9455,N_9028);
and U11404 (N_11404,N_10166,N_10007);
nor U11405 (N_11405,N_10366,N_10348);
nor U11406 (N_11406,N_9910,N_9120);
xnor U11407 (N_11407,N_9663,N_9355);
or U11408 (N_11408,N_9435,N_9285);
xnor U11409 (N_11409,N_9331,N_9342);
and U11410 (N_11410,N_9965,N_9457);
and U11411 (N_11411,N_9410,N_9712);
nor U11412 (N_11412,N_9748,N_9052);
or U11413 (N_11413,N_9314,N_10439);
or U11414 (N_11414,N_9717,N_9494);
and U11415 (N_11415,N_10000,N_9593);
and U11416 (N_11416,N_10341,N_10093);
nand U11417 (N_11417,N_10466,N_10355);
xor U11418 (N_11418,N_9676,N_10234);
nor U11419 (N_11419,N_9972,N_10319);
nand U11420 (N_11420,N_9669,N_9108);
nor U11421 (N_11421,N_10241,N_10465);
and U11422 (N_11422,N_9775,N_9154);
xor U11423 (N_11423,N_9006,N_9934);
nand U11424 (N_11424,N_9621,N_9168);
xor U11425 (N_11425,N_9703,N_10108);
and U11426 (N_11426,N_9724,N_9773);
xnor U11427 (N_11427,N_9644,N_9766);
xnor U11428 (N_11428,N_10177,N_10304);
and U11429 (N_11429,N_9112,N_9658);
xnor U11430 (N_11430,N_9005,N_9691);
and U11431 (N_11431,N_9408,N_10000);
and U11432 (N_11432,N_9665,N_9730);
xor U11433 (N_11433,N_10376,N_10378);
nand U11434 (N_11434,N_9172,N_9813);
and U11435 (N_11435,N_9816,N_9499);
and U11436 (N_11436,N_9354,N_9253);
nor U11437 (N_11437,N_10064,N_10047);
and U11438 (N_11438,N_9871,N_10138);
xor U11439 (N_11439,N_9622,N_9468);
or U11440 (N_11440,N_9050,N_9151);
nand U11441 (N_11441,N_9936,N_10257);
and U11442 (N_11442,N_10127,N_9900);
nand U11443 (N_11443,N_9668,N_9120);
nand U11444 (N_11444,N_9613,N_9780);
nor U11445 (N_11445,N_9513,N_9090);
xor U11446 (N_11446,N_10171,N_9323);
xnor U11447 (N_11447,N_9452,N_9589);
and U11448 (N_11448,N_9104,N_9209);
or U11449 (N_11449,N_10349,N_9886);
or U11450 (N_11450,N_9825,N_9208);
and U11451 (N_11451,N_9573,N_9337);
or U11452 (N_11452,N_9811,N_10037);
and U11453 (N_11453,N_9383,N_9651);
or U11454 (N_11454,N_9767,N_9074);
or U11455 (N_11455,N_10188,N_9516);
nand U11456 (N_11456,N_10276,N_9822);
xor U11457 (N_11457,N_9484,N_10321);
or U11458 (N_11458,N_10362,N_9162);
or U11459 (N_11459,N_10250,N_9428);
or U11460 (N_11460,N_9806,N_10134);
and U11461 (N_11461,N_9270,N_9957);
nor U11462 (N_11462,N_10428,N_10496);
nand U11463 (N_11463,N_9139,N_10174);
or U11464 (N_11464,N_9237,N_9273);
nand U11465 (N_11465,N_9150,N_9944);
xor U11466 (N_11466,N_9549,N_9103);
nand U11467 (N_11467,N_10113,N_10196);
xor U11468 (N_11468,N_9091,N_10329);
nand U11469 (N_11469,N_9932,N_10373);
xor U11470 (N_11470,N_10081,N_9535);
and U11471 (N_11471,N_9751,N_10329);
nor U11472 (N_11472,N_10480,N_9145);
and U11473 (N_11473,N_9030,N_10497);
nor U11474 (N_11474,N_9736,N_9610);
xor U11475 (N_11475,N_9404,N_10258);
nor U11476 (N_11476,N_9948,N_10088);
and U11477 (N_11477,N_9590,N_9485);
xnor U11478 (N_11478,N_10456,N_9569);
or U11479 (N_11479,N_9335,N_9936);
and U11480 (N_11480,N_9602,N_9798);
and U11481 (N_11481,N_9423,N_10481);
or U11482 (N_11482,N_10294,N_9610);
or U11483 (N_11483,N_10036,N_9758);
and U11484 (N_11484,N_9653,N_10464);
xor U11485 (N_11485,N_9613,N_9218);
or U11486 (N_11486,N_9776,N_9220);
or U11487 (N_11487,N_9680,N_9797);
or U11488 (N_11488,N_9535,N_9258);
xor U11489 (N_11489,N_9425,N_9619);
and U11490 (N_11490,N_9262,N_10056);
xor U11491 (N_11491,N_9135,N_10361);
xnor U11492 (N_11492,N_9468,N_10454);
nand U11493 (N_11493,N_9399,N_9987);
xor U11494 (N_11494,N_10042,N_9330);
and U11495 (N_11495,N_9806,N_10127);
nand U11496 (N_11496,N_10141,N_9577);
and U11497 (N_11497,N_9872,N_9072);
nor U11498 (N_11498,N_10031,N_9785);
nand U11499 (N_11499,N_9820,N_9180);
nand U11500 (N_11500,N_9749,N_9079);
xor U11501 (N_11501,N_10060,N_9932);
xnor U11502 (N_11502,N_9736,N_9357);
xnor U11503 (N_11503,N_9649,N_10011);
nor U11504 (N_11504,N_10169,N_9010);
or U11505 (N_11505,N_10050,N_10059);
xor U11506 (N_11506,N_9602,N_9179);
nand U11507 (N_11507,N_10102,N_9529);
and U11508 (N_11508,N_10391,N_9920);
nand U11509 (N_11509,N_9321,N_9404);
nor U11510 (N_11510,N_9113,N_9402);
nor U11511 (N_11511,N_9641,N_10278);
nor U11512 (N_11512,N_9299,N_9145);
nor U11513 (N_11513,N_9093,N_10062);
and U11514 (N_11514,N_9337,N_9233);
and U11515 (N_11515,N_9689,N_9760);
xor U11516 (N_11516,N_10190,N_10081);
nor U11517 (N_11517,N_9270,N_9950);
nor U11518 (N_11518,N_9896,N_9101);
xor U11519 (N_11519,N_9371,N_9267);
and U11520 (N_11520,N_9573,N_9053);
nor U11521 (N_11521,N_9603,N_9545);
nand U11522 (N_11522,N_9812,N_9031);
and U11523 (N_11523,N_9708,N_9841);
xnor U11524 (N_11524,N_9749,N_9816);
and U11525 (N_11525,N_9009,N_9471);
nor U11526 (N_11526,N_9976,N_9728);
xor U11527 (N_11527,N_10106,N_10094);
nor U11528 (N_11528,N_9131,N_9458);
nand U11529 (N_11529,N_10333,N_10252);
xnor U11530 (N_11530,N_10292,N_9110);
xor U11531 (N_11531,N_9068,N_9385);
xnor U11532 (N_11532,N_9690,N_9249);
and U11533 (N_11533,N_9203,N_9308);
nor U11534 (N_11534,N_10296,N_9927);
and U11535 (N_11535,N_9040,N_9803);
nor U11536 (N_11536,N_9938,N_9463);
or U11537 (N_11537,N_10174,N_9076);
xnor U11538 (N_11538,N_9442,N_9755);
or U11539 (N_11539,N_10411,N_9450);
or U11540 (N_11540,N_9894,N_9174);
nand U11541 (N_11541,N_10286,N_10205);
xor U11542 (N_11542,N_9401,N_9794);
xnor U11543 (N_11543,N_9183,N_9895);
and U11544 (N_11544,N_9809,N_10005);
and U11545 (N_11545,N_9932,N_9889);
nand U11546 (N_11546,N_9256,N_9349);
nand U11547 (N_11547,N_9343,N_9448);
nand U11548 (N_11548,N_10278,N_9020);
and U11549 (N_11549,N_10061,N_9592);
and U11550 (N_11550,N_10337,N_10185);
nor U11551 (N_11551,N_10485,N_10422);
xnor U11552 (N_11552,N_9152,N_10402);
nor U11553 (N_11553,N_9004,N_10096);
nor U11554 (N_11554,N_10116,N_9847);
xnor U11555 (N_11555,N_9600,N_10486);
nor U11556 (N_11556,N_9002,N_9954);
or U11557 (N_11557,N_10353,N_9542);
xor U11558 (N_11558,N_9620,N_10114);
xor U11559 (N_11559,N_10212,N_9610);
xor U11560 (N_11560,N_9267,N_9477);
nor U11561 (N_11561,N_9900,N_9005);
xor U11562 (N_11562,N_9278,N_9721);
or U11563 (N_11563,N_10301,N_9058);
nor U11564 (N_11564,N_9127,N_9600);
nor U11565 (N_11565,N_9315,N_9660);
nand U11566 (N_11566,N_9046,N_9237);
xor U11567 (N_11567,N_10084,N_9213);
nand U11568 (N_11568,N_9447,N_9921);
or U11569 (N_11569,N_9446,N_9846);
nor U11570 (N_11570,N_9090,N_10257);
and U11571 (N_11571,N_9097,N_9231);
nand U11572 (N_11572,N_10267,N_9926);
or U11573 (N_11573,N_9502,N_9495);
or U11574 (N_11574,N_9718,N_10453);
nor U11575 (N_11575,N_9632,N_9964);
nor U11576 (N_11576,N_9851,N_9022);
and U11577 (N_11577,N_10230,N_9256);
nor U11578 (N_11578,N_9647,N_10293);
xor U11579 (N_11579,N_9967,N_9425);
or U11580 (N_11580,N_9129,N_9181);
and U11581 (N_11581,N_9199,N_10227);
or U11582 (N_11582,N_9564,N_10346);
xnor U11583 (N_11583,N_10493,N_9951);
and U11584 (N_11584,N_10262,N_10407);
nor U11585 (N_11585,N_10148,N_9793);
or U11586 (N_11586,N_10121,N_10433);
nor U11587 (N_11587,N_9571,N_9787);
nand U11588 (N_11588,N_10044,N_9794);
or U11589 (N_11589,N_10211,N_10024);
xor U11590 (N_11590,N_10106,N_10476);
or U11591 (N_11591,N_10399,N_9524);
xor U11592 (N_11592,N_9387,N_9919);
nor U11593 (N_11593,N_9348,N_10311);
or U11594 (N_11594,N_9182,N_9131);
nand U11595 (N_11595,N_9803,N_9712);
xnor U11596 (N_11596,N_9313,N_9443);
nand U11597 (N_11597,N_10331,N_9372);
and U11598 (N_11598,N_9698,N_9891);
and U11599 (N_11599,N_9817,N_9654);
xor U11600 (N_11600,N_9420,N_9566);
and U11601 (N_11601,N_10196,N_9117);
xnor U11602 (N_11602,N_10388,N_9345);
xor U11603 (N_11603,N_9013,N_10414);
and U11604 (N_11604,N_9791,N_10322);
nor U11605 (N_11605,N_9942,N_9561);
xnor U11606 (N_11606,N_9105,N_10406);
nand U11607 (N_11607,N_9755,N_10015);
nor U11608 (N_11608,N_10463,N_9140);
nand U11609 (N_11609,N_10229,N_9304);
and U11610 (N_11610,N_10354,N_10214);
nor U11611 (N_11611,N_9414,N_9057);
xor U11612 (N_11612,N_10043,N_9402);
nand U11613 (N_11613,N_10232,N_10185);
or U11614 (N_11614,N_9093,N_9528);
xor U11615 (N_11615,N_10233,N_10016);
and U11616 (N_11616,N_9650,N_9845);
nor U11617 (N_11617,N_9581,N_10047);
nand U11618 (N_11618,N_10480,N_9276);
or U11619 (N_11619,N_9355,N_9265);
and U11620 (N_11620,N_10140,N_10093);
or U11621 (N_11621,N_10424,N_10404);
and U11622 (N_11622,N_10314,N_10253);
or U11623 (N_11623,N_10443,N_9137);
or U11624 (N_11624,N_9087,N_9802);
and U11625 (N_11625,N_9805,N_9701);
xnor U11626 (N_11626,N_9758,N_9573);
nand U11627 (N_11627,N_10094,N_9475);
nor U11628 (N_11628,N_9013,N_10465);
nor U11629 (N_11629,N_9968,N_10401);
nand U11630 (N_11630,N_9374,N_10304);
nor U11631 (N_11631,N_9408,N_9489);
nand U11632 (N_11632,N_9807,N_9640);
or U11633 (N_11633,N_10246,N_9886);
nand U11634 (N_11634,N_9129,N_9099);
xor U11635 (N_11635,N_9334,N_10259);
or U11636 (N_11636,N_9186,N_9519);
nand U11637 (N_11637,N_9658,N_10450);
and U11638 (N_11638,N_9053,N_10043);
xnor U11639 (N_11639,N_10128,N_9204);
nand U11640 (N_11640,N_9740,N_9317);
xor U11641 (N_11641,N_9230,N_9633);
and U11642 (N_11642,N_10262,N_10280);
xnor U11643 (N_11643,N_9974,N_10338);
nor U11644 (N_11644,N_9369,N_9992);
nand U11645 (N_11645,N_9069,N_10161);
nor U11646 (N_11646,N_9795,N_10187);
or U11647 (N_11647,N_9943,N_10060);
xnor U11648 (N_11648,N_10144,N_10075);
or U11649 (N_11649,N_9773,N_9147);
or U11650 (N_11650,N_9372,N_10173);
or U11651 (N_11651,N_9037,N_9008);
nor U11652 (N_11652,N_10184,N_9581);
nand U11653 (N_11653,N_9897,N_10332);
nand U11654 (N_11654,N_9971,N_9531);
nor U11655 (N_11655,N_9040,N_10094);
nand U11656 (N_11656,N_9385,N_9979);
nand U11657 (N_11657,N_9350,N_9417);
xnor U11658 (N_11658,N_10401,N_10273);
nand U11659 (N_11659,N_10083,N_10379);
nor U11660 (N_11660,N_9883,N_10197);
nand U11661 (N_11661,N_9809,N_10085);
xor U11662 (N_11662,N_10439,N_10005);
and U11663 (N_11663,N_10384,N_9596);
nand U11664 (N_11664,N_9781,N_10005);
and U11665 (N_11665,N_10203,N_10233);
and U11666 (N_11666,N_9635,N_9278);
or U11667 (N_11667,N_9802,N_9261);
nor U11668 (N_11668,N_9797,N_9704);
nand U11669 (N_11669,N_10207,N_10463);
or U11670 (N_11670,N_10065,N_9684);
xor U11671 (N_11671,N_9769,N_9391);
or U11672 (N_11672,N_10348,N_10374);
nand U11673 (N_11673,N_10118,N_9755);
or U11674 (N_11674,N_10491,N_9010);
or U11675 (N_11675,N_9323,N_9454);
nor U11676 (N_11676,N_9079,N_10207);
nand U11677 (N_11677,N_9951,N_9680);
nand U11678 (N_11678,N_9013,N_9545);
or U11679 (N_11679,N_10495,N_9479);
nor U11680 (N_11680,N_9570,N_10067);
nand U11681 (N_11681,N_10352,N_9205);
or U11682 (N_11682,N_10090,N_9756);
and U11683 (N_11683,N_10129,N_9637);
or U11684 (N_11684,N_9257,N_10161);
xnor U11685 (N_11685,N_9776,N_9026);
and U11686 (N_11686,N_10289,N_9564);
xnor U11687 (N_11687,N_9882,N_9187);
nand U11688 (N_11688,N_9450,N_9226);
or U11689 (N_11689,N_9457,N_9267);
or U11690 (N_11690,N_9914,N_10330);
nor U11691 (N_11691,N_9407,N_9274);
nor U11692 (N_11692,N_10013,N_10054);
nor U11693 (N_11693,N_9838,N_9303);
xnor U11694 (N_11694,N_10484,N_9277);
nor U11695 (N_11695,N_9945,N_9842);
or U11696 (N_11696,N_9864,N_10442);
nand U11697 (N_11697,N_9402,N_9852);
or U11698 (N_11698,N_9491,N_9781);
and U11699 (N_11699,N_10426,N_10264);
and U11700 (N_11700,N_9885,N_10271);
nand U11701 (N_11701,N_9132,N_9303);
and U11702 (N_11702,N_9746,N_9429);
and U11703 (N_11703,N_9343,N_9048);
nand U11704 (N_11704,N_9875,N_9331);
nor U11705 (N_11705,N_10046,N_9423);
nand U11706 (N_11706,N_10220,N_9815);
nand U11707 (N_11707,N_9777,N_9280);
nand U11708 (N_11708,N_10043,N_9687);
or U11709 (N_11709,N_10372,N_10224);
or U11710 (N_11710,N_10361,N_9924);
nor U11711 (N_11711,N_9073,N_9049);
or U11712 (N_11712,N_10478,N_9344);
and U11713 (N_11713,N_10260,N_9135);
or U11714 (N_11714,N_10199,N_10309);
and U11715 (N_11715,N_10357,N_9899);
or U11716 (N_11716,N_10400,N_10198);
and U11717 (N_11717,N_10397,N_10498);
nor U11718 (N_11718,N_9690,N_10469);
xnor U11719 (N_11719,N_10075,N_9770);
and U11720 (N_11720,N_9456,N_10242);
and U11721 (N_11721,N_9517,N_9675);
nand U11722 (N_11722,N_10405,N_10211);
and U11723 (N_11723,N_10114,N_9602);
nand U11724 (N_11724,N_10022,N_10130);
nand U11725 (N_11725,N_9982,N_9827);
xnor U11726 (N_11726,N_10221,N_9896);
nand U11727 (N_11727,N_9127,N_10410);
and U11728 (N_11728,N_9895,N_10464);
nor U11729 (N_11729,N_10341,N_10002);
nor U11730 (N_11730,N_10077,N_9958);
xnor U11731 (N_11731,N_9087,N_9530);
nand U11732 (N_11732,N_9642,N_9017);
nor U11733 (N_11733,N_9010,N_9376);
xnor U11734 (N_11734,N_9029,N_9643);
or U11735 (N_11735,N_10201,N_9764);
and U11736 (N_11736,N_10298,N_9799);
or U11737 (N_11737,N_9905,N_9156);
and U11738 (N_11738,N_9246,N_10453);
xor U11739 (N_11739,N_9823,N_9297);
xnor U11740 (N_11740,N_9140,N_9142);
nor U11741 (N_11741,N_10447,N_10477);
and U11742 (N_11742,N_9440,N_10171);
xor U11743 (N_11743,N_10446,N_10045);
xor U11744 (N_11744,N_9857,N_9137);
xnor U11745 (N_11745,N_10274,N_9400);
and U11746 (N_11746,N_9638,N_9421);
nand U11747 (N_11747,N_9779,N_9587);
and U11748 (N_11748,N_9229,N_9759);
and U11749 (N_11749,N_9178,N_10264);
or U11750 (N_11750,N_9403,N_9430);
or U11751 (N_11751,N_9044,N_9053);
and U11752 (N_11752,N_10319,N_9498);
xnor U11753 (N_11753,N_10026,N_9140);
or U11754 (N_11754,N_9328,N_9544);
and U11755 (N_11755,N_10149,N_10300);
and U11756 (N_11756,N_9070,N_9142);
or U11757 (N_11757,N_9597,N_9426);
xor U11758 (N_11758,N_9681,N_9828);
or U11759 (N_11759,N_9857,N_9834);
and U11760 (N_11760,N_9640,N_10443);
nand U11761 (N_11761,N_10030,N_9591);
nor U11762 (N_11762,N_9203,N_9543);
or U11763 (N_11763,N_9796,N_10235);
and U11764 (N_11764,N_9496,N_10110);
nand U11765 (N_11765,N_10177,N_9527);
or U11766 (N_11766,N_9393,N_9320);
or U11767 (N_11767,N_10132,N_9236);
and U11768 (N_11768,N_9795,N_9762);
nor U11769 (N_11769,N_9558,N_9471);
nor U11770 (N_11770,N_10488,N_9870);
xnor U11771 (N_11771,N_9417,N_9383);
or U11772 (N_11772,N_10349,N_9002);
nor U11773 (N_11773,N_9478,N_10240);
and U11774 (N_11774,N_10243,N_10012);
nand U11775 (N_11775,N_9946,N_10062);
nand U11776 (N_11776,N_9624,N_9462);
nor U11777 (N_11777,N_9151,N_9974);
xnor U11778 (N_11778,N_9577,N_10497);
nand U11779 (N_11779,N_10236,N_9154);
nor U11780 (N_11780,N_10387,N_9321);
nor U11781 (N_11781,N_10234,N_9299);
xnor U11782 (N_11782,N_9661,N_9672);
or U11783 (N_11783,N_9088,N_9310);
nand U11784 (N_11784,N_9546,N_9127);
or U11785 (N_11785,N_10472,N_9724);
nor U11786 (N_11786,N_10180,N_10271);
and U11787 (N_11787,N_9808,N_9641);
nand U11788 (N_11788,N_9049,N_9769);
or U11789 (N_11789,N_9384,N_9142);
xor U11790 (N_11790,N_9897,N_9420);
xnor U11791 (N_11791,N_9808,N_9799);
or U11792 (N_11792,N_10368,N_10028);
nand U11793 (N_11793,N_9035,N_10299);
nor U11794 (N_11794,N_9656,N_10060);
nor U11795 (N_11795,N_10306,N_9456);
nand U11796 (N_11796,N_9724,N_9799);
or U11797 (N_11797,N_9481,N_10191);
nor U11798 (N_11798,N_9880,N_9890);
nand U11799 (N_11799,N_9738,N_10191);
nand U11800 (N_11800,N_9491,N_9107);
nor U11801 (N_11801,N_10102,N_10274);
or U11802 (N_11802,N_9316,N_10119);
nand U11803 (N_11803,N_9576,N_9755);
xor U11804 (N_11804,N_9351,N_9345);
and U11805 (N_11805,N_9218,N_9744);
and U11806 (N_11806,N_10071,N_10355);
xor U11807 (N_11807,N_10183,N_9456);
or U11808 (N_11808,N_9229,N_10163);
xnor U11809 (N_11809,N_10119,N_10306);
xnor U11810 (N_11810,N_9549,N_9709);
xor U11811 (N_11811,N_9783,N_9688);
nor U11812 (N_11812,N_10415,N_9466);
nor U11813 (N_11813,N_9963,N_9972);
nand U11814 (N_11814,N_10341,N_10424);
nor U11815 (N_11815,N_9212,N_9455);
nand U11816 (N_11816,N_9833,N_10160);
xnor U11817 (N_11817,N_9400,N_9922);
nand U11818 (N_11818,N_9996,N_9573);
or U11819 (N_11819,N_10038,N_9127);
and U11820 (N_11820,N_9777,N_9705);
or U11821 (N_11821,N_9744,N_9198);
or U11822 (N_11822,N_9109,N_9358);
nand U11823 (N_11823,N_9878,N_10331);
or U11824 (N_11824,N_9309,N_9426);
xnor U11825 (N_11825,N_9679,N_9639);
and U11826 (N_11826,N_9907,N_9874);
or U11827 (N_11827,N_9516,N_10100);
nor U11828 (N_11828,N_10156,N_10302);
and U11829 (N_11829,N_10229,N_9267);
xnor U11830 (N_11830,N_10111,N_9933);
xor U11831 (N_11831,N_10176,N_9132);
nor U11832 (N_11832,N_10498,N_9419);
nand U11833 (N_11833,N_9065,N_9556);
nand U11834 (N_11834,N_10452,N_10026);
nand U11835 (N_11835,N_9263,N_9935);
or U11836 (N_11836,N_10425,N_10080);
nand U11837 (N_11837,N_9990,N_9960);
or U11838 (N_11838,N_10359,N_10330);
nor U11839 (N_11839,N_9961,N_10302);
nand U11840 (N_11840,N_10309,N_10234);
or U11841 (N_11841,N_9761,N_10435);
nand U11842 (N_11842,N_9507,N_9227);
xnor U11843 (N_11843,N_10055,N_10454);
nor U11844 (N_11844,N_10253,N_9532);
xor U11845 (N_11845,N_10242,N_9708);
or U11846 (N_11846,N_9003,N_9640);
xnor U11847 (N_11847,N_9780,N_9969);
nand U11848 (N_11848,N_10335,N_9972);
xor U11849 (N_11849,N_9293,N_9614);
nor U11850 (N_11850,N_10385,N_9066);
or U11851 (N_11851,N_10277,N_9164);
xnor U11852 (N_11852,N_9312,N_9339);
and U11853 (N_11853,N_9937,N_10332);
xnor U11854 (N_11854,N_9604,N_9954);
nor U11855 (N_11855,N_10139,N_9142);
or U11856 (N_11856,N_9670,N_9513);
or U11857 (N_11857,N_9039,N_9188);
or U11858 (N_11858,N_10083,N_10290);
or U11859 (N_11859,N_9240,N_10413);
or U11860 (N_11860,N_10185,N_9039);
nand U11861 (N_11861,N_9432,N_9354);
nor U11862 (N_11862,N_10469,N_9430);
nand U11863 (N_11863,N_10121,N_9956);
xnor U11864 (N_11864,N_9210,N_9251);
nand U11865 (N_11865,N_9703,N_10464);
and U11866 (N_11866,N_10184,N_9897);
and U11867 (N_11867,N_10395,N_10008);
and U11868 (N_11868,N_9212,N_10405);
nand U11869 (N_11869,N_10224,N_10132);
nor U11870 (N_11870,N_9211,N_10410);
and U11871 (N_11871,N_10435,N_10075);
and U11872 (N_11872,N_9501,N_10199);
xor U11873 (N_11873,N_9434,N_9607);
nand U11874 (N_11874,N_9409,N_9653);
nand U11875 (N_11875,N_9534,N_9839);
and U11876 (N_11876,N_9022,N_9916);
nor U11877 (N_11877,N_10375,N_10257);
nand U11878 (N_11878,N_9758,N_9059);
nand U11879 (N_11879,N_9218,N_9420);
and U11880 (N_11880,N_9118,N_9955);
nor U11881 (N_11881,N_10369,N_9704);
and U11882 (N_11882,N_9531,N_9980);
nand U11883 (N_11883,N_9402,N_10103);
nor U11884 (N_11884,N_10175,N_9917);
or U11885 (N_11885,N_10202,N_9534);
and U11886 (N_11886,N_9459,N_9851);
and U11887 (N_11887,N_9027,N_9501);
or U11888 (N_11888,N_9560,N_9099);
or U11889 (N_11889,N_9735,N_9964);
nand U11890 (N_11890,N_10336,N_9109);
xnor U11891 (N_11891,N_9421,N_9056);
xor U11892 (N_11892,N_10436,N_10167);
xor U11893 (N_11893,N_9984,N_9970);
and U11894 (N_11894,N_9077,N_9993);
xor U11895 (N_11895,N_9361,N_9750);
xnor U11896 (N_11896,N_10062,N_9696);
nand U11897 (N_11897,N_10459,N_9850);
nor U11898 (N_11898,N_9364,N_10472);
nor U11899 (N_11899,N_9605,N_9302);
nand U11900 (N_11900,N_10362,N_9264);
nor U11901 (N_11901,N_9255,N_9523);
and U11902 (N_11902,N_9458,N_9271);
or U11903 (N_11903,N_10179,N_10482);
and U11904 (N_11904,N_9383,N_9882);
or U11905 (N_11905,N_9994,N_9466);
xor U11906 (N_11906,N_9648,N_10074);
xnor U11907 (N_11907,N_10119,N_10477);
xnor U11908 (N_11908,N_9664,N_10267);
nand U11909 (N_11909,N_9552,N_9233);
nor U11910 (N_11910,N_9304,N_9427);
nand U11911 (N_11911,N_10309,N_9538);
xor U11912 (N_11912,N_10092,N_9742);
xnor U11913 (N_11913,N_10204,N_9784);
nor U11914 (N_11914,N_9768,N_9786);
or U11915 (N_11915,N_9138,N_10022);
xor U11916 (N_11916,N_9392,N_9993);
nor U11917 (N_11917,N_9600,N_9494);
nand U11918 (N_11918,N_10304,N_9890);
and U11919 (N_11919,N_9405,N_10132);
nor U11920 (N_11920,N_10016,N_9148);
xor U11921 (N_11921,N_9521,N_9112);
xnor U11922 (N_11922,N_10288,N_10404);
xor U11923 (N_11923,N_10135,N_9405);
or U11924 (N_11924,N_9781,N_9147);
nand U11925 (N_11925,N_10489,N_9270);
nand U11926 (N_11926,N_9815,N_10351);
nand U11927 (N_11927,N_10123,N_10495);
or U11928 (N_11928,N_9767,N_10106);
nand U11929 (N_11929,N_9763,N_9639);
and U11930 (N_11930,N_10157,N_9282);
xor U11931 (N_11931,N_10371,N_9052);
and U11932 (N_11932,N_10266,N_9186);
nor U11933 (N_11933,N_9727,N_9721);
nand U11934 (N_11934,N_10314,N_9064);
xnor U11935 (N_11935,N_9208,N_9428);
and U11936 (N_11936,N_10056,N_10363);
nor U11937 (N_11937,N_10168,N_10133);
or U11938 (N_11938,N_10088,N_10114);
nand U11939 (N_11939,N_9270,N_9923);
nor U11940 (N_11940,N_9283,N_10358);
xnor U11941 (N_11941,N_9183,N_10179);
or U11942 (N_11942,N_10479,N_10202);
and U11943 (N_11943,N_9077,N_9920);
and U11944 (N_11944,N_9028,N_9200);
or U11945 (N_11945,N_10394,N_9724);
xor U11946 (N_11946,N_9080,N_9849);
or U11947 (N_11947,N_9610,N_9546);
and U11948 (N_11948,N_10357,N_9502);
or U11949 (N_11949,N_9367,N_9778);
and U11950 (N_11950,N_10221,N_9663);
nor U11951 (N_11951,N_10075,N_9840);
nand U11952 (N_11952,N_10119,N_9381);
xor U11953 (N_11953,N_9204,N_10280);
and U11954 (N_11954,N_9836,N_9066);
nor U11955 (N_11955,N_9515,N_9812);
nor U11956 (N_11956,N_9312,N_9954);
or U11957 (N_11957,N_9381,N_9100);
nand U11958 (N_11958,N_9760,N_10288);
and U11959 (N_11959,N_9157,N_9270);
and U11960 (N_11960,N_10404,N_9044);
or U11961 (N_11961,N_10102,N_9370);
nand U11962 (N_11962,N_9508,N_9672);
or U11963 (N_11963,N_9739,N_10403);
xnor U11964 (N_11964,N_9449,N_9902);
xnor U11965 (N_11965,N_9644,N_10035);
xor U11966 (N_11966,N_10173,N_9707);
nor U11967 (N_11967,N_9225,N_9272);
and U11968 (N_11968,N_9700,N_9623);
and U11969 (N_11969,N_9197,N_10001);
nor U11970 (N_11970,N_9285,N_9635);
nand U11971 (N_11971,N_9108,N_10252);
xnor U11972 (N_11972,N_9664,N_9969);
or U11973 (N_11973,N_9070,N_10176);
nand U11974 (N_11974,N_10005,N_9540);
nor U11975 (N_11975,N_9048,N_10288);
nand U11976 (N_11976,N_10107,N_9523);
xor U11977 (N_11977,N_9091,N_9537);
and U11978 (N_11978,N_9914,N_9938);
or U11979 (N_11979,N_9978,N_9234);
xnor U11980 (N_11980,N_10385,N_9164);
xor U11981 (N_11981,N_10107,N_9049);
xor U11982 (N_11982,N_10070,N_10443);
nor U11983 (N_11983,N_10199,N_9969);
nand U11984 (N_11984,N_10356,N_10346);
xor U11985 (N_11985,N_10385,N_9139);
nor U11986 (N_11986,N_9188,N_9537);
nand U11987 (N_11987,N_9286,N_9928);
xor U11988 (N_11988,N_10041,N_9060);
nand U11989 (N_11989,N_9736,N_10125);
nor U11990 (N_11990,N_9325,N_9165);
nor U11991 (N_11991,N_9953,N_9143);
or U11992 (N_11992,N_9897,N_9639);
or U11993 (N_11993,N_9660,N_9220);
xor U11994 (N_11994,N_9978,N_9067);
nor U11995 (N_11995,N_9393,N_10157);
or U11996 (N_11996,N_10364,N_10333);
or U11997 (N_11997,N_9710,N_9245);
nor U11998 (N_11998,N_10266,N_10212);
and U11999 (N_11999,N_10035,N_9663);
or U12000 (N_12000,N_11530,N_10765);
xnor U12001 (N_12001,N_11957,N_11855);
or U12002 (N_12002,N_11579,N_10564);
and U12003 (N_12003,N_11978,N_11129);
xnor U12004 (N_12004,N_11370,N_11410);
nor U12005 (N_12005,N_10995,N_10788);
and U12006 (N_12006,N_10710,N_11954);
nor U12007 (N_12007,N_11486,N_10639);
xor U12008 (N_12008,N_11171,N_11895);
nor U12009 (N_12009,N_11438,N_11427);
and U12010 (N_12010,N_11386,N_11284);
nand U12011 (N_12011,N_10735,N_11613);
or U12012 (N_12012,N_10692,N_11392);
nand U12013 (N_12013,N_10634,N_11545);
nand U12014 (N_12014,N_10928,N_11909);
nor U12015 (N_12015,N_11308,N_11040);
and U12016 (N_12016,N_11341,N_11583);
nor U12017 (N_12017,N_11446,N_11749);
xnor U12018 (N_12018,N_11272,N_11698);
or U12019 (N_12019,N_11282,N_11226);
xnor U12020 (N_12020,N_11679,N_11873);
and U12021 (N_12021,N_11373,N_10570);
nor U12022 (N_12022,N_11293,N_11290);
or U12023 (N_12023,N_11215,N_10610);
xnor U12024 (N_12024,N_11696,N_10693);
and U12025 (N_12025,N_11300,N_11629);
or U12026 (N_12026,N_11585,N_11265);
or U12027 (N_12027,N_10559,N_11607);
xnor U12028 (N_12028,N_10591,N_10526);
xor U12029 (N_12029,N_11317,N_11376);
and U12030 (N_12030,N_11510,N_11221);
and U12031 (N_12031,N_11884,N_11405);
or U12032 (N_12032,N_11496,N_11952);
xor U12033 (N_12033,N_10757,N_11224);
or U12034 (N_12034,N_11866,N_11720);
or U12035 (N_12035,N_11563,N_11186);
or U12036 (N_12036,N_11925,N_10956);
nor U12037 (N_12037,N_10912,N_11942);
nor U12038 (N_12038,N_11092,N_11628);
nor U12039 (N_12039,N_10791,N_11707);
xor U12040 (N_12040,N_11469,N_10764);
nor U12041 (N_12041,N_11618,N_10797);
nand U12042 (N_12042,N_11258,N_11653);
xnor U12043 (N_12043,N_11702,N_11677);
nand U12044 (N_12044,N_11437,N_11649);
and U12045 (N_12045,N_11753,N_11595);
nand U12046 (N_12046,N_11366,N_11149);
or U12047 (N_12047,N_11087,N_10961);
or U12048 (N_12048,N_11778,N_10923);
xor U12049 (N_12049,N_10958,N_11984);
nor U12050 (N_12050,N_11274,N_11870);
nand U12051 (N_12051,N_10972,N_11908);
or U12052 (N_12052,N_10677,N_11935);
nand U12053 (N_12053,N_11863,N_10608);
nor U12054 (N_12054,N_11097,N_11923);
nand U12055 (N_12055,N_11192,N_10846);
nand U12056 (N_12056,N_11830,N_11104);
or U12057 (N_12057,N_11448,N_11782);
nor U12058 (N_12058,N_11736,N_11632);
nand U12059 (N_12059,N_10770,N_11877);
nand U12060 (N_12060,N_10986,N_11899);
or U12061 (N_12061,N_11795,N_11523);
or U12062 (N_12062,N_10720,N_11304);
xor U12063 (N_12063,N_10784,N_11671);
and U12064 (N_12064,N_11881,N_11484);
nor U12065 (N_12065,N_10800,N_10992);
xor U12066 (N_12066,N_11587,N_10704);
xor U12067 (N_12067,N_11350,N_11540);
or U12068 (N_12068,N_11959,N_11663);
or U12069 (N_12069,N_10857,N_11703);
nor U12070 (N_12070,N_11482,N_11344);
and U12071 (N_12071,N_10917,N_11686);
nor U12072 (N_12072,N_11754,N_11497);
nand U12073 (N_12073,N_10563,N_10707);
nand U12074 (N_12074,N_11651,N_11614);
or U12075 (N_12075,N_10970,N_11483);
nor U12076 (N_12076,N_10867,N_11365);
or U12077 (N_12077,N_11139,N_11385);
or U12078 (N_12078,N_10853,N_10967);
and U12079 (N_12079,N_10814,N_11478);
or U12080 (N_12080,N_11112,N_10924);
and U12081 (N_12081,N_11006,N_11283);
xor U12082 (N_12082,N_11231,N_10577);
nor U12083 (N_12083,N_11612,N_11352);
nor U12084 (N_12084,N_11023,N_11557);
or U12085 (N_12085,N_11126,N_10776);
nand U12086 (N_12086,N_10925,N_10687);
xor U12087 (N_12087,N_11460,N_11211);
nand U12088 (N_12088,N_10521,N_11177);
xor U12089 (N_12089,N_10511,N_11903);
xnor U12090 (N_12090,N_11603,N_11644);
or U12091 (N_12091,N_11569,N_11798);
and U12092 (N_12092,N_10531,N_11291);
xnor U12093 (N_12093,N_10843,N_11475);
xor U12094 (N_12094,N_11159,N_11277);
xor U12095 (N_12095,N_11132,N_10918);
nor U12096 (N_12096,N_11039,N_11229);
nor U12097 (N_12097,N_10840,N_11154);
nand U12098 (N_12098,N_11489,N_11916);
nand U12099 (N_12099,N_10805,N_10790);
nand U12100 (N_12100,N_10848,N_11917);
xnor U12101 (N_12101,N_11787,N_11025);
or U12102 (N_12102,N_11718,N_10562);
nand U12103 (N_12103,N_11334,N_11145);
nand U12104 (N_12104,N_11941,N_10951);
and U12105 (N_12105,N_10860,N_11044);
or U12106 (N_12106,N_11416,N_11988);
xnor U12107 (N_12107,N_11289,N_11592);
nor U12108 (N_12108,N_10502,N_10593);
or U12109 (N_12109,N_11577,N_10963);
or U12110 (N_12110,N_11180,N_11949);
nor U12111 (N_12111,N_10982,N_10506);
xnor U12112 (N_12112,N_11528,N_11424);
nor U12113 (N_12113,N_11161,N_10510);
nand U12114 (N_12114,N_10609,N_10754);
xnor U12115 (N_12115,N_11374,N_11433);
xnor U12116 (N_12116,N_11281,N_10618);
nor U12117 (N_12117,N_11826,N_11989);
nand U12118 (N_12118,N_10552,N_11662);
or U12119 (N_12119,N_11306,N_11885);
xnor U12120 (N_12120,N_11355,N_11791);
nand U12121 (N_12121,N_11425,N_10883);
nor U12122 (N_12122,N_11847,N_10786);
and U12123 (N_12123,N_10539,N_10603);
or U12124 (N_12124,N_10695,N_11983);
nor U12125 (N_12125,N_11522,N_11999);
or U12126 (N_12126,N_11635,N_10597);
xor U12127 (N_12127,N_10568,N_11248);
xor U12128 (N_12128,N_11889,N_10650);
nand U12129 (N_12129,N_11393,N_11359);
nor U12130 (N_12130,N_10894,N_11319);
or U12131 (N_12131,N_11842,N_10755);
or U12132 (N_12132,N_11368,N_11075);
nor U12133 (N_12133,N_11774,N_11403);
or U12134 (N_12134,N_10738,N_11953);
nor U12135 (N_12135,N_10761,N_10689);
nor U12136 (N_12136,N_11656,N_11764);
xnor U12137 (N_12137,N_10922,N_11822);
nor U12138 (N_12138,N_11252,N_11314);
xnor U12139 (N_12139,N_11046,N_11975);
or U12140 (N_12140,N_11750,N_11426);
nor U12141 (N_12141,N_11580,N_11914);
nor U12142 (N_12142,N_11665,N_11088);
nand U12143 (N_12143,N_11067,N_11198);
or U12144 (N_12144,N_11835,N_11379);
nor U12145 (N_12145,N_10808,N_10512);
nand U12146 (N_12146,N_10914,N_11115);
or U12147 (N_12147,N_11806,N_11553);
or U12148 (N_12148,N_10891,N_11387);
nor U12149 (N_12149,N_10777,N_11243);
nor U12150 (N_12150,N_11779,N_10582);
nand U12151 (N_12151,N_10719,N_11167);
nand U12152 (N_12152,N_10679,N_11449);
or U12153 (N_12153,N_11737,N_11467);
nor U12154 (N_12154,N_11432,N_11071);
and U12155 (N_12155,N_10826,N_11270);
and U12156 (N_12156,N_11105,N_10709);
and U12157 (N_12157,N_10850,N_11652);
xnor U12158 (N_12158,N_10722,N_11819);
or U12159 (N_12159,N_10642,N_11814);
or U12160 (N_12160,N_10876,N_10927);
nand U12161 (N_12161,N_11588,N_10561);
nand U12162 (N_12162,N_11458,N_11054);
xor U12163 (N_12163,N_10994,N_11372);
nor U12164 (N_12164,N_11242,N_11173);
xor U12165 (N_12165,N_11454,N_11421);
or U12166 (N_12166,N_11584,N_10630);
and U12167 (N_12167,N_11758,N_10999);
and U12168 (N_12168,N_11148,N_11709);
or U12169 (N_12169,N_11578,N_11419);
and U12170 (N_12170,N_11951,N_11896);
nor U12171 (N_12171,N_10783,N_11943);
and U12172 (N_12172,N_10656,N_11086);
nand U12173 (N_12173,N_10533,N_11622);
or U12174 (N_12174,N_11422,N_10955);
nor U12175 (N_12175,N_10948,N_11253);
or U12176 (N_12176,N_11381,N_11061);
nand U12177 (N_12177,N_11843,N_10964);
xnor U12178 (N_12178,N_11768,N_11364);
and U12179 (N_12179,N_11331,N_10872);
or U12180 (N_12180,N_11049,N_10515);
and U12181 (N_12181,N_11945,N_11727);
and U12182 (N_12182,N_11269,N_11853);
xor U12183 (N_12183,N_11207,N_11670);
nand U12184 (N_12184,N_10910,N_11028);
or U12185 (N_12185,N_11190,N_11034);
or U12186 (N_12186,N_10694,N_11157);
xnor U12187 (N_12187,N_10688,N_11911);
and U12188 (N_12188,N_11800,N_11770);
or U12189 (N_12189,N_11777,N_11122);
or U12190 (N_12190,N_11986,N_10621);
and U12191 (N_12191,N_11982,N_11558);
nor U12192 (N_12192,N_10648,N_11659);
and U12193 (N_12193,N_10957,N_11803);
and U12194 (N_12194,N_11719,N_11815);
xnor U12195 (N_12195,N_10904,N_11246);
xor U12196 (N_12196,N_11055,N_11078);
nand U12197 (N_12197,N_11776,N_11820);
nand U12198 (N_12198,N_11222,N_10852);
nand U12199 (N_12199,N_11333,N_11928);
or U12200 (N_12200,N_10638,N_11516);
and U12201 (N_12201,N_10525,N_11851);
nor U12202 (N_12202,N_11195,N_10941);
nor U12203 (N_12203,N_10553,N_11623);
xor U12204 (N_12204,N_11546,N_11029);
and U12205 (N_12205,N_11409,N_10520);
and U12206 (N_12206,N_10571,N_10595);
or U12207 (N_12207,N_11840,N_10729);
and U12208 (N_12208,N_11008,N_11176);
nor U12209 (N_12209,N_11919,N_11309);
and U12210 (N_12210,N_10641,N_11763);
nand U12211 (N_12211,N_11690,N_10888);
nand U12212 (N_12212,N_11726,N_11429);
nor U12213 (N_12213,N_11940,N_11748);
or U12214 (N_12214,N_11048,N_11996);
and U12215 (N_12215,N_11642,N_10815);
nand U12216 (N_12216,N_10979,N_11133);
nand U12217 (N_12217,N_11094,N_11450);
nor U12218 (N_12218,N_10816,N_10651);
and U12219 (N_12219,N_11538,N_11435);
or U12220 (N_12220,N_10858,N_11712);
nor U12221 (N_12221,N_11453,N_11684);
or U12222 (N_12222,N_10943,N_11031);
nor U12223 (N_12223,N_11688,N_11116);
nand U12224 (N_12224,N_11481,N_11856);
or U12225 (N_12225,N_11608,N_10991);
and U12226 (N_12226,N_11414,N_10885);
xnor U12227 (N_12227,N_11339,N_11152);
xor U12228 (N_12228,N_11740,N_11747);
and U12229 (N_12229,N_11692,N_10529);
and U12230 (N_12230,N_11020,N_11883);
and U12231 (N_12231,N_11428,N_10793);
nor U12232 (N_12232,N_11871,N_11893);
xnor U12233 (N_12233,N_10895,N_11415);
xor U12234 (N_12234,N_10551,N_11168);
nand U12235 (N_12235,N_11160,N_11490);
nand U12236 (N_12236,N_11328,N_11643);
xor U12237 (N_12237,N_11661,N_11135);
and U12238 (N_12238,N_11199,N_11297);
nand U12239 (N_12239,N_11637,N_11348);
nand U12240 (N_12240,N_11600,N_11487);
nor U12241 (N_12241,N_11119,N_10589);
and U12242 (N_12242,N_10817,N_10574);
nor U12243 (N_12243,N_10949,N_10666);
and U12244 (N_12244,N_10897,N_11236);
nand U12245 (N_12245,N_10792,N_11107);
nand U12246 (N_12246,N_11744,N_11461);
nand U12247 (N_12247,N_11804,N_11706);
and U12248 (N_12248,N_11839,N_11205);
and U12249 (N_12249,N_11302,N_11465);
xnor U12250 (N_12250,N_10717,N_11194);
and U12251 (N_12251,N_11441,N_10643);
nand U12252 (N_12252,N_11861,N_11468);
xor U12253 (N_12253,N_10600,N_11455);
and U12254 (N_12254,N_11687,N_10960);
nor U12255 (N_12255,N_10683,N_11743);
nor U12256 (N_12256,N_10810,N_11369);
xor U12257 (N_12257,N_11247,N_11756);
nand U12258 (N_12258,N_10742,N_11052);
and U12259 (N_12259,N_11666,N_11882);
xnor U12260 (N_12260,N_11164,N_11858);
nor U12261 (N_12261,N_11346,N_10624);
nand U12262 (N_12262,N_11472,N_10973);
nand U12263 (N_12263,N_11683,N_11298);
nor U12264 (N_12264,N_10522,N_11412);
and U12265 (N_12265,N_11930,N_10833);
or U12266 (N_12266,N_10708,N_11110);
and U12267 (N_12267,N_11664,N_11491);
xnor U12268 (N_12268,N_11638,N_10746);
nand U12269 (N_12269,N_10567,N_11076);
xnor U12270 (N_12270,N_11203,N_11144);
and U12271 (N_12271,N_10803,N_10959);
nor U12272 (N_12272,N_10987,N_11509);
nand U12273 (N_12273,N_11358,N_11728);
xor U12274 (N_12274,N_11069,N_10845);
nor U12275 (N_12275,N_10988,N_11009);
nand U12276 (N_12276,N_11033,N_10901);
nor U12277 (N_12277,N_11431,N_10580);
nand U12278 (N_12278,N_11507,N_11760);
or U12279 (N_12279,N_11762,N_11811);
or U12280 (N_12280,N_11556,N_11354);
or U12281 (N_12281,N_10727,N_11675);
nor U12282 (N_12282,N_11479,N_11193);
nor U12283 (N_12283,N_11170,N_10716);
xor U12284 (N_12284,N_10646,N_11977);
nor U12285 (N_12285,N_11485,N_11147);
and U12286 (N_12286,N_11506,N_10818);
nor U12287 (N_12287,N_11375,N_10667);
nor U12288 (N_12288,N_11011,N_11402);
nor U12289 (N_12289,N_10737,N_11775);
and U12290 (N_12290,N_11920,N_11615);
xor U12291 (N_12291,N_10665,N_10605);
and U12292 (N_12292,N_10745,N_11138);
xnor U12293 (N_12293,N_10534,N_11322);
nor U12294 (N_12294,N_10940,N_11705);
nand U12295 (N_12295,N_11827,N_10601);
nand U12296 (N_12296,N_10868,N_11567);
xnor U12297 (N_12297,N_10678,N_11464);
xnor U12298 (N_12298,N_10753,N_11810);
xor U12299 (N_12299,N_11970,N_10756);
and U12300 (N_12300,N_11178,N_10513);
xor U12301 (N_12301,N_11275,N_10696);
and U12302 (N_12302,N_11910,N_11561);
nand U12303 (N_12303,N_10664,N_11095);
nand U12304 (N_12304,N_10977,N_10732);
nand U12305 (N_12305,N_11751,N_11947);
nand U12306 (N_12306,N_10996,N_11459);
nor U12307 (N_12307,N_10806,N_11276);
xnor U12308 (N_12308,N_10544,N_10887);
and U12309 (N_12309,N_11723,N_10906);
xnor U12310 (N_12310,N_10673,N_11807);
or U12311 (N_12311,N_11278,N_11257);
and U12312 (N_12312,N_10637,N_11058);
nor U12313 (N_12313,N_11016,N_11267);
or U12314 (N_12314,N_11394,N_11197);
nand U12315 (N_12315,N_11239,N_10975);
xor U12316 (N_12316,N_10672,N_11150);
xor U12317 (N_12317,N_10881,N_10557);
nor U12318 (N_12318,N_11955,N_10911);
nor U12319 (N_12319,N_10950,N_11508);
or U12320 (N_12320,N_11525,N_10590);
nand U12321 (N_12321,N_11901,N_11254);
nor U12322 (N_12322,N_10524,N_10532);
or U12323 (N_12323,N_11013,N_10844);
and U12324 (N_12324,N_10863,N_11187);
nor U12325 (N_12325,N_10985,N_11003);
or U12326 (N_12326,N_11624,N_11792);
nor U12327 (N_12327,N_11127,N_10527);
nor U12328 (N_12328,N_11733,N_10538);
or U12329 (N_12329,N_11445,N_11788);
and U12330 (N_12330,N_10584,N_10581);
and U12331 (N_12331,N_11539,N_11141);
nor U12332 (N_12332,N_10825,N_11391);
and U12333 (N_12333,N_10938,N_10890);
nor U12334 (N_12334,N_10997,N_10744);
xor U12335 (N_12335,N_11109,N_11918);
nor U12336 (N_12336,N_10668,N_11351);
nor U12337 (N_12337,N_11336,N_10715);
and U12338 (N_12338,N_11862,N_10530);
or U12339 (N_12339,N_10655,N_11555);
or U12340 (N_12340,N_10620,N_11596);
nor U12341 (N_12341,N_11759,N_11695);
nor U12342 (N_12342,N_11413,N_11010);
nand U12343 (N_12343,N_11390,N_11828);
and U12344 (N_12344,N_11256,N_11238);
xnor U12345 (N_12345,N_11301,N_11906);
or U12346 (N_12346,N_11627,N_10705);
and U12347 (N_12347,N_11059,N_11832);
and U12348 (N_12348,N_11090,N_11262);
and U12349 (N_12349,N_10774,N_10751);
or U12350 (N_12350,N_11991,N_11174);
xnor U12351 (N_12351,N_10896,N_11140);
or U12352 (N_12352,N_10905,N_10962);
nor U12353 (N_12353,N_11755,N_11724);
xnor U12354 (N_12354,N_11880,N_11681);
or U12355 (N_12355,N_11565,N_11500);
nor U12356 (N_12356,N_11316,N_11227);
xnor U12357 (N_12357,N_11400,N_11879);
and U12358 (N_12358,N_10821,N_10528);
nand U12359 (N_12359,N_11401,N_11691);
nor U12360 (N_12360,N_11844,N_10886);
and U12361 (N_12361,N_11047,N_11206);
nand U12362 (N_12362,N_11700,N_11713);
nand U12363 (N_12363,N_11674,N_11717);
or U12364 (N_12364,N_11566,N_10739);
xor U12365 (N_12365,N_11273,N_10752);
nand U12366 (N_12366,N_11096,N_11318);
and U12367 (N_12367,N_11255,N_10615);
xor U12368 (N_12368,N_11225,N_10795);
and U12369 (N_12369,N_11846,N_11894);
and U12370 (N_12370,N_11151,N_10965);
nand U12371 (N_12371,N_11590,N_11418);
nor U12372 (N_12372,N_11646,N_10837);
xor U12373 (N_12373,N_11241,N_10968);
and U12374 (N_12374,N_11022,N_11406);
nand U12375 (N_12375,N_10781,N_11867);
nor U12376 (N_12376,N_11451,N_11915);
or U12377 (N_12377,N_11905,N_11388);
nand U12378 (N_12378,N_10907,N_11572);
nor U12379 (N_12379,N_11377,N_10789);
or U12380 (N_12380,N_11630,N_10594);
xnor U12381 (N_12381,N_10546,N_11956);
xnor U12382 (N_12382,N_11875,N_11992);
nor U12383 (N_12383,N_11968,N_10658);
xor U12384 (N_12384,N_10542,N_11074);
nor U12385 (N_12385,N_10903,N_11136);
nor U12386 (N_12386,N_11515,N_10983);
nor U12387 (N_12387,N_10588,N_11601);
xor U12388 (N_12388,N_11347,N_11650);
and U12389 (N_12389,N_11594,N_11101);
nor U12390 (N_12390,N_11974,N_11120);
nand U12391 (N_12391,N_11188,N_11326);
or U12392 (N_12392,N_11605,N_11250);
nor U12393 (N_12393,N_11361,N_11311);
nand U12394 (N_12394,N_11710,N_10740);
nor U12395 (N_12395,N_11362,N_11155);
and U12396 (N_12396,N_11073,N_11327);
nand U12397 (N_12397,N_11480,N_11384);
nand U12398 (N_12398,N_11837,N_11091);
nor U12399 (N_12399,N_10750,N_11551);
nor U12400 (N_12400,N_10933,N_10700);
nor U12401 (N_12401,N_11548,N_10697);
xnor U12402 (N_12402,N_10640,N_11541);
xor U12403 (N_12403,N_10856,N_10909);
or U12404 (N_12404,N_10782,N_10878);
or U12405 (N_12405,N_11876,N_11019);
nor U12406 (N_12406,N_10550,N_11746);
or U12407 (N_12407,N_11493,N_10935);
nor U12408 (N_12408,N_10686,N_10766);
nand U12409 (N_12409,N_10760,N_10902);
and U12410 (N_12410,N_11654,N_11156);
xor U12411 (N_12411,N_10623,N_11153);
and U12412 (N_12412,N_11018,N_10939);
xnor U12413 (N_12413,N_11823,N_10644);
or U12414 (N_12414,N_11473,N_10827);
and U12415 (N_12415,N_11817,N_10811);
and U12416 (N_12416,N_11244,N_10645);
nand U12417 (N_12417,N_10990,N_10587);
or U12418 (N_12418,N_11868,N_10952);
xor U12419 (N_12419,N_11179,N_11320);
and U12420 (N_12420,N_11589,N_11564);
and U12421 (N_12421,N_11356,N_10505);
nand U12422 (N_12422,N_10734,N_10796);
nor U12423 (N_12423,N_11985,N_11735);
nor U12424 (N_12424,N_11602,N_11442);
nand U12425 (N_12425,N_10543,N_11694);
and U12426 (N_12426,N_10824,N_11398);
xnor U12427 (N_12427,N_11371,N_11002);
nor U12428 (N_12428,N_11172,N_11345);
nor U12429 (N_12429,N_11338,N_11471);
or U12430 (N_12430,N_11738,N_11793);
or U12431 (N_12431,N_11066,N_10675);
or U12432 (N_12432,N_11447,N_11444);
nor U12433 (N_12433,N_11813,N_11617);
xor U12434 (N_12434,N_10947,N_11032);
nor U12435 (N_12435,N_11072,N_11980);
nand U12436 (N_12436,N_10540,N_11981);
nand U12437 (N_12437,N_10676,N_10978);
xor U12438 (N_12438,N_11685,N_10743);
nand U12439 (N_12439,N_11382,N_11891);
and U12440 (N_12440,N_11079,N_11730);
nand U12441 (N_12441,N_11513,N_11669);
xnor U12442 (N_12442,N_11268,N_11201);
or U12443 (N_12443,N_11850,N_10976);
xnor U12444 (N_12444,N_11969,N_11597);
nor U12445 (N_12445,N_10613,N_11315);
or U12446 (N_12446,N_11944,N_11781);
and U12447 (N_12447,N_11783,N_10578);
or U12448 (N_12448,N_11900,N_11537);
nor U12449 (N_12449,N_11640,N_10864);
nand U12450 (N_12450,N_11544,N_10920);
nand U12451 (N_12451,N_11208,N_11734);
and U12452 (N_12452,N_10617,N_10627);
nand U12453 (N_12453,N_10839,N_10779);
and U12454 (N_12454,N_10622,N_11294);
nor U12455 (N_12455,N_11488,N_11082);
nor U12456 (N_12456,N_11216,N_11964);
or U12457 (N_12457,N_10579,N_10998);
or U12458 (N_12458,N_11125,N_11801);
xnor U12459 (N_12459,N_11742,N_11950);
or U12460 (N_12460,N_10892,N_11196);
nor U12461 (N_12461,N_10865,N_10565);
nor U12462 (N_12462,N_10701,N_10820);
and U12463 (N_12463,N_11799,N_11098);
nor U12464 (N_12464,N_11307,N_11474);
or U12465 (N_12465,N_11568,N_10741);
nand U12466 (N_12466,N_10758,N_10780);
nand U12467 (N_12467,N_10984,N_11083);
xnor U12468 (N_12468,N_10851,N_11611);
nand U12469 (N_12469,N_11816,N_10969);
xnor U12470 (N_12470,N_11535,N_11030);
and U12471 (N_12471,N_11062,N_11360);
nand U12472 (N_12472,N_11921,N_11864);
xnor U12473 (N_12473,N_10953,N_11021);
nor U12474 (N_12474,N_11542,N_11505);
and U12475 (N_12475,N_11404,N_11966);
or U12476 (N_12476,N_10893,N_11926);
nand U12477 (N_12477,N_11521,N_11305);
and U12478 (N_12478,N_10736,N_11299);
nand U12479 (N_12479,N_10592,N_11693);
nor U12480 (N_12480,N_11860,N_11765);
xor U12481 (N_12481,N_11027,N_10616);
or U12482 (N_12482,N_11869,N_10828);
and U12483 (N_12483,N_11184,N_10849);
nor U12484 (N_12484,N_10931,N_11007);
nor U12485 (N_12485,N_11796,N_11279);
nor U12486 (N_12486,N_11708,N_11888);
nand U12487 (N_12487,N_11210,N_10822);
xor U12488 (N_12488,N_11439,N_10596);
or U12489 (N_12489,N_11859,N_11310);
and U12490 (N_12490,N_11731,N_11068);
xor U12491 (N_12491,N_11631,N_11503);
nor U12492 (N_12492,N_10768,N_11518);
nand U12493 (N_12493,N_11619,N_10921);
nor U12494 (N_12494,N_11367,N_11939);
xnor U12495 (N_12495,N_11892,N_10611);
xor U12496 (N_12496,N_11288,N_11128);
nand U12497 (N_12497,N_11220,N_10898);
and U12498 (N_12498,N_11053,N_11845);
and U12499 (N_12499,N_11504,N_10838);
xnor U12500 (N_12500,N_11938,N_11111);
xor U12501 (N_12501,N_10554,N_11610);
xor U12502 (N_12502,N_11263,N_11636);
nor U12503 (N_12503,N_11045,N_11245);
xnor U12504 (N_12504,N_11711,N_10971);
nand U12505 (N_12505,N_10674,N_10670);
nand U12506 (N_12506,N_10682,N_11961);
xnor U12507 (N_12507,N_11958,N_11051);
nor U12508 (N_12508,N_10547,N_11993);
and U12509 (N_12509,N_10749,N_11704);
nor U12510 (N_12510,N_11492,N_11934);
and U12511 (N_12511,N_11181,N_10555);
nand U12512 (N_12512,N_11434,N_11142);
or U12513 (N_12513,N_11185,N_11233);
or U12514 (N_12514,N_11794,N_11000);
and U12515 (N_12515,N_11946,N_11511);
xor U12516 (N_12516,N_10787,N_11512);
and U12517 (N_12517,N_11499,N_11552);
and U12518 (N_12518,N_11532,N_10718);
nor U12519 (N_12519,N_10929,N_10871);
or U12520 (N_12520,N_10514,N_11162);
nand U12521 (N_12521,N_11324,N_11189);
xnor U12522 (N_12522,N_10807,N_11353);
nand U12523 (N_12523,N_11634,N_10767);
and U12524 (N_12524,N_10874,N_11739);
nor U12525 (N_12525,N_11990,N_11725);
nor U12526 (N_12526,N_11621,N_10647);
nand U12527 (N_12527,N_10813,N_10945);
xnor U12528 (N_12528,N_10763,N_11312);
or U12529 (N_12529,N_11056,N_10930);
or U12530 (N_12530,N_11191,N_11829);
or U12531 (N_12531,N_10919,N_11036);
and U12532 (N_12532,N_11886,N_10536);
nor U12533 (N_12533,N_11337,N_11824);
nand U12534 (N_12534,N_10775,N_11080);
nor U12535 (N_12535,N_11085,N_11536);
xor U12536 (N_12536,N_11280,N_11838);
xnor U12537 (N_12537,N_11772,N_11113);
nor U12538 (N_12538,N_10632,N_11924);
xor U12539 (N_12539,N_10836,N_11100);
xnor U12540 (N_12540,N_11395,N_11766);
or U12541 (N_12541,N_11099,N_11012);
nand U12542 (N_12542,N_11714,N_10690);
nand U12543 (N_12543,N_11527,N_11213);
or U12544 (N_12544,N_11531,N_11645);
nand U12545 (N_12545,N_10569,N_11854);
and U12546 (N_12546,N_11626,N_10660);
nand U12547 (N_12547,N_11330,N_10944);
nand U12548 (N_12548,N_10516,N_10654);
nor U12549 (N_12549,N_11604,N_10908);
or U12550 (N_12550,N_10733,N_11780);
and U12551 (N_12551,N_10915,N_11495);
or U12552 (N_12552,N_10832,N_11973);
xnor U12553 (N_12553,N_11502,N_10942);
and U12554 (N_12554,N_10572,N_10875);
nor U12555 (N_12555,N_10604,N_10989);
or U12556 (N_12556,N_11785,N_11466);
or U12557 (N_12557,N_10537,N_11907);
nor U12558 (N_12558,N_11108,N_10711);
and U12559 (N_12559,N_11689,N_10669);
and U12560 (N_12560,N_11575,N_11084);
or U12561 (N_12561,N_11209,N_11633);
xnor U12562 (N_12562,N_11722,N_11929);
xnor U12563 (N_12563,N_10771,N_10649);
xor U12564 (N_12564,N_11967,N_10862);
xnor U12565 (N_12565,N_11560,N_11660);
xor U12566 (N_12566,N_11325,N_11463);
nand U12567 (N_12567,N_11976,N_11573);
or U12568 (N_12568,N_10517,N_11303);
and U12569 (N_12569,N_11070,N_10798);
xnor U12570 (N_12570,N_11625,N_11285);
xor U12571 (N_12571,N_10794,N_10713);
xor U12572 (N_12572,N_11332,N_11313);
xnor U12573 (N_12573,N_11146,N_10819);
nand U12574 (N_12574,N_10772,N_10731);
and U12575 (N_12575,N_11223,N_11732);
nor U12576 (N_12576,N_11103,N_10831);
nand U12577 (N_12577,N_10899,N_11790);
nand U12578 (N_12578,N_11658,N_11296);
or U12579 (N_12579,N_11004,N_11962);
nand U12580 (N_12580,N_10566,N_11060);
xnor U12581 (N_12581,N_10804,N_10834);
and U12582 (N_12582,N_11936,N_11219);
nand U12583 (N_12583,N_10631,N_10652);
nand U12584 (N_12584,N_10954,N_11037);
nor U12585 (N_12585,N_10628,N_11834);
nor U12586 (N_12586,N_11874,N_11784);
nand U12587 (N_12587,N_10981,N_11606);
nand U12588 (N_12588,N_10680,N_10598);
nor U12589 (N_12589,N_11240,N_11163);
and U12590 (N_12590,N_10812,N_11821);
nor U12591 (N_12591,N_11647,N_10869);
or U12592 (N_12592,N_10873,N_11802);
nand U12593 (N_12593,N_11549,N_11571);
xor U12594 (N_12594,N_11857,N_10712);
nand U12595 (N_12595,N_10653,N_11134);
nor U12596 (N_12596,N_10635,N_11931);
or U12597 (N_12597,N_11972,N_11890);
nor U12598 (N_12598,N_10799,N_10535);
and U12599 (N_12599,N_11043,N_11524);
nor U12600 (N_12600,N_11699,N_11378);
and U12601 (N_12601,N_11797,N_11357);
or U12602 (N_12602,N_10866,N_10671);
xor U12603 (N_12603,N_11639,N_11081);
and U12604 (N_12604,N_11232,N_10835);
or U12605 (N_12605,N_11234,N_11836);
xnor U12606 (N_12606,N_10507,N_11015);
or U12607 (N_12607,N_10558,N_11897);
xor U12608 (N_12608,N_10607,N_11898);
and U12609 (N_12609,N_11202,N_11825);
and U12610 (N_12610,N_11494,N_11065);
xnor U12611 (N_12611,N_11477,N_11729);
xnor U12612 (N_12612,N_11716,N_10859);
nand U12613 (N_12613,N_10785,N_10974);
or U12614 (N_12614,N_10636,N_10934);
and U12615 (N_12615,N_10681,N_10662);
and U12616 (N_12616,N_10993,N_11912);
and U12617 (N_12617,N_11715,N_10585);
nor U12618 (N_12618,N_11786,N_10870);
or U12619 (N_12619,N_11554,N_11214);
nand U12620 (N_12620,N_11057,N_11570);
nor U12621 (N_12621,N_11559,N_11809);
or U12622 (N_12622,N_10659,N_10619);
and U12623 (N_12623,N_11411,N_10916);
nand U12624 (N_12624,N_11841,N_10633);
xnor U12625 (N_12625,N_10606,N_11657);
nand U12626 (N_12626,N_10877,N_11808);
or U12627 (N_12627,N_11865,N_11230);
nand U12628 (N_12628,N_11960,N_11342);
xnor U12629 (N_12629,N_11251,N_11038);
xor U12630 (N_12630,N_10854,N_11063);
and U12631 (N_12631,N_11158,N_11831);
and U12632 (N_12632,N_10809,N_10889);
xor U12633 (N_12633,N_10913,N_11833);
nor U12634 (N_12634,N_11848,N_11593);
nand U12635 (N_12635,N_11423,N_11457);
xnor U12636 (N_12636,N_11456,N_10801);
xnor U12637 (N_12637,N_11417,N_11678);
xor U12638 (N_12638,N_11121,N_11872);
nand U12639 (N_12639,N_11102,N_10691);
nor U12640 (N_12640,N_11767,N_11235);
nand U12641 (N_12641,N_11212,N_11165);
nand U12642 (N_12642,N_11264,N_11042);
nor U12643 (N_12643,N_11237,N_10830);
and U12644 (N_12644,N_11562,N_10509);
nor U12645 (N_12645,N_10657,N_11323);
and U12646 (N_12646,N_11547,N_11389);
and U12647 (N_12647,N_11948,N_10841);
nor U12648 (N_12648,N_11286,N_11260);
and U12649 (N_12649,N_11397,N_11576);
xor U12650 (N_12650,N_11363,N_11093);
nor U12651 (N_12651,N_11550,N_11878);
nor U12652 (N_12652,N_10847,N_11887);
and U12653 (N_12653,N_11517,N_10599);
xor U12654 (N_12654,N_11745,N_10698);
nor U12655 (N_12655,N_11430,N_11443);
nand U12656 (N_12656,N_11757,N_11470);
nor U12657 (N_12657,N_11396,N_10946);
xnor U12658 (N_12658,N_11064,N_10549);
xor U12659 (N_12659,N_11591,N_11979);
xor U12660 (N_12660,N_11131,N_10728);
nor U12661 (N_12661,N_10602,N_11380);
and U12662 (N_12662,N_11526,N_11721);
nor U12663 (N_12663,N_11680,N_11266);
xnor U12664 (N_12664,N_11752,N_11620);
nor U12665 (N_12665,N_11520,N_11200);
and U12666 (N_12666,N_10730,N_10703);
and U12667 (N_12667,N_11574,N_10560);
xnor U12668 (N_12668,N_10882,N_11024);
or U12669 (N_12669,N_11124,N_11697);
or U12670 (N_12670,N_11995,N_10501);
and U12671 (N_12671,N_10504,N_11183);
nand U12672 (N_12672,N_11217,N_10884);
nor U12673 (N_12673,N_10612,N_11436);
xnor U12674 (N_12674,N_11963,N_10900);
or U12675 (N_12675,N_10626,N_11769);
nor U12676 (N_12676,N_10575,N_11329);
or U12677 (N_12677,N_11041,N_11249);
and U12678 (N_12678,N_11137,N_11913);
or U12679 (N_12679,N_11655,N_10802);
or U12680 (N_12680,N_10823,N_11789);
xnor U12681 (N_12681,N_10684,N_11998);
and U12682 (N_12682,N_11295,N_11673);
xnor U12683 (N_12683,N_11335,N_11452);
nand U12684 (N_12684,N_11169,N_11287);
or U12685 (N_12685,N_10699,N_11001);
and U12686 (N_12686,N_11228,N_11701);
nor U12687 (N_12687,N_11932,N_10614);
nor U12688 (N_12688,N_10663,N_10721);
nor U12689 (N_12689,N_10926,N_10936);
or U12690 (N_12690,N_11672,N_10503);
nor U12691 (N_12691,N_10519,N_11581);
xor U12692 (N_12692,N_11994,N_11462);
and U12693 (N_12693,N_11166,N_10541);
and U12694 (N_12694,N_10759,N_11399);
xnor U12695 (N_12695,N_11771,N_11118);
and U12696 (N_12696,N_11271,N_10625);
nor U12697 (N_12697,N_10769,N_11514);
or U12698 (N_12698,N_11582,N_11476);
xnor U12699 (N_12699,N_11543,N_11407);
or U12700 (N_12700,N_11519,N_10556);
or U12701 (N_12701,N_11997,N_11741);
nand U12702 (N_12702,N_10723,N_11321);
nor U12703 (N_12703,N_10726,N_11408);
or U12704 (N_12704,N_11676,N_11218);
xor U12705 (N_12705,N_10629,N_10932);
or U12706 (N_12706,N_10702,N_11130);
nor U12707 (N_12707,N_11641,N_10583);
or U12708 (N_12708,N_11383,N_11014);
xor U12709 (N_12709,N_11182,N_10545);
nor U12710 (N_12710,N_11852,N_10725);
xor U12711 (N_12711,N_10500,N_11616);
nor U12712 (N_12712,N_10937,N_11077);
or U12713 (N_12713,N_11005,N_11501);
nor U12714 (N_12714,N_10980,N_11668);
nand U12715 (N_12715,N_11026,N_10706);
or U12716 (N_12716,N_10879,N_11599);
nand U12717 (N_12717,N_11904,N_10829);
xnor U12718 (N_12718,N_11965,N_10576);
nand U12719 (N_12719,N_11343,N_11667);
and U12720 (N_12720,N_11204,N_10747);
xnor U12721 (N_12721,N_11106,N_10586);
or U12722 (N_12722,N_11529,N_11609);
nor U12723 (N_12723,N_11682,N_11586);
and U12724 (N_12724,N_11175,N_10508);
xor U12725 (N_12725,N_10714,N_11440);
and U12726 (N_12726,N_11292,N_10685);
nor U12727 (N_12727,N_10880,N_10724);
nor U12728 (N_12728,N_11017,N_11114);
nor U12729 (N_12729,N_11761,N_10573);
xnor U12730 (N_12730,N_11089,N_11933);
or U12731 (N_12731,N_11420,N_11805);
nor U12732 (N_12732,N_11498,N_11340);
nor U12733 (N_12733,N_11598,N_11259);
nand U12734 (N_12734,N_11971,N_10548);
or U12735 (N_12735,N_11648,N_11534);
or U12736 (N_12736,N_10855,N_11050);
and U12737 (N_12737,N_11349,N_11123);
and U12738 (N_12738,N_11812,N_11773);
nand U12739 (N_12739,N_10861,N_11117);
and U12740 (N_12740,N_10773,N_10762);
nor U12741 (N_12741,N_10748,N_11937);
nand U12742 (N_12742,N_10518,N_11533);
xnor U12743 (N_12743,N_10661,N_11035);
or U12744 (N_12744,N_11927,N_10842);
nand U12745 (N_12745,N_11902,N_11987);
nand U12746 (N_12746,N_11261,N_11922);
or U12747 (N_12747,N_11849,N_11818);
xnor U12748 (N_12748,N_10966,N_11143);
nor U12749 (N_12749,N_10778,N_10523);
nand U12750 (N_12750,N_11672,N_11048);
or U12751 (N_12751,N_11305,N_11399);
xnor U12752 (N_12752,N_11279,N_11047);
xnor U12753 (N_12753,N_11331,N_10605);
xor U12754 (N_12754,N_11536,N_10510);
nand U12755 (N_12755,N_11164,N_10532);
and U12756 (N_12756,N_10685,N_11919);
nor U12757 (N_12757,N_10569,N_10547);
or U12758 (N_12758,N_11232,N_10525);
nand U12759 (N_12759,N_10678,N_10919);
or U12760 (N_12760,N_11672,N_11749);
or U12761 (N_12761,N_11648,N_11786);
nor U12762 (N_12762,N_10741,N_11746);
or U12763 (N_12763,N_11242,N_11256);
and U12764 (N_12764,N_11343,N_11214);
nand U12765 (N_12765,N_11188,N_11317);
or U12766 (N_12766,N_11132,N_10983);
nand U12767 (N_12767,N_11450,N_10572);
or U12768 (N_12768,N_10625,N_10511);
or U12769 (N_12769,N_11072,N_11050);
and U12770 (N_12770,N_10894,N_11527);
nor U12771 (N_12771,N_10879,N_11614);
and U12772 (N_12772,N_11826,N_11521);
nor U12773 (N_12773,N_11849,N_10758);
and U12774 (N_12774,N_11927,N_10744);
nand U12775 (N_12775,N_11285,N_11333);
nand U12776 (N_12776,N_10943,N_11861);
and U12777 (N_12777,N_11807,N_10756);
nand U12778 (N_12778,N_11698,N_10812);
or U12779 (N_12779,N_10860,N_11294);
nor U12780 (N_12780,N_11566,N_11856);
or U12781 (N_12781,N_11198,N_11433);
nor U12782 (N_12782,N_10948,N_11818);
nand U12783 (N_12783,N_11767,N_11029);
and U12784 (N_12784,N_10840,N_10576);
xnor U12785 (N_12785,N_10737,N_11355);
and U12786 (N_12786,N_11448,N_11758);
nor U12787 (N_12787,N_11738,N_10947);
and U12788 (N_12788,N_11040,N_10993);
nand U12789 (N_12789,N_10813,N_11184);
xnor U12790 (N_12790,N_10603,N_11571);
xor U12791 (N_12791,N_10653,N_10658);
and U12792 (N_12792,N_10624,N_10563);
nand U12793 (N_12793,N_11961,N_10767);
xnor U12794 (N_12794,N_10868,N_10928);
xor U12795 (N_12795,N_10676,N_11358);
nand U12796 (N_12796,N_11842,N_11249);
or U12797 (N_12797,N_10678,N_10689);
nor U12798 (N_12798,N_11779,N_11590);
xor U12799 (N_12799,N_11559,N_11242);
nand U12800 (N_12800,N_10873,N_11934);
or U12801 (N_12801,N_11137,N_10593);
or U12802 (N_12802,N_10997,N_11788);
nor U12803 (N_12803,N_11199,N_11349);
xnor U12804 (N_12804,N_11960,N_11303);
and U12805 (N_12805,N_11249,N_10707);
nor U12806 (N_12806,N_10699,N_11936);
or U12807 (N_12807,N_11382,N_11406);
xnor U12808 (N_12808,N_10619,N_11928);
xnor U12809 (N_12809,N_11266,N_11487);
nand U12810 (N_12810,N_11820,N_11940);
or U12811 (N_12811,N_11180,N_11489);
or U12812 (N_12812,N_11912,N_11724);
nand U12813 (N_12813,N_10515,N_11811);
and U12814 (N_12814,N_11255,N_10515);
xor U12815 (N_12815,N_10640,N_11732);
and U12816 (N_12816,N_10894,N_11414);
or U12817 (N_12817,N_10519,N_11325);
nor U12818 (N_12818,N_11810,N_10555);
and U12819 (N_12819,N_11497,N_10959);
and U12820 (N_12820,N_11643,N_10846);
and U12821 (N_12821,N_10930,N_10715);
xnor U12822 (N_12822,N_10915,N_10726);
and U12823 (N_12823,N_11814,N_10665);
or U12824 (N_12824,N_10572,N_11052);
nand U12825 (N_12825,N_11890,N_11243);
nand U12826 (N_12826,N_11128,N_11764);
or U12827 (N_12827,N_11373,N_10534);
xor U12828 (N_12828,N_11693,N_11894);
nand U12829 (N_12829,N_11090,N_10742);
xor U12830 (N_12830,N_11082,N_11592);
nand U12831 (N_12831,N_11370,N_10584);
xnor U12832 (N_12832,N_11319,N_11979);
and U12833 (N_12833,N_11907,N_10855);
and U12834 (N_12834,N_11320,N_10697);
and U12835 (N_12835,N_11659,N_11527);
nand U12836 (N_12836,N_11530,N_11609);
or U12837 (N_12837,N_11099,N_11334);
xnor U12838 (N_12838,N_11968,N_11784);
xor U12839 (N_12839,N_10680,N_10705);
and U12840 (N_12840,N_10575,N_10623);
xnor U12841 (N_12841,N_11908,N_11404);
nor U12842 (N_12842,N_10515,N_11095);
xor U12843 (N_12843,N_11518,N_11840);
and U12844 (N_12844,N_11340,N_11072);
or U12845 (N_12845,N_10673,N_10952);
and U12846 (N_12846,N_10522,N_11020);
nor U12847 (N_12847,N_10869,N_11898);
and U12848 (N_12848,N_11166,N_11943);
nand U12849 (N_12849,N_10829,N_10764);
nor U12850 (N_12850,N_10887,N_11630);
or U12851 (N_12851,N_10851,N_10605);
or U12852 (N_12852,N_11286,N_11712);
or U12853 (N_12853,N_11421,N_11316);
nand U12854 (N_12854,N_11920,N_11212);
nand U12855 (N_12855,N_11076,N_11849);
or U12856 (N_12856,N_11163,N_10703);
xor U12857 (N_12857,N_11228,N_11787);
or U12858 (N_12858,N_11412,N_10889);
nand U12859 (N_12859,N_10900,N_10500);
and U12860 (N_12860,N_11484,N_10769);
or U12861 (N_12861,N_10513,N_11963);
nor U12862 (N_12862,N_11377,N_10963);
xnor U12863 (N_12863,N_11239,N_11601);
nand U12864 (N_12864,N_10854,N_11181);
nor U12865 (N_12865,N_11467,N_11310);
nor U12866 (N_12866,N_10884,N_10975);
and U12867 (N_12867,N_11418,N_11294);
or U12868 (N_12868,N_11014,N_11841);
or U12869 (N_12869,N_10500,N_11800);
and U12870 (N_12870,N_11611,N_11350);
xnor U12871 (N_12871,N_11620,N_11985);
or U12872 (N_12872,N_11026,N_10594);
nor U12873 (N_12873,N_11511,N_11844);
nand U12874 (N_12874,N_10522,N_11194);
and U12875 (N_12875,N_11993,N_11508);
and U12876 (N_12876,N_10922,N_11359);
xor U12877 (N_12877,N_10690,N_11231);
xor U12878 (N_12878,N_11948,N_11336);
nor U12879 (N_12879,N_10792,N_11939);
xnor U12880 (N_12880,N_11911,N_11550);
xor U12881 (N_12881,N_11884,N_11174);
and U12882 (N_12882,N_11625,N_11399);
nor U12883 (N_12883,N_11762,N_11596);
nor U12884 (N_12884,N_11323,N_11268);
or U12885 (N_12885,N_11014,N_11999);
nor U12886 (N_12886,N_11228,N_11921);
nand U12887 (N_12887,N_10815,N_11957);
or U12888 (N_12888,N_10732,N_11632);
nand U12889 (N_12889,N_10964,N_11914);
nor U12890 (N_12890,N_10644,N_11678);
nand U12891 (N_12891,N_11373,N_11554);
and U12892 (N_12892,N_11279,N_11982);
xor U12893 (N_12893,N_11575,N_10653);
xnor U12894 (N_12894,N_10853,N_11859);
or U12895 (N_12895,N_10903,N_11352);
nand U12896 (N_12896,N_11075,N_11843);
nand U12897 (N_12897,N_10696,N_10915);
nor U12898 (N_12898,N_11528,N_11797);
nand U12899 (N_12899,N_11712,N_11190);
and U12900 (N_12900,N_10929,N_11769);
nand U12901 (N_12901,N_11077,N_11837);
and U12902 (N_12902,N_11655,N_11222);
xnor U12903 (N_12903,N_10620,N_11974);
and U12904 (N_12904,N_11063,N_11657);
nand U12905 (N_12905,N_10689,N_11330);
and U12906 (N_12906,N_11084,N_11529);
and U12907 (N_12907,N_11447,N_11266);
nor U12908 (N_12908,N_11760,N_11658);
nor U12909 (N_12909,N_11115,N_10935);
nand U12910 (N_12910,N_11759,N_11841);
or U12911 (N_12911,N_11925,N_11908);
nand U12912 (N_12912,N_11220,N_11516);
xnor U12913 (N_12913,N_10815,N_10608);
and U12914 (N_12914,N_11924,N_10547);
xnor U12915 (N_12915,N_10930,N_11888);
xnor U12916 (N_12916,N_11795,N_11684);
and U12917 (N_12917,N_11087,N_10780);
and U12918 (N_12918,N_10792,N_10590);
xor U12919 (N_12919,N_11158,N_11582);
xnor U12920 (N_12920,N_10924,N_10684);
or U12921 (N_12921,N_11802,N_11528);
nor U12922 (N_12922,N_11829,N_11551);
or U12923 (N_12923,N_11870,N_11678);
and U12924 (N_12924,N_10743,N_11935);
nand U12925 (N_12925,N_10804,N_11891);
nor U12926 (N_12926,N_10631,N_11038);
nand U12927 (N_12927,N_11013,N_11825);
xnor U12928 (N_12928,N_11549,N_11664);
xor U12929 (N_12929,N_11585,N_11728);
or U12930 (N_12930,N_11815,N_11620);
nand U12931 (N_12931,N_11694,N_10943);
and U12932 (N_12932,N_11683,N_11971);
nor U12933 (N_12933,N_11430,N_11886);
xnor U12934 (N_12934,N_11038,N_10620);
nand U12935 (N_12935,N_10586,N_11754);
and U12936 (N_12936,N_11878,N_10909);
nor U12937 (N_12937,N_11545,N_11092);
nor U12938 (N_12938,N_11655,N_11153);
xnor U12939 (N_12939,N_11460,N_10987);
nand U12940 (N_12940,N_11395,N_11461);
xor U12941 (N_12941,N_10853,N_11413);
nor U12942 (N_12942,N_11047,N_11341);
and U12943 (N_12943,N_11430,N_10545);
or U12944 (N_12944,N_11748,N_10879);
nor U12945 (N_12945,N_10885,N_11585);
or U12946 (N_12946,N_11338,N_11607);
and U12947 (N_12947,N_11812,N_11259);
and U12948 (N_12948,N_11269,N_10828);
nor U12949 (N_12949,N_11438,N_10914);
and U12950 (N_12950,N_10636,N_11148);
nand U12951 (N_12951,N_11931,N_11703);
nor U12952 (N_12952,N_11869,N_11136);
or U12953 (N_12953,N_11937,N_11808);
nand U12954 (N_12954,N_11176,N_11386);
nand U12955 (N_12955,N_11027,N_11396);
and U12956 (N_12956,N_11225,N_10712);
nand U12957 (N_12957,N_11037,N_11852);
or U12958 (N_12958,N_10527,N_11180);
and U12959 (N_12959,N_10790,N_10918);
nor U12960 (N_12960,N_11339,N_11504);
nand U12961 (N_12961,N_11017,N_11078);
nor U12962 (N_12962,N_10898,N_10687);
nand U12963 (N_12963,N_10747,N_10678);
or U12964 (N_12964,N_11390,N_11883);
nor U12965 (N_12965,N_11573,N_11392);
nor U12966 (N_12966,N_11356,N_11838);
or U12967 (N_12967,N_10516,N_10548);
xnor U12968 (N_12968,N_10605,N_11326);
xor U12969 (N_12969,N_11897,N_11224);
or U12970 (N_12970,N_11799,N_11597);
xnor U12971 (N_12971,N_10756,N_10936);
nor U12972 (N_12972,N_10805,N_11793);
nand U12973 (N_12973,N_10728,N_11651);
nor U12974 (N_12974,N_11233,N_11729);
or U12975 (N_12975,N_10627,N_11890);
or U12976 (N_12976,N_11225,N_11129);
xnor U12977 (N_12977,N_10623,N_11790);
or U12978 (N_12978,N_10914,N_10579);
nand U12979 (N_12979,N_11411,N_11847);
or U12980 (N_12980,N_10604,N_11535);
nand U12981 (N_12981,N_11843,N_10902);
or U12982 (N_12982,N_11784,N_11372);
or U12983 (N_12983,N_10512,N_10573);
nor U12984 (N_12984,N_11740,N_11033);
and U12985 (N_12985,N_10886,N_11115);
nand U12986 (N_12986,N_11577,N_10500);
or U12987 (N_12987,N_11009,N_10972);
xnor U12988 (N_12988,N_10708,N_10794);
nand U12989 (N_12989,N_11914,N_11720);
nor U12990 (N_12990,N_11199,N_11335);
nor U12991 (N_12991,N_11509,N_11167);
xnor U12992 (N_12992,N_10576,N_11917);
xor U12993 (N_12993,N_11366,N_11018);
nand U12994 (N_12994,N_10674,N_10513);
nor U12995 (N_12995,N_11842,N_11609);
nand U12996 (N_12996,N_11972,N_11240);
and U12997 (N_12997,N_11569,N_11038);
nand U12998 (N_12998,N_10714,N_11426);
or U12999 (N_12999,N_10720,N_11829);
or U13000 (N_13000,N_11820,N_11157);
or U13001 (N_13001,N_10929,N_11164);
xnor U13002 (N_13002,N_10692,N_11558);
nor U13003 (N_13003,N_10747,N_11289);
nor U13004 (N_13004,N_11177,N_11996);
or U13005 (N_13005,N_11627,N_11645);
or U13006 (N_13006,N_11948,N_10574);
nand U13007 (N_13007,N_11781,N_11024);
xor U13008 (N_13008,N_11312,N_11479);
and U13009 (N_13009,N_11633,N_11439);
nand U13010 (N_13010,N_11369,N_11041);
nor U13011 (N_13011,N_11098,N_11345);
or U13012 (N_13012,N_11542,N_11339);
and U13013 (N_13013,N_11693,N_10648);
nand U13014 (N_13014,N_11674,N_10654);
and U13015 (N_13015,N_11523,N_10723);
and U13016 (N_13016,N_10886,N_11041);
and U13017 (N_13017,N_11705,N_11499);
nor U13018 (N_13018,N_10986,N_10660);
and U13019 (N_13019,N_11816,N_10613);
and U13020 (N_13020,N_10661,N_10685);
or U13021 (N_13021,N_10816,N_10890);
or U13022 (N_13022,N_11444,N_10998);
or U13023 (N_13023,N_10742,N_11667);
and U13024 (N_13024,N_10743,N_11546);
nand U13025 (N_13025,N_11184,N_10594);
xnor U13026 (N_13026,N_11092,N_11337);
nand U13027 (N_13027,N_11685,N_11999);
or U13028 (N_13028,N_11270,N_11237);
or U13029 (N_13029,N_10883,N_11313);
or U13030 (N_13030,N_11990,N_11195);
and U13031 (N_13031,N_11533,N_11928);
nor U13032 (N_13032,N_11665,N_11502);
nor U13033 (N_13033,N_10851,N_10830);
or U13034 (N_13034,N_10578,N_11725);
or U13035 (N_13035,N_10629,N_10872);
or U13036 (N_13036,N_11380,N_11112);
nand U13037 (N_13037,N_11987,N_11566);
or U13038 (N_13038,N_11483,N_11579);
xnor U13039 (N_13039,N_11317,N_10940);
xnor U13040 (N_13040,N_11621,N_10708);
or U13041 (N_13041,N_11582,N_10966);
nand U13042 (N_13042,N_11248,N_11928);
nand U13043 (N_13043,N_11435,N_11897);
xnor U13044 (N_13044,N_10987,N_10738);
or U13045 (N_13045,N_10678,N_11236);
nor U13046 (N_13046,N_11186,N_11237);
xnor U13047 (N_13047,N_10884,N_11016);
or U13048 (N_13048,N_10825,N_11871);
or U13049 (N_13049,N_10998,N_11320);
xnor U13050 (N_13050,N_10868,N_11216);
and U13051 (N_13051,N_11365,N_10850);
nand U13052 (N_13052,N_10743,N_11285);
nand U13053 (N_13053,N_11756,N_11061);
nor U13054 (N_13054,N_11812,N_10909);
and U13055 (N_13055,N_11015,N_11001);
nand U13056 (N_13056,N_11853,N_10800);
or U13057 (N_13057,N_11984,N_10557);
xor U13058 (N_13058,N_11645,N_11084);
xnor U13059 (N_13059,N_11323,N_11491);
xnor U13060 (N_13060,N_11134,N_10842);
or U13061 (N_13061,N_10715,N_11008);
or U13062 (N_13062,N_11110,N_11589);
and U13063 (N_13063,N_11051,N_10886);
nand U13064 (N_13064,N_10806,N_11489);
xor U13065 (N_13065,N_11520,N_11836);
or U13066 (N_13066,N_11580,N_10719);
nand U13067 (N_13067,N_11000,N_10967);
xor U13068 (N_13068,N_10809,N_10850);
nand U13069 (N_13069,N_10625,N_11172);
or U13070 (N_13070,N_11799,N_11036);
xnor U13071 (N_13071,N_11329,N_11912);
nand U13072 (N_13072,N_11649,N_11830);
nor U13073 (N_13073,N_10990,N_11234);
and U13074 (N_13074,N_11350,N_11723);
xor U13075 (N_13075,N_10964,N_11832);
nor U13076 (N_13076,N_10667,N_11947);
nand U13077 (N_13077,N_11230,N_11156);
nand U13078 (N_13078,N_10731,N_11101);
nand U13079 (N_13079,N_10661,N_11560);
and U13080 (N_13080,N_11329,N_11895);
or U13081 (N_13081,N_10959,N_11192);
and U13082 (N_13082,N_11926,N_11797);
nor U13083 (N_13083,N_10653,N_11613);
nor U13084 (N_13084,N_11868,N_11483);
or U13085 (N_13085,N_11085,N_11168);
nor U13086 (N_13086,N_11434,N_10842);
xor U13087 (N_13087,N_11701,N_11556);
nor U13088 (N_13088,N_11765,N_10911);
xor U13089 (N_13089,N_10706,N_11117);
xor U13090 (N_13090,N_10949,N_11231);
xor U13091 (N_13091,N_10890,N_11345);
nand U13092 (N_13092,N_11060,N_11188);
or U13093 (N_13093,N_10937,N_11750);
xnor U13094 (N_13094,N_11047,N_10803);
xor U13095 (N_13095,N_11481,N_11142);
nand U13096 (N_13096,N_11365,N_10540);
nor U13097 (N_13097,N_11513,N_11782);
or U13098 (N_13098,N_10881,N_11264);
or U13099 (N_13099,N_11357,N_10615);
nand U13100 (N_13100,N_10692,N_11517);
xnor U13101 (N_13101,N_10920,N_10725);
or U13102 (N_13102,N_11718,N_10567);
or U13103 (N_13103,N_11455,N_11496);
nand U13104 (N_13104,N_11991,N_10543);
nand U13105 (N_13105,N_11968,N_11613);
or U13106 (N_13106,N_11953,N_11011);
xnor U13107 (N_13107,N_10864,N_10597);
xor U13108 (N_13108,N_11015,N_11351);
xnor U13109 (N_13109,N_11326,N_10732);
nor U13110 (N_13110,N_11629,N_11607);
or U13111 (N_13111,N_10579,N_11047);
nand U13112 (N_13112,N_11707,N_11527);
and U13113 (N_13113,N_11642,N_11641);
nor U13114 (N_13114,N_10807,N_11386);
or U13115 (N_13115,N_10613,N_11974);
and U13116 (N_13116,N_11007,N_11419);
xnor U13117 (N_13117,N_11801,N_11317);
and U13118 (N_13118,N_11696,N_11248);
nor U13119 (N_13119,N_11896,N_11238);
nor U13120 (N_13120,N_11718,N_11904);
or U13121 (N_13121,N_10928,N_10511);
nor U13122 (N_13122,N_10923,N_10855);
nand U13123 (N_13123,N_11761,N_11460);
and U13124 (N_13124,N_11261,N_11894);
nor U13125 (N_13125,N_10548,N_11346);
nand U13126 (N_13126,N_11740,N_11035);
nand U13127 (N_13127,N_11506,N_11832);
nor U13128 (N_13128,N_11626,N_10590);
nor U13129 (N_13129,N_11372,N_11031);
nor U13130 (N_13130,N_11269,N_10890);
and U13131 (N_13131,N_11225,N_10862);
and U13132 (N_13132,N_11418,N_10984);
nor U13133 (N_13133,N_10510,N_10747);
nor U13134 (N_13134,N_11534,N_10503);
and U13135 (N_13135,N_11015,N_11520);
or U13136 (N_13136,N_10505,N_11751);
nor U13137 (N_13137,N_11836,N_11145);
xor U13138 (N_13138,N_11771,N_11024);
and U13139 (N_13139,N_11188,N_11636);
and U13140 (N_13140,N_11607,N_11344);
or U13141 (N_13141,N_11570,N_10546);
nor U13142 (N_13142,N_10570,N_11525);
nor U13143 (N_13143,N_11459,N_11347);
xnor U13144 (N_13144,N_10890,N_10737);
nor U13145 (N_13145,N_11610,N_10829);
nor U13146 (N_13146,N_11796,N_10610);
nand U13147 (N_13147,N_11800,N_11989);
and U13148 (N_13148,N_11644,N_11858);
xnor U13149 (N_13149,N_10669,N_10881);
and U13150 (N_13150,N_11621,N_10603);
and U13151 (N_13151,N_11642,N_11571);
and U13152 (N_13152,N_11137,N_11268);
or U13153 (N_13153,N_10846,N_11709);
xnor U13154 (N_13154,N_11175,N_10864);
and U13155 (N_13155,N_11716,N_11310);
and U13156 (N_13156,N_10768,N_10578);
xnor U13157 (N_13157,N_11310,N_10876);
nand U13158 (N_13158,N_10842,N_10659);
xor U13159 (N_13159,N_11816,N_10522);
and U13160 (N_13160,N_10872,N_10829);
nand U13161 (N_13161,N_11660,N_11569);
or U13162 (N_13162,N_10982,N_10980);
or U13163 (N_13163,N_11573,N_10573);
nor U13164 (N_13164,N_11197,N_11412);
xor U13165 (N_13165,N_11270,N_11466);
and U13166 (N_13166,N_10832,N_11283);
nor U13167 (N_13167,N_11951,N_11321);
or U13168 (N_13168,N_11947,N_11807);
nand U13169 (N_13169,N_11793,N_11795);
and U13170 (N_13170,N_11149,N_11850);
or U13171 (N_13171,N_10600,N_11050);
nand U13172 (N_13172,N_10679,N_11922);
xnor U13173 (N_13173,N_11693,N_11602);
or U13174 (N_13174,N_11651,N_11792);
xnor U13175 (N_13175,N_11556,N_11561);
nor U13176 (N_13176,N_10750,N_11542);
and U13177 (N_13177,N_11464,N_11878);
xor U13178 (N_13178,N_10769,N_10601);
xor U13179 (N_13179,N_11094,N_11623);
nor U13180 (N_13180,N_10517,N_11610);
nor U13181 (N_13181,N_10505,N_10545);
nor U13182 (N_13182,N_11811,N_10911);
nand U13183 (N_13183,N_11973,N_11019);
nand U13184 (N_13184,N_10917,N_11388);
nand U13185 (N_13185,N_11102,N_10704);
and U13186 (N_13186,N_11764,N_10837);
and U13187 (N_13187,N_11114,N_10957);
and U13188 (N_13188,N_10564,N_11899);
or U13189 (N_13189,N_11484,N_11863);
or U13190 (N_13190,N_11453,N_11177);
nor U13191 (N_13191,N_11293,N_11389);
or U13192 (N_13192,N_11819,N_11477);
xor U13193 (N_13193,N_11934,N_10882);
nor U13194 (N_13194,N_11360,N_10546);
nor U13195 (N_13195,N_10715,N_11687);
nand U13196 (N_13196,N_10775,N_10715);
or U13197 (N_13197,N_10522,N_11015);
nor U13198 (N_13198,N_11782,N_11328);
nor U13199 (N_13199,N_11140,N_11273);
nand U13200 (N_13200,N_10703,N_11362);
xor U13201 (N_13201,N_11640,N_10632);
xor U13202 (N_13202,N_11327,N_10782);
xor U13203 (N_13203,N_10757,N_11539);
xor U13204 (N_13204,N_11882,N_11873);
or U13205 (N_13205,N_10866,N_11925);
nand U13206 (N_13206,N_10933,N_11127);
and U13207 (N_13207,N_11087,N_11067);
xor U13208 (N_13208,N_11098,N_11685);
xor U13209 (N_13209,N_10633,N_11363);
nand U13210 (N_13210,N_10962,N_11490);
nand U13211 (N_13211,N_11856,N_11647);
nand U13212 (N_13212,N_11201,N_11152);
nand U13213 (N_13213,N_10620,N_10614);
xor U13214 (N_13214,N_10509,N_10954);
or U13215 (N_13215,N_11596,N_11122);
and U13216 (N_13216,N_11715,N_11644);
and U13217 (N_13217,N_11134,N_10525);
nand U13218 (N_13218,N_10824,N_11567);
or U13219 (N_13219,N_10765,N_11887);
or U13220 (N_13220,N_11649,N_11563);
nor U13221 (N_13221,N_11061,N_11986);
nand U13222 (N_13222,N_11633,N_11173);
nand U13223 (N_13223,N_10888,N_11787);
xor U13224 (N_13224,N_10588,N_11388);
nor U13225 (N_13225,N_11118,N_11289);
or U13226 (N_13226,N_11911,N_11969);
or U13227 (N_13227,N_11302,N_10823);
nand U13228 (N_13228,N_10768,N_11923);
xor U13229 (N_13229,N_11819,N_10765);
xor U13230 (N_13230,N_10685,N_10674);
and U13231 (N_13231,N_11784,N_11457);
xor U13232 (N_13232,N_11814,N_11005);
nand U13233 (N_13233,N_11688,N_11439);
xor U13234 (N_13234,N_11423,N_11554);
nand U13235 (N_13235,N_11752,N_10564);
and U13236 (N_13236,N_10671,N_10978);
nor U13237 (N_13237,N_11663,N_11518);
nor U13238 (N_13238,N_11257,N_11772);
or U13239 (N_13239,N_10542,N_11207);
and U13240 (N_13240,N_11950,N_10693);
or U13241 (N_13241,N_11135,N_11884);
and U13242 (N_13242,N_11684,N_11273);
or U13243 (N_13243,N_11115,N_11639);
nor U13244 (N_13244,N_10784,N_11338);
or U13245 (N_13245,N_11718,N_11857);
or U13246 (N_13246,N_11246,N_10632);
nand U13247 (N_13247,N_11815,N_11256);
nor U13248 (N_13248,N_10728,N_11895);
nand U13249 (N_13249,N_10843,N_11361);
nand U13250 (N_13250,N_11182,N_10908);
nand U13251 (N_13251,N_11606,N_10954);
nor U13252 (N_13252,N_10520,N_11541);
nand U13253 (N_13253,N_11084,N_10617);
and U13254 (N_13254,N_11205,N_10911);
and U13255 (N_13255,N_11217,N_11696);
nand U13256 (N_13256,N_11720,N_10711);
nor U13257 (N_13257,N_10783,N_11398);
nand U13258 (N_13258,N_10770,N_11031);
or U13259 (N_13259,N_10710,N_11093);
nand U13260 (N_13260,N_11468,N_11286);
xor U13261 (N_13261,N_10951,N_11269);
xor U13262 (N_13262,N_11361,N_10891);
or U13263 (N_13263,N_11924,N_11840);
xnor U13264 (N_13264,N_10984,N_11767);
or U13265 (N_13265,N_11477,N_11356);
and U13266 (N_13266,N_11384,N_11897);
nand U13267 (N_13267,N_11871,N_11251);
nor U13268 (N_13268,N_11589,N_10624);
and U13269 (N_13269,N_11804,N_11584);
nor U13270 (N_13270,N_11890,N_10659);
and U13271 (N_13271,N_10922,N_11698);
nor U13272 (N_13272,N_11254,N_11036);
xor U13273 (N_13273,N_11685,N_10954);
xnor U13274 (N_13274,N_11282,N_11371);
nor U13275 (N_13275,N_10995,N_11435);
nor U13276 (N_13276,N_11050,N_11650);
xnor U13277 (N_13277,N_10720,N_11370);
and U13278 (N_13278,N_11116,N_10906);
or U13279 (N_13279,N_11340,N_10684);
nand U13280 (N_13280,N_11649,N_10683);
xor U13281 (N_13281,N_10830,N_10796);
xor U13282 (N_13282,N_11299,N_11098);
nor U13283 (N_13283,N_11417,N_10708);
nand U13284 (N_13284,N_11896,N_10568);
and U13285 (N_13285,N_11606,N_11274);
xnor U13286 (N_13286,N_11838,N_11403);
nor U13287 (N_13287,N_11161,N_11582);
nor U13288 (N_13288,N_11296,N_11613);
xor U13289 (N_13289,N_10869,N_11137);
or U13290 (N_13290,N_10848,N_11401);
xor U13291 (N_13291,N_11759,N_10898);
and U13292 (N_13292,N_10730,N_10971);
xor U13293 (N_13293,N_11648,N_11220);
xor U13294 (N_13294,N_10944,N_11697);
nand U13295 (N_13295,N_10870,N_11766);
and U13296 (N_13296,N_11231,N_11230);
nor U13297 (N_13297,N_10586,N_10571);
and U13298 (N_13298,N_11531,N_10693);
xor U13299 (N_13299,N_10887,N_10993);
nand U13300 (N_13300,N_10736,N_11413);
or U13301 (N_13301,N_11932,N_11059);
xor U13302 (N_13302,N_11443,N_11261);
or U13303 (N_13303,N_11196,N_10717);
and U13304 (N_13304,N_11608,N_11165);
nand U13305 (N_13305,N_10963,N_11906);
and U13306 (N_13306,N_10564,N_10537);
and U13307 (N_13307,N_10984,N_10838);
or U13308 (N_13308,N_10590,N_11416);
xor U13309 (N_13309,N_11901,N_10583);
xor U13310 (N_13310,N_11659,N_11606);
nand U13311 (N_13311,N_11436,N_10704);
or U13312 (N_13312,N_10952,N_10605);
nand U13313 (N_13313,N_11826,N_11370);
xnor U13314 (N_13314,N_10777,N_10886);
xnor U13315 (N_13315,N_11949,N_10679);
xor U13316 (N_13316,N_11611,N_11364);
xor U13317 (N_13317,N_11358,N_11719);
or U13318 (N_13318,N_11128,N_11436);
and U13319 (N_13319,N_11034,N_11984);
or U13320 (N_13320,N_11642,N_11975);
nor U13321 (N_13321,N_11099,N_11701);
nand U13322 (N_13322,N_11784,N_11433);
and U13323 (N_13323,N_10513,N_10541);
nand U13324 (N_13324,N_11124,N_10718);
nor U13325 (N_13325,N_11150,N_11833);
or U13326 (N_13326,N_11872,N_10665);
nand U13327 (N_13327,N_11822,N_11182);
or U13328 (N_13328,N_10583,N_11016);
nand U13329 (N_13329,N_11699,N_11350);
xnor U13330 (N_13330,N_11156,N_10705);
xnor U13331 (N_13331,N_10771,N_11512);
or U13332 (N_13332,N_10952,N_11240);
nor U13333 (N_13333,N_10761,N_11728);
nor U13334 (N_13334,N_11777,N_10796);
or U13335 (N_13335,N_10933,N_10849);
and U13336 (N_13336,N_10708,N_11852);
xnor U13337 (N_13337,N_11462,N_11288);
or U13338 (N_13338,N_10889,N_11111);
nor U13339 (N_13339,N_10591,N_10873);
and U13340 (N_13340,N_10925,N_11425);
nor U13341 (N_13341,N_10936,N_11813);
or U13342 (N_13342,N_11611,N_11812);
and U13343 (N_13343,N_10660,N_10517);
xnor U13344 (N_13344,N_10620,N_11520);
and U13345 (N_13345,N_10704,N_11953);
or U13346 (N_13346,N_11295,N_10518);
nand U13347 (N_13347,N_10512,N_11273);
and U13348 (N_13348,N_11530,N_11671);
xnor U13349 (N_13349,N_10848,N_10998);
nand U13350 (N_13350,N_10730,N_11367);
and U13351 (N_13351,N_11946,N_11596);
and U13352 (N_13352,N_10948,N_11679);
or U13353 (N_13353,N_10652,N_11275);
xor U13354 (N_13354,N_11117,N_10996);
nor U13355 (N_13355,N_10974,N_11587);
or U13356 (N_13356,N_11217,N_10931);
xnor U13357 (N_13357,N_11062,N_11609);
and U13358 (N_13358,N_11547,N_11798);
xnor U13359 (N_13359,N_11433,N_10805);
xor U13360 (N_13360,N_11520,N_10826);
xnor U13361 (N_13361,N_11750,N_10818);
nand U13362 (N_13362,N_11829,N_11987);
nand U13363 (N_13363,N_10715,N_11004);
nor U13364 (N_13364,N_10527,N_10817);
nand U13365 (N_13365,N_11085,N_11880);
and U13366 (N_13366,N_11204,N_10699);
and U13367 (N_13367,N_11199,N_10668);
nand U13368 (N_13368,N_11170,N_11943);
xnor U13369 (N_13369,N_10851,N_11244);
nor U13370 (N_13370,N_10772,N_11470);
nand U13371 (N_13371,N_10717,N_11317);
nor U13372 (N_13372,N_10569,N_11966);
nand U13373 (N_13373,N_11257,N_10544);
or U13374 (N_13374,N_10837,N_11120);
or U13375 (N_13375,N_11773,N_10805);
and U13376 (N_13376,N_11856,N_11447);
xnor U13377 (N_13377,N_11625,N_11517);
or U13378 (N_13378,N_11477,N_11091);
and U13379 (N_13379,N_10713,N_11957);
nand U13380 (N_13380,N_11726,N_10557);
nor U13381 (N_13381,N_11907,N_11176);
nand U13382 (N_13382,N_11590,N_11309);
xor U13383 (N_13383,N_10936,N_11558);
and U13384 (N_13384,N_11376,N_11281);
xor U13385 (N_13385,N_11002,N_11154);
and U13386 (N_13386,N_11523,N_10779);
nand U13387 (N_13387,N_10634,N_11845);
and U13388 (N_13388,N_11059,N_11179);
and U13389 (N_13389,N_11019,N_11621);
nand U13390 (N_13390,N_10833,N_11471);
or U13391 (N_13391,N_10853,N_10565);
nor U13392 (N_13392,N_10581,N_11857);
nor U13393 (N_13393,N_11552,N_11361);
and U13394 (N_13394,N_11252,N_11724);
and U13395 (N_13395,N_11810,N_10559);
xnor U13396 (N_13396,N_10802,N_10670);
nand U13397 (N_13397,N_10830,N_11923);
nor U13398 (N_13398,N_11490,N_11348);
nand U13399 (N_13399,N_11982,N_10849);
nor U13400 (N_13400,N_11286,N_11070);
nand U13401 (N_13401,N_11161,N_11362);
and U13402 (N_13402,N_10976,N_11601);
or U13403 (N_13403,N_11528,N_10688);
nand U13404 (N_13404,N_11816,N_11446);
nand U13405 (N_13405,N_10702,N_11299);
or U13406 (N_13406,N_11373,N_11099);
xnor U13407 (N_13407,N_11781,N_11428);
xor U13408 (N_13408,N_11443,N_10582);
xor U13409 (N_13409,N_11975,N_11363);
xnor U13410 (N_13410,N_10741,N_11534);
nor U13411 (N_13411,N_11991,N_10684);
nor U13412 (N_13412,N_11530,N_11880);
xor U13413 (N_13413,N_11175,N_11586);
or U13414 (N_13414,N_10788,N_11967);
and U13415 (N_13415,N_11363,N_11819);
and U13416 (N_13416,N_10708,N_11605);
nand U13417 (N_13417,N_11470,N_10895);
xor U13418 (N_13418,N_11177,N_10561);
nor U13419 (N_13419,N_11497,N_11468);
and U13420 (N_13420,N_11523,N_11888);
nand U13421 (N_13421,N_11519,N_10573);
nor U13422 (N_13422,N_11080,N_11432);
nand U13423 (N_13423,N_11614,N_11053);
nor U13424 (N_13424,N_11815,N_10821);
nor U13425 (N_13425,N_11293,N_10851);
xor U13426 (N_13426,N_11146,N_11401);
nor U13427 (N_13427,N_11596,N_11444);
and U13428 (N_13428,N_10728,N_11877);
and U13429 (N_13429,N_11506,N_11472);
nor U13430 (N_13430,N_11728,N_11383);
nor U13431 (N_13431,N_10802,N_10676);
xnor U13432 (N_13432,N_11702,N_11829);
xor U13433 (N_13433,N_11436,N_11122);
xnor U13434 (N_13434,N_11180,N_11815);
nor U13435 (N_13435,N_11343,N_10826);
and U13436 (N_13436,N_11705,N_11202);
or U13437 (N_13437,N_10979,N_11523);
nor U13438 (N_13438,N_10502,N_11765);
or U13439 (N_13439,N_10711,N_10773);
or U13440 (N_13440,N_11057,N_10947);
nor U13441 (N_13441,N_11115,N_10888);
nand U13442 (N_13442,N_10869,N_11922);
or U13443 (N_13443,N_10910,N_11464);
and U13444 (N_13444,N_11125,N_10653);
and U13445 (N_13445,N_10776,N_11056);
nor U13446 (N_13446,N_11311,N_10949);
xnor U13447 (N_13447,N_11995,N_11712);
nand U13448 (N_13448,N_11028,N_10540);
xor U13449 (N_13449,N_11326,N_10536);
nor U13450 (N_13450,N_11621,N_10584);
and U13451 (N_13451,N_11368,N_10701);
nand U13452 (N_13452,N_11648,N_11982);
nor U13453 (N_13453,N_11992,N_11673);
nand U13454 (N_13454,N_11769,N_11713);
xor U13455 (N_13455,N_11366,N_11219);
and U13456 (N_13456,N_11976,N_11469);
nor U13457 (N_13457,N_11950,N_10723);
or U13458 (N_13458,N_11632,N_11953);
nor U13459 (N_13459,N_11512,N_11129);
nor U13460 (N_13460,N_10858,N_10899);
nand U13461 (N_13461,N_11671,N_10586);
or U13462 (N_13462,N_10729,N_11848);
nor U13463 (N_13463,N_11860,N_11375);
nor U13464 (N_13464,N_10885,N_10818);
and U13465 (N_13465,N_11395,N_11124);
xor U13466 (N_13466,N_11828,N_11832);
and U13467 (N_13467,N_10687,N_11695);
and U13468 (N_13468,N_11584,N_11852);
xor U13469 (N_13469,N_11006,N_11458);
and U13470 (N_13470,N_10781,N_11244);
and U13471 (N_13471,N_11745,N_11476);
nand U13472 (N_13472,N_11094,N_11203);
and U13473 (N_13473,N_11336,N_11701);
or U13474 (N_13474,N_10624,N_10616);
and U13475 (N_13475,N_11847,N_11542);
or U13476 (N_13476,N_11881,N_11083);
or U13477 (N_13477,N_11425,N_10769);
nand U13478 (N_13478,N_11355,N_11738);
xnor U13479 (N_13479,N_10579,N_11900);
nor U13480 (N_13480,N_11300,N_11607);
nand U13481 (N_13481,N_11593,N_11827);
and U13482 (N_13482,N_11910,N_10529);
nand U13483 (N_13483,N_10679,N_11424);
and U13484 (N_13484,N_10591,N_11859);
nand U13485 (N_13485,N_11583,N_10550);
and U13486 (N_13486,N_11135,N_11043);
and U13487 (N_13487,N_11696,N_11573);
and U13488 (N_13488,N_11844,N_10977);
nor U13489 (N_13489,N_10718,N_10817);
or U13490 (N_13490,N_10998,N_11599);
nor U13491 (N_13491,N_10931,N_11067);
nor U13492 (N_13492,N_10942,N_10965);
nor U13493 (N_13493,N_11907,N_10832);
nor U13494 (N_13494,N_11422,N_10668);
nand U13495 (N_13495,N_11102,N_11650);
and U13496 (N_13496,N_10687,N_10507);
nor U13497 (N_13497,N_11823,N_11224);
and U13498 (N_13498,N_11241,N_11987);
xnor U13499 (N_13499,N_11580,N_11325);
nor U13500 (N_13500,N_12976,N_13471);
nand U13501 (N_13501,N_13236,N_12619);
xnor U13502 (N_13502,N_12109,N_13126);
nor U13503 (N_13503,N_12610,N_13488);
nor U13504 (N_13504,N_13159,N_12186);
nand U13505 (N_13505,N_13454,N_13343);
and U13506 (N_13506,N_13341,N_13180);
nand U13507 (N_13507,N_13167,N_12150);
xor U13508 (N_13508,N_13214,N_12641);
and U13509 (N_13509,N_12541,N_12993);
xnor U13510 (N_13510,N_13456,N_12810);
and U13511 (N_13511,N_12622,N_12921);
and U13512 (N_13512,N_12489,N_13018);
xnor U13513 (N_13513,N_12323,N_12973);
nor U13514 (N_13514,N_12889,N_12819);
nor U13515 (N_13515,N_12594,N_12532);
or U13516 (N_13516,N_12146,N_12542);
or U13517 (N_13517,N_13345,N_13349);
nand U13518 (N_13518,N_12788,N_12488);
nand U13519 (N_13519,N_13242,N_12683);
and U13520 (N_13520,N_12691,N_13333);
xnor U13521 (N_13521,N_13472,N_13469);
xor U13522 (N_13522,N_12706,N_13417);
and U13523 (N_13523,N_12848,N_12593);
xor U13524 (N_13524,N_12236,N_12509);
nand U13525 (N_13525,N_13478,N_13119);
or U13526 (N_13526,N_12590,N_12799);
or U13527 (N_13527,N_12733,N_12855);
nand U13528 (N_13528,N_12475,N_13385);
or U13529 (N_13529,N_12714,N_13161);
or U13530 (N_13530,N_12721,N_12241);
nor U13531 (N_13531,N_12115,N_12493);
nand U13532 (N_13532,N_12661,N_13303);
and U13533 (N_13533,N_12046,N_12937);
or U13534 (N_13534,N_12245,N_12010);
and U13535 (N_13535,N_13389,N_12329);
nor U13536 (N_13536,N_12379,N_12098);
nand U13537 (N_13537,N_12203,N_12292);
or U13538 (N_13538,N_12125,N_12777);
xnor U13539 (N_13539,N_13444,N_12082);
xnor U13540 (N_13540,N_13332,N_13379);
nand U13541 (N_13541,N_13081,N_13044);
or U13542 (N_13542,N_12100,N_12992);
and U13543 (N_13543,N_12740,N_12213);
xor U13544 (N_13544,N_13066,N_12999);
or U13545 (N_13545,N_13377,N_12798);
nor U13546 (N_13546,N_12291,N_12206);
nand U13547 (N_13547,N_13075,N_12633);
nor U13548 (N_13548,N_12429,N_12580);
nand U13549 (N_13549,N_13468,N_12214);
xor U13550 (N_13550,N_12219,N_12222);
or U13551 (N_13551,N_12045,N_13154);
xnor U13552 (N_13552,N_12195,N_12658);
nand U13553 (N_13553,N_12118,N_13411);
nand U13554 (N_13554,N_13482,N_12880);
or U13555 (N_13555,N_12751,N_12899);
or U13556 (N_13556,N_13193,N_13493);
and U13557 (N_13557,N_13145,N_12831);
nor U13558 (N_13558,N_12561,N_12709);
nand U13559 (N_13559,N_12579,N_12916);
nand U13560 (N_13560,N_12998,N_13295);
nand U13561 (N_13561,N_12638,N_13270);
or U13562 (N_13562,N_13105,N_12469);
and U13563 (N_13563,N_12237,N_13179);
or U13564 (N_13564,N_12602,N_13185);
xor U13565 (N_13565,N_12192,N_12576);
and U13566 (N_13566,N_12570,N_12005);
nor U13567 (N_13567,N_12085,N_13293);
xnor U13568 (N_13568,N_13116,N_13036);
xnor U13569 (N_13569,N_12101,N_12764);
or U13570 (N_13570,N_12261,N_12060);
or U13571 (N_13571,N_13334,N_12169);
nand U13572 (N_13572,N_13133,N_12745);
xnor U13573 (N_13573,N_12523,N_13291);
nand U13574 (N_13574,N_12158,N_12900);
nand U13575 (N_13575,N_12103,N_12491);
nor U13576 (N_13576,N_13003,N_12464);
nand U13577 (N_13577,N_12736,N_13353);
or U13578 (N_13578,N_12828,N_12436);
and U13579 (N_13579,N_12161,N_13225);
xnor U13580 (N_13580,N_13302,N_12107);
nor U13581 (N_13581,N_12556,N_12263);
nand U13582 (N_13582,N_13048,N_12587);
or U13583 (N_13583,N_13326,N_12494);
nor U13584 (N_13584,N_13191,N_12823);
nand U13585 (N_13585,N_12316,N_13307);
or U13586 (N_13586,N_13011,N_12813);
and U13587 (N_13587,N_12412,N_13442);
xnor U13588 (N_13588,N_13376,N_12164);
nand U13589 (N_13589,N_12334,N_13285);
nand U13590 (N_13590,N_12967,N_12907);
and U13591 (N_13591,N_12024,N_12586);
nand U13592 (N_13592,N_12856,N_13182);
nand U13593 (N_13593,N_13336,N_12088);
and U13594 (N_13594,N_12378,N_13323);
or U13595 (N_13595,N_12552,N_12416);
nor U13596 (N_13596,N_12875,N_12618);
and U13597 (N_13597,N_12212,N_12824);
and U13598 (N_13598,N_12652,N_12159);
xor U13599 (N_13599,N_12168,N_12722);
and U13600 (N_13600,N_12019,N_12351);
nor U13601 (N_13601,N_13097,N_12853);
nor U13602 (N_13602,N_13380,N_13390);
nor U13603 (N_13603,N_12965,N_12187);
xnor U13604 (N_13604,N_13210,N_12924);
nor U13605 (N_13605,N_12194,N_13288);
xor U13606 (N_13606,N_12560,N_12271);
and U13607 (N_13607,N_12180,N_12400);
xnor U13608 (N_13608,N_12735,N_13477);
xor U13609 (N_13609,N_13490,N_12966);
or U13610 (N_13610,N_12707,N_13368);
or U13611 (N_13611,N_12634,N_12969);
and U13612 (N_13612,N_12632,N_12444);
nand U13613 (N_13613,N_12435,N_12104);
or U13614 (N_13614,N_12871,N_12275);
or U13615 (N_13615,N_12269,N_13221);
or U13616 (N_13616,N_12309,N_12346);
or U13617 (N_13617,N_13231,N_13200);
nor U13618 (N_13618,N_12787,N_12496);
xor U13619 (N_13619,N_13452,N_12226);
xor U13620 (N_13620,N_12314,N_12595);
and U13621 (N_13621,N_12256,N_12918);
nand U13622 (N_13622,N_13050,N_13207);
or U13623 (N_13623,N_13260,N_13250);
nor U13624 (N_13624,N_13294,N_12616);
and U13625 (N_13625,N_12336,N_13117);
nor U13626 (N_13626,N_12403,N_12270);
xor U13627 (N_13627,N_13004,N_13370);
and U13628 (N_13628,N_13234,N_12859);
xnor U13629 (N_13629,N_12179,N_13022);
nand U13630 (N_13630,N_12018,N_12507);
nand U13631 (N_13631,N_12093,N_13272);
nand U13632 (N_13632,N_12356,N_13283);
and U13633 (N_13633,N_12233,N_12569);
or U13634 (N_13634,N_13318,N_13346);
nand U13635 (N_13635,N_12811,N_13264);
xnor U13636 (N_13636,N_13078,N_13329);
nor U13637 (N_13637,N_12427,N_12487);
and U13638 (N_13638,N_12850,N_13095);
xor U13639 (N_13639,N_12132,N_12303);
xor U13640 (N_13640,N_12762,N_12317);
nor U13641 (N_13641,N_12386,N_13073);
xor U13642 (N_13642,N_12742,N_12779);
nor U13643 (N_13643,N_12202,N_12264);
xor U13644 (N_13644,N_12753,N_12295);
nor U13645 (N_13645,N_12081,N_12963);
or U13646 (N_13646,N_13113,N_13392);
and U13647 (N_13647,N_12348,N_13110);
nand U13648 (N_13648,N_12534,N_13339);
nand U13649 (N_13649,N_13311,N_12796);
xnor U13650 (N_13650,N_12422,N_13172);
and U13651 (N_13651,N_12328,N_12315);
xnor U13652 (N_13652,N_12766,N_12009);
or U13653 (N_13653,N_12841,N_12337);
and U13654 (N_13654,N_12131,N_12234);
nand U13655 (N_13655,N_12077,N_12845);
and U13656 (N_13656,N_13362,N_13451);
nor U13657 (N_13657,N_13181,N_13282);
nand U13658 (N_13658,N_12957,N_13164);
nor U13659 (N_13659,N_12204,N_12769);
and U13660 (N_13660,N_12761,N_12763);
nor U13661 (N_13661,N_13413,N_12364);
nand U13662 (N_13662,N_12703,N_12952);
nand U13663 (N_13663,N_13271,N_13374);
nor U13664 (N_13664,N_13122,N_12913);
xnor U13665 (N_13665,N_13278,N_12228);
nor U13666 (N_13666,N_12861,N_12613);
and U13667 (N_13667,N_12680,N_13287);
and U13668 (N_13668,N_12384,N_13175);
or U13669 (N_13669,N_12719,N_13408);
nor U13670 (N_13670,N_13094,N_13176);
and U13671 (N_13671,N_13254,N_12011);
nand U13672 (N_13672,N_12734,N_13423);
nor U13673 (N_13673,N_12106,N_12227);
nor U13674 (N_13674,N_12962,N_13013);
or U13675 (N_13675,N_13049,N_13330);
xor U13676 (N_13676,N_12837,N_12694);
nor U13677 (N_13677,N_13223,N_12182);
nand U13678 (N_13678,N_12419,N_12663);
nor U13679 (N_13679,N_13183,N_12954);
nand U13680 (N_13680,N_12426,N_13059);
nand U13681 (N_13681,N_12445,N_13258);
nand U13682 (N_13682,N_13047,N_12370);
nand U13683 (N_13683,N_13170,N_12760);
xnor U13684 (N_13684,N_12020,N_12770);
nand U13685 (N_13685,N_12262,N_13280);
nor U13686 (N_13686,N_12743,N_12800);
nor U13687 (N_13687,N_13496,N_13204);
nand U13688 (N_13688,N_12394,N_12588);
or U13689 (N_13689,N_12991,N_12756);
and U13690 (N_13690,N_13249,N_13429);
xor U13691 (N_13691,N_13089,N_13057);
nand U13692 (N_13692,N_13099,N_12790);
and U13693 (N_13693,N_12781,N_12301);
xor U13694 (N_13694,N_12113,N_12341);
nand U13695 (N_13695,N_13373,N_12514);
xor U13696 (N_13696,N_12332,N_12350);
nor U13697 (N_13697,N_13247,N_12276);
nor U13698 (N_13698,N_13243,N_12050);
and U13699 (N_13699,N_12340,N_12460);
xnor U13700 (N_13700,N_12660,N_12806);
and U13701 (N_13701,N_12879,N_12327);
nand U13702 (N_13702,N_12216,N_12512);
xnor U13703 (N_13703,N_12723,N_12597);
or U13704 (N_13704,N_12655,N_12997);
nor U13705 (N_13705,N_13202,N_12319);
and U13706 (N_13706,N_12905,N_12648);
nor U13707 (N_13707,N_12758,N_12198);
xor U13708 (N_13708,N_12865,N_12930);
and U13709 (N_13709,N_12543,N_12895);
or U13710 (N_13710,N_12657,N_13216);
and U13711 (N_13711,N_13268,N_12732);
xnor U13712 (N_13712,N_12479,N_13196);
xnor U13713 (N_13713,N_13188,N_13267);
and U13714 (N_13714,N_12814,N_12151);
nand U13715 (N_13715,N_13153,N_12155);
and U13716 (N_13716,N_12869,N_12649);
xnor U13717 (N_13717,N_13331,N_12369);
xor U13718 (N_13718,N_12955,N_12910);
nand U13719 (N_13719,N_13218,N_12897);
nand U13720 (N_13720,N_12432,N_12883);
xor U13721 (N_13721,N_13042,N_12359);
xor U13722 (N_13722,N_12036,N_12152);
xnor U13723 (N_13723,N_13024,N_12473);
nand U13724 (N_13724,N_12135,N_12160);
or U13725 (N_13725,N_13124,N_13100);
or U13726 (N_13726,N_12728,N_12324);
or U13727 (N_13727,N_12140,N_13152);
and U13728 (N_13728,N_13449,N_13098);
xor U13729 (N_13729,N_12451,N_12274);
or U13730 (N_13730,N_12573,N_12858);
xnor U13731 (N_13731,N_13051,N_12371);
or U13732 (N_13732,N_12934,N_12389);
nor U13733 (N_13733,N_13256,N_12027);
xor U13734 (N_13734,N_12844,N_13103);
and U13735 (N_13735,N_13498,N_13029);
or U13736 (N_13736,N_12970,N_12071);
or U13737 (N_13737,N_13222,N_13383);
xor U13738 (N_13738,N_12960,N_13014);
nor U13739 (N_13739,N_13080,N_12574);
or U13740 (N_13740,N_12345,N_12977);
nor U13741 (N_13741,N_12362,N_12670);
and U13742 (N_13742,N_13150,N_12792);
or U13743 (N_13743,N_13284,N_12529);
nor U13744 (N_13744,N_12840,N_13450);
and U13745 (N_13745,N_12189,N_13091);
or U13746 (N_13746,N_12067,N_12134);
nand U13747 (N_13747,N_12247,N_13273);
xnor U13748 (N_13748,N_13151,N_13286);
xnor U13749 (N_13749,N_13173,N_13206);
and U13750 (N_13750,N_12860,N_13002);
or U13751 (N_13751,N_12842,N_13101);
xnor U13752 (N_13752,N_13178,N_13396);
nor U13753 (N_13753,N_12749,N_12253);
xnor U13754 (N_13754,N_12016,N_12017);
and U13755 (N_13755,N_13483,N_12502);
nor U13756 (N_13756,N_12108,N_12197);
or U13757 (N_13757,N_12443,N_13261);
nor U13758 (N_13758,N_12640,N_12218);
nor U13759 (N_13759,N_13229,N_12912);
and U13760 (N_13760,N_12300,N_12437);
xor U13761 (N_13761,N_12874,N_13056);
nand U13762 (N_13762,N_12083,N_12058);
nor U13763 (N_13763,N_13226,N_12053);
xor U13764 (N_13764,N_12785,N_12456);
xor U13765 (N_13765,N_13365,N_13000);
nor U13766 (N_13766,N_13348,N_13443);
nand U13767 (N_13767,N_13420,N_12626);
and U13768 (N_13768,N_12091,N_12805);
xor U13769 (N_13769,N_12747,N_12133);
nor U13770 (N_13770,N_12682,N_12490);
xor U13771 (N_13771,N_13129,N_12958);
and U13772 (N_13772,N_12231,N_12166);
nor U13773 (N_13773,N_13025,N_12625);
nor U13774 (N_13774,N_13030,N_12668);
or U13775 (N_13775,N_13171,N_12387);
and U13776 (N_13776,N_12925,N_13463);
or U13777 (N_13777,N_13292,N_13359);
xnor U13778 (N_13778,N_12225,N_13475);
nor U13779 (N_13779,N_12903,N_13131);
or U13780 (N_13780,N_12390,N_12636);
and U13781 (N_13781,N_12637,N_12395);
and U13782 (N_13782,N_12409,N_13195);
xor U13783 (N_13783,N_12620,N_12931);
nand U13784 (N_13784,N_12731,N_12522);
nor U13785 (N_13785,N_12510,N_12405);
and U13786 (N_13786,N_12789,N_13015);
nor U13787 (N_13787,N_13055,N_13134);
or U13788 (N_13788,N_12688,N_12553);
or U13789 (N_13789,N_13064,N_12671);
nor U13790 (N_13790,N_12679,N_12368);
nand U13791 (N_13791,N_13354,N_12000);
and U13792 (N_13792,N_12410,N_12235);
nand U13793 (N_13793,N_12313,N_12834);
nand U13794 (N_13794,N_12922,N_12450);
nor U13795 (N_13795,N_13088,N_13404);
nor U13796 (N_13796,N_13426,N_13371);
nand U13797 (N_13797,N_12056,N_13010);
and U13798 (N_13798,N_12557,N_12535);
or U13799 (N_13799,N_12294,N_12447);
xor U13800 (N_13800,N_13084,N_13263);
nand U13801 (N_13801,N_13019,N_12477);
and U13802 (N_13802,N_12944,N_13065);
and U13803 (N_13803,N_12181,N_12217);
nor U13804 (N_13804,N_13240,N_12190);
nor U13805 (N_13805,N_13074,N_12374);
or U13806 (N_13806,N_12248,N_12035);
or U13807 (N_13807,N_12326,N_13069);
nor U13808 (N_13808,N_12839,N_13315);
and U13809 (N_13809,N_12442,N_12457);
nor U13810 (N_13810,N_12074,N_12196);
xnor U13811 (N_13811,N_13464,N_12041);
nor U13812 (N_13812,N_12486,N_13158);
and U13813 (N_13813,N_13155,N_12408);
nor U13814 (N_13814,N_12028,N_12515);
or U13815 (N_13815,N_12628,N_12564);
nor U13816 (N_13816,N_12376,N_13037);
xnor U13817 (N_13817,N_13357,N_12354);
nand U13818 (N_13818,N_12675,N_13470);
nor U13819 (N_13819,N_12746,N_12978);
and U13820 (N_13820,N_12695,N_12791);
nor U13821 (N_13821,N_13149,N_12145);
nand U13822 (N_13822,N_13197,N_12304);
or U13823 (N_13823,N_12372,N_12755);
and U13824 (N_13824,N_13405,N_12305);
xnor U13825 (N_13825,N_12531,N_12984);
xor U13826 (N_13826,N_12778,N_13440);
nor U13827 (N_13827,N_12037,N_12273);
nor U13828 (N_13828,N_12193,N_12175);
or U13829 (N_13829,N_13143,N_13412);
nor U13830 (N_13830,N_13424,N_13304);
or U13831 (N_13831,N_13312,N_12849);
or U13832 (N_13832,N_12873,N_12006);
nor U13833 (N_13833,N_12268,N_12406);
xnor U13834 (N_13834,N_12127,N_12049);
or U13835 (N_13835,N_12544,N_12885);
nor U13836 (N_13836,N_12829,N_12872);
and U13837 (N_13837,N_12012,N_12673);
xnor U13838 (N_13838,N_12566,N_13448);
xor U13839 (N_13839,N_12545,N_13061);
or U13840 (N_13840,N_12210,N_12627);
and U13841 (N_13841,N_12908,N_13156);
or U13842 (N_13842,N_12068,N_12748);
nand U13843 (N_13843,N_12563,N_12882);
or U13844 (N_13844,N_12730,N_12985);
nor U13845 (N_13845,N_12928,N_12794);
or U13846 (N_13846,N_12232,N_12783);
and U13847 (N_13847,N_12996,N_12047);
nand U13848 (N_13848,N_12147,N_12951);
xor U13849 (N_13849,N_12308,N_12765);
or U13850 (N_13850,N_13480,N_12835);
xor U13851 (N_13851,N_12759,N_12177);
nor U13852 (N_13852,N_12495,N_12591);
nor U13853 (N_13853,N_12418,N_12650);
and U13854 (N_13854,N_12741,N_12130);
and U13855 (N_13855,N_13040,N_12286);
nor U13856 (N_13856,N_13135,N_13212);
nor U13857 (N_13857,N_12826,N_12307);
nand U13858 (N_13858,N_12321,N_13104);
and U13859 (N_13859,N_13486,N_12667);
or U13860 (N_13860,N_12793,N_13208);
and U13861 (N_13861,N_13265,N_13198);
or U13862 (N_13862,N_12772,N_13123);
xnor U13863 (N_13863,N_13487,N_12526);
or U13864 (N_13864,N_12712,N_12935);
or U13865 (N_13865,N_13457,N_13281);
nor U13866 (N_13866,N_13485,N_12920);
xnor U13867 (N_13867,N_13043,N_13313);
or U13868 (N_13868,N_12343,N_12565);
xnor U13869 (N_13869,N_12773,N_13275);
and U13870 (N_13870,N_12401,N_12430);
nand U13871 (N_13871,N_12310,N_12122);
and U13872 (N_13872,N_12360,N_12911);
and U13873 (N_13873,N_12272,N_13039);
nor U13874 (N_13874,N_13402,N_13462);
or U13875 (N_13875,N_13211,N_12003);
nor U13876 (N_13876,N_13205,N_13363);
or U13877 (N_13877,N_12710,N_12932);
nand U13878 (N_13878,N_13232,N_13174);
nand U13879 (N_13879,N_12260,N_12605);
or U13880 (N_13880,N_13360,N_13033);
nor U13881 (N_13881,N_13021,N_12174);
nand U13882 (N_13882,N_13092,N_12282);
xnor U13883 (N_13883,N_13324,N_13063);
nor U13884 (N_13884,N_12687,N_12964);
and U13885 (N_13885,N_12646,N_12681);
xor U13886 (N_13886,N_13305,N_12111);
nor U13887 (N_13887,N_12280,N_12221);
xnor U13888 (N_13888,N_12737,N_12142);
and U13889 (N_13889,N_12771,N_12827);
xnor U13890 (N_13890,N_12439,N_12804);
and U13891 (N_13891,N_13233,N_12063);
xnor U13892 (N_13892,N_12980,N_13248);
xnor U13893 (N_13893,N_13194,N_12076);
xor U13894 (N_13894,N_13499,N_13093);
nand U13895 (N_13895,N_12538,N_12939);
xor U13896 (N_13896,N_12843,N_12575);
nand U13897 (N_13897,N_13459,N_12008);
or U13898 (N_13898,N_12815,N_12578);
nor U13899 (N_13899,N_12651,N_12431);
or U13900 (N_13900,N_12143,N_12002);
or U13901 (N_13901,N_13209,N_12645);
nand U13902 (N_13902,N_12901,N_12448);
nor U13903 (N_13903,N_12629,N_13259);
or U13904 (N_13904,N_12540,N_12087);
or U13905 (N_13905,N_12119,N_12536);
nor U13906 (N_13906,N_12521,N_13121);
xnor U13907 (N_13907,N_12698,N_13005);
nand U13908 (N_13908,N_12862,N_12549);
xor U13909 (N_13909,N_13141,N_12623);
nor U13910 (N_13910,N_12267,N_12547);
nand U13911 (N_13911,N_13388,N_12229);
nor U13912 (N_13912,N_12786,N_12097);
nand U13913 (N_13913,N_13186,N_12503);
xnor U13914 (N_13914,N_13192,N_12325);
xnor U13915 (N_13915,N_12562,N_12888);
nor U13916 (N_13916,N_12600,N_12258);
nand U13917 (N_13917,N_13068,N_12809);
xor U13918 (N_13918,N_13403,N_13415);
nor U13919 (N_13919,N_12601,N_12784);
xor U13920 (N_13920,N_12669,N_13125);
xor U13921 (N_13921,N_12023,N_12801);
and U13922 (N_13922,N_12666,N_12959);
xor U13923 (N_13923,N_12867,N_12611);
and U13924 (N_13924,N_12205,N_12539);
and U13925 (N_13925,N_12554,N_13361);
nor U13926 (N_13926,N_12468,N_12363);
and U13927 (N_13927,N_13414,N_12392);
xor U13928 (N_13928,N_12884,N_12073);
xnor U13929 (N_13929,N_12385,N_12846);
nor U13930 (N_13930,N_13384,N_13438);
nand U13931 (N_13931,N_12366,N_12986);
or U13932 (N_13932,N_12022,N_13190);
or U13933 (N_13933,N_12312,N_12713);
xnor U13934 (N_13934,N_12029,N_13220);
xor U13935 (N_13935,N_13465,N_12708);
and U13936 (N_13936,N_13422,N_12767);
nand U13937 (N_13937,N_13053,N_12090);
and U13938 (N_13938,N_13077,N_12344);
nor U13939 (N_13939,N_12092,N_13474);
nor U13940 (N_13940,N_12242,N_13473);
xnor U13941 (N_13941,N_13476,N_12558);
and U13942 (N_13942,N_12176,N_12185);
nor U13943 (N_13943,N_13428,N_12411);
nand U13944 (N_13944,N_13453,N_12084);
or U13945 (N_13945,N_12462,N_12816);
and U13946 (N_13946,N_12750,N_13227);
nor U13947 (N_13947,N_13187,N_12096);
or U13948 (N_13948,N_12148,N_13199);
nand U13949 (N_13949,N_12455,N_12754);
and U13950 (N_13950,N_13118,N_12612);
xnor U13951 (N_13951,N_12171,N_12407);
nand U13952 (N_13952,N_12803,N_13219);
nand U13953 (N_13953,N_12123,N_13335);
nor U13954 (N_13954,N_12676,N_12178);
nor U13955 (N_13955,N_13441,N_12797);
nand U13956 (N_13956,N_13337,N_12705);
or U13957 (N_13957,N_12014,N_12297);
nor U13958 (N_13958,N_12454,N_12812);
or U13959 (N_13959,N_12065,N_12288);
and U13960 (N_13960,N_12320,N_13054);
nor U13961 (N_13961,N_13397,N_12040);
nand U13962 (N_13962,N_12211,N_12739);
nor U13963 (N_13963,N_12546,N_12277);
nand U13964 (N_13964,N_12201,N_12287);
xor U13965 (N_13965,N_12266,N_13203);
nor U13966 (N_13966,N_12572,N_12240);
or U13967 (N_13967,N_13421,N_13217);
or U13968 (N_13968,N_12380,N_12725);
xnor U13969 (N_13969,N_12249,N_12397);
nand U13970 (N_13970,N_12635,N_12662);
and U13971 (N_13971,N_13246,N_12141);
xor U13972 (N_13972,N_12025,N_12484);
or U13973 (N_13973,N_13355,N_12153);
nand U13974 (N_13974,N_12720,N_12015);
xnor U13975 (N_13975,N_12832,N_13008);
or U13976 (N_13976,N_12463,N_13016);
or U13977 (N_13977,N_12347,N_13382);
nor U13978 (N_13978,N_12066,N_12518);
and U13979 (N_13979,N_12654,N_12887);
and U13980 (N_13980,N_12459,N_12223);
and U13981 (N_13981,N_12007,N_12458);
nor U13982 (N_13982,N_12026,N_12738);
or U13983 (N_13983,N_12729,N_12034);
xor U13984 (N_13984,N_12551,N_13358);
xnor U13985 (N_13985,N_12631,N_12252);
nand U13986 (N_13986,N_12391,N_12355);
or U13987 (N_13987,N_12121,N_12128);
xnor U13988 (N_13988,N_12516,N_12674);
xor U13989 (N_13989,N_12039,N_12044);
nand U13990 (N_13990,N_12298,N_12517);
nand U13991 (N_13991,N_12775,N_13045);
nand U13992 (N_13992,N_12684,N_13399);
nor U13993 (N_13993,N_12686,N_13393);
and U13994 (N_13994,N_13255,N_12396);
nor U13995 (N_13995,N_13455,N_12353);
xor U13996 (N_13996,N_12434,N_12055);
xnor U13997 (N_13997,N_12877,N_12881);
xnor U13998 (N_13998,N_13460,N_13023);
xnor U13999 (N_13999,N_13072,N_12945);
nand U14000 (N_14000,N_13279,N_13127);
nor U14001 (N_14001,N_12358,N_12199);
or U14002 (N_14002,N_12377,N_13325);
and U14003 (N_14003,N_13071,N_13401);
xor U14004 (N_14004,N_13310,N_12284);
and U14005 (N_14005,N_13306,N_13046);
or U14006 (N_14006,N_13035,N_13146);
nand U14007 (N_14007,N_12157,N_12504);
xor U14008 (N_14008,N_13168,N_12038);
and U14009 (N_14009,N_12550,N_12030);
nor U14010 (N_14010,N_12520,N_13300);
xnor U14011 (N_14011,N_12296,N_12112);
and U14012 (N_14012,N_12961,N_12059);
nor U14013 (N_14013,N_13189,N_13165);
nor U14014 (N_14014,N_13266,N_12866);
nor U14015 (N_14015,N_12170,N_12365);
nor U14016 (N_14016,N_12339,N_12642);
and U14017 (N_14017,N_12555,N_12972);
nor U14018 (N_14018,N_13058,N_12246);
and U14019 (N_14019,N_12933,N_13114);
xnor U14020 (N_14020,N_12480,N_12335);
nand U14021 (N_14021,N_13262,N_13276);
nor U14022 (N_14022,N_12852,N_13257);
xnor U14023 (N_14023,N_12653,N_12870);
xnor U14024 (N_14024,N_13138,N_13147);
or U14025 (N_14025,N_13245,N_13274);
or U14026 (N_14026,N_12672,N_12822);
xor U14027 (N_14027,N_13177,N_13087);
nand U14028 (N_14028,N_12836,N_12664);
or U14029 (N_14029,N_12208,N_12333);
xor U14030 (N_14030,N_13375,N_12715);
nand U14031 (N_14031,N_13006,N_12149);
or U14032 (N_14032,N_12481,N_12117);
nor U14033 (N_14033,N_12367,N_12609);
or U14034 (N_14034,N_12424,N_12230);
nor U14035 (N_14035,N_12154,N_13425);
xnor U14036 (N_14036,N_12144,N_12678);
or U14037 (N_14037,N_13316,N_12689);
xnor U14038 (N_14038,N_12643,N_12089);
nand U14039 (N_14039,N_13430,N_12665);
or U14040 (N_14040,N_13461,N_12425);
xnor U14041 (N_14041,N_13407,N_12946);
nand U14042 (N_14042,N_13328,N_12968);
nand U14043 (N_14043,N_12979,N_12393);
xnor U14044 (N_14044,N_12820,N_13409);
nor U14045 (N_14045,N_12215,N_12505);
nor U14046 (N_14046,N_13032,N_12095);
nand U14047 (N_14047,N_13418,N_12311);
or U14048 (N_14048,N_13434,N_13427);
nand U14049 (N_14049,N_13031,N_12857);
and U14050 (N_14050,N_13239,N_12528);
or U14051 (N_14051,N_13251,N_12902);
and U14052 (N_14052,N_12876,N_12126);
nor U14053 (N_14053,N_13309,N_12079);
xnor U14054 (N_14054,N_12589,N_12941);
nor U14055 (N_14055,N_12072,N_12808);
nand U14056 (N_14056,N_12500,N_12042);
nand U14057 (N_14057,N_12624,N_13107);
xnor U14058 (N_14058,N_13111,N_12693);
nor U14059 (N_14059,N_12948,N_12656);
nor U14060 (N_14060,N_12990,N_12069);
nor U14061 (N_14061,N_13431,N_12352);
nand U14062 (N_14062,N_13215,N_12567);
xnor U14063 (N_14063,N_12598,N_13327);
and U14064 (N_14064,N_13416,N_12094);
nand U14065 (N_14065,N_12690,N_12914);
and U14066 (N_14066,N_12716,N_13387);
or U14067 (N_14067,N_12251,N_12891);
and U14068 (N_14068,N_13252,N_13038);
nor U14069 (N_14069,N_13052,N_12383);
and U14070 (N_14070,N_12893,N_12603);
or U14071 (N_14071,N_12524,N_12064);
or U14072 (N_14072,N_13369,N_13489);
nor U14073 (N_14073,N_12031,N_12940);
xnor U14074 (N_14074,N_12780,N_12950);
nand U14075 (N_14075,N_12139,N_13060);
nand U14076 (N_14076,N_12483,N_12259);
xnor U14077 (N_14077,N_12537,N_12774);
and U14078 (N_14078,N_12909,N_12582);
nand U14079 (N_14079,N_12621,N_13314);
or U14080 (N_14080,N_12375,N_12021);
nor U14081 (N_14081,N_13244,N_12004);
and U14082 (N_14082,N_13347,N_12075);
nand U14083 (N_14083,N_13301,N_12838);
nand U14084 (N_14084,N_13436,N_12607);
or U14085 (N_14085,N_13398,N_13350);
nand U14086 (N_14086,N_12250,N_12200);
nor U14087 (N_14087,N_12306,N_13070);
nand U14088 (N_14088,N_12470,N_12994);
or U14089 (N_14089,N_12257,N_13082);
nor U14090 (N_14090,N_12802,N_12807);
nand U14091 (N_14091,N_12078,N_12854);
xor U14092 (N_14092,N_13466,N_13290);
and U14093 (N_14093,N_12864,N_13130);
nor U14094 (N_14094,N_12440,N_12508);
nor U14095 (N_14095,N_13319,N_13289);
xnor U14096 (N_14096,N_12349,N_13085);
xnor U14097 (N_14097,N_13308,N_12420);
nand U14098 (N_14098,N_12124,N_12685);
and U14099 (N_14099,N_12847,N_12137);
nor U14100 (N_14100,N_12478,N_12724);
nor U14101 (N_14101,N_12238,N_13142);
xor U14102 (N_14102,N_12942,N_13169);
or U14103 (N_14103,N_12982,N_13356);
or U14104 (N_14104,N_12498,N_12988);
and U14105 (N_14105,N_12191,N_12382);
or U14106 (N_14106,N_13340,N_13017);
xor U14107 (N_14107,N_12989,N_13484);
nor U14108 (N_14108,N_12704,N_13395);
nand U14109 (N_14109,N_13269,N_12896);
or U14110 (N_14110,N_12441,N_12471);
and U14111 (N_14111,N_13317,N_13445);
or U14112 (N_14112,N_13112,N_13344);
or U14113 (N_14113,N_12482,N_13322);
and U14114 (N_14114,N_12173,N_13139);
nor U14115 (N_14115,N_12043,N_12330);
or U14116 (N_14116,N_13163,N_12584);
or U14117 (N_14117,N_12915,N_12207);
nor U14118 (N_14118,N_12165,N_12398);
or U14119 (N_14119,N_12949,N_12289);
nor U14120 (N_14120,N_13062,N_13495);
nor U14121 (N_14121,N_12559,N_13433);
xnor U14122 (N_14122,N_12449,N_12136);
or U14123 (N_14123,N_13106,N_12114);
or U14124 (N_14124,N_13109,N_12886);
nand U14125 (N_14125,N_12239,N_13410);
or U14126 (N_14126,N_12726,N_13435);
or U14127 (N_14127,N_12404,N_13128);
nand U14128 (N_14128,N_13096,N_12357);
xnor U14129 (N_14129,N_12428,N_13026);
or U14130 (N_14130,N_13479,N_12906);
nand U14131 (N_14131,N_13007,N_12244);
or U14132 (N_14132,N_12322,N_12373);
and U14133 (N_14133,N_13235,N_13184);
or U14134 (N_14134,N_12506,N_12138);
xnor U14135 (N_14135,N_12466,N_12501);
nor U14136 (N_14136,N_12279,N_12817);
nor U14137 (N_14137,N_12744,N_13237);
xnor U14138 (N_14138,N_12929,N_12863);
xnor U14139 (N_14139,N_13342,N_12062);
nand U14140 (N_14140,N_12898,N_12833);
xnor U14141 (N_14141,N_12110,N_13439);
or U14142 (N_14142,N_13497,N_12953);
or U14143 (N_14143,N_12414,N_13253);
or U14144 (N_14144,N_12571,N_12116);
and U14145 (N_14145,N_12894,N_13381);
or U14146 (N_14146,N_13079,N_13120);
or U14147 (N_14147,N_12172,N_12492);
xnor U14148 (N_14148,N_13378,N_12696);
or U14149 (N_14149,N_13090,N_12318);
nand U14150 (N_14150,N_12465,N_12583);
xor U14151 (N_14151,N_13027,N_12830);
or U14152 (N_14152,N_12120,N_13366);
nor U14153 (N_14153,N_13467,N_12604);
nand U14154 (N_14154,N_12080,N_13372);
xnor U14155 (N_14155,N_12825,N_12220);
xor U14156 (N_14156,N_12254,N_12699);
or U14157 (N_14157,N_12904,N_13437);
and U14158 (N_14158,N_13086,N_13001);
or U14159 (N_14159,N_13491,N_12013);
or U14160 (N_14160,N_12057,N_12302);
and U14161 (N_14161,N_13157,N_12388);
nor U14162 (N_14162,N_12474,N_12947);
and U14163 (N_14163,N_12167,N_12099);
nor U14164 (N_14164,N_13447,N_12615);
or U14165 (N_14165,N_12892,N_12467);
nor U14166 (N_14166,N_12001,N_12592);
xor U14167 (N_14167,N_13391,N_12499);
and U14168 (N_14168,N_12639,N_12399);
and U14169 (N_14169,N_12452,N_12243);
and U14170 (N_14170,N_13367,N_12105);
nor U14171 (N_14171,N_12702,N_12156);
nor U14172 (N_14172,N_13238,N_12644);
xor U14173 (N_14173,N_12701,N_13136);
xnor U14174 (N_14174,N_13228,N_13102);
xor U14175 (N_14175,N_12299,N_12596);
and U14176 (N_14176,N_13108,N_13076);
or U14177 (N_14177,N_13201,N_12453);
nand U14178 (N_14178,N_12052,N_13020);
or U14179 (N_14179,N_13162,N_12525);
or U14180 (N_14180,N_12599,N_12975);
and U14181 (N_14181,N_12421,N_12919);
xor U14182 (N_14182,N_12290,N_12923);
nand U14183 (N_14183,N_13494,N_12381);
nor U14184 (N_14184,N_13230,N_12086);
xnor U14185 (N_14185,N_12981,N_12878);
and U14186 (N_14186,N_13166,N_13067);
xor U14187 (N_14187,N_13481,N_12987);
nor U14188 (N_14188,N_12423,N_13492);
and U14189 (N_14189,N_12647,N_12971);
or U14190 (N_14190,N_12163,N_13351);
nor U14191 (N_14191,N_12224,N_12983);
nor U14192 (N_14192,N_12659,N_13132);
nor U14193 (N_14193,N_13140,N_12033);
or U14194 (N_14194,N_12727,N_13352);
nand U14195 (N_14195,N_12718,N_13083);
and U14196 (N_14196,N_12209,N_12070);
or U14197 (N_14197,N_13419,N_13296);
or U14198 (N_14198,N_12614,N_12527);
nand U14199 (N_14199,N_13213,N_12183);
nand U14200 (N_14200,N_13148,N_12265);
and U14201 (N_14201,N_12338,N_13241);
xnor U14202 (N_14202,N_12818,N_12417);
xor U14203 (N_14203,N_12630,N_12278);
and U14204 (N_14204,N_12485,N_12361);
nor U14205 (N_14205,N_12255,N_13321);
nand U14206 (N_14206,N_12717,N_12577);
nor U14207 (N_14207,N_12415,N_12585);
nor U14208 (N_14208,N_13446,N_12606);
nor U14209 (N_14209,N_12776,N_12061);
or U14210 (N_14210,N_12433,N_13041);
nand U14211 (N_14211,N_12519,N_13137);
xor U14212 (N_14212,N_12032,N_12281);
nand U14213 (N_14213,N_12851,N_12890);
nand U14214 (N_14214,N_13297,N_12497);
xor U14215 (N_14215,N_12048,N_12608);
nor U14216 (N_14216,N_12581,N_12413);
nand U14217 (N_14217,N_12533,N_12476);
nand U14218 (N_14218,N_12285,N_13298);
nor U14219 (N_14219,N_13406,N_13009);
or U14220 (N_14220,N_12461,N_13028);
nand U14221 (N_14221,N_12782,N_12917);
nor U14222 (N_14222,N_12795,N_12821);
nor U14223 (N_14223,N_12438,N_13458);
nor U14224 (N_14224,N_12956,N_12530);
or U14225 (N_14225,N_12342,N_12548);
nand U14226 (N_14226,N_12974,N_12283);
xor U14227 (N_14227,N_12700,N_12927);
nand U14228 (N_14228,N_12129,N_12568);
xor U14229 (N_14229,N_12697,N_12943);
xnor U14230 (N_14230,N_12768,N_12926);
xor U14231 (N_14231,N_13144,N_13364);
xor U14232 (N_14232,N_12051,N_13320);
or U14233 (N_14233,N_12446,N_13338);
and U14234 (N_14234,N_12757,N_13394);
and U14235 (N_14235,N_12188,N_13160);
and U14236 (N_14236,N_12184,N_13224);
nand U14237 (N_14237,N_12711,N_13299);
or U14238 (N_14238,N_13277,N_12472);
or U14239 (N_14239,N_12162,N_13432);
nand U14240 (N_14240,N_12102,N_12293);
nand U14241 (N_14241,N_12692,N_13034);
or U14242 (N_14242,N_12752,N_12995);
or U14243 (N_14243,N_12331,N_12617);
xnor U14244 (N_14244,N_12513,N_13115);
nand U14245 (N_14245,N_12402,N_12938);
xnor U14246 (N_14246,N_13012,N_12677);
nand U14247 (N_14247,N_12054,N_13386);
and U14248 (N_14248,N_12511,N_12868);
nand U14249 (N_14249,N_13400,N_12936);
nand U14250 (N_14250,N_12705,N_13354);
or U14251 (N_14251,N_13448,N_12931);
xnor U14252 (N_14252,N_13069,N_13241);
nand U14253 (N_14253,N_12119,N_12535);
nor U14254 (N_14254,N_12313,N_12858);
and U14255 (N_14255,N_12708,N_12509);
or U14256 (N_14256,N_13315,N_12382);
xnor U14257 (N_14257,N_13004,N_12239);
and U14258 (N_14258,N_13330,N_12604);
xnor U14259 (N_14259,N_13489,N_12600);
or U14260 (N_14260,N_12132,N_12741);
xor U14261 (N_14261,N_13406,N_12542);
xor U14262 (N_14262,N_13392,N_12056);
nor U14263 (N_14263,N_12442,N_12447);
or U14264 (N_14264,N_13483,N_13308);
or U14265 (N_14265,N_13027,N_12022);
and U14266 (N_14266,N_13089,N_12554);
nand U14267 (N_14267,N_12204,N_13346);
and U14268 (N_14268,N_12529,N_12950);
and U14269 (N_14269,N_12484,N_13270);
or U14270 (N_14270,N_12256,N_12442);
and U14271 (N_14271,N_12229,N_12773);
nor U14272 (N_14272,N_12808,N_12353);
nand U14273 (N_14273,N_13270,N_12552);
or U14274 (N_14274,N_12953,N_13239);
or U14275 (N_14275,N_12376,N_13199);
xnor U14276 (N_14276,N_12148,N_13373);
nor U14277 (N_14277,N_13132,N_12229);
nand U14278 (N_14278,N_13371,N_13180);
and U14279 (N_14279,N_13280,N_13011);
nor U14280 (N_14280,N_13345,N_12834);
nor U14281 (N_14281,N_12333,N_13132);
xor U14282 (N_14282,N_12971,N_12538);
nor U14283 (N_14283,N_12980,N_12403);
or U14284 (N_14284,N_12336,N_12611);
nor U14285 (N_14285,N_12415,N_13027);
xor U14286 (N_14286,N_13464,N_12756);
or U14287 (N_14287,N_12584,N_12727);
xnor U14288 (N_14288,N_12240,N_13234);
and U14289 (N_14289,N_13400,N_13095);
or U14290 (N_14290,N_13323,N_13299);
and U14291 (N_14291,N_13250,N_12642);
nor U14292 (N_14292,N_13113,N_12308);
nand U14293 (N_14293,N_13372,N_12173);
xor U14294 (N_14294,N_13015,N_12736);
xor U14295 (N_14295,N_12963,N_12880);
nor U14296 (N_14296,N_13209,N_12107);
nor U14297 (N_14297,N_12372,N_12384);
nand U14298 (N_14298,N_12979,N_12831);
xor U14299 (N_14299,N_12681,N_12579);
or U14300 (N_14300,N_12309,N_12327);
nand U14301 (N_14301,N_12672,N_12514);
xnor U14302 (N_14302,N_12088,N_13472);
xnor U14303 (N_14303,N_12330,N_12632);
and U14304 (N_14304,N_12288,N_12176);
nand U14305 (N_14305,N_12325,N_13010);
xor U14306 (N_14306,N_12064,N_12822);
xor U14307 (N_14307,N_12865,N_12879);
or U14308 (N_14308,N_13069,N_13223);
and U14309 (N_14309,N_12948,N_12724);
nor U14310 (N_14310,N_12604,N_12952);
and U14311 (N_14311,N_12184,N_12246);
xnor U14312 (N_14312,N_13486,N_12865);
nand U14313 (N_14313,N_12069,N_12834);
nand U14314 (N_14314,N_12128,N_13004);
or U14315 (N_14315,N_12225,N_12617);
and U14316 (N_14316,N_12111,N_13353);
nand U14317 (N_14317,N_12057,N_12665);
nor U14318 (N_14318,N_13414,N_13363);
nand U14319 (N_14319,N_12734,N_13287);
and U14320 (N_14320,N_12601,N_13354);
xor U14321 (N_14321,N_12528,N_12204);
nor U14322 (N_14322,N_13421,N_13347);
and U14323 (N_14323,N_12658,N_12837);
or U14324 (N_14324,N_13226,N_13361);
or U14325 (N_14325,N_12230,N_12343);
and U14326 (N_14326,N_12833,N_12738);
xor U14327 (N_14327,N_13430,N_12803);
nand U14328 (N_14328,N_13218,N_13059);
nor U14329 (N_14329,N_12829,N_12491);
nand U14330 (N_14330,N_13259,N_12477);
nor U14331 (N_14331,N_13067,N_13144);
xor U14332 (N_14332,N_13246,N_12106);
or U14333 (N_14333,N_12498,N_12197);
and U14334 (N_14334,N_12634,N_12897);
nor U14335 (N_14335,N_13276,N_12835);
nor U14336 (N_14336,N_13475,N_13080);
nor U14337 (N_14337,N_12044,N_13243);
and U14338 (N_14338,N_12166,N_12047);
and U14339 (N_14339,N_13399,N_12796);
and U14340 (N_14340,N_12935,N_12440);
xor U14341 (N_14341,N_12351,N_12743);
nand U14342 (N_14342,N_13162,N_12786);
and U14343 (N_14343,N_12382,N_13279);
nor U14344 (N_14344,N_12806,N_12859);
nor U14345 (N_14345,N_12279,N_13181);
xor U14346 (N_14346,N_12856,N_12728);
and U14347 (N_14347,N_12640,N_12886);
and U14348 (N_14348,N_13371,N_12723);
or U14349 (N_14349,N_13096,N_12683);
nor U14350 (N_14350,N_12247,N_12723);
nor U14351 (N_14351,N_12097,N_12514);
nor U14352 (N_14352,N_13419,N_12894);
nand U14353 (N_14353,N_12524,N_12624);
xnor U14354 (N_14354,N_12152,N_12591);
xnor U14355 (N_14355,N_12795,N_12842);
or U14356 (N_14356,N_12862,N_12332);
xor U14357 (N_14357,N_13463,N_13211);
and U14358 (N_14358,N_12166,N_12104);
nor U14359 (N_14359,N_12629,N_13430);
or U14360 (N_14360,N_12565,N_13346);
and U14361 (N_14361,N_12970,N_13343);
and U14362 (N_14362,N_13274,N_12657);
and U14363 (N_14363,N_13223,N_13496);
xnor U14364 (N_14364,N_12442,N_13032);
and U14365 (N_14365,N_12041,N_13399);
or U14366 (N_14366,N_12440,N_12866);
or U14367 (N_14367,N_12983,N_12606);
nand U14368 (N_14368,N_12918,N_12959);
or U14369 (N_14369,N_13499,N_12848);
nor U14370 (N_14370,N_12473,N_13420);
xor U14371 (N_14371,N_13198,N_13144);
xnor U14372 (N_14372,N_12745,N_12096);
or U14373 (N_14373,N_12658,N_12358);
nand U14374 (N_14374,N_12673,N_13114);
nand U14375 (N_14375,N_13439,N_12183);
and U14376 (N_14376,N_12041,N_12293);
nand U14377 (N_14377,N_12296,N_12606);
xor U14378 (N_14378,N_12653,N_12672);
xor U14379 (N_14379,N_12008,N_13037);
nand U14380 (N_14380,N_13219,N_12922);
or U14381 (N_14381,N_12937,N_12647);
xor U14382 (N_14382,N_12089,N_13079);
xnor U14383 (N_14383,N_12866,N_12559);
xnor U14384 (N_14384,N_13155,N_13389);
or U14385 (N_14385,N_12900,N_12884);
nor U14386 (N_14386,N_13446,N_12813);
nand U14387 (N_14387,N_12157,N_12619);
and U14388 (N_14388,N_12007,N_12769);
nand U14389 (N_14389,N_12644,N_12773);
and U14390 (N_14390,N_12378,N_12904);
nand U14391 (N_14391,N_12967,N_12471);
nand U14392 (N_14392,N_13498,N_13158);
and U14393 (N_14393,N_12435,N_12252);
nand U14394 (N_14394,N_12515,N_13449);
or U14395 (N_14395,N_13118,N_12335);
or U14396 (N_14396,N_13212,N_12756);
or U14397 (N_14397,N_12255,N_12566);
nand U14398 (N_14398,N_12491,N_12051);
and U14399 (N_14399,N_13252,N_12911);
nand U14400 (N_14400,N_13021,N_12499);
and U14401 (N_14401,N_13122,N_13258);
and U14402 (N_14402,N_12422,N_12420);
or U14403 (N_14403,N_12168,N_12537);
nand U14404 (N_14404,N_12945,N_12435);
and U14405 (N_14405,N_12131,N_12600);
xor U14406 (N_14406,N_12612,N_12659);
nand U14407 (N_14407,N_13330,N_12444);
nand U14408 (N_14408,N_12682,N_12310);
or U14409 (N_14409,N_12776,N_12694);
or U14410 (N_14410,N_12085,N_12730);
and U14411 (N_14411,N_13285,N_13458);
nor U14412 (N_14412,N_12234,N_12410);
or U14413 (N_14413,N_13188,N_13234);
or U14414 (N_14414,N_13096,N_12053);
or U14415 (N_14415,N_12110,N_12780);
xor U14416 (N_14416,N_12330,N_13190);
or U14417 (N_14417,N_12758,N_12249);
or U14418 (N_14418,N_12585,N_12388);
and U14419 (N_14419,N_12457,N_12234);
and U14420 (N_14420,N_12275,N_13279);
nor U14421 (N_14421,N_12831,N_12050);
and U14422 (N_14422,N_13223,N_12071);
or U14423 (N_14423,N_12103,N_13457);
nor U14424 (N_14424,N_13450,N_13485);
nand U14425 (N_14425,N_12183,N_13384);
and U14426 (N_14426,N_12785,N_12032);
or U14427 (N_14427,N_12702,N_13290);
nor U14428 (N_14428,N_12233,N_13182);
or U14429 (N_14429,N_12387,N_13241);
and U14430 (N_14430,N_13400,N_12112);
nand U14431 (N_14431,N_13013,N_12816);
and U14432 (N_14432,N_13424,N_12085);
and U14433 (N_14433,N_12342,N_12397);
nand U14434 (N_14434,N_13210,N_12098);
xnor U14435 (N_14435,N_12290,N_13095);
or U14436 (N_14436,N_13411,N_12888);
or U14437 (N_14437,N_13170,N_12063);
nor U14438 (N_14438,N_12998,N_12634);
or U14439 (N_14439,N_12253,N_12504);
nand U14440 (N_14440,N_13047,N_13043);
xor U14441 (N_14441,N_12760,N_12104);
xnor U14442 (N_14442,N_12048,N_13334);
and U14443 (N_14443,N_12846,N_13272);
nor U14444 (N_14444,N_12154,N_13030);
nor U14445 (N_14445,N_12308,N_12552);
and U14446 (N_14446,N_12511,N_12776);
xnor U14447 (N_14447,N_12146,N_13238);
xor U14448 (N_14448,N_12412,N_13117);
or U14449 (N_14449,N_12607,N_12419);
nand U14450 (N_14450,N_12470,N_12089);
xor U14451 (N_14451,N_12345,N_12628);
nor U14452 (N_14452,N_12279,N_12816);
nor U14453 (N_14453,N_13425,N_13172);
nor U14454 (N_14454,N_12325,N_12290);
xnor U14455 (N_14455,N_13362,N_12545);
nand U14456 (N_14456,N_12651,N_12239);
nand U14457 (N_14457,N_12911,N_13026);
nand U14458 (N_14458,N_13032,N_12121);
or U14459 (N_14459,N_12644,N_13414);
and U14460 (N_14460,N_12757,N_12561);
xnor U14461 (N_14461,N_12859,N_12241);
and U14462 (N_14462,N_12627,N_12583);
nand U14463 (N_14463,N_12717,N_12125);
xor U14464 (N_14464,N_13289,N_12865);
and U14465 (N_14465,N_13331,N_12780);
nand U14466 (N_14466,N_12981,N_12009);
nor U14467 (N_14467,N_12199,N_13262);
or U14468 (N_14468,N_12933,N_12827);
and U14469 (N_14469,N_12557,N_12719);
nand U14470 (N_14470,N_12341,N_12058);
and U14471 (N_14471,N_12079,N_13139);
xor U14472 (N_14472,N_12730,N_12402);
nor U14473 (N_14473,N_13167,N_13475);
or U14474 (N_14474,N_12139,N_12789);
xnor U14475 (N_14475,N_12069,N_12505);
xor U14476 (N_14476,N_13410,N_12401);
nand U14477 (N_14477,N_13121,N_12830);
nand U14478 (N_14478,N_12377,N_12825);
nor U14479 (N_14479,N_13239,N_12031);
xor U14480 (N_14480,N_13089,N_12066);
nor U14481 (N_14481,N_13376,N_12183);
or U14482 (N_14482,N_12660,N_12470);
nand U14483 (N_14483,N_12568,N_12713);
and U14484 (N_14484,N_12246,N_13439);
or U14485 (N_14485,N_12032,N_12589);
xor U14486 (N_14486,N_12110,N_13146);
nor U14487 (N_14487,N_12264,N_12761);
xnor U14488 (N_14488,N_12879,N_12638);
and U14489 (N_14489,N_13317,N_12533);
and U14490 (N_14490,N_12193,N_12527);
xor U14491 (N_14491,N_13173,N_12460);
or U14492 (N_14492,N_12065,N_12902);
and U14493 (N_14493,N_13132,N_12190);
nor U14494 (N_14494,N_13112,N_12497);
xor U14495 (N_14495,N_12281,N_12833);
nand U14496 (N_14496,N_12823,N_12561);
or U14497 (N_14497,N_13247,N_12343);
xnor U14498 (N_14498,N_12956,N_12292);
xor U14499 (N_14499,N_12364,N_12529);
and U14500 (N_14500,N_13304,N_13148);
or U14501 (N_14501,N_13456,N_12916);
nor U14502 (N_14502,N_12623,N_12475);
nand U14503 (N_14503,N_13261,N_12493);
and U14504 (N_14504,N_12012,N_13427);
xor U14505 (N_14505,N_13035,N_13206);
xor U14506 (N_14506,N_13017,N_13028);
or U14507 (N_14507,N_12923,N_13010);
and U14508 (N_14508,N_13091,N_12419);
xnor U14509 (N_14509,N_12464,N_12024);
or U14510 (N_14510,N_13251,N_13122);
nand U14511 (N_14511,N_13023,N_13221);
nor U14512 (N_14512,N_13185,N_12246);
and U14513 (N_14513,N_12290,N_12059);
nor U14514 (N_14514,N_13155,N_12823);
xor U14515 (N_14515,N_12839,N_13433);
nand U14516 (N_14516,N_12187,N_12795);
nor U14517 (N_14517,N_13153,N_13141);
nand U14518 (N_14518,N_12924,N_12173);
and U14519 (N_14519,N_12515,N_13255);
or U14520 (N_14520,N_12065,N_12200);
nand U14521 (N_14521,N_12650,N_12473);
or U14522 (N_14522,N_12109,N_12483);
xor U14523 (N_14523,N_12616,N_12077);
xnor U14524 (N_14524,N_12959,N_12742);
xor U14525 (N_14525,N_12721,N_12656);
nand U14526 (N_14526,N_12282,N_13307);
nor U14527 (N_14527,N_12718,N_12675);
xor U14528 (N_14528,N_13142,N_12623);
nand U14529 (N_14529,N_12185,N_13452);
nand U14530 (N_14530,N_12042,N_13119);
or U14531 (N_14531,N_13018,N_12816);
nor U14532 (N_14532,N_12674,N_12701);
xnor U14533 (N_14533,N_12028,N_12485);
or U14534 (N_14534,N_12311,N_12692);
and U14535 (N_14535,N_12167,N_12497);
and U14536 (N_14536,N_13103,N_12252);
and U14537 (N_14537,N_12187,N_12614);
xnor U14538 (N_14538,N_13335,N_12934);
xnor U14539 (N_14539,N_12029,N_12580);
xor U14540 (N_14540,N_13475,N_12737);
nor U14541 (N_14541,N_12266,N_13279);
or U14542 (N_14542,N_13012,N_12804);
xnor U14543 (N_14543,N_12893,N_12967);
and U14544 (N_14544,N_13142,N_13095);
and U14545 (N_14545,N_12997,N_12328);
nor U14546 (N_14546,N_12603,N_13237);
and U14547 (N_14547,N_13454,N_12183);
nor U14548 (N_14548,N_13456,N_12185);
nand U14549 (N_14549,N_12850,N_12008);
nor U14550 (N_14550,N_12194,N_12865);
and U14551 (N_14551,N_13074,N_12854);
nand U14552 (N_14552,N_12600,N_12396);
nand U14553 (N_14553,N_12259,N_13404);
xnor U14554 (N_14554,N_12787,N_13206);
xor U14555 (N_14555,N_12407,N_12913);
xnor U14556 (N_14556,N_13232,N_13325);
or U14557 (N_14557,N_12483,N_13322);
nand U14558 (N_14558,N_13189,N_13172);
and U14559 (N_14559,N_12521,N_12383);
xor U14560 (N_14560,N_12715,N_12442);
or U14561 (N_14561,N_12068,N_13395);
nor U14562 (N_14562,N_12017,N_12035);
nand U14563 (N_14563,N_12625,N_12624);
nor U14564 (N_14564,N_12215,N_13470);
and U14565 (N_14565,N_12272,N_12164);
and U14566 (N_14566,N_13072,N_13365);
nand U14567 (N_14567,N_13314,N_12529);
nand U14568 (N_14568,N_13260,N_12176);
or U14569 (N_14569,N_12303,N_12782);
xor U14570 (N_14570,N_12529,N_12329);
nand U14571 (N_14571,N_13255,N_12964);
and U14572 (N_14572,N_12461,N_13139);
and U14573 (N_14573,N_12986,N_13187);
nor U14574 (N_14574,N_12005,N_13115);
nand U14575 (N_14575,N_13423,N_13108);
nand U14576 (N_14576,N_12383,N_12470);
nor U14577 (N_14577,N_12720,N_12974);
nand U14578 (N_14578,N_12814,N_13084);
or U14579 (N_14579,N_13316,N_13196);
nand U14580 (N_14580,N_12546,N_13085);
xnor U14581 (N_14581,N_12489,N_12832);
xor U14582 (N_14582,N_13478,N_13222);
or U14583 (N_14583,N_12450,N_13337);
nand U14584 (N_14584,N_12987,N_12766);
or U14585 (N_14585,N_12951,N_12781);
nand U14586 (N_14586,N_12094,N_12649);
and U14587 (N_14587,N_13136,N_13061);
nor U14588 (N_14588,N_12169,N_12004);
nand U14589 (N_14589,N_12770,N_12239);
and U14590 (N_14590,N_13260,N_13054);
nor U14591 (N_14591,N_13214,N_12855);
xor U14592 (N_14592,N_12573,N_12786);
nor U14593 (N_14593,N_13337,N_12451);
or U14594 (N_14594,N_13467,N_13360);
nor U14595 (N_14595,N_12876,N_12107);
xnor U14596 (N_14596,N_12236,N_12878);
xnor U14597 (N_14597,N_12141,N_13212);
and U14598 (N_14598,N_13120,N_13016);
nor U14599 (N_14599,N_12204,N_13344);
xnor U14600 (N_14600,N_13020,N_12216);
xor U14601 (N_14601,N_13205,N_12840);
nand U14602 (N_14602,N_12134,N_12531);
and U14603 (N_14603,N_12814,N_12568);
nor U14604 (N_14604,N_12311,N_12637);
nand U14605 (N_14605,N_12681,N_12175);
or U14606 (N_14606,N_12098,N_12288);
and U14607 (N_14607,N_13002,N_12753);
nor U14608 (N_14608,N_12810,N_12874);
nor U14609 (N_14609,N_12880,N_12207);
and U14610 (N_14610,N_13005,N_12230);
nand U14611 (N_14611,N_12539,N_13358);
nor U14612 (N_14612,N_12521,N_13227);
and U14613 (N_14613,N_13485,N_12729);
nor U14614 (N_14614,N_13047,N_13075);
xor U14615 (N_14615,N_12738,N_13495);
or U14616 (N_14616,N_12009,N_12603);
nor U14617 (N_14617,N_12872,N_13195);
nand U14618 (N_14618,N_12573,N_12834);
nand U14619 (N_14619,N_13474,N_12835);
xor U14620 (N_14620,N_13439,N_13329);
xnor U14621 (N_14621,N_13310,N_12754);
xnor U14622 (N_14622,N_12977,N_12284);
nor U14623 (N_14623,N_13415,N_13423);
or U14624 (N_14624,N_12639,N_13341);
or U14625 (N_14625,N_12503,N_13087);
nor U14626 (N_14626,N_12468,N_12202);
and U14627 (N_14627,N_12324,N_12837);
or U14628 (N_14628,N_12047,N_12631);
nor U14629 (N_14629,N_13481,N_12849);
nand U14630 (N_14630,N_12801,N_12184);
and U14631 (N_14631,N_12941,N_12902);
nand U14632 (N_14632,N_12198,N_13344);
and U14633 (N_14633,N_12479,N_13065);
nand U14634 (N_14634,N_12111,N_12917);
xor U14635 (N_14635,N_12197,N_12567);
nor U14636 (N_14636,N_12872,N_13383);
nand U14637 (N_14637,N_12341,N_12823);
xnor U14638 (N_14638,N_13298,N_13108);
nand U14639 (N_14639,N_12466,N_12355);
nand U14640 (N_14640,N_13029,N_12064);
or U14641 (N_14641,N_12788,N_12629);
nand U14642 (N_14642,N_13474,N_12714);
nor U14643 (N_14643,N_12107,N_12353);
nand U14644 (N_14644,N_13117,N_12005);
nor U14645 (N_14645,N_13431,N_12081);
or U14646 (N_14646,N_13110,N_13042);
or U14647 (N_14647,N_13364,N_12616);
nor U14648 (N_14648,N_13266,N_12673);
and U14649 (N_14649,N_12061,N_13322);
and U14650 (N_14650,N_12853,N_13282);
nor U14651 (N_14651,N_12630,N_13126);
xnor U14652 (N_14652,N_12025,N_12900);
nand U14653 (N_14653,N_13259,N_12859);
nor U14654 (N_14654,N_12311,N_13066);
nand U14655 (N_14655,N_12085,N_12090);
nor U14656 (N_14656,N_12624,N_12875);
nand U14657 (N_14657,N_13373,N_13154);
nor U14658 (N_14658,N_13281,N_13023);
nand U14659 (N_14659,N_12289,N_12495);
and U14660 (N_14660,N_12345,N_12816);
and U14661 (N_14661,N_12102,N_12559);
xnor U14662 (N_14662,N_12489,N_12833);
nand U14663 (N_14663,N_12981,N_12941);
nand U14664 (N_14664,N_12856,N_13378);
or U14665 (N_14665,N_13084,N_12727);
xnor U14666 (N_14666,N_12656,N_12622);
and U14667 (N_14667,N_12387,N_12800);
nor U14668 (N_14668,N_12487,N_12248);
nor U14669 (N_14669,N_12012,N_13311);
and U14670 (N_14670,N_12524,N_13133);
nor U14671 (N_14671,N_12071,N_12810);
nand U14672 (N_14672,N_12546,N_12833);
xnor U14673 (N_14673,N_13338,N_12047);
nand U14674 (N_14674,N_12790,N_12633);
nand U14675 (N_14675,N_12687,N_13176);
and U14676 (N_14676,N_12684,N_13497);
xor U14677 (N_14677,N_13360,N_13319);
nand U14678 (N_14678,N_13407,N_12383);
or U14679 (N_14679,N_12812,N_13236);
or U14680 (N_14680,N_13099,N_12228);
or U14681 (N_14681,N_13328,N_12791);
and U14682 (N_14682,N_13344,N_12291);
nor U14683 (N_14683,N_13129,N_13077);
xor U14684 (N_14684,N_13176,N_13493);
and U14685 (N_14685,N_12052,N_13334);
nand U14686 (N_14686,N_12650,N_12826);
nor U14687 (N_14687,N_12557,N_12124);
nand U14688 (N_14688,N_12840,N_13230);
xor U14689 (N_14689,N_12539,N_12620);
nor U14690 (N_14690,N_12234,N_12050);
xnor U14691 (N_14691,N_12831,N_13490);
and U14692 (N_14692,N_12672,N_12163);
nor U14693 (N_14693,N_12451,N_13063);
and U14694 (N_14694,N_13296,N_13376);
nand U14695 (N_14695,N_12333,N_12870);
and U14696 (N_14696,N_12883,N_12438);
xor U14697 (N_14697,N_12922,N_13493);
and U14698 (N_14698,N_12236,N_12152);
nor U14699 (N_14699,N_12906,N_13130);
nor U14700 (N_14700,N_12513,N_13480);
xnor U14701 (N_14701,N_12813,N_12199);
and U14702 (N_14702,N_12000,N_12172);
xnor U14703 (N_14703,N_12078,N_13183);
nand U14704 (N_14704,N_12756,N_12173);
xor U14705 (N_14705,N_13108,N_12044);
nor U14706 (N_14706,N_13016,N_12257);
or U14707 (N_14707,N_12480,N_12663);
xnor U14708 (N_14708,N_12177,N_12193);
xnor U14709 (N_14709,N_12661,N_12509);
and U14710 (N_14710,N_12335,N_13417);
nand U14711 (N_14711,N_12831,N_12846);
nand U14712 (N_14712,N_12199,N_12084);
nor U14713 (N_14713,N_13175,N_12587);
xor U14714 (N_14714,N_12608,N_12605);
or U14715 (N_14715,N_12008,N_13360);
or U14716 (N_14716,N_13194,N_13383);
or U14717 (N_14717,N_12327,N_12845);
or U14718 (N_14718,N_13260,N_12013);
xnor U14719 (N_14719,N_13001,N_12325);
and U14720 (N_14720,N_13070,N_12192);
nor U14721 (N_14721,N_13497,N_12472);
and U14722 (N_14722,N_12977,N_12565);
or U14723 (N_14723,N_13178,N_12357);
xor U14724 (N_14724,N_12542,N_13215);
nor U14725 (N_14725,N_12728,N_12051);
nor U14726 (N_14726,N_12686,N_12535);
nor U14727 (N_14727,N_12257,N_12707);
or U14728 (N_14728,N_12186,N_12745);
nor U14729 (N_14729,N_12649,N_12762);
xnor U14730 (N_14730,N_12348,N_13345);
or U14731 (N_14731,N_12998,N_13036);
xnor U14732 (N_14732,N_12490,N_12379);
xor U14733 (N_14733,N_12056,N_12178);
nor U14734 (N_14734,N_12684,N_12996);
and U14735 (N_14735,N_12354,N_13452);
xnor U14736 (N_14736,N_12145,N_13392);
and U14737 (N_14737,N_12474,N_13139);
and U14738 (N_14738,N_12167,N_13285);
nor U14739 (N_14739,N_12763,N_12040);
or U14740 (N_14740,N_12222,N_13316);
and U14741 (N_14741,N_13061,N_12420);
nand U14742 (N_14742,N_13153,N_12953);
nor U14743 (N_14743,N_12424,N_12449);
and U14744 (N_14744,N_12747,N_12205);
nand U14745 (N_14745,N_12648,N_12260);
nor U14746 (N_14746,N_13347,N_13158);
or U14747 (N_14747,N_13003,N_12773);
nand U14748 (N_14748,N_12088,N_12881);
xor U14749 (N_14749,N_13349,N_12873);
nor U14750 (N_14750,N_12337,N_13268);
nand U14751 (N_14751,N_12722,N_13333);
xor U14752 (N_14752,N_12002,N_12206);
nand U14753 (N_14753,N_12125,N_13423);
xor U14754 (N_14754,N_12412,N_13164);
and U14755 (N_14755,N_12632,N_13125);
and U14756 (N_14756,N_12570,N_13282);
nor U14757 (N_14757,N_12950,N_12877);
nor U14758 (N_14758,N_13301,N_12592);
or U14759 (N_14759,N_13062,N_12301);
nand U14760 (N_14760,N_12231,N_12592);
or U14761 (N_14761,N_12226,N_12772);
or U14762 (N_14762,N_13352,N_12646);
or U14763 (N_14763,N_12219,N_13147);
nand U14764 (N_14764,N_12421,N_13023);
nand U14765 (N_14765,N_12364,N_13023);
xnor U14766 (N_14766,N_12780,N_13314);
nor U14767 (N_14767,N_12182,N_12480);
or U14768 (N_14768,N_12862,N_12269);
or U14769 (N_14769,N_12099,N_13011);
xnor U14770 (N_14770,N_12562,N_13206);
xnor U14771 (N_14771,N_12108,N_12650);
nand U14772 (N_14772,N_12564,N_12878);
nand U14773 (N_14773,N_12699,N_12931);
nor U14774 (N_14774,N_12781,N_12799);
xnor U14775 (N_14775,N_12702,N_13087);
nor U14776 (N_14776,N_13402,N_12503);
nor U14777 (N_14777,N_13082,N_12712);
and U14778 (N_14778,N_12483,N_13422);
nor U14779 (N_14779,N_13241,N_12423);
and U14780 (N_14780,N_12065,N_13446);
xnor U14781 (N_14781,N_13170,N_12647);
xor U14782 (N_14782,N_12534,N_12175);
nor U14783 (N_14783,N_12402,N_12060);
or U14784 (N_14784,N_13073,N_12045);
xor U14785 (N_14785,N_12591,N_12100);
nor U14786 (N_14786,N_13257,N_12445);
and U14787 (N_14787,N_12325,N_12066);
nand U14788 (N_14788,N_13487,N_12861);
xor U14789 (N_14789,N_12619,N_13390);
nand U14790 (N_14790,N_12612,N_13190);
xor U14791 (N_14791,N_12223,N_13196);
nor U14792 (N_14792,N_13491,N_13381);
nor U14793 (N_14793,N_12611,N_12392);
nor U14794 (N_14794,N_13290,N_12383);
nand U14795 (N_14795,N_13199,N_12536);
nor U14796 (N_14796,N_13336,N_12215);
nand U14797 (N_14797,N_12435,N_12829);
xor U14798 (N_14798,N_12715,N_13312);
xnor U14799 (N_14799,N_12308,N_13220);
xnor U14800 (N_14800,N_13120,N_13465);
nor U14801 (N_14801,N_12370,N_13467);
xor U14802 (N_14802,N_13273,N_12661);
and U14803 (N_14803,N_13111,N_12051);
and U14804 (N_14804,N_12377,N_12151);
nand U14805 (N_14805,N_12987,N_12068);
and U14806 (N_14806,N_12873,N_12437);
and U14807 (N_14807,N_13366,N_12969);
or U14808 (N_14808,N_12218,N_12374);
or U14809 (N_14809,N_12263,N_13211);
xnor U14810 (N_14810,N_12743,N_12121);
nor U14811 (N_14811,N_12687,N_12989);
nand U14812 (N_14812,N_12013,N_13448);
xnor U14813 (N_14813,N_12487,N_13067);
and U14814 (N_14814,N_12622,N_12792);
or U14815 (N_14815,N_12237,N_12806);
nand U14816 (N_14816,N_13223,N_12908);
xnor U14817 (N_14817,N_12326,N_12800);
or U14818 (N_14818,N_12745,N_12779);
and U14819 (N_14819,N_13254,N_13366);
nor U14820 (N_14820,N_13118,N_12464);
nor U14821 (N_14821,N_12616,N_12834);
and U14822 (N_14822,N_12283,N_12194);
and U14823 (N_14823,N_13226,N_12854);
nor U14824 (N_14824,N_13275,N_13424);
or U14825 (N_14825,N_13152,N_12029);
and U14826 (N_14826,N_12250,N_13056);
or U14827 (N_14827,N_12086,N_12404);
nor U14828 (N_14828,N_12120,N_12440);
nand U14829 (N_14829,N_12597,N_12549);
xnor U14830 (N_14830,N_12576,N_12409);
and U14831 (N_14831,N_13061,N_12363);
nor U14832 (N_14832,N_13398,N_12300);
xor U14833 (N_14833,N_12426,N_13356);
or U14834 (N_14834,N_13492,N_12148);
nand U14835 (N_14835,N_12201,N_12847);
or U14836 (N_14836,N_12836,N_12102);
nor U14837 (N_14837,N_12215,N_13496);
nand U14838 (N_14838,N_12848,N_12589);
or U14839 (N_14839,N_13137,N_12035);
xor U14840 (N_14840,N_13142,N_13227);
nor U14841 (N_14841,N_13180,N_12560);
xor U14842 (N_14842,N_13399,N_12825);
or U14843 (N_14843,N_12512,N_13318);
and U14844 (N_14844,N_12963,N_13331);
or U14845 (N_14845,N_12195,N_13014);
nand U14846 (N_14846,N_12717,N_13268);
nand U14847 (N_14847,N_13223,N_12225);
nor U14848 (N_14848,N_13126,N_13284);
nand U14849 (N_14849,N_13368,N_13432);
nor U14850 (N_14850,N_12532,N_12262);
and U14851 (N_14851,N_12306,N_13287);
nor U14852 (N_14852,N_12959,N_12443);
and U14853 (N_14853,N_12001,N_13336);
xnor U14854 (N_14854,N_12824,N_13286);
and U14855 (N_14855,N_13047,N_12229);
or U14856 (N_14856,N_13486,N_13204);
nor U14857 (N_14857,N_13378,N_12698);
nor U14858 (N_14858,N_12105,N_12620);
or U14859 (N_14859,N_13287,N_13152);
nor U14860 (N_14860,N_12044,N_12466);
nor U14861 (N_14861,N_13067,N_12008);
and U14862 (N_14862,N_12411,N_13013);
and U14863 (N_14863,N_13147,N_12370);
nand U14864 (N_14864,N_12550,N_12323);
or U14865 (N_14865,N_12443,N_13152);
xor U14866 (N_14866,N_13124,N_12628);
nand U14867 (N_14867,N_13292,N_12810);
xor U14868 (N_14868,N_12472,N_12436);
and U14869 (N_14869,N_13367,N_12822);
nand U14870 (N_14870,N_13181,N_13496);
and U14871 (N_14871,N_13020,N_13166);
or U14872 (N_14872,N_12532,N_12392);
and U14873 (N_14873,N_13171,N_13437);
nand U14874 (N_14874,N_13217,N_12304);
nor U14875 (N_14875,N_12129,N_12689);
nor U14876 (N_14876,N_13159,N_12188);
nand U14877 (N_14877,N_13120,N_13499);
nand U14878 (N_14878,N_12147,N_12239);
xnor U14879 (N_14879,N_13061,N_13432);
nand U14880 (N_14880,N_12815,N_12457);
and U14881 (N_14881,N_13338,N_13045);
or U14882 (N_14882,N_13287,N_12768);
or U14883 (N_14883,N_12526,N_12217);
nor U14884 (N_14884,N_12297,N_12132);
and U14885 (N_14885,N_13290,N_12621);
or U14886 (N_14886,N_12946,N_13465);
or U14887 (N_14887,N_12042,N_12831);
or U14888 (N_14888,N_12104,N_12820);
nor U14889 (N_14889,N_12872,N_13470);
nand U14890 (N_14890,N_13215,N_12415);
and U14891 (N_14891,N_12038,N_13372);
xor U14892 (N_14892,N_13069,N_12344);
nand U14893 (N_14893,N_13382,N_13496);
xnor U14894 (N_14894,N_12300,N_12734);
nor U14895 (N_14895,N_13188,N_13118);
xnor U14896 (N_14896,N_13028,N_12024);
or U14897 (N_14897,N_13390,N_12181);
nand U14898 (N_14898,N_13127,N_12789);
or U14899 (N_14899,N_12213,N_13318);
and U14900 (N_14900,N_13239,N_12763);
nand U14901 (N_14901,N_12610,N_13207);
and U14902 (N_14902,N_12209,N_13469);
nand U14903 (N_14903,N_13076,N_13349);
nand U14904 (N_14904,N_12318,N_12697);
xnor U14905 (N_14905,N_12901,N_13473);
xnor U14906 (N_14906,N_12449,N_12151);
nor U14907 (N_14907,N_13057,N_13458);
nor U14908 (N_14908,N_13308,N_12413);
nand U14909 (N_14909,N_12110,N_13089);
and U14910 (N_14910,N_12364,N_12819);
nand U14911 (N_14911,N_12920,N_12411);
nor U14912 (N_14912,N_12585,N_12233);
xnor U14913 (N_14913,N_13088,N_12415);
and U14914 (N_14914,N_12030,N_13463);
and U14915 (N_14915,N_12800,N_12944);
or U14916 (N_14916,N_13351,N_13248);
or U14917 (N_14917,N_13327,N_12518);
xor U14918 (N_14918,N_13269,N_12387);
or U14919 (N_14919,N_12032,N_13162);
nand U14920 (N_14920,N_12706,N_12497);
and U14921 (N_14921,N_12272,N_12863);
xor U14922 (N_14922,N_13095,N_12463);
and U14923 (N_14923,N_13275,N_12985);
or U14924 (N_14924,N_12427,N_13010);
nor U14925 (N_14925,N_12365,N_12538);
or U14926 (N_14926,N_13311,N_12421);
and U14927 (N_14927,N_12525,N_12923);
or U14928 (N_14928,N_12674,N_12443);
or U14929 (N_14929,N_12626,N_13009);
or U14930 (N_14930,N_13338,N_12026);
xnor U14931 (N_14931,N_12979,N_13245);
or U14932 (N_14932,N_12206,N_12302);
and U14933 (N_14933,N_12203,N_13018);
and U14934 (N_14934,N_13259,N_12557);
nand U14935 (N_14935,N_12655,N_12585);
or U14936 (N_14936,N_13044,N_13234);
nand U14937 (N_14937,N_12991,N_12799);
or U14938 (N_14938,N_12089,N_12343);
xnor U14939 (N_14939,N_12223,N_12280);
nand U14940 (N_14940,N_12200,N_13464);
or U14941 (N_14941,N_12558,N_13242);
nand U14942 (N_14942,N_12206,N_12022);
and U14943 (N_14943,N_13208,N_12546);
and U14944 (N_14944,N_12988,N_12450);
or U14945 (N_14945,N_13011,N_12587);
or U14946 (N_14946,N_12125,N_13014);
or U14947 (N_14947,N_12371,N_12737);
and U14948 (N_14948,N_12984,N_12538);
and U14949 (N_14949,N_12341,N_12267);
and U14950 (N_14950,N_12575,N_12288);
nor U14951 (N_14951,N_12055,N_12078);
nor U14952 (N_14952,N_12140,N_12395);
nand U14953 (N_14953,N_13264,N_12602);
or U14954 (N_14954,N_12594,N_13218);
nand U14955 (N_14955,N_12123,N_12567);
nor U14956 (N_14956,N_12079,N_13146);
and U14957 (N_14957,N_12491,N_12489);
xor U14958 (N_14958,N_13186,N_12330);
xor U14959 (N_14959,N_12704,N_12372);
xnor U14960 (N_14960,N_12411,N_12113);
xor U14961 (N_14961,N_12283,N_13204);
nor U14962 (N_14962,N_13208,N_13263);
nand U14963 (N_14963,N_12369,N_13110);
xnor U14964 (N_14964,N_12305,N_12545);
or U14965 (N_14965,N_13287,N_13290);
nor U14966 (N_14966,N_12455,N_12884);
xor U14967 (N_14967,N_13025,N_12359);
or U14968 (N_14968,N_13010,N_13249);
xor U14969 (N_14969,N_12930,N_13340);
nor U14970 (N_14970,N_13037,N_13004);
or U14971 (N_14971,N_13041,N_12557);
xnor U14972 (N_14972,N_12485,N_12628);
and U14973 (N_14973,N_12366,N_12355);
nand U14974 (N_14974,N_12535,N_12977);
or U14975 (N_14975,N_13266,N_13164);
and U14976 (N_14976,N_12248,N_12099);
xor U14977 (N_14977,N_13196,N_12798);
nor U14978 (N_14978,N_13273,N_13380);
xor U14979 (N_14979,N_12013,N_13107);
or U14980 (N_14980,N_12976,N_12128);
nor U14981 (N_14981,N_13199,N_12242);
nand U14982 (N_14982,N_12656,N_12378);
xor U14983 (N_14983,N_13299,N_13283);
nor U14984 (N_14984,N_12390,N_12407);
nand U14985 (N_14985,N_12695,N_13068);
and U14986 (N_14986,N_12772,N_13167);
xnor U14987 (N_14987,N_12717,N_12618);
xnor U14988 (N_14988,N_12466,N_12581);
nor U14989 (N_14989,N_12541,N_13156);
nand U14990 (N_14990,N_12512,N_12801);
nor U14991 (N_14991,N_13381,N_12226);
nor U14992 (N_14992,N_13488,N_12270);
or U14993 (N_14993,N_12596,N_12609);
nor U14994 (N_14994,N_12050,N_12520);
nand U14995 (N_14995,N_12125,N_12910);
nand U14996 (N_14996,N_12218,N_12305);
and U14997 (N_14997,N_12749,N_13262);
and U14998 (N_14998,N_13317,N_13134);
xor U14999 (N_14999,N_12107,N_12043);
nor U15000 (N_15000,N_13681,N_13980);
nand U15001 (N_15001,N_13539,N_14737);
nor U15002 (N_15002,N_14947,N_14932);
xor U15003 (N_15003,N_13618,N_14227);
nor U15004 (N_15004,N_14255,N_14538);
or U15005 (N_15005,N_14346,N_14467);
nand U15006 (N_15006,N_14708,N_14589);
and U15007 (N_15007,N_14850,N_14048);
xnor U15008 (N_15008,N_14211,N_13550);
xor U15009 (N_15009,N_14221,N_13714);
and U15010 (N_15010,N_14109,N_13928);
and U15011 (N_15011,N_13802,N_14067);
nor U15012 (N_15012,N_14481,N_14466);
nand U15013 (N_15013,N_14974,N_14855);
xor U15014 (N_15014,N_14331,N_13638);
or U15015 (N_15015,N_14123,N_14229);
or U15016 (N_15016,N_14875,N_13865);
nand U15017 (N_15017,N_14012,N_14925);
nand U15018 (N_15018,N_14540,N_14282);
nand U15019 (N_15019,N_14535,N_13741);
xor U15020 (N_15020,N_14070,N_14408);
nand U15021 (N_15021,N_14018,N_14715);
or U15022 (N_15022,N_14185,N_14507);
xor U15023 (N_15023,N_14370,N_14645);
or U15024 (N_15024,N_14004,N_14399);
xnor U15025 (N_15025,N_13876,N_14612);
nand U15026 (N_15026,N_13705,N_14834);
or U15027 (N_15027,N_13636,N_14684);
and U15028 (N_15028,N_14972,N_14877);
xnor U15029 (N_15029,N_14874,N_14059);
nor U15030 (N_15030,N_14889,N_14967);
nor U15031 (N_15031,N_14144,N_14456);
nor U15032 (N_15032,N_13855,N_13576);
xor U15033 (N_15033,N_14147,N_14579);
nor U15034 (N_15034,N_14573,N_14624);
nor U15035 (N_15035,N_13611,N_13505);
nand U15036 (N_15036,N_13686,N_13597);
or U15037 (N_15037,N_14117,N_14712);
or U15038 (N_15038,N_14438,N_14750);
and U15039 (N_15039,N_14561,N_14701);
and U15040 (N_15040,N_14280,N_13748);
and U15041 (N_15041,N_14388,N_14598);
xor U15042 (N_15042,N_14577,N_14631);
and U15043 (N_15043,N_14361,N_13557);
nand U15044 (N_15044,N_14541,N_14544);
nor U15045 (N_15045,N_14494,N_13879);
xnor U15046 (N_15046,N_14909,N_14757);
and U15047 (N_15047,N_14262,N_14093);
nor U15048 (N_15048,N_13946,N_13915);
and U15049 (N_15049,N_14851,N_13640);
and U15050 (N_15050,N_13944,N_14263);
and U15051 (N_15051,N_14574,N_13656);
and U15052 (N_15052,N_14417,N_13782);
xnor U15053 (N_15053,N_14862,N_14790);
nor U15054 (N_15054,N_14818,N_14375);
nor U15055 (N_15055,N_13588,N_14349);
xor U15056 (N_15056,N_13767,N_13892);
and U15057 (N_15057,N_14509,N_14813);
and U15058 (N_15058,N_14977,N_14114);
nor U15059 (N_15059,N_14521,N_14023);
or U15060 (N_15060,N_13589,N_13911);
and U15061 (N_15061,N_14901,N_14415);
xor U15062 (N_15062,N_13540,N_13533);
xnor U15063 (N_15063,N_13757,N_13871);
nor U15064 (N_15064,N_14188,N_14215);
or U15065 (N_15065,N_13961,N_14040);
nand U15066 (N_15066,N_13722,N_13524);
xor U15067 (N_15067,N_14213,N_14697);
or U15068 (N_15068,N_14127,N_13942);
or U15069 (N_15069,N_14333,N_13937);
or U15070 (N_15070,N_14665,N_13662);
nor U15071 (N_15071,N_13695,N_13858);
or U15072 (N_15072,N_14603,N_14582);
and U15073 (N_15073,N_13659,N_14195);
nand U15074 (N_15074,N_13812,N_14892);
nand U15075 (N_15075,N_13771,N_14590);
xor U15076 (N_15076,N_13828,N_14395);
nand U15077 (N_15077,N_14209,N_14578);
nor U15078 (N_15078,N_14196,N_14869);
nand U15079 (N_15079,N_13700,N_13545);
nand U15080 (N_15080,N_14134,N_13793);
xnor U15081 (N_15081,N_14774,N_13926);
nor U15082 (N_15082,N_14105,N_13718);
or U15083 (N_15083,N_13956,N_14106);
and U15084 (N_15084,N_14381,N_13668);
nor U15085 (N_15085,N_13500,N_14452);
nor U15086 (N_15086,N_13848,N_13507);
nor U15087 (N_15087,N_13555,N_13979);
nor U15088 (N_15088,N_14946,N_14672);
nand U15089 (N_15089,N_13822,N_13606);
xor U15090 (N_15090,N_14557,N_13627);
xor U15091 (N_15091,N_14652,N_13970);
nand U15092 (N_15092,N_13586,N_14170);
nor U15093 (N_15093,N_14091,N_14780);
or U15094 (N_15094,N_13584,N_13963);
and U15095 (N_15095,N_13610,N_14725);
xnor U15096 (N_15096,N_14576,N_13951);
and U15097 (N_15097,N_14896,N_14938);
and U15098 (N_15098,N_13508,N_13502);
nand U15099 (N_15099,N_14998,N_13836);
xor U15100 (N_15100,N_14788,N_14753);
or U15101 (N_15101,N_14128,N_14219);
nor U15102 (N_15102,N_14823,N_14001);
nor U15103 (N_15103,N_14228,N_14250);
nand U15104 (N_15104,N_14198,N_13780);
nor U15105 (N_15105,N_14657,N_14824);
xor U15106 (N_15106,N_14762,N_13805);
xor U15107 (N_15107,N_14190,N_14667);
and U15108 (N_15108,N_13845,N_13725);
nand U15109 (N_15109,N_13929,N_14181);
xnor U15110 (N_15110,N_14880,N_14898);
nor U15111 (N_15111,N_13740,N_14251);
and U15112 (N_15112,N_14843,N_13752);
nor U15113 (N_15113,N_13719,N_14095);
and U15114 (N_15114,N_14794,N_13582);
xor U15115 (N_15115,N_14118,N_14024);
and U15116 (N_15116,N_14107,N_13632);
nand U15117 (N_15117,N_14944,N_13934);
nand U15118 (N_15118,N_14642,N_14427);
and U15119 (N_15119,N_14656,N_14845);
nor U15120 (N_15120,N_14635,N_13673);
xnor U15121 (N_15121,N_14797,N_13666);
and U15122 (N_15122,N_14044,N_14055);
and U15123 (N_15123,N_13885,N_14513);
xnor U15124 (N_15124,N_13893,N_14177);
and U15125 (N_15125,N_14063,N_14277);
and U15126 (N_15126,N_13736,N_14311);
or U15127 (N_15127,N_14424,N_13841);
nor U15128 (N_15128,N_14945,N_13528);
and U15129 (N_15129,N_13578,N_14168);
and U15130 (N_15130,N_14274,N_14726);
xnor U15131 (N_15131,N_14478,N_13676);
nor U15132 (N_15132,N_14766,N_13823);
nand U15133 (N_15133,N_14416,N_13663);
xnor U15134 (N_15134,N_13515,N_13954);
xnor U15135 (N_15135,N_14747,N_13900);
xor U15136 (N_15136,N_14300,N_13850);
nand U15137 (N_15137,N_14137,N_13563);
and U15138 (N_15138,N_14542,N_14252);
and U15139 (N_15139,N_14899,N_14143);
xor U15140 (N_15140,N_14917,N_14992);
nand U15141 (N_15141,N_14453,N_13800);
and U15142 (N_15142,N_14679,N_14524);
and U15143 (N_15143,N_14525,N_13623);
nand U15144 (N_15144,N_13992,N_14296);
and U15145 (N_15145,N_13818,N_13556);
xnor U15146 (N_15146,N_14306,N_13947);
nand U15147 (N_15147,N_14508,N_14621);
nand U15148 (N_15148,N_14192,N_14298);
and U15149 (N_15149,N_14826,N_13962);
or U15150 (N_15150,N_14391,N_14791);
or U15151 (N_15151,N_14622,N_13733);
nand U15152 (N_15152,N_14247,N_13587);
nor U15153 (N_15153,N_14108,N_14694);
nand U15154 (N_15154,N_14552,N_13868);
and U15155 (N_15155,N_13669,N_13605);
xnor U15156 (N_15156,N_14058,N_13753);
nand U15157 (N_15157,N_14020,N_13581);
and U15158 (N_15158,N_14911,N_14152);
and U15159 (N_15159,N_14328,N_14888);
or U15160 (N_15160,N_14455,N_13774);
or U15161 (N_15161,N_14283,N_14640);
or U15162 (N_15162,N_14003,N_13991);
or U15163 (N_15163,N_14086,N_14618);
xor U15164 (N_15164,N_14596,N_14324);
xnor U15165 (N_15165,N_13595,N_14373);
or U15166 (N_15166,N_14162,N_14581);
or U15167 (N_15167,N_14560,N_14802);
nand U15168 (N_15168,N_14459,N_13861);
and U15169 (N_15169,N_14770,N_14394);
or U15170 (N_15170,N_14239,N_14852);
nor U15171 (N_15171,N_13715,N_13621);
xnor U15172 (N_15172,N_14704,N_14563);
nor U15173 (N_15173,N_14611,N_13760);
xnor U15174 (N_15174,N_14476,N_13960);
nand U15175 (N_15175,N_13974,N_13849);
nand U15176 (N_15176,N_14685,N_14900);
nand U15177 (N_15177,N_14189,N_14369);
or U15178 (N_15178,N_14545,N_14342);
nor U15179 (N_15179,N_13699,N_14919);
xnor U15180 (N_15180,N_14376,N_13986);
or U15181 (N_15181,N_14831,N_13620);
nor U15182 (N_15182,N_13927,N_14918);
nor U15183 (N_15183,N_13862,N_14275);
nand U15184 (N_15184,N_14949,N_14721);
and U15185 (N_15185,N_14960,N_14829);
and U15186 (N_15186,N_14015,N_14210);
and U15187 (N_15187,N_14191,N_14692);
nor U15188 (N_15188,N_14014,N_14223);
xor U15189 (N_15189,N_13955,N_14953);
nor U15190 (N_15190,N_14073,N_14744);
or U15191 (N_15191,N_14301,N_14194);
nor U15192 (N_15192,N_14339,N_14758);
xnor U15193 (N_15193,N_13664,N_13631);
nor U15194 (N_15194,N_13526,N_14430);
or U15195 (N_15195,N_14366,N_14979);
or U15196 (N_15196,N_14693,N_14419);
nand U15197 (N_15197,N_14836,N_14350);
xor U15198 (N_15198,N_14396,N_13895);
and U15199 (N_15199,N_13814,N_14288);
or U15200 (N_15200,N_13626,N_14230);
nand U15201 (N_15201,N_14519,N_13854);
or U15202 (N_15202,N_14668,N_13878);
nand U15203 (N_15203,N_14835,N_13792);
nor U15204 (N_15204,N_14341,N_13815);
or U15205 (N_15205,N_13601,N_14547);
nor U15206 (N_15206,N_13938,N_14516);
and U15207 (N_15207,N_14775,N_14759);
xnor U15208 (N_15208,N_14013,N_13711);
and U15209 (N_15209,N_13797,N_14987);
xor U15210 (N_15210,N_14546,N_13710);
nor U15211 (N_15211,N_14327,N_14962);
or U15212 (N_15212,N_13616,N_14201);
nor U15213 (N_15213,N_14060,N_14098);
nor U15214 (N_15214,N_14085,N_13688);
and U15215 (N_15215,N_14727,N_14267);
and U15216 (N_15216,N_14240,N_14308);
and U15217 (N_15217,N_14153,N_14043);
and U15218 (N_15218,N_14202,N_13981);
nor U15219 (N_15219,N_14890,N_14047);
or U15220 (N_15220,N_13651,N_13971);
xor U15221 (N_15221,N_14928,N_14450);
xor U15222 (N_15222,N_13503,N_14854);
or U15223 (N_15223,N_13590,N_14902);
or U15224 (N_15224,N_13566,N_14315);
xnor U15225 (N_15225,N_14723,N_13930);
and U15226 (N_15226,N_14604,N_13901);
xnor U15227 (N_15227,N_13872,N_13564);
nor U15228 (N_15228,N_13541,N_14066);
nand U15229 (N_15229,N_14207,N_13851);
or U15230 (N_15230,N_13567,N_13965);
and U15231 (N_15231,N_13538,N_14236);
and U15232 (N_15232,N_13553,N_13645);
nor U15233 (N_15233,N_14859,N_13987);
nor U15234 (N_15234,N_14752,N_13637);
nand U15235 (N_15235,N_14666,N_13770);
nor U15236 (N_15236,N_14748,N_14895);
nor U15237 (N_15237,N_14076,N_14053);
nand U15238 (N_15238,N_13609,N_14532);
nor U15239 (N_15239,N_14506,N_13830);
and U15240 (N_15240,N_13953,N_13698);
xnor U15241 (N_15241,N_14479,N_14092);
and U15242 (N_15242,N_13537,N_13561);
xor U15243 (N_15243,N_14312,N_14504);
nand U15244 (N_15244,N_14115,N_13795);
nor U15245 (N_15245,N_13808,N_14517);
nand U15246 (N_15246,N_13964,N_13829);
xnor U15247 (N_15247,N_13819,N_14695);
nand U15248 (N_15248,N_14908,N_14523);
nor U15249 (N_15249,N_14781,N_13520);
or U15250 (N_15250,N_14054,N_14100);
nor U15251 (N_15251,N_14110,N_14833);
xor U15252 (N_15252,N_13650,N_14608);
xnor U15253 (N_15253,N_13614,N_14539);
xnor U15254 (N_15254,N_14332,N_13667);
xnor U15255 (N_15255,N_14320,N_13510);
and U15256 (N_15256,N_14353,N_14948);
xor U15257 (N_15257,N_14606,N_14097);
xnor U15258 (N_15258,N_13677,N_14585);
xnor U15259 (N_15259,N_13863,N_13794);
or U15260 (N_15260,N_13891,N_14437);
nand U15261 (N_15261,N_14584,N_14907);
or U15262 (N_15262,N_14005,N_13912);
and U15263 (N_15263,N_14351,N_14597);
and U15264 (N_15264,N_14849,N_14713);
nand U15265 (N_15265,N_14261,N_14449);
xor U15266 (N_15266,N_14290,N_14903);
xnor U15267 (N_15267,N_14498,N_13720);
xnor U15268 (N_15268,N_14683,N_14646);
nor U15269 (N_15269,N_14374,N_14122);
nand U15270 (N_15270,N_13785,N_14322);
nor U15271 (N_15271,N_14310,N_14730);
xor U15272 (N_15272,N_14434,N_14971);
nor U15273 (N_15273,N_13775,N_13995);
or U15274 (N_15274,N_14555,N_14873);
and U15275 (N_15275,N_14864,N_14527);
xnor U15276 (N_15276,N_13966,N_14964);
nand U15277 (N_15277,N_14980,N_14359);
and U15278 (N_15278,N_14993,N_14777);
nor U15279 (N_15279,N_14378,N_14135);
xor U15280 (N_15280,N_13717,N_14988);
and U15281 (N_15281,N_14736,N_14812);
nor U15282 (N_15282,N_14627,N_14626);
and U15283 (N_15283,N_14056,N_13916);
and U15284 (N_15284,N_13798,N_14075);
nand U15285 (N_15285,N_14138,N_13534);
xnor U15286 (N_15286,N_14814,N_13525);
xnor U15287 (N_15287,N_14879,N_13535);
and U15288 (N_15288,N_13596,N_13709);
xnor U15289 (N_15289,N_13747,N_13531);
xor U15290 (N_15290,N_13511,N_14386);
or U15291 (N_15291,N_13936,N_13920);
or U15292 (N_15292,N_14287,N_13873);
or U15293 (N_15293,N_14077,N_14232);
xnor U15294 (N_15294,N_14856,N_13904);
xor U15295 (N_15295,N_13765,N_14245);
nor U15296 (N_15296,N_14404,N_13952);
xor U15297 (N_15297,N_14179,N_13516);
or U15298 (N_15298,N_14203,N_13749);
or U15299 (N_15299,N_14472,N_14981);
nor U15300 (N_15300,N_14528,N_13514);
nand U15301 (N_15301,N_13660,N_14676);
or U15302 (N_15302,N_13923,N_13641);
and U15303 (N_15303,N_13925,N_14164);
nor U15304 (N_15304,N_14489,N_14382);
nor U15305 (N_15305,N_13746,N_14458);
and U15306 (N_15306,N_14397,N_14571);
and U15307 (N_15307,N_13630,N_13592);
xor U15308 (N_15308,N_14924,N_14772);
and U15309 (N_15309,N_13504,N_14664);
or U15310 (N_15310,N_14619,N_14488);
and U15311 (N_15311,N_13788,N_14062);
or U15312 (N_15312,N_13512,N_14436);
and U15313 (N_15313,N_14763,N_14033);
xor U15314 (N_15314,N_14083,N_14749);
nor U15315 (N_15315,N_13523,N_13560);
nand U15316 (N_15316,N_13517,N_14553);
and U15317 (N_15317,N_13552,N_14068);
and U15318 (N_15318,N_13682,N_13776);
or U15319 (N_15319,N_13976,N_13820);
nand U15320 (N_15320,N_14496,N_14099);
xor U15321 (N_15321,N_14484,N_13513);
nor U15322 (N_15322,N_13789,N_14658);
xor U15323 (N_15323,N_14216,N_14660);
nand U15324 (N_15324,N_14805,N_14103);
and U15325 (N_15325,N_13727,N_14559);
nand U15326 (N_15326,N_14238,N_14973);
and U15327 (N_15327,N_13607,N_14041);
nand U15328 (N_15328,N_13799,N_14937);
xor U15329 (N_15329,N_14079,N_14268);
nor U15330 (N_15330,N_14113,N_14171);
xor U15331 (N_15331,N_13622,N_14817);
nor U15332 (N_15332,N_14139,N_13737);
nor U15333 (N_15333,N_13968,N_14398);
xor U15334 (N_15334,N_14187,N_13728);
nor U15335 (N_15335,N_14549,N_14620);
xor U15336 (N_15336,N_14451,N_13832);
and U15337 (N_15337,N_14554,N_14088);
nor U15338 (N_15338,N_14357,N_14858);
and U15339 (N_15339,N_13721,N_14614);
and U15340 (N_15340,N_14910,N_14687);
nand U15341 (N_15341,N_14989,N_13731);
nand U15342 (N_15342,N_14038,N_14926);
or U15343 (N_15343,N_14299,N_14564);
nand U15344 (N_15344,N_13957,N_14678);
xnor U15345 (N_15345,N_14916,N_13687);
and U15346 (N_15346,N_14051,N_14231);
or U15347 (N_15347,N_13781,N_13977);
and U15348 (N_15348,N_13672,N_13568);
nor U15349 (N_15349,N_14305,N_14343);
and U15350 (N_15350,N_14368,N_13671);
nand U15351 (N_15351,N_13867,N_14445);
and U15352 (N_15352,N_14030,N_14371);
and U15353 (N_15353,N_14625,N_13969);
nand U15354 (N_15354,N_14384,N_13763);
xnor U15355 (N_15355,N_14444,N_13978);
nor U15356 (N_15356,N_14273,N_14487);
nand U15357 (N_15357,N_13522,N_14154);
or U15358 (N_15358,N_14933,N_14126);
or U15359 (N_15359,N_13690,N_14161);
or U15360 (N_15360,N_14429,N_14957);
nand U15361 (N_15361,N_13880,N_13577);
xnor U15362 (N_15362,N_14601,N_14428);
nand U15363 (N_15363,N_13870,N_14821);
nor U15364 (N_15364,N_14362,N_13844);
and U15365 (N_15365,N_14848,N_14112);
xor U15366 (N_15366,N_14222,N_13565);
and U15367 (N_15367,N_13674,N_14206);
and U15368 (N_15368,N_14515,N_14026);
or U15369 (N_15369,N_14629,N_14008);
nor U15370 (N_15370,N_14832,N_14257);
nor U15371 (N_15371,N_14183,N_14609);
nor U15372 (N_15372,N_14558,N_14355);
nor U15373 (N_15373,N_13835,N_14286);
and U15374 (N_15374,N_13602,N_13807);
nand U15375 (N_15375,N_14591,N_14639);
xnor U15376 (N_15376,N_14304,N_14820);
xnor U15377 (N_15377,N_14876,N_14411);
or U15378 (N_15378,N_14878,N_13875);
nor U15379 (N_15379,N_14995,N_14931);
or U15380 (N_15380,N_14580,N_14413);
and U15381 (N_15381,N_13745,N_14968);
nand U15382 (N_15382,N_14819,N_14292);
and U15383 (N_15383,N_14491,N_14363);
and U15384 (N_15384,N_14344,N_14439);
nand U15385 (N_15385,N_14000,N_14148);
xnor U15386 (N_15386,N_13608,N_14991);
or U15387 (N_15387,N_13772,N_13903);
nor U15388 (N_15388,N_14199,N_14754);
or U15389 (N_15389,N_14724,N_14474);
and U15390 (N_15390,N_14769,N_14501);
and U15391 (N_15391,N_13833,N_14248);
and U15392 (N_15392,N_14915,N_13519);
or U15393 (N_15393,N_14675,N_14731);
xnor U15394 (N_15394,N_14745,N_13856);
nor U15395 (N_15395,N_14922,N_14284);
nor U15396 (N_15396,N_13993,N_14499);
and U15397 (N_15397,N_14461,N_13532);
nand U15398 (N_15398,N_14052,N_14798);
or U15399 (N_15399,N_13834,N_14688);
xor U15400 (N_15400,N_14101,N_14208);
nand U15401 (N_15401,N_13629,N_14125);
and U15402 (N_15402,N_13890,N_14010);
xnor U15403 (N_15403,N_14080,N_14816);
nand U15404 (N_15404,N_14096,N_14756);
xor U15405 (N_15405,N_14297,N_14218);
nand U15406 (N_15406,N_14163,N_14323);
and U15407 (N_15407,N_13777,N_14418);
xnor U15408 (N_15408,N_14421,N_14380);
or U15409 (N_15409,N_14716,N_14969);
or U15410 (N_15410,N_13612,N_14807);
or U15411 (N_15411,N_14550,N_14032);
or U15412 (N_15412,N_14356,N_13999);
and U15413 (N_15413,N_13827,N_14914);
nand U15414 (N_15414,N_14881,N_13933);
nand U15415 (N_15415,N_14243,N_13898);
xor U15416 (N_15416,N_13683,N_13922);
or U15417 (N_15417,N_14764,N_14242);
nand U15418 (N_15418,N_14970,N_14885);
or U15419 (N_15419,N_13661,N_13647);
or U15420 (N_15420,N_14568,N_14983);
or U15421 (N_15421,N_13983,N_13949);
and U15422 (N_15422,N_13591,N_14326);
nand U15423 (N_15423,N_14039,N_14706);
and U15424 (N_15424,N_14628,N_14317);
xnor U15425 (N_15425,N_14490,N_14178);
nor U15426 (N_15426,N_14784,N_14468);
or U15427 (N_15427,N_14462,N_14844);
nand U15428 (N_15428,N_14266,N_13558);
nand U15429 (N_15429,N_14803,N_14906);
and U15430 (N_15430,N_14840,N_14119);
xnor U15431 (N_15431,N_13910,N_13551);
nand U15432 (N_15432,N_14662,N_14533);
nor U15433 (N_15433,N_14169,N_14699);
nand U15434 (N_15434,N_14565,N_13542);
or U15435 (N_15435,N_13544,N_14160);
and U15436 (N_15436,N_14482,N_14965);
or U15437 (N_15437,N_14259,N_14529);
xor U15438 (N_15438,N_14984,N_14702);
or U15439 (N_15439,N_14082,N_13973);
or U15440 (N_15440,N_14016,N_14246);
nand U15441 (N_15441,N_14904,N_13701);
nand U15442 (N_15442,N_14718,N_14632);
nand U15443 (N_15443,N_14336,N_14330);
xor U15444 (N_15444,N_14566,N_14289);
xor U15445 (N_15445,N_14714,N_14689);
or U15446 (N_15446,N_14682,N_14929);
and U15447 (N_15447,N_14800,N_14511);
nand U15448 (N_15448,N_14838,N_13989);
xor U15449 (N_15449,N_14174,N_13562);
xnor U15450 (N_15450,N_14959,N_13806);
nor U15451 (N_15451,N_14383,N_13600);
xnor U15452 (N_15452,N_14593,N_14167);
or U15453 (N_15453,N_14432,N_14575);
and U15454 (N_15454,N_14649,N_14985);
and U15455 (N_15455,N_14409,N_14806);
and U15456 (N_15456,N_14037,N_14711);
nand U15457 (N_15457,N_14433,N_14661);
xnor U15458 (N_15458,N_13702,N_14182);
xnor U15459 (N_15459,N_14670,N_13658);
nor U15460 (N_15460,N_14279,N_14815);
nand U15461 (N_15461,N_14943,N_14912);
nand U15462 (N_15462,N_14217,N_14503);
nor U15463 (N_15463,N_13604,N_14340);
xor U15464 (N_15464,N_14145,N_13639);
nand U15465 (N_15465,N_14440,N_14707);
xnor U15466 (N_15466,N_14522,N_14810);
nor U15467 (N_15467,N_14636,N_14265);
and U15468 (N_15468,N_14734,N_13583);
and U15469 (N_15469,N_14905,N_13678);
nor U15470 (N_15470,N_14994,N_13693);
xnor U15471 (N_15471,N_14827,N_14084);
or U15472 (N_15472,N_13670,N_14367);
or U15473 (N_15473,N_13762,N_14460);
nand U15474 (N_15474,N_13972,N_14607);
and U15475 (N_15475,N_14870,N_13824);
xor U15476 (N_15476,N_14738,N_13644);
xor U15477 (N_15477,N_14307,N_14285);
nor U15478 (N_15478,N_14473,N_14935);
xor U15479 (N_15479,N_14021,N_14868);
nor U15480 (N_15480,N_14785,N_14673);
nor U15481 (N_15481,N_13685,N_13665);
nand U15482 (N_15482,N_14654,N_14761);
and U15483 (N_15483,N_13732,N_14294);
xor U15484 (N_15484,N_14743,N_14321);
xnor U15485 (N_15485,N_13804,N_13821);
nor U15486 (N_15486,N_14543,N_14886);
nor U15487 (N_15487,N_14132,N_13724);
nand U15488 (N_15488,N_14927,N_13735);
xor U15489 (N_15489,N_13931,N_14334);
xor U15490 (N_15490,N_14111,N_14776);
nand U15491 (N_15491,N_14235,N_14677);
or U15492 (N_15492,N_14955,N_14587);
and U15493 (N_15493,N_14930,N_13939);
or U15494 (N_15494,N_14782,N_13837);
xnor U15495 (N_15495,N_13887,N_13905);
nand U15496 (N_15496,N_14615,N_14028);
nor U15497 (N_15497,N_13593,N_14244);
nor U15498 (N_15498,N_14387,N_14042);
xnor U15499 (N_15499,N_14027,N_14090);
nand U15500 (N_15500,N_13874,N_13759);
nor U15501 (N_15501,N_13619,N_13743);
or U15502 (N_15502,N_14830,N_14205);
xnor U15503 (N_15503,N_14303,N_13575);
or U15504 (N_15504,N_14651,N_13860);
or U15505 (N_15505,N_13791,N_13758);
nand U15506 (N_15506,N_14441,N_14865);
and U15507 (N_15507,N_14271,N_14595);
nand U15508 (N_15508,N_13945,N_14493);
and U15509 (N_15509,N_13884,N_13739);
nand U15510 (N_15510,N_14939,N_14999);
nand U15511 (N_15511,N_14839,N_13691);
nor U15512 (N_15512,N_13751,N_14081);
nor U15513 (N_15513,N_14325,N_14696);
xnor U15514 (N_15514,N_14087,N_14200);
nor U15515 (N_15515,N_13543,N_14345);
xor U15516 (N_15516,N_14887,N_14061);
xnor U15517 (N_15517,N_14069,N_14226);
xnor U15518 (N_15518,N_14422,N_14377);
xor U15519 (N_15519,N_14124,N_14495);
or U15520 (N_15520,N_14773,N_14669);
nand U15521 (N_15521,N_14882,N_14913);
or U15522 (N_15522,N_14318,N_13883);
and U15523 (N_15523,N_14347,N_14709);
nand U15524 (N_15524,N_13646,N_13997);
or U15525 (N_15525,N_14260,N_14588);
or U15526 (N_15526,N_14986,N_14863);
nand U15527 (N_15527,N_14337,N_14884);
nand U15528 (N_15528,N_13959,N_13831);
nor U15529 (N_15529,N_14225,N_13574);
and U15530 (N_15530,N_14364,N_14956);
nor U15531 (N_15531,N_13642,N_14583);
and U15532 (N_15532,N_14897,N_14936);
nor U15533 (N_15533,N_14760,N_14505);
or U15534 (N_15534,N_14893,N_14644);
nand U15535 (N_15535,N_14329,N_13572);
nor U15536 (N_15536,N_13509,N_14613);
or U15537 (N_15537,N_14746,N_14022);
nor U15538 (N_15538,N_14141,N_14463);
or U15539 (N_15539,N_13899,N_14094);
xor U15540 (N_15540,N_14809,N_13810);
and U15541 (N_15541,N_14634,N_13706);
or U15542 (N_15542,N_14050,N_14007);
or U15543 (N_15543,N_13917,N_13501);
and U15544 (N_15544,N_14166,N_14133);
nand U15545 (N_15545,N_14872,N_14241);
nand U15546 (N_15546,N_14348,N_13990);
nor U15547 (N_15547,N_14372,N_13943);
or U15548 (N_15548,N_13921,N_13813);
and U15549 (N_15549,N_14686,N_14036);
nand U15550 (N_15550,N_13803,N_14569);
and U15551 (N_15551,N_14966,N_14978);
and U15552 (N_15552,N_14425,N_14006);
xnor U15553 (N_15553,N_14951,N_13756);
or U15554 (N_15554,N_13689,N_14175);
or U15555 (N_15555,N_13958,N_14172);
nand U15556 (N_15556,N_13694,N_14151);
and U15557 (N_15557,N_13679,N_14393);
or U15558 (N_15558,N_14420,N_14360);
or U15559 (N_15559,N_13529,N_14883);
nor U15560 (N_15560,N_14102,N_13847);
xor U15561 (N_15561,N_13594,N_14009);
or U15562 (N_15562,N_13643,N_13913);
nand U15563 (N_15563,N_14237,N_14698);
nand U15564 (N_15564,N_13726,N_14842);
xor U15565 (N_15565,N_14272,N_14562);
xnor U15566 (N_15566,N_14150,N_13906);
or U15567 (N_15567,N_14258,N_13579);
or U15568 (N_15568,N_14520,N_14729);
xor U15569 (N_15569,N_14963,N_14822);
nor U15570 (N_15570,N_14857,N_14548);
or U15571 (N_15571,N_14313,N_14990);
nor U15572 (N_15572,N_14861,N_14389);
and U15573 (N_15573,N_14392,N_14029);
and U15574 (N_15574,N_13696,N_13684);
or U15575 (N_15575,N_13729,N_13864);
and U15576 (N_15576,N_13712,N_14116);
xnor U15577 (N_15577,N_14405,N_14586);
nor U15578 (N_15578,N_14690,N_14401);
or U15579 (N_15579,N_14365,N_14064);
and U15580 (N_15580,N_14270,N_13839);
and U15581 (N_15581,N_13655,N_13809);
and U15582 (N_15582,N_13615,N_14847);
nand U15583 (N_15583,N_14801,N_14254);
xnor U15584 (N_15584,N_14319,N_14253);
and U15585 (N_15585,N_13530,N_14074);
nand U15586 (N_15586,N_14149,N_14120);
nor U15587 (N_15587,N_14131,N_13888);
nor U15588 (N_15588,N_13882,N_13950);
xor U15589 (N_15589,N_13549,N_13652);
nand U15590 (N_15590,N_14071,N_14142);
nor U15591 (N_15591,N_14435,N_14457);
xnor U15592 (N_15592,N_14846,N_14572);
nand U15593 (N_15593,N_14691,N_13769);
and U15594 (N_15594,N_14671,N_13897);
xor U15595 (N_15595,N_13967,N_14049);
xor U15596 (N_15596,N_13881,N_13624);
and U15597 (N_15597,N_14828,N_13518);
nand U15598 (N_15598,N_14786,N_13768);
nand U15599 (N_15599,N_13649,N_14471);
xor U15600 (N_15600,N_13536,N_14335);
or U15601 (N_15601,N_14256,N_14406);
nor U15602 (N_15602,N_13654,N_13734);
or U15603 (N_15603,N_14002,N_14853);
nand U15604 (N_15604,N_14659,N_14470);
xor U15605 (N_15605,N_14787,N_14610);
and U15606 (N_15606,N_14961,N_14423);
xor U15607 (N_15607,N_14537,N_14866);
or U15608 (N_15608,N_14276,N_14518);
nand U15609 (N_15609,N_14485,N_14278);
nand U15610 (N_15610,N_13723,N_14385);
and U15611 (N_15611,N_14647,N_13703);
nand U15612 (N_15612,N_14771,N_14155);
nor U15613 (N_15613,N_14121,N_13634);
or U15614 (N_15614,N_14510,N_14475);
or U15615 (N_15615,N_14796,N_13817);
and U15616 (N_15616,N_14078,N_14703);
nand U15617 (N_15617,N_14442,N_14212);
and U15618 (N_15618,N_14710,N_13941);
and U15619 (N_15619,N_14921,N_14269);
or U15620 (N_15620,N_14599,N_14765);
and U15621 (N_15621,N_14446,N_14176);
nor U15622 (N_15622,N_14783,N_14443);
and U15623 (N_15623,N_13559,N_13866);
nor U15624 (N_15624,N_13750,N_13996);
nor U15625 (N_15625,N_14825,N_14412);
nor U15626 (N_15626,N_14722,N_14616);
xnor U15627 (N_15627,N_13548,N_13988);
and U15628 (N_15628,N_14871,N_14600);
or U15629 (N_15629,N_14778,N_14728);
or U15630 (N_15630,N_14650,N_13816);
nand U15631 (N_15631,N_13599,N_14617);
nand U15632 (N_15632,N_13554,N_14072);
xor U15633 (N_15633,N_14338,N_13598);
or U15634 (N_15634,N_14674,N_14741);
nor U15635 (N_15635,N_13547,N_14799);
or U15636 (N_15636,N_13843,N_14638);
and U15637 (N_15637,N_14755,N_14249);
or U15638 (N_15638,N_13852,N_14046);
and U15639 (N_15639,N_14390,N_14486);
nand U15640 (N_15640,N_13783,N_13603);
nor U15641 (N_15641,N_13784,N_14808);
nand U15642 (N_15642,N_13580,N_13796);
nand U15643 (N_15643,N_13935,N_14309);
and U15644 (N_15644,N_14407,N_13902);
and U15645 (N_15645,N_14641,N_14740);
nand U15646 (N_15646,N_14789,N_13653);
or U15647 (N_15647,N_13680,N_13773);
nand U15648 (N_15648,N_14233,N_14531);
xnor U15649 (N_15649,N_13742,N_14551);
or U15650 (N_15650,N_13570,N_14792);
nand U15651 (N_15651,N_13730,N_14767);
xnor U15652 (N_15652,N_14952,N_13521);
nand U15653 (N_15653,N_14402,N_13761);
xor U15654 (N_15654,N_14065,N_13825);
nand U15655 (N_15655,N_14867,N_13811);
nand U15656 (N_15656,N_14136,N_13984);
or U15657 (N_15657,N_14811,N_13764);
nand U15658 (N_15658,N_13675,N_14197);
xnor U15659 (N_15659,N_14431,N_14400);
nand U15660 (N_15660,N_14264,N_14454);
nand U15661 (N_15661,N_14592,N_14891);
and U15662 (N_15662,N_14941,N_14860);
nand U15663 (N_15663,N_14920,N_13975);
and U15664 (N_15664,N_13908,N_14536);
or U15665 (N_15665,N_14958,N_14224);
xor U15666 (N_15666,N_14316,N_14293);
or U15667 (N_15667,N_13924,N_14663);
or U15668 (N_15668,N_14567,N_13766);
nand U15669 (N_15669,N_14717,N_13786);
and U15670 (N_15670,N_13985,N_14295);
xnor U15671 (N_15671,N_14804,N_13909);
nor U15672 (N_15672,N_14942,N_14637);
or U15673 (N_15673,N_14950,N_14158);
or U15674 (N_15674,N_13571,N_13754);
xor U15675 (N_15675,N_14193,N_13914);
nor U15676 (N_15676,N_14602,N_13948);
xnor U15677 (N_15677,N_13869,N_14530);
nor U15678 (N_15678,N_13918,N_14732);
xor U15679 (N_15679,N_14447,N_14841);
or U15680 (N_15680,N_13744,N_14291);
xor U15681 (N_15681,N_14403,N_14534);
nand U15682 (N_15682,N_13648,N_14129);
nor U15683 (N_15683,N_14492,N_13779);
or U15684 (N_15684,N_14184,N_14173);
xor U15685 (N_15685,N_14352,N_14483);
xor U15686 (N_15686,N_13506,N_14837);
nand U15687 (N_15687,N_13613,N_14186);
xor U15688 (N_15688,N_14655,N_14426);
nor U15689 (N_15689,N_14017,N_13919);
and U15690 (N_15690,N_14220,N_13704);
nor U15691 (N_15691,N_14140,N_14104);
and U15692 (N_15692,N_13635,N_14923);
xor U15693 (N_15693,N_14733,N_13573);
or U15694 (N_15694,N_13826,N_13940);
and U15695 (N_15695,N_13907,N_14681);
nor U15696 (N_15696,N_14700,N_13853);
xnor U15697 (N_15697,N_14680,N_14630);
xnor U15698 (N_15698,N_14045,N_14997);
xor U15699 (N_15699,N_14035,N_13738);
xor U15700 (N_15700,N_14982,N_14556);
xor U15701 (N_15701,N_14204,N_13585);
nor U15702 (N_15702,N_14410,N_14464);
nand U15703 (N_15703,N_14130,N_13857);
xnor U15704 (N_15704,N_14089,N_14643);
xor U15705 (N_15705,N_14156,N_14934);
and U15706 (N_15706,N_14735,N_13707);
nand U15707 (N_15707,N_14157,N_14623);
xor U15708 (N_15708,N_14031,N_13713);
nand U15709 (N_15709,N_13617,N_13628);
nand U15710 (N_15710,N_14025,N_14469);
and U15711 (N_15711,N_14996,N_14011);
or U15712 (N_15712,N_13838,N_14705);
nor U15713 (N_15713,N_13846,N_14358);
and U15714 (N_15714,N_14180,N_14057);
and U15715 (N_15715,N_14146,N_14719);
xnor U15716 (N_15716,N_14379,N_14234);
or U15717 (N_15717,N_14894,N_13697);
nand U15718 (N_15718,N_14720,N_14512);
nand U15719 (N_15719,N_13859,N_13657);
nor U15720 (N_15720,N_14605,N_13886);
xnor U15721 (N_15721,N_14570,N_13889);
xnor U15722 (N_15722,N_14165,N_14954);
and U15723 (N_15723,N_14514,N_13877);
or U15724 (N_15724,N_13787,N_14940);
or U15725 (N_15725,N_13842,N_13527);
xnor U15726 (N_15726,N_13998,N_14975);
xor U15727 (N_15727,N_14480,N_13625);
nand U15728 (N_15728,N_13994,N_14414);
nand U15729 (N_15729,N_13896,N_14497);
and U15730 (N_15730,N_14793,N_14314);
nand U15731 (N_15731,N_13546,N_13708);
nand U15732 (N_15732,N_14448,N_14159);
and U15733 (N_15733,N_14477,N_14742);
xnor U15734 (N_15734,N_14739,N_14653);
or U15735 (N_15735,N_14354,N_14648);
nor U15736 (N_15736,N_13840,N_14594);
nor U15737 (N_15737,N_14779,N_13633);
or U15738 (N_15738,N_13569,N_14465);
xor U15739 (N_15739,N_14500,N_14034);
nor U15740 (N_15740,N_14976,N_13982);
and U15741 (N_15741,N_13894,N_14502);
or U15742 (N_15742,N_13716,N_14795);
nand U15743 (N_15743,N_14302,N_14526);
nor U15744 (N_15744,N_14019,N_14768);
nor U15745 (N_15745,N_13755,N_13801);
and U15746 (N_15746,N_13692,N_13932);
xor U15747 (N_15747,N_14633,N_14214);
nand U15748 (N_15748,N_14751,N_13790);
xnor U15749 (N_15749,N_14281,N_13778);
and U15750 (N_15750,N_14002,N_14555);
nor U15751 (N_15751,N_14856,N_13854);
nor U15752 (N_15752,N_13771,N_13770);
xor U15753 (N_15753,N_13728,N_13770);
nand U15754 (N_15754,N_14092,N_13877);
nor U15755 (N_15755,N_14684,N_14589);
and U15756 (N_15756,N_14506,N_14549);
xnor U15757 (N_15757,N_14087,N_14599);
xor U15758 (N_15758,N_14783,N_14893);
or U15759 (N_15759,N_14139,N_14960);
and U15760 (N_15760,N_13589,N_14228);
nor U15761 (N_15761,N_13523,N_14900);
or U15762 (N_15762,N_13612,N_14046);
or U15763 (N_15763,N_14466,N_14669);
xor U15764 (N_15764,N_14092,N_14903);
and U15765 (N_15765,N_14019,N_13821);
and U15766 (N_15766,N_13717,N_14700);
xnor U15767 (N_15767,N_14746,N_14785);
or U15768 (N_15768,N_13634,N_14065);
and U15769 (N_15769,N_14625,N_14526);
nand U15770 (N_15770,N_13933,N_13743);
nand U15771 (N_15771,N_14733,N_13925);
or U15772 (N_15772,N_13989,N_13590);
or U15773 (N_15773,N_14290,N_14864);
xor U15774 (N_15774,N_13523,N_13724);
or U15775 (N_15775,N_13875,N_14474);
nand U15776 (N_15776,N_14520,N_14441);
xnor U15777 (N_15777,N_13797,N_14111);
nor U15778 (N_15778,N_13955,N_14642);
xnor U15779 (N_15779,N_13555,N_14270);
and U15780 (N_15780,N_14644,N_14086);
or U15781 (N_15781,N_14924,N_14175);
nand U15782 (N_15782,N_13588,N_14849);
nand U15783 (N_15783,N_14022,N_13989);
xor U15784 (N_15784,N_13988,N_14289);
or U15785 (N_15785,N_13564,N_14037);
and U15786 (N_15786,N_14764,N_14798);
nand U15787 (N_15787,N_13542,N_14604);
nor U15788 (N_15788,N_14605,N_13564);
nor U15789 (N_15789,N_14269,N_14101);
nand U15790 (N_15790,N_13740,N_14553);
nor U15791 (N_15791,N_14013,N_13813);
and U15792 (N_15792,N_14740,N_14803);
nand U15793 (N_15793,N_14018,N_14235);
xnor U15794 (N_15794,N_14938,N_14396);
or U15795 (N_15795,N_14211,N_13657);
and U15796 (N_15796,N_13636,N_14036);
xor U15797 (N_15797,N_14361,N_14063);
and U15798 (N_15798,N_14603,N_13705);
or U15799 (N_15799,N_14850,N_13511);
nor U15800 (N_15800,N_13999,N_14933);
nand U15801 (N_15801,N_14671,N_13820);
xnor U15802 (N_15802,N_14806,N_13656);
nand U15803 (N_15803,N_13958,N_14701);
nand U15804 (N_15804,N_14893,N_14558);
nor U15805 (N_15805,N_14924,N_13605);
nor U15806 (N_15806,N_14694,N_13856);
nand U15807 (N_15807,N_14640,N_14270);
and U15808 (N_15808,N_14598,N_14420);
or U15809 (N_15809,N_13619,N_13970);
and U15810 (N_15810,N_13859,N_14261);
or U15811 (N_15811,N_14121,N_13879);
xnor U15812 (N_15812,N_13751,N_13523);
or U15813 (N_15813,N_14458,N_13645);
and U15814 (N_15814,N_14340,N_13995);
or U15815 (N_15815,N_14020,N_13669);
nor U15816 (N_15816,N_13770,N_14673);
nor U15817 (N_15817,N_14535,N_13587);
nor U15818 (N_15818,N_13651,N_14336);
nor U15819 (N_15819,N_14046,N_14288);
and U15820 (N_15820,N_13529,N_14837);
or U15821 (N_15821,N_14683,N_14184);
and U15822 (N_15822,N_13555,N_13673);
nor U15823 (N_15823,N_14537,N_14867);
or U15824 (N_15824,N_13845,N_14388);
nor U15825 (N_15825,N_14435,N_13843);
and U15826 (N_15826,N_13920,N_14870);
xnor U15827 (N_15827,N_13527,N_14342);
xor U15828 (N_15828,N_14100,N_14907);
nand U15829 (N_15829,N_13711,N_14134);
and U15830 (N_15830,N_14766,N_13705);
nor U15831 (N_15831,N_13762,N_14949);
nand U15832 (N_15832,N_13808,N_14977);
nor U15833 (N_15833,N_14797,N_13747);
xnor U15834 (N_15834,N_14014,N_13988);
xnor U15835 (N_15835,N_13851,N_14790);
nor U15836 (N_15836,N_14528,N_13803);
or U15837 (N_15837,N_13718,N_14080);
or U15838 (N_15838,N_14747,N_14400);
xor U15839 (N_15839,N_14098,N_14367);
xor U15840 (N_15840,N_14974,N_14779);
or U15841 (N_15841,N_14148,N_13955);
and U15842 (N_15842,N_14536,N_14835);
xor U15843 (N_15843,N_14044,N_13858);
nand U15844 (N_15844,N_13549,N_14997);
nand U15845 (N_15845,N_14561,N_14161);
or U15846 (N_15846,N_13697,N_14356);
nand U15847 (N_15847,N_14155,N_14576);
xnor U15848 (N_15848,N_13830,N_14974);
nand U15849 (N_15849,N_14262,N_13712);
and U15850 (N_15850,N_14578,N_13647);
nand U15851 (N_15851,N_13582,N_13561);
or U15852 (N_15852,N_13812,N_14581);
or U15853 (N_15853,N_13847,N_13932);
nand U15854 (N_15854,N_13937,N_13661);
and U15855 (N_15855,N_14080,N_13730);
and U15856 (N_15856,N_14802,N_13500);
and U15857 (N_15857,N_13808,N_13991);
nand U15858 (N_15858,N_14573,N_13742);
and U15859 (N_15859,N_14278,N_14273);
xor U15860 (N_15860,N_14592,N_14675);
nor U15861 (N_15861,N_14410,N_14049);
nand U15862 (N_15862,N_13577,N_13816);
and U15863 (N_15863,N_14330,N_14830);
and U15864 (N_15864,N_14479,N_14399);
xnor U15865 (N_15865,N_14182,N_14066);
nand U15866 (N_15866,N_13897,N_14236);
and U15867 (N_15867,N_14146,N_13816);
and U15868 (N_15868,N_14375,N_14003);
or U15869 (N_15869,N_13880,N_14881);
nor U15870 (N_15870,N_13519,N_14454);
nand U15871 (N_15871,N_14590,N_13927);
xor U15872 (N_15872,N_13748,N_13831);
and U15873 (N_15873,N_14093,N_14141);
and U15874 (N_15874,N_13951,N_13937);
nand U15875 (N_15875,N_14917,N_14331);
nor U15876 (N_15876,N_14928,N_13999);
xnor U15877 (N_15877,N_14904,N_13892);
nor U15878 (N_15878,N_14478,N_14278);
nand U15879 (N_15879,N_13536,N_14130);
or U15880 (N_15880,N_13770,N_14490);
and U15881 (N_15881,N_13546,N_14893);
nor U15882 (N_15882,N_14394,N_13845);
nor U15883 (N_15883,N_14420,N_13870);
and U15884 (N_15884,N_14856,N_14794);
xnor U15885 (N_15885,N_14806,N_14462);
nor U15886 (N_15886,N_13861,N_14039);
or U15887 (N_15887,N_14380,N_13846);
nand U15888 (N_15888,N_13958,N_14523);
and U15889 (N_15889,N_14781,N_13953);
xor U15890 (N_15890,N_14021,N_13793);
and U15891 (N_15891,N_13847,N_14015);
nand U15892 (N_15892,N_14531,N_13962);
and U15893 (N_15893,N_14233,N_14227);
nand U15894 (N_15894,N_13782,N_14525);
or U15895 (N_15895,N_14671,N_14819);
or U15896 (N_15896,N_13533,N_14691);
nor U15897 (N_15897,N_14736,N_14161);
and U15898 (N_15898,N_14814,N_14242);
or U15899 (N_15899,N_13919,N_14628);
xnor U15900 (N_15900,N_13703,N_13817);
nor U15901 (N_15901,N_14701,N_14047);
and U15902 (N_15902,N_14830,N_14273);
and U15903 (N_15903,N_14917,N_13612);
nand U15904 (N_15904,N_14450,N_13948);
or U15905 (N_15905,N_14304,N_14398);
xnor U15906 (N_15906,N_14040,N_14486);
and U15907 (N_15907,N_13724,N_14691);
or U15908 (N_15908,N_14827,N_14554);
nand U15909 (N_15909,N_14897,N_14508);
nor U15910 (N_15910,N_14732,N_13849);
nand U15911 (N_15911,N_13970,N_14005);
nand U15912 (N_15912,N_14444,N_14547);
nor U15913 (N_15913,N_14976,N_14921);
nand U15914 (N_15914,N_14755,N_14173);
or U15915 (N_15915,N_14336,N_14293);
and U15916 (N_15916,N_14350,N_13851);
xor U15917 (N_15917,N_13933,N_14786);
xor U15918 (N_15918,N_14604,N_13654);
or U15919 (N_15919,N_14751,N_14279);
and U15920 (N_15920,N_14128,N_14268);
nor U15921 (N_15921,N_14533,N_13990);
and U15922 (N_15922,N_14941,N_14706);
xnor U15923 (N_15923,N_14339,N_14555);
nand U15924 (N_15924,N_14882,N_14620);
nand U15925 (N_15925,N_14051,N_14582);
nand U15926 (N_15926,N_13615,N_14715);
and U15927 (N_15927,N_13592,N_14515);
nor U15928 (N_15928,N_13657,N_14456);
xor U15929 (N_15929,N_14550,N_14578);
nand U15930 (N_15930,N_13579,N_14286);
nand U15931 (N_15931,N_14631,N_14897);
or U15932 (N_15932,N_13668,N_14884);
nand U15933 (N_15933,N_13689,N_13524);
xnor U15934 (N_15934,N_13839,N_13807);
nor U15935 (N_15935,N_14395,N_14736);
xor U15936 (N_15936,N_13702,N_14830);
nand U15937 (N_15937,N_13590,N_14505);
or U15938 (N_15938,N_14410,N_14756);
xor U15939 (N_15939,N_14291,N_14059);
and U15940 (N_15940,N_14351,N_14255);
or U15941 (N_15941,N_14057,N_14005);
or U15942 (N_15942,N_13537,N_13698);
xnor U15943 (N_15943,N_13557,N_13706);
and U15944 (N_15944,N_14595,N_14418);
nor U15945 (N_15945,N_14979,N_13788);
xor U15946 (N_15946,N_14208,N_14749);
and U15947 (N_15947,N_14963,N_14105);
or U15948 (N_15948,N_13935,N_14790);
nand U15949 (N_15949,N_13881,N_14994);
nand U15950 (N_15950,N_14818,N_14359);
or U15951 (N_15951,N_14653,N_14304);
nor U15952 (N_15952,N_13705,N_14344);
xor U15953 (N_15953,N_13765,N_14243);
nand U15954 (N_15954,N_13560,N_13757);
or U15955 (N_15955,N_14442,N_14986);
or U15956 (N_15956,N_13730,N_14469);
xor U15957 (N_15957,N_14512,N_13746);
and U15958 (N_15958,N_13798,N_14044);
or U15959 (N_15959,N_14217,N_14916);
or U15960 (N_15960,N_14869,N_13733);
nor U15961 (N_15961,N_13788,N_14103);
or U15962 (N_15962,N_14321,N_13700);
and U15963 (N_15963,N_13617,N_14790);
or U15964 (N_15964,N_14538,N_14724);
and U15965 (N_15965,N_14402,N_14296);
or U15966 (N_15966,N_14795,N_14051);
xor U15967 (N_15967,N_14230,N_13575);
xnor U15968 (N_15968,N_14309,N_14965);
xnor U15969 (N_15969,N_14689,N_13827);
or U15970 (N_15970,N_13954,N_14357);
and U15971 (N_15971,N_14828,N_14936);
nand U15972 (N_15972,N_13903,N_14566);
nor U15973 (N_15973,N_14879,N_14042);
xnor U15974 (N_15974,N_14010,N_14140);
or U15975 (N_15975,N_14702,N_13613);
xor U15976 (N_15976,N_13512,N_13555);
nand U15977 (N_15977,N_13674,N_14268);
nand U15978 (N_15978,N_14620,N_14274);
nand U15979 (N_15979,N_14104,N_14395);
xnor U15980 (N_15980,N_14882,N_14928);
xnor U15981 (N_15981,N_13823,N_14546);
xor U15982 (N_15982,N_14962,N_14313);
nand U15983 (N_15983,N_14066,N_14104);
nor U15984 (N_15984,N_13699,N_14594);
nor U15985 (N_15985,N_13531,N_14433);
nor U15986 (N_15986,N_13922,N_14224);
and U15987 (N_15987,N_14020,N_14240);
or U15988 (N_15988,N_14452,N_14259);
nor U15989 (N_15989,N_13559,N_14046);
nor U15990 (N_15990,N_13585,N_14493);
or U15991 (N_15991,N_13647,N_14740);
xor U15992 (N_15992,N_14547,N_14634);
or U15993 (N_15993,N_14002,N_14352);
xnor U15994 (N_15994,N_14422,N_14584);
and U15995 (N_15995,N_14275,N_14915);
xor U15996 (N_15996,N_14237,N_14361);
nand U15997 (N_15997,N_14845,N_14272);
nand U15998 (N_15998,N_13997,N_14528);
or U15999 (N_15999,N_14950,N_14524);
and U16000 (N_16000,N_14538,N_14911);
nor U16001 (N_16001,N_14785,N_13989);
nand U16002 (N_16002,N_14781,N_13684);
nor U16003 (N_16003,N_14788,N_14040);
and U16004 (N_16004,N_14549,N_14879);
nor U16005 (N_16005,N_13620,N_13827);
nor U16006 (N_16006,N_13559,N_14434);
or U16007 (N_16007,N_14670,N_14752);
xor U16008 (N_16008,N_14003,N_14200);
and U16009 (N_16009,N_14231,N_14833);
and U16010 (N_16010,N_14147,N_14404);
nand U16011 (N_16011,N_14088,N_14570);
or U16012 (N_16012,N_14705,N_14573);
or U16013 (N_16013,N_13889,N_13743);
nand U16014 (N_16014,N_14698,N_14736);
nand U16015 (N_16015,N_14412,N_14107);
nand U16016 (N_16016,N_14497,N_14724);
and U16017 (N_16017,N_13640,N_13785);
and U16018 (N_16018,N_14843,N_13952);
or U16019 (N_16019,N_14710,N_14527);
nand U16020 (N_16020,N_13952,N_13559);
xor U16021 (N_16021,N_13755,N_14921);
nor U16022 (N_16022,N_13515,N_14529);
nand U16023 (N_16023,N_14619,N_14411);
xor U16024 (N_16024,N_13677,N_13768);
xor U16025 (N_16025,N_13960,N_14623);
xor U16026 (N_16026,N_14020,N_14299);
nor U16027 (N_16027,N_14181,N_14129);
and U16028 (N_16028,N_14039,N_14877);
and U16029 (N_16029,N_13582,N_14675);
nor U16030 (N_16030,N_13895,N_13731);
xor U16031 (N_16031,N_13941,N_14662);
and U16032 (N_16032,N_14777,N_14414);
or U16033 (N_16033,N_13645,N_13883);
nand U16034 (N_16034,N_14417,N_13569);
xor U16035 (N_16035,N_14715,N_14997);
or U16036 (N_16036,N_14404,N_14980);
xnor U16037 (N_16037,N_14182,N_13782);
xor U16038 (N_16038,N_13675,N_14061);
or U16039 (N_16039,N_13862,N_14441);
nor U16040 (N_16040,N_14664,N_14566);
xnor U16041 (N_16041,N_13995,N_14108);
nand U16042 (N_16042,N_14419,N_14435);
nor U16043 (N_16043,N_13712,N_13955);
nor U16044 (N_16044,N_14325,N_14547);
nor U16045 (N_16045,N_14603,N_14977);
nand U16046 (N_16046,N_14819,N_13881);
or U16047 (N_16047,N_14433,N_14057);
nor U16048 (N_16048,N_14377,N_14795);
xor U16049 (N_16049,N_14076,N_14078);
nor U16050 (N_16050,N_13828,N_14542);
nor U16051 (N_16051,N_13650,N_14335);
nand U16052 (N_16052,N_13670,N_13859);
or U16053 (N_16053,N_13519,N_14473);
and U16054 (N_16054,N_14202,N_14679);
and U16055 (N_16055,N_14741,N_14819);
xnor U16056 (N_16056,N_13732,N_13620);
nand U16057 (N_16057,N_14418,N_14672);
or U16058 (N_16058,N_14035,N_14470);
nor U16059 (N_16059,N_14647,N_14616);
xnor U16060 (N_16060,N_14893,N_14965);
nand U16061 (N_16061,N_14096,N_14106);
or U16062 (N_16062,N_14867,N_14711);
nor U16063 (N_16063,N_14775,N_13979);
or U16064 (N_16064,N_13699,N_14872);
nand U16065 (N_16065,N_13930,N_13858);
nand U16066 (N_16066,N_13839,N_13674);
xnor U16067 (N_16067,N_14837,N_14081);
and U16068 (N_16068,N_13842,N_14589);
nand U16069 (N_16069,N_14332,N_14167);
xor U16070 (N_16070,N_13769,N_14752);
nor U16071 (N_16071,N_14871,N_14665);
or U16072 (N_16072,N_13940,N_14331);
and U16073 (N_16073,N_14306,N_14437);
and U16074 (N_16074,N_13756,N_14220);
and U16075 (N_16075,N_13657,N_14929);
nor U16076 (N_16076,N_14401,N_14976);
xnor U16077 (N_16077,N_14859,N_14188);
or U16078 (N_16078,N_14052,N_13757);
or U16079 (N_16079,N_14714,N_13762);
and U16080 (N_16080,N_13584,N_14105);
xnor U16081 (N_16081,N_14163,N_14248);
or U16082 (N_16082,N_14621,N_14297);
xor U16083 (N_16083,N_14227,N_14058);
xor U16084 (N_16084,N_13551,N_14077);
and U16085 (N_16085,N_13668,N_13828);
nand U16086 (N_16086,N_14520,N_13739);
or U16087 (N_16087,N_14140,N_14684);
or U16088 (N_16088,N_14059,N_14732);
xnor U16089 (N_16089,N_14145,N_14754);
xnor U16090 (N_16090,N_14648,N_13873);
nand U16091 (N_16091,N_13568,N_13861);
nor U16092 (N_16092,N_14351,N_14415);
xor U16093 (N_16093,N_13839,N_13753);
nand U16094 (N_16094,N_14775,N_14769);
and U16095 (N_16095,N_14626,N_13840);
and U16096 (N_16096,N_13877,N_14326);
and U16097 (N_16097,N_13832,N_13709);
and U16098 (N_16098,N_14309,N_14702);
nand U16099 (N_16099,N_14063,N_13640);
xor U16100 (N_16100,N_14304,N_13940);
and U16101 (N_16101,N_14059,N_13722);
or U16102 (N_16102,N_14196,N_13810);
nand U16103 (N_16103,N_14004,N_14979);
or U16104 (N_16104,N_14704,N_14289);
nor U16105 (N_16105,N_13992,N_13918);
nand U16106 (N_16106,N_13590,N_14265);
or U16107 (N_16107,N_13853,N_13666);
or U16108 (N_16108,N_13509,N_14378);
xnor U16109 (N_16109,N_14472,N_14041);
or U16110 (N_16110,N_13695,N_13677);
or U16111 (N_16111,N_14092,N_14040);
and U16112 (N_16112,N_14988,N_14809);
xor U16113 (N_16113,N_13573,N_14132);
and U16114 (N_16114,N_14543,N_14965);
and U16115 (N_16115,N_13865,N_14727);
nor U16116 (N_16116,N_14385,N_14663);
and U16117 (N_16117,N_14481,N_14283);
or U16118 (N_16118,N_14023,N_14722);
nand U16119 (N_16119,N_14579,N_14215);
or U16120 (N_16120,N_14295,N_13657);
nor U16121 (N_16121,N_14898,N_14405);
or U16122 (N_16122,N_14721,N_13952);
xor U16123 (N_16123,N_13745,N_14029);
or U16124 (N_16124,N_14238,N_13786);
xnor U16125 (N_16125,N_14847,N_13522);
nor U16126 (N_16126,N_13523,N_13757);
xnor U16127 (N_16127,N_14412,N_14433);
nor U16128 (N_16128,N_14398,N_13603);
xor U16129 (N_16129,N_14819,N_14431);
or U16130 (N_16130,N_13730,N_14305);
xnor U16131 (N_16131,N_14071,N_13829);
nor U16132 (N_16132,N_14560,N_13876);
nand U16133 (N_16133,N_14991,N_14042);
xnor U16134 (N_16134,N_13682,N_14679);
nand U16135 (N_16135,N_13937,N_13681);
nor U16136 (N_16136,N_14446,N_14903);
nor U16137 (N_16137,N_13623,N_14052);
nand U16138 (N_16138,N_14267,N_14744);
xnor U16139 (N_16139,N_14154,N_13596);
nor U16140 (N_16140,N_14331,N_13546);
xor U16141 (N_16141,N_14054,N_13811);
nand U16142 (N_16142,N_13908,N_14958);
nand U16143 (N_16143,N_14068,N_14450);
xor U16144 (N_16144,N_14055,N_13554);
xnor U16145 (N_16145,N_13866,N_13522);
and U16146 (N_16146,N_13907,N_14709);
xnor U16147 (N_16147,N_13875,N_13552);
xnor U16148 (N_16148,N_13822,N_14735);
nand U16149 (N_16149,N_13633,N_13574);
xnor U16150 (N_16150,N_13715,N_14149);
or U16151 (N_16151,N_14613,N_14929);
nor U16152 (N_16152,N_14347,N_14756);
or U16153 (N_16153,N_14000,N_13712);
xor U16154 (N_16154,N_14951,N_14918);
or U16155 (N_16155,N_14282,N_13751);
xor U16156 (N_16156,N_13853,N_14382);
or U16157 (N_16157,N_14229,N_14017);
nand U16158 (N_16158,N_14658,N_14650);
and U16159 (N_16159,N_14624,N_14457);
xor U16160 (N_16160,N_14576,N_14181);
and U16161 (N_16161,N_13536,N_14801);
nor U16162 (N_16162,N_14564,N_14893);
xor U16163 (N_16163,N_14519,N_13589);
nor U16164 (N_16164,N_13557,N_13548);
and U16165 (N_16165,N_13562,N_14167);
nor U16166 (N_16166,N_14572,N_14324);
or U16167 (N_16167,N_13642,N_13555);
nand U16168 (N_16168,N_14294,N_13753);
nor U16169 (N_16169,N_14042,N_13548);
or U16170 (N_16170,N_14096,N_14415);
and U16171 (N_16171,N_13772,N_14049);
and U16172 (N_16172,N_14096,N_14073);
nand U16173 (N_16173,N_14333,N_14775);
xor U16174 (N_16174,N_14777,N_13657);
or U16175 (N_16175,N_13744,N_13630);
and U16176 (N_16176,N_14567,N_14906);
and U16177 (N_16177,N_14986,N_14559);
nand U16178 (N_16178,N_14927,N_14519);
xor U16179 (N_16179,N_13969,N_14904);
xnor U16180 (N_16180,N_14762,N_13879);
or U16181 (N_16181,N_14686,N_14693);
and U16182 (N_16182,N_14433,N_14285);
xor U16183 (N_16183,N_14919,N_14562);
xor U16184 (N_16184,N_13683,N_14109);
nor U16185 (N_16185,N_14760,N_13984);
or U16186 (N_16186,N_13705,N_13815);
nand U16187 (N_16187,N_13624,N_13829);
nand U16188 (N_16188,N_13726,N_14582);
and U16189 (N_16189,N_14604,N_14690);
and U16190 (N_16190,N_14930,N_13579);
nand U16191 (N_16191,N_13535,N_14651);
or U16192 (N_16192,N_13704,N_13543);
and U16193 (N_16193,N_13676,N_14055);
or U16194 (N_16194,N_14942,N_14027);
nor U16195 (N_16195,N_13701,N_14889);
nand U16196 (N_16196,N_14574,N_14289);
xnor U16197 (N_16197,N_14183,N_13549);
nor U16198 (N_16198,N_14578,N_13869);
xor U16199 (N_16199,N_13723,N_14523);
and U16200 (N_16200,N_14702,N_14360);
or U16201 (N_16201,N_13619,N_14747);
xnor U16202 (N_16202,N_14534,N_13716);
nand U16203 (N_16203,N_13590,N_14273);
xor U16204 (N_16204,N_14220,N_14540);
xor U16205 (N_16205,N_14209,N_14070);
and U16206 (N_16206,N_14970,N_14164);
or U16207 (N_16207,N_13633,N_14179);
nand U16208 (N_16208,N_14655,N_14356);
nor U16209 (N_16209,N_14398,N_13688);
xnor U16210 (N_16210,N_13631,N_14997);
or U16211 (N_16211,N_13867,N_14950);
nor U16212 (N_16212,N_14192,N_14409);
or U16213 (N_16213,N_14160,N_13884);
or U16214 (N_16214,N_13922,N_14876);
xor U16215 (N_16215,N_13913,N_14261);
nor U16216 (N_16216,N_14713,N_14148);
or U16217 (N_16217,N_14086,N_14601);
nor U16218 (N_16218,N_13828,N_14554);
or U16219 (N_16219,N_13626,N_14680);
or U16220 (N_16220,N_14913,N_14109);
and U16221 (N_16221,N_14308,N_13906);
or U16222 (N_16222,N_14888,N_14945);
and U16223 (N_16223,N_14919,N_14798);
nor U16224 (N_16224,N_13939,N_14271);
and U16225 (N_16225,N_13638,N_14160);
or U16226 (N_16226,N_14337,N_14795);
xor U16227 (N_16227,N_14789,N_13925);
nor U16228 (N_16228,N_14002,N_14033);
or U16229 (N_16229,N_14455,N_14559);
xor U16230 (N_16230,N_13654,N_13531);
nand U16231 (N_16231,N_14696,N_14594);
or U16232 (N_16232,N_14463,N_13779);
xnor U16233 (N_16233,N_14081,N_14849);
xnor U16234 (N_16234,N_14406,N_14115);
nand U16235 (N_16235,N_13637,N_14647);
or U16236 (N_16236,N_14089,N_14242);
and U16237 (N_16237,N_14173,N_14358);
or U16238 (N_16238,N_13747,N_14449);
nor U16239 (N_16239,N_14808,N_14256);
xnor U16240 (N_16240,N_14157,N_14933);
or U16241 (N_16241,N_14425,N_14437);
nand U16242 (N_16242,N_14051,N_14036);
nand U16243 (N_16243,N_14754,N_13844);
nor U16244 (N_16244,N_14937,N_14726);
xor U16245 (N_16245,N_14896,N_13641);
nand U16246 (N_16246,N_14277,N_13511);
or U16247 (N_16247,N_14443,N_13538);
nor U16248 (N_16248,N_14356,N_13857);
xor U16249 (N_16249,N_14946,N_14035);
nor U16250 (N_16250,N_13798,N_14783);
xor U16251 (N_16251,N_14682,N_13701);
nand U16252 (N_16252,N_14192,N_13665);
nand U16253 (N_16253,N_14530,N_14322);
nor U16254 (N_16254,N_14642,N_14726);
xnor U16255 (N_16255,N_13791,N_14076);
or U16256 (N_16256,N_14648,N_14721);
nand U16257 (N_16257,N_13624,N_13842);
and U16258 (N_16258,N_14579,N_14079);
or U16259 (N_16259,N_13627,N_14630);
xor U16260 (N_16260,N_14430,N_13859);
and U16261 (N_16261,N_14856,N_14393);
and U16262 (N_16262,N_14448,N_13585);
and U16263 (N_16263,N_14492,N_14827);
nand U16264 (N_16264,N_14031,N_13777);
and U16265 (N_16265,N_14922,N_13879);
and U16266 (N_16266,N_13894,N_13804);
nand U16267 (N_16267,N_14823,N_13566);
or U16268 (N_16268,N_13893,N_14477);
nor U16269 (N_16269,N_14929,N_14794);
nand U16270 (N_16270,N_14103,N_14180);
nand U16271 (N_16271,N_13586,N_14669);
xor U16272 (N_16272,N_14931,N_14862);
and U16273 (N_16273,N_14599,N_13891);
xnor U16274 (N_16274,N_14995,N_14831);
and U16275 (N_16275,N_14576,N_13662);
and U16276 (N_16276,N_13847,N_14948);
and U16277 (N_16277,N_13522,N_14132);
xnor U16278 (N_16278,N_13722,N_14851);
nor U16279 (N_16279,N_14212,N_14839);
xor U16280 (N_16280,N_14545,N_14724);
and U16281 (N_16281,N_14643,N_14311);
and U16282 (N_16282,N_14866,N_14014);
and U16283 (N_16283,N_14210,N_14354);
and U16284 (N_16284,N_14752,N_14627);
nand U16285 (N_16285,N_13786,N_14769);
nor U16286 (N_16286,N_14262,N_14400);
nor U16287 (N_16287,N_14776,N_14576);
xor U16288 (N_16288,N_13893,N_13840);
xor U16289 (N_16289,N_14213,N_14774);
nor U16290 (N_16290,N_14650,N_13932);
or U16291 (N_16291,N_14115,N_14081);
xor U16292 (N_16292,N_14427,N_13734);
or U16293 (N_16293,N_14447,N_14273);
or U16294 (N_16294,N_14327,N_14089);
nand U16295 (N_16295,N_13719,N_13787);
nor U16296 (N_16296,N_13785,N_14906);
and U16297 (N_16297,N_14519,N_14038);
and U16298 (N_16298,N_13767,N_14575);
or U16299 (N_16299,N_14234,N_14720);
xor U16300 (N_16300,N_14279,N_13945);
or U16301 (N_16301,N_14298,N_14121);
nand U16302 (N_16302,N_14343,N_14325);
xor U16303 (N_16303,N_13628,N_13933);
xor U16304 (N_16304,N_13862,N_14321);
and U16305 (N_16305,N_14856,N_14416);
and U16306 (N_16306,N_14240,N_14533);
and U16307 (N_16307,N_14620,N_13738);
xnor U16308 (N_16308,N_14016,N_14256);
nor U16309 (N_16309,N_13708,N_13628);
nand U16310 (N_16310,N_13651,N_13931);
nor U16311 (N_16311,N_14238,N_14672);
xor U16312 (N_16312,N_14507,N_13529);
or U16313 (N_16313,N_14888,N_14861);
nor U16314 (N_16314,N_14514,N_14271);
and U16315 (N_16315,N_14953,N_13571);
nor U16316 (N_16316,N_14559,N_14539);
and U16317 (N_16317,N_14994,N_13874);
nor U16318 (N_16318,N_14961,N_14838);
nor U16319 (N_16319,N_14833,N_14710);
or U16320 (N_16320,N_14121,N_14459);
or U16321 (N_16321,N_14460,N_13827);
or U16322 (N_16322,N_14771,N_14516);
or U16323 (N_16323,N_14551,N_14281);
nor U16324 (N_16324,N_14026,N_13553);
or U16325 (N_16325,N_14386,N_14856);
nor U16326 (N_16326,N_13720,N_14596);
or U16327 (N_16327,N_14168,N_14311);
xor U16328 (N_16328,N_14214,N_14253);
or U16329 (N_16329,N_14303,N_14197);
or U16330 (N_16330,N_14571,N_14140);
nor U16331 (N_16331,N_14067,N_13623);
nand U16332 (N_16332,N_14483,N_14030);
and U16333 (N_16333,N_14065,N_13917);
or U16334 (N_16334,N_14528,N_14416);
nand U16335 (N_16335,N_14599,N_13959);
xor U16336 (N_16336,N_14544,N_14472);
nand U16337 (N_16337,N_13792,N_14454);
nor U16338 (N_16338,N_13578,N_14239);
nand U16339 (N_16339,N_13980,N_14904);
and U16340 (N_16340,N_13718,N_13855);
xnor U16341 (N_16341,N_13782,N_14524);
and U16342 (N_16342,N_13876,N_13541);
nand U16343 (N_16343,N_14547,N_14194);
xnor U16344 (N_16344,N_13977,N_14412);
and U16345 (N_16345,N_14408,N_13772);
or U16346 (N_16346,N_14551,N_13580);
or U16347 (N_16347,N_13558,N_14209);
nor U16348 (N_16348,N_14788,N_14280);
nor U16349 (N_16349,N_14684,N_14645);
and U16350 (N_16350,N_14139,N_14563);
xnor U16351 (N_16351,N_13799,N_13741);
nor U16352 (N_16352,N_14915,N_13892);
nand U16353 (N_16353,N_14940,N_14419);
nand U16354 (N_16354,N_14200,N_13995);
or U16355 (N_16355,N_14682,N_14999);
and U16356 (N_16356,N_14670,N_14951);
xor U16357 (N_16357,N_14015,N_14804);
xnor U16358 (N_16358,N_13555,N_13511);
xor U16359 (N_16359,N_14162,N_14392);
xor U16360 (N_16360,N_14988,N_13865);
xor U16361 (N_16361,N_13730,N_13926);
and U16362 (N_16362,N_13781,N_14444);
xnor U16363 (N_16363,N_14705,N_14770);
xor U16364 (N_16364,N_14439,N_13938);
and U16365 (N_16365,N_14982,N_14550);
and U16366 (N_16366,N_14140,N_14805);
nor U16367 (N_16367,N_14767,N_13752);
nor U16368 (N_16368,N_14902,N_14248);
nand U16369 (N_16369,N_14648,N_14584);
xor U16370 (N_16370,N_14757,N_14418);
and U16371 (N_16371,N_13788,N_14923);
xnor U16372 (N_16372,N_13845,N_14414);
nand U16373 (N_16373,N_14877,N_14436);
or U16374 (N_16374,N_13712,N_14306);
xor U16375 (N_16375,N_14432,N_14094);
or U16376 (N_16376,N_14195,N_14949);
nand U16377 (N_16377,N_14238,N_14093);
and U16378 (N_16378,N_13874,N_14845);
and U16379 (N_16379,N_14734,N_14072);
nand U16380 (N_16380,N_14718,N_13863);
or U16381 (N_16381,N_13967,N_14469);
xor U16382 (N_16382,N_14410,N_13578);
or U16383 (N_16383,N_14806,N_14424);
or U16384 (N_16384,N_14197,N_14897);
and U16385 (N_16385,N_14713,N_13653);
or U16386 (N_16386,N_14678,N_14506);
and U16387 (N_16387,N_14942,N_14172);
nand U16388 (N_16388,N_13888,N_14315);
and U16389 (N_16389,N_14802,N_14137);
nand U16390 (N_16390,N_14864,N_14275);
or U16391 (N_16391,N_14664,N_13965);
nand U16392 (N_16392,N_13794,N_14465);
nor U16393 (N_16393,N_14445,N_13817);
nor U16394 (N_16394,N_13742,N_13815);
nand U16395 (N_16395,N_14357,N_14448);
or U16396 (N_16396,N_13673,N_14516);
nor U16397 (N_16397,N_14620,N_14124);
nand U16398 (N_16398,N_14632,N_14521);
or U16399 (N_16399,N_13774,N_13847);
nand U16400 (N_16400,N_14363,N_14094);
or U16401 (N_16401,N_14120,N_14198);
and U16402 (N_16402,N_14770,N_14448);
nand U16403 (N_16403,N_14658,N_13842);
nand U16404 (N_16404,N_14731,N_14242);
nand U16405 (N_16405,N_14591,N_14478);
or U16406 (N_16406,N_13941,N_14838);
nand U16407 (N_16407,N_14950,N_14597);
nand U16408 (N_16408,N_14630,N_14542);
xnor U16409 (N_16409,N_14238,N_14776);
or U16410 (N_16410,N_13910,N_14528);
xnor U16411 (N_16411,N_14552,N_14356);
xnor U16412 (N_16412,N_14688,N_14180);
nor U16413 (N_16413,N_13837,N_14612);
and U16414 (N_16414,N_13909,N_14231);
nor U16415 (N_16415,N_14859,N_14501);
xnor U16416 (N_16416,N_14825,N_13644);
and U16417 (N_16417,N_14440,N_13841);
or U16418 (N_16418,N_14522,N_14753);
and U16419 (N_16419,N_14832,N_14427);
and U16420 (N_16420,N_14247,N_14947);
nor U16421 (N_16421,N_14511,N_14845);
nand U16422 (N_16422,N_14187,N_14983);
xnor U16423 (N_16423,N_14527,N_14774);
nor U16424 (N_16424,N_14475,N_13920);
nand U16425 (N_16425,N_14321,N_14145);
xnor U16426 (N_16426,N_13744,N_14111);
xnor U16427 (N_16427,N_14245,N_14698);
nand U16428 (N_16428,N_14271,N_13569);
and U16429 (N_16429,N_14864,N_14536);
nor U16430 (N_16430,N_14877,N_14055);
and U16431 (N_16431,N_14493,N_14760);
xnor U16432 (N_16432,N_14881,N_14788);
nand U16433 (N_16433,N_13856,N_13914);
nand U16434 (N_16434,N_14192,N_14347);
nor U16435 (N_16435,N_14423,N_14984);
xnor U16436 (N_16436,N_13863,N_13885);
and U16437 (N_16437,N_14068,N_13612);
or U16438 (N_16438,N_13746,N_13846);
nor U16439 (N_16439,N_14965,N_14347);
nand U16440 (N_16440,N_14074,N_14023);
nor U16441 (N_16441,N_14389,N_14330);
nand U16442 (N_16442,N_13911,N_14251);
and U16443 (N_16443,N_13736,N_14715);
xnor U16444 (N_16444,N_13834,N_14251);
or U16445 (N_16445,N_14170,N_14649);
or U16446 (N_16446,N_14515,N_13585);
or U16447 (N_16447,N_14291,N_14028);
and U16448 (N_16448,N_13640,N_13806);
xnor U16449 (N_16449,N_14291,N_13944);
or U16450 (N_16450,N_14935,N_14260);
xor U16451 (N_16451,N_13839,N_14073);
xnor U16452 (N_16452,N_13684,N_14743);
nand U16453 (N_16453,N_13655,N_13722);
or U16454 (N_16454,N_14070,N_14348);
nand U16455 (N_16455,N_13583,N_14949);
or U16456 (N_16456,N_14565,N_14510);
xor U16457 (N_16457,N_14892,N_14420);
nor U16458 (N_16458,N_13915,N_13519);
xor U16459 (N_16459,N_14791,N_14353);
nor U16460 (N_16460,N_14533,N_13536);
xnor U16461 (N_16461,N_14748,N_14602);
and U16462 (N_16462,N_14816,N_14650);
or U16463 (N_16463,N_14606,N_14397);
nor U16464 (N_16464,N_13518,N_14201);
xnor U16465 (N_16465,N_14481,N_14019);
nor U16466 (N_16466,N_13630,N_14787);
and U16467 (N_16467,N_13652,N_14451);
xnor U16468 (N_16468,N_14418,N_13743);
or U16469 (N_16469,N_14126,N_14594);
or U16470 (N_16470,N_13815,N_14274);
nand U16471 (N_16471,N_14880,N_13665);
and U16472 (N_16472,N_13962,N_14712);
and U16473 (N_16473,N_14137,N_14886);
or U16474 (N_16474,N_13690,N_14710);
xnor U16475 (N_16475,N_14394,N_13688);
xnor U16476 (N_16476,N_14434,N_14119);
nand U16477 (N_16477,N_13806,N_14079);
nand U16478 (N_16478,N_14295,N_14196);
nor U16479 (N_16479,N_14219,N_14651);
nand U16480 (N_16480,N_14154,N_14299);
xnor U16481 (N_16481,N_14808,N_14400);
or U16482 (N_16482,N_13865,N_14661);
or U16483 (N_16483,N_14447,N_13733);
and U16484 (N_16484,N_14489,N_14787);
or U16485 (N_16485,N_13675,N_14303);
xor U16486 (N_16486,N_14878,N_14730);
nor U16487 (N_16487,N_14209,N_14450);
or U16488 (N_16488,N_14310,N_13934);
or U16489 (N_16489,N_14325,N_13872);
xor U16490 (N_16490,N_14348,N_14579);
and U16491 (N_16491,N_14931,N_13537);
and U16492 (N_16492,N_14290,N_14307);
xnor U16493 (N_16493,N_14450,N_13819);
and U16494 (N_16494,N_14265,N_13569);
nor U16495 (N_16495,N_13979,N_14466);
or U16496 (N_16496,N_13851,N_13865);
nor U16497 (N_16497,N_13560,N_13926);
or U16498 (N_16498,N_14473,N_14351);
or U16499 (N_16499,N_13716,N_14626);
xor U16500 (N_16500,N_15634,N_15602);
and U16501 (N_16501,N_16300,N_15721);
nand U16502 (N_16502,N_16218,N_15352);
or U16503 (N_16503,N_15824,N_15718);
nor U16504 (N_16504,N_15029,N_15270);
xnor U16505 (N_16505,N_16270,N_15748);
xnor U16506 (N_16506,N_16335,N_15780);
xnor U16507 (N_16507,N_15669,N_15661);
nor U16508 (N_16508,N_15524,N_15781);
and U16509 (N_16509,N_15837,N_15540);
or U16510 (N_16510,N_16238,N_15910);
nor U16511 (N_16511,N_15290,N_15859);
or U16512 (N_16512,N_15695,N_16329);
and U16513 (N_16513,N_15257,N_16384);
or U16514 (N_16514,N_15100,N_15719);
xor U16515 (N_16515,N_15127,N_16129);
xor U16516 (N_16516,N_15903,N_15967);
or U16517 (N_16517,N_15348,N_15958);
xor U16518 (N_16518,N_16356,N_16282);
nand U16519 (N_16519,N_15071,N_16181);
or U16520 (N_16520,N_16370,N_15720);
and U16521 (N_16521,N_16308,N_15789);
and U16522 (N_16522,N_15849,N_15993);
or U16523 (N_16523,N_15788,N_16199);
nand U16524 (N_16524,N_15798,N_15120);
or U16525 (N_16525,N_16266,N_15950);
xnor U16526 (N_16526,N_15851,N_15298);
and U16527 (N_16527,N_15828,N_15587);
nand U16528 (N_16528,N_15553,N_15288);
nor U16529 (N_16529,N_15826,N_16399);
nor U16530 (N_16530,N_16277,N_15434);
and U16531 (N_16531,N_16034,N_15327);
nor U16532 (N_16532,N_15920,N_15782);
nand U16533 (N_16533,N_16289,N_15373);
or U16534 (N_16534,N_15992,N_15116);
and U16535 (N_16535,N_16011,N_16097);
and U16536 (N_16536,N_16193,N_15570);
and U16537 (N_16537,N_15107,N_16130);
nor U16538 (N_16538,N_16183,N_15583);
xor U16539 (N_16539,N_15916,N_16051);
and U16540 (N_16540,N_15654,N_15905);
or U16541 (N_16541,N_16336,N_15363);
and U16542 (N_16542,N_15547,N_15049);
and U16543 (N_16543,N_16404,N_15086);
nand U16544 (N_16544,N_15980,N_16026);
and U16545 (N_16545,N_16171,N_16142);
xor U16546 (N_16546,N_15513,N_15836);
nor U16547 (N_16547,N_15699,N_16231);
nand U16548 (N_16548,N_16100,N_15066);
or U16549 (N_16549,N_15221,N_15390);
nor U16550 (N_16550,N_15083,N_15237);
nand U16551 (N_16551,N_16196,N_15433);
xor U16552 (N_16552,N_16121,N_16151);
nor U16553 (N_16553,N_16488,N_15953);
nand U16554 (N_16554,N_15409,N_15263);
or U16555 (N_16555,N_15222,N_16327);
nor U16556 (N_16556,N_15504,N_15918);
xnor U16557 (N_16557,N_15364,N_16153);
nor U16558 (N_16558,N_16072,N_15907);
and U16559 (N_16559,N_15225,N_16451);
and U16560 (N_16560,N_16297,N_15114);
xor U16561 (N_16561,N_15561,N_15538);
and U16562 (N_16562,N_16145,N_15726);
nor U16563 (N_16563,N_15179,N_15472);
nor U16564 (N_16564,N_16217,N_15823);
and U16565 (N_16565,N_16163,N_15090);
and U16566 (N_16566,N_15722,N_15834);
nor U16567 (N_16567,N_16331,N_16406);
xnor U16568 (N_16568,N_15696,N_16432);
and U16569 (N_16569,N_15601,N_15186);
xnor U16570 (N_16570,N_16295,N_16273);
nand U16571 (N_16571,N_15243,N_15501);
xor U16572 (N_16572,N_15644,N_15190);
and U16573 (N_16573,N_15153,N_16111);
and U16574 (N_16574,N_16321,N_16478);
and U16575 (N_16575,N_15240,N_16002);
xor U16576 (N_16576,N_15284,N_15934);
or U16577 (N_16577,N_15974,N_15316);
or U16578 (N_16578,N_15751,N_15329);
nor U16579 (N_16579,N_15020,N_15783);
nand U16580 (N_16580,N_15450,N_16016);
or U16581 (N_16581,N_16019,N_15685);
or U16582 (N_16582,N_15737,N_16380);
nor U16583 (N_16583,N_15238,N_16446);
nor U16584 (N_16584,N_15820,N_16101);
or U16585 (N_16585,N_15733,N_15128);
xor U16586 (N_16586,N_16208,N_16303);
and U16587 (N_16587,N_16108,N_15063);
nand U16588 (N_16588,N_16080,N_15728);
and U16589 (N_16589,N_15546,N_15843);
nor U16590 (N_16590,N_16346,N_15503);
nand U16591 (N_16591,N_15692,N_15267);
and U16592 (N_16592,N_16292,N_16029);
or U16593 (N_16593,N_16400,N_15228);
or U16594 (N_16594,N_15764,N_16443);
xor U16595 (N_16595,N_16093,N_15785);
nor U16596 (N_16596,N_15088,N_15710);
nor U16597 (N_16597,N_15014,N_15527);
nand U16598 (N_16598,N_15328,N_15101);
nand U16599 (N_16599,N_15103,N_15375);
or U16600 (N_16600,N_16168,N_16147);
nor U16601 (N_16601,N_15191,N_16060);
and U16602 (N_16602,N_15314,N_16479);
or U16603 (N_16603,N_15484,N_16460);
xor U16604 (N_16604,N_16189,N_15831);
xnor U16605 (N_16605,N_15203,N_16260);
nand U16606 (N_16606,N_15972,N_15704);
or U16607 (N_16607,N_15060,N_16000);
nand U16608 (N_16608,N_15717,N_16304);
and U16609 (N_16609,N_15469,N_16049);
nand U16610 (N_16610,N_16225,N_15471);
nor U16611 (N_16611,N_15659,N_15419);
nand U16612 (N_16612,N_15911,N_15136);
nand U16613 (N_16613,N_15681,N_15896);
and U16614 (N_16614,N_15535,N_15604);
or U16615 (N_16615,N_15919,N_16069);
and U16616 (N_16616,N_16283,N_15369);
or U16617 (N_16617,N_16458,N_16039);
and U16618 (N_16618,N_15940,N_16263);
or U16619 (N_16619,N_15807,N_16195);
nor U16620 (N_16620,N_16268,N_15135);
xnor U16621 (N_16621,N_15708,N_15966);
or U16622 (N_16622,N_15456,N_16350);
nor U16623 (N_16623,N_15898,N_16472);
and U16624 (N_16624,N_16332,N_15578);
xnor U16625 (N_16625,N_16037,N_15736);
and U16626 (N_16626,N_15537,N_15817);
xnor U16627 (N_16627,N_15145,N_15625);
and U16628 (N_16628,N_15816,N_16059);
nand U16629 (N_16629,N_15742,N_15702);
xnor U16630 (N_16630,N_15070,N_16426);
nor U16631 (N_16631,N_15310,N_15425);
nand U16632 (N_16632,N_15096,N_15961);
and U16633 (N_16633,N_16481,N_15198);
nand U16634 (N_16634,N_15391,N_16190);
and U16635 (N_16635,N_15109,N_15819);
nand U16636 (N_16636,N_15342,N_15461);
xnor U16637 (N_16637,N_15232,N_15914);
nor U16638 (N_16638,N_15167,N_15489);
xor U16639 (N_16639,N_16159,N_15378);
or U16640 (N_16640,N_15856,N_15576);
and U16641 (N_16641,N_16226,N_15030);
nor U16642 (N_16642,N_15148,N_15443);
or U16643 (N_16643,N_16079,N_16342);
nor U16644 (N_16644,N_15043,N_15854);
nor U16645 (N_16645,N_15622,N_16447);
xor U16646 (N_16646,N_16213,N_15841);
nor U16647 (N_16647,N_15068,N_15852);
nor U16648 (N_16648,N_15892,N_16154);
xor U16649 (N_16649,N_16437,N_15534);
nor U16650 (N_16650,N_16062,N_15507);
nand U16651 (N_16651,N_15714,N_15387);
nand U16652 (N_16652,N_16430,N_15108);
and U16653 (N_16653,N_15832,N_16205);
xnor U16654 (N_16654,N_15763,N_16365);
and U16655 (N_16655,N_15506,N_15906);
or U16656 (N_16656,N_16280,N_15306);
nor U16657 (N_16657,N_15293,N_16264);
or U16658 (N_16658,N_15959,N_15174);
nand U16659 (N_16659,N_16025,N_16197);
nor U16660 (N_16660,N_15648,N_15229);
xor U16661 (N_16661,N_16318,N_15023);
and U16662 (N_16662,N_15286,N_16301);
xnor U16663 (N_16663,N_16261,N_15051);
nand U16664 (N_16664,N_16252,N_15052);
xor U16665 (N_16665,N_15121,N_16192);
nand U16666 (N_16666,N_15531,N_15724);
nor U16667 (N_16667,N_15765,N_15631);
and U16668 (N_16668,N_15667,N_16298);
or U16669 (N_16669,N_16024,N_15549);
nor U16670 (N_16670,N_16007,N_16279);
and U16671 (N_16671,N_15099,N_15705);
and U16672 (N_16672,N_15581,N_16017);
and U16673 (N_16673,N_16081,N_15209);
xor U16674 (N_16674,N_16211,N_15600);
nand U16675 (N_16675,N_15778,N_15358);
and U16676 (N_16676,N_15389,N_15264);
nand U16677 (N_16677,N_15303,N_15676);
nand U16678 (N_16678,N_15196,N_15872);
nor U16679 (N_16679,N_15315,N_15054);
xor U16680 (N_16680,N_15104,N_15688);
nand U16681 (N_16681,N_16265,N_15545);
and U16682 (N_16682,N_16102,N_16450);
xnor U16683 (N_16683,N_15879,N_16156);
nand U16684 (N_16684,N_15007,N_16073);
nand U16685 (N_16685,N_16232,N_15572);
nand U16686 (N_16686,N_15032,N_16347);
nor U16687 (N_16687,N_15609,N_15755);
and U16688 (N_16688,N_15244,N_15147);
nand U16689 (N_16689,N_15496,N_16240);
nand U16690 (N_16690,N_16152,N_16194);
or U16691 (N_16691,N_15889,N_15027);
nand U16692 (N_16692,N_15322,N_15183);
nand U16693 (N_16693,N_15945,N_15729);
nand U16694 (N_16694,N_16216,N_16422);
nand U16695 (N_16695,N_15124,N_16137);
xnor U16696 (N_16696,N_16187,N_15610);
xnor U16697 (N_16697,N_16306,N_16003);
nor U16698 (N_16698,N_16484,N_15666);
nand U16699 (N_16699,N_15505,N_15077);
nand U16700 (N_16700,N_16063,N_16230);
nor U16701 (N_16701,N_15215,N_15668);
or U16702 (N_16702,N_16105,N_16076);
nor U16703 (N_16703,N_16398,N_15334);
nor U16704 (N_16704,N_15424,N_16035);
or U16705 (N_16705,N_15814,N_16057);
xor U16706 (N_16706,N_15927,N_15555);
and U16707 (N_16707,N_15712,N_16055);
and U16708 (N_16708,N_15573,N_16315);
nand U16709 (N_16709,N_15414,N_16064);
or U16710 (N_16710,N_15690,N_15563);
and U16711 (N_16711,N_16421,N_15181);
nand U16712 (N_16712,N_15723,N_16053);
xnor U16713 (N_16713,N_15818,N_16424);
nor U16714 (N_16714,N_15125,N_15162);
xnor U16715 (N_16715,N_15123,N_16255);
nand U16716 (N_16716,N_16352,N_16085);
nand U16717 (N_16717,N_16385,N_15787);
or U16718 (N_16718,N_15158,N_16429);
nor U16719 (N_16719,N_15815,N_16376);
nand U16720 (N_16720,N_15300,N_15877);
xor U16721 (N_16721,N_16207,N_15899);
and U16722 (N_16722,N_15432,N_15056);
or U16723 (N_16723,N_16050,N_15309);
and U16724 (N_16724,N_15155,N_16391);
nand U16725 (N_16725,N_16392,N_16319);
or U16726 (N_16726,N_16353,N_16041);
or U16727 (N_16727,N_16470,N_16351);
xnor U16728 (N_16728,N_16054,N_15466);
nand U16729 (N_16729,N_15113,N_15241);
nand U16730 (N_16730,N_15349,N_16191);
xor U16731 (N_16731,N_15627,N_15437);
and U16732 (N_16732,N_15242,N_16014);
nand U16733 (N_16733,N_16061,N_15771);
nor U16734 (N_16734,N_15640,N_15759);
and U16735 (N_16735,N_16312,N_15394);
xor U16736 (N_16736,N_15521,N_15482);
and U16737 (N_16737,N_15848,N_15981);
nand U16738 (N_16738,N_15130,N_15577);
or U16739 (N_16739,N_16082,N_15620);
nand U16740 (N_16740,N_15812,N_15483);
or U16741 (N_16741,N_16143,N_15891);
xor U16742 (N_16742,N_16258,N_15048);
or U16743 (N_16743,N_15448,N_15672);
nor U16744 (N_16744,N_15562,N_15773);
nand U16745 (N_16745,N_15663,N_15211);
nor U16746 (N_16746,N_15642,N_16224);
nor U16747 (N_16747,N_15713,N_15189);
or U16748 (N_16748,N_15655,N_15059);
nand U16749 (N_16749,N_16468,N_15341);
nor U16750 (N_16750,N_16141,N_16490);
xnor U16751 (N_16751,N_16498,N_15182);
nand U16752 (N_16752,N_16284,N_15833);
nor U16753 (N_16753,N_15318,N_16448);
and U16754 (N_16754,N_15415,N_15395);
xor U16755 (N_16755,N_16058,N_16174);
and U16756 (N_16756,N_16349,N_15754);
or U16757 (N_16757,N_16233,N_15268);
nand U16758 (N_16758,N_15159,N_16067);
and U16759 (N_16759,N_16158,N_15404);
nand U16760 (N_16760,N_15231,N_15844);
or U16761 (N_16761,N_15684,N_16310);
nand U16762 (N_16762,N_16248,N_16473);
or U16763 (N_16763,N_15074,N_15770);
or U16764 (N_16764,N_15287,N_15633);
nand U16765 (N_16765,N_15895,N_15295);
nor U16766 (N_16766,N_16042,N_16435);
or U16767 (N_16767,N_15883,N_15957);
nor U16768 (N_16768,N_15134,N_16030);
and U16769 (N_16769,N_15830,N_15887);
nor U16770 (N_16770,N_16320,N_16241);
or U16771 (N_16771,N_15863,N_15165);
or U16772 (N_16772,N_15792,N_16317);
xor U16773 (N_16773,N_15526,N_15963);
nand U16774 (N_16774,N_15776,N_16343);
nand U16775 (N_16775,N_15876,N_15091);
nor U16776 (N_16776,N_16489,N_15291);
nor U16777 (N_16777,N_15065,N_16486);
nand U16778 (N_16778,N_16243,N_15997);
xnor U16779 (N_16779,N_16123,N_16135);
xor U16780 (N_16780,N_15554,N_15233);
and U16781 (N_16781,N_16276,N_16387);
or U16782 (N_16782,N_15336,N_15343);
nand U16783 (N_16783,N_15031,N_15650);
or U16784 (N_16784,N_16170,N_15444);
nand U16785 (N_16785,N_15492,N_15079);
nand U16786 (N_16786,N_15979,N_16229);
nor U16787 (N_16787,N_16439,N_15447);
xor U16788 (N_16788,N_15741,N_16106);
xnor U16789 (N_16789,N_16210,N_15111);
and U16790 (N_16790,N_16001,N_15260);
nor U16791 (N_16791,N_16272,N_15612);
nand U16792 (N_16792,N_15421,N_15902);
and U16793 (N_16793,N_16220,N_15042);
or U16794 (N_16794,N_16221,N_16004);
nand U16795 (N_16795,N_16325,N_15410);
nor U16796 (N_16796,N_15700,N_15998);
or U16797 (N_16797,N_15055,N_15868);
nand U16798 (N_16798,N_15550,N_15200);
nor U16799 (N_16799,N_15384,N_15013);
and U16800 (N_16800,N_15457,N_16339);
xnor U16801 (N_16801,N_16436,N_16088);
xor U16802 (N_16802,N_15913,N_15772);
xor U16803 (N_16803,N_15463,N_16456);
and U16804 (N_16804,N_15875,N_15245);
nor U16805 (N_16805,N_15632,N_15995);
nand U16806 (N_16806,N_16031,N_15975);
xor U16807 (N_16807,N_15580,N_15462);
and U16808 (N_16808,N_15952,N_15946);
and U16809 (N_16809,N_15542,N_16374);
and U16810 (N_16810,N_15008,N_15500);
or U16811 (N_16811,N_16393,N_16333);
xor U16812 (N_16812,N_16324,N_15283);
xnor U16813 (N_16813,N_15847,N_15985);
xor U16814 (N_16814,N_16418,N_15970);
xnor U16815 (N_16815,N_16294,N_16269);
nor U16816 (N_16816,N_15499,N_15586);
or U16817 (N_16817,N_15485,N_15006);
and U16818 (N_16818,N_15380,N_16291);
and U16819 (N_16819,N_16452,N_16227);
xor U16820 (N_16820,N_15035,N_16104);
nor U16821 (N_16821,N_15210,N_15294);
or U16822 (N_16822,N_16427,N_15009);
or U16823 (N_16823,N_15405,N_15138);
nor U16824 (N_16824,N_16466,N_16487);
nor U16825 (N_16825,N_16383,N_15585);
or U16826 (N_16826,N_16462,N_15971);
or U16827 (N_16827,N_15552,N_15344);
xnor U16828 (N_16828,N_15439,N_15641);
or U16829 (N_16829,N_16474,N_16408);
xnor U16830 (N_16830,N_16433,N_16412);
nor U16831 (N_16831,N_15345,N_16395);
nor U16832 (N_16832,N_15105,N_15653);
nand U16833 (N_16833,N_15272,N_15441);
or U16834 (N_16834,N_15479,N_15078);
nor U16835 (N_16835,N_15335,N_15757);
and U16836 (N_16836,N_15219,N_15853);
xnor U16837 (N_16837,N_15594,N_16247);
and U16838 (N_16838,N_15643,N_15354);
nor U16839 (N_16839,N_15734,N_16250);
and U16840 (N_16840,N_15197,N_15163);
nand U16841 (N_16841,N_15004,N_15629);
and U16842 (N_16842,N_15599,N_15022);
xnor U16843 (N_16843,N_15122,N_16122);
xnor U16844 (N_16844,N_15703,N_15399);
nor U16845 (N_16845,N_16457,N_16371);
xor U16846 (N_16846,N_15273,N_15694);
and U16847 (N_16847,N_16464,N_16491);
nand U16848 (N_16848,N_15487,N_16471);
or U16849 (N_16849,N_16095,N_15278);
and U16850 (N_16850,N_15119,N_16378);
nor U16851 (N_16851,N_15346,N_15539);
nand U16852 (N_16852,N_15445,N_15908);
xnor U16853 (N_16853,N_16047,N_16345);
or U16854 (N_16854,N_15251,N_15558);
nor U16855 (N_16855,N_16425,N_15921);
nor U16856 (N_16856,N_15249,N_15731);
nand U16857 (N_16857,N_16316,N_16012);
nand U16858 (N_16858,N_15372,N_15860);
xnor U16859 (N_16859,N_15075,N_15098);
nor U16860 (N_16860,N_15715,N_15206);
and U16861 (N_16861,N_15630,N_15234);
and U16862 (N_16862,N_16311,N_16083);
nor U16863 (N_16863,N_16056,N_15187);
nand U16864 (N_16864,N_15598,N_16444);
or U16865 (N_16865,N_15192,N_16431);
nand U16866 (N_16866,N_15350,N_15393);
nand U16867 (N_16867,N_15353,N_15677);
nand U16868 (N_16868,N_16287,N_15525);
or U16869 (N_16869,N_15960,N_16293);
xor U16870 (N_16870,N_15403,N_15156);
nand U16871 (N_16871,N_16278,N_15811);
or U16872 (N_16872,N_16157,N_15636);
and U16873 (N_16873,N_16070,N_15169);
xor U16874 (N_16874,N_15368,N_16075);
and U16875 (N_16875,N_15989,N_15084);
xnor U16876 (N_16876,N_15988,N_15431);
nand U16877 (N_16877,N_15619,N_15925);
and U16878 (N_16878,N_15280,N_16087);
nor U16879 (N_16879,N_15230,N_15365);
nand U16880 (N_16880,N_15802,N_15157);
or U16881 (N_16881,N_15607,N_16377);
nand U16882 (N_16882,N_15646,N_15796);
and U16883 (N_16883,N_15137,N_16407);
nand U16884 (N_16884,N_15085,N_16397);
xor U16885 (N_16885,N_15289,N_15850);
and U16886 (N_16886,N_15514,N_15900);
or U16887 (N_16887,N_15276,N_15184);
nor U16888 (N_16888,N_15987,N_15011);
or U16889 (N_16889,N_16360,N_15304);
xnor U16890 (N_16890,N_15686,N_15467);
xnor U16891 (N_16891,N_15606,N_15978);
and U16892 (N_16892,N_16179,N_16358);
or U16893 (N_16893,N_15161,N_15279);
xnor U16894 (N_16894,N_16359,N_16417);
xnor U16895 (N_16895,N_15126,N_15449);
nand U16896 (N_16896,N_16124,N_15246);
or U16897 (N_16897,N_15566,N_15791);
xor U16898 (N_16898,N_15422,N_16008);
nor U16899 (N_16899,N_15769,N_15888);
nor U16900 (N_16900,N_15810,N_15869);
nand U16901 (N_16901,N_15588,N_15649);
nand U16902 (N_16902,N_15797,N_15266);
nor U16903 (N_16903,N_15095,N_16242);
xor U16904 (N_16904,N_16112,N_15865);
nor U16905 (N_16905,N_15408,N_16402);
xnor U16906 (N_16906,N_15579,N_15185);
and U16907 (N_16907,N_15180,N_15711);
nand U16908 (N_16908,N_15509,N_16267);
xor U16909 (N_16909,N_15478,N_16068);
nand U16910 (N_16910,N_15532,N_15319);
nor U16911 (N_16911,N_16184,N_16065);
nand U16912 (N_16912,N_15886,N_16071);
or U16913 (N_16913,N_15878,N_16344);
nor U16914 (N_16914,N_15005,N_16096);
or U16915 (N_16915,N_15753,N_15894);
or U16916 (N_16916,N_16228,N_15308);
or U16917 (N_16917,N_16091,N_16445);
nand U16918 (N_16918,N_15697,N_16022);
nor U16919 (N_16919,N_15223,N_15459);
nand U16920 (N_16920,N_15660,N_16322);
and U16921 (N_16921,N_15417,N_15784);
or U16922 (N_16922,N_15808,N_15258);
or U16923 (N_16923,N_15675,N_16423);
nand U16924 (N_16924,N_15110,N_16257);
xor U16925 (N_16925,N_15658,N_15076);
and U16926 (N_16926,N_15647,N_16361);
nand U16927 (N_16927,N_15806,N_15645);
nor U16928 (N_16928,N_15400,N_15502);
and U16929 (N_16929,N_16150,N_15665);
nor U16930 (N_16930,N_16175,N_16396);
nor U16931 (N_16931,N_15019,N_15347);
nor U16932 (N_16932,N_16405,N_15494);
nor U16933 (N_16933,N_15285,N_15382);
and U16934 (N_16934,N_16215,N_15779);
xor U16935 (N_16935,N_15476,N_15519);
nor U16936 (N_16936,N_16419,N_16127);
and U16937 (N_16937,N_16172,N_15786);
or U16938 (N_16938,N_16116,N_16256);
or U16939 (N_16939,N_15637,N_16134);
nor U16940 (N_16940,N_16441,N_15508);
and U16941 (N_16941,N_15840,N_15935);
xnor U16942 (N_16942,N_16090,N_16212);
xnor U16943 (N_16943,N_15568,N_16052);
nor U16944 (N_16944,N_16368,N_16132);
and U16945 (N_16945,N_15638,N_15440);
and U16946 (N_16946,N_15928,N_15758);
nor U16947 (N_16947,N_15948,N_15102);
or U16948 (N_16948,N_15528,N_15693);
nor U16949 (N_16949,N_15333,N_15118);
and U16950 (N_16950,N_16251,N_15885);
nor U16951 (N_16951,N_15379,N_15220);
nor U16952 (N_16952,N_15944,N_16440);
and U16953 (N_16953,N_15028,N_16161);
or U16954 (N_16954,N_15635,N_15904);
nor U16955 (N_16955,N_16148,N_15615);
or U16956 (N_16956,N_15396,N_15442);
nand U16957 (N_16957,N_16246,N_16499);
and U16958 (N_16958,N_15436,N_15926);
nor U16959 (N_16959,N_15761,N_15202);
or U16960 (N_16960,N_15129,N_15265);
or U16961 (N_16961,N_15081,N_16477);
nand U16962 (N_16962,N_15201,N_15057);
xor U16963 (N_16963,N_15247,N_15752);
nand U16964 (N_16964,N_16115,N_15533);
nor U16965 (N_16965,N_15803,N_15991);
nor U16966 (N_16966,N_15767,N_16262);
nand U16967 (N_16967,N_16416,N_15498);
nor U16968 (N_16968,N_15605,N_15942);
nand U16969 (N_16969,N_15170,N_15397);
nand U16970 (N_16970,N_15177,N_15058);
nor U16971 (N_16971,N_16219,N_16138);
xor U16972 (N_16972,N_15657,N_16036);
xnor U16973 (N_16973,N_16084,N_15790);
nand U16974 (N_16974,N_16144,N_15541);
xor U16975 (N_16975,N_16165,N_16066);
xor U16976 (N_16976,N_15617,N_16348);
or U16977 (N_16977,N_15331,N_15510);
nor U16978 (N_16978,N_16028,N_16290);
nand U16979 (N_16979,N_16411,N_15470);
nand U16980 (N_16980,N_15093,N_15616);
and U16981 (N_16981,N_15274,N_15142);
or U16982 (N_16982,N_16203,N_15548);
nor U16983 (N_16983,N_16176,N_15567);
xor U16984 (N_16984,N_15325,N_15039);
nand U16985 (N_16985,N_15253,N_16149);
nand U16986 (N_16986,N_15296,N_16340);
and U16987 (N_16987,N_15480,N_15326);
and U16988 (N_16988,N_15464,N_15839);
nand U16989 (N_16989,N_15140,N_15034);
or U16990 (N_16990,N_15016,N_16483);
xor U16991 (N_16991,N_15398,N_15809);
nor U16992 (N_16992,N_15813,N_15064);
nor U16993 (N_16993,N_15402,N_15259);
xor U16994 (N_16994,N_15149,N_15255);
and U16995 (N_16995,N_15082,N_15679);
nand U16996 (N_16996,N_15560,N_15002);
or U16997 (N_16997,N_15701,N_16119);
nand U16998 (N_16998,N_15915,N_15678);
xor U16999 (N_16999,N_16045,N_15529);
nor U17000 (N_17000,N_15569,N_16214);
and U17001 (N_17001,N_16113,N_15520);
nand U17002 (N_17002,N_15340,N_15024);
and U17003 (N_17003,N_15488,N_15021);
and U17004 (N_17004,N_15890,N_15312);
nand U17005 (N_17005,N_16098,N_15413);
and U17006 (N_17006,N_16126,N_15582);
nand U17007 (N_17007,N_15324,N_15683);
xor U17008 (N_17008,N_15313,N_15740);
or U17009 (N_17009,N_15117,N_16077);
nor U17010 (N_17010,N_15983,N_15618);
and U17011 (N_17011,N_15611,N_16494);
nand U17012 (N_17012,N_15608,N_15451);
nand U17013 (N_17013,N_15984,N_16118);
and U17014 (N_17014,N_15999,N_15112);
or U17015 (N_17015,N_16244,N_15366);
xnor U17016 (N_17016,N_16455,N_15407);
xnor U17017 (N_17017,N_16459,N_16307);
nor U17018 (N_17018,N_16334,N_16005);
nor U17019 (N_17019,N_15962,N_16182);
or U17020 (N_17020,N_16089,N_15994);
and U17021 (N_17021,N_16239,N_16326);
or U17022 (N_17022,N_15115,N_15951);
or U17023 (N_17023,N_16309,N_16355);
and U17024 (N_17024,N_16040,N_15912);
or U17025 (N_17025,N_16117,N_16259);
nand U17026 (N_17026,N_15955,N_16469);
nor U17027 (N_17027,N_15330,N_15922);
and U17028 (N_17028,N_15271,N_15873);
nor U17029 (N_17029,N_15386,N_15614);
nand U17030 (N_17030,N_16120,N_15361);
xnor U17031 (N_17031,N_15302,N_15406);
and U17032 (N_17032,N_15332,N_16401);
xnor U17033 (N_17033,N_15939,N_16223);
nor U17034 (N_17034,N_16094,N_15426);
xnor U17035 (N_17035,N_15428,N_15574);
nand U17036 (N_17036,N_16010,N_15725);
and U17037 (N_17037,N_16043,N_16357);
or U17038 (N_17038,N_15626,N_15929);
nand U17039 (N_17039,N_15152,N_16461);
nand U17040 (N_17040,N_15392,N_15072);
xor U17041 (N_17041,N_15938,N_16131);
nand U17042 (N_17042,N_15977,N_15909);
and U17043 (N_17043,N_15575,N_16364);
or U17044 (N_17044,N_15321,N_15427);
or U17045 (N_17045,N_15212,N_16140);
and U17046 (N_17046,N_15795,N_15652);
xnor U17047 (N_17047,N_15475,N_16480);
or U17048 (N_17048,N_15982,N_15739);
nor U17049 (N_17049,N_15825,N_16363);
nand U17050 (N_17050,N_15199,N_16373);
nor U17051 (N_17051,N_15565,N_15842);
and U17052 (N_17052,N_15297,N_15292);
nand U17053 (N_17053,N_16302,N_16453);
and U17054 (N_17054,N_15045,N_15941);
nand U17055 (N_17055,N_16204,N_15261);
xor U17056 (N_17056,N_15749,N_15050);
nor U17057 (N_17057,N_15069,N_16434);
nor U17058 (N_17058,N_16420,N_16281);
nand U17059 (N_17059,N_16020,N_15143);
or U17060 (N_17060,N_16409,N_16046);
nor U17061 (N_17061,N_15846,N_15804);
or U17062 (N_17062,N_15262,N_16467);
xor U17063 (N_17063,N_16254,N_16497);
or U17064 (N_17064,N_15281,N_16375);
nand U17065 (N_17065,N_15559,N_15682);
nand U17066 (N_17066,N_15544,N_15497);
or U17067 (N_17067,N_15743,N_15164);
or U17068 (N_17068,N_15556,N_16482);
nor U17069 (N_17069,N_16245,N_15821);
nor U17070 (N_17070,N_15680,N_16485);
nand U17071 (N_17071,N_15133,N_15766);
and U17072 (N_17072,N_15277,N_15884);
or U17073 (N_17073,N_15968,N_15762);
and U17074 (N_17074,N_15338,N_15750);
or U17075 (N_17075,N_15139,N_15047);
xnor U17076 (N_17076,N_15522,N_15671);
nand U17077 (N_17077,N_15829,N_15613);
xor U17078 (N_17078,N_15323,N_15178);
or U17079 (N_17079,N_16146,N_15204);
or U17080 (N_17080,N_15511,N_15317);
nand U17081 (N_17081,N_16234,N_16015);
xnor U17082 (N_17082,N_16372,N_15990);
or U17083 (N_17083,N_16454,N_15845);
nand U17084 (N_17084,N_16032,N_15747);
and U17085 (N_17085,N_16414,N_15867);
or U17086 (N_17086,N_16114,N_15299);
or U17087 (N_17087,N_16463,N_15094);
or U17088 (N_17088,N_16038,N_15870);
or U17089 (N_17089,N_15218,N_15307);
nor U17090 (N_17090,N_15822,N_16125);
and U17091 (N_17091,N_15592,N_15732);
xnor U17092 (N_17092,N_15623,N_15460);
and U17093 (N_17093,N_15018,N_15236);
nor U17094 (N_17094,N_15517,N_16389);
nand U17095 (N_17095,N_16169,N_15275);
or U17096 (N_17096,N_15001,N_16027);
or U17097 (N_17097,N_16222,N_15976);
or U17098 (N_17098,N_15217,N_15495);
nor U17099 (N_17099,N_15423,N_16330);
xor U17100 (N_17100,N_16415,N_16381);
nor U17101 (N_17101,N_16033,N_16188);
nand U17102 (N_17102,N_15716,N_15205);
xor U17103 (N_17103,N_15473,N_15651);
and U17104 (N_17104,N_15861,N_15301);
nor U17105 (N_17105,N_16495,N_15530);
or U17106 (N_17106,N_16162,N_15381);
or U17107 (N_17107,N_15858,N_16369);
xnor U17108 (N_17108,N_15964,N_15744);
or U17109 (N_17109,N_15673,N_16492);
and U17110 (N_17110,N_15969,N_15213);
or U17111 (N_17111,N_15864,N_16382);
nor U17112 (N_17112,N_15536,N_15698);
xnor U17113 (N_17113,N_15996,N_16253);
and U17114 (N_17114,N_15518,N_15947);
xnor U17115 (N_17115,N_15000,N_16139);
or U17116 (N_17116,N_15214,N_16410);
or U17117 (N_17117,N_15917,N_16136);
or U17118 (N_17118,N_16086,N_15515);
xnor U17119 (N_17119,N_15709,N_15768);
xnor U17120 (N_17120,N_15175,N_16390);
nand U17121 (N_17121,N_16173,N_15320);
xnor U17122 (N_17122,N_15362,N_15435);
and U17123 (N_17123,N_15429,N_15689);
nor U17124 (N_17124,N_15374,N_16078);
nor U17125 (N_17125,N_15662,N_16286);
or U17126 (N_17126,N_16413,N_16236);
xnor U17127 (N_17127,N_15359,N_15282);
xor U17128 (N_17128,N_16023,N_15760);
xnor U17129 (N_17129,N_16164,N_15687);
and U17130 (N_17130,N_15551,N_15144);
nand U17131 (N_17131,N_16018,N_16367);
or U17132 (N_17132,N_15730,N_15774);
or U17133 (N_17133,N_15491,N_15691);
nand U17134 (N_17134,N_16313,N_16166);
nand U17135 (N_17135,N_16366,N_15936);
xnor U17136 (N_17136,N_16288,N_15735);
xnor U17137 (N_17137,N_15493,N_15882);
nand U17138 (N_17138,N_16428,N_15015);
xnor U17139 (N_17139,N_15195,N_16362);
nor U17140 (N_17140,N_15474,N_16299);
and U17141 (N_17141,N_15593,N_15173);
or U17142 (N_17142,N_16449,N_16305);
nand U17143 (N_17143,N_16006,N_16155);
and U17144 (N_17144,N_15010,N_16271);
xnor U17145 (N_17145,N_15250,N_15067);
nand U17146 (N_17146,N_16107,N_15351);
nor U17147 (N_17147,N_15756,N_15418);
or U17148 (N_17148,N_15357,N_15040);
and U17149 (N_17149,N_15188,N_15061);
or U17150 (N_17150,N_15092,N_15628);
or U17151 (N_17151,N_15044,N_16274);
or U17152 (N_17152,N_16496,N_16237);
or U17153 (N_17153,N_15087,N_15931);
nor U17154 (N_17154,N_16328,N_15166);
or U17155 (N_17155,N_16493,N_15481);
xor U17156 (N_17156,N_15370,N_15799);
nor U17157 (N_17157,N_15706,N_15216);
and U17158 (N_17158,N_15707,N_16476);
xor U17159 (N_17159,N_15477,N_15154);
nor U17160 (N_17160,N_15973,N_16379);
xor U17161 (N_17161,N_16109,N_15248);
and U17162 (N_17162,N_16128,N_16403);
or U17163 (N_17163,N_15965,N_15543);
xor U17164 (N_17164,N_16442,N_16198);
or U17165 (N_17165,N_15800,N_15933);
nand U17166 (N_17166,N_15420,N_15383);
nand U17167 (N_17167,N_15835,N_15897);
or U17168 (N_17168,N_15046,N_15674);
and U17169 (N_17169,N_15937,N_16177);
or U17170 (N_17170,N_15454,N_16209);
nor U17171 (N_17171,N_15207,N_15401);
nor U17172 (N_17172,N_15385,N_15458);
xor U17173 (N_17173,N_15512,N_15311);
xnor U17174 (N_17174,N_16235,N_15777);
or U17175 (N_17175,N_15624,N_15252);
xor U17176 (N_17176,N_15639,N_16296);
nor U17177 (N_17177,N_16354,N_15584);
nor U17178 (N_17178,N_15367,N_15168);
or U17179 (N_17179,N_15603,N_15452);
and U17180 (N_17180,N_16110,N_16180);
nand U17181 (N_17181,N_16133,N_15172);
and U17182 (N_17182,N_15080,N_15923);
and U17183 (N_17183,N_15664,N_15097);
nor U17184 (N_17184,N_15026,N_15656);
nand U17185 (N_17185,N_15516,N_15017);
and U17186 (N_17186,N_15801,N_15465);
xnor U17187 (N_17187,N_15557,N_15857);
nor U17188 (N_17188,N_15932,N_15171);
xor U17189 (N_17189,N_15412,N_15239);
xnor U17190 (N_17190,N_16337,N_15041);
and U17191 (N_17191,N_15595,N_15254);
and U17192 (N_17192,N_16206,N_15036);
xnor U17193 (N_17193,N_16341,N_16103);
xor U17194 (N_17194,N_15227,N_15160);
or U17195 (N_17195,N_15589,N_15235);
and U17196 (N_17196,N_15597,N_15132);
nor U17197 (N_17197,N_15727,N_15838);
nor U17198 (N_17198,N_15738,N_15438);
and U17199 (N_17199,N_16160,N_15455);
nand U17200 (N_17200,N_15356,N_15793);
or U17201 (N_17201,N_15388,N_16202);
nand U17202 (N_17202,N_15194,N_15775);
xor U17203 (N_17203,N_15176,N_16338);
xnor U17204 (N_17204,N_15151,N_16275);
nand U17205 (N_17205,N_16178,N_15430);
xnor U17206 (N_17206,N_15453,N_15924);
and U17207 (N_17207,N_15025,N_15339);
or U17208 (N_17208,N_16074,N_15416);
xor U17209 (N_17209,N_15881,N_16201);
nand U17210 (N_17210,N_15805,N_16013);
xor U17211 (N_17211,N_16249,N_15053);
nor U17212 (N_17212,N_15305,N_15446);
or U17213 (N_17213,N_15986,N_16314);
and U17214 (N_17214,N_15855,N_15745);
or U17215 (N_17215,N_15226,N_15490);
or U17216 (N_17216,N_15871,N_16021);
nor U17217 (N_17217,N_15150,N_16475);
and U17218 (N_17218,N_16438,N_15874);
nor U17219 (N_17219,N_15943,N_15073);
and U17220 (N_17220,N_15596,N_15089);
or U17221 (N_17221,N_15930,N_16167);
nand U17222 (N_17222,N_15003,N_16200);
nor U17223 (N_17223,N_15564,N_15956);
and U17224 (N_17224,N_15033,N_15256);
and U17225 (N_17225,N_15037,N_15012);
and U17226 (N_17226,N_16009,N_15621);
xnor U17227 (N_17227,N_16044,N_15193);
nand U17228 (N_17228,N_16099,N_15880);
xor U17229 (N_17229,N_15486,N_15411);
xor U17230 (N_17230,N_15571,N_15141);
xnor U17231 (N_17231,N_16186,N_15355);
or U17232 (N_17232,N_15371,N_15746);
or U17233 (N_17233,N_15360,N_16092);
nand U17234 (N_17234,N_16394,N_15062);
xor U17235 (N_17235,N_16285,N_15208);
xor U17236 (N_17236,N_16465,N_15106);
nand U17237 (N_17237,N_15376,N_16386);
and U17238 (N_17238,N_16048,N_15377);
or U17239 (N_17239,N_15146,N_15224);
nand U17240 (N_17240,N_15591,N_15954);
and U17241 (N_17241,N_15949,N_15901);
nand U17242 (N_17242,N_16323,N_16388);
and U17243 (N_17243,N_15468,N_15337);
nand U17244 (N_17244,N_15794,N_15523);
nor U17245 (N_17245,N_15893,N_15131);
and U17246 (N_17246,N_15590,N_15866);
nor U17247 (N_17247,N_15862,N_15269);
nand U17248 (N_17248,N_16185,N_15670);
nor U17249 (N_17249,N_15038,N_15827);
or U17250 (N_17250,N_15157,N_16473);
nor U17251 (N_17251,N_16012,N_15256);
nand U17252 (N_17252,N_15204,N_15085);
xor U17253 (N_17253,N_16194,N_16070);
nor U17254 (N_17254,N_15303,N_15654);
xnor U17255 (N_17255,N_15889,N_15691);
xor U17256 (N_17256,N_15606,N_16421);
nor U17257 (N_17257,N_16489,N_15538);
xnor U17258 (N_17258,N_15621,N_15708);
xor U17259 (N_17259,N_16209,N_15705);
and U17260 (N_17260,N_16034,N_16340);
nor U17261 (N_17261,N_16301,N_16023);
or U17262 (N_17262,N_16190,N_16287);
and U17263 (N_17263,N_15958,N_15122);
xor U17264 (N_17264,N_16081,N_15048);
nor U17265 (N_17265,N_15040,N_15714);
or U17266 (N_17266,N_15721,N_15039);
and U17267 (N_17267,N_15572,N_15167);
and U17268 (N_17268,N_15079,N_15357);
and U17269 (N_17269,N_15456,N_15246);
xnor U17270 (N_17270,N_16058,N_15933);
or U17271 (N_17271,N_15443,N_16224);
xnor U17272 (N_17272,N_16495,N_16028);
and U17273 (N_17273,N_15635,N_15606);
xor U17274 (N_17274,N_16288,N_16434);
xnor U17275 (N_17275,N_15080,N_15836);
xnor U17276 (N_17276,N_16086,N_15998);
or U17277 (N_17277,N_16166,N_15677);
xor U17278 (N_17278,N_16108,N_15911);
xnor U17279 (N_17279,N_16131,N_16291);
or U17280 (N_17280,N_16156,N_16151);
xor U17281 (N_17281,N_16349,N_16087);
xnor U17282 (N_17282,N_15633,N_15202);
nand U17283 (N_17283,N_15968,N_15638);
nor U17284 (N_17284,N_15467,N_15817);
nor U17285 (N_17285,N_16459,N_16078);
nor U17286 (N_17286,N_15418,N_16431);
xnor U17287 (N_17287,N_16388,N_15677);
nor U17288 (N_17288,N_16311,N_16339);
nand U17289 (N_17289,N_15909,N_15844);
nand U17290 (N_17290,N_16394,N_15378);
and U17291 (N_17291,N_15455,N_16022);
and U17292 (N_17292,N_16399,N_15598);
or U17293 (N_17293,N_15029,N_16143);
or U17294 (N_17294,N_16269,N_16455);
xor U17295 (N_17295,N_16140,N_15453);
xnor U17296 (N_17296,N_15838,N_16477);
xnor U17297 (N_17297,N_15462,N_16365);
nor U17298 (N_17298,N_16109,N_15708);
and U17299 (N_17299,N_16346,N_16106);
xnor U17300 (N_17300,N_15863,N_15614);
or U17301 (N_17301,N_15589,N_16321);
nor U17302 (N_17302,N_16493,N_15709);
or U17303 (N_17303,N_15247,N_15519);
nand U17304 (N_17304,N_15810,N_16354);
or U17305 (N_17305,N_16178,N_15115);
and U17306 (N_17306,N_16286,N_16412);
nor U17307 (N_17307,N_16274,N_16481);
nor U17308 (N_17308,N_16054,N_15916);
and U17309 (N_17309,N_15554,N_15944);
nor U17310 (N_17310,N_15432,N_15406);
nand U17311 (N_17311,N_15863,N_15088);
nor U17312 (N_17312,N_15093,N_16170);
or U17313 (N_17313,N_16035,N_15643);
xor U17314 (N_17314,N_15808,N_15098);
nor U17315 (N_17315,N_16068,N_16186);
nand U17316 (N_17316,N_15481,N_15981);
and U17317 (N_17317,N_16092,N_16266);
or U17318 (N_17318,N_16260,N_16266);
and U17319 (N_17319,N_15831,N_16089);
and U17320 (N_17320,N_15949,N_15187);
and U17321 (N_17321,N_15997,N_16344);
and U17322 (N_17322,N_16074,N_15932);
and U17323 (N_17323,N_15456,N_16018);
nand U17324 (N_17324,N_15114,N_16471);
or U17325 (N_17325,N_16465,N_15052);
xor U17326 (N_17326,N_16205,N_15901);
xnor U17327 (N_17327,N_16476,N_15997);
xnor U17328 (N_17328,N_15693,N_15073);
nand U17329 (N_17329,N_15618,N_15302);
nand U17330 (N_17330,N_15502,N_15288);
nor U17331 (N_17331,N_16369,N_15640);
xor U17332 (N_17332,N_16377,N_15777);
or U17333 (N_17333,N_16467,N_15931);
xor U17334 (N_17334,N_15234,N_16451);
or U17335 (N_17335,N_16207,N_15800);
nor U17336 (N_17336,N_15573,N_15669);
nor U17337 (N_17337,N_15118,N_15237);
or U17338 (N_17338,N_15636,N_16106);
and U17339 (N_17339,N_16178,N_16124);
nor U17340 (N_17340,N_15712,N_16239);
nor U17341 (N_17341,N_16186,N_15050);
or U17342 (N_17342,N_16196,N_16036);
nand U17343 (N_17343,N_16417,N_15363);
or U17344 (N_17344,N_16077,N_15550);
xor U17345 (N_17345,N_16064,N_15311);
nand U17346 (N_17346,N_15566,N_15772);
and U17347 (N_17347,N_16305,N_16161);
nor U17348 (N_17348,N_16011,N_16473);
or U17349 (N_17349,N_16443,N_16113);
nor U17350 (N_17350,N_15107,N_15759);
or U17351 (N_17351,N_16441,N_16237);
nand U17352 (N_17352,N_15778,N_16183);
xor U17353 (N_17353,N_15258,N_15946);
xor U17354 (N_17354,N_15947,N_15551);
or U17355 (N_17355,N_16305,N_15956);
xnor U17356 (N_17356,N_15695,N_15268);
xor U17357 (N_17357,N_15232,N_15843);
xnor U17358 (N_17358,N_16155,N_16423);
and U17359 (N_17359,N_15819,N_15278);
and U17360 (N_17360,N_15931,N_15803);
nand U17361 (N_17361,N_16144,N_15116);
nor U17362 (N_17362,N_15111,N_15732);
nor U17363 (N_17363,N_15603,N_15235);
or U17364 (N_17364,N_15814,N_15481);
nor U17365 (N_17365,N_15652,N_15941);
nand U17366 (N_17366,N_15884,N_15974);
or U17367 (N_17367,N_15368,N_15309);
and U17368 (N_17368,N_15479,N_15785);
or U17369 (N_17369,N_15611,N_15172);
xor U17370 (N_17370,N_15086,N_16075);
or U17371 (N_17371,N_16131,N_15343);
nor U17372 (N_17372,N_15591,N_15499);
or U17373 (N_17373,N_15905,N_15490);
nor U17374 (N_17374,N_15014,N_15987);
xor U17375 (N_17375,N_15970,N_15306);
and U17376 (N_17376,N_15927,N_15887);
and U17377 (N_17377,N_16341,N_15867);
and U17378 (N_17378,N_15174,N_15250);
and U17379 (N_17379,N_16036,N_15197);
nor U17380 (N_17380,N_15300,N_16329);
nand U17381 (N_17381,N_15618,N_15078);
xor U17382 (N_17382,N_15372,N_15963);
nand U17383 (N_17383,N_15927,N_15827);
nor U17384 (N_17384,N_16307,N_15178);
and U17385 (N_17385,N_15641,N_15792);
nand U17386 (N_17386,N_15908,N_15967);
xor U17387 (N_17387,N_16158,N_15245);
nor U17388 (N_17388,N_15605,N_15037);
nand U17389 (N_17389,N_15801,N_15296);
nor U17390 (N_17390,N_15140,N_15100);
or U17391 (N_17391,N_16155,N_16139);
nor U17392 (N_17392,N_16472,N_15858);
xnor U17393 (N_17393,N_16454,N_15864);
or U17394 (N_17394,N_16063,N_16175);
or U17395 (N_17395,N_15547,N_15177);
or U17396 (N_17396,N_15863,N_15623);
or U17397 (N_17397,N_16088,N_16461);
or U17398 (N_17398,N_15293,N_16086);
or U17399 (N_17399,N_15134,N_16228);
and U17400 (N_17400,N_15701,N_16174);
or U17401 (N_17401,N_15174,N_15194);
and U17402 (N_17402,N_15144,N_16438);
or U17403 (N_17403,N_15526,N_15278);
or U17404 (N_17404,N_15274,N_15824);
xor U17405 (N_17405,N_15530,N_15845);
and U17406 (N_17406,N_15749,N_15349);
or U17407 (N_17407,N_15871,N_15465);
and U17408 (N_17408,N_15539,N_15195);
nor U17409 (N_17409,N_15231,N_16384);
xor U17410 (N_17410,N_15302,N_15928);
or U17411 (N_17411,N_15887,N_15494);
nor U17412 (N_17412,N_15389,N_15557);
or U17413 (N_17413,N_16472,N_16279);
and U17414 (N_17414,N_15366,N_15627);
or U17415 (N_17415,N_15123,N_16095);
nand U17416 (N_17416,N_15320,N_16068);
xnor U17417 (N_17417,N_15476,N_15154);
and U17418 (N_17418,N_16033,N_16201);
xor U17419 (N_17419,N_15876,N_16467);
xnor U17420 (N_17420,N_15916,N_15662);
and U17421 (N_17421,N_15512,N_16389);
xnor U17422 (N_17422,N_16066,N_16186);
nor U17423 (N_17423,N_15769,N_15696);
nand U17424 (N_17424,N_15443,N_16286);
nor U17425 (N_17425,N_15897,N_15552);
xnor U17426 (N_17426,N_16020,N_15797);
nor U17427 (N_17427,N_16308,N_15932);
nand U17428 (N_17428,N_15791,N_15780);
xnor U17429 (N_17429,N_16228,N_16455);
and U17430 (N_17430,N_15760,N_15882);
nor U17431 (N_17431,N_15815,N_16124);
xnor U17432 (N_17432,N_15605,N_16106);
xnor U17433 (N_17433,N_16370,N_16336);
and U17434 (N_17434,N_15242,N_15436);
nor U17435 (N_17435,N_15532,N_16440);
nor U17436 (N_17436,N_15783,N_15467);
nand U17437 (N_17437,N_16427,N_15073);
nand U17438 (N_17438,N_15517,N_15040);
nor U17439 (N_17439,N_15477,N_15638);
nor U17440 (N_17440,N_15914,N_15310);
xor U17441 (N_17441,N_16397,N_16229);
xor U17442 (N_17442,N_15019,N_15325);
xor U17443 (N_17443,N_16222,N_15728);
or U17444 (N_17444,N_15106,N_16271);
nor U17445 (N_17445,N_16253,N_15118);
nand U17446 (N_17446,N_15415,N_15580);
xor U17447 (N_17447,N_15098,N_16359);
and U17448 (N_17448,N_15001,N_16120);
or U17449 (N_17449,N_15526,N_16161);
xor U17450 (N_17450,N_16192,N_15539);
and U17451 (N_17451,N_16330,N_15097);
xnor U17452 (N_17452,N_15737,N_16201);
nor U17453 (N_17453,N_15492,N_16436);
xor U17454 (N_17454,N_15813,N_15689);
nor U17455 (N_17455,N_16474,N_15367);
and U17456 (N_17456,N_15953,N_16007);
nand U17457 (N_17457,N_15935,N_16268);
or U17458 (N_17458,N_16134,N_15091);
or U17459 (N_17459,N_16312,N_15678);
nand U17460 (N_17460,N_15447,N_15871);
and U17461 (N_17461,N_15805,N_15179);
nand U17462 (N_17462,N_15507,N_15347);
and U17463 (N_17463,N_15960,N_15528);
xnor U17464 (N_17464,N_15456,N_16152);
nand U17465 (N_17465,N_15476,N_15640);
and U17466 (N_17466,N_15111,N_15901);
and U17467 (N_17467,N_16469,N_15125);
nor U17468 (N_17468,N_16242,N_16438);
xor U17469 (N_17469,N_15682,N_15148);
xor U17470 (N_17470,N_15644,N_16189);
or U17471 (N_17471,N_15590,N_16437);
and U17472 (N_17472,N_16148,N_15513);
nor U17473 (N_17473,N_15946,N_16425);
nand U17474 (N_17474,N_16416,N_15763);
xnor U17475 (N_17475,N_15961,N_16432);
xnor U17476 (N_17476,N_15336,N_15189);
nor U17477 (N_17477,N_15175,N_15143);
nand U17478 (N_17478,N_15681,N_16088);
nor U17479 (N_17479,N_15683,N_15156);
and U17480 (N_17480,N_15166,N_15203);
xor U17481 (N_17481,N_15003,N_15651);
nand U17482 (N_17482,N_15578,N_15150);
xor U17483 (N_17483,N_16268,N_15989);
and U17484 (N_17484,N_16017,N_15387);
nor U17485 (N_17485,N_15377,N_16397);
xor U17486 (N_17486,N_15151,N_15552);
and U17487 (N_17487,N_15110,N_15225);
xnor U17488 (N_17488,N_15509,N_16099);
and U17489 (N_17489,N_15935,N_16113);
xor U17490 (N_17490,N_15859,N_16233);
or U17491 (N_17491,N_15883,N_15328);
or U17492 (N_17492,N_15192,N_16160);
nor U17493 (N_17493,N_15862,N_16341);
xnor U17494 (N_17494,N_15409,N_16062);
and U17495 (N_17495,N_16249,N_15993);
nand U17496 (N_17496,N_15128,N_15101);
or U17497 (N_17497,N_15233,N_15249);
nor U17498 (N_17498,N_15088,N_15013);
xnor U17499 (N_17499,N_15243,N_16295);
xor U17500 (N_17500,N_15427,N_16021);
nand U17501 (N_17501,N_15444,N_16446);
nor U17502 (N_17502,N_16137,N_16002);
xnor U17503 (N_17503,N_15457,N_15041);
nor U17504 (N_17504,N_15796,N_16324);
or U17505 (N_17505,N_15014,N_16265);
xnor U17506 (N_17506,N_15371,N_15957);
and U17507 (N_17507,N_15247,N_15107);
nand U17508 (N_17508,N_16364,N_15109);
xor U17509 (N_17509,N_16120,N_15128);
nor U17510 (N_17510,N_15059,N_16478);
xnor U17511 (N_17511,N_16410,N_16069);
or U17512 (N_17512,N_15072,N_15027);
nand U17513 (N_17513,N_15589,N_15297);
nor U17514 (N_17514,N_15230,N_15135);
nor U17515 (N_17515,N_15228,N_15729);
nand U17516 (N_17516,N_16473,N_16099);
or U17517 (N_17517,N_15661,N_16357);
and U17518 (N_17518,N_15845,N_16281);
nor U17519 (N_17519,N_16420,N_15335);
and U17520 (N_17520,N_15318,N_15606);
nor U17521 (N_17521,N_15634,N_15825);
nand U17522 (N_17522,N_16385,N_15122);
xor U17523 (N_17523,N_15056,N_15937);
and U17524 (N_17524,N_16143,N_16151);
and U17525 (N_17525,N_16279,N_15490);
xor U17526 (N_17526,N_15893,N_16107);
nor U17527 (N_17527,N_15526,N_16309);
nand U17528 (N_17528,N_15979,N_15866);
and U17529 (N_17529,N_16363,N_15009);
and U17530 (N_17530,N_15380,N_16283);
nand U17531 (N_17531,N_15133,N_15065);
nand U17532 (N_17532,N_16264,N_15398);
nand U17533 (N_17533,N_15117,N_15687);
and U17534 (N_17534,N_15966,N_15692);
nor U17535 (N_17535,N_15669,N_15342);
nor U17536 (N_17536,N_16180,N_16497);
and U17537 (N_17537,N_15896,N_16388);
xor U17538 (N_17538,N_16143,N_16482);
nor U17539 (N_17539,N_15376,N_16153);
xor U17540 (N_17540,N_15576,N_15757);
nand U17541 (N_17541,N_15096,N_16134);
or U17542 (N_17542,N_15486,N_15502);
xnor U17543 (N_17543,N_16148,N_16031);
xor U17544 (N_17544,N_15200,N_15395);
or U17545 (N_17545,N_16052,N_16241);
nand U17546 (N_17546,N_16080,N_15821);
and U17547 (N_17547,N_15486,N_15796);
nand U17548 (N_17548,N_15067,N_15068);
nor U17549 (N_17549,N_16241,N_15059);
and U17550 (N_17550,N_16435,N_16085);
or U17551 (N_17551,N_16243,N_15076);
and U17552 (N_17552,N_15425,N_15796);
and U17553 (N_17553,N_15688,N_15750);
nor U17554 (N_17554,N_16356,N_15819);
nand U17555 (N_17555,N_15079,N_15637);
nor U17556 (N_17556,N_16346,N_15843);
xnor U17557 (N_17557,N_16032,N_15138);
or U17558 (N_17558,N_15419,N_16484);
or U17559 (N_17559,N_15384,N_16021);
and U17560 (N_17560,N_15518,N_15976);
or U17561 (N_17561,N_16344,N_16155);
xnor U17562 (N_17562,N_16321,N_15956);
and U17563 (N_17563,N_15821,N_15954);
and U17564 (N_17564,N_15002,N_15556);
xnor U17565 (N_17565,N_15048,N_15684);
nand U17566 (N_17566,N_15609,N_16151);
and U17567 (N_17567,N_15758,N_15769);
and U17568 (N_17568,N_15970,N_15037);
xor U17569 (N_17569,N_15758,N_15526);
xor U17570 (N_17570,N_16446,N_15808);
and U17571 (N_17571,N_16199,N_16015);
and U17572 (N_17572,N_15288,N_15109);
and U17573 (N_17573,N_15676,N_15855);
xor U17574 (N_17574,N_15251,N_15886);
xnor U17575 (N_17575,N_16410,N_15500);
nor U17576 (N_17576,N_15289,N_15505);
or U17577 (N_17577,N_15399,N_15769);
and U17578 (N_17578,N_16014,N_16498);
nor U17579 (N_17579,N_16418,N_15030);
nand U17580 (N_17580,N_15210,N_15104);
xor U17581 (N_17581,N_15447,N_15356);
nand U17582 (N_17582,N_15264,N_16062);
or U17583 (N_17583,N_15582,N_16246);
and U17584 (N_17584,N_15951,N_16204);
nor U17585 (N_17585,N_15200,N_15672);
nand U17586 (N_17586,N_15317,N_16494);
nand U17587 (N_17587,N_15949,N_16080);
nor U17588 (N_17588,N_15674,N_15763);
xor U17589 (N_17589,N_15571,N_16375);
nor U17590 (N_17590,N_16184,N_15132);
xnor U17591 (N_17591,N_15246,N_15596);
or U17592 (N_17592,N_16158,N_15906);
and U17593 (N_17593,N_16226,N_15073);
xnor U17594 (N_17594,N_15072,N_16349);
nor U17595 (N_17595,N_16410,N_16063);
xor U17596 (N_17596,N_15088,N_15382);
nor U17597 (N_17597,N_15541,N_16418);
xnor U17598 (N_17598,N_16399,N_16042);
xor U17599 (N_17599,N_15926,N_15745);
xnor U17600 (N_17600,N_16379,N_15495);
nand U17601 (N_17601,N_15600,N_16487);
xnor U17602 (N_17602,N_15591,N_16352);
or U17603 (N_17603,N_15440,N_15135);
and U17604 (N_17604,N_15399,N_15402);
xnor U17605 (N_17605,N_16179,N_16211);
xnor U17606 (N_17606,N_15124,N_15139);
and U17607 (N_17607,N_15580,N_16227);
and U17608 (N_17608,N_15649,N_15766);
xnor U17609 (N_17609,N_15460,N_15281);
xor U17610 (N_17610,N_15794,N_15719);
xnor U17611 (N_17611,N_16089,N_16269);
or U17612 (N_17612,N_16250,N_15486);
nor U17613 (N_17613,N_15787,N_16404);
nor U17614 (N_17614,N_15128,N_16458);
nor U17615 (N_17615,N_15484,N_15581);
and U17616 (N_17616,N_16021,N_16363);
xnor U17617 (N_17617,N_15258,N_15607);
xnor U17618 (N_17618,N_16475,N_16478);
or U17619 (N_17619,N_15375,N_15628);
or U17620 (N_17620,N_16285,N_16240);
xor U17621 (N_17621,N_15827,N_15982);
xor U17622 (N_17622,N_16471,N_16204);
and U17623 (N_17623,N_15681,N_16372);
nand U17624 (N_17624,N_16407,N_16492);
xnor U17625 (N_17625,N_16398,N_15834);
nor U17626 (N_17626,N_16404,N_15953);
or U17627 (N_17627,N_16037,N_15802);
xor U17628 (N_17628,N_15945,N_16241);
or U17629 (N_17629,N_15050,N_15635);
xor U17630 (N_17630,N_15028,N_15212);
xnor U17631 (N_17631,N_15235,N_16065);
nor U17632 (N_17632,N_16295,N_15938);
and U17633 (N_17633,N_16181,N_15642);
nand U17634 (N_17634,N_16309,N_15102);
nand U17635 (N_17635,N_16492,N_15013);
or U17636 (N_17636,N_15120,N_15480);
or U17637 (N_17637,N_16400,N_15573);
xnor U17638 (N_17638,N_15982,N_16049);
nor U17639 (N_17639,N_15195,N_16446);
nor U17640 (N_17640,N_16486,N_15050);
and U17641 (N_17641,N_15905,N_15629);
nand U17642 (N_17642,N_15726,N_15272);
or U17643 (N_17643,N_15367,N_15604);
or U17644 (N_17644,N_16131,N_15178);
nand U17645 (N_17645,N_16416,N_15230);
nor U17646 (N_17646,N_15593,N_16055);
or U17647 (N_17647,N_15799,N_15037);
nand U17648 (N_17648,N_15715,N_15252);
nand U17649 (N_17649,N_16277,N_15171);
xnor U17650 (N_17650,N_15603,N_16301);
or U17651 (N_17651,N_15048,N_15180);
nand U17652 (N_17652,N_16291,N_16071);
nand U17653 (N_17653,N_15096,N_15053);
nor U17654 (N_17654,N_16418,N_15561);
nor U17655 (N_17655,N_15225,N_15352);
nor U17656 (N_17656,N_15827,N_15943);
and U17657 (N_17657,N_15018,N_15711);
nor U17658 (N_17658,N_15477,N_16487);
or U17659 (N_17659,N_15051,N_15111);
or U17660 (N_17660,N_15316,N_15419);
and U17661 (N_17661,N_15167,N_15555);
nand U17662 (N_17662,N_15601,N_15870);
nand U17663 (N_17663,N_15933,N_15184);
xor U17664 (N_17664,N_16237,N_16420);
nor U17665 (N_17665,N_15346,N_16442);
xor U17666 (N_17666,N_15447,N_16256);
nor U17667 (N_17667,N_15296,N_15934);
xnor U17668 (N_17668,N_15618,N_16346);
xor U17669 (N_17669,N_16356,N_15214);
or U17670 (N_17670,N_15154,N_15720);
nor U17671 (N_17671,N_15037,N_15232);
or U17672 (N_17672,N_15690,N_15585);
nand U17673 (N_17673,N_16289,N_15231);
and U17674 (N_17674,N_15945,N_15511);
xor U17675 (N_17675,N_15452,N_15257);
xor U17676 (N_17676,N_15316,N_15425);
xor U17677 (N_17677,N_15043,N_16108);
or U17678 (N_17678,N_15502,N_16263);
or U17679 (N_17679,N_16293,N_15500);
xor U17680 (N_17680,N_15549,N_15147);
and U17681 (N_17681,N_15682,N_15667);
nand U17682 (N_17682,N_15570,N_16434);
nor U17683 (N_17683,N_15248,N_15035);
nand U17684 (N_17684,N_16137,N_15357);
and U17685 (N_17685,N_15754,N_15951);
nor U17686 (N_17686,N_16493,N_15448);
nand U17687 (N_17687,N_16187,N_15937);
nand U17688 (N_17688,N_16297,N_15767);
xor U17689 (N_17689,N_15117,N_16439);
nor U17690 (N_17690,N_15887,N_15776);
nand U17691 (N_17691,N_16464,N_15295);
and U17692 (N_17692,N_16425,N_16134);
xor U17693 (N_17693,N_16381,N_16493);
or U17694 (N_17694,N_15943,N_16057);
nand U17695 (N_17695,N_15811,N_15026);
xor U17696 (N_17696,N_15807,N_16079);
xnor U17697 (N_17697,N_15265,N_15049);
and U17698 (N_17698,N_15131,N_16226);
nor U17699 (N_17699,N_15892,N_16146);
nand U17700 (N_17700,N_15758,N_15112);
xnor U17701 (N_17701,N_15701,N_15081);
nand U17702 (N_17702,N_15854,N_16249);
nand U17703 (N_17703,N_15631,N_15455);
nor U17704 (N_17704,N_16084,N_15108);
and U17705 (N_17705,N_15931,N_15094);
nor U17706 (N_17706,N_15051,N_15215);
nand U17707 (N_17707,N_15178,N_15239);
xor U17708 (N_17708,N_16390,N_16075);
and U17709 (N_17709,N_15694,N_16143);
and U17710 (N_17710,N_15554,N_15481);
nand U17711 (N_17711,N_15673,N_15257);
nor U17712 (N_17712,N_15667,N_15950);
nor U17713 (N_17713,N_16363,N_15477);
xor U17714 (N_17714,N_15073,N_15944);
xor U17715 (N_17715,N_15210,N_15791);
nand U17716 (N_17716,N_15737,N_15833);
xor U17717 (N_17717,N_15077,N_15995);
and U17718 (N_17718,N_16407,N_16173);
and U17719 (N_17719,N_15183,N_15435);
and U17720 (N_17720,N_16268,N_15381);
and U17721 (N_17721,N_15185,N_15331);
xnor U17722 (N_17722,N_16234,N_16402);
nand U17723 (N_17723,N_15602,N_16276);
and U17724 (N_17724,N_15307,N_16488);
nor U17725 (N_17725,N_15981,N_15823);
or U17726 (N_17726,N_16297,N_16331);
and U17727 (N_17727,N_15890,N_15946);
nor U17728 (N_17728,N_15130,N_15746);
xnor U17729 (N_17729,N_15585,N_15843);
xnor U17730 (N_17730,N_15558,N_15517);
and U17731 (N_17731,N_15733,N_15721);
nor U17732 (N_17732,N_15337,N_15243);
and U17733 (N_17733,N_15301,N_15299);
xnor U17734 (N_17734,N_16057,N_15995);
nor U17735 (N_17735,N_16464,N_16334);
xnor U17736 (N_17736,N_15087,N_15520);
or U17737 (N_17737,N_15655,N_15167);
xnor U17738 (N_17738,N_15313,N_15966);
nor U17739 (N_17739,N_15611,N_16154);
xor U17740 (N_17740,N_15383,N_16240);
nand U17741 (N_17741,N_15473,N_15627);
and U17742 (N_17742,N_15177,N_15943);
xor U17743 (N_17743,N_15764,N_15691);
xor U17744 (N_17744,N_15733,N_15386);
or U17745 (N_17745,N_15867,N_16178);
xor U17746 (N_17746,N_15047,N_16396);
nand U17747 (N_17747,N_15326,N_16312);
and U17748 (N_17748,N_15603,N_15320);
and U17749 (N_17749,N_16064,N_15796);
and U17750 (N_17750,N_16239,N_15575);
nand U17751 (N_17751,N_15468,N_16078);
nor U17752 (N_17752,N_16341,N_16328);
nor U17753 (N_17753,N_15233,N_15036);
or U17754 (N_17754,N_15640,N_15029);
or U17755 (N_17755,N_16091,N_15497);
xor U17756 (N_17756,N_15339,N_16099);
nor U17757 (N_17757,N_16312,N_15548);
xor U17758 (N_17758,N_15749,N_15361);
or U17759 (N_17759,N_15801,N_15504);
and U17760 (N_17760,N_15696,N_15139);
or U17761 (N_17761,N_15344,N_15815);
or U17762 (N_17762,N_15205,N_15728);
nand U17763 (N_17763,N_15907,N_15947);
nand U17764 (N_17764,N_16336,N_16356);
and U17765 (N_17765,N_15700,N_15330);
or U17766 (N_17766,N_15532,N_15855);
xor U17767 (N_17767,N_15563,N_16064);
nor U17768 (N_17768,N_16221,N_15114);
nor U17769 (N_17769,N_16354,N_15738);
xor U17770 (N_17770,N_16341,N_16238);
nand U17771 (N_17771,N_15994,N_16360);
and U17772 (N_17772,N_16328,N_15534);
nand U17773 (N_17773,N_15085,N_15867);
xnor U17774 (N_17774,N_15969,N_15241);
and U17775 (N_17775,N_16370,N_15737);
and U17776 (N_17776,N_15001,N_15162);
nand U17777 (N_17777,N_15407,N_16186);
and U17778 (N_17778,N_15903,N_15135);
nor U17779 (N_17779,N_15175,N_15957);
nor U17780 (N_17780,N_15476,N_15301);
or U17781 (N_17781,N_16486,N_15850);
or U17782 (N_17782,N_16405,N_15047);
nand U17783 (N_17783,N_16392,N_15320);
and U17784 (N_17784,N_15266,N_16208);
nor U17785 (N_17785,N_15764,N_15663);
and U17786 (N_17786,N_15250,N_15247);
and U17787 (N_17787,N_16283,N_15673);
nor U17788 (N_17788,N_15910,N_15972);
and U17789 (N_17789,N_15475,N_15711);
nor U17790 (N_17790,N_15154,N_16043);
and U17791 (N_17791,N_15486,N_15862);
nand U17792 (N_17792,N_16312,N_16324);
or U17793 (N_17793,N_15268,N_15505);
nand U17794 (N_17794,N_15272,N_16243);
nand U17795 (N_17795,N_15979,N_15738);
or U17796 (N_17796,N_15541,N_15582);
nand U17797 (N_17797,N_15737,N_15514);
nor U17798 (N_17798,N_16240,N_16421);
nand U17799 (N_17799,N_15944,N_16305);
xor U17800 (N_17800,N_15907,N_15630);
nor U17801 (N_17801,N_15271,N_16419);
xnor U17802 (N_17802,N_16238,N_16053);
and U17803 (N_17803,N_16188,N_15396);
xnor U17804 (N_17804,N_16387,N_16073);
xor U17805 (N_17805,N_16026,N_15285);
nor U17806 (N_17806,N_15359,N_15365);
xnor U17807 (N_17807,N_16120,N_15554);
or U17808 (N_17808,N_15238,N_15032);
and U17809 (N_17809,N_15312,N_15268);
nand U17810 (N_17810,N_15921,N_15516);
and U17811 (N_17811,N_16422,N_15296);
nor U17812 (N_17812,N_15191,N_15693);
nor U17813 (N_17813,N_15206,N_15734);
nand U17814 (N_17814,N_16175,N_15170);
or U17815 (N_17815,N_16072,N_15377);
xnor U17816 (N_17816,N_16288,N_15487);
and U17817 (N_17817,N_16265,N_16037);
and U17818 (N_17818,N_15055,N_16447);
nor U17819 (N_17819,N_15554,N_16495);
or U17820 (N_17820,N_15906,N_15306);
or U17821 (N_17821,N_16278,N_16169);
or U17822 (N_17822,N_15396,N_15839);
and U17823 (N_17823,N_16484,N_15744);
and U17824 (N_17824,N_15866,N_15374);
xor U17825 (N_17825,N_15699,N_15151);
and U17826 (N_17826,N_16479,N_15877);
nand U17827 (N_17827,N_15442,N_16347);
xnor U17828 (N_17828,N_15192,N_16230);
nor U17829 (N_17829,N_16231,N_16068);
nor U17830 (N_17830,N_15165,N_15198);
xnor U17831 (N_17831,N_16256,N_15052);
and U17832 (N_17832,N_15721,N_15024);
and U17833 (N_17833,N_15812,N_15554);
and U17834 (N_17834,N_15729,N_15405);
nor U17835 (N_17835,N_15200,N_15409);
nor U17836 (N_17836,N_16175,N_15218);
xnor U17837 (N_17837,N_15570,N_15823);
nand U17838 (N_17838,N_15573,N_15991);
or U17839 (N_17839,N_15980,N_15001);
xnor U17840 (N_17840,N_15283,N_15884);
nand U17841 (N_17841,N_16164,N_15553);
nor U17842 (N_17842,N_15865,N_16268);
nor U17843 (N_17843,N_15503,N_16311);
nor U17844 (N_17844,N_15792,N_15407);
nor U17845 (N_17845,N_15969,N_15423);
and U17846 (N_17846,N_16244,N_15103);
or U17847 (N_17847,N_15900,N_16155);
nand U17848 (N_17848,N_16008,N_15160);
nand U17849 (N_17849,N_15902,N_15805);
nor U17850 (N_17850,N_15042,N_15531);
nand U17851 (N_17851,N_15983,N_15458);
and U17852 (N_17852,N_15523,N_16202);
or U17853 (N_17853,N_15923,N_16028);
or U17854 (N_17854,N_15323,N_15601);
xnor U17855 (N_17855,N_15183,N_16089);
and U17856 (N_17856,N_15239,N_16136);
or U17857 (N_17857,N_16302,N_15048);
nand U17858 (N_17858,N_16176,N_15731);
or U17859 (N_17859,N_16455,N_16412);
or U17860 (N_17860,N_15604,N_16460);
nand U17861 (N_17861,N_16052,N_16211);
nor U17862 (N_17862,N_15045,N_16246);
or U17863 (N_17863,N_15947,N_15394);
and U17864 (N_17864,N_16079,N_15899);
nand U17865 (N_17865,N_16452,N_15595);
xnor U17866 (N_17866,N_15179,N_15971);
nand U17867 (N_17867,N_16142,N_16114);
or U17868 (N_17868,N_15734,N_15574);
nand U17869 (N_17869,N_15298,N_16080);
and U17870 (N_17870,N_16451,N_15174);
nor U17871 (N_17871,N_15363,N_15814);
xor U17872 (N_17872,N_15140,N_15699);
nor U17873 (N_17873,N_15704,N_15639);
nor U17874 (N_17874,N_15344,N_15094);
and U17875 (N_17875,N_15681,N_15426);
nand U17876 (N_17876,N_16365,N_15110);
and U17877 (N_17877,N_15660,N_16108);
nand U17878 (N_17878,N_15276,N_16344);
xnor U17879 (N_17879,N_15433,N_15324);
nor U17880 (N_17880,N_16469,N_15029);
xor U17881 (N_17881,N_15502,N_15804);
nand U17882 (N_17882,N_16079,N_15847);
and U17883 (N_17883,N_15014,N_15285);
and U17884 (N_17884,N_16208,N_15840);
xnor U17885 (N_17885,N_15780,N_15511);
and U17886 (N_17886,N_15200,N_15213);
nand U17887 (N_17887,N_15287,N_15465);
xor U17888 (N_17888,N_15738,N_15613);
nand U17889 (N_17889,N_15304,N_16486);
and U17890 (N_17890,N_15327,N_15188);
nand U17891 (N_17891,N_16131,N_16080);
xor U17892 (N_17892,N_16387,N_16247);
xor U17893 (N_17893,N_16030,N_15404);
nand U17894 (N_17894,N_15782,N_16076);
xor U17895 (N_17895,N_15251,N_16477);
nor U17896 (N_17896,N_16036,N_15766);
xor U17897 (N_17897,N_16408,N_16422);
or U17898 (N_17898,N_15650,N_15061);
nor U17899 (N_17899,N_15144,N_16237);
nor U17900 (N_17900,N_15840,N_15034);
and U17901 (N_17901,N_15756,N_15750);
and U17902 (N_17902,N_15132,N_16334);
or U17903 (N_17903,N_16236,N_15755);
and U17904 (N_17904,N_15393,N_15255);
and U17905 (N_17905,N_15846,N_15443);
nand U17906 (N_17906,N_15390,N_16274);
nand U17907 (N_17907,N_16197,N_15742);
nor U17908 (N_17908,N_16465,N_16142);
xor U17909 (N_17909,N_16362,N_15377);
nor U17910 (N_17910,N_16124,N_16312);
nor U17911 (N_17911,N_15280,N_15437);
nor U17912 (N_17912,N_15197,N_16097);
nand U17913 (N_17913,N_15558,N_16003);
or U17914 (N_17914,N_15799,N_15068);
or U17915 (N_17915,N_15501,N_16323);
and U17916 (N_17916,N_16456,N_15797);
and U17917 (N_17917,N_15947,N_16306);
nand U17918 (N_17918,N_15378,N_15461);
nand U17919 (N_17919,N_15827,N_16243);
nor U17920 (N_17920,N_15841,N_15873);
nand U17921 (N_17921,N_15655,N_15358);
nand U17922 (N_17922,N_15682,N_15263);
or U17923 (N_17923,N_16434,N_15406);
xnor U17924 (N_17924,N_16476,N_15700);
xnor U17925 (N_17925,N_16434,N_15044);
nor U17926 (N_17926,N_15315,N_15034);
or U17927 (N_17927,N_15096,N_15671);
nand U17928 (N_17928,N_16323,N_15605);
or U17929 (N_17929,N_15595,N_15938);
nor U17930 (N_17930,N_16295,N_15928);
nor U17931 (N_17931,N_16207,N_16165);
nor U17932 (N_17932,N_15389,N_15096);
and U17933 (N_17933,N_16446,N_15225);
xnor U17934 (N_17934,N_16485,N_16166);
nor U17935 (N_17935,N_16463,N_15185);
and U17936 (N_17936,N_15460,N_15781);
nor U17937 (N_17937,N_15710,N_15232);
or U17938 (N_17938,N_15413,N_15824);
nor U17939 (N_17939,N_16240,N_16030);
and U17940 (N_17940,N_15257,N_16291);
nand U17941 (N_17941,N_15285,N_16293);
xnor U17942 (N_17942,N_16164,N_15390);
or U17943 (N_17943,N_16270,N_15732);
xor U17944 (N_17944,N_16067,N_16244);
xor U17945 (N_17945,N_16064,N_16304);
and U17946 (N_17946,N_16459,N_16082);
nor U17947 (N_17947,N_16414,N_16389);
nand U17948 (N_17948,N_15049,N_15125);
and U17949 (N_17949,N_15822,N_15767);
and U17950 (N_17950,N_15989,N_15383);
nor U17951 (N_17951,N_15112,N_15838);
and U17952 (N_17952,N_15610,N_16060);
or U17953 (N_17953,N_15241,N_15302);
nor U17954 (N_17954,N_16454,N_15697);
nand U17955 (N_17955,N_15293,N_15306);
nor U17956 (N_17956,N_15754,N_15933);
or U17957 (N_17957,N_16049,N_16017);
and U17958 (N_17958,N_15064,N_15229);
and U17959 (N_17959,N_16178,N_16241);
xor U17960 (N_17960,N_15050,N_16242);
nor U17961 (N_17961,N_15737,N_15245);
nand U17962 (N_17962,N_15608,N_16398);
and U17963 (N_17963,N_15487,N_16068);
and U17964 (N_17964,N_15187,N_15026);
or U17965 (N_17965,N_15288,N_16100);
or U17966 (N_17966,N_15310,N_15024);
xnor U17967 (N_17967,N_15056,N_16493);
and U17968 (N_17968,N_15133,N_15076);
xnor U17969 (N_17969,N_16172,N_15277);
nor U17970 (N_17970,N_16320,N_15027);
nor U17971 (N_17971,N_16313,N_16323);
xor U17972 (N_17972,N_15998,N_15888);
xnor U17973 (N_17973,N_15504,N_16294);
nor U17974 (N_17974,N_15109,N_15784);
or U17975 (N_17975,N_15108,N_16335);
nor U17976 (N_17976,N_15614,N_15886);
or U17977 (N_17977,N_15991,N_15711);
and U17978 (N_17978,N_15682,N_16459);
or U17979 (N_17979,N_15336,N_16313);
nor U17980 (N_17980,N_16397,N_15203);
nor U17981 (N_17981,N_15262,N_16299);
and U17982 (N_17982,N_15678,N_16309);
and U17983 (N_17983,N_16289,N_15497);
or U17984 (N_17984,N_16120,N_15443);
nand U17985 (N_17985,N_15229,N_15681);
nand U17986 (N_17986,N_16241,N_15716);
and U17987 (N_17987,N_15332,N_15194);
nor U17988 (N_17988,N_15018,N_16039);
xor U17989 (N_17989,N_16384,N_15455);
xnor U17990 (N_17990,N_16172,N_16044);
nand U17991 (N_17991,N_16443,N_15897);
nand U17992 (N_17992,N_15281,N_15024);
nand U17993 (N_17993,N_15124,N_16319);
and U17994 (N_17994,N_15299,N_15721);
nand U17995 (N_17995,N_16044,N_15128);
nand U17996 (N_17996,N_15790,N_16384);
nand U17997 (N_17997,N_15397,N_16460);
and U17998 (N_17998,N_15117,N_16110);
nor U17999 (N_17999,N_16318,N_16475);
nand U18000 (N_18000,N_17920,N_17673);
or U18001 (N_18001,N_17741,N_16503);
or U18002 (N_18002,N_17164,N_17902);
nor U18003 (N_18003,N_16945,N_17692);
or U18004 (N_18004,N_17691,N_16588);
or U18005 (N_18005,N_17680,N_16891);
and U18006 (N_18006,N_17955,N_17355);
nor U18007 (N_18007,N_17874,N_17236);
nor U18008 (N_18008,N_17634,N_16923);
and U18009 (N_18009,N_17951,N_16708);
xor U18010 (N_18010,N_16640,N_16686);
or U18011 (N_18011,N_16541,N_16632);
and U18012 (N_18012,N_17319,N_17036);
or U18013 (N_18013,N_16739,N_16723);
xnor U18014 (N_18014,N_17128,N_17986);
nor U18015 (N_18015,N_16918,N_17081);
or U18016 (N_18016,N_17817,N_17767);
nand U18017 (N_18017,N_17743,N_17681);
xor U18018 (N_18018,N_17672,N_16556);
and U18019 (N_18019,N_17287,N_16715);
and U18020 (N_18020,N_16719,N_17478);
xor U18021 (N_18021,N_17099,N_17985);
xnor U18022 (N_18022,N_17602,N_16969);
or U18023 (N_18023,N_17948,N_16873);
nor U18024 (N_18024,N_17199,N_17538);
xor U18025 (N_18025,N_17086,N_17001);
or U18026 (N_18026,N_17092,N_16879);
nand U18027 (N_18027,N_16865,N_17658);
and U18028 (N_18028,N_16591,N_17548);
and U18029 (N_18029,N_16652,N_17089);
or U18030 (N_18030,N_16593,N_16724);
and U18031 (N_18031,N_16621,N_17305);
nor U18032 (N_18032,N_17712,N_17555);
or U18033 (N_18033,N_16960,N_17542);
nor U18034 (N_18034,N_16695,N_17540);
xnor U18035 (N_18035,N_16603,N_17091);
or U18036 (N_18036,N_17158,N_17491);
xnor U18037 (N_18037,N_17911,N_17374);
or U18038 (N_18038,N_17077,N_16505);
nor U18039 (N_18039,N_17150,N_17040);
or U18040 (N_18040,N_17313,N_17282);
xor U18041 (N_18041,N_16731,N_16849);
xor U18042 (N_18042,N_17061,N_17957);
nand U18043 (N_18043,N_16911,N_16792);
nor U18044 (N_18044,N_17775,N_16757);
and U18045 (N_18045,N_16906,N_17293);
and U18046 (N_18046,N_17172,N_17290);
nor U18047 (N_18047,N_17119,N_17849);
xor U18048 (N_18048,N_17567,N_16617);
and U18049 (N_18049,N_17472,N_16942);
or U18050 (N_18050,N_16905,N_16678);
or U18051 (N_18051,N_16675,N_17873);
and U18052 (N_18052,N_17746,N_17505);
nand U18053 (N_18053,N_17580,N_17812);
or U18054 (N_18054,N_16705,N_16784);
and U18055 (N_18055,N_17689,N_17460);
nand U18056 (N_18056,N_17552,N_16627);
xor U18057 (N_18057,N_17255,N_16579);
nand U18058 (N_18058,N_17262,N_17071);
or U18059 (N_18059,N_17582,N_16530);
nor U18060 (N_18060,N_17605,N_17063);
or U18061 (N_18061,N_16882,N_16733);
nand U18062 (N_18062,N_17385,N_16573);
nor U18063 (N_18063,N_17932,N_17659);
and U18064 (N_18064,N_17346,N_17393);
nor U18065 (N_18065,N_17517,N_17095);
and U18066 (N_18066,N_17576,N_17894);
xnor U18067 (N_18067,N_17926,N_17131);
and U18068 (N_18068,N_17760,N_17772);
nand U18069 (N_18069,N_16963,N_17843);
or U18070 (N_18070,N_17992,N_16880);
or U18071 (N_18071,N_17660,N_16629);
xnor U18072 (N_18072,N_17151,N_17525);
and U18073 (N_18073,N_16990,N_16657);
and U18074 (N_18074,N_17954,N_17773);
xnor U18075 (N_18075,N_17541,N_17882);
xnor U18076 (N_18076,N_17578,N_17014);
xor U18077 (N_18077,N_16894,N_16779);
or U18078 (N_18078,N_17802,N_17280);
nor U18079 (N_18079,N_16718,N_17807);
nand U18080 (N_18080,N_17982,N_17237);
and U18081 (N_18081,N_17766,N_17581);
xor U18082 (N_18082,N_17011,N_16997);
nand U18083 (N_18083,N_17279,N_17976);
nor U18084 (N_18084,N_17936,N_17345);
nand U18085 (N_18085,N_17209,N_16871);
xor U18086 (N_18086,N_17832,N_17546);
and U18087 (N_18087,N_17154,N_16562);
and U18088 (N_18088,N_16806,N_17571);
xnor U18089 (N_18089,N_16798,N_16580);
and U18090 (N_18090,N_17075,N_17575);
nor U18091 (N_18091,N_16890,N_16743);
xnor U18092 (N_18092,N_17499,N_16720);
nand U18093 (N_18093,N_17443,N_17211);
and U18094 (N_18094,N_16722,N_17550);
nand U18095 (N_18095,N_17267,N_16977);
and U18096 (N_18096,N_17904,N_16878);
nor U18097 (N_18097,N_17340,N_17858);
nand U18098 (N_18098,N_16655,N_17713);
nand U18099 (N_18099,N_17875,N_17501);
nor U18100 (N_18100,N_17852,N_17429);
nand U18101 (N_18101,N_17514,N_16677);
and U18102 (N_18102,N_16927,N_17600);
nand U18103 (N_18103,N_17927,N_17591);
nor U18104 (N_18104,N_16851,N_17225);
and U18105 (N_18105,N_16932,N_17263);
or U18106 (N_18106,N_17844,N_17379);
xor U18107 (N_18107,N_17959,N_17776);
or U18108 (N_18108,N_17376,N_17108);
xnor U18109 (N_18109,N_16807,N_16740);
or U18110 (N_18110,N_17815,N_16800);
nand U18111 (N_18111,N_16864,N_16998);
or U18112 (N_18112,N_17958,N_17984);
nor U18113 (N_18113,N_17603,N_17761);
or U18114 (N_18114,N_17436,N_16525);
or U18115 (N_18115,N_16786,N_17899);
nand U18116 (N_18116,N_17019,N_16809);
and U18117 (N_18117,N_16701,N_17922);
xor U18118 (N_18118,N_16512,N_16707);
nand U18119 (N_18119,N_16665,N_17228);
xor U18120 (N_18120,N_16544,N_17022);
nor U18121 (N_18121,N_16673,N_16915);
and U18122 (N_18122,N_17448,N_17521);
xnor U18123 (N_18123,N_17928,N_17269);
nor U18124 (N_18124,N_16860,N_17881);
and U18125 (N_18125,N_17284,N_17895);
nand U18126 (N_18126,N_17921,N_17117);
or U18127 (N_18127,N_16558,N_16528);
and U18128 (N_18128,N_16616,N_16821);
or U18129 (N_18129,N_17333,N_17683);
xnor U18130 (N_18130,N_16978,N_17424);
nand U18131 (N_18131,N_16926,N_17097);
nand U18132 (N_18132,N_17068,N_16670);
nand U18133 (N_18133,N_17141,N_17388);
nor U18134 (N_18134,N_17822,N_16728);
and U18135 (N_18135,N_17532,N_17855);
nand U18136 (N_18136,N_17406,N_17711);
or U18137 (N_18137,N_16703,N_17260);
nand U18138 (N_18138,N_17656,N_16826);
nor U18139 (N_18139,N_17023,N_17777);
nor U18140 (N_18140,N_17993,N_17868);
or U18141 (N_18141,N_17122,N_16683);
nand U18142 (N_18142,N_17836,N_17477);
xor U18143 (N_18143,N_17695,N_17737);
or U18144 (N_18144,N_16529,N_17239);
nor U18145 (N_18145,N_17918,N_16518);
nand U18146 (N_18146,N_16856,N_16599);
and U18147 (N_18147,N_17130,N_16790);
xnor U18148 (N_18148,N_16537,N_17915);
nand U18149 (N_18149,N_17980,N_16622);
and U18150 (N_18150,N_17411,N_16714);
nor U18151 (N_18151,N_16958,N_17662);
and U18152 (N_18152,N_17139,N_16630);
nand U18153 (N_18153,N_17268,N_17784);
and U18154 (N_18154,N_17961,N_16870);
nor U18155 (N_18155,N_16964,N_17048);
xnor U18156 (N_18156,N_17184,N_17021);
nand U18157 (N_18157,N_16660,N_17870);
or U18158 (N_18158,N_17314,N_17988);
nor U18159 (N_18159,N_17467,N_17618);
nor U18160 (N_18160,N_16506,N_16702);
nand U18161 (N_18161,N_16534,N_16750);
and U18162 (N_18162,N_17781,N_16837);
and U18163 (N_18163,N_17872,N_17206);
nor U18164 (N_18164,N_17352,N_17408);
nand U18165 (N_18165,N_16572,N_17087);
xnor U18166 (N_18166,N_17892,N_17685);
nand U18167 (N_18167,N_17360,N_17939);
and U18168 (N_18168,N_17487,N_16565);
or U18169 (N_18169,N_17450,N_17572);
nor U18170 (N_18170,N_17426,N_17213);
xnor U18171 (N_18171,N_17805,N_16748);
nor U18172 (N_18172,N_17967,N_17465);
or U18173 (N_18173,N_17190,N_17794);
and U18174 (N_18174,N_17811,N_17965);
or U18175 (N_18175,N_17787,N_17964);
nand U18176 (N_18176,N_17337,N_17729);
nand U18177 (N_18177,N_17447,N_17297);
nand U18178 (N_18178,N_17029,N_17381);
and U18179 (N_18179,N_16568,N_16966);
and U18180 (N_18180,N_16754,N_17718);
and U18181 (N_18181,N_17226,N_17528);
xor U18182 (N_18182,N_17930,N_17179);
and U18183 (N_18183,N_17455,N_17281);
xnor U18184 (N_18184,N_17938,N_17088);
nand U18185 (N_18185,N_17235,N_16884);
or U18186 (N_18186,N_17728,N_17057);
and U18187 (N_18187,N_16609,N_16853);
or U18188 (N_18188,N_17181,N_17842);
or U18189 (N_18189,N_16547,N_16758);
or U18190 (N_18190,N_17367,N_17702);
nor U18191 (N_18191,N_16698,N_17944);
nor U18192 (N_18192,N_17007,N_17624);
and U18193 (N_18193,N_16578,N_17800);
or U18194 (N_18194,N_17744,N_17474);
or U18195 (N_18195,N_17302,N_17891);
nand U18196 (N_18196,N_17142,N_17304);
nand U18197 (N_18197,N_17511,N_17035);
and U18198 (N_18198,N_16581,N_17249);
nor U18199 (N_18199,N_17299,N_16532);
nor U18200 (N_18200,N_17963,N_17459);
nand U18201 (N_18201,N_16667,N_16862);
or U18202 (N_18202,N_17339,N_16727);
and U18203 (N_18203,N_16676,N_17537);
and U18204 (N_18204,N_17522,N_17292);
nor U18205 (N_18205,N_17286,N_17682);
xnor U18206 (N_18206,N_17661,N_17869);
nor U18207 (N_18207,N_17277,N_16624);
and U18208 (N_18208,N_17318,N_17900);
nor U18209 (N_18209,N_17167,N_17278);
xor U18210 (N_18210,N_16858,N_17405);
nand U18211 (N_18211,N_17101,N_17136);
and U18212 (N_18212,N_17203,N_17752);
xnor U18213 (N_18213,N_17303,N_17608);
xor U18214 (N_18214,N_16938,N_17826);
xnor U18215 (N_18215,N_17419,N_17733);
nand U18216 (N_18216,N_17977,N_16623);
nor U18217 (N_18217,N_17909,N_17774);
and U18218 (N_18218,N_16540,N_16876);
or U18219 (N_18219,N_16931,N_17952);
xor U18220 (N_18220,N_17722,N_17905);
nor U18221 (N_18221,N_17753,N_17422);
nand U18222 (N_18222,N_16820,N_17845);
and U18223 (N_18223,N_17912,N_16612);
nand U18224 (N_18224,N_17748,N_17613);
and U18225 (N_18225,N_17543,N_16764);
xor U18226 (N_18226,N_17193,N_17125);
nor U18227 (N_18227,N_17182,N_17594);
nor U18228 (N_18228,N_16606,N_17867);
or U18229 (N_18229,N_16638,N_17013);
xor U18230 (N_18230,N_17536,N_16551);
nor U18231 (N_18231,N_16545,N_16682);
and U18232 (N_18232,N_16561,N_17641);
nand U18233 (N_18233,N_17326,N_16608);
nand U18234 (N_18234,N_17960,N_17378);
and U18235 (N_18235,N_17336,N_16649);
nor U18236 (N_18236,N_16937,N_17883);
nand U18237 (N_18237,N_16797,N_17224);
and U18238 (N_18238,N_16704,N_17910);
nand U18239 (N_18239,N_17082,N_17783);
nand U18240 (N_18240,N_16611,N_16751);
or U18241 (N_18241,N_17464,N_17549);
nand U18242 (N_18242,N_17551,N_17454);
and U18243 (N_18243,N_17338,N_17923);
or U18244 (N_18244,N_17327,N_17598);
and U18245 (N_18245,N_16514,N_17207);
xor U18246 (N_18246,N_17569,N_17573);
nor U18247 (N_18247,N_17169,N_17710);
nor U18248 (N_18248,N_17100,N_17435);
or U18249 (N_18249,N_17851,N_16737);
nor U18250 (N_18250,N_16916,N_17390);
and U18251 (N_18251,N_16895,N_17165);
nand U18252 (N_18252,N_16671,N_17451);
xor U18253 (N_18253,N_17749,N_17740);
nand U18254 (N_18254,N_17504,N_17968);
and U18255 (N_18255,N_16597,N_17577);
xor U18256 (N_18256,N_17901,N_17362);
and U18257 (N_18257,N_16590,N_17386);
xnor U18258 (N_18258,N_17322,N_17045);
and U18259 (N_18259,N_17606,N_17137);
nand U18260 (N_18260,N_17757,N_17078);
nand U18261 (N_18261,N_17859,N_17524);
and U18262 (N_18262,N_17469,N_16953);
nand U18263 (N_18263,N_16818,N_17820);
and U18264 (N_18264,N_16986,N_17545);
nor U18265 (N_18265,N_16583,N_16600);
and U18266 (N_18266,N_17442,N_17865);
and U18267 (N_18267,N_17486,N_17159);
or U18268 (N_18268,N_17186,N_17444);
nand U18269 (N_18269,N_16634,N_17298);
and U18270 (N_18270,N_17679,N_16713);
nor U18271 (N_18271,N_17717,N_17970);
and U18272 (N_18272,N_16582,N_16929);
nand U18273 (N_18273,N_16808,N_17413);
and U18274 (N_18274,N_17925,N_17067);
or U18275 (N_18275,N_16653,N_17990);
nand U18276 (N_18276,N_17003,N_17046);
xor U18277 (N_18277,N_17132,N_17372);
and U18278 (N_18278,N_17462,N_17719);
nor U18279 (N_18279,N_17017,N_17126);
and U18280 (N_18280,N_17898,N_17566);
and U18281 (N_18281,N_16507,N_17694);
nand U18282 (N_18282,N_16753,N_17838);
and U18283 (N_18283,N_16699,N_16888);
and U18284 (N_18284,N_16557,N_16825);
nor U18285 (N_18285,N_16542,N_17354);
nor U18286 (N_18286,N_17171,N_17621);
nand U18287 (N_18287,N_17888,N_16531);
xnor U18288 (N_18288,N_17198,N_16955);
or U18289 (N_18289,N_17368,N_17956);
nor U18290 (N_18290,N_17770,N_17789);
and U18291 (N_18291,N_17759,N_17107);
xnor U18292 (N_18292,N_17589,N_17509);
nand U18293 (N_18293,N_17166,N_16946);
nand U18294 (N_18294,N_17696,N_16552);
or U18295 (N_18295,N_16840,N_16988);
xnor U18296 (N_18296,N_16789,N_16635);
or U18297 (N_18297,N_17227,N_17220);
and U18298 (N_18298,N_17009,N_17330);
or U18299 (N_18299,N_17649,N_17173);
nand U18300 (N_18300,N_17792,N_17051);
and U18301 (N_18301,N_16883,N_16996);
xor U18302 (N_18302,N_17428,N_17991);
or U18303 (N_18303,N_16976,N_17008);
or U18304 (N_18304,N_16885,N_16995);
nand U18305 (N_18305,N_17535,N_17627);
nor U18306 (N_18306,N_16548,N_16538);
or U18307 (N_18307,N_17294,N_17863);
or U18308 (N_18308,N_17275,N_16761);
or U18309 (N_18309,N_16510,N_17331);
xnor U18310 (N_18310,N_16515,N_17312);
nand U18311 (N_18311,N_16625,N_16989);
or U18312 (N_18312,N_16838,N_16661);
nand U18313 (N_18313,N_17989,N_17244);
and U18314 (N_18314,N_16913,N_16650);
nand U18315 (N_18315,N_17060,N_17473);
nor U18316 (N_18316,N_17079,N_17796);
or U18317 (N_18317,N_17389,N_17430);
nand U18318 (N_18318,N_16824,N_17183);
xnor U18319 (N_18319,N_16971,N_17636);
and U18320 (N_18320,N_16717,N_17468);
or U18321 (N_18321,N_17324,N_17369);
nor U18322 (N_18322,N_16907,N_17265);
xor U18323 (N_18323,N_16567,N_17885);
nor U18324 (N_18324,N_17519,N_17457);
or U18325 (N_18325,N_17026,N_17560);
xnor U18326 (N_18326,N_17846,N_16794);
or U18327 (N_18327,N_17847,N_17876);
xnor U18328 (N_18328,N_17392,N_16857);
xor U18329 (N_18329,N_17848,N_17808);
nand U18330 (N_18330,N_16633,N_16815);
or U18331 (N_18331,N_17098,N_16684);
nor U18332 (N_18332,N_17937,N_16975);
nand U18333 (N_18333,N_17052,N_17234);
and U18334 (N_18334,N_17671,N_17147);
nand U18335 (N_18335,N_17357,N_16787);
nor U18336 (N_18336,N_16520,N_16968);
nand U18337 (N_18337,N_17670,N_17053);
nand U18338 (N_18338,N_17096,N_17231);
xnor U18339 (N_18339,N_17622,N_16680);
nor U18340 (N_18340,N_16762,N_16850);
nor U18341 (N_18341,N_17720,N_17270);
xnor U18342 (N_18342,N_17177,N_17252);
and U18343 (N_18343,N_17332,N_16993);
nor U18344 (N_18344,N_16877,N_16767);
and U18345 (N_18345,N_17410,N_17837);
xnor U18346 (N_18346,N_16760,N_17738);
nor U18347 (N_18347,N_17084,N_17497);
or U18348 (N_18348,N_17697,N_17754);
nand U18349 (N_18349,N_17187,N_17397);
nor U18350 (N_18350,N_17348,N_17431);
nor U18351 (N_18351,N_17438,N_16994);
xnor U18352 (N_18352,N_16829,N_17246);
or U18353 (N_18353,N_17440,N_17109);
or U18354 (N_18354,N_17050,N_17635);
xnor U18355 (N_18355,N_17655,N_17599);
and U18356 (N_18356,N_16711,N_17375);
or U18357 (N_18357,N_17706,N_17160);
and U18358 (N_18358,N_17854,N_17197);
nor U18359 (N_18359,N_17601,N_16559);
and U18360 (N_18360,N_16636,N_17768);
xnor U18361 (N_18361,N_17156,N_17884);
nand U18362 (N_18362,N_17590,N_17423);
or U18363 (N_18363,N_17420,N_17809);
nand U18364 (N_18364,N_17643,N_17000);
or U18365 (N_18365,N_17795,N_17913);
nor U18366 (N_18366,N_16774,N_16536);
and U18367 (N_18367,N_16553,N_16972);
and U18368 (N_18368,N_17349,N_16859);
xnor U18369 (N_18369,N_17018,N_16613);
or U18370 (N_18370,N_16984,N_17983);
nor U18371 (N_18371,N_16811,N_17507);
or U18372 (N_18372,N_17476,N_17359);
or U18373 (N_18373,N_17105,N_16844);
nor U18374 (N_18374,N_16898,N_16941);
nand U18375 (N_18375,N_17996,N_17684);
or U18376 (N_18376,N_16663,N_17445);
or U18377 (N_18377,N_17121,N_16940);
xnor U18378 (N_18378,N_17306,N_17291);
nand U18379 (N_18379,N_17083,N_17138);
nand U18380 (N_18380,N_17929,N_17202);
or U18381 (N_18381,N_16706,N_16517);
or U18382 (N_18382,N_17219,N_17033);
xor U18383 (N_18383,N_17174,N_16745);
nor U18384 (N_18384,N_16812,N_17508);
nand U18385 (N_18385,N_16516,N_17637);
nand U18386 (N_18386,N_17371,N_16901);
or U18387 (N_18387,N_17821,N_17633);
or U18388 (N_18388,N_17607,N_17002);
nor U18389 (N_18389,N_17295,N_17343);
xor U18390 (N_18390,N_17334,N_16991);
and U18391 (N_18391,N_16816,N_16928);
xnor U18392 (N_18392,N_16763,N_17004);
xnor U18393 (N_18393,N_17810,N_16620);
xor U18394 (N_18394,N_16666,N_16967);
xor U18395 (N_18395,N_17678,N_16626);
xor U18396 (N_18396,N_16845,N_17437);
and U18397 (N_18397,N_17878,N_17488);
and U18398 (N_18398,N_17129,N_17449);
xnor U18399 (N_18399,N_17638,N_17654);
nand U18400 (N_18400,N_16725,N_17625);
xnor U18401 (N_18401,N_17401,N_16791);
or U18402 (N_18402,N_16965,N_16933);
nor U18403 (N_18403,N_16999,N_16914);
or U18404 (N_18404,N_17663,N_16846);
nor U18405 (N_18405,N_17785,N_17341);
or U18406 (N_18406,N_17316,N_16726);
and U18407 (N_18407,N_17818,N_17479);
or U18408 (N_18408,N_16773,N_16560);
nor U18409 (N_18409,N_17495,N_16687);
or U18410 (N_18410,N_17947,N_17258);
xnor U18411 (N_18411,N_17049,N_17750);
nand U18412 (N_18412,N_16604,N_17645);
nor U18413 (N_18413,N_17726,N_17490);
or U18414 (N_18414,N_17118,N_17971);
and U18415 (N_18415,N_17919,N_17840);
xnor U18416 (N_18416,N_17688,N_17946);
and U18417 (N_18417,N_16951,N_17651);
nor U18418 (N_18418,N_17588,N_17853);
nor U18419 (N_18419,N_16902,N_16742);
and U18420 (N_18420,N_17834,N_17315);
or U18421 (N_18421,N_17272,N_16654);
and U18422 (N_18422,N_17221,N_16904);
nand U18423 (N_18423,N_16692,N_17188);
and U18424 (N_18424,N_16519,N_17038);
nand U18425 (N_18425,N_16747,N_17148);
or U18426 (N_18426,N_17416,N_17631);
xnor U18427 (N_18427,N_17667,N_17877);
nor U18428 (N_18428,N_16527,N_17502);
nand U18429 (N_18429,N_17526,N_17778);
nor U18430 (N_18430,N_17288,N_17028);
or U18431 (N_18431,N_17042,N_16674);
nand U18432 (N_18432,N_17686,N_16892);
or U18433 (N_18433,N_17358,N_17257);
nor U18434 (N_18434,N_16508,N_17714);
and U18435 (N_18435,N_16917,N_17168);
and U18436 (N_18436,N_17391,N_17403);
nand U18437 (N_18437,N_16783,N_17253);
xor U18438 (N_18438,N_17987,N_17310);
and U18439 (N_18439,N_17398,N_17639);
and U18440 (N_18440,N_17751,N_17797);
nand U18441 (N_18441,N_17604,N_17162);
xor U18442 (N_18442,N_17112,N_16841);
nand U18443 (N_18443,N_16772,N_16852);
nand U18444 (N_18444,N_17276,N_16924);
nor U18445 (N_18445,N_17981,N_17969);
nor U18446 (N_18446,N_17407,N_17155);
or U18447 (N_18447,N_17835,N_17563);
nor U18448 (N_18448,N_17782,N_17062);
nor U18449 (N_18449,N_17243,N_16823);
or U18450 (N_18450,N_17144,N_17758);
nor U18451 (N_18451,N_17736,N_16690);
nand U18452 (N_18452,N_17300,N_17646);
or U18453 (N_18453,N_17103,N_16819);
or U18454 (N_18454,N_16668,N_17134);
and U18455 (N_18455,N_16781,N_17212);
xor U18456 (N_18456,N_17283,N_16575);
nand U18457 (N_18457,N_17123,N_17534);
nor U18458 (N_18458,N_17072,N_16983);
or U18459 (N_18459,N_16637,N_17700);
and U18460 (N_18460,N_17069,N_17344);
xor U18461 (N_18461,N_17841,N_17180);
nand U18462 (N_18462,N_16749,N_17579);
nor U18463 (N_18463,N_17034,N_17361);
nand U18464 (N_18464,N_17065,N_17801);
nor U18465 (N_18465,N_17323,N_16521);
or U18466 (N_18466,N_16589,N_17041);
nor U18467 (N_18467,N_17570,N_16974);
and U18468 (N_18468,N_16697,N_16755);
nor U18469 (N_18469,N_17115,N_16944);
nor U18470 (N_18470,N_17178,N_16832);
or U18471 (N_18471,N_17425,N_17565);
xnor U18472 (N_18472,N_17020,N_17248);
nand U18473 (N_18473,N_17196,N_16896);
nand U18474 (N_18474,N_17723,N_17616);
or U18475 (N_18475,N_16833,N_17494);
or U18476 (N_18476,N_16689,N_17666);
nand U18477 (N_18477,N_16778,N_17030);
nand U18478 (N_18478,N_16566,N_17975);
nand U18479 (N_18479,N_17953,N_16768);
nand U18480 (N_18480,N_16709,N_16881);
nor U18481 (N_18481,N_17597,N_17974);
or U18482 (N_18482,N_17074,N_17195);
xor U18483 (N_18483,N_16736,N_17309);
xnor U18484 (N_18484,N_17005,N_17626);
nand U18485 (N_18485,N_17145,N_17617);
nand U18486 (N_18486,N_16549,N_16685);
nor U18487 (N_18487,N_17215,N_17725);
nor U18488 (N_18488,N_17483,N_17311);
nor U18489 (N_18489,N_17995,N_16756);
and U18490 (N_18490,N_17871,N_17675);
and U18491 (N_18491,N_17113,N_16641);
or U18492 (N_18492,N_17328,N_17149);
and U18493 (N_18493,N_17819,N_16672);
xor U18494 (N_18494,N_16522,N_17619);
or U18495 (N_18495,N_16691,N_17764);
nand U18496 (N_18496,N_17755,N_17648);
nand U18497 (N_18497,N_17031,N_16651);
or U18498 (N_18498,N_16866,N_17427);
nand U18499 (N_18499,N_16586,N_17471);
xnor U18500 (N_18500,N_16771,N_17321);
nand U18501 (N_18501,N_17039,N_16992);
nor U18502 (N_18502,N_16730,N_17831);
and U18503 (N_18503,N_17903,N_16788);
nand U18504 (N_18504,N_17516,N_17308);
or U18505 (N_18505,N_16863,N_17140);
nand U18506 (N_18506,N_16546,N_17492);
nor U18507 (N_18507,N_16872,N_17241);
and U18508 (N_18508,N_17110,N_17073);
xnor U18509 (N_18509,N_17596,N_17734);
and U18510 (N_18510,N_17503,N_16839);
nand U18511 (N_18511,N_17701,N_17254);
or U18512 (N_18512,N_17146,N_17529);
or U18513 (N_18513,N_16602,N_17256);
nand U18514 (N_18514,N_16869,N_17015);
and U18515 (N_18515,N_17044,N_17730);
nor U18516 (N_18516,N_17245,N_17793);
nand U18517 (N_18517,N_16664,N_17273);
or U18518 (N_18518,N_17886,N_16775);
xor U18519 (N_18519,N_17676,N_17289);
and U18520 (N_18520,N_16569,N_17715);
nand U18521 (N_18521,N_17553,N_17642);
or U18522 (N_18522,N_17480,N_16732);
nor U18523 (N_18523,N_17907,N_17674);
nand U18524 (N_18524,N_17644,N_17630);
nor U18525 (N_18525,N_16954,N_17623);
nor U18526 (N_18526,N_16939,N_16574);
nor U18527 (N_18527,N_17556,N_16741);
and U18528 (N_18528,N_17771,N_17612);
or U18529 (N_18529,N_17043,N_16947);
nor U18530 (N_18530,N_17012,N_16601);
nand U18531 (N_18531,N_16899,N_17880);
or U18532 (N_18532,N_17271,N_17827);
or U18533 (N_18533,N_16959,N_16822);
or U18534 (N_18534,N_17064,N_17587);
and U18535 (N_18535,N_17238,N_16681);
and U18536 (N_18536,N_17924,N_16867);
or U18537 (N_18537,N_17561,N_17506);
nor U18538 (N_18538,N_17531,N_17716);
nor U18539 (N_18539,N_16961,N_17482);
and U18540 (N_18540,N_17942,N_17940);
or U18541 (N_18541,N_17916,N_16694);
nand U18542 (N_18542,N_17489,N_17978);
or U18543 (N_18543,N_16843,N_16770);
or U18544 (N_18544,N_17583,N_17214);
nand U18545 (N_18545,N_16943,N_16576);
nor U18546 (N_18546,N_16526,N_17152);
and U18547 (N_18547,N_16563,N_16813);
or U18548 (N_18548,N_16908,N_17432);
xor U18549 (N_18549,N_16628,N_17453);
and U18550 (N_18550,N_17027,N_16607);
and U18551 (N_18551,N_17054,N_17402);
nor U18552 (N_18552,N_17370,N_17461);
nand U18553 (N_18553,N_16639,N_17414);
nor U18554 (N_18554,N_16631,N_17935);
xnor U18555 (N_18555,N_16716,N_17979);
nand U18556 (N_18556,N_17512,N_16889);
and U18557 (N_18557,N_17363,N_17493);
and U18558 (N_18558,N_17135,N_17615);
xnor U18559 (N_18559,N_17966,N_17564);
xor U18560 (N_18560,N_17931,N_17409);
nor U18561 (N_18561,N_17780,N_16729);
xnor U18562 (N_18562,N_16903,N_17724);
xor U18563 (N_18563,N_17301,N_17047);
or U18564 (N_18564,N_16584,N_17415);
or U18565 (N_18565,N_16533,N_17839);
nor U18566 (N_18566,N_17317,N_17475);
or U18567 (N_18567,N_16746,N_17699);
and U18568 (N_18568,N_16847,N_16615);
nor U18569 (N_18569,N_17189,N_16827);
xnor U18570 (N_18570,N_17208,N_17024);
or U18571 (N_18571,N_16643,N_16535);
nand U18572 (N_18572,N_16776,N_16605);
xnor U18573 (N_18573,N_17163,N_17698);
nand U18574 (N_18574,N_17223,N_17058);
nor U18575 (N_18575,N_17703,N_17803);
and U18576 (N_18576,N_17210,N_16550);
nand U18577 (N_18577,N_17804,N_16614);
xnor U18578 (N_18578,N_17704,N_17747);
xor U18579 (N_18579,N_17914,N_16956);
nor U18580 (N_18580,N_16836,N_17412);
xor U18581 (N_18581,N_17335,N_16577);
nor U18582 (N_18582,N_17353,N_16886);
or U18583 (N_18583,N_17261,N_17693);
and U18584 (N_18584,N_17400,N_17554);
nor U18585 (N_18585,N_17104,N_17157);
or U18586 (N_18586,N_17647,N_17568);
or U18587 (N_18587,N_17366,N_17595);
or U18588 (N_18588,N_16752,N_16912);
or U18589 (N_18589,N_17161,N_17404);
nand U18590 (N_18590,N_17185,N_17285);
xnor U18591 (N_18591,N_17788,N_17204);
and U18592 (N_18592,N_16814,N_17394);
xnor U18593 (N_18593,N_17527,N_16817);
xor U18594 (N_18594,N_16828,N_17170);
xnor U18595 (N_18595,N_17094,N_17350);
nand U18596 (N_18596,N_17828,N_17347);
and U18597 (N_18597,N_17233,N_17708);
and U18598 (N_18598,N_17373,N_16922);
nor U18599 (N_18599,N_17857,N_17264);
and U18600 (N_18600,N_17574,N_16982);
xor U18601 (N_18601,N_17106,N_17325);
or U18602 (N_18602,N_17798,N_17342);
and U18603 (N_18603,N_17814,N_17176);
or U18604 (N_18604,N_16759,N_16909);
xor U18605 (N_18605,N_17879,N_17153);
or U18606 (N_18606,N_17949,N_17791);
nand U18607 (N_18607,N_17732,N_17102);
xor U18608 (N_18608,N_17653,N_17090);
and U18609 (N_18609,N_16782,N_17889);
and U18610 (N_18610,N_17830,N_16669);
and U18611 (N_18611,N_16744,N_16950);
nand U18612 (N_18612,N_17893,N_17470);
or U18613 (N_18613,N_16970,N_16648);
nor U18614 (N_18614,N_16555,N_17259);
or U18615 (N_18615,N_17890,N_17510);
nand U18616 (N_18616,N_17668,N_17456);
nand U18617 (N_18617,N_17786,N_17640);
nand U18618 (N_18618,N_17620,N_16921);
nor U18619 (N_18619,N_17066,N_17111);
xnor U18620 (N_18620,N_17191,N_17143);
nor U18621 (N_18621,N_17055,N_17523);
nor U18622 (N_18622,N_17650,N_17080);
nand U18623 (N_18623,N_17250,N_17395);
xor U18624 (N_18624,N_17611,N_16848);
or U18625 (N_18625,N_17377,N_16659);
xor U18626 (N_18626,N_16874,N_16793);
and U18627 (N_18627,N_17742,N_17823);
or U18628 (N_18628,N_16766,N_16930);
or U18629 (N_18629,N_16642,N_17593);
nand U18630 (N_18630,N_17518,N_17941);
and U18631 (N_18631,N_17120,N_17544);
nand U18632 (N_18632,N_17652,N_17559);
nand U18633 (N_18633,N_16598,N_16679);
xnor U18634 (N_18634,N_17421,N_17240);
or U18635 (N_18635,N_17887,N_17896);
xor U18636 (N_18636,N_17439,N_16662);
nand U18637 (N_18637,N_16868,N_16981);
nor U18638 (N_18638,N_16925,N_17833);
nand U18639 (N_18639,N_16897,N_17779);
xor U18640 (N_18640,N_17498,N_17687);
nor U18641 (N_18641,N_17387,N_16805);
nor U18642 (N_18642,N_16952,N_17945);
and U18643 (N_18643,N_17962,N_16920);
nand U18644 (N_18644,N_17307,N_16948);
xnor U18645 (N_18645,N_16543,N_16962);
and U18646 (N_18646,N_17533,N_17765);
xnor U18647 (N_18647,N_17707,N_17562);
and U18648 (N_18648,N_17709,N_17799);
nor U18649 (N_18649,N_17356,N_17365);
and U18650 (N_18650,N_16610,N_17632);
nor U18651 (N_18651,N_16587,N_17973);
xor U18652 (N_18652,N_17756,N_16987);
or U18653 (N_18653,N_17628,N_17351);
or U18654 (N_18654,N_17218,N_17481);
xnor U18655 (N_18655,N_17943,N_17557);
nand U18656 (N_18656,N_16596,N_17558);
nor U18657 (N_18657,N_16735,N_17006);
xor U18658 (N_18658,N_16696,N_17547);
and U18659 (N_18659,N_17266,N_17790);
nand U18660 (N_18660,N_16985,N_17762);
nor U18661 (N_18661,N_17485,N_16796);
nor U18662 (N_18662,N_17093,N_17175);
nor U18663 (N_18663,N_17229,N_17657);
and U18664 (N_18664,N_17433,N_17908);
nand U18665 (N_18665,N_17769,N_17320);
nor U18666 (N_18666,N_17484,N_17463);
or U18667 (N_18667,N_16688,N_17296);
xor U18668 (N_18668,N_16646,N_16831);
nor U18669 (N_18669,N_17274,N_16887);
and U18670 (N_18670,N_17530,N_16799);
xnor U18671 (N_18671,N_16810,N_17824);
nand U18672 (N_18672,N_17829,N_16738);
xnor U18673 (N_18673,N_17721,N_16513);
nor U18674 (N_18674,N_17862,N_16973);
xor U18675 (N_18675,N_17382,N_16501);
or U18676 (N_18676,N_17592,N_17133);
xnor U18677 (N_18677,N_16500,N_17364);
xnor U18678 (N_18678,N_16785,N_17194);
and U18679 (N_18679,N_16592,N_16524);
nor U18680 (N_18680,N_17850,N_16802);
xnor U18681 (N_18681,N_17677,N_16893);
nand U18682 (N_18682,N_17037,N_17016);
and U18683 (N_18683,N_16619,N_16980);
nand U18684 (N_18684,N_17380,N_17998);
or U18685 (N_18685,N_17192,N_16919);
nand U18686 (N_18686,N_16647,N_17127);
xor U18687 (N_18687,N_16861,N_17860);
nand U18688 (N_18688,N_17114,N_16934);
or U18689 (N_18689,N_17972,N_16855);
xnor U18690 (N_18690,N_17329,N_17124);
nand U18691 (N_18691,N_17727,N_17897);
nand U18692 (N_18692,N_17396,N_16834);
or U18693 (N_18693,N_17520,N_17917);
or U18694 (N_18694,N_16721,N_16734);
nor U18695 (N_18695,N_16656,N_16804);
and U18696 (N_18696,N_17383,N_16502);
nand U18697 (N_18697,N_16511,N_16585);
or U18698 (N_18698,N_17418,N_16618);
xor U18699 (N_18699,N_17866,N_17861);
and U18700 (N_18700,N_17864,N_16777);
nor U18701 (N_18701,N_16780,N_16595);
nor U18702 (N_18702,N_17217,N_17906);
nand U18703 (N_18703,N_16509,N_16801);
nand U18704 (N_18704,N_17232,N_17997);
or U18705 (N_18705,N_17664,N_16564);
or U18706 (N_18706,N_17539,N_16769);
or U18707 (N_18707,N_17070,N_16957);
nand U18708 (N_18708,N_16700,N_17059);
nor U18709 (N_18709,N_16835,N_17205);
xor U18710 (N_18710,N_16571,N_16693);
and U18711 (N_18711,N_17513,N_17586);
nor U18712 (N_18712,N_17441,N_16594);
nand U18713 (N_18713,N_17032,N_17999);
or U18714 (N_18714,N_17934,N_17085);
or U18715 (N_18715,N_16765,N_17739);
xnor U18716 (N_18716,N_16539,N_17399);
and U18717 (N_18717,N_17614,N_16645);
xor U18718 (N_18718,N_16523,N_17806);
nand U18719 (N_18719,N_17242,N_16554);
and U18720 (N_18720,N_17247,N_17735);
or U18721 (N_18721,N_17584,N_17010);
and U18722 (N_18722,N_17515,N_17994);
nand U18723 (N_18723,N_17610,N_17731);
nor U18724 (N_18724,N_17025,N_17856);
or U18725 (N_18725,N_16949,N_16570);
nand U18726 (N_18726,N_17417,N_17452);
xnor U18727 (N_18727,N_16644,N_17585);
nand U18728 (N_18728,N_17116,N_16936);
and U18729 (N_18729,N_17816,N_17434);
nand U18730 (N_18730,N_17216,N_17933);
nor U18731 (N_18731,N_17222,N_17056);
and U18732 (N_18732,N_16854,N_16900);
nor U18733 (N_18733,N_16710,N_16979);
nand U18734 (N_18734,N_16803,N_17230);
nor U18735 (N_18735,N_17500,N_17705);
or U18736 (N_18736,N_17200,N_17825);
nand U18737 (N_18737,N_17629,N_16795);
nand U18738 (N_18738,N_16875,N_17076);
or U18739 (N_18739,N_17813,N_17251);
nand U18740 (N_18740,N_17690,N_16830);
or U18741 (N_18741,N_17384,N_16910);
nand U18742 (N_18742,N_17458,N_17669);
or U18743 (N_18743,N_17466,N_16712);
nor U18744 (N_18744,N_17950,N_16935);
and U18745 (N_18745,N_17446,N_17763);
and U18746 (N_18746,N_17665,N_16504);
xor U18747 (N_18747,N_17201,N_17496);
and U18748 (N_18748,N_17609,N_17745);
or U18749 (N_18749,N_16658,N_16842);
nand U18750 (N_18750,N_17053,N_16955);
nand U18751 (N_18751,N_16634,N_17210);
and U18752 (N_18752,N_16869,N_16852);
nand U18753 (N_18753,N_16592,N_16654);
or U18754 (N_18754,N_16832,N_17874);
and U18755 (N_18755,N_17968,N_16572);
or U18756 (N_18756,N_17937,N_17146);
nand U18757 (N_18757,N_17811,N_17786);
nor U18758 (N_18758,N_17561,N_17190);
nor U18759 (N_18759,N_16920,N_17826);
nand U18760 (N_18760,N_17678,N_17216);
and U18761 (N_18761,N_17106,N_16590);
nand U18762 (N_18762,N_17954,N_17970);
or U18763 (N_18763,N_17956,N_17354);
and U18764 (N_18764,N_17205,N_17518);
nor U18765 (N_18765,N_17391,N_17431);
nand U18766 (N_18766,N_17711,N_16914);
and U18767 (N_18767,N_16603,N_16553);
xnor U18768 (N_18768,N_17865,N_17438);
nor U18769 (N_18769,N_17961,N_16836);
and U18770 (N_18770,N_17367,N_17859);
nand U18771 (N_18771,N_16709,N_17242);
or U18772 (N_18772,N_17354,N_17942);
nand U18773 (N_18773,N_17327,N_17165);
nor U18774 (N_18774,N_16894,N_17387);
nand U18775 (N_18775,N_17235,N_16579);
nand U18776 (N_18776,N_17528,N_16788);
xnor U18777 (N_18777,N_16801,N_16751);
nand U18778 (N_18778,N_17627,N_17275);
or U18779 (N_18779,N_16832,N_17726);
nand U18780 (N_18780,N_17442,N_17797);
or U18781 (N_18781,N_16672,N_16924);
xor U18782 (N_18782,N_16733,N_17944);
and U18783 (N_18783,N_16871,N_17503);
nand U18784 (N_18784,N_17520,N_17905);
and U18785 (N_18785,N_17559,N_17192);
and U18786 (N_18786,N_17223,N_16821);
xor U18787 (N_18787,N_17960,N_17341);
or U18788 (N_18788,N_17223,N_17429);
nand U18789 (N_18789,N_17393,N_17719);
or U18790 (N_18790,N_17067,N_17447);
nor U18791 (N_18791,N_17752,N_17317);
nand U18792 (N_18792,N_17198,N_17590);
xnor U18793 (N_18793,N_16929,N_17941);
or U18794 (N_18794,N_17848,N_16890);
and U18795 (N_18795,N_17008,N_17335);
or U18796 (N_18796,N_16770,N_17775);
nor U18797 (N_18797,N_17106,N_16554);
and U18798 (N_18798,N_17703,N_16692);
nor U18799 (N_18799,N_16683,N_17240);
xnor U18800 (N_18800,N_16682,N_17770);
nor U18801 (N_18801,N_16728,N_17858);
xnor U18802 (N_18802,N_16782,N_17027);
xor U18803 (N_18803,N_16803,N_17663);
or U18804 (N_18804,N_16694,N_17361);
nand U18805 (N_18805,N_16809,N_17611);
nor U18806 (N_18806,N_17647,N_16853);
xnor U18807 (N_18807,N_16904,N_17577);
xor U18808 (N_18808,N_16801,N_17772);
nor U18809 (N_18809,N_17944,N_17644);
nor U18810 (N_18810,N_16544,N_17272);
xor U18811 (N_18811,N_16853,N_17668);
nand U18812 (N_18812,N_17914,N_16532);
or U18813 (N_18813,N_16779,N_17496);
nand U18814 (N_18814,N_17923,N_17593);
nand U18815 (N_18815,N_17955,N_17642);
and U18816 (N_18816,N_17269,N_17892);
and U18817 (N_18817,N_17606,N_17413);
and U18818 (N_18818,N_17775,N_17907);
xnor U18819 (N_18819,N_16562,N_17711);
or U18820 (N_18820,N_16890,N_16565);
or U18821 (N_18821,N_17434,N_17300);
or U18822 (N_18822,N_17901,N_17394);
nor U18823 (N_18823,N_17019,N_17401);
xnor U18824 (N_18824,N_16582,N_16789);
or U18825 (N_18825,N_17054,N_17927);
and U18826 (N_18826,N_16767,N_17971);
nand U18827 (N_18827,N_16833,N_17067);
or U18828 (N_18828,N_16780,N_16565);
nand U18829 (N_18829,N_16950,N_17667);
and U18830 (N_18830,N_16677,N_17409);
nand U18831 (N_18831,N_17155,N_17934);
xor U18832 (N_18832,N_17289,N_16927);
and U18833 (N_18833,N_16540,N_17271);
or U18834 (N_18834,N_17980,N_16845);
xor U18835 (N_18835,N_17098,N_17385);
xnor U18836 (N_18836,N_17361,N_17599);
xor U18837 (N_18837,N_17059,N_17472);
nor U18838 (N_18838,N_16505,N_17442);
xor U18839 (N_18839,N_16993,N_17898);
xor U18840 (N_18840,N_16848,N_17866);
or U18841 (N_18841,N_16544,N_16704);
nand U18842 (N_18842,N_16887,N_17338);
xnor U18843 (N_18843,N_17402,N_17231);
and U18844 (N_18844,N_17793,N_17813);
or U18845 (N_18845,N_17582,N_17273);
and U18846 (N_18846,N_16798,N_17858);
or U18847 (N_18847,N_16666,N_17079);
nor U18848 (N_18848,N_17334,N_17773);
and U18849 (N_18849,N_17669,N_16538);
nand U18850 (N_18850,N_16747,N_16595);
and U18851 (N_18851,N_17932,N_17850);
xnor U18852 (N_18852,N_16533,N_16583);
xor U18853 (N_18853,N_17218,N_16528);
and U18854 (N_18854,N_17530,N_17009);
xnor U18855 (N_18855,N_17134,N_16769);
and U18856 (N_18856,N_17156,N_17431);
nand U18857 (N_18857,N_17354,N_16690);
xor U18858 (N_18858,N_17677,N_17716);
nor U18859 (N_18859,N_17998,N_17814);
or U18860 (N_18860,N_17856,N_17075);
and U18861 (N_18861,N_17374,N_17430);
xor U18862 (N_18862,N_17483,N_16953);
or U18863 (N_18863,N_16701,N_17068);
or U18864 (N_18864,N_17727,N_17478);
or U18865 (N_18865,N_16890,N_16993);
and U18866 (N_18866,N_16641,N_16899);
xnor U18867 (N_18867,N_17473,N_17359);
nand U18868 (N_18868,N_17340,N_16927);
nand U18869 (N_18869,N_17362,N_17052);
nand U18870 (N_18870,N_17710,N_17938);
or U18871 (N_18871,N_17130,N_17229);
nand U18872 (N_18872,N_17329,N_17823);
nor U18873 (N_18873,N_17167,N_17924);
nand U18874 (N_18874,N_17506,N_16702);
and U18875 (N_18875,N_17264,N_17899);
nor U18876 (N_18876,N_16604,N_16535);
nand U18877 (N_18877,N_16738,N_17506);
nand U18878 (N_18878,N_16789,N_16977);
xnor U18879 (N_18879,N_17224,N_16667);
and U18880 (N_18880,N_16906,N_17478);
and U18881 (N_18881,N_17560,N_17201);
nor U18882 (N_18882,N_17250,N_16776);
nor U18883 (N_18883,N_16542,N_17362);
and U18884 (N_18884,N_17517,N_17877);
or U18885 (N_18885,N_16786,N_17553);
xor U18886 (N_18886,N_17129,N_16924);
and U18887 (N_18887,N_17450,N_17866);
and U18888 (N_18888,N_17505,N_17784);
nand U18889 (N_18889,N_16803,N_17697);
nor U18890 (N_18890,N_17499,N_17670);
or U18891 (N_18891,N_17869,N_16718);
xnor U18892 (N_18892,N_17198,N_16833);
and U18893 (N_18893,N_16758,N_17190);
nand U18894 (N_18894,N_16902,N_17128);
nand U18895 (N_18895,N_17249,N_16991);
nand U18896 (N_18896,N_16808,N_17957);
nand U18897 (N_18897,N_17674,N_17078);
and U18898 (N_18898,N_17300,N_17436);
nor U18899 (N_18899,N_17231,N_17505);
xor U18900 (N_18900,N_17188,N_16749);
xor U18901 (N_18901,N_17303,N_17540);
and U18902 (N_18902,N_16965,N_17148);
or U18903 (N_18903,N_16864,N_16637);
nor U18904 (N_18904,N_17581,N_16879);
and U18905 (N_18905,N_17767,N_17538);
nand U18906 (N_18906,N_17165,N_16629);
or U18907 (N_18907,N_17019,N_17292);
and U18908 (N_18908,N_16849,N_17817);
nand U18909 (N_18909,N_17569,N_16711);
xor U18910 (N_18910,N_16785,N_17071);
or U18911 (N_18911,N_16741,N_17877);
xnor U18912 (N_18912,N_17104,N_16772);
nor U18913 (N_18913,N_17323,N_16916);
and U18914 (N_18914,N_16740,N_17704);
or U18915 (N_18915,N_16654,N_17040);
xnor U18916 (N_18916,N_17645,N_17959);
nor U18917 (N_18917,N_16865,N_17184);
or U18918 (N_18918,N_16722,N_16656);
or U18919 (N_18919,N_17443,N_16710);
nor U18920 (N_18920,N_17420,N_17891);
or U18921 (N_18921,N_17469,N_17509);
nand U18922 (N_18922,N_16794,N_17737);
nor U18923 (N_18923,N_17700,N_17578);
and U18924 (N_18924,N_17570,N_16736);
and U18925 (N_18925,N_17715,N_17266);
or U18926 (N_18926,N_17383,N_16529);
and U18927 (N_18927,N_16641,N_17820);
xnor U18928 (N_18928,N_17124,N_16682);
or U18929 (N_18929,N_17425,N_17480);
nand U18930 (N_18930,N_17993,N_16929);
nor U18931 (N_18931,N_17480,N_17551);
nor U18932 (N_18932,N_16931,N_16827);
nor U18933 (N_18933,N_17378,N_17903);
and U18934 (N_18934,N_17664,N_16976);
xnor U18935 (N_18935,N_17487,N_17497);
and U18936 (N_18936,N_16930,N_17046);
xor U18937 (N_18937,N_17676,N_16573);
and U18938 (N_18938,N_17878,N_17368);
or U18939 (N_18939,N_17029,N_17510);
nor U18940 (N_18940,N_17214,N_17325);
nand U18941 (N_18941,N_17081,N_17857);
and U18942 (N_18942,N_17873,N_17641);
or U18943 (N_18943,N_16690,N_16961);
nand U18944 (N_18944,N_17972,N_17751);
nor U18945 (N_18945,N_16575,N_17750);
xor U18946 (N_18946,N_17020,N_17889);
and U18947 (N_18947,N_17665,N_16548);
and U18948 (N_18948,N_17908,N_17020);
nand U18949 (N_18949,N_17085,N_17357);
nor U18950 (N_18950,N_17782,N_17136);
and U18951 (N_18951,N_17466,N_16766);
xor U18952 (N_18952,N_17460,N_17440);
or U18953 (N_18953,N_17741,N_17257);
nand U18954 (N_18954,N_17883,N_17041);
nand U18955 (N_18955,N_17854,N_17312);
and U18956 (N_18956,N_16738,N_16524);
nor U18957 (N_18957,N_16755,N_16505);
and U18958 (N_18958,N_16801,N_17630);
nand U18959 (N_18959,N_17948,N_16561);
nor U18960 (N_18960,N_17736,N_17771);
or U18961 (N_18961,N_16685,N_17696);
nand U18962 (N_18962,N_17474,N_17859);
xnor U18963 (N_18963,N_16957,N_17892);
nor U18964 (N_18964,N_17205,N_17681);
xnor U18965 (N_18965,N_17467,N_16863);
nor U18966 (N_18966,N_17932,N_17574);
xor U18967 (N_18967,N_17764,N_17060);
and U18968 (N_18968,N_17555,N_16697);
or U18969 (N_18969,N_17600,N_17334);
and U18970 (N_18970,N_17587,N_17031);
and U18971 (N_18971,N_17590,N_17212);
xnor U18972 (N_18972,N_17365,N_17332);
or U18973 (N_18973,N_17826,N_17044);
or U18974 (N_18974,N_17436,N_16721);
nor U18975 (N_18975,N_17865,N_17506);
nand U18976 (N_18976,N_17699,N_16751);
or U18977 (N_18977,N_17989,N_17590);
nor U18978 (N_18978,N_16577,N_16739);
xnor U18979 (N_18979,N_17351,N_17214);
nor U18980 (N_18980,N_17587,N_17207);
nand U18981 (N_18981,N_17371,N_16738);
nand U18982 (N_18982,N_16977,N_17138);
nor U18983 (N_18983,N_16858,N_17299);
xnor U18984 (N_18984,N_17758,N_17557);
nor U18985 (N_18985,N_17126,N_16995);
and U18986 (N_18986,N_17155,N_16597);
xor U18987 (N_18987,N_17571,N_17734);
and U18988 (N_18988,N_16582,N_16947);
or U18989 (N_18989,N_16929,N_16840);
xnor U18990 (N_18990,N_17966,N_17300);
nor U18991 (N_18991,N_17751,N_17369);
nor U18992 (N_18992,N_16758,N_17367);
nand U18993 (N_18993,N_16867,N_17103);
xnor U18994 (N_18994,N_16759,N_17065);
xor U18995 (N_18995,N_17983,N_17849);
nand U18996 (N_18996,N_17218,N_16749);
and U18997 (N_18997,N_17999,N_16729);
and U18998 (N_18998,N_17365,N_17764);
or U18999 (N_18999,N_17522,N_16660);
or U19000 (N_19000,N_17730,N_16833);
nand U19001 (N_19001,N_17460,N_16989);
xnor U19002 (N_19002,N_16708,N_17751);
nor U19003 (N_19003,N_17735,N_17588);
xor U19004 (N_19004,N_16928,N_16919);
and U19005 (N_19005,N_17528,N_17703);
or U19006 (N_19006,N_16711,N_17834);
and U19007 (N_19007,N_17458,N_17613);
xor U19008 (N_19008,N_16565,N_17149);
xor U19009 (N_19009,N_17619,N_16794);
nor U19010 (N_19010,N_17737,N_17998);
nor U19011 (N_19011,N_17145,N_17214);
nor U19012 (N_19012,N_17050,N_17286);
nand U19013 (N_19013,N_17904,N_17267);
nor U19014 (N_19014,N_16671,N_17738);
or U19015 (N_19015,N_17045,N_17920);
or U19016 (N_19016,N_16664,N_17586);
and U19017 (N_19017,N_16772,N_16519);
and U19018 (N_19018,N_16559,N_17207);
or U19019 (N_19019,N_16593,N_17391);
nand U19020 (N_19020,N_17686,N_17333);
xor U19021 (N_19021,N_17037,N_17139);
nand U19022 (N_19022,N_16615,N_16995);
nand U19023 (N_19023,N_17805,N_16788);
nor U19024 (N_19024,N_17283,N_16844);
and U19025 (N_19025,N_16931,N_17922);
or U19026 (N_19026,N_17034,N_17153);
xor U19027 (N_19027,N_17877,N_17147);
or U19028 (N_19028,N_17758,N_17542);
nor U19029 (N_19029,N_17702,N_16835);
or U19030 (N_19030,N_17310,N_16767);
and U19031 (N_19031,N_17693,N_17790);
or U19032 (N_19032,N_17875,N_16846);
or U19033 (N_19033,N_17748,N_17371);
or U19034 (N_19034,N_17718,N_17190);
and U19035 (N_19035,N_17607,N_17111);
and U19036 (N_19036,N_16765,N_16540);
nand U19037 (N_19037,N_16539,N_16642);
and U19038 (N_19038,N_17267,N_17110);
or U19039 (N_19039,N_17868,N_17369);
nand U19040 (N_19040,N_17700,N_17161);
nand U19041 (N_19041,N_17450,N_17162);
nand U19042 (N_19042,N_17284,N_17512);
or U19043 (N_19043,N_17689,N_17157);
xnor U19044 (N_19044,N_17746,N_17044);
xnor U19045 (N_19045,N_17612,N_16538);
and U19046 (N_19046,N_16674,N_16500);
and U19047 (N_19047,N_17618,N_16728);
nand U19048 (N_19048,N_17776,N_16888);
or U19049 (N_19049,N_17713,N_17454);
nand U19050 (N_19050,N_16843,N_17442);
and U19051 (N_19051,N_17417,N_17790);
and U19052 (N_19052,N_17973,N_16539);
nor U19053 (N_19053,N_17273,N_16813);
and U19054 (N_19054,N_17967,N_16638);
nand U19055 (N_19055,N_17082,N_16735);
nand U19056 (N_19056,N_17552,N_16501);
xor U19057 (N_19057,N_16665,N_17323);
or U19058 (N_19058,N_16867,N_17258);
nand U19059 (N_19059,N_17047,N_17388);
xnor U19060 (N_19060,N_17012,N_17321);
nand U19061 (N_19061,N_17369,N_17014);
xnor U19062 (N_19062,N_16650,N_16619);
xnor U19063 (N_19063,N_17471,N_17681);
or U19064 (N_19064,N_17753,N_16875);
and U19065 (N_19065,N_16851,N_16837);
and U19066 (N_19066,N_17416,N_17198);
xnor U19067 (N_19067,N_16787,N_17602);
and U19068 (N_19068,N_17160,N_17467);
xor U19069 (N_19069,N_17377,N_17056);
or U19070 (N_19070,N_16952,N_16933);
and U19071 (N_19071,N_17174,N_17111);
xor U19072 (N_19072,N_17198,N_17387);
and U19073 (N_19073,N_17527,N_16639);
or U19074 (N_19074,N_17742,N_17908);
xnor U19075 (N_19075,N_17498,N_17316);
nor U19076 (N_19076,N_17408,N_17339);
or U19077 (N_19077,N_17518,N_17760);
nor U19078 (N_19078,N_17485,N_16627);
and U19079 (N_19079,N_17936,N_16990);
xnor U19080 (N_19080,N_17751,N_17437);
xor U19081 (N_19081,N_17372,N_17893);
or U19082 (N_19082,N_17895,N_17208);
and U19083 (N_19083,N_16541,N_17167);
nor U19084 (N_19084,N_17126,N_17968);
nor U19085 (N_19085,N_17467,N_17597);
xnor U19086 (N_19086,N_17712,N_17085);
nor U19087 (N_19087,N_16877,N_17520);
nand U19088 (N_19088,N_17255,N_17269);
xor U19089 (N_19089,N_16775,N_16563);
xor U19090 (N_19090,N_16959,N_17121);
xnor U19091 (N_19091,N_17753,N_17088);
and U19092 (N_19092,N_17233,N_17852);
and U19093 (N_19093,N_16594,N_16824);
and U19094 (N_19094,N_16520,N_17028);
xnor U19095 (N_19095,N_17388,N_17890);
or U19096 (N_19096,N_17103,N_16713);
or U19097 (N_19097,N_16955,N_16944);
xnor U19098 (N_19098,N_16674,N_17781);
xor U19099 (N_19099,N_16596,N_16774);
nand U19100 (N_19100,N_17168,N_17309);
xor U19101 (N_19101,N_16544,N_17399);
nand U19102 (N_19102,N_17284,N_17400);
nor U19103 (N_19103,N_17253,N_17056);
and U19104 (N_19104,N_16594,N_17266);
and U19105 (N_19105,N_16701,N_16924);
nand U19106 (N_19106,N_17602,N_17720);
or U19107 (N_19107,N_17678,N_17935);
nand U19108 (N_19108,N_17194,N_17680);
or U19109 (N_19109,N_16909,N_17315);
nor U19110 (N_19110,N_17583,N_16833);
or U19111 (N_19111,N_16773,N_17632);
nor U19112 (N_19112,N_17568,N_17128);
xor U19113 (N_19113,N_17873,N_16993);
nor U19114 (N_19114,N_17946,N_17325);
nor U19115 (N_19115,N_16550,N_17692);
or U19116 (N_19116,N_17316,N_17462);
nand U19117 (N_19117,N_17964,N_17744);
or U19118 (N_19118,N_17964,N_17148);
nand U19119 (N_19119,N_17134,N_16745);
and U19120 (N_19120,N_17042,N_16937);
nand U19121 (N_19121,N_16888,N_17333);
xnor U19122 (N_19122,N_17778,N_17387);
and U19123 (N_19123,N_16883,N_16616);
nand U19124 (N_19124,N_17882,N_17115);
nor U19125 (N_19125,N_17642,N_16918);
and U19126 (N_19126,N_17458,N_16845);
xnor U19127 (N_19127,N_17091,N_16947);
nand U19128 (N_19128,N_17238,N_17081);
nor U19129 (N_19129,N_17264,N_17909);
nor U19130 (N_19130,N_16792,N_16727);
and U19131 (N_19131,N_17451,N_17974);
or U19132 (N_19132,N_16771,N_16699);
and U19133 (N_19133,N_16952,N_16654);
xor U19134 (N_19134,N_16557,N_16743);
nor U19135 (N_19135,N_17904,N_17463);
xor U19136 (N_19136,N_17390,N_17645);
and U19137 (N_19137,N_17119,N_17935);
and U19138 (N_19138,N_17086,N_16863);
nand U19139 (N_19139,N_17771,N_17056);
nand U19140 (N_19140,N_17077,N_17637);
and U19141 (N_19141,N_16592,N_17514);
xor U19142 (N_19142,N_16712,N_16558);
nor U19143 (N_19143,N_16616,N_16730);
nor U19144 (N_19144,N_17450,N_17632);
nand U19145 (N_19145,N_16781,N_17160);
and U19146 (N_19146,N_17555,N_16517);
xnor U19147 (N_19147,N_17987,N_16862);
xor U19148 (N_19148,N_17385,N_17343);
xor U19149 (N_19149,N_17690,N_17531);
nand U19150 (N_19150,N_17324,N_16545);
nand U19151 (N_19151,N_16503,N_17652);
xnor U19152 (N_19152,N_17668,N_16518);
and U19153 (N_19153,N_16521,N_16857);
and U19154 (N_19154,N_16527,N_17505);
or U19155 (N_19155,N_16569,N_17362);
and U19156 (N_19156,N_16536,N_16901);
xor U19157 (N_19157,N_16731,N_17491);
nand U19158 (N_19158,N_17714,N_16880);
or U19159 (N_19159,N_17741,N_16675);
and U19160 (N_19160,N_17377,N_17100);
or U19161 (N_19161,N_17346,N_17504);
nor U19162 (N_19162,N_16954,N_17904);
xor U19163 (N_19163,N_17858,N_17310);
nor U19164 (N_19164,N_17286,N_17394);
or U19165 (N_19165,N_17625,N_17228);
and U19166 (N_19166,N_17018,N_17516);
and U19167 (N_19167,N_17895,N_16831);
nand U19168 (N_19168,N_16603,N_17638);
xor U19169 (N_19169,N_17628,N_17213);
or U19170 (N_19170,N_17773,N_17424);
or U19171 (N_19171,N_17564,N_17356);
nor U19172 (N_19172,N_17919,N_16596);
nand U19173 (N_19173,N_17172,N_16841);
nor U19174 (N_19174,N_17758,N_17845);
or U19175 (N_19175,N_17731,N_16598);
and U19176 (N_19176,N_17320,N_16823);
nand U19177 (N_19177,N_16630,N_16654);
nand U19178 (N_19178,N_17355,N_17886);
nor U19179 (N_19179,N_16658,N_16799);
nand U19180 (N_19180,N_17999,N_17059);
or U19181 (N_19181,N_16933,N_17051);
nor U19182 (N_19182,N_17425,N_17810);
nand U19183 (N_19183,N_16875,N_17847);
nand U19184 (N_19184,N_16589,N_17535);
xnor U19185 (N_19185,N_16879,N_17284);
nand U19186 (N_19186,N_17211,N_17752);
nor U19187 (N_19187,N_16724,N_17823);
and U19188 (N_19188,N_17449,N_17119);
nor U19189 (N_19189,N_16591,N_16559);
or U19190 (N_19190,N_16755,N_17865);
nor U19191 (N_19191,N_17205,N_17793);
nand U19192 (N_19192,N_16887,N_16654);
nand U19193 (N_19193,N_16869,N_17346);
xor U19194 (N_19194,N_16652,N_16625);
and U19195 (N_19195,N_17763,N_17796);
nor U19196 (N_19196,N_17342,N_17594);
xnor U19197 (N_19197,N_16628,N_17733);
xnor U19198 (N_19198,N_17435,N_16553);
or U19199 (N_19199,N_16818,N_16620);
nor U19200 (N_19200,N_17501,N_16793);
or U19201 (N_19201,N_17877,N_17889);
and U19202 (N_19202,N_17817,N_17270);
nor U19203 (N_19203,N_17836,N_17633);
nor U19204 (N_19204,N_17877,N_17046);
and U19205 (N_19205,N_16506,N_16959);
or U19206 (N_19206,N_17492,N_17630);
nor U19207 (N_19207,N_17667,N_17610);
and U19208 (N_19208,N_17673,N_17743);
or U19209 (N_19209,N_17316,N_16636);
nand U19210 (N_19210,N_17476,N_16905);
nand U19211 (N_19211,N_17596,N_17868);
or U19212 (N_19212,N_17877,N_17374);
or U19213 (N_19213,N_17372,N_16749);
and U19214 (N_19214,N_17255,N_17231);
nor U19215 (N_19215,N_16737,N_16953);
or U19216 (N_19216,N_17569,N_17143);
nor U19217 (N_19217,N_16548,N_17241);
or U19218 (N_19218,N_16753,N_16771);
nand U19219 (N_19219,N_17291,N_17575);
or U19220 (N_19220,N_17396,N_16732);
xor U19221 (N_19221,N_17428,N_17089);
nor U19222 (N_19222,N_17406,N_16916);
xnor U19223 (N_19223,N_16649,N_17517);
xor U19224 (N_19224,N_17767,N_16596);
nor U19225 (N_19225,N_17404,N_17243);
xor U19226 (N_19226,N_17628,N_17932);
nor U19227 (N_19227,N_16981,N_17870);
xnor U19228 (N_19228,N_16944,N_16956);
nand U19229 (N_19229,N_16971,N_17275);
nand U19230 (N_19230,N_17291,N_16731);
xor U19231 (N_19231,N_17979,N_17352);
nor U19232 (N_19232,N_16760,N_17598);
and U19233 (N_19233,N_17463,N_17690);
or U19234 (N_19234,N_17381,N_17021);
nor U19235 (N_19235,N_17156,N_17955);
and U19236 (N_19236,N_17127,N_17804);
nor U19237 (N_19237,N_16509,N_16791);
or U19238 (N_19238,N_17095,N_16542);
and U19239 (N_19239,N_17771,N_17884);
and U19240 (N_19240,N_16994,N_17799);
nand U19241 (N_19241,N_17403,N_17380);
and U19242 (N_19242,N_17743,N_17960);
or U19243 (N_19243,N_17067,N_17547);
xnor U19244 (N_19244,N_17423,N_17611);
xor U19245 (N_19245,N_16931,N_17745);
xor U19246 (N_19246,N_17645,N_17838);
nor U19247 (N_19247,N_16956,N_17072);
nand U19248 (N_19248,N_17238,N_16532);
nand U19249 (N_19249,N_16849,N_16992);
nand U19250 (N_19250,N_17483,N_16854);
xnor U19251 (N_19251,N_17241,N_17819);
or U19252 (N_19252,N_16689,N_17417);
or U19253 (N_19253,N_17335,N_17762);
nand U19254 (N_19254,N_16876,N_16635);
or U19255 (N_19255,N_17971,N_17986);
nand U19256 (N_19256,N_17104,N_17214);
and U19257 (N_19257,N_17736,N_17907);
and U19258 (N_19258,N_16872,N_16600);
nor U19259 (N_19259,N_17812,N_17405);
nor U19260 (N_19260,N_16824,N_16675);
or U19261 (N_19261,N_17721,N_16745);
xor U19262 (N_19262,N_16501,N_17288);
nor U19263 (N_19263,N_16688,N_16919);
nor U19264 (N_19264,N_17103,N_17942);
nand U19265 (N_19265,N_17844,N_16721);
nand U19266 (N_19266,N_16812,N_17131);
nand U19267 (N_19267,N_16602,N_17085);
xnor U19268 (N_19268,N_17631,N_17360);
or U19269 (N_19269,N_17104,N_17547);
xnor U19270 (N_19270,N_16703,N_17851);
and U19271 (N_19271,N_16635,N_17481);
nor U19272 (N_19272,N_16522,N_17924);
xnor U19273 (N_19273,N_17765,N_16632);
or U19274 (N_19274,N_17556,N_16859);
nand U19275 (N_19275,N_16937,N_16535);
xnor U19276 (N_19276,N_17452,N_16606);
nor U19277 (N_19277,N_17432,N_16678);
xnor U19278 (N_19278,N_17814,N_17325);
and U19279 (N_19279,N_17617,N_16739);
or U19280 (N_19280,N_16816,N_17508);
and U19281 (N_19281,N_17833,N_17013);
xnor U19282 (N_19282,N_17504,N_16676);
or U19283 (N_19283,N_17279,N_16725);
xor U19284 (N_19284,N_17464,N_17540);
nor U19285 (N_19285,N_17014,N_17500);
nand U19286 (N_19286,N_17414,N_16892);
xnor U19287 (N_19287,N_17632,N_16538);
nand U19288 (N_19288,N_17385,N_16843);
and U19289 (N_19289,N_17912,N_16896);
xor U19290 (N_19290,N_17387,N_17038);
and U19291 (N_19291,N_16810,N_17168);
and U19292 (N_19292,N_17624,N_17754);
and U19293 (N_19293,N_17079,N_17354);
xnor U19294 (N_19294,N_17005,N_16961);
or U19295 (N_19295,N_17134,N_17768);
nand U19296 (N_19296,N_17219,N_16662);
or U19297 (N_19297,N_16822,N_17621);
or U19298 (N_19298,N_16593,N_16711);
xor U19299 (N_19299,N_17272,N_17507);
nor U19300 (N_19300,N_16962,N_17822);
or U19301 (N_19301,N_17057,N_17968);
nor U19302 (N_19302,N_16751,N_16890);
and U19303 (N_19303,N_17368,N_17906);
nor U19304 (N_19304,N_17559,N_16859);
or U19305 (N_19305,N_16511,N_16535);
or U19306 (N_19306,N_17878,N_17469);
or U19307 (N_19307,N_16654,N_16677);
xnor U19308 (N_19308,N_16683,N_17822);
and U19309 (N_19309,N_17654,N_17823);
xnor U19310 (N_19310,N_17842,N_16596);
and U19311 (N_19311,N_16764,N_16822);
or U19312 (N_19312,N_16518,N_16827);
xor U19313 (N_19313,N_16764,N_17716);
nor U19314 (N_19314,N_16581,N_16547);
nand U19315 (N_19315,N_16680,N_17511);
and U19316 (N_19316,N_17047,N_16588);
nand U19317 (N_19317,N_17823,N_17426);
or U19318 (N_19318,N_17883,N_17969);
nor U19319 (N_19319,N_16813,N_17223);
nand U19320 (N_19320,N_17520,N_17838);
and U19321 (N_19321,N_17144,N_17529);
xnor U19322 (N_19322,N_16769,N_16725);
xnor U19323 (N_19323,N_17758,N_16800);
and U19324 (N_19324,N_17414,N_16802);
nand U19325 (N_19325,N_17590,N_17123);
xnor U19326 (N_19326,N_17637,N_17327);
nor U19327 (N_19327,N_16726,N_17586);
nand U19328 (N_19328,N_16703,N_16770);
nor U19329 (N_19329,N_17748,N_17743);
or U19330 (N_19330,N_17172,N_17566);
nand U19331 (N_19331,N_17546,N_17031);
and U19332 (N_19332,N_17810,N_17933);
or U19333 (N_19333,N_17878,N_17904);
nor U19334 (N_19334,N_17815,N_17363);
nor U19335 (N_19335,N_16935,N_17329);
and U19336 (N_19336,N_17380,N_16768);
or U19337 (N_19337,N_16505,N_16868);
xnor U19338 (N_19338,N_17172,N_16789);
nand U19339 (N_19339,N_16700,N_17082);
nand U19340 (N_19340,N_17430,N_16881);
and U19341 (N_19341,N_17381,N_17712);
nand U19342 (N_19342,N_17492,N_17262);
or U19343 (N_19343,N_17848,N_16664);
or U19344 (N_19344,N_17824,N_16724);
and U19345 (N_19345,N_16558,N_17949);
or U19346 (N_19346,N_16510,N_16930);
and U19347 (N_19347,N_17526,N_17923);
nand U19348 (N_19348,N_17564,N_17941);
or U19349 (N_19349,N_17937,N_16801);
or U19350 (N_19350,N_17506,N_17446);
xor U19351 (N_19351,N_16795,N_17070);
or U19352 (N_19352,N_17836,N_17750);
or U19353 (N_19353,N_17807,N_16630);
xor U19354 (N_19354,N_17475,N_17384);
xnor U19355 (N_19355,N_17423,N_17451);
and U19356 (N_19356,N_17660,N_16758);
nor U19357 (N_19357,N_17741,N_17462);
and U19358 (N_19358,N_17533,N_16694);
and U19359 (N_19359,N_17049,N_16792);
xnor U19360 (N_19360,N_17487,N_17035);
and U19361 (N_19361,N_17192,N_17826);
nand U19362 (N_19362,N_17933,N_17347);
and U19363 (N_19363,N_16610,N_16970);
nor U19364 (N_19364,N_17878,N_16900);
xnor U19365 (N_19365,N_17714,N_16942);
or U19366 (N_19366,N_16820,N_16984);
xnor U19367 (N_19367,N_17563,N_17337);
or U19368 (N_19368,N_17400,N_17089);
or U19369 (N_19369,N_16678,N_17897);
nand U19370 (N_19370,N_16633,N_17246);
and U19371 (N_19371,N_17562,N_17382);
or U19372 (N_19372,N_17864,N_17451);
and U19373 (N_19373,N_16819,N_16809);
xnor U19374 (N_19374,N_16941,N_16541);
nand U19375 (N_19375,N_17361,N_17638);
and U19376 (N_19376,N_17374,N_16833);
nand U19377 (N_19377,N_17646,N_17848);
or U19378 (N_19378,N_17220,N_17633);
and U19379 (N_19379,N_17626,N_17828);
xnor U19380 (N_19380,N_17754,N_17511);
nor U19381 (N_19381,N_16977,N_17017);
xor U19382 (N_19382,N_17689,N_17128);
nand U19383 (N_19383,N_17940,N_17778);
nand U19384 (N_19384,N_17801,N_17770);
and U19385 (N_19385,N_16652,N_16728);
or U19386 (N_19386,N_16606,N_17940);
and U19387 (N_19387,N_16784,N_17097);
nand U19388 (N_19388,N_17785,N_17457);
xnor U19389 (N_19389,N_17467,N_17030);
nand U19390 (N_19390,N_17852,N_17287);
nand U19391 (N_19391,N_17582,N_17474);
nor U19392 (N_19392,N_17689,N_16772);
and U19393 (N_19393,N_16751,N_17610);
and U19394 (N_19394,N_17031,N_17895);
nor U19395 (N_19395,N_17669,N_17307);
or U19396 (N_19396,N_17970,N_17390);
nor U19397 (N_19397,N_17567,N_16862);
or U19398 (N_19398,N_17451,N_17745);
or U19399 (N_19399,N_16623,N_17461);
xnor U19400 (N_19400,N_17318,N_17092);
and U19401 (N_19401,N_17285,N_17475);
and U19402 (N_19402,N_17803,N_17769);
nand U19403 (N_19403,N_17943,N_16614);
xor U19404 (N_19404,N_16971,N_16876);
nor U19405 (N_19405,N_17125,N_17290);
xnor U19406 (N_19406,N_17251,N_16548);
nor U19407 (N_19407,N_16654,N_16770);
nor U19408 (N_19408,N_17725,N_17990);
xor U19409 (N_19409,N_17839,N_16984);
and U19410 (N_19410,N_16691,N_17020);
nor U19411 (N_19411,N_17952,N_17090);
and U19412 (N_19412,N_16656,N_16866);
nor U19413 (N_19413,N_16900,N_17396);
and U19414 (N_19414,N_16544,N_16634);
xnor U19415 (N_19415,N_17190,N_17631);
nor U19416 (N_19416,N_17919,N_17331);
or U19417 (N_19417,N_16562,N_17746);
nand U19418 (N_19418,N_17537,N_17048);
and U19419 (N_19419,N_17461,N_17081);
or U19420 (N_19420,N_17651,N_17915);
xor U19421 (N_19421,N_17579,N_17377);
or U19422 (N_19422,N_17257,N_17154);
and U19423 (N_19423,N_17568,N_17698);
xor U19424 (N_19424,N_16629,N_17571);
nand U19425 (N_19425,N_16986,N_16567);
xnor U19426 (N_19426,N_17745,N_17065);
nand U19427 (N_19427,N_17479,N_16796);
or U19428 (N_19428,N_17966,N_17778);
xor U19429 (N_19429,N_17366,N_17785);
or U19430 (N_19430,N_16832,N_17996);
and U19431 (N_19431,N_17701,N_16582);
nand U19432 (N_19432,N_17069,N_17057);
and U19433 (N_19433,N_17587,N_17858);
xnor U19434 (N_19434,N_17412,N_16527);
or U19435 (N_19435,N_17005,N_17283);
or U19436 (N_19436,N_17743,N_17185);
nor U19437 (N_19437,N_17836,N_16773);
or U19438 (N_19438,N_17420,N_17259);
and U19439 (N_19439,N_16874,N_16967);
xor U19440 (N_19440,N_17045,N_17329);
or U19441 (N_19441,N_17200,N_17571);
nand U19442 (N_19442,N_17183,N_17656);
nand U19443 (N_19443,N_17470,N_17652);
xor U19444 (N_19444,N_17406,N_17631);
xnor U19445 (N_19445,N_17223,N_17681);
and U19446 (N_19446,N_17162,N_17565);
or U19447 (N_19447,N_17256,N_17060);
xnor U19448 (N_19448,N_16842,N_16613);
or U19449 (N_19449,N_16644,N_16656);
nand U19450 (N_19450,N_16855,N_17994);
or U19451 (N_19451,N_17679,N_17217);
or U19452 (N_19452,N_16813,N_17987);
or U19453 (N_19453,N_16615,N_16651);
or U19454 (N_19454,N_17475,N_17061);
and U19455 (N_19455,N_17528,N_17524);
xor U19456 (N_19456,N_16638,N_16945);
or U19457 (N_19457,N_17201,N_16590);
or U19458 (N_19458,N_16546,N_17370);
xnor U19459 (N_19459,N_17147,N_16849);
nand U19460 (N_19460,N_17223,N_17932);
nand U19461 (N_19461,N_17067,N_17514);
nor U19462 (N_19462,N_17687,N_17442);
or U19463 (N_19463,N_17064,N_17577);
xnor U19464 (N_19464,N_17962,N_17136);
and U19465 (N_19465,N_17399,N_16525);
and U19466 (N_19466,N_17989,N_16993);
nand U19467 (N_19467,N_16695,N_16869);
and U19468 (N_19468,N_16535,N_16978);
nor U19469 (N_19469,N_16878,N_17701);
nor U19470 (N_19470,N_17291,N_17431);
nor U19471 (N_19471,N_16536,N_16546);
nand U19472 (N_19472,N_17400,N_17280);
xor U19473 (N_19473,N_16961,N_17192);
xnor U19474 (N_19474,N_17571,N_17905);
and U19475 (N_19475,N_17518,N_17299);
or U19476 (N_19476,N_16857,N_16591);
nor U19477 (N_19477,N_16865,N_17525);
or U19478 (N_19478,N_17169,N_17554);
nand U19479 (N_19479,N_17808,N_16570);
and U19480 (N_19480,N_17385,N_17643);
or U19481 (N_19481,N_16952,N_17321);
nor U19482 (N_19482,N_17722,N_16905);
nand U19483 (N_19483,N_17709,N_16626);
and U19484 (N_19484,N_17809,N_17542);
nor U19485 (N_19485,N_17899,N_16901);
nand U19486 (N_19486,N_17712,N_17239);
and U19487 (N_19487,N_16602,N_16541);
or U19488 (N_19488,N_17895,N_16525);
nor U19489 (N_19489,N_17898,N_17188);
nand U19490 (N_19490,N_17881,N_16546);
or U19491 (N_19491,N_17511,N_17408);
xor U19492 (N_19492,N_17933,N_17427);
xor U19493 (N_19493,N_16923,N_16822);
xnor U19494 (N_19494,N_17267,N_17242);
nor U19495 (N_19495,N_16999,N_17605);
nand U19496 (N_19496,N_16917,N_16588);
xor U19497 (N_19497,N_16594,N_17327);
xnor U19498 (N_19498,N_17406,N_16645);
nand U19499 (N_19499,N_17498,N_17547);
and U19500 (N_19500,N_19087,N_18999);
or U19501 (N_19501,N_19141,N_19355);
xor U19502 (N_19502,N_18649,N_18804);
or U19503 (N_19503,N_19222,N_18602);
xnor U19504 (N_19504,N_18903,N_19429);
xnor U19505 (N_19505,N_19293,N_18078);
nand U19506 (N_19506,N_18071,N_18878);
nor U19507 (N_19507,N_18982,N_19108);
nor U19508 (N_19508,N_19367,N_18597);
nor U19509 (N_19509,N_18292,N_18591);
nand U19510 (N_19510,N_18509,N_19122);
xor U19511 (N_19511,N_18065,N_19482);
or U19512 (N_19512,N_18733,N_18297);
or U19513 (N_19513,N_18949,N_18623);
xnor U19514 (N_19514,N_18988,N_18951);
xnor U19515 (N_19515,N_19464,N_18407);
nor U19516 (N_19516,N_19033,N_19458);
xor U19517 (N_19517,N_19387,N_18183);
or U19518 (N_19518,N_18437,N_18717);
and U19519 (N_19519,N_18286,N_18149);
nor U19520 (N_19520,N_19342,N_18059);
xor U19521 (N_19521,N_19104,N_18116);
nor U19522 (N_19522,N_18004,N_19343);
xor U19523 (N_19523,N_18567,N_19148);
nand U19524 (N_19524,N_18352,N_18685);
and U19525 (N_19525,N_19045,N_18941);
and U19526 (N_19526,N_18443,N_19074);
xnor U19527 (N_19527,N_18690,N_18898);
nor U19528 (N_19528,N_18748,N_18674);
nand U19529 (N_19529,N_19176,N_18897);
nor U19530 (N_19530,N_18222,N_19016);
or U19531 (N_19531,N_18267,N_19421);
or U19532 (N_19532,N_19219,N_18345);
nor U19533 (N_19533,N_18115,N_19195);
nor U19534 (N_19534,N_18232,N_19172);
nor U19535 (N_19535,N_19204,N_19339);
or U19536 (N_19536,N_19182,N_18155);
or U19537 (N_19537,N_18347,N_18608);
nand U19538 (N_19538,N_18844,N_18343);
xor U19539 (N_19539,N_18719,N_18566);
xnor U19540 (N_19540,N_18138,N_18854);
xnor U19541 (N_19541,N_19466,N_18507);
xor U19542 (N_19542,N_18032,N_19375);
nand U19543 (N_19543,N_18745,N_19410);
nand U19544 (N_19544,N_18764,N_18360);
xor U19545 (N_19545,N_18819,N_19288);
nand U19546 (N_19546,N_19334,N_18724);
nand U19547 (N_19547,N_18568,N_18760);
xor U19548 (N_19548,N_18372,N_19450);
and U19549 (N_19549,N_18017,N_18758);
nor U19550 (N_19550,N_19237,N_18009);
or U19551 (N_19551,N_19143,N_18436);
or U19552 (N_19552,N_19208,N_18657);
nand U19553 (N_19553,N_18454,N_18179);
nor U19554 (N_19554,N_18508,N_18167);
or U19555 (N_19555,N_18787,N_18626);
or U19556 (N_19556,N_18850,N_18376);
nand U19557 (N_19557,N_18329,N_19457);
nor U19558 (N_19558,N_18170,N_18980);
xor U19559 (N_19559,N_19018,N_18381);
xnor U19560 (N_19560,N_19323,N_19459);
nand U19561 (N_19561,N_19191,N_19215);
or U19562 (N_19562,N_18575,N_18090);
or U19563 (N_19563,N_18186,N_19496);
or U19564 (N_19564,N_19202,N_18704);
and U19565 (N_19565,N_18853,N_18767);
or U19566 (N_19566,N_19260,N_18204);
nand U19567 (N_19567,N_18351,N_18257);
nor U19568 (N_19568,N_19242,N_18452);
or U19569 (N_19569,N_18755,N_19371);
and U19570 (N_19570,N_19370,N_18645);
xor U19571 (N_19571,N_19212,N_19118);
nor U19572 (N_19572,N_18293,N_19365);
and U19573 (N_19573,N_18556,N_18741);
and U19574 (N_19574,N_18814,N_19052);
nor U19575 (N_19575,N_19054,N_18552);
nor U19576 (N_19576,N_19093,N_18506);
nor U19577 (N_19577,N_19360,N_18934);
nor U19578 (N_19578,N_19063,N_18073);
or U19579 (N_19579,N_19325,N_18132);
nand U19580 (N_19580,N_18652,N_18650);
nor U19581 (N_19581,N_18024,N_19340);
xor U19582 (N_19582,N_18875,N_18808);
xor U19583 (N_19583,N_18963,N_18423);
and U19584 (N_19584,N_18694,N_18364);
and U19585 (N_19585,N_18341,N_19394);
or U19586 (N_19586,N_19043,N_18256);
or U19587 (N_19587,N_18890,N_18049);
and U19588 (N_19588,N_18740,N_18813);
nor U19589 (N_19589,N_19412,N_18832);
nor U19590 (N_19590,N_18043,N_18863);
nor U19591 (N_19591,N_19442,N_18069);
xnor U19592 (N_19592,N_18228,N_18405);
nor U19593 (N_19593,N_18722,N_18581);
xor U19594 (N_19594,N_18504,N_18203);
and U19595 (N_19595,N_19377,N_18448);
nand U19596 (N_19596,N_18205,N_19167);
or U19597 (N_19597,N_19249,N_19026);
xnor U19598 (N_19598,N_19292,N_18389);
xnor U19599 (N_19599,N_18337,N_18046);
nand U19600 (N_19600,N_18091,N_18783);
nor U19601 (N_19601,N_18060,N_18849);
nor U19602 (N_19602,N_18614,N_18265);
or U19603 (N_19603,N_18493,N_19432);
xor U19604 (N_19604,N_18971,N_18350);
nor U19605 (N_19605,N_18611,N_19161);
nor U19606 (N_19606,N_18595,N_18751);
xor U19607 (N_19607,N_19336,N_19356);
nand U19608 (N_19608,N_18217,N_18829);
nor U19609 (N_19609,N_19324,N_18672);
or U19610 (N_19610,N_18857,N_18089);
nand U19611 (N_19611,N_19048,N_18342);
xor U19612 (N_19612,N_18395,N_19424);
or U19613 (N_19613,N_18625,N_18646);
or U19614 (N_19614,N_18100,N_18867);
nand U19615 (N_19615,N_19477,N_18637);
xnor U19616 (N_19616,N_18632,N_18139);
or U19617 (N_19617,N_19083,N_19149);
nand U19618 (N_19618,N_18263,N_18067);
nand U19619 (N_19619,N_18268,N_18102);
or U19620 (N_19620,N_18770,N_18037);
and U19621 (N_19621,N_18831,N_18956);
and U19622 (N_19622,N_18369,N_18955);
nand U19623 (N_19623,N_19051,N_18848);
nand U19624 (N_19624,N_18413,N_18366);
xnor U19625 (N_19625,N_18430,N_18533);
or U19626 (N_19626,N_19270,N_18785);
nand U19627 (N_19627,N_18451,N_18280);
nor U19628 (N_19628,N_18230,N_18975);
nand U19629 (N_19629,N_18531,N_18406);
xnor U19630 (N_19630,N_19497,N_18966);
nand U19631 (N_19631,N_18334,N_18708);
nand U19632 (N_19632,N_18573,N_19453);
nand U19633 (N_19633,N_18207,N_19107);
nor U19634 (N_19634,N_18211,N_18972);
and U19635 (N_19635,N_18441,N_18718);
nand U19636 (N_19636,N_18696,N_19452);
and U19637 (N_19637,N_19455,N_18585);
xnor U19638 (N_19638,N_18039,N_18092);
xnor U19639 (N_19639,N_18969,N_18396);
xor U19640 (N_19640,N_18312,N_18712);
or U19641 (N_19641,N_19271,N_19247);
nand U19642 (N_19642,N_18750,N_19177);
nand U19643 (N_19643,N_19463,N_19368);
or U19644 (N_19644,N_19413,N_18492);
nor U19645 (N_19645,N_18553,N_19255);
nand U19646 (N_19646,N_18094,N_19447);
nor U19647 (N_19647,N_18475,N_19006);
or U19648 (N_19648,N_18148,N_18388);
or U19649 (N_19649,N_19162,N_18221);
nor U19650 (N_19650,N_19011,N_19337);
and U19651 (N_19651,N_19199,N_19160);
or U19652 (N_19652,N_18974,N_18066);
nand U19653 (N_19653,N_18001,N_18619);
and U19654 (N_19654,N_18855,N_18056);
xor U19655 (N_19655,N_18541,N_18973);
and U19656 (N_19656,N_18868,N_19415);
nor U19657 (N_19657,N_19192,N_19138);
nand U19658 (N_19658,N_19183,N_18803);
nor U19659 (N_19659,N_18140,N_19481);
or U19660 (N_19660,N_18296,N_18497);
nand U19661 (N_19661,N_18869,N_18737);
xnor U19662 (N_19662,N_19303,N_18308);
or U19663 (N_19663,N_18882,N_18738);
and U19664 (N_19664,N_18258,N_18251);
xnor U19665 (N_19665,N_18348,N_18911);
or U19666 (N_19666,N_18996,N_19042);
or U19667 (N_19667,N_18301,N_18967);
and U19668 (N_19668,N_18417,N_18404);
and U19669 (N_19669,N_18749,N_18387);
nand U19670 (N_19670,N_18599,N_19443);
and U19671 (N_19671,N_18466,N_18727);
nor U19672 (N_19672,N_18798,N_18261);
nand U19673 (N_19673,N_18063,N_18881);
nor U19674 (N_19674,N_18572,N_19210);
xnor U19675 (N_19675,N_18130,N_19297);
or U19676 (N_19676,N_19251,N_18768);
and U19677 (N_19677,N_18473,N_18682);
nor U19678 (N_19678,N_19099,N_19250);
xnor U19679 (N_19679,N_19446,N_18002);
or U19680 (N_19680,N_18047,N_18476);
xor U19681 (N_19681,N_18845,N_18870);
nor U19682 (N_19682,N_19106,N_18962);
nand U19683 (N_19683,N_18693,N_18933);
nor U19684 (N_19684,N_19475,N_19123);
xnor U19685 (N_19685,N_19105,N_19332);
nor U19686 (N_19686,N_19078,N_19069);
and U19687 (N_19687,N_18281,N_18784);
nor U19688 (N_19688,N_18121,N_18838);
or U19689 (N_19689,N_18333,N_18587);
xnor U19690 (N_19690,N_18182,N_18377);
nand U19691 (N_19691,N_19479,N_18805);
nor U19692 (N_19692,N_18948,N_18648);
or U19693 (N_19693,N_18924,N_18535);
nand U19694 (N_19694,N_19416,N_19312);
nor U19695 (N_19695,N_18335,N_18695);
nor U19696 (N_19696,N_19384,N_18667);
or U19697 (N_19697,N_18117,N_18519);
and U19698 (N_19698,N_18208,N_19163);
or U19699 (N_19699,N_18526,N_18841);
nand U19700 (N_19700,N_18467,N_18555);
and U19701 (N_19701,N_18818,N_18253);
and U19702 (N_19702,N_18926,N_18126);
and U19703 (N_19703,N_18311,N_18375);
nor U19704 (N_19704,N_18330,N_18422);
nor U19705 (N_19705,N_18057,N_19471);
and U19706 (N_19706,N_18615,N_18213);
or U19707 (N_19707,N_19094,N_18431);
and U19708 (N_19708,N_18522,N_19198);
and U19709 (N_19709,N_18198,N_18669);
xnor U19710 (N_19710,N_18936,N_18174);
or U19711 (N_19711,N_19351,N_18666);
and U19712 (N_19712,N_19281,N_19300);
and U19713 (N_19713,N_18282,N_18912);
nand U19714 (N_19714,N_18432,N_19248);
or U19715 (N_19715,N_18896,N_18639);
xnor U19716 (N_19716,N_19059,N_18363);
or U19717 (N_19717,N_19200,N_18630);
and U19718 (N_19718,N_18665,N_19269);
and U19719 (N_19719,N_19140,N_18970);
and U19720 (N_19720,N_18122,N_18013);
xor U19721 (N_19721,N_18479,N_18321);
xnor U19722 (N_19722,N_18763,N_19029);
and U19723 (N_19723,N_18252,N_18569);
or U19724 (N_19724,N_18921,N_18411);
xor U19725 (N_19725,N_19001,N_18144);
nand U19726 (N_19726,N_18908,N_19275);
or U19727 (N_19727,N_19493,N_18420);
or U19728 (N_19728,N_18496,N_18922);
xor U19729 (N_19729,N_18284,N_18168);
nand U19730 (N_19730,N_19154,N_19444);
xnor U19731 (N_19731,N_18447,N_18905);
xor U19732 (N_19732,N_18919,N_19056);
and U19733 (N_19733,N_19433,N_18275);
nand U19734 (N_19734,N_19430,N_18336);
nor U19735 (N_19735,N_19080,N_18302);
nor U19736 (N_19736,N_18914,N_19484);
nand U19737 (N_19737,N_18815,N_19346);
xor U19738 (N_19738,N_18641,N_18661);
nand U19739 (N_19739,N_19378,N_18414);
or U19740 (N_19740,N_19409,N_18861);
or U19741 (N_19741,N_19486,N_18033);
nand U19742 (N_19742,N_18817,N_18772);
nor U19743 (N_19743,N_18243,N_18957);
nor U19744 (N_19744,N_18344,N_18083);
and U19745 (N_19745,N_18673,N_18229);
nand U19746 (N_19746,N_19185,N_18315);
nor U19747 (N_19747,N_18513,N_18368);
nand U19748 (N_19748,N_18987,N_19091);
nor U19749 (N_19749,N_18491,N_18823);
nand U19750 (N_19750,N_18698,N_19095);
xor U19751 (N_19751,N_18021,N_18378);
or U19752 (N_19752,N_19025,N_18607);
and U19753 (N_19753,N_19012,N_18030);
xor U19754 (N_19754,N_18716,N_19400);
xor U19755 (N_19755,N_18393,N_19057);
nand U19756 (N_19756,N_18400,N_18548);
xor U19757 (N_19757,N_18754,N_19419);
nand U19758 (N_19758,N_19483,N_18482);
nor U19759 (N_19759,N_19448,N_18710);
nand U19760 (N_19760,N_18778,N_18169);
nand U19761 (N_19761,N_19239,N_19165);
nand U19762 (N_19762,N_18166,N_18899);
xor U19763 (N_19763,N_18088,N_18952);
xnor U19764 (N_19764,N_18384,N_18358);
nand U19765 (N_19765,N_18680,N_18574);
nand U19766 (N_19766,N_18821,N_18997);
nand U19767 (N_19767,N_18459,N_18495);
nor U19768 (N_19768,N_19285,N_18224);
xnor U19769 (N_19769,N_18559,N_18816);
or U19770 (N_19770,N_18489,N_19490);
nor U19771 (N_19771,N_18540,N_19120);
and U19772 (N_19772,N_18254,N_18040);
xor U19773 (N_19773,N_19206,N_19321);
or U19774 (N_19774,N_18488,N_18468);
and U19775 (N_19775,N_18285,N_19020);
or U19776 (N_19776,N_19358,N_19338);
nand U19777 (N_19777,N_19349,N_19014);
nand U19778 (N_19778,N_18291,N_18237);
nor U19779 (N_19779,N_19427,N_18000);
and U19780 (N_19780,N_18147,N_18199);
or U19781 (N_19781,N_18795,N_19456);
nor U19782 (N_19782,N_19070,N_19153);
nand U19783 (N_19783,N_19102,N_18189);
and U19784 (N_19784,N_18445,N_18739);
nand U19785 (N_19785,N_18554,N_18564);
nor U19786 (N_19786,N_19173,N_19060);
nor U19787 (N_19787,N_19273,N_19227);
nor U19788 (N_19788,N_18233,N_18686);
and U19789 (N_19789,N_18458,N_18915);
xnor U19790 (N_19790,N_19067,N_19175);
or U19791 (N_19791,N_18605,N_19041);
or U19792 (N_19792,N_18593,N_19055);
xor U19793 (N_19793,N_18723,N_18516);
xor U19794 (N_19794,N_18119,N_18141);
nand U19795 (N_19795,N_19276,N_18003);
or U19796 (N_19796,N_18391,N_19266);
nand U19797 (N_19797,N_18703,N_19372);
xnor U19798 (N_19798,N_19388,N_18638);
or U19799 (N_19799,N_19225,N_18779);
xnor U19800 (N_19800,N_18769,N_18108);
nor U19801 (N_19801,N_18429,N_19174);
nand U19802 (N_19802,N_19137,N_19000);
or U19803 (N_19803,N_18530,N_19119);
and U19804 (N_19804,N_18706,N_18434);
and U19805 (N_19805,N_18310,N_18631);
nand U19806 (N_19806,N_19362,N_18215);
nand U19807 (N_19807,N_18571,N_18048);
and U19808 (N_19808,N_19231,N_19470);
xnor U19809 (N_19809,N_18470,N_19098);
or U19810 (N_19810,N_18606,N_19142);
nor U19811 (N_19811,N_19385,N_18271);
and U19812 (N_19812,N_19036,N_18833);
nand U19813 (N_19813,N_18113,N_18676);
and U19814 (N_19814,N_18660,N_18227);
xor U19815 (N_19815,N_18807,N_18206);
xnor U19816 (N_19816,N_19401,N_19311);
nor U19817 (N_19817,N_18544,N_19217);
or U19818 (N_19818,N_18136,N_18181);
nand U19819 (N_19819,N_18220,N_19492);
and U19820 (N_19820,N_19062,N_18361);
nand U19821 (N_19821,N_19386,N_18156);
nand U19822 (N_19822,N_18986,N_18137);
or U19823 (N_19823,N_18025,N_18551);
nand U19824 (N_19824,N_19201,N_18776);
nor U19825 (N_19825,N_19193,N_18093);
nor U19826 (N_19826,N_18901,N_19309);
nand U19827 (N_19827,N_18886,N_19407);
and U19828 (N_19828,N_18225,N_18766);
nand U19829 (N_19829,N_18403,N_18339);
or U19830 (N_19830,N_18486,N_18762);
nor U19831 (N_19831,N_18985,N_19302);
or U19832 (N_19832,N_18323,N_19021);
nand U19833 (N_19833,N_19425,N_19007);
xnor U19834 (N_19834,N_19019,N_18386);
nor U19835 (N_19835,N_19478,N_19034);
nand U19836 (N_19836,N_18965,N_19079);
nor U19837 (N_19837,N_19090,N_18157);
xnor U19838 (N_19838,N_18129,N_18075);
nand U19839 (N_19839,N_19096,N_19053);
and U19840 (N_19840,N_18775,N_18190);
nor U19841 (N_19841,N_18523,N_18465);
or U19842 (N_19842,N_18994,N_19013);
nand U19843 (N_19843,N_18086,N_18629);
nand U19844 (N_19844,N_19115,N_18678);
and U19845 (N_19845,N_19223,N_19047);
xor U19846 (N_19846,N_18022,N_18702);
xnor U19847 (N_19847,N_18563,N_19254);
xnor U19848 (N_19848,N_18082,N_19030);
nand U19849 (N_19849,N_19218,N_19319);
or U19850 (N_19850,N_18528,N_18928);
nor U19851 (N_19851,N_18883,N_18027);
xor U19852 (N_19852,N_19329,N_18596);
xnor U19853 (N_19853,N_19129,N_18487);
nand U19854 (N_19854,N_19406,N_19272);
xor U19855 (N_19855,N_19116,N_19071);
or U19856 (N_19856,N_19089,N_18771);
nand U19857 (N_19857,N_19396,N_18683);
and U19858 (N_19858,N_18761,N_18565);
or U19859 (N_19859,N_18195,N_19188);
and U19860 (N_19860,N_18353,N_19044);
xnor U19861 (N_19861,N_19274,N_19414);
xnor U19862 (N_19862,N_18124,N_18537);
xnor U19863 (N_19863,N_18011,N_19124);
nand U19864 (N_19864,N_18991,N_18278);
xor U19865 (N_19865,N_18111,N_18610);
and U19866 (N_19866,N_18421,N_18651);
and U19867 (N_19867,N_19315,N_18038);
xnor U19868 (N_19868,N_19474,N_18185);
or U19869 (N_19869,N_19245,N_18884);
and U19870 (N_19870,N_19135,N_19305);
and U19871 (N_19871,N_19485,N_18735);
nand U19872 (N_19872,N_18120,N_18643);
and U19873 (N_19873,N_18520,N_19005);
nor U19874 (N_19874,N_18028,N_18549);
xnor U19875 (N_19875,N_19064,N_18159);
and U19876 (N_19876,N_19333,N_19263);
nand U19877 (N_19877,N_18354,N_19155);
nand U19878 (N_19878,N_18142,N_18677);
or U19879 (N_19879,N_18442,N_18932);
xnor U19880 (N_19880,N_18663,N_18759);
or U19881 (N_19881,N_18053,N_18154);
and U19882 (N_19882,N_18501,N_18864);
nand U19883 (N_19883,N_18438,N_19491);
xnor U19884 (N_19884,N_19133,N_18408);
nand U19885 (N_19885,N_18981,N_18834);
or U19886 (N_19886,N_18992,N_18462);
nor U19887 (N_19887,N_18907,N_18958);
nand U19888 (N_19888,N_19279,N_18357);
or U19889 (N_19889,N_18654,N_18484);
nand U19890 (N_19890,N_18542,N_18711);
or U19891 (N_19891,N_18847,N_18409);
nand U19892 (N_19892,N_18918,N_18675);
nor U19893 (N_19893,N_18945,N_19437);
or U19894 (N_19894,N_18525,N_18397);
nand U19895 (N_19895,N_18192,N_18830);
nor U19896 (N_19896,N_18791,N_19075);
and U19897 (N_19897,N_19328,N_18212);
nand U19898 (N_19898,N_19134,N_18913);
nand U19899 (N_19899,N_18692,N_19207);
or U19900 (N_19900,N_18008,N_19436);
and U19901 (N_19901,N_18527,N_19357);
nor U19902 (N_19902,N_19262,N_18960);
nor U19903 (N_19903,N_18536,N_18150);
or U19904 (N_19904,N_18935,N_19366);
and U19905 (N_19905,N_18782,N_18856);
nor U19906 (N_19906,N_18076,N_19258);
nand U19907 (N_19907,N_18852,N_18196);
and U19908 (N_19908,N_18515,N_18457);
nor U19909 (N_19909,N_19015,N_18440);
and U19910 (N_19910,N_19213,N_18968);
nor U19911 (N_19911,N_18790,N_18872);
nand U19912 (N_19912,N_19435,N_19289);
nor U19913 (N_19913,N_19441,N_19113);
nor U19914 (N_19914,N_18734,N_18664);
nor U19915 (N_19915,N_19345,N_18792);
xor U19916 (N_19916,N_18054,N_18172);
xor U19917 (N_19917,N_19128,N_19422);
and U19918 (N_19918,N_18604,N_18435);
nand U19919 (N_19919,N_18729,N_19290);
xnor U19920 (N_19920,N_18052,N_18382);
nor U19921 (N_19921,N_18401,N_19352);
and U19922 (N_19922,N_18851,N_18930);
xor U19923 (N_19923,N_18731,N_18780);
nor U19924 (N_19924,N_18290,N_19170);
or U19925 (N_19925,N_19379,N_18846);
or U19926 (N_19926,N_18545,N_18444);
and U19927 (N_19927,N_18107,N_18240);
nor U19928 (N_19928,N_19405,N_18586);
xor U19929 (N_19929,N_19283,N_18300);
nor U19930 (N_19930,N_18305,N_19296);
or U19931 (N_19931,N_18977,N_19299);
or U19932 (N_19932,N_18103,N_19027);
and U19933 (N_19933,N_18550,N_18662);
xor U19934 (N_19934,N_18627,N_19114);
nand U19935 (N_19935,N_18316,N_18180);
xor U19936 (N_19936,N_18720,N_18946);
or U19937 (N_19937,N_19348,N_18072);
xor U19938 (N_19938,N_19420,N_19194);
nand U19939 (N_19939,N_18356,N_18035);
and U19940 (N_19940,N_18279,N_18655);
and U19941 (N_19941,N_18510,N_19159);
and U19942 (N_19942,N_19390,N_18894);
xnor U19943 (N_19943,N_18023,N_18490);
xor U19944 (N_19944,N_18288,N_18295);
and U19945 (N_19945,N_19423,N_18416);
xor U19946 (N_19946,N_19028,N_19130);
nor U19947 (N_19947,N_18561,N_18026);
and U19948 (N_19948,N_19264,N_18029);
nor U19949 (N_19949,N_18609,N_18101);
or U19950 (N_19950,N_19278,N_18502);
nand U19951 (N_19951,N_18226,N_19327);
or U19952 (N_19952,N_18112,N_18270);
xor U19953 (N_19953,N_19449,N_18809);
xnor U19954 (N_19954,N_19313,N_18014);
xor U19955 (N_19955,N_19487,N_19009);
nand U19956 (N_19956,N_19181,N_18349);
or U19957 (N_19957,N_18244,N_18097);
or U19958 (N_19958,N_19139,N_18880);
and U19959 (N_19959,N_18276,N_18133);
and U19960 (N_19960,N_18633,N_18837);
nand U19961 (N_19961,N_18367,N_18178);
xnor U19962 (N_19962,N_18031,N_18151);
and U19963 (N_19963,N_18463,N_19039);
or U19964 (N_19964,N_19037,N_18560);
xor U19965 (N_19965,N_18653,N_18193);
nand U19966 (N_19966,N_18939,N_19151);
nand U19967 (N_19967,N_19232,N_18820);
nor U19968 (N_19968,N_18984,N_19010);
xor U19969 (N_19969,N_18732,N_18621);
nand U19970 (N_19970,N_19205,N_18681);
nand U19971 (N_19971,N_19438,N_19002);
xor U19972 (N_19972,N_19280,N_19180);
xnor U19973 (N_19973,N_19428,N_19284);
and U19974 (N_19974,N_18412,N_18892);
nor U19975 (N_19975,N_18505,N_18691);
nor U19976 (N_19976,N_18235,N_19373);
or U19977 (N_19977,N_19361,N_18248);
xnor U19978 (N_19978,N_18152,N_19032);
xnor U19979 (N_19979,N_19178,N_19197);
xor U19980 (N_19980,N_18143,N_18893);
nand U19981 (N_19981,N_18976,N_19439);
and U19982 (N_19982,N_19046,N_18659);
nand U19983 (N_19983,N_19168,N_18983);
or U19984 (N_19984,N_18843,N_18231);
or U19985 (N_19985,N_18472,N_18327);
xnor U19986 (N_19986,N_19434,N_18810);
nor U19987 (N_19987,N_18041,N_18383);
nor U19988 (N_19988,N_18398,N_18799);
nor U19989 (N_19989,N_18274,N_19101);
nor U19990 (N_19990,N_19189,N_19066);
or U19991 (N_19991,N_19469,N_18736);
nor U19992 (N_19992,N_19084,N_18579);
xnor U19993 (N_19993,N_19008,N_18162);
nand U19994 (N_19994,N_19224,N_19196);
nand U19995 (N_19995,N_18773,N_18616);
or U19996 (N_19996,N_19267,N_18765);
nand U19997 (N_19997,N_18188,N_18558);
or U19998 (N_19998,N_18415,N_18287);
xor U19999 (N_19999,N_18730,N_19150);
and U20000 (N_20000,N_18324,N_18824);
or U20001 (N_20001,N_18920,N_18910);
nand U20002 (N_20002,N_18862,N_19022);
xnor U20003 (N_20003,N_19341,N_18517);
nand U20004 (N_20004,N_18640,N_18061);
or U20005 (N_20005,N_18428,N_18889);
nand U20006 (N_20006,N_18427,N_18806);
nand U20007 (N_20007,N_18840,N_18828);
nor U20008 (N_20008,N_19461,N_19317);
nand U20009 (N_20009,N_19291,N_18464);
nand U20010 (N_20010,N_18583,N_18707);
nor U20011 (N_20011,N_18171,N_18697);
or U20012 (N_20012,N_18018,N_18449);
and U20013 (N_20013,N_18601,N_18929);
and U20014 (N_20014,N_18684,N_19476);
nand U20015 (N_20015,N_18410,N_19038);
or U20016 (N_20016,N_18216,N_18070);
and U20017 (N_20017,N_18995,N_18394);
nor U20018 (N_20018,N_18532,N_19145);
or U20019 (N_20019,N_19146,N_19144);
nor U20020 (N_20020,N_19229,N_19331);
nand U20021 (N_20021,N_18238,N_19017);
and U20022 (N_20022,N_18153,N_18392);
or U20023 (N_20023,N_18483,N_18455);
nor U20024 (N_20024,N_18954,N_19203);
nor U20025 (N_20025,N_18788,N_18104);
xor U20026 (N_20026,N_18209,N_19399);
xnor U20027 (N_20027,N_19049,N_19426);
or U20028 (N_20028,N_19209,N_18309);
nor U20029 (N_20029,N_18131,N_18084);
nand U20030 (N_20030,N_19326,N_18670);
nor U20031 (N_20031,N_18825,N_18628);
nor U20032 (N_20032,N_18570,N_18827);
nand U20033 (N_20033,N_19286,N_19294);
nor U20034 (N_20034,N_19076,N_19383);
nor U20035 (N_20035,N_18099,N_18953);
nor U20036 (N_20036,N_18603,N_18294);
nand U20037 (N_20037,N_18461,N_18580);
or U20038 (N_20038,N_19277,N_18744);
and U20039 (N_20039,N_18547,N_19480);
and U20040 (N_20040,N_18993,N_19003);
and U20041 (N_20041,N_18007,N_19156);
nand U20042 (N_20042,N_18546,N_18592);
xnor U20043 (N_20043,N_19228,N_18241);
and U20044 (N_20044,N_18636,N_18273);
nor U20045 (N_20045,N_18135,N_18106);
or U20046 (N_20046,N_18715,N_18647);
or U20047 (N_20047,N_18622,N_19082);
or U20048 (N_20048,N_18998,N_18051);
nor U20049 (N_20049,N_18259,N_18887);
xor U20050 (N_20050,N_18481,N_18752);
nand U20051 (N_20051,N_19152,N_18264);
xor U20052 (N_20052,N_19035,N_18642);
xor U20053 (N_20053,N_19023,N_19040);
nor U20054 (N_20054,N_19184,N_19179);
nor U20055 (N_20055,N_18689,N_18365);
and U20056 (N_20056,N_18362,N_18927);
xor U20057 (N_20057,N_18424,N_18098);
and U20058 (N_20058,N_18794,N_18010);
nand U20059 (N_20059,N_19240,N_18518);
and U20060 (N_20060,N_18266,N_19403);
xnor U20061 (N_20061,N_18277,N_19445);
nor U20062 (N_20062,N_19402,N_18865);
nor U20063 (N_20063,N_18786,N_18906);
or U20064 (N_20064,N_19088,N_18923);
and U20065 (N_20065,N_18223,N_19498);
xor U20066 (N_20066,N_18774,N_18164);
or U20067 (N_20067,N_19330,N_18811);
or U20068 (N_20068,N_18635,N_19220);
and U20069 (N_20069,N_18426,N_18080);
or U20070 (N_20070,N_19126,N_19253);
and U20071 (N_20071,N_19235,N_18524);
nor U20072 (N_20072,N_19131,N_19233);
or U20073 (N_20073,N_19127,N_18317);
and U20074 (N_20074,N_18283,N_18331);
nand U20075 (N_20075,N_18081,N_18521);
or U20076 (N_20076,N_19353,N_18726);
nor U20077 (N_20077,N_18634,N_18247);
nor U20078 (N_20078,N_19316,N_19221);
xor U20079 (N_20079,N_18990,N_19190);
nor U20080 (N_20080,N_18019,N_18909);
nor U20081 (N_20081,N_19374,N_18503);
or U20082 (N_20082,N_18163,N_18842);
xnor U20083 (N_20083,N_18118,N_19308);
nand U20084 (N_20084,N_18068,N_18200);
and U20085 (N_20085,N_18860,N_18836);
nand U20086 (N_20086,N_19454,N_18624);
xnor U20087 (N_20087,N_18015,N_19304);
nand U20088 (N_20088,N_18239,N_18658);
xnor U20089 (N_20089,N_18402,N_18006);
and U20090 (N_20090,N_18876,N_19230);
or U20091 (N_20091,N_18218,N_18879);
and U20092 (N_20092,N_19499,N_19241);
or U20093 (N_20093,N_19295,N_19359);
and U20094 (N_20094,N_18781,N_19214);
nand U20095 (N_20095,N_19468,N_18757);
and U20096 (N_20096,N_18399,N_19136);
nor U20097 (N_20097,N_18557,N_18020);
and U20098 (N_20098,N_18858,N_18161);
xor U20099 (N_20099,N_19467,N_19268);
and U20100 (N_20100,N_19320,N_18777);
nand U20101 (N_20101,N_18989,N_18700);
nand U20102 (N_20102,N_18979,N_18874);
nor U20103 (N_20103,N_19100,N_18789);
nand U20104 (N_20104,N_18456,N_18793);
and U20105 (N_20105,N_18346,N_19252);
xnor U20106 (N_20106,N_19397,N_18134);
nor U20107 (N_20107,N_19169,N_18425);
and U20108 (N_20108,N_19246,N_18687);
xnor U20109 (N_20109,N_18871,N_18679);
nand U20110 (N_20110,N_18045,N_18562);
xnor U20111 (N_20111,N_18314,N_19301);
nor U20112 (N_20112,N_19440,N_18197);
or U20113 (N_20113,N_18477,N_19259);
xor U20114 (N_20114,N_18618,N_19363);
or U20115 (N_20115,N_18110,N_18146);
nor U20116 (N_20116,N_18902,N_18801);
xnor U20117 (N_20117,N_18688,N_19211);
and U20118 (N_20118,N_18714,N_19097);
or U20119 (N_20119,N_18937,N_18797);
xnor U20120 (N_20120,N_19472,N_18313);
xnor U20121 (N_20121,N_19236,N_18877);
or U20122 (N_20122,N_19318,N_18042);
nand U20123 (N_20123,N_19494,N_18600);
or U20124 (N_20124,N_19226,N_18371);
nor U20125 (N_20125,N_19171,N_18105);
nand U20126 (N_20126,N_18584,N_18613);
xor U20127 (N_20127,N_18590,N_18187);
and U20128 (N_20128,N_18594,N_19418);
and U20129 (N_20129,N_19382,N_18538);
and U20130 (N_20130,N_19489,N_18917);
nor U20131 (N_20131,N_18380,N_19369);
xor U20132 (N_20132,N_18034,N_19347);
xnor U20133 (N_20133,N_18753,N_18055);
or U20134 (N_20134,N_18320,N_18262);
or U20135 (N_20135,N_18184,N_19376);
xor U20136 (N_20136,N_18742,N_18620);
xor U20137 (N_20137,N_19166,N_19404);
xnor U20138 (N_20138,N_18176,N_18701);
xor U20139 (N_20139,N_18474,N_19081);
xor U20140 (N_20140,N_18328,N_18539);
and U20141 (N_20141,N_19391,N_18900);
nor U20142 (N_20142,N_19073,N_19310);
or U20143 (N_20143,N_18885,N_18866);
nor U20144 (N_20144,N_18500,N_19109);
xor U20145 (N_20145,N_18895,N_19132);
xnor U20146 (N_20146,N_18298,N_18096);
nand U20147 (N_20147,N_18450,N_19065);
nor U20148 (N_20148,N_18095,N_18125);
nor U20149 (N_20149,N_18077,N_18191);
nor U20150 (N_20150,N_18165,N_18940);
or U20151 (N_20151,N_18127,N_18577);
and U20152 (N_20152,N_18644,N_18576);
nand U20153 (N_20153,N_18812,N_18289);
or U20154 (N_20154,N_19495,N_18950);
nand U20155 (N_20155,N_18756,N_19186);
xor U20156 (N_20156,N_18419,N_18160);
nand U20157 (N_20157,N_18123,N_18446);
nand U20158 (N_20158,N_18891,N_18058);
nor U20159 (N_20159,N_19158,N_18085);
nor U20160 (N_20160,N_19261,N_18534);
or U20161 (N_20161,N_18699,N_19187);
xnor U20162 (N_20162,N_19110,N_18036);
nand U20163 (N_20163,N_18938,N_18826);
xor U20164 (N_20164,N_18978,N_19354);
nor U20165 (N_20165,N_19111,N_19117);
and U20166 (N_20166,N_18005,N_19086);
xnor U20167 (N_20167,N_19488,N_19335);
xor U20168 (N_20168,N_18947,N_18234);
nor U20169 (N_20169,N_18322,N_19395);
or U20170 (N_20170,N_19314,N_19216);
xnor U20171 (N_20171,N_18210,N_18325);
nor U20172 (N_20172,N_18109,N_18873);
nand U20173 (N_20173,N_18390,N_18959);
or U20174 (N_20174,N_19381,N_19451);
and U20175 (N_20175,N_19103,N_19238);
nor U20176 (N_20176,N_18433,N_19004);
nor U20177 (N_20177,N_19431,N_18064);
nand U20178 (N_20178,N_18725,N_18249);
nor U20179 (N_20179,N_18074,N_18385);
nand U20180 (N_20180,N_18469,N_19072);
and U20181 (N_20181,N_19462,N_19408);
xnor U20182 (N_20182,N_19465,N_18326);
nor U20183 (N_20183,N_19244,N_19322);
or U20184 (N_20184,N_18050,N_18859);
nor U20185 (N_20185,N_19298,N_18272);
and U20186 (N_20186,N_19306,N_19350);
or U20187 (N_20187,N_18964,N_18529);
and U20188 (N_20188,N_18012,N_18478);
nand U20189 (N_20189,N_18016,N_18318);
and U20190 (N_20190,N_18177,N_18194);
and U20191 (N_20191,N_18839,N_18904);
nand U20192 (N_20192,N_18338,N_18485);
nand U20193 (N_20193,N_18668,N_19380);
and U20194 (N_20194,N_18418,N_18471);
nor U20195 (N_20195,N_18582,N_18079);
xnor U20196 (N_20196,N_18480,N_18944);
and U20197 (N_20197,N_19344,N_18747);
xor U20198 (N_20198,N_18511,N_18822);
xor U20199 (N_20199,N_19092,N_18514);
xnor U20200 (N_20200,N_18269,N_18460);
and U20201 (N_20201,N_18304,N_19050);
xor U20202 (N_20202,N_19125,N_18588);
nor U20203 (N_20203,N_19389,N_18671);
or U20204 (N_20204,N_19460,N_18961);
xnor U20205 (N_20205,N_18589,N_18543);
nand U20206 (N_20206,N_18114,N_18340);
or U20207 (N_20207,N_18373,N_18796);
and U20208 (N_20208,N_18925,N_18236);
and U20209 (N_20209,N_18374,N_19061);
nand U20210 (N_20210,N_19392,N_18512);
xnor U20211 (N_20211,N_18800,N_18219);
or U20212 (N_20212,N_19068,N_19085);
xnor U20213 (N_20213,N_19257,N_18728);
or U20214 (N_20214,N_19307,N_19287);
or U20215 (N_20215,N_18453,N_18370);
nor U20216 (N_20216,N_18612,N_18260);
and U20217 (N_20217,N_18743,N_19164);
or U20218 (N_20218,N_19024,N_18498);
nor U20219 (N_20219,N_18158,N_18598);
xor U20220 (N_20220,N_18943,N_18250);
and U20221 (N_20221,N_18245,N_19234);
or U20222 (N_20222,N_18128,N_18303);
or U20223 (N_20223,N_18617,N_19411);
or U20224 (N_20224,N_18379,N_18246);
and U20225 (N_20225,N_18494,N_18802);
or U20226 (N_20226,N_18705,N_18242);
or U20227 (N_20227,N_19265,N_19473);
xor U20228 (N_20228,N_18746,N_19157);
or U20229 (N_20229,N_19256,N_18319);
xor U20230 (N_20230,N_18439,N_18307);
nand U20231 (N_20231,N_19031,N_18359);
xor U20232 (N_20232,N_18299,N_18835);
or U20233 (N_20233,N_18044,N_19058);
xnor U20234 (N_20234,N_18332,N_19398);
or U20235 (N_20235,N_18656,N_18175);
and U20236 (N_20236,N_18201,N_18255);
and U20237 (N_20237,N_19243,N_19077);
and U20238 (N_20238,N_18931,N_18888);
nand U20239 (N_20239,N_19147,N_18087);
nor U20240 (N_20240,N_18499,N_18916);
xor U20241 (N_20241,N_19282,N_18942);
and U20242 (N_20242,N_19417,N_18173);
or U20243 (N_20243,N_18721,N_18713);
xnor U20244 (N_20244,N_19393,N_19112);
nor U20245 (N_20245,N_18214,N_19364);
nand U20246 (N_20246,N_18202,N_19121);
nor U20247 (N_20247,N_18709,N_18306);
and U20248 (N_20248,N_18355,N_18062);
and U20249 (N_20249,N_18578,N_18145);
nor U20250 (N_20250,N_19028,N_19267);
xor U20251 (N_20251,N_18100,N_18765);
nor U20252 (N_20252,N_18725,N_18232);
nand U20253 (N_20253,N_18778,N_18159);
or U20254 (N_20254,N_18872,N_18874);
or U20255 (N_20255,N_18502,N_19012);
nand U20256 (N_20256,N_18838,N_18977);
nor U20257 (N_20257,N_19189,N_18863);
and U20258 (N_20258,N_18317,N_19257);
nand U20259 (N_20259,N_18214,N_18387);
xor U20260 (N_20260,N_19092,N_19362);
xnor U20261 (N_20261,N_18659,N_19084);
or U20262 (N_20262,N_18680,N_18464);
or U20263 (N_20263,N_19429,N_19285);
nor U20264 (N_20264,N_18699,N_18877);
xnor U20265 (N_20265,N_18675,N_18204);
and U20266 (N_20266,N_18572,N_18292);
nor U20267 (N_20267,N_18972,N_18913);
xor U20268 (N_20268,N_18226,N_18054);
xnor U20269 (N_20269,N_18154,N_18874);
nand U20270 (N_20270,N_18607,N_18502);
xnor U20271 (N_20271,N_19240,N_19475);
and U20272 (N_20272,N_19261,N_18859);
xnor U20273 (N_20273,N_18224,N_18722);
nor U20274 (N_20274,N_18874,N_18533);
nand U20275 (N_20275,N_18655,N_19072);
xor U20276 (N_20276,N_18197,N_19458);
xnor U20277 (N_20277,N_18233,N_18840);
and U20278 (N_20278,N_19477,N_19023);
nor U20279 (N_20279,N_18200,N_19469);
xnor U20280 (N_20280,N_19382,N_18650);
xor U20281 (N_20281,N_18847,N_19059);
nor U20282 (N_20282,N_19205,N_18868);
and U20283 (N_20283,N_19228,N_18882);
and U20284 (N_20284,N_19035,N_18498);
and U20285 (N_20285,N_19010,N_18744);
nor U20286 (N_20286,N_18057,N_18534);
and U20287 (N_20287,N_18660,N_18929);
xor U20288 (N_20288,N_18814,N_18605);
nor U20289 (N_20289,N_18580,N_19036);
and U20290 (N_20290,N_19449,N_19499);
or U20291 (N_20291,N_18699,N_18193);
nand U20292 (N_20292,N_19059,N_18086);
xor U20293 (N_20293,N_19412,N_18703);
xnor U20294 (N_20294,N_18094,N_18045);
nand U20295 (N_20295,N_18570,N_18900);
nand U20296 (N_20296,N_18736,N_18094);
or U20297 (N_20297,N_18648,N_18079);
nand U20298 (N_20298,N_18676,N_18585);
nor U20299 (N_20299,N_18912,N_18567);
or U20300 (N_20300,N_18331,N_19416);
or U20301 (N_20301,N_18193,N_18606);
xor U20302 (N_20302,N_19301,N_18086);
nor U20303 (N_20303,N_18866,N_18187);
or U20304 (N_20304,N_19266,N_19349);
nor U20305 (N_20305,N_18000,N_19196);
and U20306 (N_20306,N_18644,N_19416);
xnor U20307 (N_20307,N_18796,N_18009);
nor U20308 (N_20308,N_19053,N_18233);
and U20309 (N_20309,N_18729,N_19233);
xor U20310 (N_20310,N_19282,N_19468);
xnor U20311 (N_20311,N_18743,N_18803);
or U20312 (N_20312,N_18281,N_18844);
nand U20313 (N_20313,N_19413,N_18616);
and U20314 (N_20314,N_18115,N_19061);
nand U20315 (N_20315,N_18745,N_18267);
or U20316 (N_20316,N_18817,N_19492);
and U20317 (N_20317,N_18674,N_18206);
nand U20318 (N_20318,N_18864,N_19331);
nand U20319 (N_20319,N_18099,N_18113);
nor U20320 (N_20320,N_18025,N_18084);
or U20321 (N_20321,N_19444,N_18132);
or U20322 (N_20322,N_18434,N_18679);
xor U20323 (N_20323,N_19484,N_18591);
nand U20324 (N_20324,N_19099,N_19322);
xnor U20325 (N_20325,N_19359,N_19196);
and U20326 (N_20326,N_19415,N_18150);
and U20327 (N_20327,N_19307,N_19090);
xor U20328 (N_20328,N_19200,N_18758);
nand U20329 (N_20329,N_18773,N_18530);
nand U20330 (N_20330,N_18085,N_18152);
xnor U20331 (N_20331,N_18172,N_18648);
and U20332 (N_20332,N_19218,N_18888);
nor U20333 (N_20333,N_18815,N_18479);
or U20334 (N_20334,N_18917,N_18272);
or U20335 (N_20335,N_18990,N_19072);
or U20336 (N_20336,N_18573,N_18858);
and U20337 (N_20337,N_18265,N_18658);
xnor U20338 (N_20338,N_18217,N_19222);
xor U20339 (N_20339,N_18270,N_18416);
nor U20340 (N_20340,N_19034,N_18481);
nor U20341 (N_20341,N_18247,N_18606);
or U20342 (N_20342,N_18607,N_18294);
xnor U20343 (N_20343,N_19220,N_18946);
or U20344 (N_20344,N_18477,N_18118);
or U20345 (N_20345,N_18877,N_19169);
and U20346 (N_20346,N_18284,N_18623);
nor U20347 (N_20347,N_19366,N_18436);
nor U20348 (N_20348,N_18321,N_18406);
xor U20349 (N_20349,N_19366,N_19373);
nor U20350 (N_20350,N_19401,N_18898);
xor U20351 (N_20351,N_18746,N_19124);
nand U20352 (N_20352,N_19197,N_19441);
and U20353 (N_20353,N_18028,N_19213);
and U20354 (N_20354,N_19463,N_19413);
nor U20355 (N_20355,N_18466,N_18815);
nand U20356 (N_20356,N_19226,N_18031);
and U20357 (N_20357,N_18657,N_18459);
nor U20358 (N_20358,N_18522,N_19338);
xor U20359 (N_20359,N_19309,N_18735);
and U20360 (N_20360,N_19212,N_19007);
and U20361 (N_20361,N_18765,N_18041);
xnor U20362 (N_20362,N_18958,N_18098);
and U20363 (N_20363,N_18473,N_18815);
nor U20364 (N_20364,N_18766,N_19126);
nor U20365 (N_20365,N_19427,N_18939);
nor U20366 (N_20366,N_19379,N_18778);
or U20367 (N_20367,N_18530,N_18924);
and U20368 (N_20368,N_18054,N_18474);
or U20369 (N_20369,N_19349,N_18533);
nor U20370 (N_20370,N_18690,N_18826);
nand U20371 (N_20371,N_19334,N_18560);
nand U20372 (N_20372,N_19496,N_18344);
or U20373 (N_20373,N_19367,N_19364);
nand U20374 (N_20374,N_19113,N_18880);
nor U20375 (N_20375,N_18958,N_19181);
nor U20376 (N_20376,N_18623,N_19174);
nand U20377 (N_20377,N_18584,N_18902);
nand U20378 (N_20378,N_18969,N_19323);
xor U20379 (N_20379,N_18729,N_18007);
nand U20380 (N_20380,N_18191,N_19266);
and U20381 (N_20381,N_18667,N_18832);
and U20382 (N_20382,N_18151,N_19390);
nand U20383 (N_20383,N_19399,N_19178);
nor U20384 (N_20384,N_18887,N_18715);
nand U20385 (N_20385,N_19275,N_18894);
or U20386 (N_20386,N_18439,N_18096);
nand U20387 (N_20387,N_18527,N_18778);
xnor U20388 (N_20388,N_18031,N_18120);
and U20389 (N_20389,N_18497,N_18160);
nor U20390 (N_20390,N_19225,N_19323);
and U20391 (N_20391,N_18113,N_19008);
or U20392 (N_20392,N_19397,N_18252);
nand U20393 (N_20393,N_18041,N_19013);
and U20394 (N_20394,N_19036,N_19206);
nor U20395 (N_20395,N_19083,N_19206);
and U20396 (N_20396,N_18460,N_18457);
nand U20397 (N_20397,N_18354,N_18522);
nor U20398 (N_20398,N_19463,N_19235);
and U20399 (N_20399,N_18239,N_19349);
xnor U20400 (N_20400,N_18514,N_19130);
or U20401 (N_20401,N_19471,N_18008);
or U20402 (N_20402,N_18710,N_19052);
and U20403 (N_20403,N_18473,N_18303);
nand U20404 (N_20404,N_18833,N_19151);
nand U20405 (N_20405,N_18511,N_18480);
nand U20406 (N_20406,N_19131,N_19174);
nand U20407 (N_20407,N_19487,N_19017);
and U20408 (N_20408,N_18916,N_19270);
nor U20409 (N_20409,N_18500,N_19489);
and U20410 (N_20410,N_18088,N_19431);
and U20411 (N_20411,N_18196,N_18531);
nand U20412 (N_20412,N_19481,N_18862);
nand U20413 (N_20413,N_18069,N_18462);
and U20414 (N_20414,N_18554,N_19125);
and U20415 (N_20415,N_18335,N_18384);
and U20416 (N_20416,N_18799,N_18857);
and U20417 (N_20417,N_19063,N_19078);
xnor U20418 (N_20418,N_19048,N_18660);
or U20419 (N_20419,N_19475,N_19137);
nor U20420 (N_20420,N_18205,N_19040);
nand U20421 (N_20421,N_18591,N_19144);
nand U20422 (N_20422,N_18052,N_19254);
nand U20423 (N_20423,N_18252,N_19110);
and U20424 (N_20424,N_19284,N_19417);
and U20425 (N_20425,N_18349,N_18742);
nor U20426 (N_20426,N_18214,N_18204);
nand U20427 (N_20427,N_18039,N_18082);
nor U20428 (N_20428,N_18850,N_19117);
or U20429 (N_20429,N_19132,N_19498);
xnor U20430 (N_20430,N_18282,N_19319);
or U20431 (N_20431,N_18411,N_18203);
xnor U20432 (N_20432,N_18628,N_18028);
xnor U20433 (N_20433,N_19061,N_19406);
and U20434 (N_20434,N_18320,N_19201);
or U20435 (N_20435,N_18243,N_18698);
nor U20436 (N_20436,N_18636,N_18872);
nand U20437 (N_20437,N_18514,N_18091);
nand U20438 (N_20438,N_18833,N_18921);
xnor U20439 (N_20439,N_18551,N_19333);
xor U20440 (N_20440,N_18411,N_18467);
or U20441 (N_20441,N_18946,N_19295);
or U20442 (N_20442,N_18343,N_19195);
or U20443 (N_20443,N_18792,N_18286);
or U20444 (N_20444,N_18554,N_18655);
xnor U20445 (N_20445,N_18972,N_19075);
nand U20446 (N_20446,N_18776,N_18169);
nand U20447 (N_20447,N_18142,N_18333);
nand U20448 (N_20448,N_18410,N_19326);
or U20449 (N_20449,N_19311,N_19198);
and U20450 (N_20450,N_18249,N_19238);
and U20451 (N_20451,N_18637,N_18427);
xor U20452 (N_20452,N_18161,N_18791);
or U20453 (N_20453,N_18155,N_18808);
nor U20454 (N_20454,N_19268,N_18749);
nand U20455 (N_20455,N_18888,N_19328);
and U20456 (N_20456,N_18896,N_18029);
nor U20457 (N_20457,N_19328,N_19467);
nor U20458 (N_20458,N_18627,N_18154);
nor U20459 (N_20459,N_19069,N_18741);
nor U20460 (N_20460,N_19208,N_18338);
and U20461 (N_20461,N_19402,N_18748);
xor U20462 (N_20462,N_18614,N_19495);
or U20463 (N_20463,N_18285,N_19494);
or U20464 (N_20464,N_18415,N_19314);
or U20465 (N_20465,N_19452,N_19268);
or U20466 (N_20466,N_18686,N_19480);
and U20467 (N_20467,N_18094,N_19323);
xnor U20468 (N_20468,N_19236,N_18927);
xor U20469 (N_20469,N_19499,N_19441);
nor U20470 (N_20470,N_18249,N_19105);
nand U20471 (N_20471,N_18356,N_18548);
nand U20472 (N_20472,N_18407,N_18675);
and U20473 (N_20473,N_19354,N_18557);
nand U20474 (N_20474,N_19063,N_18245);
nor U20475 (N_20475,N_18022,N_19190);
xor U20476 (N_20476,N_18886,N_19255);
nand U20477 (N_20477,N_18653,N_18197);
nor U20478 (N_20478,N_19430,N_19462);
xnor U20479 (N_20479,N_18842,N_18815);
nand U20480 (N_20480,N_19191,N_18747);
xnor U20481 (N_20481,N_19083,N_18235);
and U20482 (N_20482,N_18338,N_18236);
nor U20483 (N_20483,N_18307,N_18172);
and U20484 (N_20484,N_18772,N_18479);
or U20485 (N_20485,N_18041,N_18882);
xnor U20486 (N_20486,N_19067,N_18296);
nor U20487 (N_20487,N_18387,N_18170);
or U20488 (N_20488,N_18008,N_18004);
nor U20489 (N_20489,N_18628,N_19057);
or U20490 (N_20490,N_18062,N_18807);
nand U20491 (N_20491,N_19028,N_18874);
and U20492 (N_20492,N_19042,N_19093);
nor U20493 (N_20493,N_19131,N_18742);
nor U20494 (N_20494,N_18892,N_18772);
nand U20495 (N_20495,N_18733,N_18234);
nand U20496 (N_20496,N_18313,N_19460);
xnor U20497 (N_20497,N_18231,N_19301);
nor U20498 (N_20498,N_19464,N_18854);
nand U20499 (N_20499,N_18009,N_18820);
nor U20500 (N_20500,N_18544,N_18668);
and U20501 (N_20501,N_19138,N_18862);
nor U20502 (N_20502,N_18551,N_18697);
or U20503 (N_20503,N_19388,N_18528);
nand U20504 (N_20504,N_18723,N_18431);
and U20505 (N_20505,N_18163,N_18601);
nor U20506 (N_20506,N_19036,N_18743);
or U20507 (N_20507,N_19080,N_19009);
or U20508 (N_20508,N_18934,N_18424);
nand U20509 (N_20509,N_19316,N_19137);
nor U20510 (N_20510,N_18253,N_18498);
or U20511 (N_20511,N_18873,N_18610);
nand U20512 (N_20512,N_18065,N_18319);
nor U20513 (N_20513,N_18554,N_18993);
or U20514 (N_20514,N_18055,N_19232);
xnor U20515 (N_20515,N_19277,N_18633);
and U20516 (N_20516,N_18658,N_18550);
and U20517 (N_20517,N_18687,N_18050);
or U20518 (N_20518,N_18770,N_19266);
xnor U20519 (N_20519,N_18856,N_18348);
and U20520 (N_20520,N_19093,N_18355);
and U20521 (N_20521,N_18842,N_18373);
xor U20522 (N_20522,N_18015,N_18945);
and U20523 (N_20523,N_19013,N_18222);
and U20524 (N_20524,N_18259,N_19410);
xnor U20525 (N_20525,N_19020,N_18017);
xor U20526 (N_20526,N_18934,N_18037);
and U20527 (N_20527,N_18069,N_18420);
nor U20528 (N_20528,N_18363,N_18696);
or U20529 (N_20529,N_18536,N_18518);
or U20530 (N_20530,N_18700,N_18360);
xor U20531 (N_20531,N_19382,N_19185);
xor U20532 (N_20532,N_18193,N_18072);
nor U20533 (N_20533,N_18574,N_19405);
nor U20534 (N_20534,N_18376,N_19138);
or U20535 (N_20535,N_18744,N_18201);
nand U20536 (N_20536,N_18790,N_18130);
xor U20537 (N_20537,N_19440,N_19100);
xnor U20538 (N_20538,N_18554,N_18479);
and U20539 (N_20539,N_19333,N_19304);
nand U20540 (N_20540,N_18305,N_19340);
nor U20541 (N_20541,N_18584,N_18784);
nand U20542 (N_20542,N_18752,N_18727);
and U20543 (N_20543,N_18371,N_18190);
and U20544 (N_20544,N_19484,N_19166);
nand U20545 (N_20545,N_18465,N_18818);
nor U20546 (N_20546,N_19392,N_18811);
nor U20547 (N_20547,N_18760,N_19292);
nand U20548 (N_20548,N_18425,N_18748);
and U20549 (N_20549,N_18744,N_18729);
or U20550 (N_20550,N_19343,N_19176);
nor U20551 (N_20551,N_18538,N_18560);
nand U20552 (N_20552,N_18776,N_19205);
nand U20553 (N_20553,N_18232,N_18110);
and U20554 (N_20554,N_19397,N_18542);
nand U20555 (N_20555,N_18987,N_19127);
or U20556 (N_20556,N_19310,N_18530);
nand U20557 (N_20557,N_19235,N_19278);
nand U20558 (N_20558,N_18878,N_18787);
or U20559 (N_20559,N_18118,N_18696);
nand U20560 (N_20560,N_18740,N_18285);
and U20561 (N_20561,N_18302,N_18394);
and U20562 (N_20562,N_19127,N_18055);
and U20563 (N_20563,N_18862,N_18062);
nand U20564 (N_20564,N_18211,N_18988);
nor U20565 (N_20565,N_19158,N_18733);
nor U20566 (N_20566,N_19347,N_18392);
nor U20567 (N_20567,N_18296,N_19402);
nor U20568 (N_20568,N_18460,N_18945);
nor U20569 (N_20569,N_18476,N_18959);
xnor U20570 (N_20570,N_19188,N_19212);
nand U20571 (N_20571,N_18103,N_18641);
or U20572 (N_20572,N_18922,N_19126);
nand U20573 (N_20573,N_18201,N_18036);
or U20574 (N_20574,N_19383,N_18513);
and U20575 (N_20575,N_18008,N_19078);
xor U20576 (N_20576,N_19046,N_19008);
and U20577 (N_20577,N_19291,N_18536);
nor U20578 (N_20578,N_19396,N_18627);
nor U20579 (N_20579,N_19138,N_19209);
nand U20580 (N_20580,N_18168,N_19143);
nand U20581 (N_20581,N_19346,N_19005);
nor U20582 (N_20582,N_18753,N_18512);
or U20583 (N_20583,N_18123,N_19285);
nor U20584 (N_20584,N_18841,N_18158);
xnor U20585 (N_20585,N_18688,N_19498);
nand U20586 (N_20586,N_18202,N_18516);
and U20587 (N_20587,N_18762,N_18029);
nor U20588 (N_20588,N_18929,N_18477);
nor U20589 (N_20589,N_18987,N_19088);
nor U20590 (N_20590,N_18366,N_19334);
or U20591 (N_20591,N_19345,N_18507);
or U20592 (N_20592,N_19420,N_18516);
nor U20593 (N_20593,N_18388,N_18219);
xor U20594 (N_20594,N_18367,N_18248);
and U20595 (N_20595,N_18857,N_18944);
xnor U20596 (N_20596,N_18441,N_19430);
nor U20597 (N_20597,N_18198,N_18822);
and U20598 (N_20598,N_18689,N_19316);
nand U20599 (N_20599,N_19222,N_18957);
and U20600 (N_20600,N_18257,N_18719);
nor U20601 (N_20601,N_19439,N_19077);
nor U20602 (N_20602,N_18854,N_19277);
nand U20603 (N_20603,N_19376,N_18164);
or U20604 (N_20604,N_18153,N_18113);
nor U20605 (N_20605,N_18932,N_18637);
or U20606 (N_20606,N_18237,N_18419);
nand U20607 (N_20607,N_18740,N_18094);
xor U20608 (N_20608,N_19246,N_19033);
and U20609 (N_20609,N_18198,N_18724);
xor U20610 (N_20610,N_18203,N_18784);
nand U20611 (N_20611,N_19389,N_18473);
nor U20612 (N_20612,N_19216,N_19151);
or U20613 (N_20613,N_18295,N_18177);
or U20614 (N_20614,N_18042,N_18573);
and U20615 (N_20615,N_18058,N_19123);
xnor U20616 (N_20616,N_18222,N_18653);
and U20617 (N_20617,N_18639,N_18455);
nand U20618 (N_20618,N_18291,N_18315);
and U20619 (N_20619,N_18007,N_18770);
xnor U20620 (N_20620,N_18436,N_18409);
xor U20621 (N_20621,N_18551,N_18645);
and U20622 (N_20622,N_19209,N_18680);
nand U20623 (N_20623,N_18296,N_18926);
xnor U20624 (N_20624,N_18470,N_19172);
nor U20625 (N_20625,N_18531,N_18083);
and U20626 (N_20626,N_18292,N_18229);
and U20627 (N_20627,N_18579,N_18306);
nor U20628 (N_20628,N_18903,N_18960);
nor U20629 (N_20629,N_18057,N_18319);
nor U20630 (N_20630,N_18518,N_18538);
or U20631 (N_20631,N_19478,N_19050);
xnor U20632 (N_20632,N_19053,N_19331);
nand U20633 (N_20633,N_18373,N_18652);
and U20634 (N_20634,N_18122,N_19306);
nor U20635 (N_20635,N_18027,N_19003);
xor U20636 (N_20636,N_19462,N_19071);
and U20637 (N_20637,N_18020,N_18451);
or U20638 (N_20638,N_18867,N_18290);
or U20639 (N_20639,N_19253,N_18134);
xor U20640 (N_20640,N_19275,N_18601);
nand U20641 (N_20641,N_19173,N_19261);
and U20642 (N_20642,N_18555,N_19059);
xnor U20643 (N_20643,N_18832,N_18795);
or U20644 (N_20644,N_19390,N_19448);
or U20645 (N_20645,N_18197,N_18722);
nand U20646 (N_20646,N_18846,N_18877);
nand U20647 (N_20647,N_18866,N_18717);
nor U20648 (N_20648,N_18353,N_18852);
xnor U20649 (N_20649,N_19166,N_18422);
nor U20650 (N_20650,N_18693,N_19025);
or U20651 (N_20651,N_19296,N_18805);
nor U20652 (N_20652,N_18395,N_18067);
xor U20653 (N_20653,N_19211,N_18514);
xor U20654 (N_20654,N_18559,N_18703);
xnor U20655 (N_20655,N_19409,N_19310);
or U20656 (N_20656,N_18999,N_18916);
and U20657 (N_20657,N_19185,N_18269);
or U20658 (N_20658,N_18410,N_18880);
and U20659 (N_20659,N_18016,N_19005);
xor U20660 (N_20660,N_18107,N_18953);
and U20661 (N_20661,N_19445,N_18644);
xor U20662 (N_20662,N_19144,N_19348);
and U20663 (N_20663,N_18100,N_19148);
nor U20664 (N_20664,N_19110,N_18367);
and U20665 (N_20665,N_18847,N_18179);
nor U20666 (N_20666,N_19054,N_18369);
and U20667 (N_20667,N_18740,N_18107);
nor U20668 (N_20668,N_18851,N_18343);
nand U20669 (N_20669,N_19283,N_18494);
nor U20670 (N_20670,N_18162,N_18203);
nor U20671 (N_20671,N_18061,N_19104);
or U20672 (N_20672,N_18798,N_19164);
xnor U20673 (N_20673,N_18308,N_18146);
nor U20674 (N_20674,N_18390,N_18847);
and U20675 (N_20675,N_18588,N_18979);
or U20676 (N_20676,N_18356,N_19130);
and U20677 (N_20677,N_19418,N_19395);
or U20678 (N_20678,N_18318,N_19037);
xor U20679 (N_20679,N_19106,N_18686);
nand U20680 (N_20680,N_18171,N_19154);
nand U20681 (N_20681,N_18602,N_18069);
xor U20682 (N_20682,N_18245,N_18491);
or U20683 (N_20683,N_18674,N_18520);
nand U20684 (N_20684,N_18079,N_18964);
nor U20685 (N_20685,N_18912,N_18403);
and U20686 (N_20686,N_18329,N_18307);
xor U20687 (N_20687,N_18980,N_18376);
xor U20688 (N_20688,N_19395,N_18742);
nand U20689 (N_20689,N_18394,N_18291);
nor U20690 (N_20690,N_18485,N_19232);
nor U20691 (N_20691,N_19395,N_19357);
or U20692 (N_20692,N_18336,N_18059);
nor U20693 (N_20693,N_18178,N_19123);
or U20694 (N_20694,N_18391,N_18978);
and U20695 (N_20695,N_19484,N_18380);
or U20696 (N_20696,N_18142,N_18676);
and U20697 (N_20697,N_19263,N_18572);
nand U20698 (N_20698,N_18868,N_18380);
and U20699 (N_20699,N_18032,N_18435);
or U20700 (N_20700,N_18243,N_19002);
or U20701 (N_20701,N_18968,N_18256);
and U20702 (N_20702,N_18729,N_19253);
xor U20703 (N_20703,N_18846,N_18565);
nor U20704 (N_20704,N_18806,N_19150);
and U20705 (N_20705,N_19163,N_18144);
and U20706 (N_20706,N_18464,N_18231);
or U20707 (N_20707,N_19438,N_18194);
and U20708 (N_20708,N_18079,N_18000);
and U20709 (N_20709,N_19062,N_18541);
xnor U20710 (N_20710,N_19114,N_18443);
nand U20711 (N_20711,N_19239,N_18179);
nand U20712 (N_20712,N_19192,N_18657);
or U20713 (N_20713,N_18895,N_19039);
nor U20714 (N_20714,N_18152,N_18552);
xor U20715 (N_20715,N_18148,N_18905);
nand U20716 (N_20716,N_18438,N_19483);
and U20717 (N_20717,N_18835,N_18534);
nor U20718 (N_20718,N_19157,N_19346);
nor U20719 (N_20719,N_18635,N_18376);
xnor U20720 (N_20720,N_19089,N_18464);
xor U20721 (N_20721,N_19198,N_18978);
or U20722 (N_20722,N_19281,N_19088);
and U20723 (N_20723,N_19457,N_19043);
xor U20724 (N_20724,N_18206,N_18358);
xnor U20725 (N_20725,N_18051,N_18731);
nand U20726 (N_20726,N_18912,N_18993);
nand U20727 (N_20727,N_18360,N_18842);
and U20728 (N_20728,N_18360,N_18529);
nor U20729 (N_20729,N_19184,N_18273);
nor U20730 (N_20730,N_19190,N_18914);
nor U20731 (N_20731,N_18198,N_18582);
or U20732 (N_20732,N_18027,N_18997);
nor U20733 (N_20733,N_18792,N_18595);
or U20734 (N_20734,N_19264,N_19183);
or U20735 (N_20735,N_19075,N_18117);
or U20736 (N_20736,N_18721,N_18750);
or U20737 (N_20737,N_18729,N_18584);
nor U20738 (N_20738,N_18358,N_19397);
nand U20739 (N_20739,N_18835,N_18439);
and U20740 (N_20740,N_19490,N_18685);
or U20741 (N_20741,N_18816,N_18794);
nand U20742 (N_20742,N_19069,N_18734);
or U20743 (N_20743,N_18448,N_18433);
nor U20744 (N_20744,N_18718,N_18561);
nand U20745 (N_20745,N_18956,N_19428);
or U20746 (N_20746,N_18593,N_18111);
xnor U20747 (N_20747,N_18352,N_18925);
nor U20748 (N_20748,N_18954,N_18189);
or U20749 (N_20749,N_19139,N_18683);
and U20750 (N_20750,N_18836,N_18180);
or U20751 (N_20751,N_19486,N_18077);
and U20752 (N_20752,N_18399,N_19006);
xnor U20753 (N_20753,N_18327,N_19219);
xor U20754 (N_20754,N_18752,N_18137);
and U20755 (N_20755,N_19040,N_18071);
nor U20756 (N_20756,N_18459,N_19092);
xor U20757 (N_20757,N_18982,N_18042);
and U20758 (N_20758,N_18519,N_19063);
or U20759 (N_20759,N_19037,N_18064);
or U20760 (N_20760,N_19261,N_18739);
xor U20761 (N_20761,N_18972,N_18183);
or U20762 (N_20762,N_18512,N_19079);
nand U20763 (N_20763,N_18940,N_19420);
or U20764 (N_20764,N_18218,N_19335);
nor U20765 (N_20765,N_19211,N_18956);
and U20766 (N_20766,N_18314,N_19304);
xnor U20767 (N_20767,N_18580,N_18667);
and U20768 (N_20768,N_18694,N_18067);
nor U20769 (N_20769,N_18206,N_19188);
xor U20770 (N_20770,N_18703,N_18821);
and U20771 (N_20771,N_18660,N_18397);
nor U20772 (N_20772,N_19479,N_19140);
nand U20773 (N_20773,N_19171,N_18905);
or U20774 (N_20774,N_18474,N_18693);
xnor U20775 (N_20775,N_18035,N_19031);
or U20776 (N_20776,N_18972,N_18921);
nand U20777 (N_20777,N_18847,N_18724);
nand U20778 (N_20778,N_18220,N_18614);
or U20779 (N_20779,N_18791,N_18520);
nand U20780 (N_20780,N_18629,N_19394);
xnor U20781 (N_20781,N_19304,N_18597);
and U20782 (N_20782,N_19157,N_18201);
and U20783 (N_20783,N_18880,N_18765);
and U20784 (N_20784,N_18370,N_18213);
nor U20785 (N_20785,N_18484,N_18196);
nor U20786 (N_20786,N_18344,N_18263);
xor U20787 (N_20787,N_19375,N_18785);
and U20788 (N_20788,N_19403,N_18979);
nand U20789 (N_20789,N_19006,N_18407);
xor U20790 (N_20790,N_18768,N_19293);
nor U20791 (N_20791,N_19207,N_19156);
or U20792 (N_20792,N_19301,N_18830);
nor U20793 (N_20793,N_19294,N_18413);
or U20794 (N_20794,N_18008,N_18749);
or U20795 (N_20795,N_18292,N_18811);
nor U20796 (N_20796,N_18474,N_18475);
nor U20797 (N_20797,N_18382,N_18082);
nor U20798 (N_20798,N_18110,N_19290);
and U20799 (N_20799,N_19253,N_18816);
and U20800 (N_20800,N_18784,N_18488);
nand U20801 (N_20801,N_18267,N_18127);
nand U20802 (N_20802,N_18955,N_18244);
nand U20803 (N_20803,N_18117,N_18872);
nand U20804 (N_20804,N_18426,N_19388);
and U20805 (N_20805,N_18341,N_18004);
nand U20806 (N_20806,N_19168,N_18546);
and U20807 (N_20807,N_18409,N_19291);
nand U20808 (N_20808,N_18003,N_18446);
nand U20809 (N_20809,N_18636,N_18026);
xor U20810 (N_20810,N_18892,N_19053);
xor U20811 (N_20811,N_18909,N_18537);
xor U20812 (N_20812,N_18681,N_19465);
xor U20813 (N_20813,N_18316,N_19017);
and U20814 (N_20814,N_19458,N_19392);
or U20815 (N_20815,N_18139,N_19329);
nand U20816 (N_20816,N_19358,N_18542);
nand U20817 (N_20817,N_19233,N_18293);
or U20818 (N_20818,N_18955,N_18156);
xor U20819 (N_20819,N_19134,N_18529);
or U20820 (N_20820,N_18782,N_19049);
and U20821 (N_20821,N_18919,N_18306);
nand U20822 (N_20822,N_18187,N_18816);
xnor U20823 (N_20823,N_18948,N_19459);
xnor U20824 (N_20824,N_19398,N_18019);
nor U20825 (N_20825,N_18856,N_18953);
xor U20826 (N_20826,N_18118,N_19020);
nor U20827 (N_20827,N_18191,N_18053);
nor U20828 (N_20828,N_18584,N_18472);
xor U20829 (N_20829,N_19253,N_18932);
and U20830 (N_20830,N_19213,N_18428);
and U20831 (N_20831,N_18011,N_18736);
and U20832 (N_20832,N_18468,N_18963);
and U20833 (N_20833,N_18715,N_19010);
nand U20834 (N_20834,N_18336,N_18869);
xor U20835 (N_20835,N_19203,N_18897);
and U20836 (N_20836,N_18980,N_18936);
nand U20837 (N_20837,N_18631,N_19161);
nand U20838 (N_20838,N_18509,N_18784);
nor U20839 (N_20839,N_18861,N_18835);
or U20840 (N_20840,N_19277,N_18240);
xor U20841 (N_20841,N_18068,N_18447);
xor U20842 (N_20842,N_18380,N_19193);
and U20843 (N_20843,N_18325,N_19320);
and U20844 (N_20844,N_19179,N_19227);
nor U20845 (N_20845,N_18923,N_18050);
nor U20846 (N_20846,N_19044,N_18613);
and U20847 (N_20847,N_19137,N_18333);
nor U20848 (N_20848,N_19275,N_18241);
and U20849 (N_20849,N_18827,N_18398);
or U20850 (N_20850,N_19188,N_18102);
xor U20851 (N_20851,N_18123,N_18892);
xnor U20852 (N_20852,N_19208,N_19202);
nand U20853 (N_20853,N_18557,N_18619);
or U20854 (N_20854,N_18070,N_18950);
or U20855 (N_20855,N_19421,N_19083);
or U20856 (N_20856,N_18271,N_19060);
and U20857 (N_20857,N_18747,N_18606);
xnor U20858 (N_20858,N_18490,N_18119);
nand U20859 (N_20859,N_18468,N_18800);
and U20860 (N_20860,N_19354,N_18455);
nor U20861 (N_20861,N_18922,N_19166);
nor U20862 (N_20862,N_18379,N_18352);
nor U20863 (N_20863,N_19218,N_18113);
nand U20864 (N_20864,N_18534,N_18635);
nand U20865 (N_20865,N_18561,N_18454);
nand U20866 (N_20866,N_18764,N_18834);
nand U20867 (N_20867,N_18799,N_19017);
nand U20868 (N_20868,N_18286,N_18423);
xnor U20869 (N_20869,N_18445,N_18485);
or U20870 (N_20870,N_18353,N_19024);
or U20871 (N_20871,N_18989,N_18886);
nand U20872 (N_20872,N_18680,N_18570);
xnor U20873 (N_20873,N_18114,N_19304);
nor U20874 (N_20874,N_18340,N_19370);
xnor U20875 (N_20875,N_19309,N_18071);
and U20876 (N_20876,N_18972,N_18717);
nor U20877 (N_20877,N_18002,N_18070);
nor U20878 (N_20878,N_18541,N_19006);
nor U20879 (N_20879,N_18801,N_18379);
or U20880 (N_20880,N_18599,N_18797);
nand U20881 (N_20881,N_19491,N_19027);
and U20882 (N_20882,N_18649,N_19406);
xnor U20883 (N_20883,N_19296,N_18268);
nand U20884 (N_20884,N_19352,N_18796);
xnor U20885 (N_20885,N_19186,N_18861);
nor U20886 (N_20886,N_19054,N_19336);
or U20887 (N_20887,N_18491,N_19403);
or U20888 (N_20888,N_19241,N_19345);
nor U20889 (N_20889,N_19414,N_19269);
and U20890 (N_20890,N_18061,N_18882);
nand U20891 (N_20891,N_19007,N_18380);
nor U20892 (N_20892,N_18629,N_18923);
nor U20893 (N_20893,N_18364,N_18690);
xor U20894 (N_20894,N_19234,N_19486);
xor U20895 (N_20895,N_18724,N_18955);
nand U20896 (N_20896,N_18731,N_18928);
nor U20897 (N_20897,N_18725,N_18356);
nand U20898 (N_20898,N_18351,N_18518);
nor U20899 (N_20899,N_18051,N_18138);
or U20900 (N_20900,N_18974,N_18242);
nor U20901 (N_20901,N_19337,N_19362);
or U20902 (N_20902,N_18046,N_18071);
or U20903 (N_20903,N_18015,N_19330);
nor U20904 (N_20904,N_18749,N_18453);
nor U20905 (N_20905,N_18567,N_18263);
or U20906 (N_20906,N_19316,N_18735);
nand U20907 (N_20907,N_18652,N_18683);
nand U20908 (N_20908,N_19145,N_18936);
and U20909 (N_20909,N_18739,N_18456);
nor U20910 (N_20910,N_18860,N_18808);
or U20911 (N_20911,N_19136,N_18321);
nand U20912 (N_20912,N_18273,N_18629);
xnor U20913 (N_20913,N_18074,N_18751);
nand U20914 (N_20914,N_19486,N_18836);
nand U20915 (N_20915,N_19086,N_19064);
or U20916 (N_20916,N_18216,N_18283);
nor U20917 (N_20917,N_18315,N_19329);
and U20918 (N_20918,N_19329,N_18346);
xor U20919 (N_20919,N_19037,N_18664);
nor U20920 (N_20920,N_18185,N_18288);
xnor U20921 (N_20921,N_18583,N_19424);
or U20922 (N_20922,N_18925,N_19224);
and U20923 (N_20923,N_18489,N_18304);
nor U20924 (N_20924,N_18663,N_18468);
nand U20925 (N_20925,N_18954,N_18001);
nand U20926 (N_20926,N_19195,N_18716);
xor U20927 (N_20927,N_18565,N_18682);
nand U20928 (N_20928,N_18917,N_18279);
xor U20929 (N_20929,N_18236,N_18115);
or U20930 (N_20930,N_19106,N_18651);
and U20931 (N_20931,N_18987,N_18018);
or U20932 (N_20932,N_18045,N_18047);
xor U20933 (N_20933,N_18022,N_18505);
or U20934 (N_20934,N_18234,N_18977);
and U20935 (N_20935,N_18268,N_18565);
nor U20936 (N_20936,N_18179,N_19309);
and U20937 (N_20937,N_18682,N_18431);
xor U20938 (N_20938,N_18475,N_19453);
or U20939 (N_20939,N_19454,N_18445);
and U20940 (N_20940,N_18000,N_18018);
and U20941 (N_20941,N_19248,N_19075);
or U20942 (N_20942,N_18160,N_19428);
nand U20943 (N_20943,N_18598,N_19346);
or U20944 (N_20944,N_19229,N_18710);
xnor U20945 (N_20945,N_18393,N_18186);
nor U20946 (N_20946,N_18582,N_19086);
xor U20947 (N_20947,N_19154,N_19224);
nor U20948 (N_20948,N_19215,N_19287);
xor U20949 (N_20949,N_19277,N_19356);
or U20950 (N_20950,N_18548,N_18651);
nor U20951 (N_20951,N_18642,N_18423);
nand U20952 (N_20952,N_19351,N_19052);
xor U20953 (N_20953,N_19040,N_18332);
nand U20954 (N_20954,N_19484,N_18926);
xor U20955 (N_20955,N_19128,N_19200);
xnor U20956 (N_20956,N_18314,N_18012);
nand U20957 (N_20957,N_18350,N_19000);
nand U20958 (N_20958,N_18754,N_19139);
or U20959 (N_20959,N_18119,N_19301);
xnor U20960 (N_20960,N_19286,N_19017);
nor U20961 (N_20961,N_18907,N_18688);
xor U20962 (N_20962,N_19084,N_18155);
and U20963 (N_20963,N_19258,N_18595);
or U20964 (N_20964,N_18856,N_18722);
nor U20965 (N_20965,N_18407,N_19295);
and U20966 (N_20966,N_18152,N_19011);
nand U20967 (N_20967,N_19042,N_18820);
xnor U20968 (N_20968,N_18750,N_18187);
or U20969 (N_20969,N_19436,N_19429);
or U20970 (N_20970,N_18761,N_18968);
nor U20971 (N_20971,N_18868,N_18946);
nor U20972 (N_20972,N_18208,N_19372);
nor U20973 (N_20973,N_18395,N_18315);
or U20974 (N_20974,N_18579,N_18534);
and U20975 (N_20975,N_19080,N_18305);
nor U20976 (N_20976,N_18068,N_19294);
nand U20977 (N_20977,N_18525,N_19096);
nand U20978 (N_20978,N_18958,N_18272);
or U20979 (N_20979,N_19235,N_19068);
nor U20980 (N_20980,N_18158,N_19484);
and U20981 (N_20981,N_18921,N_18859);
nor U20982 (N_20982,N_18250,N_19275);
and U20983 (N_20983,N_19179,N_18949);
xnor U20984 (N_20984,N_19483,N_19282);
and U20985 (N_20985,N_18283,N_18326);
and U20986 (N_20986,N_18034,N_18895);
nand U20987 (N_20987,N_18113,N_18738);
and U20988 (N_20988,N_18821,N_18440);
xnor U20989 (N_20989,N_19296,N_18864);
nor U20990 (N_20990,N_18733,N_18163);
nand U20991 (N_20991,N_18334,N_19397);
or U20992 (N_20992,N_19019,N_19260);
xor U20993 (N_20993,N_18896,N_19156);
and U20994 (N_20994,N_18385,N_18379);
and U20995 (N_20995,N_18896,N_19057);
nor U20996 (N_20996,N_19436,N_18235);
xnor U20997 (N_20997,N_19293,N_18931);
nor U20998 (N_20998,N_18427,N_18568);
nand U20999 (N_20999,N_19095,N_18928);
and U21000 (N_21000,N_19895,N_20748);
and U21001 (N_21001,N_20689,N_20629);
or U21002 (N_21002,N_19735,N_20188);
nor U21003 (N_21003,N_20347,N_20128);
xor U21004 (N_21004,N_19559,N_20270);
and U21005 (N_21005,N_20134,N_20093);
or U21006 (N_21006,N_20789,N_19812);
xor U21007 (N_21007,N_20126,N_19564);
nor U21008 (N_21008,N_20353,N_20011);
nor U21009 (N_21009,N_20842,N_20465);
nand U21010 (N_21010,N_20266,N_19623);
nand U21011 (N_21011,N_19641,N_20478);
and U21012 (N_21012,N_19971,N_20358);
xnor U21013 (N_21013,N_20575,N_20250);
xor U21014 (N_21014,N_20161,N_20367);
xor U21015 (N_21015,N_19916,N_20096);
and U21016 (N_21016,N_19508,N_20074);
nor U21017 (N_21017,N_19960,N_20483);
xnor U21018 (N_21018,N_19813,N_20534);
xnor U21019 (N_21019,N_19590,N_19838);
xnor U21020 (N_21020,N_20166,N_19532);
and U21021 (N_21021,N_20809,N_19968);
or U21022 (N_21022,N_20245,N_19789);
nor U21023 (N_21023,N_19702,N_19665);
xnor U21024 (N_21024,N_20261,N_20766);
nor U21025 (N_21025,N_20762,N_19673);
nor U21026 (N_21026,N_19739,N_20094);
nand U21027 (N_21027,N_19900,N_19983);
and U21028 (N_21028,N_19818,N_19915);
and U21029 (N_21029,N_19951,N_20324);
nor U21030 (N_21030,N_20743,N_19531);
nor U21031 (N_21031,N_19638,N_19529);
nand U21032 (N_21032,N_20559,N_20217);
or U21033 (N_21033,N_19947,N_19829);
nor U21034 (N_21034,N_20476,N_19862);
xnor U21035 (N_21035,N_20276,N_20426);
nor U21036 (N_21036,N_20060,N_19886);
nand U21037 (N_21037,N_19930,N_20573);
nor U21038 (N_21038,N_20236,N_20514);
xor U21039 (N_21039,N_20089,N_20572);
xnor U21040 (N_21040,N_20558,N_20860);
xnor U21041 (N_21041,N_20969,N_20893);
nor U21042 (N_21042,N_20830,N_20964);
and U21043 (N_21043,N_20551,N_20764);
nor U21044 (N_21044,N_20899,N_20741);
and U21045 (N_21045,N_20008,N_20907);
nand U21046 (N_21046,N_20658,N_19845);
nor U21047 (N_21047,N_20308,N_20158);
xnor U21048 (N_21048,N_20117,N_20695);
and U21049 (N_21049,N_20460,N_20888);
or U21050 (N_21050,N_19978,N_20628);
nor U21051 (N_21051,N_19633,N_20780);
and U21052 (N_21052,N_20040,N_20756);
nor U21053 (N_21053,N_20090,N_20186);
and U21054 (N_21054,N_19686,N_19897);
xnor U21055 (N_21055,N_20585,N_19676);
nand U21056 (N_21056,N_19893,N_20344);
nor U21057 (N_21057,N_19626,N_20804);
nor U21058 (N_21058,N_20816,N_19890);
or U21059 (N_21059,N_20920,N_19899);
nand U21060 (N_21060,N_20970,N_20211);
nor U21061 (N_21061,N_19803,N_20337);
or U21062 (N_21062,N_20726,N_20277);
xnor U21063 (N_21063,N_20199,N_20148);
and U21064 (N_21064,N_20475,N_19589);
and U21065 (N_21065,N_20909,N_20535);
xor U21066 (N_21066,N_20336,N_20009);
or U21067 (N_21067,N_19699,N_19577);
and U21068 (N_21068,N_19985,N_20740);
nor U21069 (N_21069,N_19627,N_20256);
nand U21070 (N_21070,N_19567,N_19811);
or U21071 (N_21071,N_20796,N_20872);
and U21072 (N_21072,N_20889,N_19668);
nand U21073 (N_21073,N_20870,N_19745);
nor U21074 (N_21074,N_19613,N_20316);
nand U21075 (N_21075,N_19658,N_19720);
nand U21076 (N_21076,N_19840,N_19763);
or U21077 (N_21077,N_20698,N_19849);
nand U21078 (N_21078,N_20461,N_20732);
and U21079 (N_21079,N_20233,N_19989);
or U21080 (N_21080,N_20521,N_20007);
or U21081 (N_21081,N_20806,N_19859);
or U21082 (N_21082,N_20058,N_20976);
and U21083 (N_21083,N_20263,N_20023);
and U21084 (N_21084,N_19966,N_20714);
nand U21085 (N_21085,N_19857,N_20063);
and U21086 (N_21086,N_19856,N_20634);
xnor U21087 (N_21087,N_20073,N_20530);
nor U21088 (N_21088,N_20583,N_20003);
xor U21089 (N_21089,N_20010,N_20578);
and U21090 (N_21090,N_20002,N_19536);
and U21091 (N_21091,N_19621,N_19680);
nor U21092 (N_21092,N_19996,N_19674);
nor U21093 (N_21093,N_20605,N_19693);
or U21094 (N_21094,N_20654,N_20371);
xnor U21095 (N_21095,N_20280,N_20127);
nand U21096 (N_21096,N_19756,N_19500);
nor U21097 (N_21097,N_20749,N_19656);
nand U21098 (N_21098,N_19663,N_20581);
and U21099 (N_21099,N_19751,N_20987);
nand U21100 (N_21100,N_19504,N_20129);
nand U21101 (N_21101,N_20502,N_20052);
nor U21102 (N_21102,N_20998,N_20231);
or U21103 (N_21103,N_19692,N_19814);
or U21104 (N_21104,N_19952,N_20602);
nor U21105 (N_21105,N_20702,N_20232);
or U21106 (N_21106,N_20321,N_20792);
nor U21107 (N_21107,N_19622,N_20297);
nand U21108 (N_21108,N_20862,N_20850);
and U21109 (N_21109,N_20683,N_19644);
nor U21110 (N_21110,N_19765,N_20779);
nand U21111 (N_21111,N_19687,N_20712);
nor U21112 (N_21112,N_20497,N_20501);
or U21113 (N_21113,N_20482,N_19624);
and U21114 (N_21114,N_19993,N_20931);
nor U21115 (N_21115,N_20473,N_19837);
xor U21116 (N_21116,N_20390,N_20776);
or U21117 (N_21117,N_20278,N_20045);
nor U21118 (N_21118,N_19917,N_20294);
or U21119 (N_21119,N_20782,N_20917);
or U21120 (N_21120,N_20924,N_20286);
xnor U21121 (N_21121,N_20391,N_20189);
or U21122 (N_21122,N_20996,N_19880);
or U21123 (N_21123,N_20835,N_20464);
or U21124 (N_21124,N_20092,N_19939);
nand U21125 (N_21125,N_20921,N_20962);
or U21126 (N_21126,N_20638,N_20301);
and U21127 (N_21127,N_20119,N_20554);
nor U21128 (N_21128,N_20623,N_20584);
nand U21129 (N_21129,N_20662,N_20216);
and U21130 (N_21130,N_19772,N_20744);
or U21131 (N_21131,N_19652,N_20159);
xnor U21132 (N_21132,N_19706,N_20339);
xor U21133 (N_21133,N_20098,N_20494);
or U21134 (N_21134,N_20151,N_20840);
and U21135 (N_21135,N_20370,N_20704);
nand U21136 (N_21136,N_20386,N_19884);
and U21137 (N_21137,N_20095,N_20361);
nand U21138 (N_21138,N_19660,N_20257);
xor U21139 (N_21139,N_20863,N_20240);
nand U21140 (N_21140,N_20515,N_20382);
or U21141 (N_21141,N_20100,N_20427);
xnor U21142 (N_21142,N_20018,N_20847);
or U21143 (N_21143,N_20420,N_20462);
or U21144 (N_21144,N_19614,N_19933);
and U21145 (N_21145,N_19544,N_20680);
nand U21146 (N_21146,N_20647,N_20728);
nand U21147 (N_21147,N_20014,N_20925);
nor U21148 (N_21148,N_20739,N_20771);
and U21149 (N_21149,N_20984,N_20611);
or U21150 (N_21150,N_19640,N_20430);
nor U21151 (N_21151,N_19832,N_20725);
nand U21152 (N_21152,N_20088,N_20657);
nand U21153 (N_21153,N_20723,N_20318);
nor U21154 (N_21154,N_19846,N_20099);
xor U21155 (N_21155,N_20954,N_20833);
or U21156 (N_21156,N_19969,N_19848);
nand U21157 (N_21157,N_19861,N_19601);
nand U21158 (N_21158,N_19690,N_20503);
xnor U21159 (N_21159,N_20179,N_20980);
nor U21160 (N_21160,N_19860,N_20242);
nand U21161 (N_21161,N_20388,N_20223);
nand U21162 (N_21162,N_19740,N_19736);
nor U21163 (N_21163,N_19888,N_20633);
and U21164 (N_21164,N_19817,N_19908);
and U21165 (N_21165,N_19510,N_19649);
or U21166 (N_21166,N_20120,N_19501);
or U21167 (N_21167,N_19999,N_19545);
nor U21168 (N_21168,N_19773,N_19858);
or U21169 (N_21169,N_20262,N_20408);
and U21170 (N_21170,N_19598,N_19518);
nor U21171 (N_21171,N_20978,N_20315);
nor U21172 (N_21172,N_20195,N_20356);
nor U21173 (N_21173,N_20152,N_20691);
nor U21174 (N_21174,N_20220,N_20802);
nor U21175 (N_21175,N_20275,N_19546);
xnor U21176 (N_21176,N_19587,N_20822);
nor U21177 (N_21177,N_20400,N_19974);
and U21178 (N_21178,N_20857,N_20772);
or U21179 (N_21179,N_19920,N_19825);
or U21180 (N_21180,N_20729,N_19870);
or U21181 (N_21181,N_20171,N_20251);
nand U21182 (N_21182,N_20273,N_20184);
nor U21183 (N_21183,N_20259,N_19551);
or U21184 (N_21184,N_20373,N_20660);
and U21185 (N_21185,N_20387,N_19572);
and U21186 (N_21186,N_20507,N_19724);
xor U21187 (N_21187,N_20834,N_19790);
nand U21188 (N_21188,N_20168,N_20364);
nand U21189 (N_21189,N_19843,N_19921);
and U21190 (N_21190,N_19946,N_20130);
or U21191 (N_21191,N_20136,N_20908);
nand U21192 (N_21192,N_20209,N_20167);
and U21193 (N_21193,N_20661,N_20604);
nor U21194 (N_21194,N_19863,N_20035);
xor U21195 (N_21195,N_20950,N_19678);
and U21196 (N_21196,N_20989,N_20856);
or U21197 (N_21197,N_20773,N_19512);
or U21198 (N_21198,N_20360,N_19723);
and U21199 (N_21199,N_19617,N_19516);
nand U21200 (N_21200,N_20428,N_20309);
and U21201 (N_21201,N_20006,N_20225);
nor U21202 (N_21202,N_20879,N_20593);
or U21203 (N_21203,N_19535,N_19753);
and U21204 (N_21204,N_19620,N_20653);
xor U21205 (N_21205,N_19557,N_19569);
or U21206 (N_21206,N_19798,N_20610);
and U21207 (N_21207,N_20936,N_20380);
xor U21208 (N_21208,N_20330,N_20667);
or U21209 (N_21209,N_20374,N_19647);
xnor U21210 (N_21210,N_20334,N_20625);
and U21211 (N_21211,N_20971,N_20228);
and U21212 (N_21212,N_19882,N_20639);
nor U21213 (N_21213,N_20432,N_20208);
nand U21214 (N_21214,N_19851,N_19766);
nand U21215 (N_21215,N_19657,N_19833);
xnor U21216 (N_21216,N_19730,N_20902);
nand U21217 (N_21217,N_20550,N_20973);
nor U21218 (N_21218,N_20803,N_20271);
nand U21219 (N_21219,N_19963,N_19788);
xor U21220 (N_21220,N_20883,N_20307);
nor U21221 (N_21221,N_20044,N_20706);
and U21222 (N_21222,N_20753,N_20272);
nand U21223 (N_21223,N_19761,N_20734);
or U21224 (N_21224,N_20283,N_20914);
or U21225 (N_21225,N_20440,N_20291);
and U21226 (N_21226,N_20226,N_20659);
xor U21227 (N_21227,N_19961,N_20722);
or U21228 (N_21228,N_19783,N_20733);
nand U21229 (N_21229,N_20429,N_20247);
xnor U21230 (N_21230,N_20718,N_20131);
and U21231 (N_21231,N_19883,N_20929);
nand U21232 (N_21232,N_20594,N_20468);
or U21233 (N_21233,N_19926,N_20520);
nand U21234 (N_21234,N_19717,N_20851);
and U21235 (N_21235,N_20397,N_19808);
xor U21236 (N_21236,N_20222,N_19970);
and U21237 (N_21237,N_20416,N_19741);
and U21238 (N_21238,N_20531,N_20664);
and U21239 (N_21239,N_20101,N_20650);
nand U21240 (N_21240,N_20080,N_20527);
xnor U21241 (N_21241,N_20717,N_20784);
xnor U21242 (N_21242,N_20956,N_20932);
nor U21243 (N_21243,N_20113,N_20068);
nand U21244 (N_21244,N_19664,N_20446);
or U21245 (N_21245,N_20993,N_19611);
xnor U21246 (N_21246,N_20624,N_20495);
nand U21247 (N_21247,N_19584,N_20635);
nor U21248 (N_21248,N_20453,N_20812);
xor U21249 (N_21249,N_20543,N_20295);
nand U21250 (N_21250,N_19731,N_20640);
or U21251 (N_21251,N_20616,N_20681);
xnor U21252 (N_21252,N_20557,N_20174);
and U21253 (N_21253,N_20322,N_20104);
xor U21254 (N_21254,N_20891,N_20778);
nor U21255 (N_21255,N_20498,N_19697);
nor U21256 (N_21256,N_19553,N_20671);
or U21257 (N_21257,N_20431,N_20959);
xnor U21258 (N_21258,N_19956,N_20150);
nor U21259 (N_21259,N_20326,N_19734);
and U21260 (N_21260,N_20467,N_19575);
xnor U21261 (N_21261,N_19715,N_19945);
xor U21262 (N_21262,N_20791,N_20481);
xnor U21263 (N_21263,N_20258,N_20083);
or U21264 (N_21264,N_20470,N_19839);
nor U21265 (N_21265,N_20156,N_20892);
or U21266 (N_21266,N_20579,N_19733);
nand U21267 (N_21267,N_20775,N_19876);
or U21268 (N_21268,N_19526,N_19718);
nor U21269 (N_21269,N_20145,N_20051);
nor U21270 (N_21270,N_19954,N_20114);
nor U21271 (N_21271,N_20486,N_19830);
or U21272 (N_21272,N_20676,N_20670);
xor U21273 (N_21273,N_19562,N_19877);
nor U21274 (N_21274,N_20532,N_20548);
and U21275 (N_21275,N_20059,N_20622);
and U21276 (N_21276,N_19659,N_20823);
nand U21277 (N_21277,N_20672,N_20210);
or U21278 (N_21278,N_20565,N_20140);
or U21279 (N_21279,N_20124,N_20958);
nand U21280 (N_21280,N_19594,N_20582);
nor U21281 (N_21281,N_20968,N_20177);
or U21282 (N_21282,N_19965,N_20617);
and U21283 (N_21283,N_20036,N_19612);
nand U21284 (N_21284,N_19714,N_20549);
nand U21285 (N_21285,N_20474,N_20895);
xnor U21286 (N_21286,N_20811,N_19514);
or U21287 (N_21287,N_19635,N_20944);
or U21288 (N_21288,N_20600,N_20965);
nand U21289 (N_21289,N_20214,N_20673);
xnor U21290 (N_21290,N_20320,N_20724);
nand U21291 (N_21291,N_19902,N_20566);
nor U21292 (N_21292,N_20831,N_20577);
nor U21293 (N_21293,N_19552,N_19958);
nand U21294 (N_21294,N_20927,N_20886);
or U21295 (N_21295,N_20071,N_20707);
nor U21296 (N_21296,N_20445,N_20346);
nand U21297 (N_21297,N_20939,N_20032);
xnor U21298 (N_21298,N_20146,N_20807);
nor U21299 (N_21299,N_20013,N_20646);
nor U21300 (N_21300,N_20916,N_19579);
xnor U21301 (N_21301,N_20518,N_19520);
nor U21302 (N_21302,N_20064,N_20564);
and U21303 (N_21303,N_19695,N_19755);
and U21304 (N_21304,N_20196,N_20894);
and U21305 (N_21305,N_19770,N_20637);
nand U21306 (N_21306,N_20621,N_20533);
nor U21307 (N_21307,N_19596,N_19637);
nand U21308 (N_21308,N_19515,N_20172);
xnor U21309 (N_21309,N_20645,N_20742);
nor U21310 (N_21310,N_20900,N_20552);
nor U21311 (N_21311,N_20999,N_20553);
nand U21312 (N_21312,N_19521,N_19655);
or U21313 (N_21313,N_20601,N_20687);
nand U21314 (N_21314,N_20028,N_19834);
and U21315 (N_21315,N_20163,N_20853);
nand U21316 (N_21316,N_20595,N_20841);
nor U21317 (N_21317,N_20340,N_19636);
nor U21318 (N_21318,N_20981,N_19600);
nor U21319 (N_21319,N_20937,N_20805);
nor U21320 (N_21320,N_20252,N_20930);
xor U21321 (N_21321,N_19738,N_19847);
nor U21322 (N_21322,N_19809,N_19605);
or U21323 (N_21323,N_20402,N_19804);
or U21324 (N_21324,N_19698,N_20281);
or U21325 (N_21325,N_20757,N_20133);
nor U21326 (N_21326,N_19855,N_20298);
nor U21327 (N_21327,N_20668,N_20864);
and U21328 (N_21328,N_20097,N_20338);
nand U21329 (N_21329,N_19691,N_20614);
or U21330 (N_21330,N_19654,N_19782);
xnor U21331 (N_21331,N_19991,N_20953);
and U21332 (N_21332,N_19704,N_20810);
or U21333 (N_21333,N_20696,N_20323);
nand U21334 (N_21334,N_19580,N_20798);
nor U21335 (N_21335,N_20938,N_19533);
xnor U21336 (N_21336,N_20919,N_19885);
and U21337 (N_21337,N_20801,N_20434);
xor U21338 (N_21338,N_20479,N_20818);
or U21339 (N_21339,N_19819,N_19904);
and U21340 (N_21340,N_20710,N_20546);
xor U21341 (N_21341,N_19524,N_19650);
and U21342 (N_21342,N_20328,N_20077);
nor U21343 (N_21343,N_20354,N_20471);
xnor U21344 (N_21344,N_20505,N_19599);
xnor U21345 (N_21345,N_19774,N_20123);
or U21346 (N_21346,N_20444,N_20441);
xor U21347 (N_21347,N_20162,N_20730);
and U21348 (N_21348,N_19540,N_19685);
nand U21349 (N_21349,N_20022,N_19962);
or U21350 (N_21350,N_20990,N_20651);
nor U21351 (N_21351,N_19648,N_20203);
xnor U21352 (N_21352,N_20963,N_20116);
and U21353 (N_21353,N_20246,N_19866);
nand U21354 (N_21354,N_20487,N_20385);
nand U21355 (N_21355,N_20824,N_19768);
nand U21356 (N_21356,N_20284,N_20966);
or U21357 (N_21357,N_20607,N_20488);
nand U21358 (N_21358,N_20761,N_19905);
or U21359 (N_21359,N_20362,N_19869);
nor U21360 (N_21360,N_20945,N_19955);
nand U21361 (N_21361,N_20849,N_20149);
or U21362 (N_21362,N_20537,N_20492);
xnor U21363 (N_21363,N_20456,N_19752);
or U21364 (N_21364,N_19871,N_19581);
and U21365 (N_21365,N_20684,N_19909);
xnor U21366 (N_21366,N_20015,N_20312);
nor U21367 (N_21367,N_20218,N_20682);
or U21368 (N_21368,N_20173,N_20241);
nand U21369 (N_21369,N_20031,N_20046);
nor U21370 (N_21370,N_20519,N_19632);
nand U21371 (N_21371,N_20613,N_19988);
and U21372 (N_21372,N_20306,N_20826);
nand U21373 (N_21373,N_20763,N_20411);
xnor U21374 (N_21374,N_20419,N_20869);
nand U21375 (N_21375,N_20922,N_20866);
nor U21376 (N_21376,N_19646,N_20844);
or U21377 (N_21377,N_20598,N_20108);
nor U21378 (N_21378,N_20800,N_19610);
xnor U21379 (N_21379,N_19992,N_20738);
xor U21380 (N_21380,N_20215,N_19940);
or U21381 (N_21381,N_19754,N_20540);
or U21382 (N_21382,N_20923,N_20181);
xor U21383 (N_21383,N_20941,N_20086);
and U21384 (N_21384,N_20731,N_19604);
nand U21385 (N_21385,N_19776,N_20255);
nor U21386 (N_21386,N_20265,N_20112);
nand U21387 (N_21387,N_19616,N_19711);
nand U21388 (N_21388,N_20694,N_19997);
xnor U21389 (N_21389,N_20260,N_20974);
nor U21390 (N_21390,N_19750,N_20235);
xnor U21391 (N_21391,N_20597,N_19998);
xor U21392 (N_21392,N_20274,N_20055);
nor U21393 (N_21393,N_20125,N_20703);
nand U21394 (N_21394,N_20053,N_20642);
nand U21395 (N_21395,N_20106,N_20913);
xor U21396 (N_21396,N_19912,N_20439);
nand U21397 (N_21397,N_20885,N_19573);
nor U21398 (N_21398,N_20062,N_20443);
or U21399 (N_21399,N_20379,N_20327);
or U21400 (N_21400,N_20911,N_20160);
xnor U21401 (N_21401,N_20606,N_20788);
nor U21402 (N_21402,N_19625,N_19710);
and U21403 (N_21403,N_19527,N_19931);
or U21404 (N_21404,N_19919,N_20845);
nand U21405 (N_21405,N_19769,N_20524);
or U21406 (N_21406,N_20643,N_19602);
and U21407 (N_21407,N_20454,N_19628);
and U21408 (N_21408,N_20227,N_19722);
nand U21409 (N_21409,N_19972,N_19791);
nor U21410 (N_21410,N_19749,N_20042);
xor U21411 (N_21411,N_20905,N_19957);
nor U21412 (N_21412,N_20375,N_20912);
xor U21413 (N_21413,N_19746,N_19976);
nor U21414 (N_21414,N_19671,N_19786);
and U21415 (N_21415,N_20865,N_20061);
xnor U21416 (N_21416,N_20943,N_20868);
nor U21417 (N_21417,N_20525,N_20302);
or U21418 (N_21418,N_19918,N_19574);
xnor U21419 (N_21419,N_20777,N_19634);
and U21420 (N_21420,N_19682,N_20770);
or U21421 (N_21421,N_19894,N_20447);
or U21422 (N_21422,N_19683,N_20632);
xor U21423 (N_21423,N_19973,N_19779);
xor U21424 (N_21424,N_20854,N_20529);
or U21425 (N_21425,N_20508,N_20352);
nor U21426 (N_21426,N_19618,N_20522);
or U21427 (N_21427,N_20588,N_20794);
nor U21428 (N_21428,N_20652,N_20693);
nor U21429 (N_21429,N_19505,N_20314);
nor U21430 (N_21430,N_19807,N_19642);
nand U21431 (N_21431,N_20193,N_19906);
and U21432 (N_21432,N_20880,N_20313);
nand U21433 (N_21433,N_20463,N_19502);
nand U21434 (N_21434,N_19593,N_20290);
xnor U21435 (N_21435,N_20679,N_19537);
nor U21436 (N_21436,N_20663,N_19949);
nor U21437 (N_21437,N_19844,N_20017);
nor U21438 (N_21438,N_20523,N_20020);
xor U21439 (N_21439,N_19875,N_19950);
and U21440 (N_21440,N_19677,N_20157);
or U21441 (N_21441,N_20197,N_20630);
nand U21442 (N_21442,N_20369,N_20781);
nor U21443 (N_21443,N_20365,N_19948);
nor U21444 (N_21444,N_20254,N_20576);
nor U21445 (N_21445,N_20620,N_20264);
nor U21446 (N_21446,N_19670,N_20627);
nand U21447 (N_21447,N_20813,N_20037);
and U21448 (N_21448,N_19548,N_19576);
xnor U21449 (N_21449,N_19603,N_20192);
and U21450 (N_21450,N_20421,N_20904);
xnor U21451 (N_21451,N_19538,N_19583);
nor U21452 (N_21452,N_20825,N_19821);
nand U21453 (N_21453,N_20001,N_20947);
or U21454 (N_21454,N_19653,N_20412);
xnor U21455 (N_21455,N_19619,N_19941);
nor U21456 (N_21456,N_19984,N_20355);
and U21457 (N_21457,N_19513,N_19523);
xor U21458 (N_21458,N_20389,N_20452);
nand U21459 (N_21459,N_19667,N_20649);
or U21460 (N_21460,N_20279,N_20985);
nor U21461 (N_21461,N_20085,N_20268);
or U21462 (N_21462,N_20674,N_19823);
nand U21463 (N_21463,N_20949,N_19585);
or U21464 (N_21464,N_20992,N_20569);
nor U21465 (N_21465,N_20450,N_20363);
xor U21466 (N_21466,N_19560,N_19712);
nand U21467 (N_21467,N_19534,N_20875);
nor U21468 (N_21468,N_20720,N_19757);
or U21469 (N_21469,N_20539,N_20066);
nand U21470 (N_21470,N_20213,N_20054);
and U21471 (N_21471,N_20752,N_20560);
nor U21472 (N_21472,N_20815,N_20433);
or U21473 (N_21473,N_20079,N_20513);
xor U21474 (N_21474,N_20995,N_20392);
xor U21475 (N_21475,N_19937,N_20983);
nor U21476 (N_21476,N_20747,N_19868);
nor U21477 (N_21477,N_20828,N_20843);
nor U21478 (N_21478,N_20542,N_20951);
nor U21479 (N_21479,N_20041,N_20768);
and U21480 (N_21480,N_19824,N_20201);
and U21481 (N_21481,N_20897,N_20563);
nor U21482 (N_21482,N_20896,N_20169);
xor U21483 (N_21483,N_20409,N_20425);
and U21484 (N_21484,N_20183,N_19630);
xnor U21485 (N_21485,N_20033,N_19519);
xnor U21486 (N_21486,N_20977,N_20500);
nor U21487 (N_21487,N_20918,N_19935);
nand U21488 (N_21488,N_20785,N_20143);
or U21489 (N_21489,N_20310,N_20952);
and U21490 (N_21490,N_20884,N_20395);
nand U21491 (N_21491,N_19828,N_19922);
nand U21492 (N_21492,N_20383,N_20288);
xnor U21493 (N_21493,N_20372,N_19570);
xnor U21494 (N_21494,N_20333,N_20121);
nor U21495 (N_21495,N_19827,N_20799);
xnor U21496 (N_21496,N_20175,N_20699);
xnor U21497 (N_21497,N_19967,N_20517);
nor U21498 (N_21498,N_19608,N_20767);
or U21499 (N_21499,N_20138,N_19758);
nand U21500 (N_21500,N_20555,N_20110);
xor U21501 (N_21501,N_20819,N_20790);
nand U21502 (N_21502,N_20876,N_19506);
xnor U21503 (N_21503,N_20396,N_20592);
nand U21504 (N_21504,N_20586,N_19525);
nor U21505 (N_21505,N_19800,N_20836);
xor U21506 (N_21506,N_20493,N_19864);
or U21507 (N_21507,N_20155,N_20568);
xnor U21508 (N_21508,N_20636,N_20615);
xnor U21509 (N_21509,N_19554,N_20655);
and U21510 (N_21510,N_19841,N_20538);
or U21511 (N_21511,N_20378,N_20736);
nor U21512 (N_21512,N_20751,N_20997);
and U21513 (N_21513,N_20901,N_20451);
or U21514 (N_21514,N_19805,N_19896);
and U21515 (N_21515,N_20504,N_19977);
xor U21516 (N_21516,N_20934,N_20437);
nor U21517 (N_21517,N_19826,N_19914);
xor U21518 (N_21518,N_20859,N_20224);
nor U21519 (N_21519,N_19987,N_19891);
and U21520 (N_21520,N_20890,N_20282);
and U21521 (N_21521,N_20349,N_20300);
or U21522 (N_21522,N_19689,N_20737);
nor U21523 (N_21523,N_20176,N_20329);
xor U21524 (N_21524,N_20935,N_19831);
nand U21525 (N_21525,N_19522,N_19592);
xnor U21526 (N_21526,N_20528,N_19901);
and U21527 (N_21527,N_20967,N_20590);
or U21528 (N_21528,N_20027,N_20940);
and U21529 (N_21529,N_20393,N_19511);
nand U21530 (N_21530,N_19822,N_20137);
nor U21531 (N_21531,N_20982,N_20377);
or U21532 (N_21532,N_20526,N_19565);
nor U21533 (N_21533,N_19539,N_20765);
nand U21534 (N_21534,N_19684,N_20331);
xor U21535 (N_21535,N_20212,N_19760);
xnor U21536 (N_21536,N_20612,N_20404);
and U21537 (N_21537,N_19923,N_20484);
or U21538 (N_21538,N_19615,N_19701);
xnor U21539 (N_21539,N_19852,N_20047);
xor U21540 (N_21540,N_20458,N_20219);
or U21541 (N_21541,N_19541,N_20004);
xor U21542 (N_21542,N_19507,N_19555);
and U21543 (N_21543,N_20496,N_20229);
nand U21544 (N_21544,N_20690,N_20038);
and U21545 (N_21545,N_20787,N_20510);
nand U21546 (N_21546,N_20858,N_19645);
nor U21547 (N_21547,N_19892,N_20039);
nor U21548 (N_21548,N_19737,N_20205);
or U21549 (N_21549,N_20903,N_19732);
or U21550 (N_21550,N_19938,N_19595);
nand U21551 (N_21551,N_20069,N_20118);
and U21552 (N_21552,N_20332,N_20979);
and U21553 (N_21553,N_20289,N_20618);
nand U21554 (N_21554,N_20745,N_20477);
nor U21555 (N_21555,N_19597,N_19784);
xor U21556 (N_21556,N_19629,N_19542);
nor U21557 (N_21557,N_20103,N_20030);
nor U21558 (N_21558,N_20499,N_19729);
and U21559 (N_21559,N_20422,N_20351);
nand U21560 (N_21560,N_20561,N_20541);
nand U21561 (N_21561,N_19586,N_20081);
and U21562 (N_21562,N_19797,N_19547);
nor U21563 (N_21563,N_20345,N_20547);
nor U21564 (N_21564,N_19986,N_20906);
nor U21565 (N_21565,N_19675,N_20403);
nand U21566 (N_21566,N_20384,N_19762);
or U21567 (N_21567,N_20248,N_20435);
nand U21568 (N_21568,N_20669,N_19990);
xnor U21569 (N_21569,N_20424,N_20933);
or U21570 (N_21570,N_20719,N_19995);
nor U21571 (N_21571,N_19606,N_20536);
or U21572 (N_21572,N_20410,N_20469);
or U21573 (N_21573,N_19764,N_19802);
or U21574 (N_21574,N_19878,N_19850);
xor U21575 (N_21575,N_20887,N_19568);
nand U21576 (N_21576,N_20820,N_20407);
nand U21577 (N_21577,N_20848,N_19679);
nor U21578 (N_21578,N_20078,N_20024);
xor U21579 (N_21579,N_20754,N_20026);
nor U21580 (N_21580,N_20760,N_19887);
nand U21581 (N_21581,N_19688,N_20303);
nand U21582 (N_21582,N_20185,N_19705);
and U21583 (N_21583,N_20012,N_20867);
nor U21584 (N_21584,N_20141,N_20111);
nor U21585 (N_21585,N_19727,N_20727);
nand U21586 (N_21586,N_19721,N_20678);
xnor U21587 (N_21587,N_19796,N_19873);
nand U21588 (N_21588,N_20821,N_19775);
or U21589 (N_21589,N_19910,N_20417);
xnor U21590 (N_21590,N_19550,N_20490);
xor U21591 (N_21591,N_20898,N_19781);
nor U21592 (N_21592,N_20877,N_19942);
nand U21593 (N_21593,N_20243,N_19672);
and U21594 (N_21594,N_19651,N_20988);
nand U21595 (N_21595,N_20459,N_20603);
or U21596 (N_21596,N_20544,N_20418);
nand U21597 (N_21597,N_19528,N_20472);
nand U21598 (N_21598,N_20599,N_20688);
and U21599 (N_21599,N_20204,N_19578);
nor U21600 (N_21600,N_20182,N_20511);
nor U21601 (N_21601,N_20244,N_20381);
and U21602 (N_21602,N_20715,N_19867);
nand U21603 (N_21603,N_20082,N_20198);
or U21604 (N_21604,N_20735,N_19744);
xnor U21605 (N_21605,N_19747,N_19964);
xnor U21606 (N_21606,N_19571,N_20135);
nor U21607 (N_21607,N_20873,N_20115);
nand U21608 (N_21608,N_19959,N_20759);
nand U21609 (N_21609,N_19716,N_20449);
nor U21610 (N_21610,N_20716,N_20253);
nor U21611 (N_21611,N_19865,N_20132);
nand U21612 (N_21612,N_20852,N_19588);
and U21613 (N_21613,N_19854,N_20194);
and U21614 (N_21614,N_19936,N_19872);
or U21615 (N_21615,N_20034,N_20405);
and U21616 (N_21616,N_19556,N_20881);
nor U21617 (N_21617,N_20855,N_20489);
and U21618 (N_21618,N_19907,N_19662);
nand U21619 (N_21619,N_20292,N_20335);
nor U21620 (N_21620,N_20644,N_20122);
and U21621 (N_21621,N_20942,N_20448);
nor U21622 (N_21622,N_20697,N_19795);
and U21623 (N_21623,N_20758,N_20139);
nor U21624 (N_21624,N_20019,N_20348);
xor U21625 (N_21625,N_20991,N_20955);
or U21626 (N_21626,N_20070,N_20102);
and U21627 (N_21627,N_20075,N_19980);
nor U21628 (N_21628,N_20341,N_20144);
xor U21629 (N_21629,N_19929,N_20829);
nand U21630 (N_21630,N_20928,N_19767);
nand U21631 (N_21631,N_20648,N_20107);
xnor U21632 (N_21632,N_20269,N_20000);
or U21633 (N_21633,N_19759,N_20234);
xnor U21634 (N_21634,N_19566,N_20368);
nor U21635 (N_21635,N_19639,N_19934);
nand U21636 (N_21636,N_19543,N_20180);
xnor U21637 (N_21637,N_20016,N_20721);
nand U21638 (N_21638,N_20304,N_19503);
nand U21639 (N_21639,N_20414,N_19713);
and U21640 (N_21640,N_19927,N_20296);
and U21641 (N_21641,N_19669,N_20631);
nand U21642 (N_21642,N_20986,N_20317);
nand U21643 (N_21643,N_20783,N_19743);
nand U21644 (N_21644,N_20915,N_20043);
and U21645 (N_21645,N_20685,N_20359);
xnor U21646 (N_21646,N_20609,N_20666);
nand U21647 (N_21647,N_20701,N_19903);
xor U21648 (N_21648,N_20677,N_20839);
or U21649 (N_21649,N_20574,N_20641);
nand U21650 (N_21650,N_19799,N_20164);
nand U21651 (N_21651,N_20206,N_19785);
nand U21652 (N_21652,N_20882,N_20705);
or U21653 (N_21653,N_20589,N_20406);
and U21654 (N_21654,N_19793,N_19787);
or U21655 (N_21655,N_20153,N_20238);
xnor U21656 (N_21656,N_19661,N_20793);
and U21657 (N_21657,N_20562,N_20711);
and U21658 (N_21658,N_20342,N_20050);
or U21659 (N_21659,N_20516,N_20343);
nand U21660 (N_21660,N_19981,N_19874);
and U21661 (N_21661,N_19806,N_20072);
or U21662 (N_21662,N_20237,N_20591);
nand U21663 (N_21663,N_19925,N_20311);
nor U21664 (N_21664,N_20960,N_20485);
xor U21665 (N_21665,N_19563,N_20994);
and U21666 (N_21666,N_20656,N_20350);
nand U21667 (N_21667,N_20399,N_20325);
and U21668 (N_21668,N_19835,N_20455);
nor U21669 (N_21669,N_20076,N_20957);
xnor U21670 (N_21670,N_20814,N_20692);
nor U21671 (N_21671,N_19810,N_20084);
nand U21672 (N_21672,N_19898,N_19709);
or U21673 (N_21673,N_20230,N_19582);
or U21674 (N_21674,N_19607,N_19944);
and U21675 (N_21675,N_19561,N_20972);
and U21676 (N_21676,N_20846,N_19879);
or U21677 (N_21677,N_20874,N_19836);
and U21678 (N_21678,N_20556,N_19792);
nand U21679 (N_21679,N_20267,N_20774);
or U21680 (N_21680,N_19794,N_19953);
xnor U21681 (N_21681,N_20567,N_20105);
or U21682 (N_21682,N_20808,N_20413);
xnor U21683 (N_21683,N_20750,N_20287);
nor U21684 (N_21684,N_19820,N_19932);
nor U21685 (N_21685,N_20457,N_20786);
or U21686 (N_21686,N_19928,N_19700);
nand U21687 (N_21687,N_20948,N_20837);
xnor U21688 (N_21688,N_20109,N_20005);
or U21689 (N_21689,N_20619,N_20946);
xor U21690 (N_21690,N_19703,N_19778);
nand U21691 (N_21691,N_20029,N_20065);
or U21692 (N_21692,N_20165,N_19631);
nor U21693 (N_21693,N_20202,N_19719);
xnor U21694 (N_21694,N_20975,N_20827);
nand U21695 (N_21695,N_20357,N_19913);
xor U21696 (N_21696,N_20491,N_20878);
nor U21697 (N_21697,N_20512,N_20401);
nor U21698 (N_21698,N_20708,N_20832);
or U21699 (N_21699,N_20170,N_20587);
xor U21700 (N_21700,N_20797,N_20675);
nand U21701 (N_21701,N_19530,N_19911);
nand U21702 (N_21702,N_20249,N_19748);
nor U21703 (N_21703,N_20713,N_19816);
nand U21704 (N_21704,N_20665,N_20466);
or U21705 (N_21705,N_20049,N_20608);
and U21706 (N_21706,N_20571,N_19777);
and U21707 (N_21707,N_20239,N_19728);
xor U21708 (N_21708,N_20769,N_20817);
nor U21709 (N_21709,N_19696,N_20709);
or U21710 (N_21710,N_20755,N_19771);
and U21711 (N_21711,N_19975,N_20091);
xnor U21712 (N_21712,N_20746,N_20838);
or U21713 (N_21713,N_20442,N_20861);
and U21714 (N_21714,N_19694,N_20187);
nand U21715 (N_21715,N_19609,N_19889);
xor U21716 (N_21716,N_20570,N_19591);
nor U21717 (N_21717,N_20394,N_20285);
xnor U21718 (N_21718,N_20191,N_20067);
nand U21719 (N_21719,N_20871,N_19815);
xnor U21720 (N_21720,N_20142,N_19881);
nand U21721 (N_21721,N_20376,N_20580);
nand U21722 (N_21722,N_20423,N_19708);
nand U21723 (N_21723,N_19801,N_20961);
and U21724 (N_21724,N_20154,N_20506);
nand U21725 (N_21725,N_20057,N_19742);
and U21726 (N_21726,N_20200,N_19707);
and U21727 (N_21727,N_20221,N_20438);
and U21728 (N_21728,N_19509,N_19726);
and U21729 (N_21729,N_20686,N_20299);
and U21730 (N_21730,N_20700,N_20910);
nand U21731 (N_21731,N_20207,N_20545);
nand U21732 (N_21732,N_19681,N_20025);
and U21733 (N_21733,N_19725,N_20147);
xnor U21734 (N_21734,N_20178,N_20626);
nand U21735 (N_21735,N_19517,N_20415);
and U21736 (N_21736,N_20480,N_20398);
xnor U21737 (N_21737,N_19666,N_20293);
or U21738 (N_21738,N_19643,N_19549);
nor U21739 (N_21739,N_20926,N_19924);
or U21740 (N_21740,N_20305,N_20509);
xor U21741 (N_21741,N_20436,N_19558);
or U21742 (N_21742,N_20048,N_19994);
nor U21743 (N_21743,N_19979,N_19780);
and U21744 (N_21744,N_20795,N_19842);
and U21745 (N_21745,N_19853,N_20087);
nand U21746 (N_21746,N_20366,N_20596);
or U21747 (N_21747,N_20190,N_20319);
nor U21748 (N_21748,N_19943,N_19982);
nand U21749 (N_21749,N_20021,N_20056);
and U21750 (N_21750,N_20595,N_20035);
nand U21751 (N_21751,N_19976,N_20466);
and U21752 (N_21752,N_20988,N_20719);
or U21753 (N_21753,N_19993,N_20664);
nor U21754 (N_21754,N_19930,N_20194);
nand U21755 (N_21755,N_19785,N_20268);
nor U21756 (N_21756,N_20729,N_19575);
nor U21757 (N_21757,N_20783,N_20099);
nor U21758 (N_21758,N_20163,N_19932);
nor U21759 (N_21759,N_20099,N_20646);
xor U21760 (N_21760,N_20661,N_20299);
xnor U21761 (N_21761,N_20159,N_20240);
and U21762 (N_21762,N_20643,N_19539);
nand U21763 (N_21763,N_20091,N_20621);
nor U21764 (N_21764,N_19669,N_19931);
and U21765 (N_21765,N_20863,N_20914);
nor U21766 (N_21766,N_19776,N_19868);
xnor U21767 (N_21767,N_20496,N_19647);
nor U21768 (N_21768,N_20120,N_20121);
or U21769 (N_21769,N_20049,N_20098);
nor U21770 (N_21770,N_19671,N_19607);
xnor U21771 (N_21771,N_19886,N_20012);
nand U21772 (N_21772,N_20924,N_20616);
and U21773 (N_21773,N_20529,N_19631);
or U21774 (N_21774,N_20099,N_20625);
and U21775 (N_21775,N_20270,N_19728);
and U21776 (N_21776,N_20144,N_20730);
xnor U21777 (N_21777,N_19827,N_19821);
nand U21778 (N_21778,N_20629,N_20362);
or U21779 (N_21779,N_19873,N_19509);
xnor U21780 (N_21780,N_20078,N_20541);
and U21781 (N_21781,N_20518,N_19914);
xor U21782 (N_21782,N_20489,N_20809);
nand U21783 (N_21783,N_20937,N_20885);
xnor U21784 (N_21784,N_20836,N_20448);
or U21785 (N_21785,N_19546,N_20130);
nor U21786 (N_21786,N_20755,N_19760);
xnor U21787 (N_21787,N_20584,N_20471);
and U21788 (N_21788,N_19728,N_20667);
or U21789 (N_21789,N_19857,N_20803);
nor U21790 (N_21790,N_19898,N_20370);
or U21791 (N_21791,N_20046,N_19833);
xor U21792 (N_21792,N_19766,N_20891);
and U21793 (N_21793,N_19533,N_20262);
xnor U21794 (N_21794,N_19681,N_19804);
xnor U21795 (N_21795,N_20779,N_20903);
and U21796 (N_21796,N_20179,N_20118);
or U21797 (N_21797,N_20288,N_20547);
or U21798 (N_21798,N_20024,N_20085);
and U21799 (N_21799,N_19691,N_20335);
nor U21800 (N_21800,N_20512,N_20551);
xor U21801 (N_21801,N_20729,N_20932);
xor U21802 (N_21802,N_19669,N_19544);
and U21803 (N_21803,N_19638,N_19783);
nor U21804 (N_21804,N_20448,N_20861);
xnor U21805 (N_21805,N_20439,N_20507);
nor U21806 (N_21806,N_19667,N_19804);
or U21807 (N_21807,N_20907,N_20824);
nand U21808 (N_21808,N_20725,N_19882);
or U21809 (N_21809,N_20241,N_19975);
or U21810 (N_21810,N_19767,N_20212);
and U21811 (N_21811,N_20463,N_20407);
and U21812 (N_21812,N_20410,N_20662);
or U21813 (N_21813,N_19970,N_20014);
or U21814 (N_21814,N_20382,N_19744);
and U21815 (N_21815,N_20528,N_20294);
and U21816 (N_21816,N_19992,N_20146);
nand U21817 (N_21817,N_20456,N_20580);
or U21818 (N_21818,N_20008,N_19988);
and U21819 (N_21819,N_20813,N_20392);
nor U21820 (N_21820,N_19696,N_20679);
and U21821 (N_21821,N_20960,N_19741);
nor U21822 (N_21822,N_20770,N_20726);
and U21823 (N_21823,N_20067,N_19969);
xor U21824 (N_21824,N_20508,N_20251);
nor U21825 (N_21825,N_20049,N_20183);
nand U21826 (N_21826,N_19504,N_19695);
xnor U21827 (N_21827,N_19654,N_19714);
nor U21828 (N_21828,N_19810,N_20045);
xnor U21829 (N_21829,N_20249,N_20510);
or U21830 (N_21830,N_20549,N_20696);
nand U21831 (N_21831,N_20604,N_19953);
nand U21832 (N_21832,N_20601,N_20075);
nor U21833 (N_21833,N_20193,N_20362);
nor U21834 (N_21834,N_20377,N_20461);
nand U21835 (N_21835,N_20233,N_20966);
xor U21836 (N_21836,N_20385,N_20978);
nor U21837 (N_21837,N_19921,N_20392);
and U21838 (N_21838,N_19734,N_19532);
and U21839 (N_21839,N_19753,N_20160);
xor U21840 (N_21840,N_20183,N_19913);
or U21841 (N_21841,N_19856,N_19881);
and U21842 (N_21842,N_20565,N_20612);
nand U21843 (N_21843,N_20858,N_20910);
nand U21844 (N_21844,N_20300,N_20289);
nor U21845 (N_21845,N_20176,N_20294);
nand U21846 (N_21846,N_20090,N_19999);
nor U21847 (N_21847,N_19532,N_20663);
xor U21848 (N_21848,N_20360,N_20378);
or U21849 (N_21849,N_20475,N_20710);
and U21850 (N_21850,N_20994,N_19896);
and U21851 (N_21851,N_20994,N_19757);
or U21852 (N_21852,N_20271,N_20119);
nor U21853 (N_21853,N_19820,N_19524);
and U21854 (N_21854,N_20812,N_20573);
nor U21855 (N_21855,N_19957,N_20551);
xnor U21856 (N_21856,N_20926,N_20023);
nor U21857 (N_21857,N_20146,N_20976);
nor U21858 (N_21858,N_20321,N_19864);
xnor U21859 (N_21859,N_20789,N_20692);
and U21860 (N_21860,N_20181,N_19524);
nand U21861 (N_21861,N_20431,N_20414);
nand U21862 (N_21862,N_20172,N_20876);
nor U21863 (N_21863,N_20961,N_20174);
or U21864 (N_21864,N_20694,N_20655);
and U21865 (N_21865,N_20660,N_19873);
nor U21866 (N_21866,N_20967,N_20442);
nor U21867 (N_21867,N_20965,N_19878);
nor U21868 (N_21868,N_20354,N_20491);
or U21869 (N_21869,N_20407,N_20137);
and U21870 (N_21870,N_19822,N_20288);
nor U21871 (N_21871,N_19648,N_19515);
nor U21872 (N_21872,N_20640,N_20843);
nor U21873 (N_21873,N_20574,N_20049);
nor U21874 (N_21874,N_20103,N_20094);
or U21875 (N_21875,N_20255,N_20165);
nand U21876 (N_21876,N_19673,N_20108);
nand U21877 (N_21877,N_20215,N_20700);
xnor U21878 (N_21878,N_20934,N_20579);
and U21879 (N_21879,N_19532,N_19919);
nand U21880 (N_21880,N_19852,N_20972);
and U21881 (N_21881,N_20243,N_20794);
or U21882 (N_21882,N_20950,N_20784);
nand U21883 (N_21883,N_20923,N_20843);
nand U21884 (N_21884,N_20956,N_20581);
xor U21885 (N_21885,N_19871,N_20010);
or U21886 (N_21886,N_20519,N_19824);
nand U21887 (N_21887,N_19670,N_20113);
nor U21888 (N_21888,N_20097,N_20506);
xor U21889 (N_21889,N_19679,N_19549);
or U21890 (N_21890,N_19699,N_19922);
xor U21891 (N_21891,N_20310,N_20007);
nor U21892 (N_21892,N_19908,N_19705);
and U21893 (N_21893,N_20289,N_20077);
nor U21894 (N_21894,N_19789,N_20266);
xnor U21895 (N_21895,N_20043,N_19533);
nor U21896 (N_21896,N_20134,N_20128);
and U21897 (N_21897,N_20916,N_20515);
or U21898 (N_21898,N_20667,N_20211);
and U21899 (N_21899,N_19624,N_19982);
nor U21900 (N_21900,N_20913,N_20546);
nand U21901 (N_21901,N_20444,N_19531);
and U21902 (N_21902,N_19584,N_19782);
or U21903 (N_21903,N_19541,N_20547);
nor U21904 (N_21904,N_19569,N_20561);
or U21905 (N_21905,N_20345,N_20033);
xor U21906 (N_21906,N_20525,N_20652);
nor U21907 (N_21907,N_20999,N_20945);
nand U21908 (N_21908,N_20391,N_19931);
nor U21909 (N_21909,N_20536,N_19785);
nand U21910 (N_21910,N_20940,N_20908);
nand U21911 (N_21911,N_19847,N_20030);
or U21912 (N_21912,N_20918,N_19606);
xnor U21913 (N_21913,N_20071,N_20369);
and U21914 (N_21914,N_20527,N_20396);
nand U21915 (N_21915,N_20086,N_20303);
or U21916 (N_21916,N_20752,N_20398);
nor U21917 (N_21917,N_20958,N_19933);
xor U21918 (N_21918,N_19515,N_19605);
or U21919 (N_21919,N_20013,N_20601);
or U21920 (N_21920,N_20344,N_20817);
nor U21921 (N_21921,N_20568,N_20603);
or U21922 (N_21922,N_19766,N_19581);
nor U21923 (N_21923,N_19544,N_20195);
nor U21924 (N_21924,N_20974,N_20659);
nor U21925 (N_21925,N_20956,N_20445);
xnor U21926 (N_21926,N_19688,N_19518);
nor U21927 (N_21927,N_20978,N_20179);
nand U21928 (N_21928,N_19569,N_19803);
nand U21929 (N_21929,N_20376,N_20301);
and U21930 (N_21930,N_20733,N_20796);
nor U21931 (N_21931,N_20599,N_20297);
nor U21932 (N_21932,N_20619,N_20880);
xor U21933 (N_21933,N_20020,N_20470);
and U21934 (N_21934,N_19601,N_20933);
nand U21935 (N_21935,N_20457,N_20248);
xor U21936 (N_21936,N_20416,N_19677);
xnor U21937 (N_21937,N_19903,N_20622);
and U21938 (N_21938,N_20851,N_20670);
nand U21939 (N_21939,N_20370,N_20338);
nor U21940 (N_21940,N_20977,N_20547);
nor U21941 (N_21941,N_19881,N_19681);
and U21942 (N_21942,N_19839,N_20750);
nor U21943 (N_21943,N_20884,N_20341);
or U21944 (N_21944,N_20287,N_20830);
or U21945 (N_21945,N_20312,N_19695);
or U21946 (N_21946,N_19739,N_19607);
or U21947 (N_21947,N_19531,N_19789);
xnor U21948 (N_21948,N_20848,N_20887);
nand U21949 (N_21949,N_19780,N_19908);
and U21950 (N_21950,N_20035,N_19656);
and U21951 (N_21951,N_20502,N_20440);
and U21952 (N_21952,N_19962,N_19517);
xnor U21953 (N_21953,N_20960,N_20333);
nand U21954 (N_21954,N_20529,N_19783);
nand U21955 (N_21955,N_20347,N_20923);
nand U21956 (N_21956,N_20511,N_20172);
or U21957 (N_21957,N_20897,N_19573);
nand U21958 (N_21958,N_20748,N_19560);
nand U21959 (N_21959,N_20634,N_19745);
or U21960 (N_21960,N_20122,N_20520);
nand U21961 (N_21961,N_20464,N_19753);
and U21962 (N_21962,N_20488,N_20576);
and U21963 (N_21963,N_20370,N_20703);
or U21964 (N_21964,N_20004,N_20921);
and U21965 (N_21965,N_19532,N_20098);
nand U21966 (N_21966,N_19954,N_20561);
nor U21967 (N_21967,N_20174,N_19811);
nor U21968 (N_21968,N_20285,N_19501);
or U21969 (N_21969,N_19669,N_20899);
and U21970 (N_21970,N_20985,N_20727);
nand U21971 (N_21971,N_20327,N_20237);
or U21972 (N_21972,N_20717,N_20212);
and U21973 (N_21973,N_20575,N_19658);
xnor U21974 (N_21974,N_20659,N_20609);
nand U21975 (N_21975,N_20529,N_19670);
nor U21976 (N_21976,N_20339,N_20686);
nand U21977 (N_21977,N_19824,N_20326);
and U21978 (N_21978,N_20184,N_20838);
xor U21979 (N_21979,N_19814,N_19808);
and U21980 (N_21980,N_20362,N_20634);
and U21981 (N_21981,N_20060,N_20518);
or U21982 (N_21982,N_20957,N_20338);
nor U21983 (N_21983,N_20275,N_19862);
and U21984 (N_21984,N_20154,N_20413);
nor U21985 (N_21985,N_19798,N_20242);
nor U21986 (N_21986,N_19500,N_20782);
or U21987 (N_21987,N_20499,N_19987);
and U21988 (N_21988,N_20452,N_19996);
or U21989 (N_21989,N_20300,N_20450);
xor U21990 (N_21990,N_20620,N_19677);
nand U21991 (N_21991,N_19950,N_19524);
and U21992 (N_21992,N_19638,N_19890);
nor U21993 (N_21993,N_20141,N_20515);
xor U21994 (N_21994,N_20327,N_20062);
and U21995 (N_21995,N_20412,N_20219);
nand U21996 (N_21996,N_20860,N_20351);
nor U21997 (N_21997,N_19996,N_20462);
nor U21998 (N_21998,N_20199,N_20584);
or U21999 (N_21999,N_20919,N_20015);
and U22000 (N_22000,N_20520,N_19845);
or U22001 (N_22001,N_19818,N_20303);
and U22002 (N_22002,N_19970,N_20580);
and U22003 (N_22003,N_20828,N_20878);
xor U22004 (N_22004,N_19534,N_19763);
or U22005 (N_22005,N_20413,N_20096);
or U22006 (N_22006,N_20829,N_20812);
or U22007 (N_22007,N_19501,N_20033);
and U22008 (N_22008,N_20932,N_19934);
or U22009 (N_22009,N_20945,N_19677);
nand U22010 (N_22010,N_19676,N_20148);
and U22011 (N_22011,N_19908,N_20918);
nand U22012 (N_22012,N_20775,N_20839);
and U22013 (N_22013,N_20891,N_20279);
nand U22014 (N_22014,N_20225,N_20955);
nor U22015 (N_22015,N_19930,N_20508);
and U22016 (N_22016,N_20868,N_20045);
xor U22017 (N_22017,N_20239,N_20737);
xnor U22018 (N_22018,N_19529,N_19881);
nand U22019 (N_22019,N_19897,N_20172);
or U22020 (N_22020,N_19597,N_20402);
and U22021 (N_22021,N_19871,N_20475);
xor U22022 (N_22022,N_20680,N_20743);
or U22023 (N_22023,N_19720,N_19596);
nand U22024 (N_22024,N_19695,N_20567);
nand U22025 (N_22025,N_20495,N_20225);
nor U22026 (N_22026,N_20308,N_20392);
nor U22027 (N_22027,N_20251,N_19890);
and U22028 (N_22028,N_19622,N_20775);
or U22029 (N_22029,N_20856,N_19759);
xnor U22030 (N_22030,N_20713,N_19811);
and U22031 (N_22031,N_20448,N_19746);
and U22032 (N_22032,N_20094,N_20825);
nand U22033 (N_22033,N_19529,N_20973);
and U22034 (N_22034,N_19536,N_19883);
or U22035 (N_22035,N_20440,N_20830);
and U22036 (N_22036,N_19755,N_20375);
nand U22037 (N_22037,N_20664,N_19524);
nor U22038 (N_22038,N_20813,N_19868);
xnor U22039 (N_22039,N_20683,N_19750);
nor U22040 (N_22040,N_20677,N_19775);
or U22041 (N_22041,N_19942,N_20803);
xor U22042 (N_22042,N_20603,N_19989);
nand U22043 (N_22043,N_20174,N_20312);
and U22044 (N_22044,N_19972,N_19592);
and U22045 (N_22045,N_19664,N_20744);
nand U22046 (N_22046,N_19825,N_20871);
xor U22047 (N_22047,N_19610,N_20048);
xnor U22048 (N_22048,N_19943,N_20451);
xnor U22049 (N_22049,N_20346,N_20432);
or U22050 (N_22050,N_19807,N_19586);
nand U22051 (N_22051,N_19939,N_20136);
and U22052 (N_22052,N_20345,N_19703);
xor U22053 (N_22053,N_20073,N_19846);
nor U22054 (N_22054,N_20064,N_19925);
nand U22055 (N_22055,N_19847,N_20045);
xnor U22056 (N_22056,N_20140,N_20324);
nand U22057 (N_22057,N_20432,N_20831);
xor U22058 (N_22058,N_20466,N_20475);
nor U22059 (N_22059,N_20443,N_20564);
or U22060 (N_22060,N_20132,N_19516);
xnor U22061 (N_22061,N_20880,N_20773);
nand U22062 (N_22062,N_20471,N_20292);
and U22063 (N_22063,N_20448,N_19769);
xnor U22064 (N_22064,N_20425,N_19972);
and U22065 (N_22065,N_20135,N_20552);
xnor U22066 (N_22066,N_20284,N_20947);
xor U22067 (N_22067,N_20444,N_20860);
nor U22068 (N_22068,N_20761,N_20952);
xnor U22069 (N_22069,N_19959,N_20982);
nor U22070 (N_22070,N_20928,N_20446);
xnor U22071 (N_22071,N_20315,N_20958);
and U22072 (N_22072,N_19746,N_20054);
xor U22073 (N_22073,N_20714,N_20042);
nor U22074 (N_22074,N_20010,N_19559);
nand U22075 (N_22075,N_19764,N_20433);
nand U22076 (N_22076,N_20837,N_19575);
and U22077 (N_22077,N_20686,N_19836);
and U22078 (N_22078,N_19607,N_19720);
nor U22079 (N_22079,N_19846,N_20549);
or U22080 (N_22080,N_20102,N_20408);
nor U22081 (N_22081,N_20234,N_20282);
nor U22082 (N_22082,N_20674,N_19533);
and U22083 (N_22083,N_20572,N_20674);
nor U22084 (N_22084,N_19775,N_20216);
and U22085 (N_22085,N_20900,N_20131);
nor U22086 (N_22086,N_20626,N_20347);
or U22087 (N_22087,N_20419,N_19656);
xnor U22088 (N_22088,N_20678,N_20290);
nor U22089 (N_22089,N_20760,N_19688);
nand U22090 (N_22090,N_20420,N_20105);
and U22091 (N_22091,N_20352,N_20787);
nor U22092 (N_22092,N_19697,N_19522);
nand U22093 (N_22093,N_20711,N_20616);
nor U22094 (N_22094,N_20218,N_19905);
and U22095 (N_22095,N_20171,N_19594);
nand U22096 (N_22096,N_19957,N_20619);
nor U22097 (N_22097,N_20807,N_20978);
nand U22098 (N_22098,N_19678,N_19861);
xor U22099 (N_22099,N_20022,N_19761);
or U22100 (N_22100,N_20099,N_19528);
xnor U22101 (N_22101,N_19607,N_20979);
nor U22102 (N_22102,N_20796,N_19735);
or U22103 (N_22103,N_20345,N_20133);
nand U22104 (N_22104,N_20363,N_20112);
nor U22105 (N_22105,N_19558,N_19586);
nand U22106 (N_22106,N_20874,N_20916);
or U22107 (N_22107,N_19868,N_20777);
or U22108 (N_22108,N_19696,N_20339);
nand U22109 (N_22109,N_20425,N_20061);
or U22110 (N_22110,N_20488,N_20454);
xnor U22111 (N_22111,N_20133,N_19687);
nor U22112 (N_22112,N_20341,N_20206);
or U22113 (N_22113,N_19533,N_20304);
nor U22114 (N_22114,N_19697,N_19904);
nor U22115 (N_22115,N_20340,N_19541);
nor U22116 (N_22116,N_20394,N_19670);
nor U22117 (N_22117,N_19865,N_19992);
and U22118 (N_22118,N_19684,N_19916);
or U22119 (N_22119,N_19879,N_20361);
and U22120 (N_22120,N_20292,N_20908);
nand U22121 (N_22121,N_19692,N_19573);
nor U22122 (N_22122,N_19503,N_19608);
nand U22123 (N_22123,N_20811,N_19549);
or U22124 (N_22124,N_19837,N_19919);
xnor U22125 (N_22125,N_19987,N_19570);
nand U22126 (N_22126,N_20295,N_19679);
nand U22127 (N_22127,N_19526,N_20561);
nand U22128 (N_22128,N_20892,N_19760);
nor U22129 (N_22129,N_20034,N_19571);
or U22130 (N_22130,N_20845,N_19581);
nand U22131 (N_22131,N_20251,N_20455);
nand U22132 (N_22132,N_20294,N_20184);
xor U22133 (N_22133,N_20162,N_19969);
or U22134 (N_22134,N_20102,N_19537);
nor U22135 (N_22135,N_20486,N_19918);
xnor U22136 (N_22136,N_19696,N_20126);
nor U22137 (N_22137,N_20058,N_20207);
nand U22138 (N_22138,N_20870,N_20075);
and U22139 (N_22139,N_19982,N_19711);
and U22140 (N_22140,N_20761,N_19910);
nand U22141 (N_22141,N_20517,N_20797);
and U22142 (N_22142,N_20223,N_20389);
and U22143 (N_22143,N_19923,N_19705);
nand U22144 (N_22144,N_20114,N_20688);
xor U22145 (N_22145,N_20614,N_20813);
and U22146 (N_22146,N_20027,N_19704);
xor U22147 (N_22147,N_20647,N_20052);
nor U22148 (N_22148,N_19765,N_20415);
xor U22149 (N_22149,N_20810,N_19870);
nand U22150 (N_22150,N_20721,N_19523);
nand U22151 (N_22151,N_20411,N_20177);
nand U22152 (N_22152,N_20796,N_20504);
nor U22153 (N_22153,N_20514,N_19587);
xnor U22154 (N_22154,N_20367,N_19905);
nor U22155 (N_22155,N_19527,N_20688);
nor U22156 (N_22156,N_20859,N_20027);
and U22157 (N_22157,N_19935,N_19633);
xnor U22158 (N_22158,N_20737,N_20294);
nand U22159 (N_22159,N_19649,N_20855);
nand U22160 (N_22160,N_20080,N_20807);
or U22161 (N_22161,N_20561,N_20984);
and U22162 (N_22162,N_19978,N_20173);
and U22163 (N_22163,N_20437,N_20150);
or U22164 (N_22164,N_20911,N_20966);
nor U22165 (N_22165,N_20280,N_19700);
nand U22166 (N_22166,N_20570,N_19696);
nor U22167 (N_22167,N_20452,N_19859);
xor U22168 (N_22168,N_20848,N_19920);
or U22169 (N_22169,N_20911,N_20092);
nor U22170 (N_22170,N_19770,N_20172);
nor U22171 (N_22171,N_20509,N_20011);
and U22172 (N_22172,N_20480,N_20165);
and U22173 (N_22173,N_20693,N_20428);
nor U22174 (N_22174,N_20480,N_20475);
nor U22175 (N_22175,N_19958,N_20964);
nand U22176 (N_22176,N_20621,N_19964);
and U22177 (N_22177,N_19628,N_19859);
xnor U22178 (N_22178,N_20776,N_20591);
nand U22179 (N_22179,N_19905,N_20967);
and U22180 (N_22180,N_19856,N_20048);
nor U22181 (N_22181,N_19901,N_19725);
nor U22182 (N_22182,N_19650,N_20476);
xor U22183 (N_22183,N_20118,N_20437);
or U22184 (N_22184,N_20063,N_19674);
or U22185 (N_22185,N_19523,N_20633);
and U22186 (N_22186,N_20098,N_19664);
xor U22187 (N_22187,N_20150,N_19804);
and U22188 (N_22188,N_20377,N_19572);
or U22189 (N_22189,N_20739,N_20443);
nor U22190 (N_22190,N_20910,N_20956);
and U22191 (N_22191,N_20480,N_20002);
nor U22192 (N_22192,N_20948,N_20669);
xnor U22193 (N_22193,N_20606,N_20827);
nand U22194 (N_22194,N_20173,N_20409);
and U22195 (N_22195,N_20945,N_20151);
xor U22196 (N_22196,N_20666,N_19841);
and U22197 (N_22197,N_19566,N_20691);
nor U22198 (N_22198,N_20061,N_20052);
nor U22199 (N_22199,N_19811,N_20516);
or U22200 (N_22200,N_20618,N_19967);
xor U22201 (N_22201,N_20561,N_20418);
or U22202 (N_22202,N_19860,N_20337);
and U22203 (N_22203,N_19519,N_20252);
and U22204 (N_22204,N_20364,N_20592);
nand U22205 (N_22205,N_19967,N_20166);
xnor U22206 (N_22206,N_19863,N_20537);
nor U22207 (N_22207,N_20353,N_20469);
xor U22208 (N_22208,N_20285,N_20017);
xnor U22209 (N_22209,N_20474,N_19993);
xor U22210 (N_22210,N_20412,N_19614);
nor U22211 (N_22211,N_20551,N_20830);
nand U22212 (N_22212,N_19775,N_20939);
xor U22213 (N_22213,N_20113,N_19952);
and U22214 (N_22214,N_19966,N_20364);
nand U22215 (N_22215,N_19829,N_20394);
xor U22216 (N_22216,N_20278,N_20581);
nor U22217 (N_22217,N_20844,N_20688);
nand U22218 (N_22218,N_20337,N_20907);
or U22219 (N_22219,N_20875,N_19914);
xor U22220 (N_22220,N_20568,N_20160);
and U22221 (N_22221,N_20883,N_19881);
or U22222 (N_22222,N_19698,N_20122);
nand U22223 (N_22223,N_20274,N_20256);
nor U22224 (N_22224,N_20253,N_19762);
or U22225 (N_22225,N_20007,N_20347);
xor U22226 (N_22226,N_20377,N_20028);
and U22227 (N_22227,N_20619,N_20138);
and U22228 (N_22228,N_20432,N_20544);
and U22229 (N_22229,N_19633,N_20431);
and U22230 (N_22230,N_20132,N_19629);
xnor U22231 (N_22231,N_19888,N_19614);
nor U22232 (N_22232,N_20311,N_20545);
nand U22233 (N_22233,N_19719,N_19705);
xor U22234 (N_22234,N_20992,N_20847);
or U22235 (N_22235,N_19792,N_20412);
and U22236 (N_22236,N_19830,N_20459);
xor U22237 (N_22237,N_20645,N_19652);
or U22238 (N_22238,N_20071,N_20854);
nand U22239 (N_22239,N_19539,N_20547);
or U22240 (N_22240,N_20157,N_19885);
nand U22241 (N_22241,N_19941,N_20005);
nand U22242 (N_22242,N_20404,N_20651);
and U22243 (N_22243,N_19501,N_20684);
or U22244 (N_22244,N_19664,N_19847);
xor U22245 (N_22245,N_19582,N_20926);
and U22246 (N_22246,N_19940,N_19931);
and U22247 (N_22247,N_20963,N_20651);
or U22248 (N_22248,N_20059,N_20813);
xnor U22249 (N_22249,N_19548,N_20619);
xnor U22250 (N_22250,N_20810,N_19818);
nor U22251 (N_22251,N_20784,N_20737);
and U22252 (N_22252,N_20277,N_19556);
and U22253 (N_22253,N_19911,N_20840);
and U22254 (N_22254,N_20875,N_19538);
and U22255 (N_22255,N_20456,N_20633);
xor U22256 (N_22256,N_20640,N_20504);
nor U22257 (N_22257,N_20656,N_20997);
and U22258 (N_22258,N_19597,N_19634);
and U22259 (N_22259,N_19726,N_19927);
xor U22260 (N_22260,N_19589,N_20914);
xor U22261 (N_22261,N_19802,N_19842);
and U22262 (N_22262,N_19544,N_20666);
xor U22263 (N_22263,N_20685,N_19894);
or U22264 (N_22264,N_20275,N_20035);
or U22265 (N_22265,N_19532,N_20990);
and U22266 (N_22266,N_20509,N_20300);
nand U22267 (N_22267,N_19925,N_20272);
xor U22268 (N_22268,N_20178,N_20295);
and U22269 (N_22269,N_19687,N_19921);
and U22270 (N_22270,N_20812,N_20651);
and U22271 (N_22271,N_19642,N_19789);
nand U22272 (N_22272,N_20271,N_19500);
or U22273 (N_22273,N_20339,N_19738);
and U22274 (N_22274,N_20222,N_20666);
nor U22275 (N_22275,N_20965,N_19894);
xnor U22276 (N_22276,N_19512,N_20440);
xnor U22277 (N_22277,N_20452,N_19866);
nand U22278 (N_22278,N_20948,N_19877);
nand U22279 (N_22279,N_19832,N_19817);
xor U22280 (N_22280,N_19981,N_20000);
xnor U22281 (N_22281,N_19867,N_19883);
and U22282 (N_22282,N_20911,N_20728);
or U22283 (N_22283,N_19612,N_19747);
nor U22284 (N_22284,N_20835,N_20075);
or U22285 (N_22285,N_20133,N_20336);
and U22286 (N_22286,N_19857,N_20207);
or U22287 (N_22287,N_20507,N_19879);
nand U22288 (N_22288,N_20502,N_20238);
nand U22289 (N_22289,N_20102,N_20819);
or U22290 (N_22290,N_19699,N_20960);
or U22291 (N_22291,N_20052,N_19997);
and U22292 (N_22292,N_19797,N_20754);
nand U22293 (N_22293,N_20915,N_20191);
and U22294 (N_22294,N_19826,N_19670);
nand U22295 (N_22295,N_19772,N_20011);
nand U22296 (N_22296,N_20101,N_20625);
and U22297 (N_22297,N_20180,N_20665);
and U22298 (N_22298,N_20550,N_19623);
xnor U22299 (N_22299,N_20593,N_20258);
xor U22300 (N_22300,N_20906,N_19973);
and U22301 (N_22301,N_20484,N_20057);
nand U22302 (N_22302,N_20701,N_20183);
and U22303 (N_22303,N_20604,N_19716);
or U22304 (N_22304,N_19803,N_19931);
nor U22305 (N_22305,N_19535,N_20864);
or U22306 (N_22306,N_20807,N_20085);
and U22307 (N_22307,N_20927,N_20265);
nor U22308 (N_22308,N_19544,N_20748);
or U22309 (N_22309,N_20225,N_19660);
xor U22310 (N_22310,N_20428,N_20828);
nor U22311 (N_22311,N_20698,N_20738);
and U22312 (N_22312,N_20711,N_20185);
nor U22313 (N_22313,N_20695,N_19854);
xor U22314 (N_22314,N_19566,N_20759);
and U22315 (N_22315,N_20662,N_20607);
or U22316 (N_22316,N_19636,N_20327);
or U22317 (N_22317,N_20992,N_20057);
xor U22318 (N_22318,N_20363,N_20415);
or U22319 (N_22319,N_19852,N_19747);
nor U22320 (N_22320,N_19996,N_19813);
xor U22321 (N_22321,N_20173,N_20482);
or U22322 (N_22322,N_19549,N_20440);
or U22323 (N_22323,N_19764,N_20207);
nor U22324 (N_22324,N_20903,N_19506);
xnor U22325 (N_22325,N_20088,N_20663);
xor U22326 (N_22326,N_19591,N_20482);
and U22327 (N_22327,N_20527,N_19629);
and U22328 (N_22328,N_19572,N_20898);
or U22329 (N_22329,N_20854,N_20538);
or U22330 (N_22330,N_19561,N_20676);
nand U22331 (N_22331,N_20954,N_20337);
or U22332 (N_22332,N_20442,N_20474);
nand U22333 (N_22333,N_20879,N_20041);
nand U22334 (N_22334,N_20788,N_19586);
nor U22335 (N_22335,N_20165,N_20174);
nor U22336 (N_22336,N_20605,N_19677);
and U22337 (N_22337,N_19603,N_19747);
or U22338 (N_22338,N_20607,N_20112);
nor U22339 (N_22339,N_19730,N_20958);
and U22340 (N_22340,N_19545,N_20920);
nand U22341 (N_22341,N_20267,N_19656);
and U22342 (N_22342,N_19995,N_19865);
xor U22343 (N_22343,N_19935,N_19824);
and U22344 (N_22344,N_19839,N_20890);
and U22345 (N_22345,N_19837,N_19681);
or U22346 (N_22346,N_20108,N_19605);
nand U22347 (N_22347,N_20856,N_19541);
or U22348 (N_22348,N_20514,N_19873);
nor U22349 (N_22349,N_19821,N_20203);
xnor U22350 (N_22350,N_20453,N_20214);
xnor U22351 (N_22351,N_20582,N_20580);
xor U22352 (N_22352,N_20627,N_20523);
and U22353 (N_22353,N_20026,N_19882);
nor U22354 (N_22354,N_20114,N_20481);
nor U22355 (N_22355,N_19768,N_20375);
nand U22356 (N_22356,N_20237,N_20049);
or U22357 (N_22357,N_20460,N_19604);
xor U22358 (N_22358,N_19842,N_20813);
and U22359 (N_22359,N_19679,N_19937);
nand U22360 (N_22360,N_19804,N_20579);
or U22361 (N_22361,N_20704,N_20235);
and U22362 (N_22362,N_20648,N_19623);
nand U22363 (N_22363,N_19928,N_20775);
nand U22364 (N_22364,N_19775,N_19512);
xnor U22365 (N_22365,N_20131,N_19623);
xor U22366 (N_22366,N_20907,N_20536);
xnor U22367 (N_22367,N_20080,N_20813);
xor U22368 (N_22368,N_20474,N_19846);
nand U22369 (N_22369,N_20689,N_20844);
or U22370 (N_22370,N_20587,N_20675);
nand U22371 (N_22371,N_20035,N_20440);
nor U22372 (N_22372,N_20302,N_20574);
xnor U22373 (N_22373,N_20827,N_20541);
xor U22374 (N_22374,N_20987,N_20902);
nand U22375 (N_22375,N_20290,N_19791);
nor U22376 (N_22376,N_19588,N_20878);
xor U22377 (N_22377,N_19921,N_19706);
xor U22378 (N_22378,N_20436,N_19656);
nand U22379 (N_22379,N_20625,N_20240);
xnor U22380 (N_22380,N_19900,N_20062);
and U22381 (N_22381,N_20251,N_20621);
nor U22382 (N_22382,N_20564,N_20979);
nor U22383 (N_22383,N_19967,N_20728);
nand U22384 (N_22384,N_20662,N_19721);
or U22385 (N_22385,N_20686,N_20882);
and U22386 (N_22386,N_20234,N_20444);
nand U22387 (N_22387,N_19705,N_19765);
nor U22388 (N_22388,N_20827,N_20018);
nand U22389 (N_22389,N_19774,N_19953);
nor U22390 (N_22390,N_19836,N_20927);
and U22391 (N_22391,N_20165,N_19823);
nand U22392 (N_22392,N_19588,N_20332);
nand U22393 (N_22393,N_19500,N_19561);
or U22394 (N_22394,N_20009,N_20339);
and U22395 (N_22395,N_19963,N_20261);
nor U22396 (N_22396,N_20644,N_20420);
and U22397 (N_22397,N_20984,N_19692);
xor U22398 (N_22398,N_19841,N_20067);
nand U22399 (N_22399,N_20863,N_19504);
nand U22400 (N_22400,N_19566,N_20125);
xnor U22401 (N_22401,N_20795,N_20110);
nand U22402 (N_22402,N_20634,N_20824);
and U22403 (N_22403,N_20302,N_20058);
nand U22404 (N_22404,N_19724,N_20227);
nand U22405 (N_22405,N_20797,N_19648);
and U22406 (N_22406,N_20322,N_19744);
or U22407 (N_22407,N_20648,N_20335);
xnor U22408 (N_22408,N_19807,N_20844);
or U22409 (N_22409,N_20969,N_19853);
xor U22410 (N_22410,N_20497,N_20502);
or U22411 (N_22411,N_20946,N_19551);
xnor U22412 (N_22412,N_19743,N_19770);
nor U22413 (N_22413,N_20802,N_20482);
and U22414 (N_22414,N_19949,N_19956);
xnor U22415 (N_22415,N_20865,N_19714);
nor U22416 (N_22416,N_20550,N_19882);
nand U22417 (N_22417,N_20766,N_20824);
nor U22418 (N_22418,N_20189,N_20493);
nand U22419 (N_22419,N_19554,N_20429);
or U22420 (N_22420,N_20788,N_19991);
nor U22421 (N_22421,N_20383,N_19998);
or U22422 (N_22422,N_20142,N_19974);
and U22423 (N_22423,N_20199,N_20273);
and U22424 (N_22424,N_19870,N_20078);
or U22425 (N_22425,N_19512,N_19930);
nor U22426 (N_22426,N_19999,N_20234);
nand U22427 (N_22427,N_20696,N_20818);
nand U22428 (N_22428,N_20098,N_20894);
xor U22429 (N_22429,N_20413,N_19850);
nand U22430 (N_22430,N_20446,N_20951);
nand U22431 (N_22431,N_20944,N_19723);
nand U22432 (N_22432,N_20803,N_20997);
or U22433 (N_22433,N_20055,N_19916);
nor U22434 (N_22434,N_20337,N_20078);
xor U22435 (N_22435,N_19714,N_20361);
or U22436 (N_22436,N_19510,N_20182);
and U22437 (N_22437,N_19726,N_19551);
or U22438 (N_22438,N_20163,N_20869);
and U22439 (N_22439,N_19582,N_20386);
nand U22440 (N_22440,N_20326,N_20085);
or U22441 (N_22441,N_19910,N_20324);
xor U22442 (N_22442,N_19989,N_19586);
nor U22443 (N_22443,N_20471,N_20577);
and U22444 (N_22444,N_20386,N_20842);
or U22445 (N_22445,N_20633,N_19947);
and U22446 (N_22446,N_20754,N_20977);
and U22447 (N_22447,N_20881,N_20593);
and U22448 (N_22448,N_19738,N_20967);
and U22449 (N_22449,N_20677,N_19875);
or U22450 (N_22450,N_20992,N_19630);
nor U22451 (N_22451,N_20040,N_20841);
nand U22452 (N_22452,N_19551,N_20622);
and U22453 (N_22453,N_20502,N_19801);
or U22454 (N_22454,N_20695,N_20064);
nand U22455 (N_22455,N_20904,N_20253);
or U22456 (N_22456,N_20568,N_20506);
or U22457 (N_22457,N_20983,N_19961);
and U22458 (N_22458,N_19703,N_19764);
xnor U22459 (N_22459,N_19623,N_19591);
nor U22460 (N_22460,N_20564,N_20974);
and U22461 (N_22461,N_20715,N_20796);
or U22462 (N_22462,N_19830,N_19856);
nor U22463 (N_22463,N_20804,N_20208);
xnor U22464 (N_22464,N_20134,N_20092);
or U22465 (N_22465,N_19693,N_19950);
xnor U22466 (N_22466,N_19692,N_20855);
nand U22467 (N_22467,N_19949,N_19751);
and U22468 (N_22468,N_19536,N_20712);
and U22469 (N_22469,N_19999,N_20488);
nand U22470 (N_22470,N_20229,N_20132);
nor U22471 (N_22471,N_20904,N_20177);
and U22472 (N_22472,N_20050,N_20533);
or U22473 (N_22473,N_19985,N_20927);
xnor U22474 (N_22474,N_20397,N_19955);
or U22475 (N_22475,N_20720,N_19964);
xnor U22476 (N_22476,N_20711,N_20042);
or U22477 (N_22477,N_19772,N_19516);
nand U22478 (N_22478,N_19944,N_20881);
xnor U22479 (N_22479,N_20427,N_19941);
xnor U22480 (N_22480,N_20302,N_20837);
and U22481 (N_22481,N_19800,N_20292);
nand U22482 (N_22482,N_20844,N_20458);
nor U22483 (N_22483,N_20452,N_19820);
nand U22484 (N_22484,N_20268,N_19597);
and U22485 (N_22485,N_20136,N_20965);
nor U22486 (N_22486,N_20389,N_20967);
or U22487 (N_22487,N_19979,N_20278);
and U22488 (N_22488,N_20780,N_19555);
xnor U22489 (N_22489,N_20084,N_20815);
xor U22490 (N_22490,N_20367,N_19949);
or U22491 (N_22491,N_19890,N_20732);
nor U22492 (N_22492,N_20683,N_20579);
or U22493 (N_22493,N_19525,N_19549);
xor U22494 (N_22494,N_20680,N_19834);
xnor U22495 (N_22495,N_20084,N_19572);
xnor U22496 (N_22496,N_19696,N_19686);
or U22497 (N_22497,N_19803,N_20280);
xnor U22498 (N_22498,N_19709,N_19837);
nor U22499 (N_22499,N_19951,N_20690);
nor U22500 (N_22500,N_22262,N_21846);
and U22501 (N_22501,N_21129,N_22087);
nand U22502 (N_22502,N_21452,N_21569);
or U22503 (N_22503,N_21494,N_21719);
nand U22504 (N_22504,N_21139,N_22094);
and U22505 (N_22505,N_22301,N_22356);
or U22506 (N_22506,N_22276,N_22225);
nor U22507 (N_22507,N_21708,N_21118);
or U22508 (N_22508,N_21369,N_21660);
or U22509 (N_22509,N_22390,N_22370);
and U22510 (N_22510,N_22347,N_21432);
nor U22511 (N_22511,N_21367,N_21389);
or U22512 (N_22512,N_21021,N_22214);
nand U22513 (N_22513,N_21518,N_22374);
and U22514 (N_22514,N_22027,N_21136);
and U22515 (N_22515,N_21277,N_21720);
nor U22516 (N_22516,N_22336,N_21767);
xor U22517 (N_22517,N_22322,N_21290);
xnor U22518 (N_22518,N_22041,N_21812);
nand U22519 (N_22519,N_21993,N_21566);
nand U22520 (N_22520,N_22070,N_21504);
xnor U22521 (N_22521,N_21605,N_21378);
nand U22522 (N_22522,N_22146,N_21878);
and U22523 (N_22523,N_21934,N_21589);
or U22524 (N_22524,N_21050,N_21687);
nor U22525 (N_22525,N_22499,N_22083);
nand U22526 (N_22526,N_21295,N_21807);
and U22527 (N_22527,N_21827,N_21222);
or U22528 (N_22528,N_21986,N_21525);
nand U22529 (N_22529,N_22335,N_22389);
nand U22530 (N_22530,N_21067,N_21076);
nor U22531 (N_22531,N_22181,N_21310);
xor U22532 (N_22532,N_21955,N_21957);
or U22533 (N_22533,N_21492,N_21113);
xnor U22534 (N_22534,N_21074,N_22427);
xor U22535 (N_22535,N_21411,N_22229);
xnor U22536 (N_22536,N_21022,N_21024);
nor U22537 (N_22537,N_21996,N_21294);
xor U22538 (N_22538,N_22025,N_21739);
xnor U22539 (N_22539,N_21051,N_22393);
and U22540 (N_22540,N_21340,N_21462);
and U22541 (N_22541,N_21166,N_21417);
and U22542 (N_22542,N_21815,N_22194);
or U22543 (N_22543,N_21880,N_21102);
xnor U22544 (N_22544,N_22040,N_22247);
xnor U22545 (N_22545,N_22031,N_21652);
or U22546 (N_22546,N_22477,N_22236);
xor U22547 (N_22547,N_21350,N_21180);
xor U22548 (N_22548,N_22450,N_22490);
nand U22549 (N_22549,N_22260,N_22168);
nand U22550 (N_22550,N_21808,N_21087);
nor U22551 (N_22551,N_22446,N_22483);
and U22552 (N_22552,N_21601,N_22482);
nand U22553 (N_22553,N_22419,N_21564);
and U22554 (N_22554,N_22350,N_21821);
or U22555 (N_22555,N_21012,N_22293);
xor U22556 (N_22556,N_21848,N_21769);
or U22557 (N_22557,N_21949,N_21543);
nand U22558 (N_22558,N_21235,N_21795);
or U22559 (N_22559,N_21321,N_22165);
nand U22560 (N_22560,N_21285,N_21304);
or U22561 (N_22561,N_21202,N_22365);
xor U22562 (N_22562,N_22445,N_22295);
nand U22563 (N_22563,N_21585,N_21635);
and U22564 (N_22564,N_22416,N_22035);
nor U22565 (N_22565,N_22269,N_21770);
xor U22566 (N_22566,N_22357,N_21834);
xor U22567 (N_22567,N_21457,N_21733);
xor U22568 (N_22568,N_21873,N_22144);
nor U22569 (N_22569,N_21555,N_22142);
nand U22570 (N_22570,N_22257,N_21962);
or U22571 (N_22571,N_21211,N_21403);
nand U22572 (N_22572,N_21864,N_22279);
and U22573 (N_22573,N_21649,N_21112);
xor U22574 (N_22574,N_21972,N_21668);
and U22575 (N_22575,N_21381,N_22136);
nor U22576 (N_22576,N_21891,N_21419);
nand U22577 (N_22577,N_21010,N_21742);
and U22578 (N_22578,N_22011,N_21453);
nand U22579 (N_22579,N_21967,N_22020);
xnor U22580 (N_22580,N_22289,N_22046);
or U22581 (N_22581,N_21695,N_21765);
nor U22582 (N_22582,N_21468,N_22329);
xor U22583 (N_22583,N_21630,N_21713);
nand U22584 (N_22584,N_21691,N_22474);
or U22585 (N_22585,N_21942,N_22428);
nor U22586 (N_22586,N_21588,N_22324);
xor U22587 (N_22587,N_22053,N_21528);
xor U22588 (N_22588,N_22263,N_22069);
and U22589 (N_22589,N_21094,N_21485);
xnor U22590 (N_22590,N_22302,N_21465);
or U22591 (N_22591,N_22413,N_21836);
nor U22592 (N_22592,N_21701,N_21308);
or U22593 (N_22593,N_22112,N_21205);
and U22594 (N_22594,N_22415,N_21643);
xor U22595 (N_22595,N_21866,N_21547);
nand U22596 (N_22596,N_21456,N_21008);
and U22597 (N_22597,N_21988,N_21265);
nor U22598 (N_22598,N_21628,N_21000);
and U22599 (N_22599,N_22084,N_22008);
or U22600 (N_22600,N_22206,N_21802);
xnor U22601 (N_22601,N_22023,N_22195);
and U22602 (N_22602,N_21317,N_21029);
nor U22603 (N_22603,N_21443,N_22108);
xnor U22604 (N_22604,N_21859,N_21521);
and U22605 (N_22605,N_21830,N_21358);
and U22606 (N_22606,N_21616,N_21667);
nor U22607 (N_22607,N_22435,N_21120);
and U22608 (N_22608,N_22323,N_21128);
xnor U22609 (N_22609,N_21374,N_22178);
nor U22610 (N_22610,N_21620,N_22352);
and U22611 (N_22611,N_22258,N_21580);
and U22612 (N_22612,N_21441,N_22326);
and U22613 (N_22613,N_22331,N_21751);
or U22614 (N_22614,N_21828,N_22185);
xor U22615 (N_22615,N_21567,N_21420);
or U22616 (N_22616,N_22126,N_21944);
nor U22617 (N_22617,N_22488,N_22368);
and U22618 (N_22618,N_22318,N_22274);
and U22619 (N_22619,N_21216,N_21207);
and U22620 (N_22620,N_21275,N_22213);
or U22621 (N_22621,N_21685,N_21759);
or U22622 (N_22622,N_22117,N_21427);
xor U22623 (N_22623,N_21762,N_21287);
and U22624 (N_22624,N_21445,N_21005);
nor U22625 (N_22625,N_21195,N_21055);
nor U22626 (N_22626,N_22438,N_22066);
xnor U22627 (N_22627,N_21268,N_21814);
and U22628 (N_22628,N_21537,N_21234);
or U22629 (N_22629,N_22306,N_22072);
and U22630 (N_22630,N_21448,N_21423);
xnor U22631 (N_22631,N_21039,N_21710);
and U22632 (N_22632,N_21263,N_21648);
nor U22633 (N_22633,N_22442,N_22086);
xnor U22634 (N_22634,N_21360,N_21338);
and U22635 (N_22635,N_21038,N_21875);
or U22636 (N_22636,N_21159,N_21231);
nor U22637 (N_22637,N_21855,N_21884);
and U22638 (N_22638,N_21831,N_21440);
or U22639 (N_22639,N_21915,N_22182);
or U22640 (N_22640,N_21261,N_21480);
and U22641 (N_22641,N_22469,N_21405);
nor U22642 (N_22642,N_21542,N_22079);
nor U22643 (N_22643,N_21326,N_21804);
nor U22644 (N_22644,N_22243,N_21519);
nor U22645 (N_22645,N_21017,N_21838);
and U22646 (N_22646,N_21653,N_22231);
nand U22647 (N_22647,N_21192,N_21458);
xnor U22648 (N_22648,N_21786,N_22264);
nand U22649 (N_22649,N_22167,N_22360);
nor U22650 (N_22650,N_21533,N_21406);
nand U22651 (N_22651,N_21318,N_21219);
nor U22652 (N_22652,N_21430,N_21396);
nor U22653 (N_22653,N_22139,N_21262);
nor U22654 (N_22654,N_22317,N_22443);
xnor U22655 (N_22655,N_22058,N_21026);
xnor U22656 (N_22656,N_22109,N_21143);
nor U22657 (N_22657,N_21204,N_22340);
nor U22658 (N_22658,N_21953,N_21157);
nand U22659 (N_22659,N_21923,N_22417);
nor U22660 (N_22660,N_21408,N_21587);
nor U22661 (N_22661,N_21945,N_21449);
and U22662 (N_22662,N_21579,N_21981);
or U22663 (N_22663,N_22463,N_21126);
or U22664 (N_22664,N_21033,N_22026);
nand U22665 (N_22665,N_21003,N_21625);
or U22666 (N_22666,N_21174,N_21645);
nor U22667 (N_22667,N_21730,N_22281);
nand U22668 (N_22668,N_21332,N_21015);
or U22669 (N_22669,N_21901,N_21048);
nor U22670 (N_22670,N_22029,N_22134);
and U22671 (N_22671,N_21886,N_21935);
xnor U22672 (N_22672,N_21897,N_21927);
nand U22673 (N_22673,N_21218,N_21930);
xnor U22674 (N_22674,N_22003,N_22275);
nand U22675 (N_22675,N_21303,N_21858);
xnor U22676 (N_22676,N_22201,N_21467);
xnor U22677 (N_22677,N_21602,N_22047);
and U22678 (N_22678,N_21345,N_21170);
nand U22679 (N_22679,N_21783,N_22158);
and U22680 (N_22680,N_21096,N_22176);
or U22681 (N_22681,N_21870,N_22400);
nand U22682 (N_22682,N_21243,N_21357);
nand U22683 (N_22683,N_21254,N_21570);
nand U22684 (N_22684,N_21178,N_21179);
and U22685 (N_22685,N_22486,N_21309);
nand U22686 (N_22686,N_21760,N_21747);
xnor U22687 (N_22687,N_21684,N_22152);
and U22688 (N_22688,N_21793,N_21172);
nand U22689 (N_22689,N_21508,N_21851);
nor U22690 (N_22690,N_21908,N_21553);
nand U22691 (N_22691,N_21737,N_22346);
nor U22692 (N_22692,N_22161,N_21711);
xnor U22693 (N_22693,N_22485,N_22454);
xnor U22694 (N_22694,N_21604,N_22191);
and U22695 (N_22695,N_21593,N_22479);
nand U22696 (N_22696,N_22385,N_22493);
xor U22697 (N_22697,N_21210,N_21249);
nor U22698 (N_22698,N_22074,N_22123);
and U22699 (N_22699,N_22044,N_21982);
xnor U22700 (N_22700,N_22437,N_22267);
and U22701 (N_22701,N_22272,N_22314);
nand U22702 (N_22702,N_21819,N_22433);
xor U22703 (N_22703,N_22291,N_21612);
or U22704 (N_22704,N_21772,N_21924);
nand U22705 (N_22705,N_21370,N_21712);
nand U22706 (N_22706,N_21557,N_21341);
or U22707 (N_22707,N_21777,N_22043);
xor U22708 (N_22708,N_21415,N_21101);
nand U22709 (N_22709,N_21946,N_22464);
nand U22710 (N_22710,N_21191,N_21284);
or U22711 (N_22711,N_22071,N_22101);
xnor U22712 (N_22712,N_21344,N_22480);
nand U22713 (N_22713,N_22177,N_21108);
and U22714 (N_22714,N_21450,N_21068);
xor U22715 (N_22715,N_21914,N_21895);
and U22716 (N_22716,N_22021,N_21572);
or U22717 (N_22717,N_22359,N_21385);
or U22718 (N_22718,N_21699,N_22160);
nor U22719 (N_22719,N_21562,N_22062);
xnor U22720 (N_22720,N_21203,N_22294);
or U22721 (N_22721,N_22197,N_22386);
and U22722 (N_22722,N_22492,N_21790);
nor U22723 (N_22723,N_21874,N_21661);
or U22724 (N_22724,N_21069,N_22384);
or U22725 (N_22725,N_21435,N_21496);
or U22726 (N_22726,N_22497,N_21619);
nor U22727 (N_22727,N_22457,N_22354);
and U22728 (N_22728,N_22494,N_22290);
nor U22729 (N_22729,N_21410,N_22406);
xor U22730 (N_22730,N_21049,N_21407);
and U22731 (N_22731,N_21577,N_21843);
nor U22732 (N_22732,N_22127,N_21912);
and U22733 (N_22733,N_21715,N_21184);
nand U22734 (N_22734,N_21266,N_22075);
nand U22735 (N_22735,N_21740,N_21288);
and U22736 (N_22736,N_21473,N_21522);
and U22737 (N_22737,N_22312,N_21200);
or U22738 (N_22738,N_22447,N_21928);
nand U22739 (N_22739,N_22371,N_21255);
nand U22740 (N_22740,N_21089,N_21847);
nand U22741 (N_22741,N_21548,N_21158);
xnor U22742 (N_22742,N_21095,N_21177);
and U22743 (N_22743,N_21488,N_21491);
or U22744 (N_22744,N_21539,N_21926);
xor U22745 (N_22745,N_21119,N_21313);
nand U22746 (N_22746,N_21745,N_22148);
xnor U22747 (N_22747,N_21165,N_21659);
xnor U22748 (N_22748,N_22407,N_22451);
nor U22749 (N_22749,N_21671,N_21489);
nor U22750 (N_22750,N_21565,N_21399);
and U22751 (N_22751,N_21214,N_21030);
nand U22752 (N_22752,N_21623,N_22078);
xnor U22753 (N_22753,N_22455,N_21330);
xor U22754 (N_22754,N_21617,N_21983);
xnor U22755 (N_22755,N_21826,N_22475);
nand U22756 (N_22756,N_21753,N_21193);
nand U22757 (N_22757,N_22064,N_21738);
or U22758 (N_22758,N_21531,N_22124);
nor U22759 (N_22759,N_21852,N_22018);
or U22760 (N_22760,N_21797,N_22284);
and U22761 (N_22761,N_21999,N_21006);
or U22762 (N_22762,N_22448,N_22458);
nand U22763 (N_22763,N_21123,N_22327);
or U22764 (N_22764,N_21868,N_21362);
nor U22765 (N_22765,N_21657,N_22296);
and U22766 (N_22766,N_21818,N_22147);
nor U22767 (N_22767,N_22280,N_21975);
xor U22768 (N_22768,N_21558,N_21434);
or U22769 (N_22769,N_21627,N_22141);
nand U22770 (N_22770,N_21142,N_21257);
or U22771 (N_22771,N_22364,N_21299);
xnor U22772 (N_22772,N_22230,N_21312);
or U22773 (N_22773,N_21887,N_21196);
nand U22774 (N_22774,N_22391,N_22246);
nor U22775 (N_22775,N_21264,N_21844);
and U22776 (N_22776,N_21798,N_21433);
nor U22777 (N_22777,N_22471,N_21991);
or U22778 (N_22778,N_21025,N_21510);
xor U22779 (N_22779,N_21272,N_22042);
nand U22780 (N_22780,N_21071,N_22200);
and U22781 (N_22781,N_21327,N_21755);
xor U22782 (N_22782,N_21757,N_21640);
or U22783 (N_22783,N_22319,N_21535);
nand U22784 (N_22784,N_21280,N_21780);
xnor U22785 (N_22785,N_22234,N_22169);
or U22786 (N_22786,N_22004,N_22399);
nor U22787 (N_22787,N_21469,N_21151);
xor U22788 (N_22788,N_21386,N_21032);
and U22789 (N_22789,N_21359,N_21692);
nand U22790 (N_22790,N_21484,N_21933);
or U22791 (N_22791,N_21938,N_22138);
xor U22792 (N_22792,N_21961,N_22355);
xor U22793 (N_22793,N_21404,N_21621);
and U22794 (N_22794,N_22221,N_21689);
xor U22795 (N_22795,N_22128,N_21801);
nor U22796 (N_22796,N_22362,N_22189);
nor U22797 (N_22797,N_21954,N_21906);
xnor U22798 (N_22798,N_21225,N_22107);
xnor U22799 (N_22799,N_22421,N_22216);
and U22800 (N_22800,N_22135,N_22220);
xnor U22801 (N_22801,N_22394,N_21850);
nor U22802 (N_22802,N_21511,N_22052);
nand U22803 (N_22803,N_22367,N_21040);
xnor U22804 (N_22804,N_21872,N_21631);
xor U22805 (N_22805,N_21590,N_22305);
nor U22806 (N_22806,N_22015,N_21086);
xor U22807 (N_22807,N_21075,N_21789);
and U22808 (N_22808,N_21431,N_22111);
nand U22809 (N_22809,N_21414,N_21976);
nor U22810 (N_22810,N_22311,N_22383);
or U22811 (N_22811,N_21822,N_21909);
nand U22812 (N_22812,N_22038,N_21883);
and U22813 (N_22813,N_21726,N_21175);
xnor U22814 (N_22814,N_22113,N_22186);
nand U22815 (N_22815,N_21810,N_22095);
or U22816 (N_22816,N_21472,N_21641);
xor U22817 (N_22817,N_21141,N_21479);
xor U22818 (N_22818,N_22478,N_21764);
or U22819 (N_22819,N_21931,N_22163);
and U22820 (N_22820,N_21232,N_21248);
xnor U22821 (N_22821,N_21238,N_21893);
or U22822 (N_22822,N_22024,N_21741);
xnor U22823 (N_22823,N_21632,N_22405);
xor U22824 (N_22824,N_21512,N_21167);
xor U22825 (N_22825,N_21352,N_21754);
or U22826 (N_22826,N_21674,N_22208);
nor U22827 (N_22827,N_21160,N_21364);
and U22828 (N_22828,N_21477,N_22174);
nand U22829 (N_22829,N_22143,N_22430);
nand U22830 (N_22830,N_22059,N_21347);
xor U22831 (N_22831,N_21995,N_21985);
xnor U22832 (N_22832,N_22204,N_21148);
or U22833 (N_22833,N_21245,N_22366);
nand U22834 (N_22834,N_21584,N_21929);
or U22835 (N_22835,N_21220,N_22097);
xor U22836 (N_22836,N_21323,N_21233);
or U22837 (N_22837,N_22106,N_21438);
nand U22838 (N_22838,N_22397,N_22233);
nor U22839 (N_22839,N_21085,N_21293);
or U22840 (N_22840,N_21824,N_21215);
or U22841 (N_22841,N_21394,N_21376);
or U22842 (N_22842,N_21446,N_21763);
and U22843 (N_22843,N_21305,N_21916);
and U22844 (N_22844,N_22104,N_21718);
nand U22845 (N_22845,N_22150,N_21125);
nand U22846 (N_22846,N_22321,N_21031);
and U22847 (N_22847,N_21375,N_22441);
or U22848 (N_22848,N_21573,N_21199);
nor U22849 (N_22849,N_21919,N_22218);
nand U22850 (N_22850,N_22432,N_21459);
nand U22851 (N_22851,N_22100,N_22209);
nor U22852 (N_22852,N_21816,N_21937);
nor U22853 (N_22853,N_22298,N_21925);
or U22854 (N_22854,N_21865,N_21273);
xnor U22855 (N_22855,N_21613,N_21292);
and U22856 (N_22856,N_21561,N_21133);
or U22857 (N_22857,N_21036,N_21529);
or U22858 (N_22858,N_21343,N_21324);
nor U22859 (N_22859,N_22116,N_21703);
nor U22860 (N_22860,N_21059,N_21839);
or U22861 (N_22861,N_21956,N_21224);
xor U22862 (N_22862,N_21781,N_21560);
nand U22863 (N_22863,N_22080,N_21092);
nand U22864 (N_22864,N_21351,N_21088);
nand U22865 (N_22865,N_21725,N_21278);
and U22866 (N_22866,N_21698,N_22422);
nor U22867 (N_22867,N_21490,N_21794);
nor U22868 (N_22868,N_21559,N_21785);
or U22869 (N_22869,N_21965,N_22122);
nor U22870 (N_22870,N_22120,N_21515);
nand U22871 (N_22871,N_21065,N_21735);
xnor U22872 (N_22872,N_22270,N_22251);
or U22873 (N_22873,N_21514,N_22105);
and U22874 (N_22874,N_22034,N_21973);
and U22875 (N_22875,N_21422,N_21958);
nor U22876 (N_22876,N_21974,N_21672);
and U22877 (N_22877,N_21892,N_21941);
xnor U22878 (N_22878,N_21451,N_21670);
or U22879 (N_22879,N_21609,N_21551);
and U22880 (N_22880,N_21888,N_21968);
nand U22881 (N_22881,N_22308,N_22103);
or U22882 (N_22882,N_21917,N_21042);
xnor U22883 (N_22883,N_21047,N_22093);
and U22884 (N_22884,N_22198,N_22363);
or U22885 (N_22885,N_21348,N_21260);
xor U22886 (N_22886,N_21329,N_21913);
nand U22887 (N_22887,N_21900,N_21549);
nor U22888 (N_22888,N_21259,N_21773);
nand U22889 (N_22889,N_22292,N_21070);
xnor U22890 (N_22890,N_22013,N_21882);
xor U22891 (N_22891,N_22090,N_21185);
nor U22892 (N_22892,N_22465,N_22248);
or U22893 (N_22893,N_21250,N_21501);
nand U22894 (N_22894,N_21610,N_21335);
nor U22895 (N_22895,N_21252,N_22408);
nand U22896 (N_22896,N_21107,N_22098);
or U22897 (N_22897,N_21817,N_22332);
nand U22898 (N_22898,N_22440,N_22330);
nand U22899 (N_22899,N_21466,N_21750);
nand U22900 (N_22900,N_21992,N_22472);
nor U22901 (N_22901,N_21534,N_21189);
nand U22902 (N_22902,N_21183,N_22050);
nand U22903 (N_22903,N_22283,N_21444);
and U22904 (N_22904,N_21655,N_21461);
or U22905 (N_22905,N_21651,N_21397);
nand U22906 (N_22906,N_22351,N_21099);
nand U22907 (N_22907,N_21806,N_21503);
nor U22908 (N_22908,N_22310,N_21586);
nand U22909 (N_22909,N_22468,N_21532);
nor U22910 (N_22910,N_21182,N_21775);
xnor U22911 (N_22911,N_21455,N_21282);
and U22912 (N_22912,N_21550,N_21083);
nor U22913 (N_22913,N_21023,N_21028);
or U22914 (N_22914,N_21731,N_21540);
nand U22915 (N_22915,N_21236,N_21857);
nand U22916 (N_22916,N_22240,N_21054);
xnor U22917 (N_22917,N_21592,N_21497);
nand U22918 (N_22918,N_21471,N_21943);
and U22919 (N_22919,N_21482,N_21948);
or U22920 (N_22920,N_21634,N_22048);
nand U22921 (N_22921,N_22166,N_21131);
nor U22922 (N_22922,N_22487,N_22156);
nor U22923 (N_22923,N_21618,N_21146);
nand U22924 (N_22924,N_21300,N_21121);
nand U22925 (N_22925,N_22207,N_21247);
or U22926 (N_22926,N_21150,N_21728);
xor U22927 (N_22927,N_21885,N_21779);
and U22928 (N_22928,N_21894,N_21899);
nand U22929 (N_22929,N_21766,N_22334);
xnor U22930 (N_22930,N_21662,N_21813);
nand U22931 (N_22931,N_21383,N_21997);
and U22932 (N_22932,N_22320,N_21354);
nand U22933 (N_22933,N_21061,N_21723);
xor U22934 (N_22934,N_21162,N_22205);
nand U22935 (N_22935,N_21756,N_21363);
nor U22936 (N_22936,N_21744,N_21498);
xor U22937 (N_22937,N_21009,N_21835);
and U22938 (N_22938,N_22085,N_21717);
nor U22939 (N_22939,N_21697,N_21073);
xor U22940 (N_22940,N_21281,N_22115);
or U22941 (N_22941,N_21366,N_21302);
or U22942 (N_22942,N_22175,N_22007);
nand U22943 (N_22943,N_21576,N_21331);
xnor U22944 (N_22944,N_21947,N_21568);
nand U22945 (N_22945,N_21483,N_21964);
or U22946 (N_22946,N_22470,N_21090);
xnor U22947 (N_22947,N_21043,N_22092);
and U22948 (N_22948,N_21987,N_22449);
or U22949 (N_22949,N_22153,N_21035);
nand U22950 (N_22950,N_21647,N_22439);
nand U22951 (N_22951,N_22155,N_22348);
xnor U22952 (N_22952,N_21306,N_21413);
nand U22953 (N_22953,N_21439,N_21681);
nand U22954 (N_22954,N_21314,N_22297);
nand U22955 (N_22955,N_22412,N_21241);
or U22956 (N_22956,N_22255,N_21861);
or U22957 (N_22957,N_22461,N_21922);
or U22958 (N_22958,N_21093,N_21007);
or U22959 (N_22959,N_21664,N_22022);
nor U22960 (N_22960,N_22287,N_21270);
nor U22961 (N_22961,N_21663,N_21732);
nand U22962 (N_22962,N_22045,N_21081);
and U22963 (N_22963,N_21709,N_21676);
nand U22964 (N_22964,N_21194,N_21680);
nor U22965 (N_22965,N_21700,N_21011);
or U22966 (N_22966,N_21907,N_21523);
and U22967 (N_22967,N_22299,N_21334);
or U22968 (N_22968,N_22496,N_22217);
xnor U22969 (N_22969,N_21212,N_21103);
and U22970 (N_22970,N_21854,N_21391);
nand U22971 (N_22971,N_21714,N_21768);
xnor U22972 (N_22972,N_22495,N_21380);
nor U22973 (N_22973,N_22219,N_21274);
xor U22974 (N_22974,N_22414,N_21989);
or U22975 (N_22975,N_21749,N_22210);
nor U22976 (N_22976,N_21368,N_21145);
xor U22977 (N_22977,N_21217,N_21600);
nand U22978 (N_22978,N_22392,N_22271);
nand U22979 (N_22979,N_21475,N_22032);
xor U22980 (N_22980,N_22222,N_21226);
nand U22981 (N_22981,N_21080,N_21229);
and U22982 (N_22982,N_21014,N_22265);
nor U22983 (N_22983,N_21704,N_21426);
nor U22984 (N_22984,N_21460,N_21436);
and U22985 (N_22985,N_21517,N_21998);
xnor U22986 (N_22986,N_22244,N_22410);
nand U22987 (N_22987,N_21582,N_22339);
nand U22988 (N_22988,N_21876,N_22001);
xnor U22989 (N_22989,N_21163,N_21476);
and U22990 (N_22990,N_21636,N_21111);
nor U22991 (N_22991,N_22379,N_21877);
nor U22992 (N_22992,N_21144,N_22211);
xnor U22993 (N_22993,N_21546,N_21791);
nor U22994 (N_22994,N_22420,N_21401);
nand U22995 (N_22995,N_22278,N_21084);
and U22996 (N_22996,N_21276,N_22017);
or U22997 (N_22997,N_21424,N_21197);
and U22998 (N_22998,N_22253,N_21116);
and U22999 (N_22999,N_21421,N_21774);
or U23000 (N_23000,N_21454,N_21656);
nand U23001 (N_23001,N_21390,N_22130);
nand U23002 (N_23002,N_21339,N_22119);
and U23003 (N_23003,N_22099,N_22466);
and U23004 (N_23004,N_22010,N_21044);
and U23005 (N_23005,N_21058,N_22114);
and U23006 (N_23006,N_22341,N_21164);
nand U23007 (N_23007,N_21500,N_21509);
nand U23008 (N_23008,N_21871,N_22353);
xor U23009 (N_23009,N_22129,N_21932);
nand U23010 (N_23010,N_22173,N_21253);
and U23011 (N_23011,N_21373,N_22467);
and U23012 (N_23012,N_21506,N_22252);
nor U23013 (N_23013,N_22387,N_21743);
xor U23014 (N_23014,N_22121,N_21820);
or U23015 (N_23015,N_22377,N_21037);
nor U23016 (N_23016,N_21881,N_21724);
nand U23017 (N_23017,N_22055,N_21615);
nand U23018 (N_23018,N_22014,N_21240);
xor U23019 (N_23019,N_21487,N_22137);
nor U23020 (N_23020,N_21538,N_21939);
xnor U23021 (N_23021,N_22005,N_22238);
and U23022 (N_23022,N_21978,N_21527);
xnor U23023 (N_23023,N_22378,N_21186);
and U23024 (N_23024,N_21437,N_21004);
and U23025 (N_23025,N_21134,N_21696);
or U23026 (N_23026,N_22159,N_21507);
xnor U23027 (N_23027,N_21062,N_21921);
nor U23028 (N_23028,N_22316,N_21898);
or U23029 (N_23029,N_21297,N_21554);
xnor U23030 (N_23030,N_22227,N_22256);
nand U23031 (N_23031,N_22381,N_21447);
nor U23032 (N_23032,N_21361,N_21638);
and U23033 (N_23033,N_21596,N_22154);
xnor U23034 (N_23034,N_21122,N_21526);
or U23035 (N_23035,N_21960,N_21155);
and U23036 (N_23036,N_21109,N_21478);
or U23037 (N_23037,N_21393,N_22193);
or U23038 (N_23038,N_21201,N_21213);
xnor U23039 (N_23039,N_21920,N_22091);
or U23040 (N_23040,N_21387,N_22456);
and U23041 (N_23041,N_22212,N_21171);
xor U23042 (N_23042,N_21106,N_21787);
nand U23043 (N_23043,N_21097,N_21187);
nand U23044 (N_23044,N_22140,N_22460);
and U23045 (N_23045,N_21778,N_21833);
nand U23046 (N_23046,N_21098,N_22402);
xnor U23047 (N_23047,N_21633,N_22125);
nor U23048 (N_23048,N_21267,N_22054);
nand U23049 (N_23049,N_21147,N_22398);
or U23050 (N_23050,N_22073,N_22049);
nand U23051 (N_23051,N_21776,N_21761);
and U23052 (N_23052,N_22325,N_21516);
nor U23053 (N_23053,N_22187,N_22288);
and U23054 (N_23054,N_21470,N_21606);
or U23055 (N_23055,N_21053,N_22061);
nand U23056 (N_23056,N_21034,N_21372);
xor U23057 (N_23057,N_21693,N_21889);
nor U23058 (N_23058,N_22285,N_21748);
or U23059 (N_23059,N_21607,N_21903);
or U23060 (N_23060,N_21442,N_22396);
and U23061 (N_23061,N_22162,N_22333);
nand U23062 (N_23062,N_21296,N_21856);
and U23063 (N_23063,N_21702,N_21355);
or U23064 (N_23064,N_22328,N_22088);
nor U23065 (N_23065,N_21682,N_21867);
nor U23066 (N_23066,N_22199,N_22403);
nand U23067 (N_23067,N_22016,N_22358);
or U23068 (N_23068,N_22081,N_21298);
nor U23069 (N_23069,N_22498,N_22453);
nor U23070 (N_23070,N_21811,N_21286);
xnor U23071 (N_23071,N_22215,N_22245);
and U23072 (N_23072,N_21486,N_21629);
and U23073 (N_23073,N_22423,N_21860);
nor U23074 (N_23074,N_22426,N_22473);
xnor U23075 (N_23075,N_21556,N_22102);
or U23076 (N_23076,N_21694,N_21409);
xor U23077 (N_23077,N_21853,N_22068);
nand U23078 (N_23078,N_22145,N_22096);
or U23079 (N_23079,N_21752,N_21966);
or U23080 (N_23080,N_21337,N_21066);
or U23081 (N_23081,N_22429,N_21400);
or U23082 (N_23082,N_22131,N_22077);
and U23083 (N_23083,N_21614,N_21328);
nor U23084 (N_23084,N_22019,N_21301);
nor U23085 (N_23085,N_22444,N_21563);
or U23086 (N_23086,N_22259,N_22273);
or U23087 (N_23087,N_22157,N_21603);
nand U23088 (N_23088,N_22409,N_21057);
nand U23089 (N_23089,N_21706,N_21002);
or U23090 (N_23090,N_22172,N_21951);
nand U23091 (N_23091,N_21223,N_21110);
or U23092 (N_23092,N_21371,N_22476);
and U23093 (N_23093,N_21505,N_21734);
xnor U23094 (N_23094,N_21896,N_22431);
or U23095 (N_23095,N_21429,N_22223);
xnor U23096 (N_23096,N_21140,N_22303);
nand U23097 (N_23097,N_22170,N_21637);
nand U23098 (N_23098,N_21918,N_22237);
xnor U23099 (N_23099,N_21130,N_21156);
nand U23100 (N_23100,N_22249,N_22345);
nand U23101 (N_23101,N_22028,N_21581);
xor U23102 (N_23102,N_21800,N_22056);
nand U23103 (N_23103,N_21019,N_21228);
xnor U23104 (N_23104,N_21425,N_21168);
nand U23105 (N_23105,N_21246,N_21677);
or U23106 (N_23106,N_21758,N_21045);
nand U23107 (N_23107,N_21654,N_22395);
nand U23108 (N_23108,N_21594,N_21127);
nand U23109 (N_23109,N_21020,N_21104);
xnor U23110 (N_23110,N_21132,N_21325);
nor U23111 (N_23111,N_21138,N_21841);
and U23112 (N_23112,N_22228,N_21198);
nand U23113 (N_23113,N_21495,N_21251);
nor U23114 (N_23114,N_21716,N_21353);
nand U23115 (N_23115,N_21673,N_22164);
or U23116 (N_23116,N_21959,N_21536);
nor U23117 (N_23117,N_21575,N_21209);
or U23118 (N_23118,N_21079,N_21552);
nor U23119 (N_23119,N_21153,N_21626);
or U23120 (N_23120,N_21994,N_22342);
or U23121 (N_23121,N_21091,N_22184);
nand U23122 (N_23122,N_21608,N_21571);
nor U23123 (N_23123,N_22033,N_22250);
and U23124 (N_23124,N_22338,N_21979);
nor U23125 (N_23125,N_21936,N_22203);
nor U23126 (N_23126,N_21825,N_22000);
xor U23127 (N_23127,N_22309,N_21052);
and U23128 (N_23128,N_21642,N_21289);
nand U23129 (N_23129,N_21072,N_22076);
and U23130 (N_23130,N_21970,N_22401);
nor U23131 (N_23131,N_22183,N_21904);
and U23132 (N_23132,N_22235,N_22242);
and U23133 (N_23133,N_21829,N_21474);
xnor U23134 (N_23134,N_21990,N_21971);
or U23135 (N_23135,N_21513,N_21591);
xnor U23136 (N_23136,N_22315,N_21271);
xor U23137 (N_23137,N_21879,N_21481);
nor U23138 (N_23138,N_21349,N_22037);
and U23139 (N_23139,N_21258,N_22300);
nor U23140 (N_23140,N_21963,N_22349);
nand U23141 (N_23141,N_22481,N_22404);
xnor U23142 (N_23142,N_21910,N_22452);
or U23143 (N_23143,N_21377,N_22030);
or U23144 (N_23144,N_22179,N_21428);
nor U23145 (N_23145,N_21721,N_21137);
or U23146 (N_23146,N_21727,N_21416);
nand U23147 (N_23147,N_21977,N_22337);
xnor U23148 (N_23148,N_21911,N_21890);
xor U23149 (N_23149,N_21412,N_21105);
xnor U23150 (N_23150,N_22313,N_22180);
nand U23151 (N_23151,N_21117,N_21863);
nor U23152 (N_23152,N_22012,N_22009);
nor U23153 (N_23153,N_21788,N_21322);
xnor U23154 (N_23154,N_22226,N_21665);
nor U23155 (N_23155,N_22051,N_21206);
nand U23156 (N_23156,N_21705,N_21574);
and U23157 (N_23157,N_21688,N_21239);
or U23158 (N_23158,N_22459,N_21545);
nor U23159 (N_23159,N_21316,N_21082);
or U23160 (N_23160,N_21356,N_22277);
nor U23161 (N_23161,N_22057,N_21060);
or U23162 (N_23162,N_21077,N_21256);
or U23163 (N_23163,N_21980,N_21837);
xor U23164 (N_23164,N_22462,N_21384);
nand U23165 (N_23165,N_22133,N_22434);
nor U23166 (N_23166,N_21869,N_21746);
and U23167 (N_23167,N_21041,N_21319);
or U23168 (N_23168,N_21392,N_21100);
xnor U23169 (N_23169,N_22171,N_21181);
or U23170 (N_23170,N_21842,N_22489);
xnor U23171 (N_23171,N_21114,N_21622);
and U23172 (N_23172,N_21611,N_21320);
and U23173 (N_23173,N_21597,N_21173);
or U23174 (N_23174,N_21650,N_21678);
or U23175 (N_23175,N_21784,N_21805);
nand U23176 (N_23176,N_22132,N_21115);
xor U23177 (N_23177,N_21524,N_22060);
and U23178 (N_23178,N_21862,N_21984);
nand U23179 (N_23179,N_22411,N_22491);
nor U23180 (N_23180,N_21063,N_21902);
nand U23181 (N_23181,N_21683,N_21001);
and U23182 (N_23182,N_22307,N_21502);
nor U23183 (N_23183,N_21690,N_22425);
nand U23184 (N_23184,N_21530,N_22304);
nand U23185 (N_23185,N_22232,N_21379);
xor U23186 (N_23186,N_22082,N_22224);
nand U23187 (N_23187,N_21027,N_21639);
nor U23188 (N_23188,N_22344,N_21124);
nand U23189 (N_23189,N_21269,N_21669);
nor U23190 (N_23190,N_21675,N_21782);
and U23191 (N_23191,N_22424,N_21064);
and U23192 (N_23192,N_22239,N_21905);
or U23193 (N_23193,N_21242,N_22372);
xnor U23194 (N_23194,N_22065,N_21722);
xnor U23195 (N_23195,N_22369,N_22376);
or U23196 (N_23196,N_21578,N_21188);
or U23197 (N_23197,N_21230,N_21823);
or U23198 (N_23198,N_21149,N_22388);
xor U23199 (N_23199,N_21599,N_21796);
nor U23200 (N_23200,N_21237,N_21644);
or U23201 (N_23201,N_22484,N_21013);
and U23202 (N_23202,N_21418,N_21598);
nor U23203 (N_23203,N_21463,N_22380);
nor U23204 (N_23204,N_21333,N_22110);
nand U23205 (N_23205,N_22089,N_21190);
nand U23206 (N_23206,N_21395,N_21940);
nor U23207 (N_23207,N_22373,N_22188);
nor U23208 (N_23208,N_22192,N_22067);
or U23209 (N_23209,N_21969,N_21464);
and U23210 (N_23210,N_22382,N_21736);
nor U23211 (N_23211,N_21849,N_22190);
nand U23212 (N_23212,N_22002,N_21952);
nand U23213 (N_23213,N_21018,N_22268);
and U23214 (N_23214,N_21346,N_22149);
nor U23215 (N_23215,N_21803,N_22241);
xnor U23216 (N_23216,N_22266,N_21365);
and U23217 (N_23217,N_21832,N_22282);
nor U23218 (N_23218,N_22343,N_22151);
nand U23219 (N_23219,N_22418,N_21046);
xnor U23220 (N_23220,N_22254,N_21382);
xor U23221 (N_23221,N_22006,N_22118);
and U23222 (N_23222,N_21845,N_21493);
nor U23223 (N_23223,N_21279,N_22286);
xor U23224 (N_23224,N_21809,N_21520);
or U23225 (N_23225,N_22261,N_21402);
or U23226 (N_23226,N_21499,N_22202);
nand U23227 (N_23227,N_21161,N_21291);
xor U23228 (N_23228,N_21221,N_21152);
xor U23229 (N_23229,N_21679,N_21799);
or U23230 (N_23230,N_21169,N_22436);
xnor U23231 (N_23231,N_21244,N_21686);
nor U23232 (N_23232,N_21658,N_22063);
or U23233 (N_23233,N_21016,N_21078);
nand U23234 (N_23234,N_21342,N_21315);
nor U23235 (N_23235,N_21154,N_21595);
nand U23236 (N_23236,N_21227,N_21283);
nand U23237 (N_23237,N_21135,N_22196);
and U23238 (N_23238,N_21388,N_21666);
and U23239 (N_23239,N_21398,N_21583);
xnor U23240 (N_23240,N_21544,N_21707);
nor U23241 (N_23241,N_21646,N_21056);
or U23242 (N_23242,N_21336,N_21840);
nor U23243 (N_23243,N_21771,N_21729);
nor U23244 (N_23244,N_21307,N_22039);
nand U23245 (N_23245,N_21208,N_22361);
xor U23246 (N_23246,N_22375,N_21311);
xnor U23247 (N_23247,N_21176,N_21624);
or U23248 (N_23248,N_21541,N_21950);
and U23249 (N_23249,N_21792,N_22036);
xor U23250 (N_23250,N_21939,N_22460);
nand U23251 (N_23251,N_21890,N_21336);
xor U23252 (N_23252,N_21647,N_21299);
nor U23253 (N_23253,N_21306,N_21844);
nor U23254 (N_23254,N_21648,N_21178);
or U23255 (N_23255,N_21385,N_22271);
nand U23256 (N_23256,N_21224,N_21866);
or U23257 (N_23257,N_22130,N_21565);
nand U23258 (N_23258,N_22234,N_22440);
xor U23259 (N_23259,N_21177,N_21297);
xor U23260 (N_23260,N_21801,N_22410);
nand U23261 (N_23261,N_21182,N_21282);
xnor U23262 (N_23262,N_21845,N_21537);
and U23263 (N_23263,N_21995,N_21361);
nand U23264 (N_23264,N_21543,N_21746);
xnor U23265 (N_23265,N_21057,N_22144);
xor U23266 (N_23266,N_21118,N_21438);
nand U23267 (N_23267,N_21188,N_21891);
or U23268 (N_23268,N_21622,N_21644);
and U23269 (N_23269,N_22270,N_21761);
or U23270 (N_23270,N_21682,N_22369);
and U23271 (N_23271,N_21179,N_21340);
or U23272 (N_23272,N_22279,N_21898);
xor U23273 (N_23273,N_21214,N_21621);
nand U23274 (N_23274,N_21931,N_21222);
and U23275 (N_23275,N_21381,N_22465);
nand U23276 (N_23276,N_21390,N_21980);
nand U23277 (N_23277,N_21228,N_21048);
nand U23278 (N_23278,N_21853,N_21653);
xor U23279 (N_23279,N_22001,N_22445);
nand U23280 (N_23280,N_21876,N_22020);
and U23281 (N_23281,N_21968,N_21253);
and U23282 (N_23282,N_22447,N_21132);
and U23283 (N_23283,N_22043,N_21451);
nand U23284 (N_23284,N_21316,N_22431);
or U23285 (N_23285,N_21461,N_21538);
nand U23286 (N_23286,N_22227,N_21563);
and U23287 (N_23287,N_21037,N_21169);
xor U23288 (N_23288,N_21724,N_21492);
and U23289 (N_23289,N_21823,N_21831);
xor U23290 (N_23290,N_21024,N_22114);
or U23291 (N_23291,N_22350,N_21264);
nand U23292 (N_23292,N_21976,N_21588);
nor U23293 (N_23293,N_21120,N_22109);
or U23294 (N_23294,N_21777,N_21893);
xor U23295 (N_23295,N_22221,N_21144);
or U23296 (N_23296,N_21524,N_22213);
nor U23297 (N_23297,N_21558,N_21137);
and U23298 (N_23298,N_21238,N_22229);
nor U23299 (N_23299,N_22308,N_21955);
nor U23300 (N_23300,N_22472,N_22056);
and U23301 (N_23301,N_21161,N_21367);
and U23302 (N_23302,N_21494,N_21412);
nand U23303 (N_23303,N_21345,N_21013);
and U23304 (N_23304,N_22198,N_22406);
or U23305 (N_23305,N_21433,N_22343);
nor U23306 (N_23306,N_21120,N_22411);
nand U23307 (N_23307,N_22065,N_21164);
nand U23308 (N_23308,N_22054,N_21495);
and U23309 (N_23309,N_22406,N_21196);
and U23310 (N_23310,N_21649,N_22473);
nor U23311 (N_23311,N_21362,N_22106);
xor U23312 (N_23312,N_21441,N_21074);
xnor U23313 (N_23313,N_21200,N_21483);
nand U23314 (N_23314,N_21438,N_22316);
xnor U23315 (N_23315,N_22326,N_22029);
xnor U23316 (N_23316,N_21208,N_22067);
nand U23317 (N_23317,N_21590,N_21557);
and U23318 (N_23318,N_22099,N_21509);
and U23319 (N_23319,N_21802,N_21231);
xnor U23320 (N_23320,N_21834,N_21692);
nand U23321 (N_23321,N_22436,N_22040);
xnor U23322 (N_23322,N_22042,N_21919);
and U23323 (N_23323,N_21597,N_21850);
and U23324 (N_23324,N_21400,N_22176);
nor U23325 (N_23325,N_21907,N_22450);
nand U23326 (N_23326,N_21696,N_21446);
or U23327 (N_23327,N_21578,N_21379);
and U23328 (N_23328,N_21648,N_21839);
nand U23329 (N_23329,N_22064,N_21045);
and U23330 (N_23330,N_21406,N_21404);
nand U23331 (N_23331,N_21809,N_22297);
xor U23332 (N_23332,N_21741,N_21248);
nor U23333 (N_23333,N_21594,N_21894);
nor U23334 (N_23334,N_22106,N_21412);
xnor U23335 (N_23335,N_21488,N_21946);
and U23336 (N_23336,N_21504,N_22432);
or U23337 (N_23337,N_21132,N_21533);
or U23338 (N_23338,N_21258,N_22388);
and U23339 (N_23339,N_21873,N_22034);
nor U23340 (N_23340,N_22354,N_21112);
nand U23341 (N_23341,N_21606,N_22460);
or U23342 (N_23342,N_21845,N_21422);
nand U23343 (N_23343,N_21944,N_21711);
nand U23344 (N_23344,N_22218,N_22355);
and U23345 (N_23345,N_21459,N_21817);
or U23346 (N_23346,N_21428,N_21895);
xor U23347 (N_23347,N_22056,N_21281);
nand U23348 (N_23348,N_21944,N_21447);
nand U23349 (N_23349,N_21913,N_21866);
nand U23350 (N_23350,N_21179,N_21166);
nand U23351 (N_23351,N_21597,N_22160);
nor U23352 (N_23352,N_22311,N_22286);
nor U23353 (N_23353,N_21072,N_22257);
or U23354 (N_23354,N_21122,N_22184);
xor U23355 (N_23355,N_22096,N_21836);
nor U23356 (N_23356,N_21563,N_21940);
nand U23357 (N_23357,N_21886,N_21493);
or U23358 (N_23358,N_21296,N_21559);
nor U23359 (N_23359,N_22260,N_21086);
nor U23360 (N_23360,N_22015,N_21597);
or U23361 (N_23361,N_22278,N_21478);
nor U23362 (N_23362,N_21113,N_21521);
or U23363 (N_23363,N_21134,N_21011);
xnor U23364 (N_23364,N_21710,N_21013);
nor U23365 (N_23365,N_21965,N_22279);
nor U23366 (N_23366,N_21396,N_21486);
and U23367 (N_23367,N_21446,N_22253);
nor U23368 (N_23368,N_21861,N_21812);
nor U23369 (N_23369,N_22450,N_21355);
or U23370 (N_23370,N_21831,N_21904);
nor U23371 (N_23371,N_21806,N_21323);
or U23372 (N_23372,N_22177,N_21582);
nand U23373 (N_23373,N_21839,N_21694);
nand U23374 (N_23374,N_21429,N_21489);
xor U23375 (N_23375,N_21801,N_21776);
and U23376 (N_23376,N_21763,N_21768);
or U23377 (N_23377,N_21101,N_22338);
and U23378 (N_23378,N_22051,N_21213);
or U23379 (N_23379,N_22064,N_22114);
nand U23380 (N_23380,N_21698,N_21916);
or U23381 (N_23381,N_21787,N_21294);
and U23382 (N_23382,N_21091,N_21215);
xor U23383 (N_23383,N_21160,N_21965);
and U23384 (N_23384,N_21003,N_21233);
nand U23385 (N_23385,N_21943,N_21317);
nor U23386 (N_23386,N_21487,N_21431);
or U23387 (N_23387,N_21609,N_21185);
and U23388 (N_23388,N_21508,N_22407);
nor U23389 (N_23389,N_22068,N_21778);
nand U23390 (N_23390,N_21588,N_21178);
xnor U23391 (N_23391,N_21732,N_21206);
nand U23392 (N_23392,N_22334,N_21787);
xnor U23393 (N_23393,N_21420,N_22494);
nand U23394 (N_23394,N_21195,N_21878);
xor U23395 (N_23395,N_21157,N_21231);
xor U23396 (N_23396,N_22333,N_21732);
nand U23397 (N_23397,N_21394,N_21702);
nor U23398 (N_23398,N_21322,N_21235);
nand U23399 (N_23399,N_21510,N_21576);
nand U23400 (N_23400,N_21447,N_21170);
nand U23401 (N_23401,N_21936,N_21392);
nor U23402 (N_23402,N_21005,N_21404);
or U23403 (N_23403,N_21191,N_21054);
nand U23404 (N_23404,N_21263,N_21050);
or U23405 (N_23405,N_21087,N_21314);
nand U23406 (N_23406,N_21225,N_21050);
nand U23407 (N_23407,N_21445,N_21393);
and U23408 (N_23408,N_21500,N_21347);
xnor U23409 (N_23409,N_22393,N_22458);
nand U23410 (N_23410,N_21368,N_22083);
nand U23411 (N_23411,N_22234,N_22401);
xnor U23412 (N_23412,N_21387,N_22299);
xor U23413 (N_23413,N_21597,N_22471);
or U23414 (N_23414,N_21202,N_22042);
and U23415 (N_23415,N_22137,N_22189);
nand U23416 (N_23416,N_21457,N_22442);
nand U23417 (N_23417,N_21614,N_21011);
nor U23418 (N_23418,N_21910,N_21847);
xor U23419 (N_23419,N_21739,N_22350);
and U23420 (N_23420,N_22143,N_21703);
and U23421 (N_23421,N_21282,N_22366);
or U23422 (N_23422,N_21121,N_22287);
or U23423 (N_23423,N_21525,N_21981);
nand U23424 (N_23424,N_21557,N_21735);
xor U23425 (N_23425,N_21320,N_22376);
and U23426 (N_23426,N_22409,N_21817);
or U23427 (N_23427,N_21609,N_21647);
nor U23428 (N_23428,N_21120,N_22175);
nand U23429 (N_23429,N_22089,N_21560);
nor U23430 (N_23430,N_21670,N_22481);
xor U23431 (N_23431,N_21544,N_22364);
xor U23432 (N_23432,N_21465,N_22484);
nand U23433 (N_23433,N_21197,N_22024);
and U23434 (N_23434,N_22190,N_22057);
nor U23435 (N_23435,N_21732,N_22398);
or U23436 (N_23436,N_21590,N_21862);
nor U23437 (N_23437,N_21420,N_22157);
nand U23438 (N_23438,N_21940,N_22008);
and U23439 (N_23439,N_21882,N_21348);
xor U23440 (N_23440,N_21006,N_21455);
or U23441 (N_23441,N_21638,N_21406);
or U23442 (N_23442,N_21835,N_22203);
xor U23443 (N_23443,N_21114,N_22481);
and U23444 (N_23444,N_21813,N_21370);
xnor U23445 (N_23445,N_22299,N_22183);
and U23446 (N_23446,N_22304,N_21992);
nand U23447 (N_23447,N_21914,N_21995);
or U23448 (N_23448,N_22379,N_22212);
or U23449 (N_23449,N_22291,N_22250);
or U23450 (N_23450,N_21370,N_21064);
nand U23451 (N_23451,N_21495,N_22430);
xnor U23452 (N_23452,N_21230,N_22353);
nand U23453 (N_23453,N_21453,N_21047);
xor U23454 (N_23454,N_21797,N_22336);
and U23455 (N_23455,N_21359,N_22085);
xnor U23456 (N_23456,N_21100,N_21628);
xnor U23457 (N_23457,N_21838,N_21021);
nand U23458 (N_23458,N_21869,N_21457);
or U23459 (N_23459,N_21855,N_21716);
xor U23460 (N_23460,N_21819,N_21525);
xnor U23461 (N_23461,N_21915,N_21963);
or U23462 (N_23462,N_21342,N_22383);
xor U23463 (N_23463,N_21775,N_21065);
nor U23464 (N_23464,N_21815,N_21929);
nand U23465 (N_23465,N_21446,N_21694);
nand U23466 (N_23466,N_21888,N_22081);
xor U23467 (N_23467,N_21683,N_21872);
nand U23468 (N_23468,N_21056,N_21885);
xnor U23469 (N_23469,N_21756,N_22439);
and U23470 (N_23470,N_21464,N_21333);
xor U23471 (N_23471,N_21644,N_22002);
xnor U23472 (N_23472,N_22139,N_21809);
and U23473 (N_23473,N_21693,N_22314);
nand U23474 (N_23474,N_21390,N_21833);
nor U23475 (N_23475,N_22395,N_21593);
xor U23476 (N_23476,N_21901,N_22177);
or U23477 (N_23477,N_21107,N_22265);
nand U23478 (N_23478,N_21659,N_22464);
nor U23479 (N_23479,N_21114,N_21409);
xnor U23480 (N_23480,N_21797,N_21199);
xor U23481 (N_23481,N_21788,N_21699);
nand U23482 (N_23482,N_22386,N_21043);
and U23483 (N_23483,N_21368,N_21802);
and U23484 (N_23484,N_21403,N_21117);
xnor U23485 (N_23485,N_21064,N_21523);
xor U23486 (N_23486,N_21103,N_21732);
nor U23487 (N_23487,N_21270,N_21112);
or U23488 (N_23488,N_21119,N_22283);
xor U23489 (N_23489,N_22129,N_22306);
nor U23490 (N_23490,N_22054,N_21505);
nor U23491 (N_23491,N_21808,N_21514);
and U23492 (N_23492,N_21102,N_21738);
and U23493 (N_23493,N_22356,N_21044);
nor U23494 (N_23494,N_21729,N_22017);
nand U23495 (N_23495,N_21475,N_22475);
and U23496 (N_23496,N_22262,N_22318);
or U23497 (N_23497,N_21859,N_22280);
xor U23498 (N_23498,N_21839,N_22232);
xnor U23499 (N_23499,N_21552,N_21438);
and U23500 (N_23500,N_22142,N_21330);
xor U23501 (N_23501,N_21993,N_21353);
nand U23502 (N_23502,N_21957,N_22461);
and U23503 (N_23503,N_21672,N_22037);
and U23504 (N_23504,N_21386,N_22303);
nand U23505 (N_23505,N_21679,N_21064);
or U23506 (N_23506,N_21239,N_21941);
nor U23507 (N_23507,N_21718,N_21273);
and U23508 (N_23508,N_21908,N_21184);
nand U23509 (N_23509,N_22376,N_21089);
xnor U23510 (N_23510,N_21769,N_21973);
or U23511 (N_23511,N_21832,N_21916);
and U23512 (N_23512,N_22350,N_22478);
xnor U23513 (N_23513,N_22292,N_21228);
or U23514 (N_23514,N_21760,N_21351);
and U23515 (N_23515,N_22465,N_21049);
xor U23516 (N_23516,N_21826,N_21242);
and U23517 (N_23517,N_22187,N_21230);
nor U23518 (N_23518,N_21565,N_21988);
and U23519 (N_23519,N_21309,N_22092);
and U23520 (N_23520,N_21642,N_21966);
or U23521 (N_23521,N_21781,N_22009);
nand U23522 (N_23522,N_22425,N_21129);
xor U23523 (N_23523,N_21444,N_21582);
xor U23524 (N_23524,N_21805,N_21138);
xnor U23525 (N_23525,N_21004,N_22379);
xor U23526 (N_23526,N_21970,N_22414);
nand U23527 (N_23527,N_21046,N_21174);
and U23528 (N_23528,N_22138,N_21249);
nor U23529 (N_23529,N_21398,N_21944);
nand U23530 (N_23530,N_22244,N_22396);
nand U23531 (N_23531,N_22077,N_21502);
xnor U23532 (N_23532,N_21619,N_21221);
and U23533 (N_23533,N_22096,N_21527);
nand U23534 (N_23534,N_22318,N_21661);
nor U23535 (N_23535,N_21553,N_22189);
and U23536 (N_23536,N_21674,N_22091);
and U23537 (N_23537,N_22012,N_22251);
xor U23538 (N_23538,N_21359,N_21937);
and U23539 (N_23539,N_22453,N_22144);
and U23540 (N_23540,N_21410,N_22015);
nor U23541 (N_23541,N_21457,N_21152);
or U23542 (N_23542,N_21099,N_21033);
or U23543 (N_23543,N_21193,N_21796);
and U23544 (N_23544,N_22081,N_21742);
xnor U23545 (N_23545,N_22156,N_21839);
nor U23546 (N_23546,N_21681,N_21708);
nor U23547 (N_23547,N_22146,N_22138);
and U23548 (N_23548,N_21492,N_21903);
xnor U23549 (N_23549,N_21759,N_21167);
or U23550 (N_23550,N_21353,N_21479);
nor U23551 (N_23551,N_21412,N_22093);
nor U23552 (N_23552,N_21322,N_21849);
and U23553 (N_23553,N_21341,N_21118);
or U23554 (N_23554,N_21380,N_21438);
xnor U23555 (N_23555,N_22278,N_22109);
xor U23556 (N_23556,N_21683,N_21023);
nor U23557 (N_23557,N_21936,N_22306);
and U23558 (N_23558,N_21846,N_21837);
nor U23559 (N_23559,N_22297,N_21791);
nor U23560 (N_23560,N_22053,N_21002);
nor U23561 (N_23561,N_22199,N_21413);
xor U23562 (N_23562,N_21178,N_22255);
nand U23563 (N_23563,N_22231,N_21314);
nor U23564 (N_23564,N_22156,N_21064);
or U23565 (N_23565,N_21266,N_22286);
and U23566 (N_23566,N_21518,N_22073);
or U23567 (N_23567,N_22261,N_21154);
and U23568 (N_23568,N_21246,N_21174);
xor U23569 (N_23569,N_21598,N_22394);
nor U23570 (N_23570,N_21303,N_21720);
xor U23571 (N_23571,N_21009,N_21354);
nand U23572 (N_23572,N_21286,N_21787);
nand U23573 (N_23573,N_22029,N_22191);
nor U23574 (N_23574,N_21648,N_21751);
and U23575 (N_23575,N_21030,N_21715);
nor U23576 (N_23576,N_22078,N_21615);
or U23577 (N_23577,N_21842,N_21740);
or U23578 (N_23578,N_22377,N_21318);
and U23579 (N_23579,N_21362,N_21117);
or U23580 (N_23580,N_21201,N_21512);
nor U23581 (N_23581,N_21730,N_22225);
and U23582 (N_23582,N_22486,N_21141);
and U23583 (N_23583,N_22001,N_21729);
nand U23584 (N_23584,N_21801,N_21632);
nand U23585 (N_23585,N_21569,N_22289);
or U23586 (N_23586,N_21002,N_21176);
xnor U23587 (N_23587,N_22277,N_22438);
xor U23588 (N_23588,N_22273,N_22018);
and U23589 (N_23589,N_21286,N_21221);
and U23590 (N_23590,N_21562,N_21004);
or U23591 (N_23591,N_21031,N_21150);
nand U23592 (N_23592,N_21473,N_21939);
nand U23593 (N_23593,N_22316,N_21079);
and U23594 (N_23594,N_22195,N_21519);
and U23595 (N_23595,N_22153,N_21994);
nand U23596 (N_23596,N_22083,N_21158);
nand U23597 (N_23597,N_21795,N_22497);
nor U23598 (N_23598,N_22364,N_21541);
and U23599 (N_23599,N_21920,N_21969);
nor U23600 (N_23600,N_21997,N_21887);
nand U23601 (N_23601,N_22493,N_22294);
and U23602 (N_23602,N_21809,N_22342);
or U23603 (N_23603,N_22355,N_21041);
and U23604 (N_23604,N_22211,N_21974);
xnor U23605 (N_23605,N_21715,N_22403);
or U23606 (N_23606,N_22395,N_22412);
nor U23607 (N_23607,N_21483,N_21695);
xnor U23608 (N_23608,N_21170,N_21174);
nor U23609 (N_23609,N_21847,N_22272);
nand U23610 (N_23610,N_22165,N_21642);
and U23611 (N_23611,N_22156,N_22323);
or U23612 (N_23612,N_22063,N_21663);
nand U23613 (N_23613,N_21169,N_21088);
nor U23614 (N_23614,N_21511,N_21175);
or U23615 (N_23615,N_21063,N_21116);
nor U23616 (N_23616,N_21503,N_22290);
and U23617 (N_23617,N_21116,N_21972);
and U23618 (N_23618,N_22269,N_21384);
or U23619 (N_23619,N_22211,N_21321);
or U23620 (N_23620,N_22385,N_21086);
or U23621 (N_23621,N_22435,N_21548);
xnor U23622 (N_23622,N_21572,N_21532);
nor U23623 (N_23623,N_21292,N_21363);
or U23624 (N_23624,N_21786,N_22278);
nor U23625 (N_23625,N_21860,N_21406);
or U23626 (N_23626,N_21006,N_21447);
nor U23627 (N_23627,N_22041,N_22160);
nand U23628 (N_23628,N_22161,N_21958);
and U23629 (N_23629,N_21822,N_21151);
nand U23630 (N_23630,N_22276,N_21121);
and U23631 (N_23631,N_22031,N_21367);
xnor U23632 (N_23632,N_22229,N_21736);
xnor U23633 (N_23633,N_21888,N_22062);
and U23634 (N_23634,N_21581,N_21688);
and U23635 (N_23635,N_21358,N_21951);
and U23636 (N_23636,N_21180,N_21511);
xnor U23637 (N_23637,N_21198,N_21833);
or U23638 (N_23638,N_21353,N_22108);
nand U23639 (N_23639,N_21138,N_21419);
nor U23640 (N_23640,N_22347,N_21550);
and U23641 (N_23641,N_21117,N_21577);
and U23642 (N_23642,N_21907,N_21432);
xnor U23643 (N_23643,N_21205,N_21398);
nand U23644 (N_23644,N_22305,N_21259);
xnor U23645 (N_23645,N_21825,N_22167);
nand U23646 (N_23646,N_21447,N_21588);
nor U23647 (N_23647,N_21167,N_22146);
xnor U23648 (N_23648,N_21664,N_21905);
or U23649 (N_23649,N_21126,N_22011);
xor U23650 (N_23650,N_22268,N_21851);
nand U23651 (N_23651,N_22013,N_21252);
or U23652 (N_23652,N_21660,N_21669);
and U23653 (N_23653,N_22383,N_21829);
nand U23654 (N_23654,N_22128,N_21259);
nor U23655 (N_23655,N_21928,N_21079);
and U23656 (N_23656,N_22366,N_22216);
or U23657 (N_23657,N_21465,N_21810);
nor U23658 (N_23658,N_21248,N_22009);
nand U23659 (N_23659,N_22070,N_21393);
or U23660 (N_23660,N_21606,N_21681);
and U23661 (N_23661,N_22080,N_22312);
nor U23662 (N_23662,N_21946,N_22219);
or U23663 (N_23663,N_22213,N_21688);
nand U23664 (N_23664,N_22172,N_22130);
xnor U23665 (N_23665,N_21015,N_21792);
or U23666 (N_23666,N_21856,N_21193);
xnor U23667 (N_23667,N_22307,N_22317);
nor U23668 (N_23668,N_21689,N_21584);
and U23669 (N_23669,N_22287,N_21745);
nand U23670 (N_23670,N_22045,N_22270);
nand U23671 (N_23671,N_21692,N_21779);
nand U23672 (N_23672,N_21180,N_21669);
nand U23673 (N_23673,N_21396,N_21950);
nor U23674 (N_23674,N_21273,N_21044);
or U23675 (N_23675,N_21925,N_22107);
nand U23676 (N_23676,N_21895,N_21785);
xnor U23677 (N_23677,N_21209,N_21386);
and U23678 (N_23678,N_21852,N_22462);
and U23679 (N_23679,N_22234,N_22331);
nand U23680 (N_23680,N_21247,N_22137);
nand U23681 (N_23681,N_21612,N_21650);
or U23682 (N_23682,N_22042,N_22422);
and U23683 (N_23683,N_21529,N_21266);
and U23684 (N_23684,N_21849,N_22265);
or U23685 (N_23685,N_21380,N_21070);
nor U23686 (N_23686,N_21162,N_21658);
nand U23687 (N_23687,N_21749,N_21941);
or U23688 (N_23688,N_21365,N_22062);
and U23689 (N_23689,N_22118,N_21740);
and U23690 (N_23690,N_21365,N_22176);
nand U23691 (N_23691,N_22345,N_21028);
nand U23692 (N_23692,N_22201,N_21314);
nor U23693 (N_23693,N_21823,N_21010);
nor U23694 (N_23694,N_21754,N_21030);
or U23695 (N_23695,N_22293,N_22397);
xnor U23696 (N_23696,N_21531,N_22144);
or U23697 (N_23697,N_21862,N_21093);
nor U23698 (N_23698,N_22362,N_21968);
xnor U23699 (N_23699,N_22270,N_21647);
and U23700 (N_23700,N_21932,N_22476);
and U23701 (N_23701,N_21307,N_21895);
nor U23702 (N_23702,N_21012,N_21950);
nor U23703 (N_23703,N_21623,N_22296);
nand U23704 (N_23704,N_22473,N_22381);
or U23705 (N_23705,N_21823,N_21768);
nor U23706 (N_23706,N_21128,N_21858);
xnor U23707 (N_23707,N_22381,N_22218);
or U23708 (N_23708,N_21833,N_22082);
and U23709 (N_23709,N_22078,N_21014);
nand U23710 (N_23710,N_21589,N_21171);
and U23711 (N_23711,N_21443,N_22167);
or U23712 (N_23712,N_21397,N_21150);
xor U23713 (N_23713,N_21832,N_21920);
nor U23714 (N_23714,N_21020,N_22223);
or U23715 (N_23715,N_21878,N_21811);
nor U23716 (N_23716,N_21279,N_22445);
and U23717 (N_23717,N_21544,N_22102);
or U23718 (N_23718,N_21862,N_22272);
or U23719 (N_23719,N_21677,N_21141);
nand U23720 (N_23720,N_21767,N_21519);
or U23721 (N_23721,N_21115,N_22020);
and U23722 (N_23722,N_21724,N_21114);
xor U23723 (N_23723,N_21248,N_21286);
nand U23724 (N_23724,N_22264,N_21573);
or U23725 (N_23725,N_21303,N_21645);
and U23726 (N_23726,N_22135,N_22277);
xnor U23727 (N_23727,N_21520,N_22030);
or U23728 (N_23728,N_22291,N_21887);
xnor U23729 (N_23729,N_22041,N_21109);
and U23730 (N_23730,N_22336,N_21663);
nand U23731 (N_23731,N_21665,N_22006);
or U23732 (N_23732,N_21448,N_21770);
nor U23733 (N_23733,N_21819,N_21735);
xnor U23734 (N_23734,N_21679,N_21542);
nor U23735 (N_23735,N_21993,N_22294);
xor U23736 (N_23736,N_21550,N_22182);
or U23737 (N_23737,N_21902,N_22194);
xnor U23738 (N_23738,N_22223,N_22252);
xor U23739 (N_23739,N_21368,N_21864);
xnor U23740 (N_23740,N_22331,N_22333);
xnor U23741 (N_23741,N_22415,N_21467);
nand U23742 (N_23742,N_22077,N_21438);
and U23743 (N_23743,N_21015,N_22377);
and U23744 (N_23744,N_21205,N_21343);
nor U23745 (N_23745,N_22109,N_21104);
and U23746 (N_23746,N_22183,N_22490);
or U23747 (N_23747,N_22159,N_21853);
xor U23748 (N_23748,N_21928,N_22227);
and U23749 (N_23749,N_21683,N_21333);
xnor U23750 (N_23750,N_21567,N_21581);
and U23751 (N_23751,N_21171,N_21425);
and U23752 (N_23752,N_21845,N_21789);
and U23753 (N_23753,N_21246,N_21787);
and U23754 (N_23754,N_21931,N_22032);
nand U23755 (N_23755,N_21367,N_21572);
and U23756 (N_23756,N_21300,N_22387);
or U23757 (N_23757,N_21154,N_22168);
or U23758 (N_23758,N_22077,N_22035);
and U23759 (N_23759,N_22315,N_21993);
and U23760 (N_23760,N_22292,N_21886);
and U23761 (N_23761,N_21896,N_21744);
or U23762 (N_23762,N_22356,N_21657);
xor U23763 (N_23763,N_21220,N_21447);
nor U23764 (N_23764,N_22452,N_21914);
nand U23765 (N_23765,N_21111,N_21704);
or U23766 (N_23766,N_22487,N_21374);
nor U23767 (N_23767,N_22245,N_21033);
xor U23768 (N_23768,N_21850,N_22006);
or U23769 (N_23769,N_22346,N_21823);
nor U23770 (N_23770,N_21748,N_22265);
and U23771 (N_23771,N_21439,N_21293);
and U23772 (N_23772,N_22059,N_22029);
and U23773 (N_23773,N_21583,N_22442);
nor U23774 (N_23774,N_21310,N_22124);
xor U23775 (N_23775,N_22078,N_21809);
and U23776 (N_23776,N_21949,N_22044);
or U23777 (N_23777,N_21730,N_22413);
and U23778 (N_23778,N_21208,N_21703);
xor U23779 (N_23779,N_21823,N_21998);
xor U23780 (N_23780,N_22177,N_21039);
nor U23781 (N_23781,N_22251,N_21685);
nand U23782 (N_23782,N_21353,N_22418);
and U23783 (N_23783,N_21226,N_21148);
and U23784 (N_23784,N_21822,N_21951);
nor U23785 (N_23785,N_21406,N_22050);
nand U23786 (N_23786,N_21674,N_21491);
nor U23787 (N_23787,N_21181,N_22485);
nand U23788 (N_23788,N_22481,N_21717);
xor U23789 (N_23789,N_21706,N_21896);
xor U23790 (N_23790,N_22367,N_21052);
nand U23791 (N_23791,N_21211,N_21795);
nand U23792 (N_23792,N_21179,N_21712);
nor U23793 (N_23793,N_21519,N_21770);
or U23794 (N_23794,N_21923,N_21329);
nand U23795 (N_23795,N_21674,N_22187);
and U23796 (N_23796,N_21546,N_22155);
or U23797 (N_23797,N_21714,N_22409);
xnor U23798 (N_23798,N_22066,N_21989);
xor U23799 (N_23799,N_21738,N_21357);
nor U23800 (N_23800,N_22297,N_22286);
nor U23801 (N_23801,N_22256,N_22245);
and U23802 (N_23802,N_21167,N_22076);
and U23803 (N_23803,N_21937,N_22264);
or U23804 (N_23804,N_22363,N_22048);
or U23805 (N_23805,N_22277,N_21120);
nand U23806 (N_23806,N_21251,N_21073);
nand U23807 (N_23807,N_21921,N_22460);
nor U23808 (N_23808,N_21360,N_21817);
nand U23809 (N_23809,N_21880,N_21968);
nor U23810 (N_23810,N_21252,N_21169);
and U23811 (N_23811,N_22299,N_21005);
xnor U23812 (N_23812,N_21459,N_22042);
xnor U23813 (N_23813,N_21453,N_22087);
nor U23814 (N_23814,N_21946,N_22091);
nand U23815 (N_23815,N_21973,N_22124);
nand U23816 (N_23816,N_22004,N_21991);
nor U23817 (N_23817,N_21730,N_21751);
or U23818 (N_23818,N_21030,N_21056);
and U23819 (N_23819,N_21758,N_22481);
nor U23820 (N_23820,N_22470,N_22384);
or U23821 (N_23821,N_21139,N_21014);
or U23822 (N_23822,N_21031,N_21780);
nand U23823 (N_23823,N_22239,N_21999);
nand U23824 (N_23824,N_21771,N_21137);
nor U23825 (N_23825,N_21261,N_21901);
nand U23826 (N_23826,N_21981,N_22386);
nand U23827 (N_23827,N_21524,N_22436);
nor U23828 (N_23828,N_22390,N_21061);
nand U23829 (N_23829,N_21334,N_22014);
or U23830 (N_23830,N_22005,N_21265);
and U23831 (N_23831,N_21331,N_22050);
nand U23832 (N_23832,N_21431,N_22171);
nand U23833 (N_23833,N_22188,N_22364);
nor U23834 (N_23834,N_21301,N_21459);
xnor U23835 (N_23835,N_21949,N_22147);
xnor U23836 (N_23836,N_21379,N_21839);
xor U23837 (N_23837,N_21112,N_22169);
nand U23838 (N_23838,N_21871,N_21413);
nor U23839 (N_23839,N_22367,N_21385);
or U23840 (N_23840,N_22322,N_21798);
or U23841 (N_23841,N_22441,N_21523);
nor U23842 (N_23842,N_21472,N_21225);
xor U23843 (N_23843,N_21777,N_22083);
nor U23844 (N_23844,N_21570,N_21464);
and U23845 (N_23845,N_21958,N_21992);
nor U23846 (N_23846,N_22424,N_21359);
xor U23847 (N_23847,N_21049,N_22423);
or U23848 (N_23848,N_21852,N_21935);
nand U23849 (N_23849,N_22071,N_21436);
nor U23850 (N_23850,N_22162,N_21741);
nor U23851 (N_23851,N_21407,N_21148);
xnor U23852 (N_23852,N_21441,N_21922);
xnor U23853 (N_23853,N_21799,N_22055);
nand U23854 (N_23854,N_21961,N_22059);
xnor U23855 (N_23855,N_22127,N_21578);
nand U23856 (N_23856,N_21065,N_21454);
or U23857 (N_23857,N_22395,N_21976);
or U23858 (N_23858,N_22073,N_21895);
or U23859 (N_23859,N_21481,N_21743);
xnor U23860 (N_23860,N_21108,N_22238);
nor U23861 (N_23861,N_21156,N_21876);
or U23862 (N_23862,N_21404,N_21275);
xnor U23863 (N_23863,N_22485,N_22005);
xor U23864 (N_23864,N_21424,N_21292);
nand U23865 (N_23865,N_22328,N_21840);
nor U23866 (N_23866,N_21934,N_21862);
nand U23867 (N_23867,N_21447,N_22233);
or U23868 (N_23868,N_21778,N_21565);
nor U23869 (N_23869,N_22181,N_21467);
nand U23870 (N_23870,N_22107,N_22365);
or U23871 (N_23871,N_21545,N_21316);
xor U23872 (N_23872,N_21033,N_21633);
nor U23873 (N_23873,N_22149,N_21655);
and U23874 (N_23874,N_21211,N_21207);
nand U23875 (N_23875,N_21792,N_22145);
xnor U23876 (N_23876,N_21948,N_21707);
and U23877 (N_23877,N_22120,N_21820);
xor U23878 (N_23878,N_21284,N_21236);
or U23879 (N_23879,N_21939,N_21222);
and U23880 (N_23880,N_21578,N_21383);
nand U23881 (N_23881,N_22039,N_21121);
nor U23882 (N_23882,N_22305,N_21907);
nor U23883 (N_23883,N_21177,N_21608);
and U23884 (N_23884,N_21905,N_22086);
xor U23885 (N_23885,N_21675,N_22198);
or U23886 (N_23886,N_21331,N_21277);
nand U23887 (N_23887,N_21506,N_22105);
nor U23888 (N_23888,N_21650,N_21086);
nor U23889 (N_23889,N_22261,N_21714);
nand U23890 (N_23890,N_21787,N_21024);
nand U23891 (N_23891,N_21601,N_21035);
nand U23892 (N_23892,N_21258,N_21611);
and U23893 (N_23893,N_21590,N_22118);
or U23894 (N_23894,N_21267,N_21728);
nor U23895 (N_23895,N_21855,N_21705);
nand U23896 (N_23896,N_22387,N_22446);
nand U23897 (N_23897,N_22465,N_21174);
nor U23898 (N_23898,N_22327,N_21018);
and U23899 (N_23899,N_21781,N_21654);
nor U23900 (N_23900,N_21183,N_22414);
nand U23901 (N_23901,N_22098,N_21188);
nor U23902 (N_23902,N_22376,N_22297);
or U23903 (N_23903,N_22299,N_21072);
nor U23904 (N_23904,N_21335,N_22313);
and U23905 (N_23905,N_21340,N_21330);
nand U23906 (N_23906,N_22348,N_22192);
xnor U23907 (N_23907,N_21470,N_21877);
xnor U23908 (N_23908,N_22260,N_21477);
xor U23909 (N_23909,N_21605,N_22394);
or U23910 (N_23910,N_22235,N_21086);
xor U23911 (N_23911,N_22127,N_21458);
or U23912 (N_23912,N_22242,N_22488);
or U23913 (N_23913,N_22275,N_21593);
xnor U23914 (N_23914,N_21316,N_21360);
and U23915 (N_23915,N_21370,N_22218);
nor U23916 (N_23916,N_21225,N_22294);
and U23917 (N_23917,N_21575,N_21750);
nand U23918 (N_23918,N_21325,N_22233);
and U23919 (N_23919,N_21855,N_21597);
xnor U23920 (N_23920,N_22199,N_22435);
xnor U23921 (N_23921,N_21934,N_21877);
nand U23922 (N_23922,N_21601,N_22183);
nor U23923 (N_23923,N_21424,N_21097);
nand U23924 (N_23924,N_22205,N_21325);
or U23925 (N_23925,N_21961,N_21705);
nor U23926 (N_23926,N_22169,N_21733);
xor U23927 (N_23927,N_21703,N_22016);
xnor U23928 (N_23928,N_21261,N_22492);
nor U23929 (N_23929,N_21000,N_22003);
or U23930 (N_23930,N_21628,N_21327);
nor U23931 (N_23931,N_21286,N_21380);
xnor U23932 (N_23932,N_21824,N_21581);
nor U23933 (N_23933,N_22121,N_21637);
and U23934 (N_23934,N_22010,N_21512);
nor U23935 (N_23935,N_21131,N_21582);
nor U23936 (N_23936,N_22389,N_21348);
xor U23937 (N_23937,N_21143,N_21431);
xnor U23938 (N_23938,N_21322,N_22231);
and U23939 (N_23939,N_21307,N_21881);
and U23940 (N_23940,N_22086,N_21440);
nor U23941 (N_23941,N_21292,N_21320);
xnor U23942 (N_23942,N_21981,N_22419);
nand U23943 (N_23943,N_21056,N_21801);
xor U23944 (N_23944,N_22483,N_21584);
or U23945 (N_23945,N_21083,N_21361);
and U23946 (N_23946,N_21858,N_21592);
or U23947 (N_23947,N_22360,N_21969);
nand U23948 (N_23948,N_21880,N_21378);
nand U23949 (N_23949,N_21567,N_21695);
nor U23950 (N_23950,N_21433,N_21434);
or U23951 (N_23951,N_21344,N_21655);
or U23952 (N_23952,N_21700,N_21974);
xnor U23953 (N_23953,N_22474,N_21418);
xnor U23954 (N_23954,N_21687,N_22178);
nand U23955 (N_23955,N_21099,N_21671);
nand U23956 (N_23956,N_21095,N_21364);
nor U23957 (N_23957,N_22442,N_21574);
nand U23958 (N_23958,N_22356,N_22323);
nand U23959 (N_23959,N_21090,N_22427);
or U23960 (N_23960,N_21143,N_22428);
or U23961 (N_23961,N_21072,N_22313);
xnor U23962 (N_23962,N_22234,N_21003);
or U23963 (N_23963,N_21873,N_21641);
nand U23964 (N_23964,N_21890,N_21947);
or U23965 (N_23965,N_22019,N_22001);
nand U23966 (N_23966,N_21137,N_21377);
nor U23967 (N_23967,N_21305,N_21942);
nor U23968 (N_23968,N_21123,N_21084);
or U23969 (N_23969,N_21559,N_21741);
or U23970 (N_23970,N_21815,N_21828);
nand U23971 (N_23971,N_21798,N_21015);
or U23972 (N_23972,N_21832,N_21572);
and U23973 (N_23973,N_21773,N_21513);
nand U23974 (N_23974,N_21301,N_22346);
nand U23975 (N_23975,N_22476,N_21937);
xor U23976 (N_23976,N_22251,N_21581);
xnor U23977 (N_23977,N_22421,N_21606);
nor U23978 (N_23978,N_21516,N_22387);
xnor U23979 (N_23979,N_21078,N_21113);
and U23980 (N_23980,N_21254,N_22057);
and U23981 (N_23981,N_21174,N_21916);
xor U23982 (N_23982,N_21732,N_21646);
nor U23983 (N_23983,N_21104,N_21113);
and U23984 (N_23984,N_22497,N_21158);
nor U23985 (N_23985,N_22145,N_21030);
or U23986 (N_23986,N_21023,N_22363);
nor U23987 (N_23987,N_21077,N_21522);
nand U23988 (N_23988,N_21994,N_21289);
xor U23989 (N_23989,N_22386,N_21424);
or U23990 (N_23990,N_21881,N_21107);
or U23991 (N_23991,N_21464,N_21584);
and U23992 (N_23992,N_22059,N_21734);
or U23993 (N_23993,N_22175,N_21508);
and U23994 (N_23994,N_21945,N_21955);
and U23995 (N_23995,N_22373,N_21716);
and U23996 (N_23996,N_21521,N_21832);
nand U23997 (N_23997,N_22324,N_21641);
xnor U23998 (N_23998,N_22229,N_22078);
and U23999 (N_23999,N_22011,N_21179);
nand U24000 (N_24000,N_23607,N_23165);
or U24001 (N_24001,N_23556,N_23678);
nor U24002 (N_24002,N_23452,N_23045);
or U24003 (N_24003,N_23094,N_22808);
nor U24004 (N_24004,N_23781,N_23601);
nand U24005 (N_24005,N_23271,N_22849);
xor U24006 (N_24006,N_23592,N_23911);
nor U24007 (N_24007,N_22714,N_22500);
or U24008 (N_24008,N_22525,N_22960);
xnor U24009 (N_24009,N_23619,N_23789);
xor U24010 (N_24010,N_23830,N_23598);
or U24011 (N_24011,N_23960,N_23267);
or U24012 (N_24012,N_23061,N_23709);
nor U24013 (N_24013,N_23160,N_23345);
and U24014 (N_24014,N_23140,N_23388);
or U24015 (N_24015,N_22939,N_22566);
nor U24016 (N_24016,N_23337,N_23643);
nand U24017 (N_24017,N_23159,N_23609);
nand U24018 (N_24018,N_23948,N_23258);
or U24019 (N_24019,N_22595,N_23145);
and U24020 (N_24020,N_23965,N_23628);
nand U24021 (N_24021,N_22619,N_22858);
xnor U24022 (N_24022,N_23172,N_22709);
xnor U24023 (N_24023,N_22701,N_23087);
nor U24024 (N_24024,N_23297,N_23921);
nand U24025 (N_24025,N_22564,N_22534);
nor U24026 (N_24026,N_22673,N_23578);
or U24027 (N_24027,N_23856,N_23176);
nor U24028 (N_24028,N_23995,N_23752);
and U24029 (N_24029,N_23180,N_22842);
xnor U24030 (N_24030,N_22519,N_23724);
and U24031 (N_24031,N_23088,N_22859);
xnor U24032 (N_24032,N_23011,N_23237);
or U24033 (N_24033,N_22834,N_23520);
xnor U24034 (N_24034,N_23116,N_23243);
nand U24035 (N_24035,N_22763,N_23440);
and U24036 (N_24036,N_23676,N_22636);
xor U24037 (N_24037,N_23875,N_23263);
xnor U24038 (N_24038,N_23371,N_23997);
or U24039 (N_24039,N_23700,N_23956);
or U24040 (N_24040,N_23408,N_23358);
or U24041 (N_24041,N_23420,N_22962);
xnor U24042 (N_24042,N_22975,N_22561);
nor U24043 (N_24043,N_22546,N_22847);
or U24044 (N_24044,N_23486,N_23222);
xnor U24045 (N_24045,N_22662,N_23025);
xnor U24046 (N_24046,N_22761,N_22514);
xnor U24047 (N_24047,N_23132,N_23500);
xnor U24048 (N_24048,N_22892,N_23369);
xor U24049 (N_24049,N_23979,N_23534);
xnor U24050 (N_24050,N_23433,N_23195);
nor U24051 (N_24051,N_23800,N_22574);
and U24052 (N_24052,N_22941,N_23078);
and U24053 (N_24053,N_23466,N_22744);
nand U24054 (N_24054,N_23108,N_23302);
xnor U24055 (N_24055,N_23234,N_22907);
nor U24056 (N_24056,N_23204,N_22584);
and U24057 (N_24057,N_23622,N_22766);
nand U24058 (N_24058,N_22789,N_23505);
nand U24059 (N_24059,N_22787,N_22646);
or U24060 (N_24060,N_23113,N_22767);
nor U24061 (N_24061,N_23317,N_23814);
xor U24062 (N_24062,N_22658,N_23014);
xnor U24063 (N_24063,N_23883,N_22924);
nor U24064 (N_24064,N_22899,N_23888);
nor U24065 (N_24065,N_22913,N_22531);
and U24066 (N_24066,N_22791,N_23522);
and U24067 (N_24067,N_23477,N_22889);
xnor U24068 (N_24068,N_23450,N_23903);
nor U24069 (N_24069,N_23121,N_22776);
xnor U24070 (N_24070,N_23435,N_23484);
or U24071 (N_24071,N_23611,N_23928);
nand U24072 (N_24072,N_23439,N_23331);
nand U24073 (N_24073,N_23646,N_22526);
and U24074 (N_24074,N_22581,N_22955);
xnor U24075 (N_24075,N_23627,N_23573);
and U24076 (N_24076,N_22737,N_22770);
or U24077 (N_24077,N_23374,N_23060);
and U24078 (N_24078,N_23654,N_23665);
xor U24079 (N_24079,N_23907,N_23315);
nor U24080 (N_24080,N_22851,N_23192);
or U24081 (N_24081,N_22857,N_23890);
and U24082 (N_24082,N_22750,N_22610);
xnor U24083 (N_24083,N_23104,N_22993);
and U24084 (N_24084,N_23436,N_23324);
xor U24085 (N_24085,N_23873,N_23931);
nand U24086 (N_24086,N_23102,N_23924);
nand U24087 (N_24087,N_23067,N_22583);
xor U24088 (N_24088,N_22586,N_23695);
xor U24089 (N_24089,N_23033,N_23207);
xnor U24090 (N_24090,N_23183,N_22832);
nand U24091 (N_24091,N_23725,N_23853);
nand U24092 (N_24092,N_22811,N_22539);
xor U24093 (N_24093,N_23095,N_23454);
and U24094 (N_24094,N_23189,N_23982);
nor U24095 (N_24095,N_22576,N_23865);
nand U24096 (N_24096,N_23815,N_23215);
nand U24097 (N_24097,N_22739,N_23082);
nor U24098 (N_24098,N_23296,N_23075);
nor U24099 (N_24099,N_23719,N_23148);
xnor U24100 (N_24100,N_22671,N_23610);
or U24101 (N_24101,N_23461,N_23984);
or U24102 (N_24102,N_22521,N_22713);
xnor U24103 (N_24103,N_23972,N_23327);
xnor U24104 (N_24104,N_23530,N_22988);
nor U24105 (N_24105,N_22677,N_22535);
or U24106 (N_24106,N_23510,N_22843);
and U24107 (N_24107,N_23981,N_23004);
or U24108 (N_24108,N_23422,N_23096);
nor U24109 (N_24109,N_23561,N_23126);
nor U24110 (N_24110,N_22800,N_23765);
or U24111 (N_24111,N_22940,N_22854);
or U24112 (N_24112,N_22772,N_23869);
xor U24113 (N_24113,N_23482,N_22505);
or U24114 (N_24114,N_23871,N_23001);
xnor U24115 (N_24115,N_23268,N_22882);
and U24116 (N_24116,N_23854,N_22589);
or U24117 (N_24117,N_23946,N_23998);
nor U24118 (N_24118,N_23012,N_23538);
and U24119 (N_24119,N_23740,N_23214);
nor U24120 (N_24120,N_23453,N_23249);
and U24121 (N_24121,N_22873,N_23872);
nand U24122 (N_24122,N_23876,N_23264);
and U24123 (N_24123,N_23567,N_23474);
or U24124 (N_24124,N_23836,N_23736);
and U24125 (N_24125,N_22792,N_23669);
nor U24126 (N_24126,N_22928,N_22659);
nand U24127 (N_24127,N_22630,N_23242);
nor U24128 (N_24128,N_22580,N_23489);
xnor U24129 (N_24129,N_23326,N_22918);
or U24130 (N_24130,N_23503,N_23506);
xor U24131 (N_24131,N_23941,N_22784);
and U24132 (N_24132,N_23687,N_23368);
nor U24133 (N_24133,N_23156,N_23109);
nand U24134 (N_24134,N_22614,N_22632);
xor U24135 (N_24135,N_23389,N_23770);
xor U24136 (N_24136,N_23127,N_22768);
xor U24137 (N_24137,N_23124,N_23198);
and U24138 (N_24138,N_23633,N_23760);
nor U24139 (N_24139,N_22694,N_23383);
xnor U24140 (N_24140,N_22528,N_23870);
nand U24141 (N_24141,N_23158,N_22641);
and U24142 (N_24142,N_22760,N_23797);
nor U24143 (N_24143,N_22951,N_23502);
and U24144 (N_24144,N_23645,N_22785);
xnor U24145 (N_24145,N_23338,N_23514);
or U24146 (N_24146,N_23634,N_22866);
and U24147 (N_24147,N_23988,N_23680);
nand U24148 (N_24148,N_22838,N_23589);
and U24149 (N_24149,N_23451,N_22805);
xnor U24150 (N_24150,N_23034,N_23714);
and U24151 (N_24151,N_22722,N_23313);
or U24152 (N_24152,N_23456,N_23166);
nand U24153 (N_24153,N_23852,N_22840);
or U24154 (N_24154,N_22991,N_23333);
nand U24155 (N_24155,N_23910,N_22769);
or U24156 (N_24156,N_22647,N_23908);
xnor U24157 (N_24157,N_23441,N_22848);
nand U24158 (N_24158,N_22700,N_22810);
nor U24159 (N_24159,N_23544,N_23959);
or U24160 (N_24160,N_22996,N_23791);
xnor U24161 (N_24161,N_22578,N_22984);
and U24162 (N_24162,N_22512,N_23220);
or U24163 (N_24163,N_22559,N_23899);
nand U24164 (N_24164,N_22781,N_23175);
and U24165 (N_24165,N_22544,N_23962);
xnor U24166 (N_24166,N_23555,N_23091);
nand U24167 (N_24167,N_23015,N_22967);
nand U24168 (N_24168,N_22634,N_23074);
and U24169 (N_24169,N_23069,N_22911);
and U24170 (N_24170,N_23518,N_22529);
or U24171 (N_24171,N_23540,N_23403);
or U24172 (N_24172,N_23100,N_23767);
or U24173 (N_24173,N_22543,N_23339);
or U24174 (N_24174,N_23392,N_23558);
nand U24175 (N_24175,N_23233,N_23901);
nand U24176 (N_24176,N_22798,N_23713);
nand U24177 (N_24177,N_23084,N_23892);
and U24178 (N_24178,N_23247,N_22891);
or U24179 (N_24179,N_23475,N_23507);
nand U24180 (N_24180,N_22821,N_22668);
xnor U24181 (N_24181,N_23275,N_23696);
xnor U24182 (N_24182,N_23837,N_23221);
nand U24183 (N_24183,N_23648,N_23462);
xor U24184 (N_24184,N_22693,N_22896);
nor U24185 (N_24185,N_22979,N_23238);
and U24186 (N_24186,N_22817,N_22856);
or U24187 (N_24187,N_23329,N_23699);
xnor U24188 (N_24188,N_22560,N_23750);
nand U24189 (N_24189,N_23787,N_23919);
xnor U24190 (N_24190,N_22683,N_23493);
nand U24191 (N_24191,N_23769,N_23318);
and U24192 (N_24192,N_22606,N_23660);
and U24193 (N_24193,N_23013,N_22601);
and U24194 (N_24194,N_22509,N_23675);
or U24195 (N_24195,N_23777,N_23656);
nand U24196 (N_24196,N_23445,N_22507);
xor U24197 (N_24197,N_23616,N_23599);
xor U24198 (N_24198,N_22549,N_23307);
or U24199 (N_24199,N_23018,N_23923);
nor U24200 (N_24200,N_22836,N_23586);
xnor U24201 (N_24201,N_23859,N_23097);
and U24202 (N_24202,N_23379,N_23753);
nand U24203 (N_24203,N_22711,N_23138);
and U24204 (N_24204,N_22537,N_23584);
xnor U24205 (N_24205,N_22890,N_23079);
nand U24206 (N_24206,N_22628,N_22973);
nor U24207 (N_24207,N_23780,N_23421);
xor U24208 (N_24208,N_22780,N_23272);
nor U24209 (N_24209,N_23808,N_23943);
nor U24210 (N_24210,N_23361,N_22689);
and U24211 (N_24211,N_23963,N_23850);
nand U24212 (N_24212,N_23277,N_23278);
nor U24213 (N_24213,N_23776,N_22845);
nor U24214 (N_24214,N_23125,N_23673);
or U24215 (N_24215,N_23036,N_23782);
nor U24216 (N_24216,N_22816,N_22598);
nand U24217 (N_24217,N_22516,N_23746);
nand U24218 (N_24218,N_22571,N_23726);
or U24219 (N_24219,N_23245,N_23716);
nand U24220 (N_24220,N_23253,N_23008);
xnor U24221 (N_24221,N_23858,N_22934);
nand U24222 (N_24222,N_23999,N_22757);
and U24223 (N_24223,N_23839,N_23527);
or U24224 (N_24224,N_23017,N_23595);
or U24225 (N_24225,N_22826,N_23975);
or U24226 (N_24226,N_22727,N_23831);
nor U24227 (N_24227,N_23691,N_23764);
nand U24228 (N_24228,N_23755,N_22977);
nor U24229 (N_24229,N_23312,N_23762);
xnor U24230 (N_24230,N_22919,N_23712);
nor U24231 (N_24231,N_23937,N_23181);
or U24232 (N_24232,N_22573,N_23194);
nand U24233 (N_24233,N_23974,N_23524);
nand U24234 (N_24234,N_23093,N_23537);
xnor U24235 (N_24235,N_22749,N_23882);
nand U24236 (N_24236,N_23038,N_23569);
or U24237 (N_24237,N_23170,N_23481);
nor U24238 (N_24238,N_23085,N_23072);
nor U24239 (N_24239,N_23838,N_23401);
xor U24240 (N_24240,N_22633,N_23142);
or U24241 (N_24241,N_22961,N_22510);
nor U24242 (N_24242,N_22865,N_23173);
nor U24243 (N_24243,N_23284,N_22720);
or U24244 (N_24244,N_22989,N_22733);
or U24245 (N_24245,N_23879,N_23218);
nor U24246 (N_24246,N_23535,N_23193);
and U24247 (N_24247,N_23940,N_22880);
and U24248 (N_24248,N_23835,N_22923);
or U24249 (N_24249,N_23874,N_22669);
nand U24250 (N_24250,N_23228,N_23229);
or U24251 (N_24251,N_22927,N_23273);
or U24252 (N_24252,N_23071,N_23040);
nand U24253 (N_24253,N_23688,N_23551);
xor U24254 (N_24254,N_22557,N_23395);
nor U24255 (N_24255,N_22912,N_23210);
xnor U24256 (N_24256,N_22685,N_23039);
xnor U24257 (N_24257,N_22864,N_23818);
or U24258 (N_24258,N_22846,N_23664);
nand U24259 (N_24259,N_23501,N_23241);
and U24260 (N_24260,N_23301,N_23343);
xnor U24261 (N_24261,N_23240,N_23355);
or U24262 (N_24262,N_23626,N_23350);
xor U24263 (N_24263,N_23064,N_22946);
nand U24264 (N_24264,N_22556,N_22547);
nor U24265 (N_24265,N_22799,N_23705);
xor U24266 (N_24266,N_23519,N_22929);
nor U24267 (N_24267,N_23196,N_23056);
nor U24268 (N_24268,N_23394,N_23260);
nand U24269 (N_24269,N_23341,N_23496);
nand U24270 (N_24270,N_23668,N_22686);
xor U24271 (N_24271,N_22697,N_22650);
nor U24272 (N_24272,N_23387,N_22540);
xnor U24273 (N_24273,N_23887,N_23734);
nor U24274 (N_24274,N_23905,N_23255);
and U24275 (N_24275,N_23840,N_23991);
or U24276 (N_24276,N_23864,N_23602);
or U24277 (N_24277,N_22932,N_23293);
nor U24278 (N_24278,N_23692,N_23157);
or U24279 (N_24279,N_23399,N_23512);
or U24280 (N_24280,N_23577,N_23944);
or U24281 (N_24281,N_22652,N_23717);
xnor U24282 (N_24282,N_23806,N_22682);
xnor U24283 (N_24283,N_22517,N_22976);
nor U24284 (N_24284,N_23969,N_23413);
nor U24285 (N_24285,N_22985,N_23063);
xnor U24286 (N_24286,N_23715,N_23495);
and U24287 (N_24287,N_22972,N_22724);
xor U24288 (N_24288,N_22883,N_23786);
xor U24289 (N_24289,N_23980,N_23532);
nand U24290 (N_24290,N_23478,N_22751);
xor U24291 (N_24291,N_23977,N_23213);
xnor U24292 (N_24292,N_23261,N_22909);
nand U24293 (N_24293,N_22860,N_22794);
and U24294 (N_24294,N_23191,N_23805);
nand U24295 (N_24295,N_23895,N_23884);
nand U24296 (N_24296,N_22582,N_22717);
and U24297 (N_24297,N_22698,N_22593);
nor U24298 (N_24298,N_23583,N_22565);
xor U24299 (N_24299,N_23428,N_22518);
and U24300 (N_24300,N_23951,N_22527);
nor U24301 (N_24301,N_22906,N_23491);
nand U24302 (N_24302,N_23322,N_22626);
xor U24303 (N_24303,N_23479,N_23135);
nor U24304 (N_24304,N_22592,N_22956);
nand U24305 (N_24305,N_23472,N_22665);
nand U24306 (N_24306,N_22833,N_22670);
nand U24307 (N_24307,N_22503,N_23902);
nor U24308 (N_24308,N_22997,N_23427);
nand U24309 (N_24309,N_23357,N_23842);
or U24310 (N_24310,N_22622,N_23226);
nor U24311 (N_24311,N_22773,N_23042);
xor U24312 (N_24312,N_23743,N_23110);
nor U24313 (N_24313,N_23576,N_23723);
nor U24314 (N_24314,N_22958,N_22532);
or U24315 (N_24315,N_23741,N_23508);
or U24316 (N_24316,N_23990,N_23370);
and U24317 (N_24317,N_23044,N_22624);
xor U24318 (N_24318,N_23605,N_23650);
xor U24319 (N_24319,N_23492,N_22831);
xnor U24320 (N_24320,N_23396,N_22520);
or U24321 (N_24321,N_23722,N_22804);
nor U24322 (N_24322,N_23244,N_23885);
nand U24323 (N_24323,N_22620,N_23287);
or U24324 (N_24324,N_22603,N_23305);
nand U24325 (N_24325,N_23163,N_23128);
or U24326 (N_24326,N_23049,N_23342);
nor U24327 (N_24327,N_22815,N_23212);
xnor U24328 (N_24328,N_23909,N_23150);
and U24329 (N_24329,N_23295,N_22705);
or U24330 (N_24330,N_23424,N_22612);
or U24331 (N_24331,N_23062,N_23847);
xnor U24332 (N_24332,N_23671,N_23702);
xnor U24333 (N_24333,N_22731,N_22548);
nand U24334 (N_24334,N_22881,N_22591);
and U24335 (N_24335,N_23168,N_23920);
and U24336 (N_24336,N_22974,N_23169);
and U24337 (N_24337,N_23103,N_23457);
and U24338 (N_24338,N_23549,N_23073);
and U24339 (N_24339,N_22953,N_23682);
nand U24340 (N_24340,N_23683,N_22830);
nor U24341 (N_24341,N_22747,N_23353);
and U24342 (N_24342,N_22806,N_23541);
or U24343 (N_24343,N_23690,N_23230);
nor U24344 (N_24344,N_23380,N_23092);
and U24345 (N_24345,N_23119,N_23531);
nand U24346 (N_24346,N_23788,N_23179);
xor U24347 (N_24347,N_23352,N_23564);
or U24348 (N_24348,N_22797,N_23086);
xnor U24349 (N_24349,N_23855,N_22600);
and U24350 (N_24350,N_23649,N_23023);
nor U24351 (N_24351,N_22947,N_22959);
and U24352 (N_24352,N_23473,N_23171);
and U24353 (N_24353,N_22638,N_23967);
nand U24354 (N_24354,N_23742,N_23807);
nor U24355 (N_24355,N_23976,N_23309);
xnor U24356 (N_24356,N_22745,N_23933);
nor U24357 (N_24357,N_23521,N_23402);
nor U24358 (N_24358,N_23798,N_23993);
nor U24359 (N_24359,N_23153,N_23662);
nand U24360 (N_24360,N_23190,N_22609);
and U24361 (N_24361,N_23199,N_23994);
xor U24362 (N_24362,N_23861,N_22627);
nor U24363 (N_24363,N_23030,N_22691);
xnor U24364 (N_24364,N_23934,N_23328);
or U24365 (N_24365,N_22986,N_22653);
nor U24366 (N_24366,N_23111,N_23711);
nand U24367 (N_24367,N_23582,N_23382);
or U24368 (N_24368,N_23224,N_23083);
and U24369 (N_24369,N_22952,N_23232);
nand U24370 (N_24370,N_22552,N_23162);
xnor U24371 (N_24371,N_23986,N_23279);
nor U24372 (N_24372,N_23351,N_23377);
and U24373 (N_24373,N_23348,N_23779);
nand U24374 (N_24374,N_23346,N_23155);
and U24375 (N_24375,N_23130,N_23659);
and U24376 (N_24376,N_23336,N_23197);
xor U24377 (N_24377,N_23672,N_23250);
and U24378 (N_24378,N_23615,N_23667);
and U24379 (N_24379,N_22734,N_23431);
nor U24380 (N_24380,N_23470,N_22596);
nand U24381 (N_24381,N_23992,N_22649);
and U24382 (N_24382,N_22703,N_23152);
and U24383 (N_24383,N_22506,N_23829);
nor U24384 (N_24384,N_22926,N_23834);
or U24385 (N_24385,N_22661,N_23332);
and U24386 (N_24386,N_23631,N_22657);
and U24387 (N_24387,N_23334,N_23335);
or U24388 (N_24388,N_22678,N_23041);
nand U24389 (N_24389,N_23310,N_22825);
nand U24390 (N_24390,N_22629,N_22684);
nor U24391 (N_24391,N_22965,N_23661);
nor U24392 (N_24392,N_23281,N_22605);
nand U24393 (N_24393,N_23409,N_22914);
nor U24394 (N_24394,N_22886,N_23529);
or U24395 (N_24395,N_22818,N_23949);
or U24396 (N_24396,N_22704,N_23131);
xor U24397 (N_24397,N_22726,N_22725);
and U24398 (N_24398,N_22895,N_23106);
and U24399 (N_24399,N_23693,N_22672);
xnor U24400 (N_24400,N_23002,N_22964);
and U24401 (N_24401,N_22504,N_22937);
or U24402 (N_24402,N_23832,N_23386);
xor U24403 (N_24403,N_22716,N_23070);
nor U24404 (N_24404,N_23099,N_22541);
and U24405 (N_24405,N_23727,N_22674);
nor U24406 (N_24406,N_23771,N_23970);
nand U24407 (N_24407,N_22654,N_23802);
and U24408 (N_24408,N_23778,N_22523);
or U24409 (N_24409,N_22692,N_23299);
nor U24410 (N_24410,N_22536,N_22998);
nor U24411 (N_24411,N_23114,N_23617);
and U24412 (N_24412,N_23446,N_22933);
nor U24413 (N_24413,N_22922,N_23423);
nor U24414 (N_24414,N_22764,N_23703);
xor U24415 (N_24415,N_23632,N_23026);
nor U24416 (N_24416,N_23323,N_23868);
nand U24417 (N_24417,N_22719,N_22680);
nand U24418 (N_24418,N_23089,N_23372);
nand U24419 (N_24419,N_22966,N_23528);
nand U24420 (N_24420,N_22908,N_23407);
nand U24421 (N_24421,N_23053,N_23543);
or U24422 (N_24422,N_23546,N_22802);
and U24423 (N_24423,N_23821,N_22795);
xnor U24424 (N_24424,N_23914,N_22796);
and U24425 (N_24425,N_22501,N_23202);
or U24426 (N_24426,N_23954,N_22994);
xnor U24427 (N_24427,N_23843,N_23397);
nor U24428 (N_24428,N_22837,N_23417);
and U24429 (N_24429,N_23294,N_23881);
or U24430 (N_24430,N_22782,N_23259);
xor U24431 (N_24431,N_22803,N_22706);
nor U24432 (N_24432,N_22900,N_22853);
and U24433 (N_24433,N_23344,N_23471);
nand U24434 (N_24434,N_23203,N_23729);
and U24435 (N_24435,N_23235,N_23846);
nand U24436 (N_24436,N_23217,N_23860);
nand U24437 (N_24437,N_22702,N_23028);
or U24438 (N_24438,N_23913,N_23927);
nor U24439 (N_24439,N_23476,N_23465);
nor U24440 (N_24440,N_22710,N_22542);
or U24441 (N_24441,N_23076,N_23112);
nor U24442 (N_24442,N_22894,N_23139);
nor U24443 (N_24443,N_22850,N_23936);
nor U24444 (N_24444,N_22572,N_23796);
nand U24445 (N_24445,N_23698,N_22824);
and U24446 (N_24446,N_22718,N_22887);
nand U24447 (N_24447,N_22651,N_23523);
and U24448 (N_24448,N_23303,N_23101);
or U24449 (N_24449,N_23205,N_22602);
nor U24450 (N_24450,N_22642,N_23657);
nand U24451 (N_24451,N_23032,N_22752);
xnor U24452 (N_24452,N_22594,N_23811);
and U24453 (N_24453,N_23708,N_23006);
or U24454 (N_24454,N_23749,N_22708);
nand U24455 (N_24455,N_23136,N_22754);
xnor U24456 (N_24456,N_23459,N_23827);
and U24457 (N_24457,N_23425,N_23046);
nor U24458 (N_24458,N_23252,N_23174);
and U24459 (N_24459,N_23460,N_22948);
xnor U24460 (N_24460,N_23587,N_23889);
nand U24461 (N_24461,N_23898,N_23239);
nand U24462 (N_24462,N_23658,N_23123);
nor U24463 (N_24463,N_22777,N_23321);
nand U24464 (N_24464,N_23251,N_22575);
nand U24465 (N_24465,N_23580,N_22730);
nand U24466 (N_24466,N_23430,N_23600);
nand U24467 (N_24467,N_22738,N_23118);
nand U24468 (N_24468,N_23005,N_22715);
xnor U24469 (N_24469,N_22625,N_23772);
xnor U24470 (N_24470,N_22511,N_23563);
xnor U24471 (N_24471,N_22978,N_23216);
nor U24472 (N_24472,N_23390,N_23904);
nand U24473 (N_24473,N_22885,N_23674);
and U24474 (N_24474,N_22839,N_23978);
nand U24475 (N_24475,N_22569,N_23973);
and U24476 (N_24476,N_22759,N_23488);
nor U24477 (N_24477,N_22758,N_23720);
or U24478 (N_24478,N_23848,N_23966);
or U24479 (N_24479,N_23122,N_23211);
or U24480 (N_24480,N_23833,N_23971);
xnor U24481 (N_24481,N_23426,N_23803);
nor U24482 (N_24482,N_23187,N_22987);
and U24483 (N_24483,N_23694,N_23637);
nand U24484 (N_24484,N_23494,N_23897);
nand U24485 (N_24485,N_22870,N_22774);
and U24486 (N_24486,N_23367,N_23306);
nand U24487 (N_24487,N_23182,N_23504);
nor U24488 (N_24488,N_22522,N_23738);
nand U24489 (N_24489,N_23756,N_22618);
or U24490 (N_24490,N_23819,N_22613);
nand U24491 (N_24491,N_23209,N_22921);
or U24492 (N_24492,N_23129,N_22587);
nand U24493 (N_24493,N_22690,N_22611);
and U24494 (N_24494,N_23432,N_23989);
and U24495 (N_24495,N_22551,N_23362);
xnor U24496 (N_24496,N_23248,N_22742);
nand U24497 (N_24497,N_23721,N_23509);
or U24498 (N_24498,N_22869,N_23449);
nand U24499 (N_24499,N_23737,N_23257);
and U24500 (N_24500,N_23363,N_23878);
nor U24501 (N_24501,N_23007,N_23571);
nand U24502 (N_24502,N_23996,N_23167);
and U24503 (N_24503,N_23133,N_23568);
and U24504 (N_24504,N_22568,N_22823);
or U24505 (N_24505,N_23670,N_23603);
nor U24506 (N_24506,N_22688,N_23464);
and U24507 (N_24507,N_23055,N_23597);
nor U24508 (N_24508,N_23283,N_22944);
nand U24509 (N_24509,N_23498,N_22878);
xnor U24510 (N_24510,N_23021,N_22778);
nor U24511 (N_24511,N_23365,N_23223);
or U24512 (N_24512,N_22712,N_22667);
xnor U24513 (N_24513,N_22513,N_23290);
and U24514 (N_24514,N_23483,N_23801);
nor U24515 (N_24515,N_22861,N_22756);
nor U24516 (N_24516,N_23047,N_23925);
and U24517 (N_24517,N_22990,N_23438);
nand U24518 (N_24518,N_23689,N_22980);
nor U24519 (N_24519,N_23866,N_23545);
and U24520 (N_24520,N_23137,N_22898);
xor U24521 (N_24521,N_23019,N_23065);
xor U24522 (N_24522,N_22786,N_23406);
nor U24523 (N_24523,N_23983,N_23706);
or U24524 (N_24524,N_22676,N_23574);
and U24525 (N_24525,N_23054,N_22852);
xor U24526 (N_24526,N_22790,N_22631);
or U24527 (N_24527,N_23285,N_22538);
xnor U24528 (N_24528,N_23236,N_22621);
nand U24529 (N_24529,N_22765,N_23641);
or U24530 (N_24530,N_22963,N_22695);
nand U24531 (N_24531,N_23647,N_23410);
nand U24532 (N_24532,N_22753,N_23024);
xor U24533 (N_24533,N_23758,N_22771);
and U24534 (N_24534,N_23912,N_23844);
xor U24535 (N_24535,N_23270,N_22707);
or U24536 (N_24536,N_22615,N_23826);
nor U24537 (N_24537,N_23490,N_23359);
xor U24538 (N_24538,N_23845,N_23059);
and U24539 (N_24539,N_22762,N_23517);
nor U24540 (N_24540,N_22735,N_23588);
or U24541 (N_24541,N_23219,N_23447);
or U24542 (N_24542,N_23414,N_23366);
nor U24543 (N_24543,N_22608,N_23434);
and U24544 (N_24544,N_23037,N_23400);
nand U24545 (N_24545,N_23164,N_23416);
nor U24546 (N_24546,N_22533,N_23655);
xor U24547 (N_24547,N_22732,N_23730);
xnor U24548 (N_24548,N_23935,N_23010);
or U24549 (N_24549,N_23896,N_23985);
xnor U24550 (N_24550,N_23677,N_22729);
nand U24551 (N_24551,N_22957,N_23795);
and U24552 (N_24552,N_23964,N_23640);
nor U24553 (N_24553,N_22874,N_23246);
or U24554 (N_24554,N_23784,N_23429);
nand U24555 (N_24555,N_22884,N_23630);
nor U24556 (N_24556,N_23566,N_22645);
and U24557 (N_24557,N_23548,N_23227);
xor U24558 (N_24558,N_23575,N_23608);
xor U24559 (N_24559,N_22558,N_23639);
nand U24560 (N_24560,N_23120,N_22644);
nor U24561 (N_24561,N_23515,N_22681);
and U24562 (N_24562,N_22935,N_23918);
nand U24563 (N_24563,N_22920,N_22954);
and U24564 (N_24564,N_23035,N_22904);
nand U24565 (N_24565,N_23300,N_23652);
nand U24566 (N_24566,N_23105,N_23644);
nand U24567 (N_24567,N_23147,N_23511);
or U24568 (N_24568,N_23141,N_23151);
and U24569 (N_24569,N_23276,N_23487);
and U24570 (N_24570,N_23554,N_22835);
xnor U24571 (N_24571,N_22801,N_23799);
or U24572 (N_24572,N_23467,N_23775);
and U24573 (N_24573,N_23448,N_22643);
or U24574 (N_24574,N_23419,N_23751);
xnor U24575 (N_24575,N_23463,N_23364);
xor U24576 (N_24576,N_23526,N_22829);
nor U24577 (N_24577,N_23590,N_23950);
xnor U24578 (N_24578,N_23718,N_23016);
or U24579 (N_24579,N_23003,N_23759);
nand U24580 (N_24580,N_22917,N_23254);
nand U24581 (N_24581,N_23381,N_23804);
xnor U24582 (N_24582,N_23384,N_23862);
xnor U24583 (N_24583,N_22550,N_22950);
xor U24584 (N_24584,N_22995,N_23812);
nor U24585 (N_24585,N_23444,N_23286);
or U24586 (N_24586,N_23810,N_23058);
nor U24587 (N_24587,N_23291,N_23915);
nand U24588 (N_24588,N_23916,N_23817);
and U24589 (N_24589,N_23437,N_23027);
or U24590 (N_24590,N_22942,N_22545);
and U24591 (N_24591,N_22812,N_22656);
nor U24592 (N_24592,N_23391,N_23653);
nor U24593 (N_24593,N_23497,N_23894);
nand U24594 (N_24594,N_23375,N_22813);
or U24595 (N_24595,N_22660,N_23614);
and U24596 (N_24596,N_23926,N_22788);
or U24597 (N_24597,N_22809,N_22819);
and U24598 (N_24598,N_23144,N_23757);
or U24599 (N_24599,N_23987,N_23149);
or U24600 (N_24600,N_22783,N_23618);
and U24601 (N_24601,N_23325,N_22648);
nand U24602 (N_24602,N_23893,N_22925);
xor U24603 (N_24603,N_23792,N_22699);
and U24604 (N_24604,N_23458,N_23330);
xor U24605 (N_24605,N_23733,N_23642);
xor U24606 (N_24606,N_23455,N_23891);
and U24607 (N_24607,N_23373,N_23090);
or U24608 (N_24608,N_23572,N_23877);
nand U24609 (N_24609,N_23208,N_23020);
and U24610 (N_24610,N_23809,N_23929);
xor U24611 (N_24611,N_23405,N_22687);
nand U24612 (N_24612,N_23955,N_23550);
or U24613 (N_24613,N_23559,N_23774);
or U24614 (N_24614,N_23347,N_23057);
xor U24615 (N_24615,N_23048,N_22867);
xnor U24616 (N_24616,N_22970,N_22696);
or U24617 (N_24617,N_23066,N_23547);
xor U24618 (N_24618,N_23728,N_23154);
and U24619 (N_24619,N_23314,N_22901);
and U24620 (N_24620,N_22841,N_23354);
nand U24621 (N_24621,N_23206,N_23900);
nand U24622 (N_24622,N_22530,N_23256);
or U24623 (N_24623,N_22607,N_22779);
nand U24624 (N_24624,N_23269,N_22968);
xnor U24625 (N_24625,N_23783,N_22553);
or U24626 (N_24626,N_23841,N_23707);
and U24627 (N_24627,N_23398,N_22515);
xor U24628 (N_24628,N_23050,N_23077);
nor U24629 (N_24629,N_23863,N_23184);
nor U24630 (N_24630,N_23262,N_22723);
nand U24631 (N_24631,N_22943,N_23525);
nand U24632 (N_24632,N_23594,N_22827);
nand U24633 (N_24633,N_23849,N_23052);
nand U24634 (N_24634,N_22577,N_23701);
or U24635 (N_24635,N_23081,N_23513);
nor U24636 (N_24636,N_23825,N_23565);
nand U24637 (N_24637,N_23651,N_23684);
or U24638 (N_24638,N_22814,N_23080);
or U24639 (N_24639,N_23824,N_23000);
nor U24640 (N_24640,N_22982,N_22828);
or U24641 (N_24641,N_23763,N_23393);
and U24642 (N_24642,N_23265,N_22793);
and U24643 (N_24643,N_23958,N_23581);
and U24644 (N_24644,N_23686,N_22938);
xor U24645 (N_24645,N_23557,N_23828);
and U24646 (N_24646,N_23917,N_23666);
nor U24647 (N_24647,N_22524,N_22945);
xor U24648 (N_24648,N_22971,N_23304);
nand U24649 (N_24649,N_23552,N_23499);
nand U24650 (N_24650,N_22897,N_23560);
nor U24651 (N_24651,N_22721,N_22915);
xnor U24652 (N_24652,N_22567,N_23266);
xor U24653 (N_24653,N_23591,N_22570);
nand U24654 (N_24654,N_23177,N_23739);
xnor U24655 (N_24655,N_22969,N_23679);
nand U24656 (N_24656,N_23360,N_22879);
xor U24657 (N_24657,N_23068,N_23930);
and U24658 (N_24658,N_23851,N_22675);
and U24659 (N_24659,N_22579,N_22748);
or U24660 (N_24660,N_23418,N_23280);
and U24661 (N_24661,N_23820,N_22822);
xnor U24662 (N_24662,N_22604,N_23768);
nor U24663 (N_24663,N_23785,N_23612);
or U24664 (N_24664,N_23790,N_23178);
or U24665 (N_24665,N_23953,N_23143);
or U24666 (N_24666,N_23480,N_23376);
nor U24667 (N_24667,N_22983,N_22888);
and U24668 (N_24668,N_23922,N_22999);
nand U24669 (N_24669,N_23022,N_23117);
and U24670 (N_24670,N_22868,N_23356);
or U24671 (N_24671,N_22905,N_23754);
nor U24672 (N_24672,N_22639,N_23685);
nand U24673 (N_24673,N_22679,N_23188);
nor U24674 (N_24674,N_23793,N_23794);
nor U24675 (N_24675,N_23663,N_22585);
nor U24676 (N_24676,N_23562,N_23311);
xnor U24677 (N_24677,N_22554,N_22555);
or U24678 (N_24678,N_22740,N_22875);
or U24679 (N_24679,N_22728,N_23031);
nor U24680 (N_24680,N_23274,N_22562);
nor U24681 (N_24681,N_23822,N_23412);
nand U24682 (N_24682,N_23231,N_23624);
nor U24683 (N_24683,N_23469,N_23051);
xnor U24684 (N_24684,N_23349,N_23625);
nand U24685 (N_24685,N_22563,N_22902);
nand U24686 (N_24686,N_23134,N_23539);
or U24687 (N_24687,N_23516,N_22617);
nor U24688 (N_24688,N_22820,N_23043);
nor U24689 (N_24689,N_23886,N_23939);
nand U24690 (N_24690,N_23316,N_22508);
and U24691 (N_24691,N_23880,N_22981);
or U24692 (N_24692,N_23593,N_23385);
xnor U24693 (N_24693,N_22876,N_22916);
and U24694 (N_24694,N_22844,N_22635);
nand U24695 (N_24695,N_22949,N_23766);
and U24696 (N_24696,N_22741,N_23570);
or U24697 (N_24697,N_22872,N_22931);
or U24698 (N_24698,N_23468,N_22862);
nor U24699 (N_24699,N_23813,N_22663);
xnor U24700 (N_24700,N_23604,N_23029);
nand U24701 (N_24701,N_23745,N_23968);
xor U24702 (N_24702,N_22775,N_23185);
nand U24703 (N_24703,N_23735,N_23201);
or U24704 (N_24704,N_23378,N_23747);
and U24705 (N_24705,N_23485,N_22992);
nor U24706 (N_24706,N_23542,N_22597);
nand U24707 (N_24707,N_22743,N_23098);
nand U24708 (N_24708,N_23773,N_22863);
or U24709 (N_24709,N_22590,N_23636);
xor U24710 (N_24710,N_23629,N_23938);
and U24711 (N_24711,N_23744,N_22877);
and U24712 (N_24712,N_22910,N_23681);
xor U24713 (N_24713,N_23225,N_23621);
nor U24714 (N_24714,N_22616,N_23404);
and U24715 (N_24715,N_23146,N_22623);
nor U24716 (N_24716,N_23115,N_23932);
xor U24717 (N_24717,N_23816,N_23442);
nand U24718 (N_24718,N_23579,N_23704);
and U24719 (N_24719,N_23732,N_22930);
xor U24720 (N_24720,N_22893,N_22855);
nor U24721 (N_24721,N_23289,N_23186);
nand U24722 (N_24722,N_23620,N_22502);
nand U24723 (N_24723,N_23340,N_22746);
nor U24724 (N_24724,N_23823,N_23533);
nor U24725 (N_24725,N_22666,N_22903);
xor U24726 (N_24726,N_23009,N_23731);
or U24727 (N_24727,N_22655,N_23443);
and U24728 (N_24728,N_23945,N_23282);
nand U24729 (N_24729,N_23107,N_23957);
xor U24730 (N_24730,N_23638,N_22640);
and U24731 (N_24731,N_23596,N_23553);
nor U24732 (N_24732,N_23697,N_23952);
nand U24733 (N_24733,N_22664,N_23319);
nand U24734 (N_24734,N_23761,N_22755);
or U24735 (N_24735,N_23947,N_23308);
or U24736 (N_24736,N_23415,N_23292);
nand U24737 (N_24737,N_22807,N_23906);
nor U24738 (N_24738,N_22588,N_23606);
nand U24739 (N_24739,N_23857,N_23411);
nand U24740 (N_24740,N_23867,N_23635);
nor U24741 (N_24741,N_23942,N_22936);
or U24742 (N_24742,N_23585,N_23613);
nand U24743 (N_24743,N_23200,N_22736);
nor U24744 (N_24744,N_23298,N_23536);
nand U24745 (N_24745,N_23961,N_23288);
or U24746 (N_24746,N_22637,N_23748);
xor U24747 (N_24747,N_22871,N_23161);
xor U24748 (N_24748,N_22599,N_23320);
xnor U24749 (N_24749,N_23623,N_23710);
xor U24750 (N_24750,N_23887,N_23773);
and U24751 (N_24751,N_23954,N_23790);
xnor U24752 (N_24752,N_23560,N_23671);
or U24753 (N_24753,N_23898,N_22848);
and U24754 (N_24754,N_23556,N_22633);
nand U24755 (N_24755,N_23923,N_22547);
nand U24756 (N_24756,N_23864,N_23336);
xnor U24757 (N_24757,N_23801,N_23080);
or U24758 (N_24758,N_23731,N_22784);
xnor U24759 (N_24759,N_22657,N_22597);
nand U24760 (N_24760,N_22914,N_22898);
nor U24761 (N_24761,N_23727,N_23048);
xor U24762 (N_24762,N_23563,N_22620);
nand U24763 (N_24763,N_23687,N_23526);
or U24764 (N_24764,N_23053,N_23452);
nand U24765 (N_24765,N_23604,N_23496);
nand U24766 (N_24766,N_22941,N_23163);
or U24767 (N_24767,N_23500,N_22864);
nand U24768 (N_24768,N_22667,N_23493);
or U24769 (N_24769,N_22608,N_23691);
or U24770 (N_24770,N_22957,N_22747);
nor U24771 (N_24771,N_23794,N_23959);
nand U24772 (N_24772,N_23957,N_23353);
nor U24773 (N_24773,N_23245,N_23156);
and U24774 (N_24774,N_23331,N_22708);
or U24775 (N_24775,N_22570,N_23584);
or U24776 (N_24776,N_23005,N_23290);
nor U24777 (N_24777,N_23895,N_23524);
or U24778 (N_24778,N_22687,N_23662);
nand U24779 (N_24779,N_23802,N_23345);
nand U24780 (N_24780,N_22713,N_22782);
nand U24781 (N_24781,N_23690,N_22760);
nand U24782 (N_24782,N_23063,N_23313);
and U24783 (N_24783,N_23205,N_22570);
nand U24784 (N_24784,N_23997,N_22621);
nand U24785 (N_24785,N_22573,N_22654);
or U24786 (N_24786,N_23454,N_23641);
xnor U24787 (N_24787,N_22946,N_23008);
nor U24788 (N_24788,N_22545,N_23374);
or U24789 (N_24789,N_23409,N_23615);
xor U24790 (N_24790,N_23038,N_23088);
or U24791 (N_24791,N_23781,N_22985);
or U24792 (N_24792,N_23650,N_22766);
nand U24793 (N_24793,N_22619,N_23533);
nor U24794 (N_24794,N_23926,N_22643);
nand U24795 (N_24795,N_23951,N_23211);
or U24796 (N_24796,N_22924,N_23466);
nor U24797 (N_24797,N_23372,N_23410);
and U24798 (N_24798,N_22916,N_22891);
and U24799 (N_24799,N_22731,N_23597);
nand U24800 (N_24800,N_23549,N_23665);
and U24801 (N_24801,N_23398,N_23145);
nand U24802 (N_24802,N_23530,N_23613);
and U24803 (N_24803,N_23337,N_22944);
nor U24804 (N_24804,N_23662,N_23218);
nor U24805 (N_24805,N_23051,N_22506);
or U24806 (N_24806,N_23051,N_22878);
nor U24807 (N_24807,N_23672,N_22966);
xor U24808 (N_24808,N_23981,N_23771);
and U24809 (N_24809,N_23068,N_22902);
nor U24810 (N_24810,N_23438,N_23939);
nor U24811 (N_24811,N_22670,N_22983);
or U24812 (N_24812,N_23147,N_23487);
nor U24813 (N_24813,N_23735,N_23400);
xnor U24814 (N_24814,N_22564,N_23323);
nor U24815 (N_24815,N_23019,N_22562);
xor U24816 (N_24816,N_22905,N_22999);
and U24817 (N_24817,N_23143,N_22588);
and U24818 (N_24818,N_23473,N_23648);
nand U24819 (N_24819,N_22955,N_23549);
or U24820 (N_24820,N_22877,N_23675);
and U24821 (N_24821,N_22717,N_22971);
nand U24822 (N_24822,N_23068,N_23512);
or U24823 (N_24823,N_23144,N_23731);
and U24824 (N_24824,N_22557,N_22551);
or U24825 (N_24825,N_23745,N_23358);
nand U24826 (N_24826,N_22944,N_23793);
xnor U24827 (N_24827,N_23779,N_22548);
xor U24828 (N_24828,N_22943,N_23087);
or U24829 (N_24829,N_22643,N_23426);
or U24830 (N_24830,N_23579,N_22834);
and U24831 (N_24831,N_23983,N_23165);
or U24832 (N_24832,N_23376,N_22926);
xor U24833 (N_24833,N_23234,N_23556);
nor U24834 (N_24834,N_22707,N_23707);
nand U24835 (N_24835,N_23456,N_23370);
or U24836 (N_24836,N_22511,N_23030);
and U24837 (N_24837,N_23322,N_22753);
xnor U24838 (N_24838,N_23141,N_23122);
nor U24839 (N_24839,N_23966,N_22968);
nand U24840 (N_24840,N_23937,N_23414);
and U24841 (N_24841,N_23755,N_23120);
xnor U24842 (N_24842,N_23929,N_23500);
nand U24843 (N_24843,N_23697,N_22654);
nor U24844 (N_24844,N_23444,N_23550);
nor U24845 (N_24845,N_23354,N_22822);
or U24846 (N_24846,N_22959,N_22515);
xnor U24847 (N_24847,N_22527,N_23145);
xor U24848 (N_24848,N_23006,N_22845);
nand U24849 (N_24849,N_23315,N_23280);
nor U24850 (N_24850,N_22627,N_23795);
xnor U24851 (N_24851,N_22624,N_22806);
or U24852 (N_24852,N_23153,N_23405);
xnor U24853 (N_24853,N_22819,N_22753);
and U24854 (N_24854,N_22828,N_23163);
xnor U24855 (N_24855,N_23811,N_22622);
nand U24856 (N_24856,N_22805,N_22893);
or U24857 (N_24857,N_23672,N_23887);
xnor U24858 (N_24858,N_23499,N_22503);
nor U24859 (N_24859,N_23030,N_23862);
nor U24860 (N_24860,N_22521,N_23548);
xor U24861 (N_24861,N_23725,N_23914);
nand U24862 (N_24862,N_22819,N_23291);
nor U24863 (N_24863,N_23423,N_22934);
and U24864 (N_24864,N_22686,N_23392);
nor U24865 (N_24865,N_23241,N_23307);
and U24866 (N_24866,N_23206,N_23382);
xor U24867 (N_24867,N_23378,N_23812);
nor U24868 (N_24868,N_23321,N_22756);
or U24869 (N_24869,N_22888,N_23356);
or U24870 (N_24870,N_23520,N_22692);
nor U24871 (N_24871,N_23030,N_22807);
nor U24872 (N_24872,N_23650,N_22991);
xnor U24873 (N_24873,N_23875,N_23454);
nand U24874 (N_24874,N_23671,N_23305);
and U24875 (N_24875,N_22852,N_22869);
nand U24876 (N_24876,N_23800,N_23238);
or U24877 (N_24877,N_23916,N_22776);
nor U24878 (N_24878,N_23306,N_23787);
xor U24879 (N_24879,N_23534,N_23169);
xor U24880 (N_24880,N_22530,N_23116);
or U24881 (N_24881,N_23906,N_22931);
xnor U24882 (N_24882,N_23777,N_23697);
nor U24883 (N_24883,N_23819,N_22566);
xnor U24884 (N_24884,N_22809,N_22611);
nand U24885 (N_24885,N_23244,N_23913);
xnor U24886 (N_24886,N_22983,N_22773);
or U24887 (N_24887,N_23163,N_22641);
nand U24888 (N_24888,N_22920,N_23271);
nand U24889 (N_24889,N_23594,N_22757);
nor U24890 (N_24890,N_23992,N_22726);
xnor U24891 (N_24891,N_23364,N_23277);
or U24892 (N_24892,N_22941,N_23269);
and U24893 (N_24893,N_23541,N_22991);
nand U24894 (N_24894,N_22717,N_23567);
xnor U24895 (N_24895,N_22955,N_23652);
nand U24896 (N_24896,N_23523,N_23076);
nand U24897 (N_24897,N_23308,N_22928);
xnor U24898 (N_24898,N_23915,N_22851);
nand U24899 (N_24899,N_22960,N_23357);
nor U24900 (N_24900,N_23520,N_23482);
xnor U24901 (N_24901,N_22589,N_23870);
xor U24902 (N_24902,N_23831,N_22769);
and U24903 (N_24903,N_23668,N_23088);
and U24904 (N_24904,N_22946,N_23595);
nor U24905 (N_24905,N_23954,N_22918);
nand U24906 (N_24906,N_23835,N_23610);
and U24907 (N_24907,N_23757,N_23030);
nor U24908 (N_24908,N_22552,N_22526);
nand U24909 (N_24909,N_22621,N_23461);
or U24910 (N_24910,N_23233,N_22880);
nand U24911 (N_24911,N_23445,N_22770);
nand U24912 (N_24912,N_23108,N_22749);
or U24913 (N_24913,N_22888,N_23280);
and U24914 (N_24914,N_23598,N_23502);
nor U24915 (N_24915,N_22985,N_22915);
nor U24916 (N_24916,N_23419,N_23783);
xor U24917 (N_24917,N_23349,N_23350);
or U24918 (N_24918,N_23039,N_22542);
and U24919 (N_24919,N_23318,N_23552);
nor U24920 (N_24920,N_22852,N_23023);
nor U24921 (N_24921,N_22988,N_23438);
nor U24922 (N_24922,N_23144,N_23602);
nand U24923 (N_24923,N_23066,N_23089);
and U24924 (N_24924,N_22883,N_22528);
or U24925 (N_24925,N_23820,N_22719);
xnor U24926 (N_24926,N_23973,N_23565);
and U24927 (N_24927,N_23641,N_22698);
or U24928 (N_24928,N_22757,N_23754);
xor U24929 (N_24929,N_23181,N_23634);
or U24930 (N_24930,N_23012,N_22635);
and U24931 (N_24931,N_23091,N_23113);
xor U24932 (N_24932,N_23680,N_23462);
and U24933 (N_24933,N_23019,N_23451);
and U24934 (N_24934,N_23123,N_23385);
nand U24935 (N_24935,N_23109,N_22998);
xor U24936 (N_24936,N_23109,N_23581);
nor U24937 (N_24937,N_22534,N_23616);
or U24938 (N_24938,N_23255,N_23488);
xor U24939 (N_24939,N_23150,N_22942);
or U24940 (N_24940,N_22513,N_23903);
and U24941 (N_24941,N_23313,N_22841);
xor U24942 (N_24942,N_22544,N_22802);
or U24943 (N_24943,N_23435,N_23413);
nor U24944 (N_24944,N_23599,N_23131);
or U24945 (N_24945,N_23473,N_23651);
nor U24946 (N_24946,N_23192,N_22830);
and U24947 (N_24947,N_23208,N_22600);
xnor U24948 (N_24948,N_23247,N_23454);
and U24949 (N_24949,N_23825,N_22724);
nand U24950 (N_24950,N_22643,N_22763);
xnor U24951 (N_24951,N_23721,N_23833);
nor U24952 (N_24952,N_22966,N_22638);
nand U24953 (N_24953,N_23893,N_22504);
xor U24954 (N_24954,N_23447,N_22582);
nor U24955 (N_24955,N_23599,N_23648);
nand U24956 (N_24956,N_22823,N_23934);
xor U24957 (N_24957,N_23134,N_23381);
nor U24958 (N_24958,N_23239,N_22848);
and U24959 (N_24959,N_23352,N_22994);
or U24960 (N_24960,N_22945,N_23451);
xor U24961 (N_24961,N_23182,N_23036);
nor U24962 (N_24962,N_23028,N_23461);
nand U24963 (N_24963,N_22871,N_23563);
nand U24964 (N_24964,N_22683,N_22978);
nand U24965 (N_24965,N_23424,N_22756);
and U24966 (N_24966,N_23131,N_23043);
and U24967 (N_24967,N_22572,N_22559);
xor U24968 (N_24968,N_22696,N_23543);
nor U24969 (N_24969,N_23257,N_23128);
nand U24970 (N_24970,N_22520,N_23296);
nand U24971 (N_24971,N_23876,N_23997);
nor U24972 (N_24972,N_23148,N_23158);
and U24973 (N_24973,N_22871,N_23464);
nor U24974 (N_24974,N_22907,N_22709);
xor U24975 (N_24975,N_23311,N_23635);
and U24976 (N_24976,N_23022,N_22530);
or U24977 (N_24977,N_22634,N_23659);
nor U24978 (N_24978,N_23585,N_22697);
and U24979 (N_24979,N_23438,N_23763);
or U24980 (N_24980,N_23027,N_23799);
or U24981 (N_24981,N_23928,N_23606);
nor U24982 (N_24982,N_23777,N_22594);
and U24983 (N_24983,N_23512,N_23355);
nor U24984 (N_24984,N_22823,N_23933);
nand U24985 (N_24985,N_23296,N_22655);
and U24986 (N_24986,N_22792,N_23572);
nand U24987 (N_24987,N_22807,N_22509);
and U24988 (N_24988,N_22594,N_23511);
xor U24989 (N_24989,N_22701,N_23394);
nand U24990 (N_24990,N_23830,N_22742);
and U24991 (N_24991,N_22647,N_22899);
xnor U24992 (N_24992,N_22533,N_23479);
or U24993 (N_24993,N_23667,N_23072);
and U24994 (N_24994,N_23083,N_23767);
nor U24995 (N_24995,N_23967,N_23748);
and U24996 (N_24996,N_23961,N_22941);
nor U24997 (N_24997,N_23374,N_23058);
and U24998 (N_24998,N_22660,N_23900);
xnor U24999 (N_24999,N_23568,N_23039);
nand U25000 (N_25000,N_23304,N_22653);
xor U25001 (N_25001,N_23632,N_23773);
and U25002 (N_25002,N_22768,N_23552);
nand U25003 (N_25003,N_23668,N_23561);
xor U25004 (N_25004,N_22803,N_22890);
or U25005 (N_25005,N_23770,N_23659);
xnor U25006 (N_25006,N_23560,N_23910);
or U25007 (N_25007,N_23454,N_23035);
nand U25008 (N_25008,N_23950,N_23956);
xor U25009 (N_25009,N_23516,N_23896);
nor U25010 (N_25010,N_23696,N_22506);
nor U25011 (N_25011,N_23118,N_23617);
or U25012 (N_25012,N_22530,N_23671);
nor U25013 (N_25013,N_23971,N_23343);
xor U25014 (N_25014,N_23223,N_23434);
nand U25015 (N_25015,N_23714,N_23426);
nand U25016 (N_25016,N_22962,N_22680);
xnor U25017 (N_25017,N_23682,N_23522);
nor U25018 (N_25018,N_23724,N_23883);
xor U25019 (N_25019,N_23935,N_22979);
and U25020 (N_25020,N_23503,N_23786);
and U25021 (N_25021,N_23802,N_22758);
and U25022 (N_25022,N_22818,N_23043);
or U25023 (N_25023,N_23590,N_23833);
and U25024 (N_25024,N_23466,N_23605);
or U25025 (N_25025,N_23563,N_23506);
nand U25026 (N_25026,N_23904,N_23048);
nor U25027 (N_25027,N_23679,N_22597);
or U25028 (N_25028,N_23934,N_23794);
and U25029 (N_25029,N_23899,N_23515);
xnor U25030 (N_25030,N_23509,N_23407);
nand U25031 (N_25031,N_23307,N_23379);
or U25032 (N_25032,N_22973,N_23821);
nor U25033 (N_25033,N_23134,N_22586);
xnor U25034 (N_25034,N_23346,N_22705);
xnor U25035 (N_25035,N_23147,N_23710);
nor U25036 (N_25036,N_23038,N_23060);
nand U25037 (N_25037,N_23306,N_22625);
nand U25038 (N_25038,N_23939,N_23170);
and U25039 (N_25039,N_22679,N_23920);
and U25040 (N_25040,N_23017,N_23707);
and U25041 (N_25041,N_23750,N_23725);
nor U25042 (N_25042,N_22853,N_23504);
or U25043 (N_25043,N_22646,N_23349);
xnor U25044 (N_25044,N_22919,N_22752);
nor U25045 (N_25045,N_23502,N_23959);
nor U25046 (N_25046,N_22869,N_23962);
and U25047 (N_25047,N_23063,N_23309);
xor U25048 (N_25048,N_23147,N_22536);
nand U25049 (N_25049,N_23570,N_23457);
nor U25050 (N_25050,N_22686,N_23147);
xnor U25051 (N_25051,N_23362,N_23129);
nor U25052 (N_25052,N_23563,N_22854);
and U25053 (N_25053,N_23215,N_22571);
nand U25054 (N_25054,N_23808,N_23390);
and U25055 (N_25055,N_22829,N_23319);
and U25056 (N_25056,N_23575,N_22543);
and U25057 (N_25057,N_23447,N_23387);
or U25058 (N_25058,N_22952,N_22908);
or U25059 (N_25059,N_23327,N_22505);
nand U25060 (N_25060,N_22861,N_23855);
nor U25061 (N_25061,N_22762,N_23124);
and U25062 (N_25062,N_23402,N_23720);
or U25063 (N_25063,N_23894,N_23133);
or U25064 (N_25064,N_23048,N_23461);
nand U25065 (N_25065,N_23834,N_23047);
or U25066 (N_25066,N_23305,N_23869);
nor U25067 (N_25067,N_23277,N_23617);
or U25068 (N_25068,N_23448,N_23415);
nand U25069 (N_25069,N_23126,N_23829);
or U25070 (N_25070,N_23983,N_23981);
and U25071 (N_25071,N_23604,N_23278);
xnor U25072 (N_25072,N_23326,N_22708);
and U25073 (N_25073,N_22761,N_22967);
xnor U25074 (N_25074,N_22533,N_23437);
and U25075 (N_25075,N_22893,N_22869);
xor U25076 (N_25076,N_22690,N_22562);
and U25077 (N_25077,N_23321,N_23318);
xor U25078 (N_25078,N_22625,N_23249);
nor U25079 (N_25079,N_23146,N_23747);
xor U25080 (N_25080,N_22830,N_23279);
xor U25081 (N_25081,N_23239,N_23224);
and U25082 (N_25082,N_23901,N_22837);
or U25083 (N_25083,N_23430,N_23058);
or U25084 (N_25084,N_23555,N_22534);
nand U25085 (N_25085,N_22587,N_23745);
nand U25086 (N_25086,N_23612,N_23841);
nand U25087 (N_25087,N_23253,N_22783);
or U25088 (N_25088,N_23269,N_22719);
or U25089 (N_25089,N_23646,N_23005);
and U25090 (N_25090,N_23553,N_22577);
or U25091 (N_25091,N_23641,N_22547);
and U25092 (N_25092,N_23605,N_22872);
and U25093 (N_25093,N_22700,N_22789);
nand U25094 (N_25094,N_23584,N_22996);
and U25095 (N_25095,N_22901,N_22586);
or U25096 (N_25096,N_23805,N_23131);
xor U25097 (N_25097,N_23776,N_23341);
or U25098 (N_25098,N_22534,N_23658);
xor U25099 (N_25099,N_23776,N_23610);
nor U25100 (N_25100,N_22677,N_23660);
or U25101 (N_25101,N_23382,N_23889);
xnor U25102 (N_25102,N_23264,N_23645);
nor U25103 (N_25103,N_22690,N_22803);
nor U25104 (N_25104,N_23709,N_23730);
xor U25105 (N_25105,N_23250,N_23192);
or U25106 (N_25106,N_23117,N_23516);
and U25107 (N_25107,N_23659,N_23541);
nor U25108 (N_25108,N_23811,N_23560);
or U25109 (N_25109,N_23979,N_23365);
nand U25110 (N_25110,N_23448,N_23390);
nand U25111 (N_25111,N_23818,N_23299);
and U25112 (N_25112,N_23157,N_23016);
nor U25113 (N_25113,N_23252,N_23171);
or U25114 (N_25114,N_23614,N_22582);
or U25115 (N_25115,N_22947,N_23749);
xnor U25116 (N_25116,N_22738,N_22658);
or U25117 (N_25117,N_23619,N_23514);
xnor U25118 (N_25118,N_23863,N_22839);
nor U25119 (N_25119,N_22563,N_22827);
nor U25120 (N_25120,N_22718,N_23382);
nand U25121 (N_25121,N_22785,N_23300);
nor U25122 (N_25122,N_22682,N_23791);
or U25123 (N_25123,N_23536,N_22615);
or U25124 (N_25124,N_22680,N_22552);
xnor U25125 (N_25125,N_22826,N_23810);
xnor U25126 (N_25126,N_23341,N_23757);
and U25127 (N_25127,N_23755,N_23138);
nand U25128 (N_25128,N_23658,N_23020);
xnor U25129 (N_25129,N_23158,N_22737);
and U25130 (N_25130,N_23786,N_22813);
nand U25131 (N_25131,N_23322,N_23337);
nand U25132 (N_25132,N_23644,N_23232);
nor U25133 (N_25133,N_23165,N_23848);
nor U25134 (N_25134,N_22956,N_23929);
or U25135 (N_25135,N_22509,N_23507);
and U25136 (N_25136,N_22597,N_22943);
xor U25137 (N_25137,N_23191,N_22711);
nand U25138 (N_25138,N_23377,N_23534);
or U25139 (N_25139,N_23909,N_22725);
xnor U25140 (N_25140,N_23728,N_22722);
nor U25141 (N_25141,N_23939,N_23577);
or U25142 (N_25142,N_23474,N_23158);
nand U25143 (N_25143,N_22591,N_22962);
nor U25144 (N_25144,N_23229,N_23963);
and U25145 (N_25145,N_23537,N_22750);
xnor U25146 (N_25146,N_23506,N_23914);
nand U25147 (N_25147,N_22776,N_23698);
or U25148 (N_25148,N_23245,N_23491);
xor U25149 (N_25149,N_22712,N_22694);
xnor U25150 (N_25150,N_23297,N_23449);
nor U25151 (N_25151,N_23349,N_23494);
or U25152 (N_25152,N_23856,N_23741);
nor U25153 (N_25153,N_23179,N_22536);
nor U25154 (N_25154,N_23275,N_23053);
and U25155 (N_25155,N_23111,N_22526);
nand U25156 (N_25156,N_22871,N_23790);
and U25157 (N_25157,N_23252,N_22703);
and U25158 (N_25158,N_23198,N_23803);
or U25159 (N_25159,N_23391,N_22879);
or U25160 (N_25160,N_22778,N_22887);
and U25161 (N_25161,N_22508,N_23531);
or U25162 (N_25162,N_23538,N_23354);
and U25163 (N_25163,N_23217,N_23289);
xor U25164 (N_25164,N_23535,N_22573);
and U25165 (N_25165,N_23407,N_23616);
nor U25166 (N_25166,N_23353,N_23713);
nor U25167 (N_25167,N_22884,N_23628);
or U25168 (N_25168,N_22533,N_23619);
nand U25169 (N_25169,N_23213,N_23586);
nor U25170 (N_25170,N_23558,N_22903);
xor U25171 (N_25171,N_23843,N_23665);
xor U25172 (N_25172,N_23659,N_23562);
nor U25173 (N_25173,N_23009,N_23733);
nor U25174 (N_25174,N_23563,N_23220);
or U25175 (N_25175,N_23476,N_23521);
xnor U25176 (N_25176,N_23978,N_23112);
nor U25177 (N_25177,N_22586,N_23744);
and U25178 (N_25178,N_23275,N_22668);
nand U25179 (N_25179,N_23905,N_23606);
and U25180 (N_25180,N_22551,N_22611);
and U25181 (N_25181,N_23708,N_23940);
nor U25182 (N_25182,N_23051,N_22796);
nor U25183 (N_25183,N_22821,N_23225);
xnor U25184 (N_25184,N_23901,N_22868);
nand U25185 (N_25185,N_23914,N_23598);
or U25186 (N_25186,N_22619,N_22724);
nor U25187 (N_25187,N_23926,N_22613);
xor U25188 (N_25188,N_23257,N_22994);
and U25189 (N_25189,N_23165,N_22521);
nor U25190 (N_25190,N_22776,N_23008);
xnor U25191 (N_25191,N_23002,N_23244);
xnor U25192 (N_25192,N_23070,N_23590);
nor U25193 (N_25193,N_22943,N_23281);
xor U25194 (N_25194,N_22907,N_23713);
nor U25195 (N_25195,N_22669,N_22666);
nand U25196 (N_25196,N_23402,N_22635);
and U25197 (N_25197,N_23783,N_23927);
nand U25198 (N_25198,N_22841,N_22794);
nor U25199 (N_25199,N_23415,N_23016);
nand U25200 (N_25200,N_22884,N_23126);
nand U25201 (N_25201,N_23717,N_23825);
nor U25202 (N_25202,N_22813,N_23490);
nor U25203 (N_25203,N_22993,N_22724);
xnor U25204 (N_25204,N_23235,N_22932);
and U25205 (N_25205,N_23628,N_23011);
xnor U25206 (N_25206,N_23322,N_22504);
and U25207 (N_25207,N_23414,N_23462);
nand U25208 (N_25208,N_23262,N_23365);
nor U25209 (N_25209,N_23698,N_22772);
nor U25210 (N_25210,N_22671,N_23869);
xor U25211 (N_25211,N_23114,N_23905);
nor U25212 (N_25212,N_23594,N_23114);
nand U25213 (N_25213,N_22589,N_23290);
xor U25214 (N_25214,N_22582,N_23138);
nand U25215 (N_25215,N_23571,N_22692);
nand U25216 (N_25216,N_22599,N_23799);
nand U25217 (N_25217,N_23437,N_22700);
and U25218 (N_25218,N_23827,N_23798);
nor U25219 (N_25219,N_23783,N_23127);
nor U25220 (N_25220,N_22623,N_23337);
and U25221 (N_25221,N_23819,N_23879);
or U25222 (N_25222,N_23182,N_23933);
or U25223 (N_25223,N_23776,N_22742);
nand U25224 (N_25224,N_23752,N_23769);
xnor U25225 (N_25225,N_23903,N_23786);
and U25226 (N_25226,N_23761,N_23363);
xor U25227 (N_25227,N_23848,N_23836);
or U25228 (N_25228,N_23056,N_23794);
nor U25229 (N_25229,N_23987,N_23567);
nand U25230 (N_25230,N_22509,N_22867);
or U25231 (N_25231,N_23546,N_22861);
nand U25232 (N_25232,N_23048,N_23805);
nand U25233 (N_25233,N_23519,N_23587);
or U25234 (N_25234,N_23335,N_22626);
and U25235 (N_25235,N_23747,N_23510);
xor U25236 (N_25236,N_22978,N_23465);
or U25237 (N_25237,N_23930,N_22885);
and U25238 (N_25238,N_23913,N_22630);
nor U25239 (N_25239,N_23049,N_22969);
xnor U25240 (N_25240,N_23951,N_23518);
and U25241 (N_25241,N_23447,N_23216);
nand U25242 (N_25242,N_22604,N_22863);
or U25243 (N_25243,N_22976,N_23859);
and U25244 (N_25244,N_23573,N_23029);
nand U25245 (N_25245,N_23888,N_22541);
xnor U25246 (N_25246,N_23447,N_23919);
or U25247 (N_25247,N_23904,N_23391);
nand U25248 (N_25248,N_23005,N_23058);
nor U25249 (N_25249,N_23265,N_23273);
and U25250 (N_25250,N_22935,N_22941);
nor U25251 (N_25251,N_23915,N_23515);
nor U25252 (N_25252,N_22759,N_23271);
xor U25253 (N_25253,N_23127,N_23720);
and U25254 (N_25254,N_23074,N_23541);
xnor U25255 (N_25255,N_23323,N_23421);
or U25256 (N_25256,N_23822,N_23646);
xor U25257 (N_25257,N_23161,N_22936);
nand U25258 (N_25258,N_22561,N_22925);
nand U25259 (N_25259,N_23709,N_22951);
nand U25260 (N_25260,N_22916,N_23111);
nor U25261 (N_25261,N_22956,N_22652);
xnor U25262 (N_25262,N_23656,N_23448);
nor U25263 (N_25263,N_23777,N_22703);
nand U25264 (N_25264,N_23109,N_23210);
xnor U25265 (N_25265,N_23100,N_22791);
nor U25266 (N_25266,N_23109,N_23707);
or U25267 (N_25267,N_23523,N_22706);
xor U25268 (N_25268,N_22688,N_22611);
xor U25269 (N_25269,N_22990,N_23270);
xnor U25270 (N_25270,N_23189,N_23374);
nand U25271 (N_25271,N_22676,N_23928);
nand U25272 (N_25272,N_23070,N_23550);
or U25273 (N_25273,N_23418,N_23345);
and U25274 (N_25274,N_23750,N_23723);
and U25275 (N_25275,N_23709,N_23850);
xor U25276 (N_25276,N_23751,N_23355);
nor U25277 (N_25277,N_22702,N_22921);
nor U25278 (N_25278,N_23721,N_22571);
nor U25279 (N_25279,N_22997,N_23952);
or U25280 (N_25280,N_23147,N_23538);
xnor U25281 (N_25281,N_22702,N_23965);
or U25282 (N_25282,N_23853,N_22607);
xor U25283 (N_25283,N_22890,N_22656);
xnor U25284 (N_25284,N_23472,N_23691);
nor U25285 (N_25285,N_23213,N_22543);
nand U25286 (N_25286,N_23437,N_22885);
or U25287 (N_25287,N_23209,N_23241);
or U25288 (N_25288,N_23728,N_23058);
and U25289 (N_25289,N_23141,N_23774);
xor U25290 (N_25290,N_23784,N_22584);
and U25291 (N_25291,N_22838,N_23764);
or U25292 (N_25292,N_22882,N_23276);
and U25293 (N_25293,N_23642,N_23112);
or U25294 (N_25294,N_22825,N_23135);
nor U25295 (N_25295,N_23675,N_23644);
nor U25296 (N_25296,N_23463,N_23680);
or U25297 (N_25297,N_22714,N_22562);
nand U25298 (N_25298,N_23049,N_22709);
nor U25299 (N_25299,N_23708,N_22566);
nand U25300 (N_25300,N_22593,N_22808);
nor U25301 (N_25301,N_23268,N_23648);
xor U25302 (N_25302,N_22914,N_23679);
nand U25303 (N_25303,N_22965,N_22781);
xnor U25304 (N_25304,N_22868,N_22856);
nor U25305 (N_25305,N_23663,N_23715);
or U25306 (N_25306,N_23668,N_23718);
or U25307 (N_25307,N_23486,N_23795);
nand U25308 (N_25308,N_23234,N_23680);
xnor U25309 (N_25309,N_22862,N_23590);
xor U25310 (N_25310,N_23051,N_23565);
or U25311 (N_25311,N_23700,N_23789);
and U25312 (N_25312,N_22636,N_22568);
nand U25313 (N_25313,N_22927,N_23305);
xnor U25314 (N_25314,N_23130,N_22681);
or U25315 (N_25315,N_23817,N_22858);
xnor U25316 (N_25316,N_23325,N_22917);
xnor U25317 (N_25317,N_23244,N_23364);
xnor U25318 (N_25318,N_23397,N_23923);
and U25319 (N_25319,N_22544,N_23255);
xor U25320 (N_25320,N_22770,N_23985);
or U25321 (N_25321,N_22715,N_23076);
and U25322 (N_25322,N_23875,N_23187);
nand U25323 (N_25323,N_23820,N_23496);
xnor U25324 (N_25324,N_22502,N_23798);
nand U25325 (N_25325,N_23332,N_22627);
or U25326 (N_25326,N_23797,N_22731);
or U25327 (N_25327,N_23092,N_22522);
xnor U25328 (N_25328,N_22764,N_22516);
xor U25329 (N_25329,N_22979,N_22839);
or U25330 (N_25330,N_23652,N_23963);
nand U25331 (N_25331,N_23369,N_23777);
nor U25332 (N_25332,N_22802,N_23986);
xnor U25333 (N_25333,N_23412,N_22883);
xnor U25334 (N_25334,N_23365,N_22739);
or U25335 (N_25335,N_23889,N_22698);
nor U25336 (N_25336,N_22777,N_23721);
nor U25337 (N_25337,N_23452,N_23226);
nand U25338 (N_25338,N_23684,N_23379);
and U25339 (N_25339,N_23201,N_22536);
nand U25340 (N_25340,N_23087,N_23675);
nor U25341 (N_25341,N_23955,N_23819);
nand U25342 (N_25342,N_23281,N_23298);
nand U25343 (N_25343,N_22794,N_22518);
nand U25344 (N_25344,N_22678,N_23309);
nor U25345 (N_25345,N_22768,N_23338);
or U25346 (N_25346,N_23241,N_23870);
and U25347 (N_25347,N_23524,N_23052);
xnor U25348 (N_25348,N_23174,N_23220);
or U25349 (N_25349,N_22842,N_22560);
nor U25350 (N_25350,N_22592,N_23047);
nor U25351 (N_25351,N_23736,N_23070);
nand U25352 (N_25352,N_23715,N_23895);
or U25353 (N_25353,N_23808,N_22664);
nand U25354 (N_25354,N_22915,N_23540);
nor U25355 (N_25355,N_23352,N_23041);
xor U25356 (N_25356,N_23715,N_23125);
or U25357 (N_25357,N_23370,N_23187);
nor U25358 (N_25358,N_23370,N_22650);
nand U25359 (N_25359,N_22673,N_23623);
nor U25360 (N_25360,N_22757,N_23071);
nor U25361 (N_25361,N_23150,N_23891);
nand U25362 (N_25362,N_23481,N_23669);
nor U25363 (N_25363,N_23599,N_23313);
and U25364 (N_25364,N_23017,N_23735);
xor U25365 (N_25365,N_22867,N_22897);
xnor U25366 (N_25366,N_22841,N_22940);
and U25367 (N_25367,N_22610,N_23489);
nor U25368 (N_25368,N_23636,N_22810);
xnor U25369 (N_25369,N_22880,N_23493);
and U25370 (N_25370,N_23436,N_23689);
or U25371 (N_25371,N_23500,N_23377);
nand U25372 (N_25372,N_23306,N_23761);
or U25373 (N_25373,N_22784,N_22936);
xnor U25374 (N_25374,N_23668,N_23104);
nor U25375 (N_25375,N_22958,N_23997);
nand U25376 (N_25376,N_23032,N_22656);
or U25377 (N_25377,N_22798,N_22761);
nand U25378 (N_25378,N_23472,N_23515);
and U25379 (N_25379,N_22892,N_23753);
nand U25380 (N_25380,N_23246,N_23484);
or U25381 (N_25381,N_23812,N_23027);
xnor U25382 (N_25382,N_22964,N_23986);
nand U25383 (N_25383,N_23458,N_23827);
nand U25384 (N_25384,N_23698,N_23700);
nor U25385 (N_25385,N_23945,N_23444);
and U25386 (N_25386,N_22947,N_23569);
xnor U25387 (N_25387,N_23750,N_22995);
and U25388 (N_25388,N_22764,N_23411);
nor U25389 (N_25389,N_23512,N_23287);
and U25390 (N_25390,N_23493,N_23052);
nor U25391 (N_25391,N_22713,N_23618);
and U25392 (N_25392,N_23209,N_23383);
nand U25393 (N_25393,N_23724,N_22920);
and U25394 (N_25394,N_23908,N_22662);
xnor U25395 (N_25395,N_23623,N_23228);
nor U25396 (N_25396,N_23326,N_23261);
nand U25397 (N_25397,N_23351,N_23904);
or U25398 (N_25398,N_23309,N_23009);
nand U25399 (N_25399,N_23576,N_22962);
nor U25400 (N_25400,N_23540,N_22686);
or U25401 (N_25401,N_23257,N_23404);
nor U25402 (N_25402,N_23316,N_23256);
nand U25403 (N_25403,N_23961,N_22515);
xor U25404 (N_25404,N_23335,N_23555);
and U25405 (N_25405,N_22576,N_22559);
xnor U25406 (N_25406,N_22502,N_23169);
xnor U25407 (N_25407,N_22583,N_23688);
nor U25408 (N_25408,N_22979,N_23800);
and U25409 (N_25409,N_23425,N_23409);
nor U25410 (N_25410,N_23389,N_23351);
nand U25411 (N_25411,N_23559,N_23061);
nand U25412 (N_25412,N_23135,N_23873);
xor U25413 (N_25413,N_23674,N_22934);
nand U25414 (N_25414,N_23234,N_22766);
xnor U25415 (N_25415,N_23522,N_23819);
xnor U25416 (N_25416,N_23953,N_23615);
nor U25417 (N_25417,N_23820,N_23190);
nand U25418 (N_25418,N_23881,N_22596);
xnor U25419 (N_25419,N_22911,N_23687);
and U25420 (N_25420,N_23603,N_23398);
nand U25421 (N_25421,N_23563,N_23866);
or U25422 (N_25422,N_22748,N_22630);
nor U25423 (N_25423,N_22956,N_22827);
and U25424 (N_25424,N_23220,N_22702);
xnor U25425 (N_25425,N_22852,N_22811);
nand U25426 (N_25426,N_23821,N_22624);
xor U25427 (N_25427,N_23351,N_22585);
and U25428 (N_25428,N_23055,N_22831);
xor U25429 (N_25429,N_22730,N_23370);
nand U25430 (N_25430,N_23859,N_22974);
xnor U25431 (N_25431,N_23270,N_23783);
nor U25432 (N_25432,N_23329,N_22718);
nor U25433 (N_25433,N_23695,N_23889);
and U25434 (N_25434,N_22721,N_23029);
or U25435 (N_25435,N_23478,N_23870);
and U25436 (N_25436,N_22758,N_23341);
nand U25437 (N_25437,N_23669,N_22559);
nand U25438 (N_25438,N_23775,N_23463);
nand U25439 (N_25439,N_23255,N_23113);
or U25440 (N_25440,N_22995,N_23113);
nand U25441 (N_25441,N_23250,N_23401);
or U25442 (N_25442,N_22819,N_22956);
nor U25443 (N_25443,N_22596,N_23343);
and U25444 (N_25444,N_22852,N_22616);
nor U25445 (N_25445,N_23313,N_23437);
and U25446 (N_25446,N_23289,N_23578);
and U25447 (N_25447,N_22622,N_23460);
xnor U25448 (N_25448,N_23009,N_23400);
nand U25449 (N_25449,N_23563,N_22642);
or U25450 (N_25450,N_22989,N_22622);
nand U25451 (N_25451,N_22560,N_23341);
xor U25452 (N_25452,N_23998,N_23129);
or U25453 (N_25453,N_23846,N_22920);
and U25454 (N_25454,N_22898,N_23792);
nor U25455 (N_25455,N_23277,N_23131);
xnor U25456 (N_25456,N_22688,N_22616);
or U25457 (N_25457,N_23839,N_23961);
and U25458 (N_25458,N_23387,N_23609);
nor U25459 (N_25459,N_23739,N_23236);
xor U25460 (N_25460,N_23582,N_23338);
xnor U25461 (N_25461,N_22670,N_22887);
nand U25462 (N_25462,N_22601,N_23769);
and U25463 (N_25463,N_22606,N_23227);
or U25464 (N_25464,N_23590,N_23319);
and U25465 (N_25465,N_23999,N_23574);
xnor U25466 (N_25466,N_22651,N_22843);
and U25467 (N_25467,N_23955,N_23563);
xor U25468 (N_25468,N_23840,N_23636);
or U25469 (N_25469,N_23198,N_23681);
nor U25470 (N_25470,N_22937,N_22724);
or U25471 (N_25471,N_23837,N_22902);
or U25472 (N_25472,N_23649,N_23533);
or U25473 (N_25473,N_23576,N_22580);
and U25474 (N_25474,N_22673,N_23342);
or U25475 (N_25475,N_22585,N_23026);
xnor U25476 (N_25476,N_22691,N_23570);
or U25477 (N_25477,N_23121,N_22837);
nor U25478 (N_25478,N_22554,N_23152);
nand U25479 (N_25479,N_23487,N_23391);
nand U25480 (N_25480,N_23638,N_22509);
or U25481 (N_25481,N_23080,N_22697);
and U25482 (N_25482,N_23947,N_23945);
or U25483 (N_25483,N_22753,N_22640);
nor U25484 (N_25484,N_23104,N_23354);
or U25485 (N_25485,N_23161,N_23659);
nand U25486 (N_25486,N_23091,N_22758);
and U25487 (N_25487,N_23716,N_22794);
and U25488 (N_25488,N_23389,N_23724);
and U25489 (N_25489,N_22762,N_22668);
xor U25490 (N_25490,N_22676,N_22709);
and U25491 (N_25491,N_22542,N_23515);
or U25492 (N_25492,N_22909,N_22982);
xnor U25493 (N_25493,N_22577,N_22821);
xnor U25494 (N_25494,N_23721,N_23271);
nand U25495 (N_25495,N_22532,N_22720);
nand U25496 (N_25496,N_23274,N_23145);
and U25497 (N_25497,N_22500,N_23149);
nand U25498 (N_25498,N_23517,N_22774);
and U25499 (N_25499,N_23796,N_22832);
xor U25500 (N_25500,N_25041,N_24411);
xnor U25501 (N_25501,N_25263,N_24882);
and U25502 (N_25502,N_24208,N_25007);
and U25503 (N_25503,N_24115,N_24087);
nor U25504 (N_25504,N_24106,N_25028);
and U25505 (N_25505,N_25421,N_24204);
or U25506 (N_25506,N_24852,N_24375);
xor U25507 (N_25507,N_25473,N_24825);
or U25508 (N_25508,N_24335,N_24812);
and U25509 (N_25509,N_24625,N_24448);
and U25510 (N_25510,N_24057,N_25110);
xor U25511 (N_25511,N_24420,N_24754);
and U25512 (N_25512,N_25207,N_25315);
nand U25513 (N_25513,N_24537,N_24376);
nand U25514 (N_25514,N_24191,N_24254);
xnor U25515 (N_25515,N_25155,N_24226);
and U25516 (N_25516,N_24035,N_25309);
nand U25517 (N_25517,N_25039,N_25058);
nand U25518 (N_25518,N_24474,N_25451);
or U25519 (N_25519,N_24171,N_24689);
nand U25520 (N_25520,N_24407,N_24011);
and U25521 (N_25521,N_25407,N_24955);
or U25522 (N_25522,N_25399,N_25459);
xor U25523 (N_25523,N_24258,N_24389);
xor U25524 (N_25524,N_25128,N_24200);
or U25525 (N_25525,N_25241,N_24347);
and U25526 (N_25526,N_25470,N_24378);
xnor U25527 (N_25527,N_24780,N_24172);
nand U25528 (N_25528,N_24458,N_24875);
or U25529 (N_25529,N_24885,N_24518);
or U25530 (N_25530,N_25096,N_24864);
and U25531 (N_25531,N_24862,N_24900);
and U25532 (N_25532,N_24657,N_25308);
nand U25533 (N_25533,N_24583,N_25424);
and U25534 (N_25534,N_24361,N_24710);
xor U25535 (N_25535,N_24270,N_25048);
nor U25536 (N_25536,N_24810,N_24703);
nand U25537 (N_25537,N_25411,N_25192);
xnor U25538 (N_25538,N_24567,N_25419);
or U25539 (N_25539,N_24014,N_25284);
nor U25540 (N_25540,N_24280,N_24205);
nand U25541 (N_25541,N_24715,N_24570);
or U25542 (N_25542,N_24916,N_24666);
nor U25543 (N_25543,N_25291,N_24991);
and U25544 (N_25544,N_24656,N_24445);
and U25545 (N_25545,N_24113,N_24234);
and U25546 (N_25546,N_24117,N_25132);
xnor U25547 (N_25547,N_24696,N_24768);
or U25548 (N_25548,N_24934,N_24738);
nor U25549 (N_25549,N_25295,N_25382);
nand U25550 (N_25550,N_24886,N_24230);
nand U25551 (N_25551,N_24995,N_24690);
and U25552 (N_25552,N_24097,N_24815);
nor U25553 (N_25553,N_24917,N_24433);
or U25554 (N_25554,N_24735,N_25397);
nor U25555 (N_25555,N_24237,N_24473);
and U25556 (N_25556,N_24783,N_24007);
or U25557 (N_25557,N_24125,N_25108);
nor U25558 (N_25558,N_25221,N_24006);
or U25559 (N_25559,N_24156,N_24465);
nand U25560 (N_25560,N_24217,N_24720);
or U25561 (N_25561,N_25133,N_25203);
or U25562 (N_25562,N_25140,N_24248);
nor U25563 (N_25563,N_24358,N_25105);
xor U25564 (N_25564,N_25233,N_25487);
and U25565 (N_25565,N_24085,N_25253);
xor U25566 (N_25566,N_24000,N_24183);
nand U25567 (N_25567,N_25197,N_24450);
xor U25568 (N_25568,N_25498,N_25019);
and U25569 (N_25569,N_25409,N_24813);
nor U25570 (N_25570,N_25301,N_24174);
nor U25571 (N_25571,N_25240,N_24578);
nor U25572 (N_25572,N_24626,N_24364);
and U25573 (N_25573,N_24402,N_24575);
nor U25574 (N_25574,N_25163,N_24419);
and U25575 (N_25575,N_24946,N_24835);
nand U25576 (N_25576,N_24950,N_24043);
xnor U25577 (N_25577,N_24344,N_24553);
and U25578 (N_25578,N_24779,N_25330);
and U25579 (N_25579,N_24409,N_24705);
and U25580 (N_25580,N_24879,N_25341);
or U25581 (N_25581,N_24963,N_24424);
nand U25582 (N_25582,N_25214,N_25115);
nand U25583 (N_25583,N_25224,N_24002);
and U25584 (N_25584,N_25120,N_24966);
nand U25585 (N_25585,N_24773,N_25003);
nor U25586 (N_25586,N_24731,N_24551);
xnor U25587 (N_25587,N_25176,N_24952);
nor U25588 (N_25588,N_24585,N_25478);
or U25589 (N_25589,N_24031,N_24186);
and U25590 (N_25590,N_24076,N_24140);
or U25591 (N_25591,N_25492,N_25405);
or U25592 (N_25592,N_25100,N_24384);
xor U25593 (N_25593,N_24173,N_24515);
or U25594 (N_25594,N_24024,N_24741);
nor U25595 (N_25595,N_25158,N_25320);
xor U25596 (N_25596,N_24047,N_24843);
nand U25597 (N_25597,N_24467,N_25194);
nand U25598 (N_25598,N_24319,N_24541);
nor U25599 (N_25599,N_25325,N_25156);
nor U25600 (N_25600,N_25056,N_24195);
nand U25601 (N_25601,N_25064,N_25204);
or U25602 (N_25602,N_24617,N_24184);
and U25603 (N_25603,N_24032,N_24844);
or U25604 (N_25604,N_25011,N_25212);
or U25605 (N_25605,N_24086,N_24374);
or U25606 (N_25606,N_24522,N_25069);
xor U25607 (N_25607,N_24037,N_24222);
nand U25608 (N_25608,N_25157,N_24382);
nand U25609 (N_25609,N_24777,N_25146);
nand U25610 (N_25610,N_24063,N_24990);
xnor U25611 (N_25611,N_24832,N_24907);
or U25612 (N_25612,N_24277,N_24138);
xnor U25613 (N_25613,N_25305,N_24330);
or U25614 (N_25614,N_24261,N_24748);
nand U25615 (N_25615,N_25274,N_24507);
nor U25616 (N_25616,N_24789,N_24803);
and U25617 (N_25617,N_24760,N_25294);
or U25618 (N_25618,N_24139,N_25228);
or U25619 (N_25619,N_24953,N_25063);
nor U25620 (N_25620,N_24727,N_25261);
or U25621 (N_25621,N_25094,N_24753);
and U25622 (N_25622,N_25017,N_24746);
nor U25623 (N_25623,N_24124,N_24143);
or U25624 (N_25624,N_24912,N_24791);
or U25625 (N_25625,N_25130,N_25489);
nor U25626 (N_25626,N_25098,N_25326);
and U25627 (N_25627,N_25499,N_24324);
nor U25628 (N_25628,N_24153,N_24732);
or U25629 (N_25629,N_24298,N_24496);
or U25630 (N_25630,N_24785,N_24137);
and U25631 (N_25631,N_24476,N_24486);
xor U25632 (N_25632,N_25125,N_25109);
nor U25633 (N_25633,N_24726,N_24333);
nor U25634 (N_25634,N_24978,N_24022);
nor U25635 (N_25635,N_25239,N_24414);
or U25636 (N_25636,N_25112,N_24615);
or U25637 (N_25637,N_24066,N_24708);
xnor U25638 (N_25638,N_24135,N_25392);
nand U25639 (N_25639,N_24463,N_24947);
and U25640 (N_25640,N_24940,N_24469);
xor U25641 (N_25641,N_24893,N_24490);
nor U25642 (N_25642,N_24104,N_25398);
or U25643 (N_25643,N_24502,N_24134);
nor U25644 (N_25644,N_24443,N_25453);
nor U25645 (N_25645,N_25209,N_24697);
and U25646 (N_25646,N_25102,N_25088);
xnor U25647 (N_25647,N_24182,N_24273);
and U25648 (N_25648,N_25393,N_24781);
nand U25649 (N_25649,N_24930,N_24403);
xnor U25650 (N_25650,N_24750,N_24269);
and U25651 (N_25651,N_24221,N_24073);
or U25652 (N_25652,N_24623,N_24488);
or U25653 (N_25653,N_25208,N_24084);
xor U25654 (N_25654,N_24152,N_24788);
nand U25655 (N_25655,N_24634,N_24009);
xnor U25656 (N_25656,N_25321,N_24307);
xor U25657 (N_25657,N_24552,N_24455);
and U25658 (N_25658,N_24704,N_24508);
nor U25659 (N_25659,N_25307,N_25450);
nor U25660 (N_25660,N_24246,N_25496);
nand U25661 (N_25661,N_24729,N_25055);
or U25662 (N_25662,N_24056,N_24480);
xnor U25663 (N_25663,N_24004,N_24855);
nand U25664 (N_25664,N_24906,N_25380);
or U25665 (N_25665,N_25304,N_24225);
nor U25666 (N_25666,N_24533,N_24756);
xnor U25667 (N_25667,N_24516,N_24668);
nor U25668 (N_25668,N_24380,N_24514);
nand U25669 (N_25669,N_25036,N_24430);
and U25670 (N_25670,N_25329,N_25099);
or U25671 (N_25671,N_24888,N_24805);
xor U25672 (N_25672,N_24994,N_24680);
nor U25673 (N_25673,N_24663,N_25089);
nand U25674 (N_25674,N_24556,N_24510);
xnor U25675 (N_25675,N_25237,N_24446);
xnor U25676 (N_25676,N_24249,N_24099);
nand U25677 (N_25677,N_24980,N_24046);
nand U25678 (N_25678,N_25455,N_24044);
or U25679 (N_25679,N_24078,N_24013);
xor U25680 (N_25680,N_24581,N_24877);
xor U25681 (N_25681,N_25369,N_24158);
nor U25682 (N_25682,N_25364,N_25231);
nand U25683 (N_25683,N_25383,N_24539);
xnor U25684 (N_25684,N_24718,N_24896);
nand U25685 (N_25685,N_24199,N_25236);
xnor U25686 (N_25686,N_25012,N_24653);
nand U25687 (N_25687,N_24986,N_25436);
and U25688 (N_25688,N_24602,N_25288);
nand U25689 (N_25689,N_24390,N_25227);
nand U25690 (N_25690,N_24712,N_25185);
nand U25691 (N_25691,N_24157,N_25287);
and U25692 (N_25692,N_24304,N_24256);
nor U25693 (N_25693,N_24548,N_24644);
xnor U25694 (N_25694,N_24426,N_24381);
and U25695 (N_25695,N_24513,N_24436);
nand U25696 (N_25696,N_24880,N_24674);
or U25697 (N_25697,N_24968,N_25493);
or U25698 (N_25698,N_24149,N_25034);
nand U25699 (N_25699,N_24650,N_24495);
nand U25700 (N_25700,N_24100,N_24758);
nand U25701 (N_25701,N_24054,N_24931);
nor U25702 (N_25702,N_24064,N_24599);
nor U25703 (N_25703,N_24676,N_24449);
nand U25704 (N_25704,N_24560,N_24102);
or U25705 (N_25705,N_24036,N_25202);
and U25706 (N_25706,N_25442,N_24829);
or U25707 (N_25707,N_25182,N_24903);
xnor U25708 (N_25708,N_24971,N_24216);
and U25709 (N_25709,N_25427,N_24196);
and U25710 (N_25710,N_25116,N_24315);
or U25711 (N_25711,N_24224,N_24105);
nand U25712 (N_25712,N_24238,N_25190);
and U25713 (N_25713,N_24526,N_24373);
nor U25714 (N_25714,N_25279,N_25218);
xnor U25715 (N_25715,N_24147,N_25251);
xnor U25716 (N_25716,N_24489,N_24253);
nand U25717 (N_25717,N_24299,N_25068);
and U25718 (N_25718,N_24154,N_25013);
or U25719 (N_25719,N_25257,N_24811);
xnor U25720 (N_25720,N_24681,N_24547);
and U25721 (N_25721,N_25004,N_24500);
and U25722 (N_25722,N_25177,N_24637);
and U25723 (N_25723,N_25490,N_25484);
nor U25724 (N_25724,N_24027,N_25440);
xnor U25725 (N_25725,N_25254,N_25142);
nor U25726 (N_25726,N_25074,N_24889);
nor U25727 (N_25727,N_24597,N_25345);
xnor U25728 (N_25728,N_24564,N_24636);
nor U25729 (N_25729,N_24447,N_24770);
or U25730 (N_25730,N_25352,N_24053);
nor U25731 (N_25731,N_24241,N_24632);
nand U25732 (N_25732,N_25370,N_24456);
or U25733 (N_25733,N_24606,N_24853);
nand U25734 (N_25734,N_25250,N_24782);
xnor U25735 (N_25735,N_24122,N_24136);
or U25736 (N_25736,N_25414,N_24268);
and U25737 (N_25737,N_24316,N_24391);
nand U25738 (N_25738,N_25181,N_24610);
xnor U25739 (N_25739,N_25277,N_24609);
nand U25740 (N_25740,N_24638,N_25358);
and U25741 (N_25741,N_24410,N_25186);
nand U25742 (N_25742,N_24519,N_24318);
and U25743 (N_25743,N_25081,N_24709);
nand U25744 (N_25744,N_25438,N_24017);
or U25745 (N_25745,N_24658,N_25077);
nand U25746 (N_25746,N_24454,N_24179);
nor U25747 (N_25747,N_25445,N_24714);
nand U25748 (N_25748,N_24821,N_25435);
and U25749 (N_25749,N_24052,N_24142);
nand U25750 (N_25750,N_25022,N_25354);
or U25751 (N_25751,N_24935,N_24568);
or U25752 (N_25752,N_24793,N_24151);
xnor U25753 (N_25753,N_24349,N_24123);
nand U25754 (N_25754,N_25126,N_24611);
and U25755 (N_25755,N_24841,N_25335);
nand U25756 (N_25756,N_25373,N_24543);
nor U25757 (N_25757,N_24594,N_24098);
xor U25758 (N_25758,N_24354,N_25031);
or U25759 (N_25759,N_24028,N_25160);
nand U25760 (N_25760,N_25395,N_24601);
or U25761 (N_25761,N_25443,N_25401);
xor U25762 (N_25762,N_24648,N_25293);
xor U25763 (N_25763,N_25374,N_24283);
or U25764 (N_25764,N_24981,N_25183);
nor U25765 (N_25765,N_25016,N_24752);
or U25766 (N_25766,N_24742,N_24440);
nor U25767 (N_25767,N_25310,N_25477);
and U25768 (N_25768,N_24997,N_24313);
nand U25769 (N_25769,N_24908,N_24187);
nand U25770 (N_25770,N_24826,N_24992);
and U25771 (N_25771,N_24540,N_25171);
and U25772 (N_25772,N_24818,N_24328);
or U25773 (N_25773,N_24077,N_24506);
or U25774 (N_25774,N_25365,N_25479);
nor U25775 (N_25775,N_24849,N_24796);
or U25776 (N_25776,N_24736,N_24161);
nor U25777 (N_25777,N_25333,N_24635);
or U25778 (N_25778,N_25215,N_24572);
or U25779 (N_25779,N_25150,N_24262);
xor U25780 (N_25780,N_25093,N_25408);
nor U25781 (N_25781,N_24901,N_24275);
xor U25782 (N_25782,N_25006,N_24008);
or U25783 (N_25783,N_24170,N_24475);
and U25784 (N_25784,N_25466,N_25226);
xor U25785 (N_25785,N_24688,N_25360);
xnor U25786 (N_25786,N_24942,N_25191);
nor U25787 (N_25787,N_24959,N_24020);
or U25788 (N_25788,N_24193,N_25119);
nor U25789 (N_25789,N_24614,N_24695);
or U25790 (N_25790,N_25047,N_24795);
and U25791 (N_25791,N_24131,N_24645);
nand U25792 (N_25792,N_25151,N_24197);
nor U25793 (N_25793,N_24797,N_24383);
nand U25794 (N_25794,N_25273,N_25271);
or U25795 (N_25795,N_25113,N_24034);
and U25796 (N_25796,N_24385,N_24452);
or U25797 (N_25797,N_25400,N_24462);
nor U25798 (N_25798,N_24080,N_24194);
nor U25799 (N_25799,N_24178,N_24786);
xor U25800 (N_25800,N_25137,N_24622);
xor U25801 (N_25801,N_24972,N_24661);
or U25802 (N_25802,N_24512,N_24218);
and U25803 (N_25803,N_25319,N_24744);
nand U25804 (N_25804,N_24929,N_25317);
or U25805 (N_25805,N_24989,N_25061);
or U25806 (N_25806,N_24001,N_25043);
or U25807 (N_25807,N_25059,N_24295);
or U25808 (N_25808,N_24557,N_24925);
and U25809 (N_25809,N_24827,N_24817);
or U25810 (N_25810,N_25302,N_24481);
nand U25811 (N_25811,N_25118,N_24483);
or U25812 (N_25812,N_24881,N_24075);
nand U25813 (N_25813,N_24251,N_24743);
and U25814 (N_25814,N_25070,N_24279);
or U25815 (N_25815,N_24721,N_25002);
nor U25816 (N_25816,N_24621,N_24717);
xor U25817 (N_25817,N_24713,N_25472);
or U25818 (N_25818,N_24033,N_24214);
nor U25819 (N_25819,N_24285,N_24363);
nand U25820 (N_25820,N_24913,N_25327);
or U25821 (N_25821,N_24902,N_24954);
and U25822 (N_25822,N_24867,N_25027);
nor U25823 (N_25823,N_25334,N_24869);
xnor U25824 (N_25824,N_24386,N_25195);
xor U25825 (N_25825,N_25362,N_24745);
nand U25826 (N_25826,N_24071,N_24023);
or U25827 (N_25827,N_24229,N_24305);
nand U25828 (N_25828,N_24607,N_24937);
nand U25829 (N_25829,N_25269,N_24492);
or U25830 (N_25830,N_24207,N_24272);
or U25831 (N_25831,N_24212,N_24164);
and U25832 (N_25832,N_24163,N_24461);
and U25833 (N_25833,N_25467,N_25020);
nand U25834 (N_25834,N_24800,N_24370);
nor U25835 (N_25835,N_24976,N_24350);
nand U25836 (N_25836,N_24175,N_25439);
nor U25837 (N_25837,N_24276,N_25391);
and U25838 (N_25838,N_24868,N_24112);
or U25839 (N_25839,N_24856,N_24220);
and U25840 (N_25840,N_24072,N_24751);
and U25841 (N_25841,N_24274,N_25429);
or U25842 (N_25842,N_24639,N_24352);
nor U25843 (N_25843,N_24939,N_25332);
or U25844 (N_25844,N_24979,N_24554);
nand U25845 (N_25845,N_24357,N_24400);
or U25846 (N_25846,N_24192,N_24616);
and U25847 (N_25847,N_24682,N_24851);
nand U25848 (N_25848,N_25187,N_24612);
and U25849 (N_25849,N_24282,N_25394);
nor U25850 (N_25850,N_24593,N_24630);
nor U25851 (N_25851,N_24517,N_24684);
xor U25852 (N_25852,N_25091,N_24442);
nor U25853 (N_25853,N_24365,N_24778);
or U25854 (N_25854,N_25433,N_24049);
xor U25855 (N_25855,N_24228,N_24126);
xor U25856 (N_25856,N_25147,N_25344);
or U25857 (N_25857,N_24905,N_25458);
xnor U25858 (N_25858,N_24546,N_25430);
or U25859 (N_25859,N_25080,N_24339);
and U25860 (N_25860,N_24730,N_24484);
nor U25861 (N_25861,N_24168,N_25406);
nor U25862 (N_25862,N_24620,N_24911);
xor U25863 (N_25863,N_25052,N_24493);
nand U25864 (N_25864,N_24891,N_24120);
nand U25865 (N_25865,N_24421,N_24595);
xor U25866 (N_25866,N_24863,N_24871);
and U25867 (N_25867,N_25270,N_24244);
nand U25868 (N_25868,N_25050,N_25454);
and U25869 (N_25869,N_25139,N_24948);
nand U25870 (N_25870,N_24904,N_25145);
nor U25871 (N_25871,N_24922,N_24956);
and U25872 (N_25872,N_24814,N_25338);
nand U25873 (N_25873,N_24858,N_24651);
nor U25874 (N_25874,N_24497,N_24866);
nand U25875 (N_25875,N_24065,N_25377);
and U25876 (N_25876,N_25322,N_24289);
nor U25877 (N_25877,N_24505,N_24015);
or U25878 (N_25878,N_25425,N_25343);
or U25879 (N_25879,N_24413,N_24340);
xnor U25880 (N_25880,N_24165,N_24263);
nand U25881 (N_25881,N_25372,N_24998);
and U25882 (N_25882,N_24771,N_24159);
xnor U25883 (N_25883,N_24603,N_24774);
and U25884 (N_25884,N_24592,N_24790);
xor U25885 (N_25885,N_24441,N_24050);
nor U25886 (N_25886,N_24404,N_25117);
or U25887 (N_25887,N_24118,N_24395);
nor U25888 (N_25888,N_25351,N_24042);
nand U25889 (N_25889,N_25432,N_25278);
and U25890 (N_25890,N_24103,N_25087);
nand U25891 (N_25891,N_24831,N_24737);
nand U25892 (N_25892,N_25211,N_24130);
xnor U25893 (N_25893,N_24646,N_25229);
and U25894 (N_25894,N_25386,N_24576);
xor U25895 (N_25895,N_24081,N_24571);
and U25896 (N_25896,N_25260,N_24687);
nor U25897 (N_25897,N_25054,N_24041);
nor U25898 (N_25898,N_25078,N_24026);
or U25899 (N_25899,N_24949,N_25086);
or U25900 (N_25900,N_24683,N_24327);
and U25901 (N_25901,N_25285,N_24189);
nand U25902 (N_25902,N_24146,N_24619);
and U25903 (N_25903,N_24794,N_25303);
and U25904 (N_25904,N_25359,N_25248);
and U25905 (N_25905,N_25385,N_24392);
nor U25906 (N_25906,N_24673,N_24494);
nor U25907 (N_25907,N_24860,N_25384);
or U25908 (N_25908,N_24999,N_25213);
nand U25909 (N_25909,N_24962,N_24671);
xnor U25910 (N_25910,N_24288,N_24890);
xnor U25911 (N_25911,N_24351,N_24366);
nand U25912 (N_25912,N_25463,N_24740);
or U25913 (N_25913,N_24247,N_24589);
nor U25914 (N_25914,N_24569,N_25420);
or U25915 (N_25915,N_24405,N_25154);
nand U25916 (N_25916,N_25410,N_24162);
and U25917 (N_25917,N_25388,N_24150);
and U25918 (N_25918,N_24439,N_24491);
xnor U25919 (N_25919,N_25245,N_24346);
nand U25920 (N_25920,N_25434,N_24565);
nand U25921 (N_25921,N_24088,N_24309);
nand U25922 (N_25922,N_25378,N_24969);
nand U25923 (N_25923,N_24355,N_25053);
and U25924 (N_25924,N_24498,N_25348);
nand U25925 (N_25925,N_24215,N_24836);
xor U25926 (N_25926,N_24928,N_25210);
nor U25927 (N_25927,N_24362,N_24096);
or U25928 (N_25928,N_25252,N_25084);
and U25929 (N_25929,N_24764,N_24711);
or U25930 (N_25930,N_24914,N_25174);
nor U25931 (N_25931,N_24242,N_25180);
and U25932 (N_25932,N_24647,N_24719);
xnor U25933 (N_25933,N_24865,N_25103);
or U25934 (N_25934,N_24534,N_25491);
and U25935 (N_25935,N_25312,N_24763);
nor U25936 (N_25936,N_24530,N_25244);
nand U25937 (N_25937,N_24308,N_24201);
xnor U25938 (N_25938,N_24377,N_24642);
nand U25939 (N_25939,N_24932,N_24368);
nand U25940 (N_25940,N_25015,N_25247);
or U25941 (N_25941,N_24640,N_24190);
xor U25942 (N_25942,N_24883,N_25044);
xor U25943 (N_25943,N_24089,N_24051);
xnor U25944 (N_25944,N_25161,N_25350);
nor U25945 (N_25945,N_24334,N_24723);
nor U25946 (N_25946,N_25469,N_24499);
nand U25947 (N_25947,N_24114,N_24550);
xor U25948 (N_25948,N_24109,N_24698);
nand U25949 (N_25949,N_25413,N_24988);
and U25950 (N_25950,N_25051,N_24665);
or U25951 (N_25951,N_24091,N_24655);
or U25952 (N_25952,N_24082,N_25040);
nand U25953 (N_25953,N_25465,N_25353);
or U25954 (N_25954,N_24679,N_25494);
and U25955 (N_25955,N_25232,N_24255);
nand U25956 (N_25956,N_24700,N_25188);
xnor U25957 (N_25957,N_25485,N_24416);
and U25958 (N_25958,N_24107,N_24025);
or U25959 (N_25959,N_24633,N_24321);
and U25960 (N_25960,N_25106,N_24982);
nand U25961 (N_25961,N_24188,N_24466);
xnor U25962 (N_25962,N_24101,N_24177);
and U25963 (N_25963,N_24240,N_24899);
nand U25964 (N_25964,N_25045,N_24521);
or U25965 (N_25965,N_24210,N_24387);
nor U25966 (N_25966,N_24290,N_24167);
xnor U25967 (N_25967,N_24524,N_24320);
and U25968 (N_25968,N_24437,N_25206);
nor U25969 (N_25969,N_25217,N_24757);
nand U25970 (N_25970,N_25495,N_25090);
nor U25971 (N_25971,N_24322,N_24343);
or U25972 (N_25972,N_24772,N_25238);
or U25973 (N_25973,N_25066,N_24920);
or U25974 (N_25974,N_25342,N_24692);
nor U25975 (N_25975,N_24643,N_24525);
nor U25976 (N_25976,N_24176,N_24974);
and U25977 (N_25977,N_25124,N_25286);
nor U25978 (N_25978,N_24435,N_24964);
nand U25979 (N_25979,N_24252,N_24667);
nand U25980 (N_25980,N_24591,N_24544);
or U25981 (N_25981,N_24271,N_25272);
nor U25982 (N_25982,N_24074,N_24693);
nand U25983 (N_25983,N_24694,N_25402);
nor U25984 (N_25984,N_24873,N_25023);
or U25985 (N_25985,N_25037,N_24686);
nor U25986 (N_25986,N_24629,N_25468);
xnor U25987 (N_25987,N_25258,N_24977);
and U25988 (N_25988,N_24965,N_25035);
and U25989 (N_25989,N_24444,N_24691);
nor U25990 (N_25990,N_24945,N_24807);
and U25991 (N_25991,N_24501,N_24582);
nand U25992 (N_25992,N_24432,N_24798);
nor U25993 (N_25993,N_25355,N_25159);
nor U25994 (N_25994,N_24527,N_24231);
and U25995 (N_25995,N_24503,N_24846);
and U25996 (N_25996,N_24477,N_25135);
nand U25997 (N_25997,N_24876,N_24749);
nand U25998 (N_25998,N_24070,N_25416);
nand U25999 (N_25999,N_24040,N_24417);
or U26000 (N_26000,N_24039,N_25281);
nand U26001 (N_26001,N_24434,N_25431);
nor U26002 (N_26002,N_25446,N_25363);
and U26003 (N_26003,N_24127,N_25357);
nor U26004 (N_26004,N_25107,N_24281);
or U26005 (N_26005,N_24702,N_24213);
xnor U26006 (N_26006,N_25390,N_24233);
and U26007 (N_26007,N_25331,N_24747);
nor U26008 (N_26008,N_24600,N_24260);
and U26009 (N_26009,N_24535,N_24975);
and U26010 (N_26010,N_24145,N_24232);
nand U26011 (N_26011,N_25033,N_25141);
or U26012 (N_26012,N_25220,N_24329);
nand U26013 (N_26013,N_24379,N_25417);
xor U26014 (N_26014,N_25111,N_24523);
nor U26015 (N_26015,N_25426,N_24759);
nor U26016 (N_26016,N_24840,N_24311);
nand U26017 (N_26017,N_24816,N_24755);
xnor U26018 (N_26018,N_24010,N_24628);
nand U26019 (N_26019,N_25375,N_24286);
nor U26020 (N_26020,N_24418,N_24326);
nor U26021 (N_26021,N_25179,N_24878);
nand U26022 (N_26022,N_24678,N_24408);
xor U26023 (N_26023,N_24306,N_25461);
nor U26024 (N_26024,N_25296,N_25057);
or U26025 (N_26025,N_24587,N_24345);
xnor U26026 (N_26026,N_24284,N_24921);
or U26027 (N_26027,N_24003,N_25367);
xor U26028 (N_26028,N_24970,N_24509);
nor U26029 (N_26029,N_24808,N_24068);
nor U26030 (N_26030,N_25104,N_25437);
or U26031 (N_26031,N_24021,N_24579);
or U26032 (N_26032,N_24059,N_25201);
xnor U26033 (N_26033,N_24093,N_25222);
and U26034 (N_26034,N_25403,N_24520);
nor U26035 (N_26035,N_25422,N_25184);
nor U26036 (N_26036,N_25482,N_25488);
or U26037 (N_26037,N_24649,N_25025);
xor U26038 (N_26038,N_24266,N_24367);
nand U26039 (N_26039,N_24300,N_25131);
and U26040 (N_26040,N_25318,N_24631);
xor U26041 (N_26041,N_24353,N_24919);
or U26042 (N_26042,N_24590,N_24180);
xnor U26043 (N_26043,N_24148,N_24401);
nor U26044 (N_26044,N_24938,N_24422);
nor U26045 (N_26045,N_25148,N_25166);
nand U26046 (N_26046,N_25021,N_25010);
xnor U26047 (N_26047,N_24427,N_25356);
or U26048 (N_26048,N_24801,N_24119);
or U26049 (N_26049,N_24819,N_25134);
xnor U26050 (N_26050,N_25167,N_24675);
and U26051 (N_26051,N_25046,N_24062);
or U26052 (N_26052,N_25480,N_24973);
xnor U26053 (N_26053,N_24239,N_24734);
or U26054 (N_26054,N_24331,N_24652);
nand U26055 (N_26055,N_24944,N_24121);
nand U26056 (N_26056,N_25387,N_24399);
xnor U26057 (N_26057,N_24356,N_25256);
or U26058 (N_26058,N_24838,N_25379);
or U26059 (N_26059,N_25144,N_24834);
and U26060 (N_26060,N_24128,N_24155);
nand U26061 (N_26061,N_24532,N_24895);
and U26062 (N_26062,N_24198,N_25276);
nor U26063 (N_26063,N_24301,N_24012);
and U26064 (N_26064,N_24018,N_25200);
or U26065 (N_26065,N_24393,N_25075);
or U26066 (N_26066,N_24485,N_25381);
and U26067 (N_26067,N_25225,N_24314);
and U26068 (N_26068,N_24542,N_24397);
xor U26069 (N_26069,N_24428,N_25173);
nor U26070 (N_26070,N_24048,N_24848);
and U26071 (N_26071,N_24769,N_24111);
nand U26072 (N_26072,N_25457,N_25418);
and U26073 (N_26073,N_25024,N_24574);
and U26074 (N_26074,N_24453,N_24809);
or U26075 (N_26075,N_25018,N_25030);
nand U26076 (N_26076,N_25483,N_25230);
nand U26077 (N_26077,N_24596,N_24884);
or U26078 (N_26078,N_24060,N_24278);
nand U26079 (N_26079,N_24479,N_25072);
nor U26080 (N_26080,N_25283,N_25198);
and U26081 (N_26081,N_24406,N_25079);
nand U26082 (N_26082,N_25164,N_24799);
nand U26083 (N_26083,N_24996,N_25481);
or U26084 (N_26084,N_25267,N_24325);
and U26085 (N_26085,N_24806,N_24926);
nor U26086 (N_26086,N_24487,N_24613);
nor U26087 (N_26087,N_24478,N_24960);
xor U26088 (N_26088,N_24894,N_24608);
or U26089 (N_26089,N_25193,N_24257);
xor U26090 (N_26090,N_24029,N_25337);
or U26091 (N_26091,N_24303,N_24584);
xor U26092 (N_26092,N_24095,N_25129);
and U26093 (N_26093,N_25062,N_24872);
xor U26094 (N_26094,N_24677,N_25415);
nand U26095 (N_26095,N_25199,N_24264);
and U26096 (N_26096,N_25292,N_25092);
or U26097 (N_26097,N_25205,N_25280);
xor U26098 (N_26098,N_24055,N_24472);
xor U26099 (N_26099,N_25474,N_25101);
nor U26100 (N_26100,N_24845,N_24558);
xnor U26101 (N_26101,N_24776,N_24369);
nor U26102 (N_26102,N_24967,N_24765);
xnor U26103 (N_26103,N_24341,N_24699);
and U26104 (N_26104,N_24297,N_25340);
or U26105 (N_26105,N_24559,N_25376);
nand U26106 (N_26106,N_25014,N_25123);
nor U26107 (N_26107,N_25475,N_25042);
nor U26108 (N_26108,N_24654,N_25152);
and U26109 (N_26109,N_25169,N_24209);
nor U26110 (N_26110,N_24739,N_25289);
nand U26111 (N_26111,N_24562,N_24429);
nor U26112 (N_26112,N_24957,N_24360);
nand U26113 (N_26113,N_24566,N_24371);
and U26114 (N_26114,N_24061,N_24604);
and U26115 (N_26115,N_24861,N_25471);
and U26116 (N_26116,N_25347,N_24983);
nand U26117 (N_26117,N_24415,N_24824);
xnor U26118 (N_26118,N_25121,N_25371);
xor U26119 (N_26119,N_24019,N_24659);
nand U26120 (N_26120,N_25366,N_24468);
nand U26121 (N_26121,N_25265,N_25114);
xor U26122 (N_26122,N_25000,N_25298);
or U26123 (N_26123,N_24332,N_25026);
nand U26124 (N_26124,N_24669,N_25009);
xnor U26125 (N_26125,N_24586,N_24372);
or U26126 (N_26126,N_24211,N_24850);
nand U26127 (N_26127,N_24067,N_24618);
xor U26128 (N_26128,N_24511,N_24302);
and U26129 (N_26129,N_24203,N_24092);
nand U26130 (N_26130,N_24605,N_25153);
nand U26131 (N_26131,N_24830,N_24038);
xor U26132 (N_26132,N_25246,N_24722);
and U26133 (N_26133,N_25235,N_24538);
and U26134 (N_26134,N_25178,N_24094);
xor U26135 (N_26135,N_24822,N_24005);
nor U26136 (N_26136,N_24144,N_25032);
nor U26137 (N_26137,N_25449,N_24292);
xnor U26138 (N_26138,N_24804,N_24662);
nor U26139 (N_26139,N_25095,N_24293);
xnor U26140 (N_26140,N_24396,N_24108);
xnor U26141 (N_26141,N_25464,N_24359);
nand U26142 (N_26142,N_25242,N_24431);
nand U26143 (N_26143,N_25486,N_24857);
nor U26144 (N_26144,N_25143,N_24141);
nand U26145 (N_26145,N_25085,N_24859);
or U26146 (N_26146,N_25172,N_25175);
nor U26147 (N_26147,N_25300,N_24936);
nor U26148 (N_26148,N_24243,N_25462);
nand U26149 (N_26149,N_24219,N_25249);
nand U26150 (N_26150,N_24181,N_25259);
or U26151 (N_26151,N_24090,N_25067);
and U26152 (N_26152,N_24660,N_25389);
nand U26153 (N_26153,N_24470,N_25262);
xor U26154 (N_26154,N_24030,N_25361);
nand U26155 (N_26155,N_25029,N_24250);
or U26156 (N_26156,N_24707,N_24531);
and U26157 (N_26157,N_24069,N_25008);
or U26158 (N_26158,N_25299,N_25122);
nor U26159 (N_26159,N_24580,N_24423);
xor U26160 (N_26160,N_24943,N_25127);
nand U26161 (N_26161,N_24129,N_24338);
xor U26162 (N_26162,N_25149,N_24733);
and U26163 (N_26163,N_25328,N_24169);
nor U26164 (N_26164,N_24624,N_24312);
xnor U26165 (N_26165,N_24854,N_25136);
or U26166 (N_26166,N_24762,N_25268);
or U26167 (N_26167,N_24045,N_24887);
xor U26168 (N_26168,N_25165,N_24504);
nand U26169 (N_26169,N_24460,N_24412);
or U26170 (N_26170,N_24438,N_24236);
and U26171 (N_26171,N_24259,N_25266);
nand U26172 (N_26172,N_24573,N_24529);
nand U26173 (N_26173,N_25255,N_25404);
and U26174 (N_26174,N_25368,N_24820);
or U26175 (N_26175,N_24116,N_25323);
and U26176 (N_26176,N_24482,N_24915);
and U26177 (N_26177,N_24227,N_25316);
or U26178 (N_26178,N_24348,N_24837);
and U26179 (N_26179,N_24701,N_24728);
or U26180 (N_26180,N_25339,N_25349);
and U26181 (N_26181,N_25336,N_25452);
nor U26182 (N_26182,N_24464,N_24588);
xnor U26183 (N_26183,N_24987,N_24909);
nor U26184 (N_26184,N_24310,N_24235);
xor U26185 (N_26185,N_25264,N_24563);
or U26186 (N_26186,N_25297,N_25189);
xnor U26187 (N_26187,N_24951,N_25065);
and U26188 (N_26188,N_24958,N_24898);
or U26189 (N_26189,N_25412,N_24627);
xnor U26190 (N_26190,N_24874,N_24294);
nand U26191 (N_26191,N_24941,N_25168);
xnor U26192 (N_26192,N_24425,N_24058);
or U26193 (N_26193,N_24536,N_24457);
and U26194 (N_26194,N_24083,N_25076);
xnor U26195 (N_26195,N_24296,N_25219);
nand U26196 (N_26196,N_24870,N_24185);
nor U26197 (N_26197,N_24725,N_24555);
xnor U26198 (N_26198,N_25243,N_25314);
xnor U26199 (N_26199,N_24337,N_24918);
nor U26200 (N_26200,N_24766,N_24923);
or U26201 (N_26201,N_25346,N_24839);
nand U26202 (N_26202,N_24847,N_24761);
nor U26203 (N_26203,N_24897,N_25423);
nand U26204 (N_26204,N_25476,N_25456);
nand U26205 (N_26205,N_25448,N_24823);
nand U26206 (N_26206,N_24336,N_25223);
nand U26207 (N_26207,N_25396,N_24892);
nor U26208 (N_26208,N_24160,N_24398);
or U26209 (N_26209,N_25311,N_24561);
nor U26210 (N_26210,N_24842,N_24287);
xnor U26211 (N_26211,N_24223,N_25097);
nor U26212 (N_26212,N_25275,N_24927);
nor U26213 (N_26213,N_24265,N_24598);
xnor U26214 (N_26214,N_25447,N_24166);
nand U26215 (N_26215,N_24079,N_25428);
nor U26216 (N_26216,N_24016,N_25162);
xnor U26217 (N_26217,N_25282,N_24672);
nor U26218 (N_26218,N_25060,N_25313);
nor U26219 (N_26219,N_24110,N_24545);
or U26220 (N_26220,N_24724,N_25071);
and U26221 (N_26221,N_24664,N_25049);
nor U26222 (N_26222,N_24706,N_24342);
or U26223 (N_26223,N_24291,N_24451);
or U26224 (N_26224,N_24132,N_24206);
xor U26225 (N_26225,N_24775,N_25497);
xor U26226 (N_26226,N_25005,N_24267);
nand U26227 (N_26227,N_25196,N_24716);
and U26228 (N_26228,N_24577,N_24985);
nor U26229 (N_26229,N_25444,N_25234);
and U26230 (N_26230,N_25324,N_24202);
nor U26231 (N_26231,N_24787,N_24528);
or U26232 (N_26232,N_25170,N_25441);
and U26233 (N_26233,N_24910,N_24641);
or U26234 (N_26234,N_24984,N_25138);
or U26235 (N_26235,N_24792,N_24394);
and U26236 (N_26236,N_24388,N_24924);
nor U26237 (N_26237,N_25073,N_25290);
and U26238 (N_26238,N_25082,N_24993);
and U26239 (N_26239,N_25216,N_24685);
nor U26240 (N_26240,N_24133,N_24828);
xor U26241 (N_26241,N_25306,N_24784);
nand U26242 (N_26242,N_24549,N_25460);
or U26243 (N_26243,N_24802,N_24833);
nand U26244 (N_26244,N_25083,N_24317);
or U26245 (N_26245,N_24767,N_24459);
or U26246 (N_26246,N_24323,N_24245);
nand U26247 (N_26247,N_24670,N_24933);
nand U26248 (N_26248,N_24471,N_25038);
nor U26249 (N_26249,N_24961,N_25001);
or U26250 (N_26250,N_24353,N_24983);
and U26251 (N_26251,N_25324,N_24621);
or U26252 (N_26252,N_24013,N_24663);
or U26253 (N_26253,N_24497,N_24659);
xor U26254 (N_26254,N_24706,N_24639);
and U26255 (N_26255,N_25425,N_24993);
nor U26256 (N_26256,N_24397,N_25175);
nor U26257 (N_26257,N_24965,N_24328);
and U26258 (N_26258,N_25291,N_24081);
nor U26259 (N_26259,N_25441,N_25200);
or U26260 (N_26260,N_24955,N_25444);
and U26261 (N_26261,N_25020,N_24383);
nand U26262 (N_26262,N_24658,N_24977);
or U26263 (N_26263,N_24466,N_24766);
xor U26264 (N_26264,N_24683,N_25002);
xor U26265 (N_26265,N_25457,N_24048);
or U26266 (N_26266,N_25175,N_25123);
xor U26267 (N_26267,N_24654,N_24931);
xor U26268 (N_26268,N_24430,N_24411);
and U26269 (N_26269,N_25275,N_25175);
nand U26270 (N_26270,N_24735,N_24080);
nand U26271 (N_26271,N_24521,N_24353);
nor U26272 (N_26272,N_24183,N_24120);
or U26273 (N_26273,N_25233,N_24734);
xor U26274 (N_26274,N_25154,N_25203);
xnor U26275 (N_26275,N_24277,N_24038);
nor U26276 (N_26276,N_25260,N_24389);
and U26277 (N_26277,N_25254,N_25132);
nor U26278 (N_26278,N_24153,N_25258);
and U26279 (N_26279,N_24486,N_24908);
or U26280 (N_26280,N_25346,N_24525);
xnor U26281 (N_26281,N_25108,N_25436);
xnor U26282 (N_26282,N_24467,N_24261);
nor U26283 (N_26283,N_24950,N_25334);
xor U26284 (N_26284,N_25412,N_24249);
nand U26285 (N_26285,N_24810,N_25027);
nand U26286 (N_26286,N_24965,N_24443);
nor U26287 (N_26287,N_24337,N_25227);
and U26288 (N_26288,N_24054,N_25248);
xnor U26289 (N_26289,N_24866,N_25107);
or U26290 (N_26290,N_25421,N_24501);
nand U26291 (N_26291,N_24422,N_24995);
and U26292 (N_26292,N_25400,N_24078);
xor U26293 (N_26293,N_24516,N_24128);
nand U26294 (N_26294,N_25348,N_24171);
xor U26295 (N_26295,N_25226,N_25235);
xor U26296 (N_26296,N_24362,N_24496);
or U26297 (N_26297,N_25056,N_24521);
xnor U26298 (N_26298,N_24130,N_25050);
xor U26299 (N_26299,N_24832,N_24496);
and U26300 (N_26300,N_24211,N_24454);
nand U26301 (N_26301,N_24014,N_25343);
and U26302 (N_26302,N_25286,N_24845);
nor U26303 (N_26303,N_24384,N_24497);
nand U26304 (N_26304,N_25248,N_24791);
xnor U26305 (N_26305,N_24302,N_25344);
or U26306 (N_26306,N_25260,N_25326);
nand U26307 (N_26307,N_24793,N_24772);
and U26308 (N_26308,N_25256,N_24258);
or U26309 (N_26309,N_24705,N_25261);
or U26310 (N_26310,N_25035,N_25088);
nand U26311 (N_26311,N_24642,N_24206);
nand U26312 (N_26312,N_25116,N_25272);
or U26313 (N_26313,N_24363,N_24375);
nor U26314 (N_26314,N_25302,N_24513);
nor U26315 (N_26315,N_25035,N_24953);
nand U26316 (N_26316,N_25429,N_24443);
xor U26317 (N_26317,N_24125,N_24187);
nand U26318 (N_26318,N_24078,N_25111);
nor U26319 (N_26319,N_24164,N_24800);
nand U26320 (N_26320,N_24036,N_25423);
nand U26321 (N_26321,N_24320,N_24050);
xor U26322 (N_26322,N_24143,N_25433);
or U26323 (N_26323,N_24840,N_24638);
nand U26324 (N_26324,N_24067,N_24881);
and U26325 (N_26325,N_24401,N_24732);
or U26326 (N_26326,N_24447,N_25191);
and U26327 (N_26327,N_24239,N_25276);
xor U26328 (N_26328,N_24616,N_24383);
and U26329 (N_26329,N_24875,N_24775);
nor U26330 (N_26330,N_25162,N_24704);
xor U26331 (N_26331,N_24987,N_24824);
or U26332 (N_26332,N_25414,N_24274);
xor U26333 (N_26333,N_24507,N_24289);
xnor U26334 (N_26334,N_25265,N_25075);
nor U26335 (N_26335,N_24012,N_24879);
xnor U26336 (N_26336,N_24091,N_24949);
nor U26337 (N_26337,N_24289,N_25120);
nand U26338 (N_26338,N_25024,N_24052);
xor U26339 (N_26339,N_25130,N_24928);
xor U26340 (N_26340,N_25455,N_24620);
nand U26341 (N_26341,N_25259,N_24258);
nand U26342 (N_26342,N_24568,N_25177);
or U26343 (N_26343,N_25121,N_24087);
nor U26344 (N_26344,N_24372,N_24425);
nand U26345 (N_26345,N_25164,N_24504);
nand U26346 (N_26346,N_24955,N_25211);
and U26347 (N_26347,N_24962,N_24167);
or U26348 (N_26348,N_24818,N_24587);
nand U26349 (N_26349,N_24857,N_25015);
nand U26350 (N_26350,N_24115,N_24762);
nand U26351 (N_26351,N_24011,N_24014);
nand U26352 (N_26352,N_24335,N_24324);
nor U26353 (N_26353,N_24619,N_24110);
and U26354 (N_26354,N_25144,N_24218);
and U26355 (N_26355,N_24954,N_24952);
xor U26356 (N_26356,N_24307,N_24674);
nand U26357 (N_26357,N_24684,N_25140);
nor U26358 (N_26358,N_24088,N_24723);
nor U26359 (N_26359,N_24282,N_25415);
or U26360 (N_26360,N_24959,N_24067);
nand U26361 (N_26361,N_24745,N_24514);
and U26362 (N_26362,N_25353,N_24592);
xnor U26363 (N_26363,N_24062,N_25143);
or U26364 (N_26364,N_25265,N_24875);
and U26365 (N_26365,N_24234,N_25177);
xor U26366 (N_26366,N_24404,N_25331);
or U26367 (N_26367,N_25385,N_25472);
or U26368 (N_26368,N_25218,N_24149);
nor U26369 (N_26369,N_25107,N_24887);
and U26370 (N_26370,N_24051,N_24896);
nor U26371 (N_26371,N_24159,N_24824);
xor U26372 (N_26372,N_24750,N_24445);
nor U26373 (N_26373,N_24974,N_24633);
nor U26374 (N_26374,N_24355,N_25310);
nand U26375 (N_26375,N_24537,N_24514);
nand U26376 (N_26376,N_24812,N_25491);
xor U26377 (N_26377,N_24506,N_24005);
nor U26378 (N_26378,N_25155,N_24868);
and U26379 (N_26379,N_24403,N_25034);
or U26380 (N_26380,N_24427,N_24944);
or U26381 (N_26381,N_24948,N_24258);
or U26382 (N_26382,N_24575,N_25410);
and U26383 (N_26383,N_25471,N_24673);
nand U26384 (N_26384,N_25112,N_24233);
and U26385 (N_26385,N_25119,N_25148);
or U26386 (N_26386,N_24514,N_25466);
nand U26387 (N_26387,N_25148,N_24119);
and U26388 (N_26388,N_25234,N_25435);
nand U26389 (N_26389,N_24126,N_24295);
and U26390 (N_26390,N_24388,N_25476);
and U26391 (N_26391,N_25137,N_25423);
and U26392 (N_26392,N_24216,N_24071);
xnor U26393 (N_26393,N_24051,N_25027);
or U26394 (N_26394,N_24447,N_24343);
and U26395 (N_26395,N_24235,N_24324);
and U26396 (N_26396,N_24529,N_24633);
and U26397 (N_26397,N_25024,N_24749);
nand U26398 (N_26398,N_24298,N_24754);
nor U26399 (N_26399,N_25497,N_24302);
xnor U26400 (N_26400,N_25369,N_24092);
and U26401 (N_26401,N_24844,N_24216);
nor U26402 (N_26402,N_24013,N_25421);
nor U26403 (N_26403,N_24260,N_24307);
xnor U26404 (N_26404,N_24715,N_24750);
xnor U26405 (N_26405,N_24091,N_25344);
nor U26406 (N_26406,N_25072,N_24335);
nor U26407 (N_26407,N_24412,N_24416);
nor U26408 (N_26408,N_24724,N_25442);
and U26409 (N_26409,N_24593,N_24085);
xor U26410 (N_26410,N_25276,N_24514);
nand U26411 (N_26411,N_24574,N_24931);
xor U26412 (N_26412,N_24929,N_24811);
and U26413 (N_26413,N_25463,N_24775);
nor U26414 (N_26414,N_24565,N_24415);
nand U26415 (N_26415,N_24930,N_24843);
or U26416 (N_26416,N_24221,N_24533);
or U26417 (N_26417,N_24846,N_25319);
xnor U26418 (N_26418,N_25484,N_25216);
and U26419 (N_26419,N_25392,N_24236);
or U26420 (N_26420,N_24962,N_25470);
and U26421 (N_26421,N_24263,N_25394);
xor U26422 (N_26422,N_25183,N_24910);
nor U26423 (N_26423,N_24637,N_24341);
and U26424 (N_26424,N_25358,N_25162);
nand U26425 (N_26425,N_24708,N_24838);
or U26426 (N_26426,N_24841,N_24338);
nand U26427 (N_26427,N_24421,N_24678);
xnor U26428 (N_26428,N_25115,N_24657);
nand U26429 (N_26429,N_24938,N_24204);
nor U26430 (N_26430,N_25097,N_24239);
nor U26431 (N_26431,N_24987,N_24701);
nor U26432 (N_26432,N_25052,N_24196);
and U26433 (N_26433,N_24225,N_24610);
or U26434 (N_26434,N_25028,N_25076);
nor U26435 (N_26435,N_24797,N_25384);
or U26436 (N_26436,N_24910,N_25001);
or U26437 (N_26437,N_24706,N_24620);
xor U26438 (N_26438,N_24065,N_24225);
and U26439 (N_26439,N_25149,N_25190);
and U26440 (N_26440,N_24001,N_24549);
nor U26441 (N_26441,N_25101,N_24991);
nand U26442 (N_26442,N_25154,N_24828);
and U26443 (N_26443,N_25305,N_24246);
or U26444 (N_26444,N_24352,N_24024);
and U26445 (N_26445,N_24125,N_25137);
nor U26446 (N_26446,N_24103,N_25014);
and U26447 (N_26447,N_25243,N_24555);
nand U26448 (N_26448,N_25352,N_24032);
xnor U26449 (N_26449,N_24497,N_24569);
xor U26450 (N_26450,N_24849,N_24129);
xnor U26451 (N_26451,N_24808,N_24014);
nor U26452 (N_26452,N_25237,N_24269);
and U26453 (N_26453,N_25211,N_24008);
xnor U26454 (N_26454,N_24117,N_24673);
and U26455 (N_26455,N_24106,N_24860);
or U26456 (N_26456,N_24366,N_25017);
xor U26457 (N_26457,N_24048,N_24396);
and U26458 (N_26458,N_25406,N_24069);
nor U26459 (N_26459,N_25007,N_24494);
nand U26460 (N_26460,N_24922,N_24301);
nand U26461 (N_26461,N_25277,N_24813);
and U26462 (N_26462,N_25280,N_24289);
or U26463 (N_26463,N_24185,N_24606);
nor U26464 (N_26464,N_24520,N_24215);
nor U26465 (N_26465,N_24558,N_24536);
and U26466 (N_26466,N_24693,N_24290);
nor U26467 (N_26467,N_25310,N_24877);
nand U26468 (N_26468,N_24708,N_24698);
nor U26469 (N_26469,N_25363,N_24206);
xor U26470 (N_26470,N_24101,N_24147);
or U26471 (N_26471,N_25471,N_25018);
and U26472 (N_26472,N_25044,N_25217);
nor U26473 (N_26473,N_24964,N_24618);
xnor U26474 (N_26474,N_24990,N_24725);
and U26475 (N_26475,N_25222,N_24818);
xor U26476 (N_26476,N_24786,N_25180);
and U26477 (N_26477,N_25284,N_25398);
xnor U26478 (N_26478,N_24721,N_24963);
xor U26479 (N_26479,N_24358,N_25295);
nor U26480 (N_26480,N_24210,N_25488);
or U26481 (N_26481,N_24218,N_24814);
or U26482 (N_26482,N_24335,N_24637);
xnor U26483 (N_26483,N_24875,N_25400);
or U26484 (N_26484,N_24891,N_24526);
or U26485 (N_26485,N_25475,N_24881);
nor U26486 (N_26486,N_24383,N_24490);
nand U26487 (N_26487,N_25172,N_24599);
and U26488 (N_26488,N_25117,N_25049);
or U26489 (N_26489,N_25166,N_24888);
xnor U26490 (N_26490,N_24441,N_24527);
nor U26491 (N_26491,N_25050,N_24394);
xnor U26492 (N_26492,N_25388,N_24000);
xnor U26493 (N_26493,N_24603,N_24202);
nand U26494 (N_26494,N_24336,N_24406);
or U26495 (N_26495,N_24518,N_25341);
xnor U26496 (N_26496,N_24696,N_24558);
nand U26497 (N_26497,N_24476,N_25326);
nand U26498 (N_26498,N_24654,N_24984);
nor U26499 (N_26499,N_24939,N_25339);
nor U26500 (N_26500,N_24193,N_24293);
nand U26501 (N_26501,N_24524,N_24295);
or U26502 (N_26502,N_24168,N_24490);
nor U26503 (N_26503,N_24371,N_24323);
nand U26504 (N_26504,N_25326,N_24198);
or U26505 (N_26505,N_25213,N_24441);
or U26506 (N_26506,N_24281,N_24291);
and U26507 (N_26507,N_25331,N_24856);
xnor U26508 (N_26508,N_24203,N_24301);
and U26509 (N_26509,N_25291,N_24777);
and U26510 (N_26510,N_25184,N_24487);
nand U26511 (N_26511,N_24108,N_25212);
xor U26512 (N_26512,N_24838,N_24955);
xnor U26513 (N_26513,N_25414,N_24000);
nor U26514 (N_26514,N_24082,N_24591);
nor U26515 (N_26515,N_24846,N_24633);
and U26516 (N_26516,N_25249,N_24149);
and U26517 (N_26517,N_24133,N_25320);
xnor U26518 (N_26518,N_24187,N_24097);
and U26519 (N_26519,N_24383,N_24674);
nand U26520 (N_26520,N_24860,N_25159);
nand U26521 (N_26521,N_24093,N_25086);
and U26522 (N_26522,N_24727,N_24457);
xnor U26523 (N_26523,N_25213,N_24473);
xnor U26524 (N_26524,N_24405,N_24961);
or U26525 (N_26525,N_24368,N_24765);
or U26526 (N_26526,N_24304,N_24459);
nand U26527 (N_26527,N_25073,N_24661);
nand U26528 (N_26528,N_24660,N_25112);
nand U26529 (N_26529,N_24962,N_25148);
or U26530 (N_26530,N_25050,N_25056);
xor U26531 (N_26531,N_24257,N_24351);
or U26532 (N_26532,N_24003,N_25489);
or U26533 (N_26533,N_25116,N_24935);
and U26534 (N_26534,N_25309,N_25247);
or U26535 (N_26535,N_25284,N_25252);
nor U26536 (N_26536,N_24404,N_24595);
and U26537 (N_26537,N_25354,N_24252);
xnor U26538 (N_26538,N_24073,N_24407);
nand U26539 (N_26539,N_25356,N_25343);
nor U26540 (N_26540,N_24315,N_24088);
and U26541 (N_26541,N_24990,N_24364);
nor U26542 (N_26542,N_24006,N_24932);
nor U26543 (N_26543,N_24633,N_25211);
or U26544 (N_26544,N_24971,N_24446);
nor U26545 (N_26545,N_24314,N_24766);
nand U26546 (N_26546,N_24983,N_25445);
or U26547 (N_26547,N_24770,N_24326);
nor U26548 (N_26548,N_24640,N_25265);
nand U26549 (N_26549,N_24159,N_24927);
and U26550 (N_26550,N_25112,N_24915);
xnor U26551 (N_26551,N_25398,N_24838);
and U26552 (N_26552,N_25111,N_24170);
xnor U26553 (N_26553,N_25185,N_24577);
or U26554 (N_26554,N_24163,N_25312);
and U26555 (N_26555,N_24772,N_24239);
nand U26556 (N_26556,N_24890,N_24143);
and U26557 (N_26557,N_25109,N_25368);
nor U26558 (N_26558,N_24559,N_24560);
xnor U26559 (N_26559,N_25412,N_25338);
and U26560 (N_26560,N_24062,N_24394);
nor U26561 (N_26561,N_25116,N_25290);
nand U26562 (N_26562,N_24575,N_24934);
xor U26563 (N_26563,N_24560,N_24125);
or U26564 (N_26564,N_24173,N_25412);
xnor U26565 (N_26565,N_24146,N_25198);
or U26566 (N_26566,N_24510,N_24112);
xnor U26567 (N_26567,N_24541,N_25414);
or U26568 (N_26568,N_24819,N_25129);
nand U26569 (N_26569,N_24981,N_25388);
nor U26570 (N_26570,N_24383,N_24488);
nor U26571 (N_26571,N_25263,N_24232);
or U26572 (N_26572,N_24154,N_24977);
xnor U26573 (N_26573,N_24094,N_24732);
nand U26574 (N_26574,N_24916,N_25309);
nand U26575 (N_26575,N_24339,N_24866);
nor U26576 (N_26576,N_24627,N_24900);
or U26577 (N_26577,N_25234,N_25269);
nor U26578 (N_26578,N_24765,N_24205);
xor U26579 (N_26579,N_25431,N_24956);
nor U26580 (N_26580,N_24513,N_24842);
nand U26581 (N_26581,N_25319,N_24541);
or U26582 (N_26582,N_25173,N_25352);
xnor U26583 (N_26583,N_24700,N_24727);
and U26584 (N_26584,N_25484,N_24595);
nor U26585 (N_26585,N_25196,N_24479);
xor U26586 (N_26586,N_24272,N_25037);
or U26587 (N_26587,N_25464,N_25425);
xnor U26588 (N_26588,N_25015,N_24498);
or U26589 (N_26589,N_24998,N_25274);
or U26590 (N_26590,N_24451,N_24100);
or U26591 (N_26591,N_24953,N_24397);
xnor U26592 (N_26592,N_24706,N_24906);
or U26593 (N_26593,N_25187,N_25152);
nor U26594 (N_26594,N_24850,N_25173);
nand U26595 (N_26595,N_24988,N_25345);
and U26596 (N_26596,N_24581,N_24192);
and U26597 (N_26597,N_24085,N_24010);
or U26598 (N_26598,N_24357,N_24570);
nand U26599 (N_26599,N_25382,N_24715);
nor U26600 (N_26600,N_24464,N_24931);
nor U26601 (N_26601,N_24399,N_25233);
or U26602 (N_26602,N_25323,N_25269);
nand U26603 (N_26603,N_24520,N_24399);
or U26604 (N_26604,N_24139,N_25155);
nand U26605 (N_26605,N_25069,N_25050);
nand U26606 (N_26606,N_24489,N_25393);
xor U26607 (N_26607,N_24626,N_24550);
xnor U26608 (N_26608,N_24872,N_24823);
nand U26609 (N_26609,N_25411,N_25266);
nand U26610 (N_26610,N_25014,N_24252);
and U26611 (N_26611,N_24619,N_25324);
xnor U26612 (N_26612,N_24004,N_24985);
or U26613 (N_26613,N_25276,N_25307);
xor U26614 (N_26614,N_24011,N_24206);
or U26615 (N_26615,N_25287,N_24556);
or U26616 (N_26616,N_24892,N_25417);
nand U26617 (N_26617,N_24364,N_24305);
nand U26618 (N_26618,N_24856,N_24737);
or U26619 (N_26619,N_24589,N_25156);
or U26620 (N_26620,N_24886,N_24477);
nor U26621 (N_26621,N_25364,N_24418);
nor U26622 (N_26622,N_25406,N_25014);
and U26623 (N_26623,N_25413,N_24002);
nor U26624 (N_26624,N_24616,N_25311);
nor U26625 (N_26625,N_25223,N_24140);
nand U26626 (N_26626,N_24991,N_25064);
nor U26627 (N_26627,N_25017,N_25327);
nor U26628 (N_26628,N_24474,N_25291);
nor U26629 (N_26629,N_25477,N_25476);
or U26630 (N_26630,N_24184,N_25190);
nor U26631 (N_26631,N_25240,N_25448);
nor U26632 (N_26632,N_24711,N_25222);
nor U26633 (N_26633,N_25434,N_24116);
xor U26634 (N_26634,N_24323,N_25232);
or U26635 (N_26635,N_25136,N_24468);
xnor U26636 (N_26636,N_24868,N_24337);
and U26637 (N_26637,N_24152,N_25248);
or U26638 (N_26638,N_24173,N_24710);
and U26639 (N_26639,N_24505,N_24250);
and U26640 (N_26640,N_25169,N_25039);
nor U26641 (N_26641,N_24660,N_24352);
nor U26642 (N_26642,N_25059,N_25066);
or U26643 (N_26643,N_24649,N_24378);
or U26644 (N_26644,N_24668,N_25356);
or U26645 (N_26645,N_24247,N_24415);
nor U26646 (N_26646,N_24075,N_24928);
nand U26647 (N_26647,N_25017,N_24943);
or U26648 (N_26648,N_24412,N_24078);
nand U26649 (N_26649,N_24260,N_24230);
nand U26650 (N_26650,N_24198,N_24115);
nor U26651 (N_26651,N_25401,N_24156);
nor U26652 (N_26652,N_24525,N_25094);
nand U26653 (N_26653,N_24139,N_25066);
nor U26654 (N_26654,N_24037,N_24913);
xnor U26655 (N_26655,N_24380,N_24178);
or U26656 (N_26656,N_24795,N_24328);
and U26657 (N_26657,N_24828,N_25270);
nor U26658 (N_26658,N_24281,N_24487);
and U26659 (N_26659,N_24430,N_24194);
and U26660 (N_26660,N_24165,N_24544);
and U26661 (N_26661,N_24646,N_25289);
and U26662 (N_26662,N_24910,N_25028);
nand U26663 (N_26663,N_24913,N_25390);
nand U26664 (N_26664,N_24891,N_24190);
or U26665 (N_26665,N_25348,N_25341);
and U26666 (N_26666,N_25388,N_24457);
nor U26667 (N_26667,N_24211,N_25058);
and U26668 (N_26668,N_24580,N_24640);
xnor U26669 (N_26669,N_25424,N_24667);
or U26670 (N_26670,N_24079,N_25237);
nor U26671 (N_26671,N_24582,N_24373);
nor U26672 (N_26672,N_24998,N_25445);
xor U26673 (N_26673,N_24179,N_24710);
nor U26674 (N_26674,N_24260,N_25006);
or U26675 (N_26675,N_24565,N_24030);
xnor U26676 (N_26676,N_25433,N_24400);
xor U26677 (N_26677,N_24517,N_24991);
or U26678 (N_26678,N_25225,N_25391);
nand U26679 (N_26679,N_24932,N_24769);
nor U26680 (N_26680,N_25248,N_24969);
or U26681 (N_26681,N_25410,N_24899);
or U26682 (N_26682,N_24349,N_24026);
or U26683 (N_26683,N_24217,N_24387);
xor U26684 (N_26684,N_24415,N_25166);
and U26685 (N_26685,N_24932,N_25294);
nor U26686 (N_26686,N_24347,N_24822);
nor U26687 (N_26687,N_24031,N_24174);
nand U26688 (N_26688,N_24032,N_24343);
xnor U26689 (N_26689,N_24012,N_24496);
and U26690 (N_26690,N_24393,N_25323);
nand U26691 (N_26691,N_24548,N_25437);
or U26692 (N_26692,N_24942,N_24318);
nand U26693 (N_26693,N_25319,N_25209);
or U26694 (N_26694,N_25234,N_24017);
or U26695 (N_26695,N_24183,N_24981);
nor U26696 (N_26696,N_24786,N_24317);
nand U26697 (N_26697,N_24545,N_25306);
nand U26698 (N_26698,N_25459,N_24069);
nand U26699 (N_26699,N_25383,N_25287);
and U26700 (N_26700,N_24838,N_25023);
xnor U26701 (N_26701,N_24450,N_24982);
nand U26702 (N_26702,N_24861,N_24126);
nor U26703 (N_26703,N_24304,N_24047);
nor U26704 (N_26704,N_24410,N_25389);
nor U26705 (N_26705,N_24856,N_24459);
nand U26706 (N_26706,N_24551,N_25126);
xnor U26707 (N_26707,N_24743,N_24452);
or U26708 (N_26708,N_24703,N_24862);
or U26709 (N_26709,N_24054,N_24288);
xnor U26710 (N_26710,N_24651,N_24001);
nor U26711 (N_26711,N_25120,N_24492);
xor U26712 (N_26712,N_24421,N_25308);
xnor U26713 (N_26713,N_24702,N_25331);
and U26714 (N_26714,N_25313,N_24916);
xnor U26715 (N_26715,N_24435,N_24840);
nor U26716 (N_26716,N_24013,N_25327);
and U26717 (N_26717,N_25269,N_24250);
and U26718 (N_26718,N_25269,N_24449);
or U26719 (N_26719,N_24197,N_24783);
or U26720 (N_26720,N_25224,N_24950);
or U26721 (N_26721,N_24762,N_24442);
nor U26722 (N_26722,N_25321,N_24004);
xnor U26723 (N_26723,N_25413,N_24893);
nor U26724 (N_26724,N_24785,N_25197);
nand U26725 (N_26725,N_24461,N_25240);
nand U26726 (N_26726,N_25413,N_24782);
nand U26727 (N_26727,N_24903,N_24150);
and U26728 (N_26728,N_24560,N_24772);
nor U26729 (N_26729,N_24521,N_24656);
and U26730 (N_26730,N_24371,N_24619);
or U26731 (N_26731,N_25194,N_24143);
and U26732 (N_26732,N_24440,N_24016);
xor U26733 (N_26733,N_24020,N_25127);
nand U26734 (N_26734,N_25128,N_24734);
xnor U26735 (N_26735,N_24951,N_24571);
nor U26736 (N_26736,N_25450,N_24015);
and U26737 (N_26737,N_25032,N_24293);
xor U26738 (N_26738,N_24372,N_25021);
and U26739 (N_26739,N_24519,N_25342);
and U26740 (N_26740,N_24958,N_25079);
xor U26741 (N_26741,N_24896,N_24165);
and U26742 (N_26742,N_24904,N_24812);
nor U26743 (N_26743,N_24620,N_24830);
nand U26744 (N_26744,N_24159,N_25339);
nand U26745 (N_26745,N_24026,N_24221);
and U26746 (N_26746,N_25249,N_24298);
and U26747 (N_26747,N_24428,N_24075);
and U26748 (N_26748,N_24208,N_24882);
xor U26749 (N_26749,N_24672,N_24036);
or U26750 (N_26750,N_24592,N_25224);
or U26751 (N_26751,N_25221,N_24627);
or U26752 (N_26752,N_24359,N_25281);
nor U26753 (N_26753,N_24598,N_25100);
nor U26754 (N_26754,N_24126,N_24008);
nor U26755 (N_26755,N_25106,N_24405);
nor U26756 (N_26756,N_24980,N_24358);
or U26757 (N_26757,N_24776,N_25074);
xnor U26758 (N_26758,N_24678,N_24163);
and U26759 (N_26759,N_24153,N_25283);
nand U26760 (N_26760,N_24689,N_24135);
xor U26761 (N_26761,N_24464,N_25495);
nor U26762 (N_26762,N_24693,N_24550);
xor U26763 (N_26763,N_24984,N_24348);
or U26764 (N_26764,N_24982,N_24656);
or U26765 (N_26765,N_24356,N_25099);
or U26766 (N_26766,N_24075,N_24251);
nand U26767 (N_26767,N_24736,N_24804);
nor U26768 (N_26768,N_24831,N_25162);
or U26769 (N_26769,N_25242,N_24004);
and U26770 (N_26770,N_24768,N_24393);
or U26771 (N_26771,N_24136,N_24403);
nor U26772 (N_26772,N_25264,N_24023);
or U26773 (N_26773,N_24745,N_24876);
nand U26774 (N_26774,N_25405,N_25204);
and U26775 (N_26775,N_24266,N_24708);
nor U26776 (N_26776,N_25133,N_24081);
xnor U26777 (N_26777,N_24421,N_24582);
and U26778 (N_26778,N_24492,N_24017);
and U26779 (N_26779,N_24683,N_24772);
and U26780 (N_26780,N_24405,N_24026);
and U26781 (N_26781,N_25058,N_24321);
or U26782 (N_26782,N_24878,N_24631);
nor U26783 (N_26783,N_24666,N_25403);
nor U26784 (N_26784,N_24484,N_24239);
nor U26785 (N_26785,N_25054,N_25199);
or U26786 (N_26786,N_24644,N_24769);
or U26787 (N_26787,N_24569,N_25477);
xor U26788 (N_26788,N_25276,N_25209);
nand U26789 (N_26789,N_24411,N_24523);
nor U26790 (N_26790,N_24371,N_25187);
nor U26791 (N_26791,N_25312,N_24042);
or U26792 (N_26792,N_25392,N_24483);
xnor U26793 (N_26793,N_24720,N_24138);
and U26794 (N_26794,N_24592,N_24595);
nor U26795 (N_26795,N_25419,N_25045);
nor U26796 (N_26796,N_25000,N_24112);
xnor U26797 (N_26797,N_24847,N_24490);
nor U26798 (N_26798,N_24448,N_24937);
xnor U26799 (N_26799,N_24516,N_25021);
or U26800 (N_26800,N_25062,N_24456);
nand U26801 (N_26801,N_25294,N_24740);
nor U26802 (N_26802,N_24421,N_25466);
nand U26803 (N_26803,N_24017,N_25139);
xor U26804 (N_26804,N_24524,N_24752);
or U26805 (N_26805,N_24839,N_24217);
xnor U26806 (N_26806,N_24719,N_25066);
nand U26807 (N_26807,N_25241,N_25044);
nor U26808 (N_26808,N_25215,N_24843);
nand U26809 (N_26809,N_25459,N_24004);
xnor U26810 (N_26810,N_24404,N_24815);
nor U26811 (N_26811,N_25040,N_25273);
nor U26812 (N_26812,N_24220,N_24323);
xnor U26813 (N_26813,N_24276,N_24048);
or U26814 (N_26814,N_24456,N_24178);
nor U26815 (N_26815,N_24362,N_24180);
and U26816 (N_26816,N_24579,N_25471);
or U26817 (N_26817,N_24103,N_24911);
xor U26818 (N_26818,N_24205,N_24130);
or U26819 (N_26819,N_24953,N_25499);
xor U26820 (N_26820,N_25141,N_25243);
nand U26821 (N_26821,N_25056,N_25018);
or U26822 (N_26822,N_25406,N_24770);
and U26823 (N_26823,N_25382,N_24799);
nand U26824 (N_26824,N_24423,N_24783);
or U26825 (N_26825,N_24393,N_24977);
nand U26826 (N_26826,N_25233,N_25314);
nand U26827 (N_26827,N_25107,N_25299);
nand U26828 (N_26828,N_25242,N_24184);
xor U26829 (N_26829,N_24718,N_25199);
or U26830 (N_26830,N_24925,N_24554);
or U26831 (N_26831,N_25385,N_24658);
nor U26832 (N_26832,N_24524,N_24564);
xnor U26833 (N_26833,N_25160,N_24419);
nand U26834 (N_26834,N_24045,N_24973);
nor U26835 (N_26835,N_24263,N_24886);
xor U26836 (N_26836,N_24912,N_24990);
nand U26837 (N_26837,N_24484,N_24441);
nand U26838 (N_26838,N_24734,N_25491);
nand U26839 (N_26839,N_24811,N_25274);
xnor U26840 (N_26840,N_24674,N_24904);
nor U26841 (N_26841,N_24377,N_25204);
nand U26842 (N_26842,N_24341,N_24250);
nand U26843 (N_26843,N_24396,N_24869);
and U26844 (N_26844,N_24088,N_25025);
xor U26845 (N_26845,N_25235,N_25320);
and U26846 (N_26846,N_24214,N_24185);
or U26847 (N_26847,N_24098,N_24166);
and U26848 (N_26848,N_24567,N_24389);
nor U26849 (N_26849,N_25138,N_24539);
and U26850 (N_26850,N_25196,N_24963);
or U26851 (N_26851,N_25387,N_24517);
xnor U26852 (N_26852,N_24280,N_24622);
or U26853 (N_26853,N_25057,N_25200);
and U26854 (N_26854,N_24351,N_24425);
or U26855 (N_26855,N_25093,N_25279);
and U26856 (N_26856,N_24775,N_24396);
nand U26857 (N_26857,N_25458,N_24584);
or U26858 (N_26858,N_24737,N_24921);
and U26859 (N_26859,N_24846,N_24921);
and U26860 (N_26860,N_24587,N_24515);
and U26861 (N_26861,N_24606,N_24145);
xnor U26862 (N_26862,N_24084,N_25028);
xnor U26863 (N_26863,N_24608,N_24911);
or U26864 (N_26864,N_24740,N_25133);
nand U26865 (N_26865,N_24345,N_25388);
and U26866 (N_26866,N_24794,N_25413);
and U26867 (N_26867,N_24184,N_24686);
or U26868 (N_26868,N_24440,N_24921);
or U26869 (N_26869,N_24096,N_25083);
nor U26870 (N_26870,N_24294,N_24526);
and U26871 (N_26871,N_24817,N_25365);
nand U26872 (N_26872,N_25011,N_24210);
nand U26873 (N_26873,N_24942,N_24365);
and U26874 (N_26874,N_24395,N_24315);
xnor U26875 (N_26875,N_25183,N_24294);
xor U26876 (N_26876,N_24031,N_24458);
nor U26877 (N_26877,N_25464,N_24920);
and U26878 (N_26878,N_24142,N_24500);
nor U26879 (N_26879,N_24049,N_24759);
nand U26880 (N_26880,N_24446,N_24209);
and U26881 (N_26881,N_25492,N_24626);
or U26882 (N_26882,N_25068,N_25161);
nor U26883 (N_26883,N_24662,N_24724);
nor U26884 (N_26884,N_25215,N_24391);
and U26885 (N_26885,N_24470,N_25359);
or U26886 (N_26886,N_24026,N_24703);
nor U26887 (N_26887,N_25411,N_24913);
nand U26888 (N_26888,N_25077,N_24324);
nand U26889 (N_26889,N_25485,N_24040);
xor U26890 (N_26890,N_25183,N_24145);
xnor U26891 (N_26891,N_24567,N_25379);
nand U26892 (N_26892,N_24804,N_25321);
or U26893 (N_26893,N_25328,N_24205);
xor U26894 (N_26894,N_24998,N_25201);
nor U26895 (N_26895,N_25372,N_24943);
xnor U26896 (N_26896,N_24268,N_24495);
nor U26897 (N_26897,N_25441,N_24345);
or U26898 (N_26898,N_25434,N_24581);
and U26899 (N_26899,N_24325,N_25044);
or U26900 (N_26900,N_25439,N_24463);
or U26901 (N_26901,N_24145,N_25195);
and U26902 (N_26902,N_25004,N_25200);
and U26903 (N_26903,N_25253,N_24766);
xor U26904 (N_26904,N_24478,N_25412);
and U26905 (N_26905,N_24140,N_25206);
xnor U26906 (N_26906,N_24830,N_24591);
nand U26907 (N_26907,N_24633,N_24020);
nand U26908 (N_26908,N_24719,N_24095);
nand U26909 (N_26909,N_25418,N_24920);
or U26910 (N_26910,N_24125,N_24245);
nand U26911 (N_26911,N_24476,N_24912);
nor U26912 (N_26912,N_25128,N_24105);
and U26913 (N_26913,N_25186,N_25135);
xnor U26914 (N_26914,N_24177,N_25177);
or U26915 (N_26915,N_24779,N_25188);
nor U26916 (N_26916,N_24081,N_25135);
and U26917 (N_26917,N_25351,N_25496);
nand U26918 (N_26918,N_25308,N_25447);
and U26919 (N_26919,N_25251,N_25160);
and U26920 (N_26920,N_24365,N_24336);
nor U26921 (N_26921,N_25191,N_24860);
xnor U26922 (N_26922,N_24920,N_25310);
nor U26923 (N_26923,N_24256,N_25177);
xor U26924 (N_26924,N_24956,N_25246);
nand U26925 (N_26925,N_24502,N_24683);
or U26926 (N_26926,N_25459,N_25009);
xnor U26927 (N_26927,N_24758,N_24500);
nand U26928 (N_26928,N_24445,N_25222);
nor U26929 (N_26929,N_25163,N_24711);
and U26930 (N_26930,N_24515,N_24119);
nand U26931 (N_26931,N_24067,N_24075);
nand U26932 (N_26932,N_24525,N_25084);
nand U26933 (N_26933,N_24506,N_24569);
xor U26934 (N_26934,N_24607,N_25436);
nand U26935 (N_26935,N_24314,N_24405);
nand U26936 (N_26936,N_25041,N_24776);
and U26937 (N_26937,N_24666,N_25410);
nand U26938 (N_26938,N_24592,N_24724);
xnor U26939 (N_26939,N_24993,N_24517);
and U26940 (N_26940,N_25145,N_24991);
or U26941 (N_26941,N_25168,N_25329);
nor U26942 (N_26942,N_25467,N_24397);
nor U26943 (N_26943,N_24714,N_25293);
or U26944 (N_26944,N_25218,N_24538);
nor U26945 (N_26945,N_25085,N_24542);
xor U26946 (N_26946,N_25179,N_25467);
and U26947 (N_26947,N_24716,N_24514);
xnor U26948 (N_26948,N_25331,N_25277);
and U26949 (N_26949,N_24599,N_24468);
nor U26950 (N_26950,N_24299,N_25302);
nand U26951 (N_26951,N_24473,N_24275);
xnor U26952 (N_26952,N_24401,N_25107);
xnor U26953 (N_26953,N_24973,N_25080);
nand U26954 (N_26954,N_25311,N_24816);
nor U26955 (N_26955,N_24791,N_25191);
or U26956 (N_26956,N_24248,N_24114);
nor U26957 (N_26957,N_25273,N_24986);
and U26958 (N_26958,N_25139,N_24245);
xor U26959 (N_26959,N_24129,N_24743);
nand U26960 (N_26960,N_24906,N_24897);
xnor U26961 (N_26961,N_25279,N_24655);
nand U26962 (N_26962,N_25069,N_25467);
or U26963 (N_26963,N_24930,N_25111);
or U26964 (N_26964,N_24289,N_24448);
or U26965 (N_26965,N_24934,N_24056);
and U26966 (N_26966,N_24786,N_24923);
xnor U26967 (N_26967,N_24879,N_25040);
xnor U26968 (N_26968,N_24132,N_25219);
or U26969 (N_26969,N_24134,N_24260);
nor U26970 (N_26970,N_24662,N_24961);
nor U26971 (N_26971,N_25133,N_24943);
or U26972 (N_26972,N_24690,N_25156);
nor U26973 (N_26973,N_24108,N_24087);
xor U26974 (N_26974,N_25054,N_24257);
xor U26975 (N_26975,N_25034,N_24837);
xnor U26976 (N_26976,N_24397,N_24180);
and U26977 (N_26977,N_24280,N_24647);
and U26978 (N_26978,N_24033,N_24790);
nor U26979 (N_26979,N_24331,N_24392);
or U26980 (N_26980,N_24656,N_25416);
or U26981 (N_26981,N_25397,N_24803);
and U26982 (N_26982,N_24856,N_24808);
and U26983 (N_26983,N_24508,N_25105);
and U26984 (N_26984,N_25311,N_24157);
and U26985 (N_26985,N_24198,N_24228);
nor U26986 (N_26986,N_24058,N_25414);
nand U26987 (N_26987,N_24594,N_24605);
xnor U26988 (N_26988,N_25092,N_24379);
nor U26989 (N_26989,N_24360,N_25279);
nand U26990 (N_26990,N_25244,N_24001);
or U26991 (N_26991,N_24261,N_24250);
xnor U26992 (N_26992,N_25116,N_24498);
nand U26993 (N_26993,N_24292,N_24801);
xnor U26994 (N_26994,N_24742,N_25193);
and U26995 (N_26995,N_24628,N_24808);
nand U26996 (N_26996,N_24671,N_25202);
nor U26997 (N_26997,N_24616,N_24808);
nor U26998 (N_26998,N_24534,N_24147);
xor U26999 (N_26999,N_25135,N_24971);
or U27000 (N_27000,N_26804,N_26546);
xor U27001 (N_27001,N_26442,N_25625);
or U27002 (N_27002,N_25646,N_26862);
and U27003 (N_27003,N_25811,N_26336);
xor U27004 (N_27004,N_26056,N_25568);
nand U27005 (N_27005,N_26491,N_26250);
and U27006 (N_27006,N_26682,N_25964);
xnor U27007 (N_27007,N_26517,N_26693);
and U27008 (N_27008,N_26438,N_26649);
nand U27009 (N_27009,N_26227,N_25543);
nand U27010 (N_27010,N_25752,N_26125);
or U27011 (N_27011,N_26267,N_25627);
nor U27012 (N_27012,N_26746,N_25609);
nor U27013 (N_27013,N_25536,N_26918);
nand U27014 (N_27014,N_25859,N_26032);
nor U27015 (N_27015,N_26779,N_26843);
xor U27016 (N_27016,N_26280,N_26194);
nor U27017 (N_27017,N_25762,N_25582);
or U27018 (N_27018,N_25677,N_26664);
xnor U27019 (N_27019,N_25841,N_25826);
nand U27020 (N_27020,N_25507,N_25660);
and U27021 (N_27021,N_26900,N_26157);
and U27022 (N_27022,N_26705,N_25516);
xor U27023 (N_27023,N_26386,N_26987);
nand U27024 (N_27024,N_25969,N_26313);
xnor U27025 (N_27025,N_26497,N_25647);
and U27026 (N_27026,N_25958,N_26257);
and U27027 (N_27027,N_25804,N_26030);
xnor U27028 (N_27028,N_26506,N_25699);
and U27029 (N_27029,N_26234,N_25670);
xor U27030 (N_27030,N_26767,N_26970);
xnor U27031 (N_27031,N_26667,N_26453);
nand U27032 (N_27032,N_26369,N_25860);
or U27033 (N_27033,N_26635,N_26008);
nand U27034 (N_27034,N_26230,N_26081);
nor U27035 (N_27035,N_26816,N_26122);
nand U27036 (N_27036,N_25888,N_26305);
xnor U27037 (N_27037,N_25922,N_26296);
or U27038 (N_27038,N_25503,N_26521);
xnor U27039 (N_27039,N_25707,N_26299);
or U27040 (N_27040,N_26284,N_26513);
or U27041 (N_27041,N_26983,N_26685);
nand U27042 (N_27042,N_25758,N_26569);
and U27043 (N_27043,N_26055,N_25626);
xnor U27044 (N_27044,N_25622,N_26264);
nand U27045 (N_27045,N_25680,N_25664);
nand U27046 (N_27046,N_26289,N_26557);
and U27047 (N_27047,N_26858,N_26728);
nor U27048 (N_27048,N_26845,N_25753);
nand U27049 (N_27049,N_25673,N_26531);
xor U27050 (N_27050,N_25994,N_26961);
xnor U27051 (N_27051,N_26205,N_26803);
and U27052 (N_27052,N_26487,N_26895);
or U27053 (N_27053,N_26066,N_26080);
nor U27054 (N_27054,N_26043,N_26880);
xor U27055 (N_27055,N_26692,N_26412);
or U27056 (N_27056,N_26168,N_26777);
or U27057 (N_27057,N_26181,N_26394);
or U27058 (N_27058,N_26347,N_26159);
nor U27059 (N_27059,N_26643,N_26238);
nor U27060 (N_27060,N_25698,N_26024);
nand U27061 (N_27061,N_25831,N_26958);
or U27062 (N_27062,N_26113,N_25945);
xor U27063 (N_27063,N_26774,N_26917);
xor U27064 (N_27064,N_26447,N_25633);
and U27065 (N_27065,N_26087,N_26818);
nand U27066 (N_27066,N_25852,N_26887);
nand U27067 (N_27067,N_26366,N_26824);
xnor U27068 (N_27068,N_26331,N_26575);
and U27069 (N_27069,N_26320,N_26076);
nand U27070 (N_27070,N_25741,N_25764);
or U27071 (N_27071,N_26171,N_26923);
and U27072 (N_27072,N_26822,N_26640);
or U27073 (N_27073,N_26458,N_26422);
nor U27074 (N_27074,N_25744,N_26536);
nor U27075 (N_27075,N_26718,N_26794);
xor U27076 (N_27076,N_25941,N_26831);
xnor U27077 (N_27077,N_26620,N_25649);
xor U27078 (N_27078,N_26545,N_26708);
and U27079 (N_27079,N_26123,N_25750);
nor U27080 (N_27080,N_25913,N_26158);
nor U27081 (N_27081,N_25828,N_26677);
and U27082 (N_27082,N_25585,N_26922);
xor U27083 (N_27083,N_26244,N_25963);
and U27084 (N_27084,N_26769,N_25573);
nand U27085 (N_27085,N_26065,N_26352);
nand U27086 (N_27086,N_25579,N_26118);
nand U27087 (N_27087,N_26503,N_26063);
and U27088 (N_27088,N_25834,N_26185);
nor U27089 (N_27089,N_26833,N_26756);
xor U27090 (N_27090,N_25930,N_26672);
nand U27091 (N_27091,N_26075,N_26594);
and U27092 (N_27092,N_26971,N_26042);
and U27093 (N_27093,N_26776,N_26015);
or U27094 (N_27094,N_25937,N_26104);
nor U27095 (N_27095,N_26499,N_26012);
and U27096 (N_27096,N_26360,N_25959);
xor U27097 (N_27097,N_26431,N_26003);
and U27098 (N_27098,N_26851,N_25902);
nor U27099 (N_27099,N_26834,N_26560);
nor U27100 (N_27100,N_25634,N_26246);
nand U27101 (N_27101,N_26763,N_26669);
nor U27102 (N_27102,N_26405,N_26696);
and U27103 (N_27103,N_26071,N_26977);
xnor U27104 (N_27104,N_26678,N_26214);
or U27105 (N_27105,N_26534,N_25993);
or U27106 (N_27106,N_26568,N_25578);
nand U27107 (N_27107,N_26460,N_26629);
nand U27108 (N_27108,N_26149,N_25950);
nor U27109 (N_27109,N_26930,N_26037);
nand U27110 (N_27110,N_26308,N_26564);
or U27111 (N_27111,N_26021,N_26975);
nand U27112 (N_27112,N_26790,N_25988);
or U27113 (N_27113,N_26239,N_25713);
nor U27114 (N_27114,N_25986,N_26092);
or U27115 (N_27115,N_25689,N_26473);
and U27116 (N_27116,N_26734,N_26663);
nor U27117 (N_27117,N_25817,N_26034);
xnor U27118 (N_27118,N_25549,N_25748);
nand U27119 (N_27119,N_26627,N_26551);
xor U27120 (N_27120,N_25749,N_25931);
or U27121 (N_27121,N_26119,N_26472);
and U27122 (N_27122,N_26179,N_26272);
nor U27123 (N_27123,N_26787,N_26590);
nor U27124 (N_27124,N_25956,N_26695);
nand U27125 (N_27125,N_26924,N_25690);
nand U27126 (N_27126,N_26111,N_25808);
or U27127 (N_27127,N_26559,N_25616);
nor U27128 (N_27128,N_25862,N_25618);
nor U27129 (N_27129,N_26407,N_26842);
and U27130 (N_27130,N_25755,N_26062);
and U27131 (N_27131,N_26941,N_26872);
and U27132 (N_27132,N_26811,N_26363);
xor U27133 (N_27133,N_26013,N_26068);
xor U27134 (N_27134,N_26143,N_25759);
and U27135 (N_27135,N_26871,N_26074);
or U27136 (N_27136,N_26539,N_25832);
or U27137 (N_27137,N_26288,N_26603);
and U27138 (N_27138,N_26595,N_26962);
xor U27139 (N_27139,N_26647,N_25592);
and U27140 (N_27140,N_26699,N_26502);
nor U27141 (N_27141,N_26825,N_26538);
or U27142 (N_27142,N_26314,N_26628);
or U27143 (N_27143,N_26249,N_26217);
nor U27144 (N_27144,N_25628,N_26617);
and U27145 (N_27145,N_25863,N_26929);
xor U27146 (N_27146,N_26578,N_26368);
or U27147 (N_27147,N_26206,N_26322);
nor U27148 (N_27148,N_25533,N_26463);
xnor U27149 (N_27149,N_26132,N_25921);
nand U27150 (N_27150,N_26697,N_25818);
nand U27151 (N_27151,N_26298,N_25676);
xor U27152 (N_27152,N_25933,N_26579);
or U27153 (N_27153,N_26203,N_26440);
xor U27154 (N_27154,N_26488,N_26417);
nor U27155 (N_27155,N_26733,N_26642);
nand U27156 (N_27156,N_26175,N_26455);
and U27157 (N_27157,N_26057,N_25500);
nand U27158 (N_27158,N_25621,N_26775);
or U27159 (N_27159,N_26046,N_26547);
or U27160 (N_27160,N_26318,N_26371);
and U27161 (N_27161,N_26651,N_25942);
or U27162 (N_27162,N_25665,N_26702);
and U27163 (N_27163,N_25606,N_26009);
or U27164 (N_27164,N_26241,N_26840);
or U27165 (N_27165,N_26372,N_26530);
xor U27166 (N_27166,N_26484,N_25757);
xnor U27167 (N_27167,N_25595,N_26465);
nor U27168 (N_27168,N_25789,N_26349);
nand U27169 (N_27169,N_25954,N_26354);
or U27170 (N_27170,N_25881,N_26064);
xor U27171 (N_27171,N_26942,N_25892);
nand U27172 (N_27172,N_25605,N_26164);
and U27173 (N_27173,N_26624,N_26144);
or U27174 (N_27174,N_25928,N_26327);
nor U27175 (N_27175,N_26020,N_25737);
and U27176 (N_27176,N_26665,N_26645);
nor U27177 (N_27177,N_26852,N_26136);
and U27178 (N_27178,N_26739,N_25989);
and U27179 (N_27179,N_26940,N_25836);
nand U27180 (N_27180,N_26928,N_25906);
nor U27181 (N_27181,N_26268,N_26380);
xor U27182 (N_27182,N_25545,N_26483);
nor U27183 (N_27183,N_26891,N_26233);
nand U27184 (N_27184,N_25730,N_26050);
nand U27185 (N_27185,N_26245,N_25919);
nor U27186 (N_27186,N_26480,N_26799);
or U27187 (N_27187,N_26124,N_26543);
xor U27188 (N_27188,N_26425,N_26969);
nor U27189 (N_27189,N_26823,N_26263);
or U27190 (N_27190,N_26556,N_26419);
nand U27191 (N_27191,N_25525,N_26886);
or U27192 (N_27192,N_25693,N_25688);
nor U27193 (N_27193,N_26294,N_26952);
nand U27194 (N_27194,N_25770,N_25920);
and U27195 (N_27195,N_26182,N_26501);
nor U27196 (N_27196,N_25645,N_25720);
or U27197 (N_27197,N_26540,N_26089);
nor U27198 (N_27198,N_25878,N_26990);
nor U27199 (N_27199,N_25765,N_26041);
or U27200 (N_27200,N_25583,N_25827);
and U27201 (N_27201,N_25521,N_26984);
and U27202 (N_27202,N_25974,N_25854);
xor U27203 (N_27203,N_26948,N_25844);
nand U27204 (N_27204,N_26078,N_26229);
and U27205 (N_27205,N_26982,N_26090);
nand U27206 (N_27206,N_26553,N_26943);
or U27207 (N_27207,N_26088,N_25637);
or U27208 (N_27208,N_26370,N_26162);
or U27209 (N_27209,N_26608,N_25619);
and U27210 (N_27210,N_26849,N_26725);
nor U27211 (N_27211,N_26385,N_26999);
nand U27212 (N_27212,N_25857,N_26029);
xnor U27213 (N_27213,N_25795,N_25564);
and U27214 (N_27214,N_26131,N_25880);
xor U27215 (N_27215,N_25802,N_25990);
or U27216 (N_27216,N_25632,N_26988);
and U27217 (N_27217,N_25916,N_26989);
or U27218 (N_27218,N_25635,N_26867);
nor U27219 (N_27219,N_25961,N_25965);
or U27220 (N_27220,N_26112,N_26985);
and U27221 (N_27221,N_25910,N_25641);
xnor U27222 (N_27222,N_25935,N_26587);
or U27223 (N_27223,N_25742,N_26896);
xor U27224 (N_27224,N_25756,N_25815);
xnor U27225 (N_27225,N_25611,N_25904);
xnor U27226 (N_27226,N_25926,N_26670);
and U27227 (N_27227,N_26186,N_26932);
nand U27228 (N_27228,N_26832,N_26637);
or U27229 (N_27229,N_26945,N_26237);
xor U27230 (N_27230,N_25780,N_26378);
nor U27231 (N_27231,N_26522,N_26716);
nand U27232 (N_27232,N_26215,N_26052);
nand U27233 (N_27233,N_25840,N_26690);
and U27234 (N_27234,N_26018,N_26964);
or U27235 (N_27235,N_25687,N_25785);
and U27236 (N_27236,N_25565,N_26646);
nor U27237 (N_27237,N_25537,N_26291);
nand U27238 (N_27238,N_26408,N_26710);
nor U27239 (N_27239,N_26992,N_25957);
nor U27240 (N_27240,N_26657,N_26140);
and U27241 (N_27241,N_26467,N_26765);
or U27242 (N_27242,N_26562,N_26615);
xnor U27243 (N_27243,N_26535,N_26901);
nand U27244 (N_27244,N_26525,N_26202);
xnor U27245 (N_27245,N_26662,N_26618);
nand U27246 (N_27246,N_25853,N_26495);
nand U27247 (N_27247,N_25515,N_26154);
xnor U27248 (N_27248,N_25777,N_26481);
nor U27249 (N_27249,N_25855,N_26793);
and U27250 (N_27250,N_25722,N_26996);
nor U27251 (N_27251,N_26884,N_25985);
nor U27252 (N_27252,N_26938,N_26002);
and U27253 (N_27253,N_26326,N_26772);
and U27254 (N_27254,N_26526,N_26749);
nor U27255 (N_27255,N_25555,N_26532);
or U27256 (N_27256,N_25640,N_26778);
xor U27257 (N_27257,N_26847,N_26743);
and U27258 (N_27258,N_26836,N_26152);
or U27259 (N_27259,N_25886,N_26666);
and U27260 (N_27260,N_25523,N_25775);
or U27261 (N_27261,N_26570,N_26888);
xor U27262 (N_27262,N_25905,N_25783);
and U27263 (N_27263,N_25820,N_26421);
and U27264 (N_27264,N_26821,N_25763);
or U27265 (N_27265,N_26196,N_26897);
xnor U27266 (N_27266,N_26599,N_26748);
xor U27267 (N_27267,N_25949,N_25875);
or U27268 (N_27268,N_26582,N_25528);
nand U27269 (N_27269,N_26683,N_26600);
xnor U27270 (N_27270,N_26729,N_26395);
and U27271 (N_27271,N_26192,N_26622);
nor U27272 (N_27272,N_25554,N_25871);
or U27273 (N_27273,N_25845,N_26648);
nor U27274 (N_27274,N_25672,N_26993);
nand U27275 (N_27275,N_26784,N_26745);
and U27276 (N_27276,N_25519,N_26219);
xor U27277 (N_27277,N_26698,N_26631);
nor U27278 (N_27278,N_26220,N_26626);
xor U27279 (N_27279,N_26814,N_25569);
nand U27280 (N_27280,N_26025,N_25653);
nor U27281 (N_27281,N_26950,N_26638);
nor U27282 (N_27282,N_26333,N_26151);
nand U27283 (N_27283,N_25970,N_26907);
nand U27284 (N_27284,N_26126,N_26486);
nand U27285 (N_27285,N_26542,N_26411);
xor U27286 (N_27286,N_26780,N_26084);
and U27287 (N_27287,N_25932,N_26931);
or U27288 (N_27288,N_26301,N_25890);
xor U27289 (N_27289,N_26554,N_26364);
or U27290 (N_27290,N_26873,N_25882);
nor U27291 (N_27291,N_26325,N_26653);
and U27292 (N_27292,N_26475,N_25900);
xnor U27293 (N_27293,N_26270,N_25768);
nor U27294 (N_27294,N_26788,N_25899);
nand U27295 (N_27295,N_26903,N_26894);
and U27296 (N_27296,N_26361,N_26266);
nand U27297 (N_27297,N_26242,N_26116);
or U27298 (N_27298,N_26040,N_26432);
xor U27299 (N_27299,N_26265,N_26340);
nand U27300 (N_27300,N_26555,N_25729);
xnor U27301 (N_27301,N_25538,N_26226);
nor U27302 (N_27302,N_26255,N_26187);
nor U27303 (N_27303,N_26796,N_26311);
and U27304 (N_27304,N_25709,N_26520);
nor U27305 (N_27305,N_26754,N_26869);
nor U27306 (N_27306,N_26414,N_26625);
and U27307 (N_27307,N_26452,N_25588);
nand U27308 (N_27308,N_26913,N_25939);
or U27309 (N_27309,N_26355,N_26576);
xor U27310 (N_27310,N_25813,N_25799);
or U27311 (N_27311,N_26719,N_26636);
and U27312 (N_27312,N_26469,N_25607);
nand U27313 (N_27313,N_26142,N_25971);
xor U27314 (N_27314,N_26771,N_26485);
nand U27315 (N_27315,N_26507,N_26070);
xor U27316 (N_27316,N_26468,N_25668);
nand U27317 (N_27317,N_26616,N_25774);
nor U27318 (N_27318,N_26519,N_25630);
nor U27319 (N_27319,N_25865,N_25524);
xnor U27320 (N_27320,N_26810,N_25591);
nand U27321 (N_27321,N_26141,N_25710);
xnor U27322 (N_27322,N_25792,N_26879);
nand U27323 (N_27323,N_26330,N_26170);
nand U27324 (N_27324,N_26813,N_25572);
nor U27325 (N_27325,N_25546,N_25502);
and U27326 (N_27326,N_26760,N_26269);
nand U27327 (N_27327,N_26006,N_26176);
or U27328 (N_27328,N_26258,N_25686);
or U27329 (N_27329,N_26954,N_26150);
nor U27330 (N_27330,N_26882,N_25566);
nand U27331 (N_27331,N_25897,N_26949);
nand U27332 (N_27332,N_26448,N_26515);
nor U27333 (N_27333,N_25651,N_26986);
nor U27334 (N_27334,N_25837,N_26429);
xnor U27335 (N_27335,N_26589,N_26462);
xnor U27336 (N_27336,N_26868,N_26367);
nand U27337 (N_27337,N_26630,N_25912);
nor U27338 (N_27338,N_26083,N_25732);
and U27339 (N_27339,N_26261,N_26039);
nand U27340 (N_27340,N_25586,N_26972);
and U27341 (N_27341,N_26049,N_26036);
or U27342 (N_27342,N_25909,N_26509);
or U27343 (N_27343,N_26359,N_26946);
xnor U27344 (N_27344,N_25821,N_25842);
or U27345 (N_27345,N_25508,N_26902);
or U27346 (N_27346,N_25798,N_26786);
or U27347 (N_27347,N_25746,N_26101);
nor U27348 (N_27348,N_25915,N_25700);
xnor U27349 (N_27349,N_26514,N_26285);
or U27350 (N_27350,N_26782,N_26671);
nand U27351 (N_27351,N_26797,N_25790);
xnor U27352 (N_27352,N_26188,N_26351);
and U27353 (N_27353,N_26802,N_26659);
nor U27354 (N_27354,N_26508,N_25929);
and U27355 (N_27355,N_26200,N_26752);
or U27356 (N_27356,N_26376,N_26623);
nand U27357 (N_27357,N_25898,N_26863);
and U27358 (N_27358,N_26365,N_26373);
xor U27359 (N_27359,N_25669,N_26820);
xor U27360 (N_27360,N_26201,N_26260);
and U27361 (N_27361,N_26121,N_26655);
or U27362 (N_27362,N_25703,N_26114);
xor U27363 (N_27363,N_26138,N_26161);
and U27364 (N_27364,N_26766,N_26650);
or U27365 (N_27365,N_25830,N_26965);
nor U27366 (N_27366,N_26434,N_26584);
and U27367 (N_27367,N_25877,N_26236);
nor U27368 (N_27368,N_26883,N_26504);
or U27369 (N_27369,N_26598,N_26957);
nand U27370 (N_27370,N_26439,N_26253);
and U27371 (N_27371,N_25782,N_26676);
and U27372 (N_27372,N_26160,N_25608);
xor U27373 (N_27373,N_25692,N_26218);
and U27374 (N_27374,N_26722,N_26981);
and U27375 (N_27375,N_26108,N_26474);
nor U27376 (N_27376,N_26817,N_25936);
nor U27377 (N_27377,N_25563,N_25711);
or U27378 (N_27378,N_25513,N_26353);
nand U27379 (N_27379,N_26905,N_26290);
or U27380 (N_27380,N_26700,N_25980);
nor U27381 (N_27381,N_26283,N_26248);
xnor U27382 (N_27382,N_26533,N_25869);
nand U27383 (N_27383,N_25858,N_26730);
nand U27384 (N_27384,N_26726,N_26614);
nand U27385 (N_27385,N_26433,N_26335);
nor U27386 (N_27386,N_26047,N_26435);
or U27387 (N_27387,N_26450,N_26956);
nand U27388 (N_27388,N_25846,N_26445);
or U27389 (N_27389,N_26027,N_26302);
xnor U27390 (N_27390,N_26328,N_25816);
nor U27391 (N_27391,N_26795,N_25570);
and U27392 (N_27392,N_26281,N_26208);
nand U27393 (N_27393,N_25867,N_25991);
or U27394 (N_27394,N_25663,N_25683);
nor U27395 (N_27395,N_26909,N_26921);
or U27396 (N_27396,N_26859,N_26190);
and U27397 (N_27397,N_25797,N_26939);
or U27398 (N_27398,N_25835,N_25812);
and U27399 (N_27399,N_25719,N_25983);
nor U27400 (N_27400,N_25751,N_26082);
nand U27401 (N_27401,N_25784,N_25678);
xor U27402 (N_27402,N_25577,N_26426);
xor U27403 (N_27403,N_26044,N_25781);
nand U27404 (N_27404,N_26714,N_26919);
or U27405 (N_27405,N_25728,N_26505);
or U27406 (N_27406,N_26023,N_26926);
xor U27407 (N_27407,N_26135,N_25544);
and U27408 (N_27408,N_25955,N_25679);
or U27409 (N_27409,N_25885,N_26740);
or U27410 (N_27410,N_26558,N_26815);
or U27411 (N_27411,N_25512,N_26994);
nand U27412 (N_27412,N_26436,N_26490);
nand U27413 (N_27413,N_25833,N_26345);
nor U27414 (N_27414,N_25560,N_25530);
nor U27415 (N_27415,N_26148,N_25873);
xor U27416 (N_27416,N_26310,N_26967);
nor U27417 (N_27417,N_26457,N_26974);
and U27418 (N_27418,N_26316,N_26881);
xnor U27419 (N_27419,N_25810,N_26607);
and U27420 (N_27420,N_26221,N_26935);
xor U27421 (N_27421,N_26271,N_26341);
and U27422 (N_27422,N_25580,N_26397);
nand U27423 (N_27423,N_26343,N_26388);
or U27424 (N_27424,N_25594,N_25776);
or U27425 (N_27425,N_26978,N_26966);
or U27426 (N_27426,N_25925,N_25705);
nand U27427 (N_27427,N_25617,N_25505);
or U27428 (N_27428,N_26128,N_26362);
or U27429 (N_27429,N_26172,N_26110);
or U27430 (N_27430,N_25940,N_26224);
nor U27431 (N_27431,N_26130,N_25725);
nand U27432 (N_27432,N_26593,N_26658);
xnor U27433 (N_27433,N_26085,N_25656);
xor U27434 (N_27434,N_25889,N_26139);
nand U27435 (N_27435,N_26944,N_25870);
xor U27436 (N_27436,N_25576,N_26955);
nor U27437 (N_27437,N_26963,N_26707);
xor U27438 (N_27438,N_25610,N_26303);
or U27439 (N_27439,N_25714,N_26512);
xnor U27440 (N_27440,N_26908,N_26529);
nand U27441 (N_27441,N_26588,N_25747);
and U27442 (N_27442,N_25981,N_26674);
xor U27443 (N_27443,N_26441,N_25599);
or U27444 (N_27444,N_25819,N_26392);
nand U27445 (N_27445,N_26997,N_26937);
and U27446 (N_27446,N_25934,N_26409);
nand U27447 (N_27447,N_26494,N_26016);
or U27448 (N_27448,N_26621,N_26240);
xor U27449 (N_27449,N_26391,N_25522);
and U27450 (N_27450,N_25553,N_26511);
and U27451 (N_27451,N_26686,N_26048);
and U27452 (N_27452,N_25953,N_26893);
or U27453 (N_27453,N_25982,N_26830);
or U27454 (N_27454,N_26033,N_25501);
nand U27455 (N_27455,N_26058,N_26864);
and U27456 (N_27456,N_25992,N_26792);
or U27457 (N_27457,N_26925,N_25996);
or U27458 (N_27458,N_25527,N_25761);
xor U27459 (N_27459,N_26552,N_26701);
and U27460 (N_27460,N_26639,N_26761);
or U27461 (N_27461,N_25740,N_26383);
nand U27462 (N_27462,N_25535,N_25895);
nand U27463 (N_27463,N_25644,N_25767);
xor U27464 (N_27464,N_26580,N_26980);
nand U27465 (N_27465,N_26004,N_26731);
and U27466 (N_27466,N_26850,N_25743);
nor U27467 (N_27467,N_25887,N_26147);
nand U27468 (N_27468,N_26606,N_26632);
nand U27469 (N_27469,N_26783,N_26611);
xor U27470 (N_27470,N_25598,N_26968);
nor U27471 (N_27471,N_26826,N_26764);
or U27472 (N_27472,N_26528,N_26844);
xnor U27473 (N_27473,N_26641,N_26410);
nand U27474 (N_27474,N_25694,N_26853);
nand U27475 (N_27475,N_26976,N_26915);
xnor U27476 (N_27476,N_26398,N_25541);
xnor U27477 (N_27477,N_25529,N_26934);
nand U27478 (N_27478,N_26273,N_25946);
or U27479 (N_27479,N_26225,N_26256);
xnor U27480 (N_27480,N_26936,N_26133);
or U27481 (N_27481,N_26482,N_25695);
and U27482 (N_27482,N_26605,N_25518);
nand U27483 (N_27483,N_26193,N_25951);
nor U27484 (N_27484,N_26694,N_26741);
nand U27485 (N_27485,N_26077,N_26262);
xor U27486 (N_27486,N_25590,N_25738);
or U27487 (N_27487,N_26315,N_26591);
nand U27488 (N_27488,N_26675,N_25718);
nor U27489 (N_27489,N_26107,N_26211);
nand U27490 (N_27490,N_26001,N_25603);
nand U27491 (N_27491,N_26846,N_26323);
nand U27492 (N_27492,N_26768,N_26757);
or U27493 (N_27493,N_26420,N_25786);
nor U27494 (N_27494,N_25893,N_26998);
xnor U27495 (N_27495,N_26183,N_25908);
or U27496 (N_27496,N_26094,N_25655);
nor U27497 (N_27497,N_26633,N_26518);
and U27498 (N_27498,N_25856,N_26155);
nor U27499 (N_27499,N_26819,N_26737);
nand U27500 (N_27500,N_26251,N_26916);
xor U27501 (N_27501,N_26758,N_26276);
nand U27502 (N_27502,N_25814,N_26602);
nor U27503 (N_27503,N_26103,N_25684);
and U27504 (N_27504,N_26773,N_26377);
xnor U27505 (N_27505,N_25734,N_26356);
xor U27506 (N_27506,N_25532,N_26073);
nor U27507 (N_27507,N_25510,N_25766);
nand U27508 (N_27508,N_26232,N_26060);
nand U27509 (N_27509,N_26145,N_25604);
nor U27510 (N_27510,N_26687,N_26750);
nor U27511 (N_27511,N_26309,N_26093);
xnor U27512 (N_27512,N_26736,N_26061);
nor U27513 (N_27513,N_25575,N_25643);
xor U27514 (N_27514,N_25947,N_26427);
nor U27515 (N_27515,N_26911,N_26876);
or U27516 (N_27516,N_26418,N_25891);
and U27517 (N_27517,N_26010,N_26091);
nand U27518 (N_27518,N_26874,N_26567);
or U27519 (N_27519,N_25975,N_25829);
nor U27520 (N_27520,N_26709,N_25624);
xnor U27521 (N_27521,N_26527,N_26344);
xor U27522 (N_27522,N_25514,N_25771);
and U27523 (N_27523,N_26295,N_25736);
or U27524 (N_27524,N_26477,N_25631);
xor U27525 (N_27525,N_25801,N_26404);
nor U27526 (N_27526,N_26231,N_26334);
or U27527 (N_27527,N_26443,N_26899);
nor U27528 (N_27528,N_26660,N_26688);
or U27529 (N_27529,N_26028,N_25806);
nand U27530 (N_27530,N_26127,N_26178);
xnor U27531 (N_27531,N_26428,N_25506);
or U27532 (N_27532,N_26293,N_25745);
or U27533 (N_27533,N_26720,N_25557);
or U27534 (N_27534,N_25601,N_25613);
nand U27535 (N_27535,N_26278,N_26174);
nand U27536 (N_27536,N_26019,N_26544);
xor U27537 (N_27537,N_25639,N_26586);
or U27538 (N_27538,N_26713,N_26223);
nor U27539 (N_27539,N_26829,N_25561);
xor U27540 (N_27540,N_25708,N_26337);
or U27541 (N_27541,N_26035,N_26097);
nand U27542 (N_27542,N_25662,N_26837);
xor U27543 (N_27543,N_25702,N_26493);
xor U27544 (N_27544,N_26459,N_26791);
and U27545 (N_27545,N_26098,N_26991);
or U27546 (N_27546,N_25872,N_25642);
nor U27547 (N_27547,N_26933,N_26210);
xor U27548 (N_27548,N_25999,N_26252);
nor U27549 (N_27549,N_26297,N_26644);
or U27550 (N_27550,N_26051,N_25938);
or U27551 (N_27551,N_26951,N_25944);
or U27552 (N_27552,N_25509,N_25978);
xnor U27553 (N_27553,N_25548,N_26109);
or U27554 (N_27554,N_26129,N_25772);
nand U27555 (N_27555,N_26199,N_26496);
or U27556 (N_27556,N_26342,N_26120);
nand U27557 (N_27557,N_26995,N_26717);
or U27558 (N_27558,N_26523,N_25773);
or U27559 (N_27559,N_26069,N_25620);
and U27560 (N_27560,N_25779,N_26715);
nor U27561 (N_27561,N_26596,N_26329);
nor U27562 (N_27562,N_25534,N_26446);
or U27563 (N_27563,N_26856,N_26189);
xnor U27564 (N_27564,N_26180,N_26571);
nand U27565 (N_27565,N_25794,N_26979);
nand U27566 (N_27566,N_26489,N_26358);
nand U27567 (N_27567,N_25567,N_26346);
nor U27568 (N_27568,N_26000,N_26742);
or U27569 (N_27569,N_26207,N_25602);
nand U27570 (N_27570,N_25825,N_26413);
and U27571 (N_27571,N_26581,N_25850);
or U27572 (N_27572,N_26835,N_25681);
xnor U27573 (N_27573,N_26393,N_25574);
or U27574 (N_27574,N_26324,N_26163);
xor U27575 (N_27575,N_26689,N_25571);
nor U27576 (N_27576,N_26054,N_26561);
nor U27577 (N_27577,N_26541,N_26759);
nand U27578 (N_27578,N_26500,N_25597);
nand U27579 (N_27579,N_26789,N_26115);
or U27580 (N_27580,N_26382,N_25701);
nand U27581 (N_27581,N_25851,N_26920);
nand U27582 (N_27582,N_26870,N_25593);
nor U27583 (N_27583,N_26279,N_26197);
or U27584 (N_27584,N_26286,N_26031);
or U27585 (N_27585,N_26548,N_26277);
nand U27586 (N_27586,N_25973,N_26634);
nand U27587 (N_27587,N_26304,N_25706);
or U27588 (N_27588,N_26601,N_26191);
nor U27589 (N_27589,N_26808,N_25918);
xnor U27590 (N_27590,N_26885,N_26524);
or U27591 (N_27591,N_26007,N_25581);
xnor U27592 (N_27592,N_25952,N_25715);
and U27593 (N_27593,N_26332,N_25788);
or U27594 (N_27594,N_25697,N_26684);
nand U27595 (N_27595,N_25809,N_25866);
or U27596 (N_27596,N_25778,N_25927);
or U27597 (N_27597,N_26597,N_25807);
nand U27598 (N_27598,N_26681,N_26102);
or U27599 (N_27599,N_25823,N_26134);
nand U27600 (N_27600,N_26400,N_26389);
and U27601 (N_27601,N_25520,N_25979);
or U27602 (N_27602,N_26724,N_26339);
and U27603 (N_27603,N_26566,N_26451);
nand U27604 (N_27604,N_26195,N_26204);
nand U27605 (N_27605,N_25661,N_25612);
xnor U27606 (N_27606,N_26865,N_26476);
nand U27607 (N_27607,N_25623,N_25542);
nor U27608 (N_27608,N_26166,N_26732);
and U27609 (N_27609,N_26613,N_26723);
nor U27610 (N_27610,N_25997,N_25754);
or U27611 (N_27611,N_26423,N_26738);
and U27612 (N_27612,N_25511,N_26727);
xor U27613 (N_27613,N_26464,N_26011);
xnor U27614 (N_27614,N_25903,N_25559);
nor U27615 (N_27615,N_25769,N_26259);
or U27616 (N_27616,N_26574,N_25838);
nor U27617 (N_27617,N_26307,N_26668);
or U27618 (N_27618,N_25962,N_25716);
or U27619 (N_27619,N_26106,N_25712);
nor U27620 (N_27620,N_26892,N_26374);
nand U27621 (N_27621,N_26857,N_25861);
and U27622 (N_27622,N_26510,N_26387);
nand U27623 (N_27623,N_26338,N_26809);
nor U27624 (N_27624,N_26228,N_25696);
nand U27625 (N_27625,N_25659,N_26572);
and U27626 (N_27626,N_25551,N_26022);
nand U27627 (N_27627,N_26396,N_25864);
or U27628 (N_27628,N_26292,N_25896);
nand U27629 (N_27629,N_25876,N_26100);
and U27630 (N_27630,N_25739,N_26747);
or U27631 (N_27631,N_26711,N_26592);
nor U27632 (N_27632,N_26319,N_25675);
xnor U27633 (N_27633,N_26454,N_25724);
nand U27634 (N_27634,N_25504,N_25735);
and U27635 (N_27635,N_25539,N_26661);
nand U27636 (N_27636,N_26275,N_26079);
nor U27637 (N_27637,N_26177,N_26801);
nand U27638 (N_27638,N_26953,N_25674);
nand U27639 (N_27639,N_26466,N_25638);
or U27640 (N_27640,N_26679,N_25966);
nand U27641 (N_27641,N_26479,N_26744);
and U27642 (N_27642,N_25587,N_26384);
and U27643 (N_27643,N_25726,N_26216);
nor U27644 (N_27644,N_26444,N_26375);
xnor U27645 (N_27645,N_26086,N_26096);
nand U27646 (N_27646,N_26403,N_26017);
nor U27647 (N_27647,N_26583,N_26348);
and U27648 (N_27648,N_26712,N_25995);
and U27649 (N_27649,N_26321,N_26424);
or U27650 (N_27650,N_25911,N_25883);
or U27651 (N_27651,N_26243,N_26704);
and U27652 (N_27652,N_26105,N_26904);
and U27653 (N_27653,N_26184,N_26828);
nand U27654 (N_27654,N_26721,N_25657);
nand U27655 (N_27655,N_26312,N_26800);
xor U27656 (N_27656,N_26827,N_25943);
xor U27657 (N_27657,N_26673,N_25526);
or U27658 (N_27658,N_26753,N_25671);
nand U27659 (N_27659,N_26947,N_26213);
nand U27660 (N_27660,N_26492,N_25948);
or U27661 (N_27661,N_26585,N_25972);
and U27662 (N_27662,N_26254,N_26399);
and U27663 (N_27663,N_26838,N_26430);
or U27664 (N_27664,N_25721,N_26026);
xor U27665 (N_27665,N_25760,N_26461);
or U27666 (N_27666,N_25787,N_26173);
or U27667 (N_27667,N_26890,N_26806);
xor U27668 (N_27668,N_25977,N_25849);
xor U27669 (N_27669,N_25614,N_25848);
and U27670 (N_27670,N_25879,N_26563);
nor U27671 (N_27671,N_25805,N_26906);
xnor U27672 (N_27672,N_26401,N_25901);
nor U27673 (N_27673,N_25652,N_26610);
xnor U27674 (N_27674,N_25667,N_25917);
nor U27675 (N_27675,N_26478,N_25596);
or U27676 (N_27676,N_26350,N_25960);
or U27677 (N_27677,N_25531,N_26549);
xnor U27678 (N_27678,N_26379,N_26470);
nor U27679 (N_27679,N_26878,N_25658);
and U27680 (N_27680,N_26067,N_25803);
or U27681 (N_27681,N_25998,N_26807);
nand U27682 (N_27682,N_26072,N_26212);
nor U27683 (N_27683,N_26169,N_26877);
nor U27684 (N_27684,N_26550,N_25884);
nand U27685 (N_27685,N_25636,N_26014);
nor U27686 (N_27686,N_26839,N_26959);
or U27687 (N_27687,N_26095,N_26406);
xor U27688 (N_27688,N_26153,N_25967);
xor U27689 (N_27689,N_25648,N_26812);
or U27690 (N_27690,N_26848,N_26137);
and U27691 (N_27691,N_26573,N_26973);
and U27692 (N_27692,N_26516,N_25629);
nor U27693 (N_27693,N_25682,N_26604);
nand U27694 (N_27694,N_25894,N_26274);
and U27695 (N_27695,N_25968,N_26045);
and U27696 (N_27696,N_26053,N_26282);
xor U27697 (N_27697,N_25874,N_26861);
or U27698 (N_27698,N_25650,N_26402);
nand U27699 (N_27699,N_26306,N_25685);
nand U27700 (N_27700,N_26167,N_26146);
nor U27701 (N_27701,N_26038,N_25796);
nor U27702 (N_27702,N_26914,N_26866);
nand U27703 (N_27703,N_26287,N_25914);
nand U27704 (N_27704,N_25843,N_26117);
or U27705 (N_27705,N_26652,N_26691);
nor U27706 (N_27706,N_25615,N_25800);
nand U27707 (N_27707,N_25723,N_25654);
nand U27708 (N_27708,N_26751,N_26222);
xor U27709 (N_27709,N_25984,N_26381);
nand U27710 (N_27710,N_25976,N_26198);
and U27711 (N_27711,N_26854,N_26449);
and U27712 (N_27712,N_26357,N_26654);
nand U27713 (N_27713,N_25907,N_25589);
xor U27714 (N_27714,N_25822,N_25839);
nand U27715 (N_27715,N_26912,N_26235);
and U27716 (N_27716,N_26889,N_26209);
nand U27717 (N_27717,N_26656,N_26537);
xnor U27718 (N_27718,N_25600,N_26456);
or U27719 (N_27719,N_25727,N_25550);
or U27720 (N_27720,N_26680,N_25584);
and U27721 (N_27721,N_26785,N_26565);
and U27722 (N_27722,N_26781,N_26706);
nand U27723 (N_27723,N_26099,N_25552);
or U27724 (N_27724,N_26416,N_26612);
nor U27725 (N_27725,N_25562,N_26855);
and U27726 (N_27726,N_26390,N_26415);
xor U27727 (N_27727,N_25824,N_26165);
or U27728 (N_27728,N_26317,N_25793);
and U27729 (N_27729,N_26910,N_26247);
xnor U27730 (N_27730,N_26609,N_26860);
and U27731 (N_27731,N_25847,N_26577);
nor U27732 (N_27732,N_25868,N_25691);
nor U27733 (N_27733,N_26841,N_25987);
or U27734 (N_27734,N_25547,N_26762);
xnor U27735 (N_27735,N_26960,N_26437);
and U27736 (N_27736,N_26875,N_26059);
nor U27737 (N_27737,N_25923,N_26798);
and U27738 (N_27738,N_25704,N_26471);
nor U27739 (N_27739,N_26898,N_25517);
and U27740 (N_27740,N_25731,N_26498);
or U27741 (N_27741,N_26300,N_25717);
and U27742 (N_27742,N_25540,N_25558);
nor U27743 (N_27743,N_26619,N_25733);
or U27744 (N_27744,N_26735,N_26927);
nand U27745 (N_27745,N_25924,N_26703);
nor U27746 (N_27746,N_26770,N_25791);
and U27747 (N_27747,N_26005,N_25556);
or U27748 (N_27748,N_26755,N_26805);
and U27749 (N_27749,N_25666,N_26156);
and U27750 (N_27750,N_25571,N_26082);
and U27751 (N_27751,N_26440,N_26710);
nor U27752 (N_27752,N_26220,N_26581);
xnor U27753 (N_27753,N_26274,N_25586);
nor U27754 (N_27754,N_26335,N_26464);
or U27755 (N_27755,N_25609,N_26638);
xor U27756 (N_27756,N_26698,N_26153);
or U27757 (N_27757,N_26208,N_25970);
nor U27758 (N_27758,N_26293,N_26811);
xor U27759 (N_27759,N_26142,N_26836);
xor U27760 (N_27760,N_25914,N_26233);
xnor U27761 (N_27761,N_26853,N_25948);
nor U27762 (N_27762,N_26866,N_25939);
and U27763 (N_27763,N_26847,N_26878);
or U27764 (N_27764,N_26579,N_26793);
xor U27765 (N_27765,N_25520,N_25981);
xor U27766 (N_27766,N_26015,N_25985);
xor U27767 (N_27767,N_26953,N_25585);
nand U27768 (N_27768,N_25778,N_26856);
and U27769 (N_27769,N_26278,N_25596);
nor U27770 (N_27770,N_26969,N_26142);
and U27771 (N_27771,N_26471,N_25522);
and U27772 (N_27772,N_26043,N_25938);
or U27773 (N_27773,N_26283,N_25659);
xor U27774 (N_27774,N_25937,N_26180);
nand U27775 (N_27775,N_25858,N_25625);
xnor U27776 (N_27776,N_26846,N_25595);
xnor U27777 (N_27777,N_26673,N_26935);
nor U27778 (N_27778,N_26442,N_26412);
and U27779 (N_27779,N_26619,N_25633);
nor U27780 (N_27780,N_25501,N_25610);
xnor U27781 (N_27781,N_26462,N_26050);
nor U27782 (N_27782,N_26324,N_26570);
and U27783 (N_27783,N_26888,N_26567);
xor U27784 (N_27784,N_26853,N_25973);
or U27785 (N_27785,N_26820,N_26685);
and U27786 (N_27786,N_26336,N_26091);
or U27787 (N_27787,N_25652,N_25934);
nor U27788 (N_27788,N_26271,N_26811);
or U27789 (N_27789,N_26596,N_26406);
nand U27790 (N_27790,N_26355,N_26310);
xor U27791 (N_27791,N_26105,N_26532);
and U27792 (N_27792,N_26458,N_26939);
nand U27793 (N_27793,N_26485,N_26544);
nor U27794 (N_27794,N_26465,N_26912);
and U27795 (N_27795,N_26493,N_25739);
nor U27796 (N_27796,N_25539,N_26329);
nor U27797 (N_27797,N_25605,N_25745);
or U27798 (N_27798,N_26879,N_26529);
and U27799 (N_27799,N_25531,N_25777);
or U27800 (N_27800,N_26500,N_26398);
xnor U27801 (N_27801,N_25982,N_26795);
nand U27802 (N_27802,N_26132,N_26442);
or U27803 (N_27803,N_26197,N_25837);
nand U27804 (N_27804,N_26631,N_25577);
nor U27805 (N_27805,N_26896,N_25946);
and U27806 (N_27806,N_26465,N_26447);
xnor U27807 (N_27807,N_25557,N_26366);
and U27808 (N_27808,N_26120,N_25569);
xor U27809 (N_27809,N_26571,N_26812);
nand U27810 (N_27810,N_26037,N_25734);
nand U27811 (N_27811,N_26362,N_26977);
and U27812 (N_27812,N_26862,N_26752);
or U27813 (N_27813,N_26752,N_26527);
or U27814 (N_27814,N_26708,N_26505);
nand U27815 (N_27815,N_26896,N_26796);
nor U27816 (N_27816,N_26238,N_25822);
nand U27817 (N_27817,N_26766,N_26561);
or U27818 (N_27818,N_26554,N_26927);
nor U27819 (N_27819,N_25884,N_25912);
and U27820 (N_27820,N_26137,N_25901);
and U27821 (N_27821,N_25862,N_26081);
xnor U27822 (N_27822,N_26014,N_26288);
or U27823 (N_27823,N_26784,N_26911);
nand U27824 (N_27824,N_25505,N_26659);
nand U27825 (N_27825,N_26762,N_26601);
nor U27826 (N_27826,N_26648,N_26154);
and U27827 (N_27827,N_26436,N_26386);
xor U27828 (N_27828,N_26201,N_25653);
xor U27829 (N_27829,N_25599,N_26272);
xnor U27830 (N_27830,N_26068,N_25738);
nor U27831 (N_27831,N_25853,N_25989);
nor U27832 (N_27832,N_25702,N_25819);
and U27833 (N_27833,N_25685,N_25838);
or U27834 (N_27834,N_26460,N_26618);
or U27835 (N_27835,N_26805,N_26629);
xnor U27836 (N_27836,N_25788,N_25765);
and U27837 (N_27837,N_26502,N_25919);
nor U27838 (N_27838,N_26842,N_26208);
and U27839 (N_27839,N_26414,N_25714);
xor U27840 (N_27840,N_26642,N_26060);
or U27841 (N_27841,N_26279,N_26181);
xnor U27842 (N_27842,N_26692,N_25792);
nor U27843 (N_27843,N_25705,N_26573);
or U27844 (N_27844,N_26270,N_25809);
xnor U27845 (N_27845,N_25730,N_25623);
and U27846 (N_27846,N_26207,N_25700);
or U27847 (N_27847,N_26627,N_26118);
and U27848 (N_27848,N_26426,N_25779);
nor U27849 (N_27849,N_26482,N_26593);
and U27850 (N_27850,N_25514,N_25510);
nor U27851 (N_27851,N_26830,N_25902);
nor U27852 (N_27852,N_25896,N_26764);
xnor U27853 (N_27853,N_26103,N_26707);
nand U27854 (N_27854,N_26975,N_26118);
xnor U27855 (N_27855,N_26003,N_26121);
xor U27856 (N_27856,N_25750,N_26203);
or U27857 (N_27857,N_26506,N_26520);
or U27858 (N_27858,N_26635,N_25638);
nor U27859 (N_27859,N_25980,N_26160);
xor U27860 (N_27860,N_26969,N_25831);
nor U27861 (N_27861,N_26648,N_25782);
and U27862 (N_27862,N_26364,N_26040);
and U27863 (N_27863,N_26739,N_25645);
nor U27864 (N_27864,N_25500,N_25537);
xnor U27865 (N_27865,N_26656,N_26940);
or U27866 (N_27866,N_26967,N_25988);
xnor U27867 (N_27867,N_26844,N_26059);
xnor U27868 (N_27868,N_25581,N_26149);
nor U27869 (N_27869,N_26461,N_25585);
nand U27870 (N_27870,N_26216,N_26704);
or U27871 (N_27871,N_26807,N_26587);
or U27872 (N_27872,N_26998,N_26065);
nand U27873 (N_27873,N_26916,N_26133);
and U27874 (N_27874,N_25617,N_26590);
nor U27875 (N_27875,N_26285,N_26978);
or U27876 (N_27876,N_25782,N_25750);
nand U27877 (N_27877,N_26302,N_26994);
or U27878 (N_27878,N_26663,N_26863);
nor U27879 (N_27879,N_26487,N_26698);
nand U27880 (N_27880,N_26290,N_26816);
or U27881 (N_27881,N_26483,N_26699);
nand U27882 (N_27882,N_26048,N_26987);
and U27883 (N_27883,N_26602,N_26754);
xor U27884 (N_27884,N_25699,N_26463);
and U27885 (N_27885,N_26383,N_25534);
or U27886 (N_27886,N_25673,N_26632);
and U27887 (N_27887,N_26082,N_26377);
nand U27888 (N_27888,N_25902,N_25988);
or U27889 (N_27889,N_26972,N_26454);
xor U27890 (N_27890,N_26589,N_26332);
nor U27891 (N_27891,N_26465,N_26118);
nand U27892 (N_27892,N_25651,N_25979);
nand U27893 (N_27893,N_25625,N_26932);
or U27894 (N_27894,N_26687,N_25691);
nor U27895 (N_27895,N_26496,N_25845);
nor U27896 (N_27896,N_26013,N_26127);
nand U27897 (N_27897,N_26245,N_26399);
and U27898 (N_27898,N_26646,N_26187);
nor U27899 (N_27899,N_26051,N_25675);
nand U27900 (N_27900,N_26256,N_25551);
or U27901 (N_27901,N_25578,N_25796);
xnor U27902 (N_27902,N_26892,N_25901);
or U27903 (N_27903,N_25814,N_26842);
xor U27904 (N_27904,N_26069,N_25635);
nand U27905 (N_27905,N_25823,N_26629);
xnor U27906 (N_27906,N_26879,N_25839);
nor U27907 (N_27907,N_26532,N_26125);
xor U27908 (N_27908,N_26574,N_25538);
or U27909 (N_27909,N_26863,N_25588);
xnor U27910 (N_27910,N_25676,N_25874);
nand U27911 (N_27911,N_25801,N_26449);
xor U27912 (N_27912,N_25674,N_25796);
nor U27913 (N_27913,N_26310,N_26093);
nor U27914 (N_27914,N_26654,N_25900);
nor U27915 (N_27915,N_26976,N_25794);
nand U27916 (N_27916,N_26309,N_25908);
nor U27917 (N_27917,N_26570,N_26875);
or U27918 (N_27918,N_25738,N_26510);
or U27919 (N_27919,N_26493,N_26472);
or U27920 (N_27920,N_26109,N_26836);
xor U27921 (N_27921,N_26744,N_26563);
xor U27922 (N_27922,N_26200,N_26441);
nand U27923 (N_27923,N_26172,N_25750);
xor U27924 (N_27924,N_25614,N_26022);
or U27925 (N_27925,N_26109,N_26488);
or U27926 (N_27926,N_26247,N_25655);
xnor U27927 (N_27927,N_26921,N_26284);
or U27928 (N_27928,N_26726,N_26649);
nor U27929 (N_27929,N_26203,N_25865);
and U27930 (N_27930,N_26815,N_26346);
nor U27931 (N_27931,N_26077,N_26316);
nand U27932 (N_27932,N_26214,N_25779);
or U27933 (N_27933,N_26581,N_26606);
or U27934 (N_27934,N_25514,N_26129);
or U27935 (N_27935,N_26123,N_26636);
nand U27936 (N_27936,N_25539,N_26457);
and U27937 (N_27937,N_26736,N_26991);
xor U27938 (N_27938,N_25957,N_26082);
nor U27939 (N_27939,N_25500,N_25815);
nand U27940 (N_27940,N_26422,N_25671);
or U27941 (N_27941,N_25912,N_26511);
nor U27942 (N_27942,N_26564,N_26056);
nand U27943 (N_27943,N_25713,N_26841);
or U27944 (N_27944,N_26937,N_26538);
nor U27945 (N_27945,N_26519,N_25834);
nor U27946 (N_27946,N_25802,N_26419);
nand U27947 (N_27947,N_26108,N_26730);
nor U27948 (N_27948,N_26887,N_25924);
or U27949 (N_27949,N_26775,N_25774);
nand U27950 (N_27950,N_26432,N_26398);
xnor U27951 (N_27951,N_25895,N_25711);
and U27952 (N_27952,N_26683,N_26206);
and U27953 (N_27953,N_26718,N_26210);
xor U27954 (N_27954,N_26174,N_26823);
nand U27955 (N_27955,N_26249,N_25655);
and U27956 (N_27956,N_26398,N_25795);
nor U27957 (N_27957,N_26139,N_26206);
xor U27958 (N_27958,N_26682,N_25864);
or U27959 (N_27959,N_26349,N_25715);
nor U27960 (N_27960,N_26992,N_25687);
nor U27961 (N_27961,N_26247,N_26032);
nor U27962 (N_27962,N_26696,N_25824);
nor U27963 (N_27963,N_25832,N_26746);
nor U27964 (N_27964,N_25696,N_25662);
nor U27965 (N_27965,N_26460,N_26186);
or U27966 (N_27966,N_26750,N_26395);
or U27967 (N_27967,N_25504,N_26840);
nor U27968 (N_27968,N_26786,N_25913);
nand U27969 (N_27969,N_25641,N_25840);
xor U27970 (N_27970,N_26746,N_26066);
and U27971 (N_27971,N_26616,N_25968);
and U27972 (N_27972,N_25865,N_26384);
nand U27973 (N_27973,N_25731,N_26308);
nand U27974 (N_27974,N_26468,N_26702);
nor U27975 (N_27975,N_26011,N_26515);
xnor U27976 (N_27976,N_25888,N_26293);
xnor U27977 (N_27977,N_26502,N_26406);
nand U27978 (N_27978,N_25863,N_26431);
nand U27979 (N_27979,N_25875,N_26474);
nand U27980 (N_27980,N_26433,N_25978);
nor U27981 (N_27981,N_25564,N_25893);
nor U27982 (N_27982,N_26132,N_26403);
or U27983 (N_27983,N_25852,N_25549);
or U27984 (N_27984,N_26867,N_25634);
nor U27985 (N_27985,N_25625,N_25911);
nor U27986 (N_27986,N_26588,N_26893);
and U27987 (N_27987,N_25938,N_26086);
or U27988 (N_27988,N_25828,N_26410);
xnor U27989 (N_27989,N_26655,N_26739);
nor U27990 (N_27990,N_26673,N_25568);
nor U27991 (N_27991,N_26852,N_25550);
or U27992 (N_27992,N_26986,N_25667);
and U27993 (N_27993,N_26359,N_25997);
or U27994 (N_27994,N_26812,N_26293);
xor U27995 (N_27995,N_25718,N_25861);
and U27996 (N_27996,N_26425,N_25622);
or U27997 (N_27997,N_26744,N_26444);
and U27998 (N_27998,N_26350,N_26218);
nor U27999 (N_27999,N_25880,N_25934);
nand U28000 (N_28000,N_26096,N_25860);
nor U28001 (N_28001,N_25591,N_25715);
nand U28002 (N_28002,N_25698,N_25901);
or U28003 (N_28003,N_26097,N_26326);
xnor U28004 (N_28004,N_26986,N_25557);
nand U28005 (N_28005,N_26556,N_26660);
nor U28006 (N_28006,N_25697,N_25848);
and U28007 (N_28007,N_26067,N_26469);
nor U28008 (N_28008,N_26987,N_26303);
or U28009 (N_28009,N_25707,N_26872);
xor U28010 (N_28010,N_25794,N_26195);
xor U28011 (N_28011,N_26457,N_26512);
nor U28012 (N_28012,N_26970,N_26178);
and U28013 (N_28013,N_26583,N_26249);
and U28014 (N_28014,N_26905,N_26715);
xor U28015 (N_28015,N_25584,N_26339);
or U28016 (N_28016,N_25525,N_25709);
xnor U28017 (N_28017,N_26854,N_26837);
nor U28018 (N_28018,N_25890,N_25563);
nor U28019 (N_28019,N_26046,N_26896);
or U28020 (N_28020,N_25653,N_26931);
xor U28021 (N_28021,N_26512,N_25754);
or U28022 (N_28022,N_26812,N_26487);
nand U28023 (N_28023,N_26116,N_26893);
nand U28024 (N_28024,N_26422,N_25594);
or U28025 (N_28025,N_26847,N_26221);
xnor U28026 (N_28026,N_26185,N_26300);
nor U28027 (N_28027,N_25586,N_25929);
and U28028 (N_28028,N_25777,N_25891);
and U28029 (N_28029,N_26816,N_26944);
nand U28030 (N_28030,N_26596,N_26327);
xnor U28031 (N_28031,N_25687,N_26512);
and U28032 (N_28032,N_26150,N_25500);
or U28033 (N_28033,N_26483,N_26050);
nand U28034 (N_28034,N_26221,N_25675);
xnor U28035 (N_28035,N_25628,N_26229);
or U28036 (N_28036,N_26391,N_26898);
and U28037 (N_28037,N_25635,N_26306);
xnor U28038 (N_28038,N_25539,N_25528);
nand U28039 (N_28039,N_26020,N_26255);
xor U28040 (N_28040,N_26763,N_26371);
xnor U28041 (N_28041,N_25732,N_25605);
xnor U28042 (N_28042,N_25998,N_25526);
or U28043 (N_28043,N_26335,N_26449);
xnor U28044 (N_28044,N_26297,N_25888);
and U28045 (N_28045,N_26856,N_26509);
or U28046 (N_28046,N_26381,N_25880);
nor U28047 (N_28047,N_25797,N_26737);
and U28048 (N_28048,N_25702,N_25952);
nand U28049 (N_28049,N_26003,N_26019);
xor U28050 (N_28050,N_25773,N_26778);
xor U28051 (N_28051,N_26667,N_26954);
xnor U28052 (N_28052,N_26638,N_25685);
xnor U28053 (N_28053,N_26803,N_25610);
nand U28054 (N_28054,N_26031,N_25971);
nand U28055 (N_28055,N_26963,N_26524);
and U28056 (N_28056,N_26718,N_26615);
xnor U28057 (N_28057,N_25882,N_26946);
or U28058 (N_28058,N_25896,N_26011);
nor U28059 (N_28059,N_26178,N_26383);
xnor U28060 (N_28060,N_26482,N_25685);
and U28061 (N_28061,N_25735,N_26544);
or U28062 (N_28062,N_26051,N_26384);
and U28063 (N_28063,N_26052,N_25878);
and U28064 (N_28064,N_25643,N_26660);
xnor U28065 (N_28065,N_25937,N_26414);
xnor U28066 (N_28066,N_26367,N_26472);
xor U28067 (N_28067,N_26961,N_26425);
and U28068 (N_28068,N_25676,N_25582);
nor U28069 (N_28069,N_26210,N_25942);
nor U28070 (N_28070,N_25577,N_26086);
or U28071 (N_28071,N_26484,N_26258);
nand U28072 (N_28072,N_25945,N_26978);
nor U28073 (N_28073,N_25808,N_26036);
nor U28074 (N_28074,N_25999,N_25723);
and U28075 (N_28075,N_25661,N_25513);
or U28076 (N_28076,N_26882,N_26807);
or U28077 (N_28077,N_26261,N_25922);
nand U28078 (N_28078,N_26689,N_26713);
nand U28079 (N_28079,N_25891,N_26848);
and U28080 (N_28080,N_25615,N_25532);
xor U28081 (N_28081,N_26545,N_25501);
or U28082 (N_28082,N_26198,N_26573);
nor U28083 (N_28083,N_26266,N_26828);
or U28084 (N_28084,N_26453,N_26191);
and U28085 (N_28085,N_25514,N_26914);
or U28086 (N_28086,N_26872,N_25581);
xnor U28087 (N_28087,N_26635,N_25839);
nand U28088 (N_28088,N_26751,N_25858);
xnor U28089 (N_28089,N_26241,N_26135);
and U28090 (N_28090,N_25904,N_25991);
xor U28091 (N_28091,N_25865,N_26843);
nand U28092 (N_28092,N_26087,N_26540);
or U28093 (N_28093,N_26177,N_25962);
and U28094 (N_28094,N_25664,N_26193);
nor U28095 (N_28095,N_25587,N_26391);
or U28096 (N_28096,N_26916,N_26661);
xnor U28097 (N_28097,N_26492,N_26672);
nor U28098 (N_28098,N_26177,N_26758);
or U28099 (N_28099,N_26965,N_26011);
or U28100 (N_28100,N_26739,N_25977);
or U28101 (N_28101,N_25800,N_25873);
or U28102 (N_28102,N_25929,N_25860);
or U28103 (N_28103,N_26680,N_25736);
or U28104 (N_28104,N_25634,N_26221);
nand U28105 (N_28105,N_26147,N_26121);
xnor U28106 (N_28106,N_26692,N_26389);
or U28107 (N_28107,N_25517,N_26992);
xnor U28108 (N_28108,N_26750,N_26067);
nand U28109 (N_28109,N_26235,N_25915);
nor U28110 (N_28110,N_25943,N_26143);
nand U28111 (N_28111,N_25975,N_25599);
xor U28112 (N_28112,N_26312,N_26482);
or U28113 (N_28113,N_25682,N_26665);
or U28114 (N_28114,N_26463,N_26488);
xnor U28115 (N_28115,N_25557,N_26319);
nor U28116 (N_28116,N_25874,N_26546);
or U28117 (N_28117,N_26480,N_26375);
xor U28118 (N_28118,N_26994,N_25711);
or U28119 (N_28119,N_26076,N_26215);
xnor U28120 (N_28120,N_25621,N_25784);
xor U28121 (N_28121,N_26705,N_26238);
or U28122 (N_28122,N_25562,N_26102);
nor U28123 (N_28123,N_26354,N_25836);
nand U28124 (N_28124,N_25547,N_25604);
and U28125 (N_28125,N_26683,N_26297);
or U28126 (N_28126,N_26743,N_25704);
nand U28127 (N_28127,N_26886,N_26207);
nor U28128 (N_28128,N_26867,N_26502);
or U28129 (N_28129,N_26576,N_25713);
or U28130 (N_28130,N_26765,N_26986);
and U28131 (N_28131,N_25516,N_26888);
xnor U28132 (N_28132,N_26180,N_26495);
nand U28133 (N_28133,N_25629,N_25957);
nand U28134 (N_28134,N_25768,N_26848);
nand U28135 (N_28135,N_25912,N_25533);
nand U28136 (N_28136,N_26833,N_26348);
nor U28137 (N_28137,N_26799,N_25822);
or U28138 (N_28138,N_26488,N_25886);
nor U28139 (N_28139,N_25625,N_25830);
or U28140 (N_28140,N_25629,N_26942);
or U28141 (N_28141,N_26308,N_26028);
nor U28142 (N_28142,N_26449,N_26697);
nor U28143 (N_28143,N_26113,N_25791);
nor U28144 (N_28144,N_26485,N_26174);
or U28145 (N_28145,N_26142,N_25675);
or U28146 (N_28146,N_26849,N_26930);
nand U28147 (N_28147,N_26618,N_26822);
and U28148 (N_28148,N_26355,N_26337);
nand U28149 (N_28149,N_25753,N_26760);
and U28150 (N_28150,N_25594,N_26540);
or U28151 (N_28151,N_25978,N_25575);
nor U28152 (N_28152,N_25765,N_25537);
nand U28153 (N_28153,N_26071,N_26848);
nor U28154 (N_28154,N_26391,N_26066);
nand U28155 (N_28155,N_26862,N_26300);
or U28156 (N_28156,N_26995,N_25963);
or U28157 (N_28157,N_25526,N_25798);
nand U28158 (N_28158,N_25859,N_26634);
nor U28159 (N_28159,N_26176,N_26178);
xnor U28160 (N_28160,N_26560,N_25756);
nand U28161 (N_28161,N_26348,N_25510);
nor U28162 (N_28162,N_26782,N_26881);
nor U28163 (N_28163,N_25742,N_26053);
nand U28164 (N_28164,N_26324,N_26369);
or U28165 (N_28165,N_26930,N_25627);
nand U28166 (N_28166,N_26090,N_26190);
or U28167 (N_28167,N_26909,N_26610);
or U28168 (N_28168,N_26110,N_25917);
nor U28169 (N_28169,N_26811,N_26270);
nand U28170 (N_28170,N_26046,N_26972);
xnor U28171 (N_28171,N_26008,N_26029);
nor U28172 (N_28172,N_25753,N_26170);
and U28173 (N_28173,N_26331,N_25745);
or U28174 (N_28174,N_25565,N_25892);
nand U28175 (N_28175,N_25653,N_26307);
xor U28176 (N_28176,N_25922,N_26704);
and U28177 (N_28177,N_26008,N_26299);
nor U28178 (N_28178,N_26007,N_25761);
nand U28179 (N_28179,N_26341,N_26775);
nand U28180 (N_28180,N_26460,N_26446);
nor U28181 (N_28181,N_26902,N_26342);
xnor U28182 (N_28182,N_25910,N_26782);
nor U28183 (N_28183,N_26894,N_26840);
or U28184 (N_28184,N_25566,N_26533);
xor U28185 (N_28185,N_26424,N_25844);
nor U28186 (N_28186,N_25939,N_25931);
xnor U28187 (N_28187,N_26474,N_25595);
xor U28188 (N_28188,N_26972,N_25671);
nor U28189 (N_28189,N_26572,N_25806);
nand U28190 (N_28190,N_25529,N_26013);
xor U28191 (N_28191,N_26989,N_25533);
nand U28192 (N_28192,N_25851,N_26266);
nor U28193 (N_28193,N_25951,N_26921);
xor U28194 (N_28194,N_26774,N_25763);
nand U28195 (N_28195,N_26702,N_26055);
nand U28196 (N_28196,N_26709,N_25845);
or U28197 (N_28197,N_25800,N_26075);
nand U28198 (N_28198,N_25829,N_25593);
and U28199 (N_28199,N_26554,N_25677);
nor U28200 (N_28200,N_25968,N_26775);
or U28201 (N_28201,N_26258,N_26588);
and U28202 (N_28202,N_25683,N_26191);
nand U28203 (N_28203,N_26219,N_25864);
xor U28204 (N_28204,N_26574,N_26206);
nand U28205 (N_28205,N_25783,N_25925);
and U28206 (N_28206,N_26686,N_25986);
nand U28207 (N_28207,N_26086,N_26284);
or U28208 (N_28208,N_26211,N_26626);
nor U28209 (N_28209,N_26002,N_26598);
and U28210 (N_28210,N_26638,N_26389);
xor U28211 (N_28211,N_26520,N_26261);
or U28212 (N_28212,N_26783,N_26792);
nand U28213 (N_28213,N_25756,N_25693);
nand U28214 (N_28214,N_26037,N_26305);
and U28215 (N_28215,N_25577,N_26959);
nor U28216 (N_28216,N_25904,N_26068);
nand U28217 (N_28217,N_25851,N_26169);
xnor U28218 (N_28218,N_25927,N_25977);
and U28219 (N_28219,N_26982,N_26925);
nor U28220 (N_28220,N_26926,N_25842);
xnor U28221 (N_28221,N_26265,N_25748);
and U28222 (N_28222,N_26926,N_26474);
xor U28223 (N_28223,N_26156,N_26625);
nor U28224 (N_28224,N_26801,N_26016);
and U28225 (N_28225,N_26951,N_25685);
or U28226 (N_28226,N_26587,N_26793);
and U28227 (N_28227,N_26029,N_25585);
and U28228 (N_28228,N_25571,N_25909);
or U28229 (N_28229,N_26260,N_25559);
nor U28230 (N_28230,N_26082,N_26442);
nand U28231 (N_28231,N_25779,N_26557);
nor U28232 (N_28232,N_26656,N_26621);
nand U28233 (N_28233,N_25919,N_26737);
nor U28234 (N_28234,N_26162,N_26879);
or U28235 (N_28235,N_25655,N_26362);
nand U28236 (N_28236,N_25586,N_26722);
and U28237 (N_28237,N_26058,N_26540);
nor U28238 (N_28238,N_26246,N_26882);
nand U28239 (N_28239,N_25885,N_25565);
or U28240 (N_28240,N_26430,N_26969);
and U28241 (N_28241,N_26411,N_25957);
nor U28242 (N_28242,N_26864,N_26051);
and U28243 (N_28243,N_26695,N_25997);
xor U28244 (N_28244,N_26962,N_26505);
nand U28245 (N_28245,N_26710,N_25742);
nor U28246 (N_28246,N_25957,N_26823);
xor U28247 (N_28247,N_26850,N_26205);
nor U28248 (N_28248,N_26653,N_26644);
xnor U28249 (N_28249,N_26831,N_26215);
nor U28250 (N_28250,N_26370,N_26914);
xnor U28251 (N_28251,N_25979,N_26908);
and U28252 (N_28252,N_25917,N_26953);
nand U28253 (N_28253,N_26940,N_25704);
xnor U28254 (N_28254,N_26119,N_26452);
or U28255 (N_28255,N_26646,N_26307);
and U28256 (N_28256,N_26791,N_26261);
nor U28257 (N_28257,N_26118,N_25573);
xor U28258 (N_28258,N_26844,N_26033);
or U28259 (N_28259,N_25868,N_25875);
xnor U28260 (N_28260,N_25741,N_25625);
or U28261 (N_28261,N_25880,N_26983);
nor U28262 (N_28262,N_25829,N_26994);
or U28263 (N_28263,N_26317,N_26324);
or U28264 (N_28264,N_26605,N_26003);
or U28265 (N_28265,N_25857,N_25908);
or U28266 (N_28266,N_26121,N_26498);
nand U28267 (N_28267,N_26019,N_26200);
nand U28268 (N_28268,N_26792,N_25567);
nand U28269 (N_28269,N_25868,N_26608);
xor U28270 (N_28270,N_26142,N_25838);
xor U28271 (N_28271,N_26613,N_25768);
nand U28272 (N_28272,N_26262,N_26716);
xnor U28273 (N_28273,N_26879,N_26265);
nand U28274 (N_28274,N_26046,N_26269);
and U28275 (N_28275,N_26516,N_25661);
xor U28276 (N_28276,N_25507,N_26966);
and U28277 (N_28277,N_26275,N_26919);
nor U28278 (N_28278,N_26351,N_25638);
xor U28279 (N_28279,N_26278,N_26771);
nand U28280 (N_28280,N_26806,N_26521);
xor U28281 (N_28281,N_26102,N_26899);
or U28282 (N_28282,N_25542,N_26668);
and U28283 (N_28283,N_26798,N_26253);
nor U28284 (N_28284,N_26502,N_25602);
nand U28285 (N_28285,N_25677,N_25868);
and U28286 (N_28286,N_25730,N_26515);
or U28287 (N_28287,N_26442,N_26809);
nand U28288 (N_28288,N_25873,N_26955);
xor U28289 (N_28289,N_26038,N_26556);
and U28290 (N_28290,N_26582,N_25954);
and U28291 (N_28291,N_25942,N_25679);
nand U28292 (N_28292,N_25835,N_26667);
nor U28293 (N_28293,N_25748,N_26458);
xnor U28294 (N_28294,N_26081,N_26053);
nor U28295 (N_28295,N_25941,N_26529);
nand U28296 (N_28296,N_26569,N_26338);
and U28297 (N_28297,N_26406,N_26669);
nor U28298 (N_28298,N_26806,N_26450);
xnor U28299 (N_28299,N_25973,N_26695);
and U28300 (N_28300,N_26847,N_26242);
and U28301 (N_28301,N_26495,N_25740);
xnor U28302 (N_28302,N_26218,N_26988);
or U28303 (N_28303,N_26208,N_25966);
or U28304 (N_28304,N_25971,N_26322);
nor U28305 (N_28305,N_26377,N_26989);
nor U28306 (N_28306,N_25676,N_26199);
nand U28307 (N_28307,N_26875,N_26213);
or U28308 (N_28308,N_26614,N_25786);
nor U28309 (N_28309,N_26353,N_25702);
and U28310 (N_28310,N_25795,N_26306);
nand U28311 (N_28311,N_25762,N_25765);
xnor U28312 (N_28312,N_25866,N_25752);
nor U28313 (N_28313,N_26059,N_26747);
nand U28314 (N_28314,N_26343,N_26348);
nor U28315 (N_28315,N_25909,N_26434);
or U28316 (N_28316,N_25739,N_26562);
nand U28317 (N_28317,N_26517,N_26630);
xor U28318 (N_28318,N_26529,N_25699);
and U28319 (N_28319,N_26098,N_26317);
and U28320 (N_28320,N_26921,N_26613);
nand U28321 (N_28321,N_26699,N_25502);
xnor U28322 (N_28322,N_25983,N_26769);
and U28323 (N_28323,N_26039,N_26203);
nand U28324 (N_28324,N_26655,N_26381);
xor U28325 (N_28325,N_26917,N_25935);
and U28326 (N_28326,N_25622,N_25746);
xnor U28327 (N_28327,N_25744,N_25953);
nand U28328 (N_28328,N_26038,N_25867);
xnor U28329 (N_28329,N_25745,N_26112);
xnor U28330 (N_28330,N_26232,N_26507);
nand U28331 (N_28331,N_26110,N_25799);
nor U28332 (N_28332,N_26507,N_25758);
nor U28333 (N_28333,N_26834,N_25536);
nor U28334 (N_28334,N_26370,N_25732);
nand U28335 (N_28335,N_25558,N_25776);
or U28336 (N_28336,N_26552,N_26362);
nand U28337 (N_28337,N_26184,N_26867);
or U28338 (N_28338,N_26802,N_25559);
or U28339 (N_28339,N_25646,N_26001);
nand U28340 (N_28340,N_25785,N_26868);
nand U28341 (N_28341,N_25986,N_26894);
and U28342 (N_28342,N_26998,N_26171);
and U28343 (N_28343,N_26554,N_26190);
xnor U28344 (N_28344,N_26931,N_25516);
nor U28345 (N_28345,N_25628,N_26058);
xnor U28346 (N_28346,N_25983,N_25882);
and U28347 (N_28347,N_25717,N_25952);
nor U28348 (N_28348,N_26825,N_26080);
nand U28349 (N_28349,N_25745,N_25984);
nand U28350 (N_28350,N_26422,N_25755);
or U28351 (N_28351,N_25778,N_26871);
nor U28352 (N_28352,N_26299,N_26841);
and U28353 (N_28353,N_26069,N_26103);
and U28354 (N_28354,N_26368,N_25935);
xnor U28355 (N_28355,N_26285,N_26088);
and U28356 (N_28356,N_25693,N_25815);
nand U28357 (N_28357,N_25620,N_26215);
nor U28358 (N_28358,N_26468,N_25940);
or U28359 (N_28359,N_26338,N_25546);
or U28360 (N_28360,N_26992,N_26168);
or U28361 (N_28361,N_25917,N_26147);
or U28362 (N_28362,N_25660,N_26128);
xor U28363 (N_28363,N_26594,N_26288);
and U28364 (N_28364,N_26180,N_26411);
xor U28365 (N_28365,N_26566,N_26979);
nor U28366 (N_28366,N_25725,N_26335);
and U28367 (N_28367,N_25988,N_26891);
or U28368 (N_28368,N_26038,N_26931);
xor U28369 (N_28369,N_26544,N_26220);
xnor U28370 (N_28370,N_26706,N_26659);
nor U28371 (N_28371,N_26646,N_25836);
or U28372 (N_28372,N_25932,N_26401);
and U28373 (N_28373,N_26722,N_26457);
or U28374 (N_28374,N_25586,N_26913);
and U28375 (N_28375,N_26475,N_25624);
or U28376 (N_28376,N_26609,N_26021);
and U28377 (N_28377,N_26692,N_26216);
nand U28378 (N_28378,N_25906,N_25566);
and U28379 (N_28379,N_26685,N_26649);
and U28380 (N_28380,N_26250,N_25863);
or U28381 (N_28381,N_26583,N_26246);
xor U28382 (N_28382,N_26543,N_26292);
nor U28383 (N_28383,N_25860,N_25810);
nor U28384 (N_28384,N_25780,N_26729);
and U28385 (N_28385,N_25803,N_26779);
or U28386 (N_28386,N_25774,N_26333);
nor U28387 (N_28387,N_26673,N_26182);
or U28388 (N_28388,N_25671,N_26123);
nor U28389 (N_28389,N_26190,N_26255);
and U28390 (N_28390,N_26515,N_26966);
nand U28391 (N_28391,N_26835,N_26064);
or U28392 (N_28392,N_26702,N_26901);
or U28393 (N_28393,N_26360,N_25652);
or U28394 (N_28394,N_26726,N_26096);
nor U28395 (N_28395,N_26302,N_26150);
and U28396 (N_28396,N_26173,N_26489);
or U28397 (N_28397,N_26338,N_26222);
nor U28398 (N_28398,N_26375,N_26009);
and U28399 (N_28399,N_26781,N_25818);
nor U28400 (N_28400,N_26472,N_26322);
and U28401 (N_28401,N_26353,N_26883);
nor U28402 (N_28402,N_26376,N_26937);
xor U28403 (N_28403,N_25675,N_26191);
and U28404 (N_28404,N_25963,N_26060);
and U28405 (N_28405,N_26623,N_26109);
nand U28406 (N_28406,N_25901,N_26577);
nor U28407 (N_28407,N_25656,N_26542);
nand U28408 (N_28408,N_26771,N_26078);
xnor U28409 (N_28409,N_26077,N_26892);
and U28410 (N_28410,N_25703,N_25607);
nand U28411 (N_28411,N_26268,N_26756);
nand U28412 (N_28412,N_25847,N_26923);
and U28413 (N_28413,N_26950,N_26776);
or U28414 (N_28414,N_26287,N_25898);
xor U28415 (N_28415,N_26653,N_25569);
nand U28416 (N_28416,N_26399,N_26749);
and U28417 (N_28417,N_25567,N_26706);
or U28418 (N_28418,N_25912,N_26075);
or U28419 (N_28419,N_26796,N_25830);
xor U28420 (N_28420,N_26012,N_25675);
nand U28421 (N_28421,N_26856,N_26045);
or U28422 (N_28422,N_26021,N_26899);
nand U28423 (N_28423,N_25740,N_25726);
or U28424 (N_28424,N_26059,N_26975);
and U28425 (N_28425,N_26406,N_25655);
xor U28426 (N_28426,N_26573,N_26666);
nor U28427 (N_28427,N_26642,N_26452);
nor U28428 (N_28428,N_25619,N_25929);
or U28429 (N_28429,N_26850,N_26996);
nand U28430 (N_28430,N_26480,N_26255);
nand U28431 (N_28431,N_26653,N_26888);
or U28432 (N_28432,N_26914,N_25538);
nand U28433 (N_28433,N_25546,N_26489);
or U28434 (N_28434,N_26261,N_26487);
and U28435 (N_28435,N_25634,N_26539);
and U28436 (N_28436,N_26661,N_26348);
and U28437 (N_28437,N_26880,N_26793);
or U28438 (N_28438,N_26058,N_25880);
xnor U28439 (N_28439,N_26726,N_26399);
nand U28440 (N_28440,N_25505,N_26026);
xor U28441 (N_28441,N_26346,N_26511);
nand U28442 (N_28442,N_26734,N_25926);
and U28443 (N_28443,N_26838,N_26847);
and U28444 (N_28444,N_25755,N_25929);
xnor U28445 (N_28445,N_26410,N_26134);
and U28446 (N_28446,N_26379,N_26554);
and U28447 (N_28447,N_26328,N_26977);
and U28448 (N_28448,N_26028,N_26323);
nor U28449 (N_28449,N_25697,N_25869);
xor U28450 (N_28450,N_26273,N_25575);
nand U28451 (N_28451,N_26886,N_26123);
and U28452 (N_28452,N_25731,N_25684);
or U28453 (N_28453,N_25891,N_26203);
nor U28454 (N_28454,N_26655,N_26633);
xnor U28455 (N_28455,N_26992,N_26012);
and U28456 (N_28456,N_26790,N_26333);
and U28457 (N_28457,N_26685,N_26989);
nand U28458 (N_28458,N_26144,N_25973);
xnor U28459 (N_28459,N_26869,N_25821);
nand U28460 (N_28460,N_25754,N_25772);
nand U28461 (N_28461,N_26001,N_25842);
and U28462 (N_28462,N_26808,N_26910);
or U28463 (N_28463,N_26521,N_25977);
xnor U28464 (N_28464,N_25939,N_26597);
or U28465 (N_28465,N_26422,N_26196);
xnor U28466 (N_28466,N_25893,N_26775);
and U28467 (N_28467,N_26168,N_26284);
nor U28468 (N_28468,N_25943,N_26415);
nor U28469 (N_28469,N_25803,N_26655);
or U28470 (N_28470,N_26872,N_26003);
nand U28471 (N_28471,N_26295,N_26203);
nand U28472 (N_28472,N_25574,N_26880);
or U28473 (N_28473,N_26945,N_26393);
and U28474 (N_28474,N_26090,N_26386);
nor U28475 (N_28475,N_26148,N_25741);
nand U28476 (N_28476,N_26962,N_26082);
xor U28477 (N_28477,N_25569,N_26782);
and U28478 (N_28478,N_26818,N_26243);
or U28479 (N_28479,N_26958,N_25782);
nor U28480 (N_28480,N_26446,N_25672);
or U28481 (N_28481,N_25672,N_25953);
and U28482 (N_28482,N_26812,N_26113);
nand U28483 (N_28483,N_25522,N_26128);
and U28484 (N_28484,N_26800,N_26522);
or U28485 (N_28485,N_26545,N_26377);
or U28486 (N_28486,N_26025,N_26492);
nand U28487 (N_28487,N_26109,N_26698);
and U28488 (N_28488,N_26885,N_25890);
nor U28489 (N_28489,N_25527,N_25525);
xor U28490 (N_28490,N_26163,N_26147);
nand U28491 (N_28491,N_26804,N_26983);
and U28492 (N_28492,N_26097,N_26147);
nor U28493 (N_28493,N_26833,N_26330);
xor U28494 (N_28494,N_26810,N_25903);
or U28495 (N_28495,N_26981,N_25891);
and U28496 (N_28496,N_25797,N_26734);
nand U28497 (N_28497,N_25730,N_26656);
or U28498 (N_28498,N_25870,N_26197);
and U28499 (N_28499,N_26821,N_26327);
or U28500 (N_28500,N_27317,N_27304);
and U28501 (N_28501,N_27024,N_27508);
nor U28502 (N_28502,N_28394,N_27445);
and U28503 (N_28503,N_27268,N_27142);
nand U28504 (N_28504,N_27090,N_27307);
or U28505 (N_28505,N_27745,N_27099);
nand U28506 (N_28506,N_27237,N_28444);
and U28507 (N_28507,N_27935,N_27644);
nor U28508 (N_28508,N_27302,N_27920);
nand U28509 (N_28509,N_27426,N_28225);
and U28510 (N_28510,N_28038,N_27983);
xnor U28511 (N_28511,N_27507,N_27805);
nand U28512 (N_28512,N_27200,N_28323);
or U28513 (N_28513,N_28020,N_27741);
nand U28514 (N_28514,N_28180,N_27564);
xnor U28515 (N_28515,N_28239,N_27886);
nor U28516 (N_28516,N_27325,N_28227);
xnor U28517 (N_28517,N_27976,N_28399);
and U28518 (N_28518,N_28216,N_27377);
xnor U28519 (N_28519,N_27216,N_27893);
nor U28520 (N_28520,N_27381,N_27670);
xnor U28521 (N_28521,N_27846,N_27136);
nand U28522 (N_28522,N_28260,N_27500);
xnor U28523 (N_28523,N_27206,N_28390);
and U28524 (N_28524,N_28460,N_27406);
nand U28525 (N_28525,N_27750,N_28073);
or U28526 (N_28526,N_27281,N_27392);
nor U28527 (N_28527,N_27947,N_28302);
and U28528 (N_28528,N_28206,N_28379);
and U28529 (N_28529,N_27835,N_27737);
nor U28530 (N_28530,N_27581,N_28172);
and U28531 (N_28531,N_27316,N_27075);
xor U28532 (N_28532,N_27424,N_28226);
or U28533 (N_28533,N_27273,N_28035);
and U28534 (N_28534,N_27818,N_27039);
and U28535 (N_28535,N_27702,N_28032);
nand U28536 (N_28536,N_28418,N_28300);
or U28537 (N_28537,N_27554,N_27995);
or U28538 (N_28538,N_28343,N_28425);
nor U28539 (N_28539,N_28223,N_28437);
and U28540 (N_28540,N_27765,N_27472);
or U28541 (N_28541,N_28426,N_27997);
nand U28542 (N_28542,N_27116,N_28337);
nor U28543 (N_28543,N_28339,N_27952);
nor U28544 (N_28544,N_28064,N_28334);
nor U28545 (N_28545,N_28107,N_27149);
xor U28546 (N_28546,N_27402,N_27885);
nor U28547 (N_28547,N_28371,N_28449);
or U28548 (N_28548,N_28238,N_28123);
xor U28549 (N_28549,N_27459,N_28283);
xnor U28550 (N_28550,N_28276,N_27026);
and U28551 (N_28551,N_27719,N_28205);
and U28552 (N_28552,N_27964,N_27296);
nor U28553 (N_28553,N_27816,N_27861);
nand U28554 (N_28554,N_27855,N_27884);
or U28555 (N_28555,N_28374,N_27336);
or U28556 (N_28556,N_28469,N_27904);
xor U28557 (N_28557,N_28474,N_27235);
xor U28558 (N_28558,N_28433,N_28256);
nand U28559 (N_28559,N_28243,N_27486);
xnor U28560 (N_28560,N_28110,N_27608);
and U28561 (N_28561,N_28349,N_28413);
nor U28562 (N_28562,N_27594,N_27686);
nand U28563 (N_28563,N_28023,N_28146);
nor U28564 (N_28564,N_28295,N_27308);
and U28565 (N_28565,N_27263,N_28310);
nand U28566 (N_28566,N_27938,N_27673);
nand U28567 (N_28567,N_27771,N_27321);
xnor U28568 (N_28568,N_28489,N_27157);
and U28569 (N_28569,N_28196,N_27658);
nor U28570 (N_28570,N_27772,N_27433);
nand U28571 (N_28571,N_27191,N_27261);
nor U28572 (N_28572,N_27262,N_27298);
nor U28573 (N_28573,N_27159,N_27867);
and U28574 (N_28574,N_28287,N_27485);
nor U28575 (N_28575,N_28457,N_27796);
and U28576 (N_28576,N_27405,N_28076);
nor U28577 (N_28577,N_27172,N_27657);
nand U28578 (N_28578,N_27479,N_27731);
nand U28579 (N_28579,N_27397,N_27269);
or U28580 (N_28580,N_27088,N_27450);
xor U28581 (N_28581,N_27919,N_27990);
xnor U28582 (N_28582,N_27502,N_27797);
and U28583 (N_28583,N_27119,N_28497);
or U28584 (N_28584,N_28383,N_27044);
nand U28585 (N_28585,N_28048,N_27549);
and U28586 (N_28586,N_28067,N_27553);
and U28587 (N_28587,N_27637,N_27696);
nand U28588 (N_28588,N_27709,N_27066);
or U28589 (N_28589,N_27094,N_27160);
and U28590 (N_28590,N_27081,N_27877);
and U28591 (N_28591,N_27587,N_28100);
and U28592 (N_28592,N_28044,N_28347);
and U28593 (N_28593,N_27333,N_27738);
or U28594 (N_28594,N_28376,N_27453);
or U28595 (N_28595,N_27348,N_27106);
and U28596 (N_28596,N_28057,N_27084);
xor U28597 (N_28597,N_27277,N_27539);
xor U28598 (N_28598,N_27649,N_27386);
or U28599 (N_28599,N_28017,N_27889);
nor U28600 (N_28600,N_28309,N_28125);
and U28601 (N_28601,N_27064,N_28031);
xor U28602 (N_28602,N_27661,N_27188);
nand U28603 (N_28603,N_27598,N_27948);
and U28604 (N_28604,N_28273,N_28423);
or U28605 (N_28605,N_27408,N_27220);
or U28606 (N_28606,N_27838,N_27186);
and U28607 (N_28607,N_28106,N_28293);
xnor U28608 (N_28608,N_28414,N_27945);
nor U28609 (N_28609,N_28246,N_28094);
nor U28610 (N_28610,N_28463,N_27435);
nand U28611 (N_28611,N_28403,N_27175);
and U28612 (N_28612,N_27561,N_27833);
or U28613 (N_28613,N_27596,N_27312);
xnor U28614 (N_28614,N_27444,N_27028);
and U28615 (N_28615,N_27586,N_28289);
nor U28616 (N_28616,N_27461,N_27565);
nor U28617 (N_28617,N_27568,N_27937);
and U28618 (N_28618,N_27869,N_27556);
and U28619 (N_28619,N_27001,N_27437);
nor U28620 (N_28620,N_27866,N_27233);
nand U28621 (N_28621,N_27783,N_27624);
nor U28622 (N_28622,N_28422,N_27045);
or U28623 (N_28623,N_28159,N_28145);
or U28624 (N_28624,N_27591,N_27966);
or U28625 (N_28625,N_27132,N_27671);
nor U28626 (N_28626,N_27101,N_27258);
or U28627 (N_28627,N_28113,N_27848);
xor U28628 (N_28628,N_27830,N_27894);
or U28629 (N_28629,N_28454,N_27270);
nor U28630 (N_28630,N_27739,N_28191);
xor U28631 (N_28631,N_28492,N_28404);
and U28632 (N_28632,N_28452,N_27802);
nor U28633 (N_28633,N_27680,N_27713);
nand U28634 (N_28634,N_27943,N_27899);
or U28635 (N_28635,N_27449,N_28236);
xor U28636 (N_28636,N_27681,N_27463);
nand U28637 (N_28637,N_27700,N_28152);
xnor U28638 (N_28638,N_27354,N_28372);
or U28639 (N_28639,N_27842,N_27143);
and U28640 (N_28640,N_27369,N_27432);
and U28641 (N_28641,N_28292,N_27718);
and U28642 (N_28642,N_27641,N_28007);
and U28643 (N_28643,N_28075,N_28131);
and U28644 (N_28644,N_27616,N_27740);
and U28645 (N_28645,N_27197,N_28090);
and U28646 (N_28646,N_27653,N_27626);
nand U28647 (N_28647,N_27398,N_27388);
or U28648 (N_28648,N_27525,N_27240);
and U28649 (N_28649,N_27015,N_27743);
or U28650 (N_28650,N_27609,N_27895);
xor U28651 (N_28651,N_27213,N_27788);
nor U28652 (N_28652,N_28061,N_28315);
and U28653 (N_28653,N_28409,N_27120);
nand U28654 (N_28654,N_27870,N_28137);
and U28655 (N_28655,N_27394,N_28201);
nand U28656 (N_28656,N_27313,N_28173);
xnor U28657 (N_28657,N_28440,N_27823);
or U28658 (N_28658,N_28010,N_28391);
and U28659 (N_28659,N_28088,N_28290);
and U28660 (N_28660,N_28118,N_27786);
nor U28661 (N_28661,N_27847,N_27138);
or U28662 (N_28662,N_27462,N_27859);
or U28663 (N_28663,N_27036,N_28465);
nand U28664 (N_28664,N_27271,N_27151);
and U28665 (N_28665,N_27009,N_28208);
nand U28666 (N_28666,N_28326,N_28428);
or U28667 (N_28667,N_27247,N_28228);
or U28668 (N_28668,N_27560,N_27399);
nand U28669 (N_28669,N_28015,N_28411);
and U28670 (N_28670,N_28164,N_28194);
and U28671 (N_28671,N_27016,N_28156);
and U28672 (N_28672,N_27621,N_28401);
xor U28673 (N_28673,N_27495,N_27425);
nand U28674 (N_28674,N_27559,N_27601);
xor U28675 (N_28675,N_28219,N_27589);
nor U28676 (N_28676,N_28144,N_28186);
nand U28677 (N_28677,N_28298,N_28265);
xnor U28678 (N_28678,N_27496,N_28108);
or U28679 (N_28679,N_27518,N_28467);
and U28680 (N_28680,N_28338,N_27791);
and U28681 (N_28681,N_27804,N_28001);
nor U28682 (N_28682,N_28456,N_28091);
or U28683 (N_28683,N_27536,N_28365);
and U28684 (N_28684,N_27575,N_27178);
nor U28685 (N_28685,N_27625,N_27506);
nor U28686 (N_28686,N_27253,N_28360);
or U28687 (N_28687,N_27732,N_27431);
nor U28688 (N_28688,N_27865,N_27639);
and U28689 (N_28689,N_28491,N_28033);
xnor U28690 (N_28690,N_28024,N_27335);
nand U28691 (N_28691,N_27972,N_27027);
xor U28692 (N_28692,N_27953,N_27675);
nand U28693 (N_28693,N_28478,N_28011);
or U28694 (N_28694,N_27647,N_27611);
nor U28695 (N_28695,N_27887,N_28170);
xor U28696 (N_28696,N_27930,N_27668);
and U28697 (N_28697,N_27366,N_27008);
nor U28698 (N_28698,N_28441,N_27949);
xor U28699 (N_28699,N_27828,N_27470);
or U28700 (N_28700,N_28451,N_27141);
nand U28701 (N_28701,N_27295,N_27655);
nand U28702 (N_28702,N_27280,N_27734);
and U28703 (N_28703,N_27544,N_27767);
or U28704 (N_28704,N_28342,N_28357);
or U28705 (N_28705,N_27056,N_27717);
nand U28706 (N_28706,N_27513,N_28427);
or U28707 (N_28707,N_27613,N_27134);
nand U28708 (N_28708,N_27965,N_27455);
or U28709 (N_28709,N_28249,N_28112);
nand U28710 (N_28710,N_28060,N_27465);
nand U28711 (N_28711,N_27257,N_27697);
nor U28712 (N_28712,N_27708,N_27950);
nand U28713 (N_28713,N_27288,N_27819);
nor U28714 (N_28714,N_28340,N_28255);
nand U28715 (N_28715,N_27722,N_27092);
xnor U28716 (N_28716,N_27474,N_27249);
xor U28717 (N_28717,N_27002,N_27493);
or U28718 (N_28718,N_28192,N_28368);
nand U28719 (N_28719,N_27762,N_27127);
nand U28720 (N_28720,N_27057,N_27692);
xor U28721 (N_28721,N_27769,N_27211);
nand U28722 (N_28722,N_27020,N_27751);
and U28723 (N_28723,N_27688,N_27416);
or U28724 (N_28724,N_27382,N_27108);
xor U28725 (N_28725,N_27290,N_27289);
and U28726 (N_28726,N_27117,N_28079);
and U28727 (N_28727,N_27652,N_27597);
nor U28728 (N_28728,N_28188,N_27748);
nor U28729 (N_28729,N_27808,N_27391);
and U28730 (N_28730,N_27622,N_27969);
xor U28731 (N_28731,N_27892,N_27933);
xnor U28732 (N_28732,N_27636,N_27375);
nor U28733 (N_28733,N_27523,N_27994);
and U28734 (N_28734,N_27633,N_28153);
and U28735 (N_28735,N_27883,N_28138);
and U28736 (N_28736,N_27404,N_27152);
nand U28737 (N_28737,N_27729,N_27401);
nor U28738 (N_28738,N_27684,N_28495);
nand U28739 (N_28739,N_27961,N_27936);
nand U28740 (N_28740,N_28448,N_27774);
or U28741 (N_28741,N_27097,N_27993);
xnor U28742 (N_28742,N_27098,N_28461);
xor U28743 (N_28743,N_27590,N_27464);
nor U28744 (N_28744,N_27873,N_28183);
or U28745 (N_28745,N_27096,N_27519);
nor U28746 (N_28746,N_27103,N_28353);
xnor U28747 (N_28747,N_27113,N_27931);
and U28748 (N_28748,N_27730,N_27407);
or U28749 (N_28749,N_27475,N_27501);
and U28750 (N_28750,N_28417,N_27856);
nor U28751 (N_28751,N_27156,N_27198);
or U28752 (N_28752,N_27635,N_27775);
nand U28753 (N_28753,N_27987,N_27543);
nand U28754 (N_28754,N_28050,N_28373);
xnor U28755 (N_28755,N_28042,N_28080);
and U28756 (N_28756,N_27839,N_27293);
xor U28757 (N_28757,N_28412,N_28447);
or U28758 (N_28758,N_27139,N_27114);
and U28759 (N_28759,N_28286,N_27801);
or U28760 (N_28760,N_27980,N_27538);
or U28761 (N_28761,N_27022,N_28065);
and U28762 (N_28762,N_27572,N_27292);
nand U28763 (N_28763,N_28299,N_28092);
xor U28764 (N_28764,N_28204,N_27758);
nor U28765 (N_28765,N_27082,N_27358);
nand U28766 (N_28766,N_27588,N_27913);
or U28767 (N_28767,N_27996,N_27306);
xnor U28768 (N_28768,N_27612,N_27355);
xnor U28769 (N_28769,N_27315,N_27309);
or U28770 (N_28770,N_28455,N_28154);
nor U28771 (N_28771,N_28139,N_28301);
or U28772 (N_28772,N_28132,N_27787);
and U28773 (N_28773,N_27215,N_27778);
or U28774 (N_28774,N_27569,N_27605);
or U28775 (N_28775,N_28259,N_27939);
xnor U28776 (N_28776,N_27107,N_27442);
xor U28777 (N_28777,N_27524,N_28251);
and U28778 (N_28778,N_28013,N_27574);
or U28779 (N_28779,N_28378,N_27115);
nand U28780 (N_28780,N_28285,N_27194);
xor U28781 (N_28781,N_28415,N_27222);
xnor U28782 (N_28782,N_28335,N_27104);
nor U28783 (N_28783,N_27050,N_27468);
xor U28784 (N_28784,N_27580,N_27048);
and U28785 (N_28785,N_28278,N_28096);
nor U28786 (N_28786,N_27441,N_28271);
and U28787 (N_28787,N_27343,N_28482);
or U28788 (N_28788,N_28332,N_27322);
xor U28789 (N_28789,N_27164,N_27725);
nor U28790 (N_28790,N_28052,N_28071);
or U28791 (N_28791,N_28479,N_28483);
xnor U28792 (N_28792,N_27779,N_27212);
or U28793 (N_28793,N_27168,N_27109);
xnor U28794 (N_28794,N_28000,N_27390);
xor U28795 (N_28795,N_27422,N_28199);
nor U28796 (N_28796,N_28250,N_28135);
nand U28797 (N_28797,N_28361,N_27959);
or U28798 (N_28798,N_27339,N_27192);
or U28799 (N_28799,N_27723,N_28158);
nor U28800 (N_28800,N_27267,N_27534);
nand U28801 (N_28801,N_27360,N_27807);
xnor U28802 (N_28802,N_28389,N_28136);
nor U28803 (N_28803,N_27578,N_27225);
and U28804 (N_28804,N_28410,N_28179);
nand U28805 (N_28805,N_28329,N_28367);
nand U28806 (N_28806,N_28066,N_28439);
and U28807 (N_28807,N_27032,N_28036);
and U28808 (N_28808,N_28258,N_27509);
or U28809 (N_28809,N_27478,N_27439);
nor U28810 (N_28810,N_28117,N_28025);
and U28811 (N_28811,N_27144,N_28224);
or U28812 (N_28812,N_27085,N_28321);
and U28813 (N_28813,N_27476,N_27025);
or U28814 (N_28814,N_27438,N_27126);
nand U28815 (N_28815,N_28009,N_28473);
nor U28816 (N_28816,N_28161,N_27409);
nand U28817 (N_28817,N_28476,N_27691);
nand U28818 (N_28818,N_27654,N_27914);
nand U28819 (N_28819,N_27790,N_27196);
and U28820 (N_28820,N_27060,N_27971);
nor U28821 (N_28821,N_28237,N_28459);
xor U28822 (N_28822,N_27412,N_27185);
nand U28823 (N_28823,N_27849,N_28450);
xnor U28824 (N_28824,N_28234,N_27037);
nor U28825 (N_28825,N_27676,N_27434);
nor U28826 (N_28826,N_28486,N_27916);
nor U28827 (N_28827,N_27121,N_27874);
and U28828 (N_28828,N_27323,N_27137);
xnor U28829 (N_28829,N_27182,N_28129);
xor U28830 (N_28830,N_28244,N_27687);
xnor U28831 (N_28831,N_28037,N_27630);
nor U28832 (N_28832,N_27881,N_27733);
or U28833 (N_28833,N_27146,N_27667);
xnor U28834 (N_28834,N_27130,N_27456);
and U28835 (N_28835,N_28466,N_28307);
nor U28836 (N_28836,N_28253,N_27190);
nor U28837 (N_28837,N_27248,N_27551);
nand U28838 (N_28838,N_27367,N_28174);
and U28839 (N_28839,N_27042,N_28214);
and U28840 (N_28840,N_27571,N_27773);
or U28841 (N_28841,N_27863,N_27794);
nor U28842 (N_28842,N_27150,N_28014);
or U28843 (N_28843,N_28317,N_27579);
nand U28844 (N_28844,N_27034,N_27970);
and U28845 (N_28845,N_27857,N_28430);
and U28846 (N_28846,N_28281,N_28041);
or U28847 (N_28847,N_27582,N_27825);
nand U28848 (N_28848,N_27875,N_27954);
nor U28849 (N_28849,N_28093,N_28324);
and U28850 (N_28850,N_27843,N_28443);
or U28851 (N_28851,N_27690,N_27577);
nor U28852 (N_28852,N_27204,N_27195);
xnor U28853 (N_28853,N_28045,N_27299);
xnor U28854 (N_28854,N_28406,N_27926);
nor U28855 (N_28855,N_28083,N_27068);
or U28856 (N_28856,N_27753,N_27078);
nor U28857 (N_28857,N_28493,N_27837);
xnor U28858 (N_28858,N_28026,N_28097);
xnor U28859 (N_28859,N_27557,N_27202);
nor U28860 (N_28860,N_27076,N_27728);
xnor U28861 (N_28861,N_27166,N_28318);
nand U28862 (N_28862,N_27759,N_27207);
nand U28863 (N_28863,N_27891,N_27595);
nand U28864 (N_28864,N_27457,N_27614);
and U28865 (N_28865,N_27129,N_27246);
or U28866 (N_28866,N_28082,N_27357);
nand U28867 (N_28867,N_27642,N_28058);
xnor U28868 (N_28868,N_27736,N_28470);
or U28869 (N_28869,N_28217,N_27054);
or U28870 (N_28870,N_28344,N_27419);
and U28871 (N_28871,N_27189,N_27944);
nand U28872 (N_28872,N_28182,N_27545);
nor U28873 (N_28873,N_27698,N_27041);
or U28874 (N_28874,N_28322,N_28345);
nor U28875 (N_28875,N_27365,N_28356);
and U28876 (N_28876,N_27985,N_28220);
or U28877 (N_28877,N_27634,N_27726);
and U28878 (N_28878,N_27010,N_27297);
nand U28879 (N_28879,N_28316,N_27558);
nor U28880 (N_28880,N_28016,N_27324);
xor U28881 (N_28881,N_27678,N_27451);
xor U28882 (N_28882,N_28130,N_27570);
nand U28883 (N_28883,N_27283,N_27845);
nor U28884 (N_28884,N_27087,N_28084);
or U28885 (N_28885,N_28438,N_28006);
nor U28886 (N_28886,N_27537,N_27260);
nor U28887 (N_28887,N_27040,N_28421);
xor U28888 (N_28888,N_27006,N_27327);
xnor U28889 (N_28889,N_27757,N_27917);
or U28890 (N_28890,N_27706,N_27467);
nor U28891 (N_28891,N_27962,N_28304);
nand U28892 (N_28892,N_27862,N_27907);
nor U28893 (N_28893,N_27984,N_27466);
nand U28894 (N_28894,N_27173,N_27694);
nor U28895 (N_28895,N_28364,N_28103);
and U28896 (N_28896,N_27573,N_28176);
xnor U28897 (N_28897,N_27529,N_27111);
xor U28898 (N_28898,N_28375,N_27413);
or U28899 (N_28899,N_28116,N_27666);
or U28900 (N_28900,N_27811,N_28054);
nor U28901 (N_28901,N_28069,N_27303);
or U28902 (N_28902,N_28102,N_27527);
nor U28903 (N_28903,N_27430,N_28148);
nor U28904 (N_28904,N_28056,N_27209);
nor U28905 (N_28905,N_27023,N_28140);
or U28906 (N_28906,N_28346,N_27515);
or U28907 (N_28907,N_28397,N_27429);
nor U28908 (N_28908,N_28126,N_27603);
and U28909 (N_28909,N_27361,N_27902);
or U28910 (N_28910,N_28046,N_27817);
nand U28911 (N_28911,N_27683,N_27448);
nand U28912 (N_28912,N_28330,N_27311);
nand U28913 (N_28913,N_27440,N_27380);
nor U28914 (N_28914,N_27223,N_27359);
nand U28915 (N_28915,N_27344,N_27682);
and U28916 (N_28916,N_27427,N_27208);
xnor U28917 (N_28917,N_27793,N_27494);
nor U28918 (N_28918,N_27770,N_28215);
and U28919 (N_28919,N_27827,N_28222);
nand U28920 (N_28920,N_27338,N_27925);
and U28921 (N_28921,N_28232,N_27091);
and U28922 (N_28922,N_28157,N_28178);
or U28923 (N_28923,N_27393,N_27876);
or U28924 (N_28924,N_28351,N_27033);
nand U28925 (N_28925,N_27319,N_27704);
and U28926 (N_28926,N_27318,N_27803);
or U28927 (N_28927,N_27287,N_28008);
nand U28928 (N_28928,N_28218,N_27177);
xnor U28929 (N_28929,N_27231,N_27238);
or U28930 (N_28930,N_28162,N_27656);
nand U28931 (N_28931,N_27989,N_28143);
xor U28932 (N_28932,N_27662,N_27148);
and U28933 (N_28933,N_28099,N_28085);
xor U28934 (N_28934,N_27498,N_28257);
nand U28935 (N_28935,N_27715,N_27403);
xor U28936 (N_28936,N_27284,N_27294);
or U28937 (N_28937,N_27535,N_28072);
or U28938 (N_28938,N_27062,N_27777);
nor U28939 (N_28939,N_27880,N_27242);
and U28940 (N_28940,N_27526,N_27968);
nor U28941 (N_28941,N_27005,N_27232);
nor U28942 (N_28942,N_28121,N_27888);
xor U28943 (N_28943,N_28328,N_27973);
or U28944 (N_28944,N_28193,N_27712);
xnor U28945 (N_28945,N_27255,N_28169);
nor U28946 (N_28946,N_27105,N_28419);
nand U28947 (N_28947,N_28384,N_28086);
and U28948 (N_28948,N_27620,N_27615);
or U28949 (N_28949,N_28034,N_27305);
nand U28950 (N_28950,N_28348,N_27999);
and U28951 (N_28951,N_27915,N_27245);
xnor U28952 (N_28952,N_27070,N_27711);
nor U28953 (N_28953,N_27266,N_27370);
xnor U28954 (N_28954,N_27593,N_27224);
nand U28955 (N_28955,N_27176,N_27004);
nor U28956 (N_28956,N_27850,N_27013);
and U28957 (N_28957,N_27555,N_27163);
and U28958 (N_28958,N_28053,N_27443);
and U28959 (N_28959,N_27533,N_27960);
nor U28960 (N_28960,N_27286,N_28078);
nor U28961 (N_28961,N_28280,N_27038);
or U28962 (N_28962,N_28279,N_28398);
nor U28963 (N_28963,N_28210,N_28475);
nand U28964 (N_28964,N_28101,N_28494);
and U28965 (N_28965,N_27840,N_27051);
nor U28966 (N_28966,N_27912,N_28231);
and U28967 (N_28967,N_28319,N_27083);
nand U28968 (N_28968,N_28387,N_27187);
and U28969 (N_28969,N_27351,N_28233);
or U28970 (N_28970,N_27617,N_27900);
and U28971 (N_28971,N_27184,N_27860);
and U28972 (N_28972,N_28336,N_28021);
nor U28973 (N_28973,N_27063,N_27218);
nor U28974 (N_28974,N_27784,N_28262);
and U28975 (N_28975,N_27362,N_27274);
nor U28976 (N_28976,N_27145,N_27607);
or U28977 (N_28977,N_27781,N_27170);
and U28978 (N_28978,N_27679,N_28471);
nor U28979 (N_28979,N_28354,N_27073);
nor U28980 (N_28980,N_27724,N_28277);
xnor U28981 (N_28981,N_28370,N_27963);
or U28982 (N_28982,N_28120,N_28163);
and U28983 (N_28983,N_28077,N_27659);
nor U28984 (N_28984,N_27147,N_27714);
xor U28985 (N_28985,N_27396,N_27623);
nor U28986 (N_28986,N_27065,N_28040);
nand U28987 (N_28987,N_28039,N_27368);
nand U28988 (N_28988,N_28355,N_28264);
nor U28989 (N_28989,N_28458,N_27584);
or U28990 (N_28990,N_27505,N_27499);
nor U28991 (N_28991,N_27940,N_28481);
nor U28992 (N_28992,N_27924,N_27489);
xor U28993 (N_28993,N_27019,N_28030);
or U28994 (N_28994,N_27632,N_28119);
and U28995 (N_28995,N_27086,N_27095);
xor U28996 (N_28996,N_27744,N_28377);
nand U28997 (N_28997,N_27125,N_28147);
xnor U28998 (N_28998,N_28175,N_27118);
nand U28999 (N_28999,N_27764,N_27516);
and U29000 (N_29000,N_27974,N_28095);
xor U29001 (N_29001,N_28181,N_28122);
xnor U29002 (N_29002,N_28267,N_27436);
nand U29003 (N_29003,N_28029,N_27254);
nor U29004 (N_29004,N_28104,N_27243);
or U29005 (N_29005,N_27872,N_27167);
and U29006 (N_29006,N_27908,N_27956);
nor U29007 (N_29007,N_28424,N_27812);
xor U29008 (N_29008,N_28151,N_27530);
and U29009 (N_29009,N_27473,N_27279);
and U29010 (N_29010,N_27922,N_27768);
or U29011 (N_29011,N_27821,N_28089);
nor U29012 (N_29012,N_27007,N_27932);
or U29013 (N_29013,N_27606,N_28221);
xnor U29014 (N_29014,N_28059,N_27490);
xnor U29015 (N_29015,N_27992,N_27824);
nor U29016 (N_29016,N_27341,N_27552);
nor U29017 (N_29017,N_27858,N_27660);
or U29018 (N_29018,N_27665,N_27663);
nand U29019 (N_29019,N_27183,N_27514);
nor U29020 (N_29020,N_27820,N_27058);
and U29021 (N_29021,N_27052,N_27331);
or U29022 (N_29022,N_27721,N_28213);
nor U29023 (N_29023,N_27131,N_27929);
xnor U29024 (N_29024,N_28429,N_27909);
nor U29025 (N_29025,N_27522,N_28247);
nand U29026 (N_29026,N_27646,N_28420);
nand U29027 (N_29027,N_27521,N_27227);
or U29028 (N_29028,N_28312,N_27799);
or U29029 (N_29029,N_27766,N_27735);
or U29030 (N_29030,N_28477,N_28165);
or U29031 (N_29031,N_27049,N_27205);
nand U29032 (N_29032,N_27193,N_28134);
nand U29033 (N_29033,N_28268,N_27967);
nand U29034 (N_29034,N_28266,N_28068);
nor U29035 (N_29035,N_27447,N_27179);
and U29036 (N_29036,N_27898,N_28124);
or U29037 (N_29037,N_27854,N_28184);
and U29038 (N_29038,N_27077,N_28115);
or U29039 (N_29039,N_27174,N_27648);
nor U29040 (N_29040,N_28386,N_27776);
nand U29041 (N_29041,N_27806,N_28109);
or U29042 (N_29042,N_28229,N_27003);
xor U29043 (N_29043,N_27251,N_27927);
nor U29044 (N_29044,N_27428,N_28245);
xor U29045 (N_29045,N_27853,N_27763);
or U29046 (N_29046,N_27328,N_27955);
nor U29047 (N_29047,N_27746,N_28488);
xor U29048 (N_29048,N_28185,N_28171);
nor U29049 (N_29049,N_28294,N_28002);
nor U29050 (N_29050,N_27664,N_27510);
and U29051 (N_29051,N_28149,N_27813);
and U29052 (N_29052,N_28369,N_28027);
or U29053 (N_29053,N_27975,N_28446);
or U29054 (N_29054,N_27878,N_27385);
or U29055 (N_29055,N_27497,N_27046);
and U29056 (N_29056,N_27345,N_28070);
xor U29057 (N_29057,N_28333,N_27000);
and U29058 (N_29058,N_27979,N_27342);
or U29059 (N_29059,N_28313,N_27901);
nand U29060 (N_29060,N_28388,N_28019);
or U29061 (N_29061,N_28269,N_27282);
and U29062 (N_29062,N_28062,N_28200);
and U29063 (N_29063,N_27030,N_27102);
nor U29064 (N_29064,N_28189,N_28142);
or U29065 (N_29065,N_27320,N_27483);
nor U29066 (N_29066,N_28407,N_27689);
and U29067 (N_29067,N_27374,N_28308);
or U29068 (N_29068,N_27563,N_27517);
nand U29069 (N_29069,N_27710,N_27203);
or U29070 (N_29070,N_28445,N_27600);
nor U29071 (N_29071,N_28453,N_28240);
nor U29072 (N_29072,N_27701,N_28063);
nand U29073 (N_29073,N_28203,N_27452);
nor U29074 (N_29074,N_27080,N_27171);
nor U29075 (N_29075,N_27420,N_27110);
or U29076 (N_29076,N_28381,N_27981);
nand U29077 (N_29077,N_28435,N_27411);
or U29078 (N_29078,N_27252,N_27800);
xnor U29079 (N_29079,N_28498,N_27014);
xnor U29080 (N_29080,N_27592,N_27998);
xor U29081 (N_29081,N_27511,N_27844);
xnor U29082 (N_29082,N_27562,N_27165);
xor U29083 (N_29083,N_27782,N_27350);
nor U29084 (N_29084,N_27669,N_28400);
nor U29085 (N_29085,N_28395,N_28382);
or U29086 (N_29086,N_28022,N_27749);
nand U29087 (N_29087,N_27378,N_27481);
xnor U29088 (N_29088,N_27155,N_27460);
xor U29089 (N_29089,N_27789,N_28402);
and U29090 (N_29090,N_27123,N_27384);
nand U29091 (N_29091,N_28150,N_27072);
nand U29092 (N_29092,N_28288,N_28254);
nand U29093 (N_29093,N_27228,N_27415);
nand U29094 (N_29094,N_27055,N_27079);
xnor U29095 (N_29095,N_27941,N_27067);
nor U29096 (N_29096,N_27035,N_27583);
or U29097 (N_29097,N_27239,N_28464);
nor U29098 (N_29098,N_27346,N_28074);
or U29099 (N_29099,N_27256,N_28270);
nor U29100 (N_29100,N_27071,N_27410);
or U29101 (N_29101,N_27018,N_28392);
and U29102 (N_29102,N_28408,N_27285);
or U29103 (N_29103,N_27214,N_28472);
xor U29104 (N_29104,N_27011,N_27868);
or U29105 (N_29105,N_27334,N_28496);
and U29106 (N_29106,N_27471,N_27373);
or U29107 (N_29107,N_27353,N_27792);
nor U29108 (N_29108,N_28081,N_27069);
xor U29109 (N_29109,N_28314,N_27903);
xor U29110 (N_29110,N_28385,N_27531);
or U29111 (N_29111,N_27133,N_28190);
nor U29112 (N_29112,N_27761,N_27798);
xnor U29113 (N_29113,N_27376,N_27484);
nand U29114 (N_29114,N_28127,N_27836);
nand U29115 (N_29115,N_27332,N_28468);
nand U29116 (N_29116,N_28480,N_27550);
and U29117 (N_29117,N_27153,N_27259);
or U29118 (N_29118,N_27504,N_27905);
nor U29119 (N_29119,N_27918,N_28003);
and U29120 (N_29120,N_27414,N_27275);
or U29121 (N_29121,N_27879,N_27928);
nor U29122 (N_29122,N_27566,N_28209);
nor U29123 (N_29123,N_27389,N_27988);
or U29124 (N_29124,N_28242,N_27951);
or U29125 (N_29125,N_27301,N_28111);
nand U29126 (N_29126,N_27112,N_27815);
nand U29127 (N_29127,N_27264,N_27423);
nor U29128 (N_29128,N_27851,N_27640);
xnor U29129 (N_29129,N_27512,N_28352);
nand U29130 (N_29130,N_27244,N_28168);
xnor U29131 (N_29131,N_27180,N_27978);
nand U29132 (N_29132,N_27832,N_27528);
xor U29133 (N_29133,N_28284,N_27541);
and U29134 (N_29134,N_27982,N_27400);
nor U29135 (N_29135,N_28275,N_27379);
and U29136 (N_29136,N_27674,N_28128);
xnor U29137 (N_29137,N_28049,N_27540);
nand U29138 (N_29138,N_28098,N_27610);
or U29139 (N_29139,N_27795,N_28490);
nor U29140 (N_29140,N_28320,N_27747);
and U29141 (N_29141,N_27074,N_27387);
nor U29142 (N_29142,N_28341,N_28272);
xnor U29143 (N_29143,N_27576,N_28087);
and U29144 (N_29144,N_27326,N_27542);
and U29145 (N_29145,N_27651,N_28485);
nand U29146 (N_29146,N_27754,N_27469);
xnor U29147 (N_29147,N_28166,N_27124);
nor U29148 (N_29148,N_28442,N_28012);
nor U29149 (N_29149,N_27602,N_27241);
nand U29150 (N_29150,N_28028,N_27631);
nand U29151 (N_29151,N_27643,N_27629);
or U29152 (N_29152,N_27314,N_27991);
and U29153 (N_29153,N_27089,N_28261);
nand U29154 (N_29154,N_27477,N_27672);
xnor U29155 (N_29155,N_27520,N_27645);
and U29156 (N_29156,N_27201,N_28396);
nor U29157 (N_29157,N_27012,N_27546);
or U29158 (N_29158,N_27356,N_28291);
or U29159 (N_29159,N_28114,N_27871);
nand U29160 (N_29160,N_28462,N_28197);
xor U29161 (N_29161,N_27337,N_28362);
and U29162 (N_29162,N_27363,N_27488);
nand U29163 (N_29163,N_27760,N_27921);
nor U29164 (N_29164,N_27219,N_27547);
xor U29165 (N_29165,N_27229,N_27061);
nor U29166 (N_29166,N_28297,N_27716);
xnor U29167 (N_29167,N_28331,N_28207);
or U29168 (N_29168,N_27210,N_28047);
nor U29169 (N_29169,N_28311,N_27421);
nor U29170 (N_29170,N_27154,N_28198);
or U29171 (N_29171,N_27896,N_27140);
nand U29172 (N_29172,N_27480,N_28434);
nor U29173 (N_29173,N_28187,N_27977);
or U29174 (N_29174,N_28306,N_27650);
nor U29175 (N_29175,N_27230,N_27910);
and U29176 (N_29176,N_27169,N_27882);
nor U29177 (N_29177,N_27628,N_28230);
nand U29178 (N_29178,N_28350,N_27785);
or U29179 (N_29179,N_28252,N_27372);
and U29180 (N_29180,N_27059,N_28358);
xor U29181 (N_29181,N_27503,N_27250);
xnor U29182 (N_29182,N_27705,N_27329);
nor U29183 (N_29183,N_27162,N_27829);
nand U29184 (N_29184,N_27826,N_27492);
or U29185 (N_29185,N_28055,N_27199);
and U29186 (N_29186,N_27300,N_28380);
nor U29187 (N_29187,N_27364,N_27707);
or U29188 (N_29188,N_27278,N_27236);
xnor U29189 (N_29189,N_27567,N_28018);
or U29190 (N_29190,N_28363,N_27418);
or U29191 (N_29191,N_27371,N_27599);
nand U29192 (N_29192,N_27482,N_28105);
or U29193 (N_29193,N_27685,N_27619);
or U29194 (N_29194,N_27695,N_27677);
xor U29195 (N_29195,N_27890,N_27135);
xor U29196 (N_29196,N_27946,N_27417);
xor U29197 (N_29197,N_28043,N_28416);
nor U29198 (N_29198,N_28051,N_27053);
or U29199 (N_29199,N_27330,N_28499);
nor U29200 (N_29200,N_27349,N_27310);
nand U29201 (N_29201,N_27161,N_27395);
and U29202 (N_29202,N_27755,N_28274);
xnor U29203 (N_29203,N_27958,N_28202);
nor U29204 (N_29204,N_27029,N_27834);
nor U29205 (N_29205,N_27809,N_27221);
and U29206 (N_29206,N_28155,N_27934);
nand U29207 (N_29207,N_27780,N_27923);
xor U29208 (N_29208,N_28235,N_27727);
or U29209 (N_29209,N_28005,N_27548);
and U29210 (N_29210,N_28432,N_28160);
and U29211 (N_29211,N_27841,N_27276);
or U29212 (N_29212,N_27226,N_27458);
or U29213 (N_29213,N_27383,N_28405);
nor U29214 (N_29214,N_28133,N_28484);
nand U29215 (N_29215,N_28327,N_27852);
and U29216 (N_29216,N_27752,N_28393);
xor U29217 (N_29217,N_27699,N_27720);
nor U29218 (N_29218,N_28296,N_27814);
xnor U29219 (N_29219,N_28431,N_28167);
and U29220 (N_29220,N_27234,N_28177);
and U29221 (N_29221,N_27864,N_28359);
nand U29222 (N_29222,N_27291,N_27265);
nand U29223 (N_29223,N_27942,N_27822);
nor U29224 (N_29224,N_27446,N_27272);
and U29225 (N_29225,N_27017,N_27831);
or U29226 (N_29226,N_27986,N_28211);
nor U29227 (N_29227,N_27618,N_27122);
xnor U29228 (N_29228,N_27100,N_27487);
or U29229 (N_29229,N_27756,N_28263);
nand U29230 (N_29230,N_27911,N_27347);
xor U29231 (N_29231,N_27693,N_27957);
xor U29232 (N_29232,N_27491,N_27158);
and U29233 (N_29233,N_27742,N_27454);
nor U29234 (N_29234,N_27352,N_28305);
xnor U29235 (N_29235,N_27021,N_28248);
or U29236 (N_29236,N_27031,N_27897);
xor U29237 (N_29237,N_28282,N_28325);
nand U29238 (N_29238,N_27047,N_28436);
or U29239 (N_29239,N_28195,N_28004);
or U29240 (N_29240,N_28303,N_27043);
nand U29241 (N_29241,N_27604,N_28487);
xor U29242 (N_29242,N_28241,N_27217);
or U29243 (N_29243,N_27181,N_27638);
or U29244 (N_29244,N_27532,N_27585);
nand U29245 (N_29245,N_27093,N_27627);
nor U29246 (N_29246,N_28141,N_27810);
nor U29247 (N_29247,N_28212,N_27906);
xnor U29248 (N_29248,N_27128,N_27340);
nand U29249 (N_29249,N_28366,N_27703);
nor U29250 (N_29250,N_27834,N_27628);
and U29251 (N_29251,N_28454,N_28390);
and U29252 (N_29252,N_27025,N_27521);
nand U29253 (N_29253,N_27266,N_27601);
nand U29254 (N_29254,N_28152,N_28219);
and U29255 (N_29255,N_27275,N_28267);
and U29256 (N_29256,N_27597,N_27540);
nand U29257 (N_29257,N_28286,N_28241);
nor U29258 (N_29258,N_28316,N_27442);
and U29259 (N_29259,N_27373,N_28016);
nor U29260 (N_29260,N_27498,N_27792);
and U29261 (N_29261,N_27011,N_27467);
or U29262 (N_29262,N_27236,N_27268);
nor U29263 (N_29263,N_27994,N_27915);
or U29264 (N_29264,N_27088,N_27145);
nand U29265 (N_29265,N_27105,N_28107);
or U29266 (N_29266,N_27192,N_27101);
nor U29267 (N_29267,N_27110,N_27688);
nor U29268 (N_29268,N_28061,N_27349);
and U29269 (N_29269,N_27892,N_28225);
xor U29270 (N_29270,N_28456,N_27978);
or U29271 (N_29271,N_27083,N_27782);
and U29272 (N_29272,N_27471,N_27730);
or U29273 (N_29273,N_28232,N_27365);
xnor U29274 (N_29274,N_27617,N_27168);
or U29275 (N_29275,N_27801,N_27110);
nor U29276 (N_29276,N_28318,N_27662);
nand U29277 (N_29277,N_27273,N_28400);
nor U29278 (N_29278,N_28025,N_27460);
nor U29279 (N_29279,N_27657,N_28191);
xor U29280 (N_29280,N_27491,N_27389);
and U29281 (N_29281,N_28141,N_27493);
and U29282 (N_29282,N_28155,N_27700);
or U29283 (N_29283,N_27497,N_27131);
xor U29284 (N_29284,N_27999,N_28378);
or U29285 (N_29285,N_28084,N_28376);
and U29286 (N_29286,N_28197,N_27582);
or U29287 (N_29287,N_27955,N_27952);
nand U29288 (N_29288,N_27694,N_27780);
and U29289 (N_29289,N_27591,N_27655);
nand U29290 (N_29290,N_27691,N_27696);
nand U29291 (N_29291,N_27142,N_28208);
xnor U29292 (N_29292,N_28041,N_28095);
xor U29293 (N_29293,N_28282,N_27648);
xnor U29294 (N_29294,N_28120,N_27060);
nor U29295 (N_29295,N_28253,N_27109);
or U29296 (N_29296,N_27146,N_27459);
xnor U29297 (N_29297,N_27150,N_27872);
nor U29298 (N_29298,N_27407,N_28001);
and U29299 (N_29299,N_28226,N_27694);
or U29300 (N_29300,N_27117,N_28291);
and U29301 (N_29301,N_28045,N_28426);
nand U29302 (N_29302,N_27516,N_27918);
nand U29303 (N_29303,N_27965,N_27059);
nor U29304 (N_29304,N_27763,N_28173);
nor U29305 (N_29305,N_28184,N_27503);
nand U29306 (N_29306,N_28443,N_27073);
and U29307 (N_29307,N_28428,N_27696);
xnor U29308 (N_29308,N_28182,N_27855);
and U29309 (N_29309,N_28245,N_27404);
or U29310 (N_29310,N_27295,N_28127);
or U29311 (N_29311,N_27386,N_27852);
nand U29312 (N_29312,N_28320,N_28136);
or U29313 (N_29313,N_27988,N_27266);
and U29314 (N_29314,N_27195,N_27746);
nand U29315 (N_29315,N_27684,N_27107);
xor U29316 (N_29316,N_27379,N_27613);
and U29317 (N_29317,N_27209,N_28157);
and U29318 (N_29318,N_27691,N_28125);
or U29319 (N_29319,N_27889,N_27586);
or U29320 (N_29320,N_27958,N_27673);
nand U29321 (N_29321,N_27013,N_27179);
or U29322 (N_29322,N_28146,N_27142);
nand U29323 (N_29323,N_27336,N_27801);
nand U29324 (N_29324,N_27484,N_27171);
or U29325 (N_29325,N_27522,N_28145);
or U29326 (N_29326,N_27612,N_27127);
xnor U29327 (N_29327,N_27413,N_27390);
or U29328 (N_29328,N_27849,N_27339);
xor U29329 (N_29329,N_27194,N_27141);
nor U29330 (N_29330,N_27762,N_27921);
nand U29331 (N_29331,N_28122,N_27707);
nand U29332 (N_29332,N_27754,N_27918);
xnor U29333 (N_29333,N_28192,N_27068);
or U29334 (N_29334,N_27676,N_27011);
and U29335 (N_29335,N_28303,N_27348);
xnor U29336 (N_29336,N_28222,N_27675);
nand U29337 (N_29337,N_27597,N_27936);
xnor U29338 (N_29338,N_28389,N_28278);
or U29339 (N_29339,N_28484,N_28357);
nor U29340 (N_29340,N_27313,N_27929);
nand U29341 (N_29341,N_28314,N_27253);
or U29342 (N_29342,N_27992,N_28464);
nand U29343 (N_29343,N_28430,N_27392);
and U29344 (N_29344,N_27479,N_28355);
nand U29345 (N_29345,N_27388,N_28029);
or U29346 (N_29346,N_27033,N_28357);
nor U29347 (N_29347,N_27365,N_27684);
and U29348 (N_29348,N_27501,N_27261);
nor U29349 (N_29349,N_27958,N_27335);
and U29350 (N_29350,N_28300,N_27608);
nand U29351 (N_29351,N_28299,N_27398);
nor U29352 (N_29352,N_28184,N_27490);
nor U29353 (N_29353,N_28264,N_27754);
xor U29354 (N_29354,N_27576,N_27946);
nor U29355 (N_29355,N_27910,N_27622);
nor U29356 (N_29356,N_28466,N_27460);
or U29357 (N_29357,N_27823,N_27400);
nor U29358 (N_29358,N_28036,N_27084);
nor U29359 (N_29359,N_27686,N_27156);
nor U29360 (N_29360,N_27499,N_28370);
or U29361 (N_29361,N_27104,N_27379);
nand U29362 (N_29362,N_27719,N_28407);
xnor U29363 (N_29363,N_27753,N_28260);
nand U29364 (N_29364,N_27278,N_27768);
nand U29365 (N_29365,N_27984,N_27965);
nand U29366 (N_29366,N_27251,N_27935);
xnor U29367 (N_29367,N_28216,N_27165);
xor U29368 (N_29368,N_27892,N_28123);
nand U29369 (N_29369,N_27860,N_27697);
nor U29370 (N_29370,N_27880,N_28065);
or U29371 (N_29371,N_27167,N_28012);
nand U29372 (N_29372,N_28053,N_28118);
nand U29373 (N_29373,N_27595,N_28392);
xnor U29374 (N_29374,N_27986,N_27167);
nor U29375 (N_29375,N_28235,N_27450);
nor U29376 (N_29376,N_27277,N_27807);
or U29377 (N_29377,N_27958,N_27350);
xor U29378 (N_29378,N_28232,N_27504);
xor U29379 (N_29379,N_27800,N_27476);
nand U29380 (N_29380,N_27666,N_27525);
nor U29381 (N_29381,N_27869,N_27824);
and U29382 (N_29382,N_28131,N_28005);
and U29383 (N_29383,N_27389,N_28430);
and U29384 (N_29384,N_27077,N_28395);
xnor U29385 (N_29385,N_27868,N_27068);
xor U29386 (N_29386,N_27686,N_27231);
or U29387 (N_29387,N_28022,N_27321);
and U29388 (N_29388,N_27705,N_28009);
or U29389 (N_29389,N_27318,N_27321);
xnor U29390 (N_29390,N_27370,N_28131);
or U29391 (N_29391,N_27289,N_28390);
xnor U29392 (N_29392,N_27867,N_28487);
nor U29393 (N_29393,N_28239,N_27451);
or U29394 (N_29394,N_27410,N_27168);
and U29395 (N_29395,N_28331,N_28249);
or U29396 (N_29396,N_27537,N_27212);
and U29397 (N_29397,N_27391,N_27662);
and U29398 (N_29398,N_28470,N_27455);
nor U29399 (N_29399,N_27134,N_27403);
and U29400 (N_29400,N_27016,N_27977);
or U29401 (N_29401,N_27876,N_27106);
nand U29402 (N_29402,N_28221,N_28075);
and U29403 (N_29403,N_28035,N_27447);
or U29404 (N_29404,N_28239,N_27384);
nor U29405 (N_29405,N_28150,N_27769);
nor U29406 (N_29406,N_27414,N_27544);
or U29407 (N_29407,N_27835,N_27802);
xor U29408 (N_29408,N_28032,N_27877);
xnor U29409 (N_29409,N_27835,N_28079);
xor U29410 (N_29410,N_28334,N_27540);
nor U29411 (N_29411,N_28309,N_27755);
xor U29412 (N_29412,N_28202,N_28206);
nor U29413 (N_29413,N_27401,N_27275);
nand U29414 (N_29414,N_27199,N_28197);
or U29415 (N_29415,N_27228,N_28006);
or U29416 (N_29416,N_27688,N_27382);
xnor U29417 (N_29417,N_27880,N_28244);
nand U29418 (N_29418,N_28344,N_28146);
or U29419 (N_29419,N_27957,N_27240);
xor U29420 (N_29420,N_27149,N_27966);
xnor U29421 (N_29421,N_27798,N_28331);
and U29422 (N_29422,N_27386,N_27097);
nand U29423 (N_29423,N_27927,N_28235);
nand U29424 (N_29424,N_27398,N_27114);
nor U29425 (N_29425,N_27432,N_27749);
nor U29426 (N_29426,N_27354,N_28274);
nand U29427 (N_29427,N_27952,N_27698);
and U29428 (N_29428,N_27894,N_27613);
nand U29429 (N_29429,N_27217,N_28174);
nand U29430 (N_29430,N_28468,N_28334);
xnor U29431 (N_29431,N_27792,N_28168);
or U29432 (N_29432,N_27120,N_27714);
nor U29433 (N_29433,N_27334,N_28088);
and U29434 (N_29434,N_28240,N_27360);
or U29435 (N_29435,N_27432,N_27889);
nor U29436 (N_29436,N_28087,N_28407);
nand U29437 (N_29437,N_27994,N_27167);
xor U29438 (N_29438,N_27548,N_27374);
and U29439 (N_29439,N_27276,N_27887);
xnor U29440 (N_29440,N_27625,N_28070);
xnor U29441 (N_29441,N_27169,N_27138);
and U29442 (N_29442,N_28077,N_27285);
nor U29443 (N_29443,N_28209,N_27204);
and U29444 (N_29444,N_28119,N_27066);
and U29445 (N_29445,N_27715,N_27661);
nand U29446 (N_29446,N_27882,N_27994);
or U29447 (N_29447,N_27044,N_27138);
and U29448 (N_29448,N_28032,N_27325);
xnor U29449 (N_29449,N_27432,N_27992);
xor U29450 (N_29450,N_28315,N_27178);
xnor U29451 (N_29451,N_28051,N_27042);
xor U29452 (N_29452,N_27961,N_27099);
nor U29453 (N_29453,N_27661,N_28411);
or U29454 (N_29454,N_27027,N_28341);
and U29455 (N_29455,N_27467,N_27104);
nor U29456 (N_29456,N_27217,N_28219);
or U29457 (N_29457,N_27044,N_27173);
or U29458 (N_29458,N_28452,N_27896);
and U29459 (N_29459,N_28285,N_28395);
nand U29460 (N_29460,N_27416,N_27759);
nor U29461 (N_29461,N_27259,N_28104);
xnor U29462 (N_29462,N_27990,N_27006);
nor U29463 (N_29463,N_28473,N_27331);
nand U29464 (N_29464,N_27175,N_27255);
xnor U29465 (N_29465,N_27140,N_27445);
and U29466 (N_29466,N_27324,N_27726);
or U29467 (N_29467,N_27690,N_28314);
nand U29468 (N_29468,N_28440,N_27805);
nand U29469 (N_29469,N_27840,N_28256);
nor U29470 (N_29470,N_27229,N_27527);
and U29471 (N_29471,N_27592,N_28426);
xor U29472 (N_29472,N_28119,N_28275);
xor U29473 (N_29473,N_27348,N_27069);
nand U29474 (N_29474,N_28373,N_27754);
and U29475 (N_29475,N_27850,N_27544);
or U29476 (N_29476,N_27483,N_27190);
nor U29477 (N_29477,N_27850,N_27699);
and U29478 (N_29478,N_27902,N_27107);
xnor U29479 (N_29479,N_27705,N_27099);
xnor U29480 (N_29480,N_28075,N_27319);
and U29481 (N_29481,N_27855,N_27079);
nand U29482 (N_29482,N_28107,N_28113);
nor U29483 (N_29483,N_27891,N_27709);
nor U29484 (N_29484,N_27943,N_27370);
and U29485 (N_29485,N_27672,N_27919);
nor U29486 (N_29486,N_27820,N_27245);
or U29487 (N_29487,N_28081,N_27407);
and U29488 (N_29488,N_27671,N_27804);
or U29489 (N_29489,N_28438,N_27863);
or U29490 (N_29490,N_27112,N_28377);
nand U29491 (N_29491,N_27794,N_28431);
xor U29492 (N_29492,N_27802,N_28414);
xor U29493 (N_29493,N_27004,N_27119);
and U29494 (N_29494,N_28303,N_28409);
nor U29495 (N_29495,N_27361,N_27688);
nor U29496 (N_29496,N_27718,N_28275);
or U29497 (N_29497,N_27311,N_27893);
or U29498 (N_29498,N_27285,N_28447);
nand U29499 (N_29499,N_27107,N_27141);
xor U29500 (N_29500,N_27584,N_27344);
or U29501 (N_29501,N_28275,N_27657);
nand U29502 (N_29502,N_28441,N_27200);
nor U29503 (N_29503,N_27859,N_27906);
xor U29504 (N_29504,N_28058,N_27173);
nor U29505 (N_29505,N_27454,N_27407);
or U29506 (N_29506,N_28374,N_28359);
xor U29507 (N_29507,N_27479,N_27430);
xor U29508 (N_29508,N_27259,N_27269);
nor U29509 (N_29509,N_27783,N_27749);
and U29510 (N_29510,N_27154,N_28425);
xor U29511 (N_29511,N_27970,N_28202);
or U29512 (N_29512,N_27827,N_27976);
nand U29513 (N_29513,N_28495,N_28036);
nand U29514 (N_29514,N_28271,N_28415);
nor U29515 (N_29515,N_28099,N_27445);
nand U29516 (N_29516,N_27050,N_27423);
or U29517 (N_29517,N_27971,N_27062);
xor U29518 (N_29518,N_27130,N_27316);
and U29519 (N_29519,N_27644,N_27179);
xor U29520 (N_29520,N_27397,N_27085);
nand U29521 (N_29521,N_27915,N_28136);
and U29522 (N_29522,N_28018,N_27169);
xor U29523 (N_29523,N_27423,N_28005);
or U29524 (N_29524,N_27818,N_28173);
nand U29525 (N_29525,N_27309,N_27338);
xor U29526 (N_29526,N_27043,N_27957);
nand U29527 (N_29527,N_27726,N_28054);
or U29528 (N_29528,N_27909,N_27639);
and U29529 (N_29529,N_27636,N_28324);
and U29530 (N_29530,N_27547,N_27561);
and U29531 (N_29531,N_27945,N_28411);
nand U29532 (N_29532,N_27018,N_28444);
and U29533 (N_29533,N_28031,N_27659);
nand U29534 (N_29534,N_27877,N_27398);
xnor U29535 (N_29535,N_27794,N_27705);
nor U29536 (N_29536,N_27362,N_27313);
or U29537 (N_29537,N_27141,N_27599);
xor U29538 (N_29538,N_27184,N_27180);
or U29539 (N_29539,N_27697,N_28444);
and U29540 (N_29540,N_27243,N_28383);
xor U29541 (N_29541,N_27314,N_27732);
or U29542 (N_29542,N_27496,N_27281);
nand U29543 (N_29543,N_28300,N_28136);
and U29544 (N_29544,N_28066,N_28398);
and U29545 (N_29545,N_27009,N_27759);
xnor U29546 (N_29546,N_28349,N_28126);
nor U29547 (N_29547,N_28056,N_27201);
nor U29548 (N_29548,N_27013,N_27260);
and U29549 (N_29549,N_27847,N_27371);
or U29550 (N_29550,N_28276,N_27241);
or U29551 (N_29551,N_28431,N_27775);
nand U29552 (N_29552,N_27574,N_27248);
xor U29553 (N_29553,N_28152,N_28471);
nand U29554 (N_29554,N_27020,N_27265);
and U29555 (N_29555,N_27663,N_28190);
or U29556 (N_29556,N_27676,N_27586);
nor U29557 (N_29557,N_27841,N_27810);
and U29558 (N_29558,N_27291,N_28481);
and U29559 (N_29559,N_27089,N_28402);
xnor U29560 (N_29560,N_27634,N_27618);
nor U29561 (N_29561,N_28246,N_27932);
and U29562 (N_29562,N_28202,N_27675);
xnor U29563 (N_29563,N_27430,N_27721);
and U29564 (N_29564,N_27124,N_27609);
nor U29565 (N_29565,N_27104,N_27992);
xor U29566 (N_29566,N_28295,N_27429);
nand U29567 (N_29567,N_27398,N_27557);
nor U29568 (N_29568,N_27592,N_28221);
and U29569 (N_29569,N_27317,N_28298);
nor U29570 (N_29570,N_28363,N_28279);
nor U29571 (N_29571,N_27961,N_27199);
xnor U29572 (N_29572,N_28134,N_27040);
xor U29573 (N_29573,N_27806,N_27735);
nand U29574 (N_29574,N_28148,N_27204);
xnor U29575 (N_29575,N_27950,N_27294);
and U29576 (N_29576,N_27472,N_27496);
nand U29577 (N_29577,N_27578,N_27112);
or U29578 (N_29578,N_28051,N_28159);
nand U29579 (N_29579,N_27554,N_28110);
and U29580 (N_29580,N_27260,N_28067);
xnor U29581 (N_29581,N_27730,N_28066);
nor U29582 (N_29582,N_28048,N_27337);
and U29583 (N_29583,N_27139,N_27967);
or U29584 (N_29584,N_28211,N_27680);
nand U29585 (N_29585,N_28327,N_27544);
nand U29586 (N_29586,N_28069,N_28101);
nor U29587 (N_29587,N_27827,N_27955);
and U29588 (N_29588,N_27020,N_27450);
and U29589 (N_29589,N_28193,N_27503);
nor U29590 (N_29590,N_27942,N_27640);
and U29591 (N_29591,N_27949,N_28016);
nor U29592 (N_29592,N_27821,N_28097);
or U29593 (N_29593,N_27243,N_27221);
nand U29594 (N_29594,N_27551,N_27981);
nor U29595 (N_29595,N_27153,N_27593);
xor U29596 (N_29596,N_28310,N_27040);
nor U29597 (N_29597,N_27322,N_28334);
nand U29598 (N_29598,N_27983,N_27313);
or U29599 (N_29599,N_28432,N_27822);
xnor U29600 (N_29600,N_27248,N_28493);
xor U29601 (N_29601,N_27606,N_28176);
and U29602 (N_29602,N_28146,N_28038);
and U29603 (N_29603,N_27602,N_27341);
nand U29604 (N_29604,N_27952,N_28099);
or U29605 (N_29605,N_27386,N_28042);
xor U29606 (N_29606,N_27740,N_27920);
or U29607 (N_29607,N_27919,N_27311);
or U29608 (N_29608,N_27120,N_27787);
or U29609 (N_29609,N_27619,N_27624);
nand U29610 (N_29610,N_28148,N_28413);
nand U29611 (N_29611,N_27587,N_28254);
nor U29612 (N_29612,N_28125,N_27608);
nor U29613 (N_29613,N_27338,N_28426);
xor U29614 (N_29614,N_27858,N_28000);
or U29615 (N_29615,N_27092,N_27339);
and U29616 (N_29616,N_27403,N_27040);
or U29617 (N_29617,N_27823,N_27913);
nand U29618 (N_29618,N_28428,N_28224);
and U29619 (N_29619,N_27971,N_27702);
and U29620 (N_29620,N_27994,N_27324);
nor U29621 (N_29621,N_27491,N_27574);
xor U29622 (N_29622,N_27865,N_27463);
nand U29623 (N_29623,N_27724,N_27108);
and U29624 (N_29624,N_27999,N_27362);
or U29625 (N_29625,N_27511,N_27491);
nor U29626 (N_29626,N_27035,N_28269);
or U29627 (N_29627,N_27508,N_27086);
and U29628 (N_29628,N_28387,N_28322);
or U29629 (N_29629,N_27884,N_27526);
nand U29630 (N_29630,N_27275,N_27460);
or U29631 (N_29631,N_28228,N_28077);
or U29632 (N_29632,N_28301,N_28032);
nor U29633 (N_29633,N_27478,N_28201);
xor U29634 (N_29634,N_27717,N_27077);
nor U29635 (N_29635,N_28347,N_28477);
nand U29636 (N_29636,N_27583,N_28306);
nor U29637 (N_29637,N_27448,N_28344);
nand U29638 (N_29638,N_27919,N_28451);
and U29639 (N_29639,N_27741,N_27711);
nor U29640 (N_29640,N_27700,N_27466);
and U29641 (N_29641,N_27093,N_27012);
or U29642 (N_29642,N_27533,N_27774);
and U29643 (N_29643,N_27199,N_27782);
nor U29644 (N_29644,N_27742,N_27007);
and U29645 (N_29645,N_27799,N_27775);
nor U29646 (N_29646,N_27559,N_28012);
nor U29647 (N_29647,N_27786,N_27609);
nand U29648 (N_29648,N_27944,N_27078);
xnor U29649 (N_29649,N_27930,N_27421);
or U29650 (N_29650,N_28188,N_27821);
nor U29651 (N_29651,N_27059,N_27858);
nor U29652 (N_29652,N_27843,N_27947);
nor U29653 (N_29653,N_27499,N_27938);
and U29654 (N_29654,N_28263,N_27666);
xor U29655 (N_29655,N_28135,N_27694);
nor U29656 (N_29656,N_27275,N_27481);
nand U29657 (N_29657,N_27468,N_27202);
nand U29658 (N_29658,N_27030,N_28235);
nor U29659 (N_29659,N_28451,N_27109);
or U29660 (N_29660,N_27406,N_27646);
nand U29661 (N_29661,N_28104,N_27642);
and U29662 (N_29662,N_28254,N_28262);
or U29663 (N_29663,N_27955,N_27432);
xnor U29664 (N_29664,N_28293,N_27751);
xnor U29665 (N_29665,N_27467,N_27982);
nor U29666 (N_29666,N_28306,N_27509);
or U29667 (N_29667,N_28243,N_27093);
or U29668 (N_29668,N_28199,N_27756);
or U29669 (N_29669,N_28388,N_27857);
and U29670 (N_29670,N_27221,N_27522);
nand U29671 (N_29671,N_28058,N_28431);
xnor U29672 (N_29672,N_27988,N_27857);
nand U29673 (N_29673,N_27229,N_28278);
xor U29674 (N_29674,N_28327,N_27394);
or U29675 (N_29675,N_28015,N_27546);
and U29676 (N_29676,N_27619,N_28123);
and U29677 (N_29677,N_27408,N_27280);
nand U29678 (N_29678,N_27991,N_27139);
nand U29679 (N_29679,N_27300,N_27576);
nor U29680 (N_29680,N_27765,N_27977);
xnor U29681 (N_29681,N_27091,N_28429);
xnor U29682 (N_29682,N_27682,N_28184);
and U29683 (N_29683,N_27295,N_27210);
nand U29684 (N_29684,N_27930,N_28425);
and U29685 (N_29685,N_28335,N_27644);
nand U29686 (N_29686,N_27068,N_27926);
and U29687 (N_29687,N_28453,N_27791);
and U29688 (N_29688,N_27488,N_27076);
nor U29689 (N_29689,N_27260,N_27174);
xnor U29690 (N_29690,N_27033,N_27690);
and U29691 (N_29691,N_27241,N_27502);
nand U29692 (N_29692,N_28099,N_27903);
xor U29693 (N_29693,N_28388,N_27788);
or U29694 (N_29694,N_27766,N_28284);
nand U29695 (N_29695,N_27325,N_27509);
xnor U29696 (N_29696,N_27862,N_27009);
and U29697 (N_29697,N_27165,N_28018);
nand U29698 (N_29698,N_27211,N_27134);
xor U29699 (N_29699,N_27187,N_28126);
nor U29700 (N_29700,N_27515,N_27916);
nor U29701 (N_29701,N_27821,N_28240);
and U29702 (N_29702,N_27942,N_27673);
or U29703 (N_29703,N_27426,N_27065);
and U29704 (N_29704,N_27316,N_28257);
nand U29705 (N_29705,N_27636,N_28041);
nor U29706 (N_29706,N_27320,N_27849);
or U29707 (N_29707,N_27532,N_27255);
or U29708 (N_29708,N_27065,N_28047);
xor U29709 (N_29709,N_28419,N_27881);
or U29710 (N_29710,N_27907,N_28335);
nand U29711 (N_29711,N_27735,N_28056);
or U29712 (N_29712,N_27698,N_28491);
nor U29713 (N_29713,N_28211,N_28018);
nand U29714 (N_29714,N_27753,N_27669);
xnor U29715 (N_29715,N_27101,N_27678);
and U29716 (N_29716,N_28399,N_28228);
and U29717 (N_29717,N_27688,N_27570);
or U29718 (N_29718,N_27374,N_27053);
xor U29719 (N_29719,N_27900,N_28212);
xor U29720 (N_29720,N_28405,N_28018);
nand U29721 (N_29721,N_28058,N_27558);
nor U29722 (N_29722,N_28183,N_27278);
nor U29723 (N_29723,N_28146,N_27056);
nor U29724 (N_29724,N_27898,N_27375);
or U29725 (N_29725,N_27941,N_27862);
nand U29726 (N_29726,N_28478,N_27499);
xnor U29727 (N_29727,N_27854,N_27412);
nor U29728 (N_29728,N_28420,N_28082);
or U29729 (N_29729,N_27418,N_27010);
xnor U29730 (N_29730,N_28054,N_28098);
nand U29731 (N_29731,N_27316,N_27500);
and U29732 (N_29732,N_27553,N_28453);
and U29733 (N_29733,N_28147,N_27997);
xor U29734 (N_29734,N_28480,N_28395);
nand U29735 (N_29735,N_28358,N_27054);
nor U29736 (N_29736,N_27037,N_27725);
nand U29737 (N_29737,N_27075,N_27913);
or U29738 (N_29738,N_27930,N_28291);
nand U29739 (N_29739,N_28050,N_27854);
xnor U29740 (N_29740,N_27258,N_27000);
nand U29741 (N_29741,N_27692,N_28234);
and U29742 (N_29742,N_28103,N_27068);
nand U29743 (N_29743,N_27495,N_28135);
nand U29744 (N_29744,N_27077,N_27161);
or U29745 (N_29745,N_27987,N_27757);
or U29746 (N_29746,N_28328,N_27191);
nand U29747 (N_29747,N_27994,N_27495);
nor U29748 (N_29748,N_27851,N_27834);
or U29749 (N_29749,N_27539,N_27244);
nor U29750 (N_29750,N_27415,N_27063);
xnor U29751 (N_29751,N_27353,N_27386);
or U29752 (N_29752,N_28387,N_27768);
nand U29753 (N_29753,N_28194,N_27752);
nor U29754 (N_29754,N_28332,N_28018);
nand U29755 (N_29755,N_28156,N_27939);
or U29756 (N_29756,N_28106,N_27272);
nand U29757 (N_29757,N_27157,N_27341);
xor U29758 (N_29758,N_27276,N_27243);
xnor U29759 (N_29759,N_27639,N_27200);
or U29760 (N_29760,N_27462,N_27413);
or U29761 (N_29761,N_27619,N_28205);
and U29762 (N_29762,N_27828,N_28263);
or U29763 (N_29763,N_27698,N_27025);
nand U29764 (N_29764,N_27666,N_27939);
nor U29765 (N_29765,N_28338,N_28048);
or U29766 (N_29766,N_27518,N_28120);
xor U29767 (N_29767,N_28154,N_27435);
nor U29768 (N_29768,N_27632,N_28101);
xnor U29769 (N_29769,N_28131,N_28054);
nor U29770 (N_29770,N_28105,N_27252);
and U29771 (N_29771,N_27678,N_27289);
or U29772 (N_29772,N_28334,N_27728);
xor U29773 (N_29773,N_27456,N_27732);
nor U29774 (N_29774,N_28116,N_28265);
and U29775 (N_29775,N_27203,N_27982);
nor U29776 (N_29776,N_27569,N_28315);
nor U29777 (N_29777,N_27605,N_27105);
nor U29778 (N_29778,N_27177,N_27745);
nor U29779 (N_29779,N_28393,N_27197);
nor U29780 (N_29780,N_27665,N_27785);
xor U29781 (N_29781,N_27873,N_27668);
xor U29782 (N_29782,N_28246,N_28016);
and U29783 (N_29783,N_27882,N_27108);
or U29784 (N_29784,N_28403,N_27397);
nor U29785 (N_29785,N_27708,N_27811);
or U29786 (N_29786,N_27740,N_27282);
or U29787 (N_29787,N_28042,N_28300);
nand U29788 (N_29788,N_27051,N_28364);
and U29789 (N_29789,N_28321,N_27770);
and U29790 (N_29790,N_27463,N_27938);
nand U29791 (N_29791,N_27407,N_27228);
xor U29792 (N_29792,N_27642,N_28401);
nand U29793 (N_29793,N_28090,N_27229);
nand U29794 (N_29794,N_27786,N_27989);
nor U29795 (N_29795,N_27793,N_27858);
nand U29796 (N_29796,N_28324,N_27006);
nor U29797 (N_29797,N_27626,N_27586);
or U29798 (N_29798,N_28254,N_27282);
or U29799 (N_29799,N_28302,N_27027);
xor U29800 (N_29800,N_28031,N_27352);
and U29801 (N_29801,N_28186,N_27159);
xnor U29802 (N_29802,N_28315,N_28063);
and U29803 (N_29803,N_28275,N_27826);
or U29804 (N_29804,N_27978,N_27144);
and U29805 (N_29805,N_28149,N_27845);
xor U29806 (N_29806,N_28065,N_27412);
nor U29807 (N_29807,N_28274,N_27478);
xnor U29808 (N_29808,N_28245,N_27967);
and U29809 (N_29809,N_27741,N_27797);
nor U29810 (N_29810,N_27910,N_27822);
nand U29811 (N_29811,N_27473,N_27604);
xor U29812 (N_29812,N_28082,N_28059);
nor U29813 (N_29813,N_28076,N_27620);
or U29814 (N_29814,N_27865,N_27385);
nor U29815 (N_29815,N_27326,N_27217);
and U29816 (N_29816,N_27224,N_28012);
nor U29817 (N_29817,N_27158,N_28203);
and U29818 (N_29818,N_27415,N_28054);
or U29819 (N_29819,N_28444,N_27308);
or U29820 (N_29820,N_27259,N_27396);
and U29821 (N_29821,N_27308,N_28134);
xor U29822 (N_29822,N_28116,N_28458);
or U29823 (N_29823,N_27114,N_27943);
nor U29824 (N_29824,N_27385,N_27343);
xor U29825 (N_29825,N_27819,N_28201);
nor U29826 (N_29826,N_27700,N_27200);
nor U29827 (N_29827,N_27744,N_28101);
and U29828 (N_29828,N_27744,N_28193);
xnor U29829 (N_29829,N_27026,N_27326);
or U29830 (N_29830,N_27740,N_27166);
nor U29831 (N_29831,N_27520,N_27453);
nor U29832 (N_29832,N_28215,N_27083);
nand U29833 (N_29833,N_27584,N_27704);
nor U29834 (N_29834,N_27273,N_27855);
or U29835 (N_29835,N_28442,N_27439);
nand U29836 (N_29836,N_28039,N_28077);
nor U29837 (N_29837,N_27241,N_27037);
nor U29838 (N_29838,N_28076,N_27911);
and U29839 (N_29839,N_27305,N_27884);
and U29840 (N_29840,N_27618,N_27112);
or U29841 (N_29841,N_27422,N_27959);
nor U29842 (N_29842,N_27677,N_28185);
nor U29843 (N_29843,N_27690,N_27496);
xnor U29844 (N_29844,N_27487,N_27844);
nor U29845 (N_29845,N_28004,N_28383);
and U29846 (N_29846,N_27884,N_28253);
nor U29847 (N_29847,N_27055,N_28345);
nor U29848 (N_29848,N_28127,N_27841);
xor U29849 (N_29849,N_28470,N_27676);
nor U29850 (N_29850,N_27736,N_28159);
or U29851 (N_29851,N_27499,N_28328);
nor U29852 (N_29852,N_27041,N_27938);
nand U29853 (N_29853,N_27850,N_27751);
nand U29854 (N_29854,N_27771,N_28165);
or U29855 (N_29855,N_27880,N_27768);
nand U29856 (N_29856,N_27451,N_28299);
nand U29857 (N_29857,N_28194,N_28435);
and U29858 (N_29858,N_28113,N_27989);
and U29859 (N_29859,N_27237,N_27962);
and U29860 (N_29860,N_28472,N_27244);
and U29861 (N_29861,N_27541,N_27619);
and U29862 (N_29862,N_28003,N_27783);
xor U29863 (N_29863,N_28247,N_28157);
and U29864 (N_29864,N_27236,N_27128);
nor U29865 (N_29865,N_27093,N_27394);
xor U29866 (N_29866,N_27430,N_27216);
or U29867 (N_29867,N_27879,N_27450);
xnor U29868 (N_29868,N_27011,N_28202);
or U29869 (N_29869,N_27055,N_27477);
or U29870 (N_29870,N_27669,N_27482);
nor U29871 (N_29871,N_28303,N_27061);
or U29872 (N_29872,N_27210,N_27725);
nor U29873 (N_29873,N_28074,N_28308);
nand U29874 (N_29874,N_27530,N_27234);
or U29875 (N_29875,N_27898,N_27864);
nand U29876 (N_29876,N_27514,N_27347);
or U29877 (N_29877,N_27264,N_27124);
and U29878 (N_29878,N_27727,N_27432);
xnor U29879 (N_29879,N_27188,N_27914);
and U29880 (N_29880,N_27041,N_28474);
nand U29881 (N_29881,N_28400,N_27050);
or U29882 (N_29882,N_28427,N_28144);
xnor U29883 (N_29883,N_27292,N_27108);
xnor U29884 (N_29884,N_27647,N_27430);
nor U29885 (N_29885,N_27624,N_27116);
nor U29886 (N_29886,N_27311,N_28464);
xnor U29887 (N_29887,N_27598,N_27715);
xor U29888 (N_29888,N_28226,N_27269);
nor U29889 (N_29889,N_27395,N_27030);
and U29890 (N_29890,N_27879,N_27570);
nand U29891 (N_29891,N_27273,N_27323);
nand U29892 (N_29892,N_27326,N_27396);
nand U29893 (N_29893,N_27527,N_27491);
or U29894 (N_29894,N_27994,N_27253);
or U29895 (N_29895,N_27084,N_28182);
xnor U29896 (N_29896,N_27050,N_27660);
nand U29897 (N_29897,N_27826,N_28010);
xnor U29898 (N_29898,N_27621,N_27100);
nor U29899 (N_29899,N_27342,N_27180);
nor U29900 (N_29900,N_27791,N_27332);
or U29901 (N_29901,N_27983,N_27821);
nor U29902 (N_29902,N_27811,N_28405);
nor U29903 (N_29903,N_27776,N_27550);
nand U29904 (N_29904,N_27124,N_27584);
xor U29905 (N_29905,N_27387,N_27122);
or U29906 (N_29906,N_28022,N_27746);
nand U29907 (N_29907,N_27802,N_27142);
nor U29908 (N_29908,N_27584,N_27719);
xnor U29909 (N_29909,N_27920,N_27824);
and U29910 (N_29910,N_28378,N_28047);
nor U29911 (N_29911,N_28052,N_27549);
xnor U29912 (N_29912,N_27658,N_27536);
or U29913 (N_29913,N_27220,N_27375);
nor U29914 (N_29914,N_28066,N_28330);
nand U29915 (N_29915,N_27202,N_27965);
or U29916 (N_29916,N_27109,N_27706);
and U29917 (N_29917,N_27904,N_27039);
nor U29918 (N_29918,N_28449,N_27670);
nand U29919 (N_29919,N_28202,N_28176);
xnor U29920 (N_29920,N_27704,N_27318);
and U29921 (N_29921,N_28086,N_28240);
and U29922 (N_29922,N_28030,N_28400);
and U29923 (N_29923,N_28185,N_28016);
nand U29924 (N_29924,N_28024,N_28049);
nor U29925 (N_29925,N_28154,N_28460);
or U29926 (N_29926,N_27516,N_27941);
or U29927 (N_29927,N_27704,N_27636);
nand U29928 (N_29928,N_27222,N_27346);
and U29929 (N_29929,N_27758,N_27847);
and U29930 (N_29930,N_27649,N_27571);
nand U29931 (N_29931,N_27685,N_28023);
xor U29932 (N_29932,N_27010,N_27967);
xnor U29933 (N_29933,N_27000,N_28370);
and U29934 (N_29934,N_28420,N_28029);
or U29935 (N_29935,N_27495,N_28422);
xor U29936 (N_29936,N_27869,N_27214);
nand U29937 (N_29937,N_27445,N_27433);
nand U29938 (N_29938,N_27674,N_28100);
or U29939 (N_29939,N_27140,N_27689);
nor U29940 (N_29940,N_27570,N_27674);
or U29941 (N_29941,N_28337,N_27239);
nor U29942 (N_29942,N_27132,N_27654);
nor U29943 (N_29943,N_28337,N_27274);
or U29944 (N_29944,N_27309,N_28151);
or U29945 (N_29945,N_27912,N_28004);
nand U29946 (N_29946,N_27219,N_28029);
and U29947 (N_29947,N_28292,N_28110);
and U29948 (N_29948,N_28343,N_28401);
or U29949 (N_29949,N_28334,N_27361);
nand U29950 (N_29950,N_28410,N_27616);
nor U29951 (N_29951,N_28251,N_28386);
nand U29952 (N_29952,N_27926,N_27809);
nor U29953 (N_29953,N_27790,N_27736);
or U29954 (N_29954,N_27824,N_28172);
nor U29955 (N_29955,N_27427,N_28405);
or U29956 (N_29956,N_27546,N_27022);
nand U29957 (N_29957,N_28493,N_28305);
or U29958 (N_29958,N_27155,N_27895);
nor U29959 (N_29959,N_28143,N_27488);
or U29960 (N_29960,N_27482,N_27083);
or U29961 (N_29961,N_28061,N_27546);
or U29962 (N_29962,N_27489,N_28035);
or U29963 (N_29963,N_28308,N_27951);
or U29964 (N_29964,N_27995,N_27129);
and U29965 (N_29965,N_28149,N_27573);
and U29966 (N_29966,N_28073,N_27422);
nand U29967 (N_29967,N_27741,N_27519);
and U29968 (N_29968,N_27650,N_27903);
nor U29969 (N_29969,N_27925,N_27847);
or U29970 (N_29970,N_28091,N_27379);
and U29971 (N_29971,N_27890,N_27517);
and U29972 (N_29972,N_28004,N_27044);
nor U29973 (N_29973,N_27529,N_28047);
or U29974 (N_29974,N_27299,N_28109);
and U29975 (N_29975,N_27608,N_27685);
and U29976 (N_29976,N_27014,N_27892);
xor U29977 (N_29977,N_27434,N_27924);
xor U29978 (N_29978,N_27791,N_28144);
xnor U29979 (N_29979,N_27214,N_27356);
or U29980 (N_29980,N_27129,N_28120);
nand U29981 (N_29981,N_27603,N_28044);
and U29982 (N_29982,N_28049,N_27152);
and U29983 (N_29983,N_28354,N_27121);
and U29984 (N_29984,N_27479,N_27728);
and U29985 (N_29985,N_28458,N_28074);
nand U29986 (N_29986,N_27514,N_27600);
and U29987 (N_29987,N_27200,N_27307);
or U29988 (N_29988,N_28337,N_27347);
and U29989 (N_29989,N_27500,N_27679);
and U29990 (N_29990,N_27895,N_27352);
nor U29991 (N_29991,N_28263,N_28000);
xnor U29992 (N_29992,N_27708,N_27753);
or U29993 (N_29993,N_27779,N_28298);
nor U29994 (N_29994,N_27767,N_27811);
nand U29995 (N_29995,N_27231,N_28479);
xor U29996 (N_29996,N_27185,N_27880);
and U29997 (N_29997,N_27801,N_27314);
nand U29998 (N_29998,N_28330,N_27726);
nand U29999 (N_29999,N_27568,N_27063);
nand UO_0 (O_0,N_29166,N_29458);
or UO_1 (O_1,N_29586,N_29472);
nor UO_2 (O_2,N_28911,N_28538);
xnor UO_3 (O_3,N_29289,N_29482);
nor UO_4 (O_4,N_29639,N_29025);
xnor UO_5 (O_5,N_28716,N_29009);
xnor UO_6 (O_6,N_29741,N_29031);
or UO_7 (O_7,N_29450,N_28600);
nand UO_8 (O_8,N_28929,N_29777);
and UO_9 (O_9,N_28525,N_28815);
and UO_10 (O_10,N_29814,N_28517);
nor UO_11 (O_11,N_28833,N_28996);
xor UO_12 (O_12,N_29567,N_29818);
xnor UO_13 (O_13,N_29965,N_29211);
and UO_14 (O_14,N_29863,N_29996);
or UO_15 (O_15,N_29614,N_29561);
xor UO_16 (O_16,N_29419,N_29983);
or UO_17 (O_17,N_29109,N_28798);
xnor UO_18 (O_18,N_29684,N_29615);
nand UO_19 (O_19,N_29620,N_29499);
nand UO_20 (O_20,N_29445,N_29296);
or UO_21 (O_21,N_29701,N_29210);
nand UO_22 (O_22,N_28763,N_28635);
nor UO_23 (O_23,N_28808,N_29149);
nand UO_24 (O_24,N_29518,N_28662);
or UO_25 (O_25,N_29007,N_29866);
xnor UO_26 (O_26,N_29401,N_29422);
nand UO_27 (O_27,N_29033,N_29093);
or UO_28 (O_28,N_28947,N_28645);
and UO_29 (O_29,N_28641,N_29354);
nor UO_30 (O_30,N_29562,N_29541);
and UO_31 (O_31,N_29893,N_29896);
nand UO_32 (O_32,N_28725,N_28785);
xor UO_33 (O_33,N_29871,N_29105);
or UO_34 (O_34,N_29012,N_28856);
or UO_35 (O_35,N_28521,N_28807);
or UO_36 (O_36,N_29408,N_28570);
and UO_37 (O_37,N_29432,N_28657);
or UO_38 (O_38,N_28864,N_28842);
xor UO_39 (O_39,N_28787,N_29589);
nor UO_40 (O_40,N_29810,N_28784);
nor UO_41 (O_41,N_29717,N_28670);
or UO_42 (O_42,N_29125,N_28540);
nor UO_43 (O_43,N_29321,N_28762);
xnor UO_44 (O_44,N_29867,N_28953);
and UO_45 (O_45,N_29591,N_29413);
and UO_46 (O_46,N_29569,N_29100);
nand UO_47 (O_47,N_29629,N_29968);
or UO_48 (O_48,N_29427,N_29503);
nor UO_49 (O_49,N_29351,N_29074);
nor UO_50 (O_50,N_29170,N_29207);
or UO_51 (O_51,N_29146,N_29512);
nor UO_52 (O_52,N_28861,N_29409);
nor UO_53 (O_53,N_29131,N_29740);
or UO_54 (O_54,N_29295,N_29570);
nand UO_55 (O_55,N_29449,N_29440);
nand UO_56 (O_56,N_29302,N_28562);
and UO_57 (O_57,N_29221,N_29737);
nor UO_58 (O_58,N_29193,N_29697);
nor UO_59 (O_59,N_28544,N_29693);
nor UO_60 (O_60,N_28943,N_28745);
xor UO_61 (O_61,N_28906,N_28898);
or UO_62 (O_62,N_29659,N_29935);
and UO_63 (O_63,N_28971,N_28897);
and UO_64 (O_64,N_28862,N_29127);
and UO_65 (O_65,N_29997,N_29218);
xnor UO_66 (O_66,N_28688,N_29682);
or UO_67 (O_67,N_29575,N_28620);
or UO_68 (O_68,N_29635,N_29936);
xor UO_69 (O_69,N_29673,N_29085);
xor UO_70 (O_70,N_29494,N_29601);
nand UO_71 (O_71,N_29200,N_29714);
or UO_72 (O_72,N_28537,N_28788);
nor UO_73 (O_73,N_29642,N_29164);
or UO_74 (O_74,N_28919,N_28520);
nor UO_75 (O_75,N_28790,N_28847);
and UO_76 (O_76,N_28868,N_29630);
xnor UO_77 (O_77,N_29305,N_28758);
nand UO_78 (O_78,N_28951,N_29485);
xor UO_79 (O_79,N_28749,N_28841);
and UO_80 (O_80,N_29593,N_29262);
xnor UO_81 (O_81,N_29869,N_28985);
and UO_82 (O_82,N_29424,N_29725);
and UO_83 (O_83,N_29126,N_29830);
nand UO_84 (O_84,N_29515,N_29229);
or UO_85 (O_85,N_29723,N_29201);
or UO_86 (O_86,N_29197,N_28984);
nand UO_87 (O_87,N_29055,N_29568);
and UO_88 (O_88,N_28849,N_29802);
and UO_89 (O_89,N_29312,N_29969);
or UO_90 (O_90,N_29666,N_28845);
nand UO_91 (O_91,N_29395,N_29791);
nand UO_92 (O_92,N_29758,N_29045);
xor UO_93 (O_93,N_29124,N_29358);
and UO_94 (O_94,N_29719,N_29636);
and UO_95 (O_95,N_29171,N_29784);
and UO_96 (O_96,N_28902,N_29828);
or UO_97 (O_97,N_29405,N_28903);
and UO_98 (O_98,N_29683,N_28814);
or UO_99 (O_99,N_29751,N_28974);
and UO_100 (O_100,N_29939,N_28826);
or UO_101 (O_101,N_29565,N_29792);
or UO_102 (O_102,N_29334,N_29444);
xnor UO_103 (O_103,N_29026,N_29577);
and UO_104 (O_104,N_29469,N_29911);
xnor UO_105 (O_105,N_29471,N_28793);
nor UO_106 (O_106,N_28772,N_28811);
xnor UO_107 (O_107,N_28748,N_28939);
and UO_108 (O_108,N_29342,N_28590);
nor UO_109 (O_109,N_29613,N_29011);
or UO_110 (O_110,N_29744,N_29970);
nor UO_111 (O_111,N_29418,N_28873);
nor UO_112 (O_112,N_28977,N_28595);
nand UO_113 (O_113,N_29198,N_28923);
xor UO_114 (O_114,N_29677,N_29977);
xnor UO_115 (O_115,N_29195,N_29581);
and UO_116 (O_116,N_29919,N_28559);
or UO_117 (O_117,N_29319,N_29750);
or UO_118 (O_118,N_29648,N_29006);
nor UO_119 (O_119,N_29078,N_29436);
xor UO_120 (O_120,N_28764,N_29088);
nor UO_121 (O_121,N_29196,N_29550);
nor UO_122 (O_122,N_29769,N_28844);
and UO_123 (O_123,N_29098,N_29442);
nand UO_124 (O_124,N_29715,N_28970);
or UO_125 (O_125,N_28752,N_29421);
or UO_126 (O_126,N_29024,N_28846);
xnor UO_127 (O_127,N_29510,N_29584);
nor UO_128 (O_128,N_28995,N_29158);
xnor UO_129 (O_129,N_28778,N_29688);
and UO_130 (O_130,N_29174,N_29331);
nor UO_131 (O_131,N_29813,N_28742);
or UO_132 (O_132,N_28552,N_29580);
nand UO_133 (O_133,N_29803,N_28722);
nand UO_134 (O_134,N_28555,N_28687);
xor UO_135 (O_135,N_29689,N_28750);
and UO_136 (O_136,N_28805,N_29492);
nand UO_137 (O_137,N_28589,N_28816);
and UO_138 (O_138,N_29437,N_28770);
xnor UO_139 (O_139,N_29579,N_28592);
nand UO_140 (O_140,N_29854,N_29535);
xor UO_141 (O_141,N_29699,N_28850);
or UO_142 (O_142,N_28957,N_29256);
nand UO_143 (O_143,N_29459,N_28596);
xnor UO_144 (O_144,N_29900,N_28863);
nand UO_145 (O_145,N_29644,N_29425);
nor UO_146 (O_146,N_28606,N_29721);
nor UO_147 (O_147,N_29794,N_29379);
xor UO_148 (O_148,N_29215,N_29299);
or UO_149 (O_149,N_29861,N_29314);
nand UO_150 (O_150,N_29142,N_29381);
xor UO_151 (O_151,N_29003,N_29940);
and UO_152 (O_152,N_28536,N_29364);
or UO_153 (O_153,N_28693,N_28765);
xor UO_154 (O_154,N_29691,N_29129);
or UO_155 (O_155,N_29770,N_29778);
or UO_156 (O_156,N_29576,N_29343);
nor UO_157 (O_157,N_28691,N_29637);
xor UO_158 (O_158,N_28604,N_28678);
nor UO_159 (O_159,N_29353,N_28634);
nand UO_160 (O_160,N_28879,N_29134);
nor UO_161 (O_161,N_28619,N_29539);
and UO_162 (O_162,N_29764,N_29916);
and UO_163 (O_163,N_29806,N_28578);
and UO_164 (O_164,N_29999,N_29907);
or UO_165 (O_165,N_29044,N_29456);
xor UO_166 (O_166,N_29357,N_29759);
xnor UO_167 (O_167,N_29891,N_29558);
nor UO_168 (O_168,N_29220,N_28535);
or UO_169 (O_169,N_28932,N_29313);
and UO_170 (O_170,N_29847,N_28771);
nor UO_171 (O_171,N_29235,N_29527);
and UO_172 (O_172,N_29301,N_29671);
nor UO_173 (O_173,N_29141,N_28575);
and UO_174 (O_174,N_28505,N_29322);
and UO_175 (O_175,N_29300,N_29117);
xnor UO_176 (O_176,N_28777,N_29604);
nand UO_177 (O_177,N_29915,N_28918);
nand UO_178 (O_178,N_28603,N_28853);
xor UO_179 (O_179,N_29116,N_28551);
nand UO_180 (O_180,N_28999,N_29051);
nor UO_181 (O_181,N_28820,N_29260);
and UO_182 (O_182,N_29859,N_29955);
nand UO_183 (O_183,N_28727,N_29795);
and UO_184 (O_184,N_29392,N_29175);
and UO_185 (O_185,N_29731,N_28618);
or UO_186 (O_186,N_29239,N_29528);
nand UO_187 (O_187,N_28936,N_29611);
nand UO_188 (O_188,N_28528,N_29619);
and UO_189 (O_189,N_28924,N_29821);
and UO_190 (O_190,N_29061,N_29058);
xor UO_191 (O_191,N_28757,N_29933);
nand UO_192 (O_192,N_29360,N_29548);
xnor UO_193 (O_193,N_28602,N_28665);
or UO_194 (O_194,N_28891,N_28683);
nand UO_195 (O_195,N_29898,N_29243);
xnor UO_196 (O_196,N_29153,N_28900);
xor UO_197 (O_197,N_29797,N_29929);
or UO_198 (O_198,N_28714,N_28822);
and UO_199 (O_199,N_28515,N_29768);
nor UO_200 (O_200,N_29920,N_28741);
or UO_201 (O_201,N_29502,N_29836);
and UO_202 (O_202,N_28699,N_29519);
nand UO_203 (O_203,N_28531,N_29948);
or UO_204 (O_204,N_28534,N_29115);
or UO_205 (O_205,N_29206,N_29804);
and UO_206 (O_206,N_29530,N_28511);
nand UO_207 (O_207,N_28802,N_29678);
or UO_208 (O_208,N_28673,N_29441);
or UO_209 (O_209,N_29598,N_29038);
nor UO_210 (O_210,N_29888,N_28648);
xnor UO_211 (O_211,N_29367,N_29323);
and UO_212 (O_212,N_29008,N_29780);
nand UO_213 (O_213,N_28715,N_28663);
and UO_214 (O_214,N_28782,N_29909);
and UO_215 (O_215,N_29189,N_29255);
or UO_216 (O_216,N_29749,N_29724);
xnor UO_217 (O_217,N_29382,N_29934);
xnor UO_218 (O_218,N_29140,N_28940);
nor UO_219 (O_219,N_28610,N_29612);
nor UO_220 (O_220,N_29557,N_29698);
or UO_221 (O_221,N_28899,N_29692);
nand UO_222 (O_222,N_28712,N_29742);
and UO_223 (O_223,N_28916,N_28709);
xnor UO_224 (O_224,N_29583,N_29159);
nor UO_225 (O_225,N_29030,N_29710);
nand UO_226 (O_226,N_29087,N_29960);
and UO_227 (O_227,N_29374,N_29022);
nor UO_228 (O_228,N_28875,N_29798);
or UO_229 (O_229,N_29118,N_29230);
nor UO_230 (O_230,N_29138,N_29521);
or UO_231 (O_231,N_29549,N_28976);
nor UO_232 (O_232,N_29812,N_28956);
nor UO_233 (O_233,N_28866,N_28659);
xor UO_234 (O_234,N_29027,N_28732);
nor UO_235 (O_235,N_28871,N_28608);
or UO_236 (O_236,N_29417,N_29573);
or UO_237 (O_237,N_29820,N_29004);
or UO_238 (O_238,N_29001,N_29533);
or UO_239 (O_239,N_29137,N_29252);
and UO_240 (O_240,N_29873,N_29479);
nand UO_241 (O_241,N_29309,N_29407);
or UO_242 (O_242,N_28968,N_29973);
nand UO_243 (O_243,N_28708,N_29862);
nand UO_244 (O_244,N_29976,N_28622);
or UO_245 (O_245,N_29466,N_28859);
xor UO_246 (O_246,N_29212,N_29377);
nor UO_247 (O_247,N_28840,N_29059);
xnor UO_248 (O_248,N_29834,N_28692);
and UO_249 (O_249,N_28827,N_29028);
nor UO_250 (O_250,N_28623,N_29597);
or UO_251 (O_251,N_28804,N_29148);
xnor UO_252 (O_252,N_29072,N_29623);
nand UO_253 (O_253,N_29771,N_29506);
and UO_254 (O_254,N_29157,N_28768);
nand UO_255 (O_255,N_29853,N_29857);
or UO_256 (O_256,N_28931,N_29039);
or UO_257 (O_257,N_28601,N_28944);
xor UO_258 (O_258,N_29728,N_29464);
and UO_259 (O_259,N_29885,N_29345);
xor UO_260 (O_260,N_29776,N_29653);
and UO_261 (O_261,N_29040,N_29455);
or UO_262 (O_262,N_28955,N_29773);
nand UO_263 (O_263,N_29307,N_29881);
nand UO_264 (O_264,N_29297,N_29130);
and UO_265 (O_265,N_28605,N_29278);
and UO_266 (O_266,N_29236,N_29808);
xnor UO_267 (O_267,N_29480,N_29348);
and UO_268 (O_268,N_29186,N_28935);
nand UO_269 (O_269,N_28922,N_29978);
or UO_270 (O_270,N_29384,N_29216);
xnor UO_271 (O_271,N_29429,N_28626);
or UO_272 (O_272,N_28921,N_29981);
nor UO_273 (O_273,N_29414,N_28574);
or UO_274 (O_274,N_29416,N_28513);
xor UO_275 (O_275,N_28860,N_29048);
nand UO_276 (O_276,N_29602,N_29679);
xnor UO_277 (O_277,N_28576,N_29089);
or UO_278 (O_278,N_28834,N_28887);
nor UO_279 (O_279,N_29700,N_29020);
nand UO_280 (O_280,N_28746,N_29617);
xnor UO_281 (O_281,N_29905,N_29766);
and UO_282 (O_282,N_29320,N_29918);
or UO_283 (O_283,N_28567,N_29095);
nand UO_284 (O_284,N_29757,N_29546);
and UO_285 (O_285,N_28915,N_29498);
nand UO_286 (O_286,N_29035,N_29283);
nand UO_287 (O_287,N_29694,N_29075);
nand UO_288 (O_288,N_29280,N_29961);
xnor UO_289 (O_289,N_29041,N_29454);
nand UO_290 (O_290,N_29014,N_29476);
nand UO_291 (O_291,N_28829,N_28877);
and UO_292 (O_292,N_29036,N_29327);
xor UO_293 (O_293,N_29463,N_29178);
or UO_294 (O_294,N_28883,N_29362);
or UO_295 (O_295,N_28710,N_29966);
nand UO_296 (O_296,N_28509,N_29281);
nand UO_297 (O_297,N_28945,N_29560);
xor UO_298 (O_298,N_28658,N_29091);
nor UO_299 (O_299,N_28754,N_28653);
nor UO_300 (O_300,N_28823,N_29308);
nor UO_301 (O_301,N_29956,N_29361);
xor UO_302 (O_302,N_29254,N_29288);
xor UO_303 (O_303,N_29690,N_29002);
or UO_304 (O_304,N_28783,N_29423);
or UO_305 (O_305,N_28967,N_29340);
nand UO_306 (O_306,N_29641,N_29034);
nor UO_307 (O_307,N_29021,N_29258);
nor UO_308 (O_308,N_28813,N_29815);
and UO_309 (O_309,N_29344,N_29337);
nor UO_310 (O_310,N_29073,N_28656);
or UO_311 (O_311,N_28809,N_28726);
or UO_312 (O_312,N_29858,N_28774);
and UO_313 (O_313,N_29160,N_29120);
and UO_314 (O_314,N_29964,N_29649);
nor UO_315 (O_315,N_29133,N_28577);
nor UO_316 (O_316,N_29925,N_29203);
nor UO_317 (O_317,N_29056,N_29662);
nor UO_318 (O_318,N_28655,N_29128);
xor UO_319 (O_319,N_29667,N_28848);
and UO_320 (O_320,N_29366,N_29788);
xnor UO_321 (O_321,N_29453,N_29669);
or UO_322 (O_322,N_29655,N_29523);
or UO_323 (O_323,N_28594,N_29015);
or UO_324 (O_324,N_28743,N_29588);
nand UO_325 (O_325,N_28920,N_29660);
xor UO_326 (O_326,N_28686,N_29225);
or UO_327 (O_327,N_29447,N_29057);
or UO_328 (O_328,N_29277,N_29988);
nand UO_329 (O_329,N_28707,N_28832);
nand UO_330 (O_330,N_29722,N_29595);
xnor UO_331 (O_331,N_29248,N_29946);
nand UO_332 (O_332,N_29292,N_29325);
nand UO_333 (O_333,N_29202,N_28507);
nand UO_334 (O_334,N_29712,N_29191);
xnor UO_335 (O_335,N_28588,N_29428);
and UO_336 (O_336,N_28880,N_29762);
nor UO_337 (O_337,N_29356,N_29261);
or UO_338 (O_338,N_28529,N_29681);
nor UO_339 (O_339,N_28800,N_29805);
and UO_340 (O_340,N_29578,N_29163);
nand UO_341 (O_341,N_29420,N_28991);
or UO_342 (O_342,N_29555,N_29801);
or UO_343 (O_343,N_28616,N_28934);
and UO_344 (O_344,N_29101,N_29214);
or UO_345 (O_345,N_28773,N_28780);
and UO_346 (O_346,N_28583,N_29460);
xor UO_347 (O_347,N_29668,N_29328);
nor UO_348 (O_348,N_29904,N_29716);
nor UO_349 (O_349,N_28865,N_29897);
nor UO_350 (O_350,N_29910,N_29989);
or UO_351 (O_351,N_28597,N_29930);
nor UO_352 (O_352,N_28516,N_29083);
or UO_353 (O_353,N_29746,N_29224);
and UO_354 (O_354,N_29554,N_29107);
and UO_355 (O_355,N_29540,N_29832);
nand UO_356 (O_356,N_29979,N_29470);
nand UO_357 (O_357,N_29587,N_29086);
nand UO_358 (O_358,N_29650,N_29259);
or UO_359 (O_359,N_28679,N_29103);
or UO_360 (O_360,N_29410,N_29906);
or UO_361 (O_361,N_28652,N_28512);
nand UO_362 (O_362,N_29290,N_29856);
nand UO_363 (O_363,N_29448,N_29609);
nor UO_364 (O_364,N_28735,N_29504);
and UO_365 (O_365,N_28851,N_28913);
nor UO_366 (O_366,N_29860,N_28950);
and UO_367 (O_367,N_29227,N_28744);
xnor UO_368 (O_368,N_28959,N_29396);
nor UO_369 (O_369,N_29706,N_29023);
and UO_370 (O_370,N_29373,N_29135);
nand UO_371 (O_371,N_29298,N_28893);
nor UO_372 (O_372,N_29508,N_28522);
xnor UO_373 (O_373,N_28837,N_28839);
xor UO_374 (O_374,N_29657,N_29542);
nor UO_375 (O_375,N_29825,N_29709);
xor UO_376 (O_376,N_29475,N_29372);
xnor UO_377 (O_377,N_29685,N_28792);
and UO_378 (O_378,N_28625,N_29627);
nand UO_379 (O_379,N_29231,N_29182);
nor UO_380 (O_380,N_29537,N_29664);
or UO_381 (O_381,N_28905,N_29349);
and UO_382 (O_382,N_28994,N_29286);
xnor UO_383 (O_383,N_29005,N_28628);
xnor UO_384 (O_384,N_28649,N_28642);
or UO_385 (O_385,N_29501,N_28609);
nor UO_386 (O_386,N_29238,N_29799);
xor UO_387 (O_387,N_29213,N_29285);
nor UO_388 (O_388,N_28591,N_29110);
or UO_389 (O_389,N_29434,N_29790);
or UO_390 (O_390,N_29921,N_29845);
and UO_391 (O_391,N_29192,N_28627);
nand UO_392 (O_392,N_29081,N_28682);
nand UO_393 (O_393,N_29947,N_28504);
xnor UO_394 (O_394,N_28704,N_29270);
xnor UO_395 (O_395,N_28542,N_29855);
and UO_396 (O_396,N_28527,N_28526);
xor UO_397 (O_397,N_29446,N_28556);
and UO_398 (O_398,N_28914,N_29651);
and UO_399 (O_399,N_29495,N_29412);
xor UO_400 (O_400,N_29743,N_29816);
xnor UO_401 (O_401,N_29923,N_28801);
or UO_402 (O_402,N_28779,N_28753);
nor UO_403 (O_403,N_29346,N_28684);
or UO_404 (O_404,N_28724,N_29901);
and UO_405 (O_405,N_29071,N_29811);
or UO_406 (O_406,N_29917,N_29894);
nor UO_407 (O_407,N_28983,N_29179);
or UO_408 (O_408,N_29938,N_29462);
xor UO_409 (O_409,N_29849,N_29739);
xnor UO_410 (O_410,N_29084,N_29104);
xor UO_411 (O_411,N_28987,N_29532);
nand UO_412 (O_412,N_29605,N_29984);
nand UO_413 (O_413,N_29177,N_29250);
or UO_414 (O_414,N_29199,N_29350);
xnor UO_415 (O_415,N_29047,N_29594);
xor UO_416 (O_416,N_29241,N_29054);
or UO_417 (O_417,N_29781,N_28549);
nand UO_418 (O_418,N_29266,N_29730);
xnor UO_419 (O_419,N_28639,N_28917);
and UO_420 (O_420,N_29877,N_29718);
nand UO_421 (O_421,N_29132,N_29332);
or UO_422 (O_422,N_29912,N_29500);
xor UO_423 (O_423,N_29851,N_28736);
nor UO_424 (O_424,N_28756,N_29665);
or UO_425 (O_425,N_28926,N_28740);
and UO_426 (O_426,N_29121,N_29272);
and UO_427 (O_427,N_29995,N_28907);
nor UO_428 (O_428,N_29406,N_28857);
and UO_429 (O_429,N_29176,N_29108);
nand UO_430 (O_430,N_29807,N_28889);
or UO_431 (O_431,N_29950,N_29112);
xnor UO_432 (O_432,N_28964,N_29145);
nor UO_433 (O_433,N_28791,N_29079);
xor UO_434 (O_434,N_29632,N_29247);
nor UO_435 (O_435,N_29046,N_29000);
and UO_436 (O_436,N_29335,N_29010);
and UO_437 (O_437,N_28614,N_29809);
nor UO_438 (O_438,N_29707,N_29887);
xor UO_439 (O_439,N_29150,N_29094);
xnor UO_440 (O_440,N_29545,N_29874);
nor UO_441 (O_441,N_28993,N_28696);
or UO_442 (O_442,N_28607,N_28988);
and UO_443 (O_443,N_28766,N_29068);
nand UO_444 (O_444,N_28794,N_28508);
nand UO_445 (O_445,N_29754,N_29782);
nor UO_446 (O_446,N_29435,N_28884);
xnor UO_447 (O_447,N_29151,N_29926);
or UO_448 (O_448,N_28667,N_29876);
nand UO_449 (O_449,N_28675,N_28569);
nand UO_450 (O_450,N_29793,N_28828);
nor UO_451 (O_451,N_29439,N_29329);
nor UO_452 (O_452,N_28661,N_29275);
nor UO_453 (O_453,N_29333,N_29378);
and UO_454 (O_454,N_29551,N_29779);
nor UO_455 (O_455,N_29638,N_29204);
nand UO_456 (O_456,N_29172,N_28980);
and UO_457 (O_457,N_29941,N_28737);
or UO_458 (O_458,N_29738,N_28781);
xnor UO_459 (O_459,N_29720,N_28817);
xnor UO_460 (O_460,N_28633,N_29147);
and UO_461 (O_461,N_29355,N_28519);
or UO_462 (O_462,N_29080,N_28835);
nand UO_463 (O_463,N_29067,N_28587);
nand UO_464 (O_464,N_29829,N_28671);
and UO_465 (O_465,N_29488,N_29631);
or UO_466 (O_466,N_28580,N_29843);
nand UO_467 (O_467,N_28677,N_29553);
or UO_468 (O_468,N_29365,N_28717);
xnor UO_469 (O_469,N_28598,N_28982);
and UO_470 (O_470,N_29398,N_29842);
nand UO_471 (O_471,N_29237,N_28581);
or UO_472 (O_472,N_28539,N_29431);
xnor UO_473 (O_473,N_29526,N_29616);
or UO_474 (O_474,N_29747,N_29070);
nor UO_475 (O_475,N_29774,N_28908);
nand UO_476 (O_476,N_29680,N_29330);
nand UO_477 (O_477,N_29119,N_28930);
or UO_478 (O_478,N_29732,N_29886);
or UO_479 (O_479,N_29013,N_29363);
nand UO_480 (O_480,N_29209,N_28894);
xor UO_481 (O_481,N_29986,N_29388);
nand UO_482 (O_482,N_28599,N_29574);
or UO_483 (O_483,N_28755,N_28909);
xor UO_484 (O_484,N_29696,N_29063);
or UO_485 (O_485,N_28613,N_29890);
and UO_486 (O_486,N_29242,N_29474);
nor UO_487 (O_487,N_29082,N_28901);
and UO_488 (O_488,N_29525,N_29161);
and UO_489 (O_489,N_29490,N_29824);
xnor UO_490 (O_490,N_29403,N_29908);
nand UO_491 (O_491,N_29092,N_29123);
or UO_492 (O_492,N_29391,N_29992);
and UO_493 (O_493,N_29234,N_29143);
or UO_494 (O_494,N_29251,N_29957);
xnor UO_495 (O_495,N_28941,N_28869);
or UO_496 (O_496,N_28797,N_29536);
xnor UO_497 (O_497,N_29652,N_28546);
nor UO_498 (O_498,N_28876,N_28561);
nor UO_499 (O_499,N_28506,N_29924);
or UO_500 (O_500,N_28664,N_28925);
nor UO_501 (O_501,N_28646,N_28998);
or UO_502 (O_502,N_29433,N_29228);
or UO_503 (O_503,N_29658,N_29457);
nand UO_504 (O_504,N_28582,N_29385);
or UO_505 (O_505,N_29018,N_29647);
nand UO_506 (O_506,N_28819,N_29461);
or UO_507 (O_507,N_29183,N_29663);
or UO_508 (O_508,N_28566,N_29571);
or UO_509 (O_509,N_28812,N_29324);
or UO_510 (O_510,N_29370,N_28571);
or UO_511 (O_511,N_28963,N_29233);
nand UO_512 (O_512,N_28870,N_29341);
xor UO_513 (O_513,N_29060,N_29982);
or UO_514 (O_514,N_28711,N_29282);
nand UO_515 (O_515,N_28824,N_29878);
and UO_516 (O_516,N_28706,N_28796);
or UO_517 (O_517,N_29389,N_28701);
nand UO_518 (O_518,N_28500,N_28978);
and UO_519 (O_519,N_28681,N_29538);
or UO_520 (O_520,N_29572,N_29624);
xnor UO_521 (O_521,N_29397,N_29352);
nand UO_522 (O_522,N_29451,N_29772);
nor UO_523 (O_523,N_29522,N_29371);
and UO_524 (O_524,N_29625,N_29800);
and UO_525 (O_525,N_29443,N_29823);
nand UO_526 (O_526,N_29264,N_29265);
or UO_527 (O_527,N_28703,N_29099);
nor UO_528 (O_528,N_28503,N_29954);
nor UO_529 (O_529,N_28647,N_28533);
or UO_530 (O_530,N_29922,N_28721);
or UO_531 (O_531,N_29052,N_28518);
xor UO_532 (O_532,N_29687,N_29733);
or UO_533 (O_533,N_28510,N_29547);
nor UO_534 (O_534,N_29156,N_28700);
and UO_535 (O_535,N_29895,N_29531);
or UO_536 (O_536,N_29838,N_29656);
xnor UO_537 (O_537,N_29076,N_29672);
or UO_538 (O_538,N_28689,N_29154);
or UO_539 (O_539,N_29670,N_29315);
xor UO_540 (O_540,N_29646,N_29339);
and UO_541 (O_541,N_29990,N_28666);
and UO_542 (O_542,N_28912,N_28952);
or UO_543 (O_543,N_28733,N_29980);
or UO_544 (O_544,N_29534,N_28776);
or UO_545 (O_545,N_29267,N_28986);
or UO_546 (O_546,N_28731,N_29287);
nand UO_547 (O_547,N_29944,N_29902);
or UO_548 (O_548,N_28593,N_29763);
nand UO_549 (O_549,N_29184,N_29168);
and UO_550 (O_550,N_28572,N_29654);
or UO_551 (O_551,N_29394,N_29042);
nor UO_552 (O_552,N_29155,N_28818);
or UO_553 (O_553,N_28654,N_29276);
or UO_554 (O_554,N_28532,N_28674);
and UO_555 (O_555,N_28502,N_28821);
nand UO_556 (O_556,N_29049,N_29491);
and UO_557 (O_557,N_29544,N_29380);
nor UO_558 (O_558,N_29111,N_29053);
and UO_559 (O_559,N_28612,N_28557);
nor UO_560 (O_560,N_29852,N_28651);
or UO_561 (O_561,N_28972,N_28730);
and UO_562 (O_562,N_29483,N_29481);
and UO_563 (O_563,N_29643,N_28718);
or UO_564 (O_564,N_28680,N_28759);
xor UO_565 (O_565,N_29144,N_29819);
xnor UO_566 (O_566,N_29686,N_28545);
nor UO_567 (O_567,N_29253,N_29755);
nor UO_568 (O_568,N_28895,N_29257);
and UO_569 (O_569,N_29486,N_29606);
and UO_570 (O_570,N_28568,N_28672);
nand UO_571 (O_571,N_29438,N_29993);
nor UO_572 (O_572,N_29066,N_29304);
or UO_573 (O_573,N_29705,N_28713);
xnor UO_574 (O_574,N_29338,N_29293);
or UO_575 (O_575,N_29870,N_29559);
nor UO_576 (O_576,N_28836,N_29937);
and UO_577 (O_577,N_28874,N_28739);
or UO_578 (O_578,N_29493,N_28888);
nor UO_579 (O_579,N_28867,N_28501);
or UO_580 (O_580,N_29240,N_28668);
nand UO_581 (O_581,N_29043,N_28969);
nor UO_582 (O_582,N_29566,N_29745);
nor UO_583 (O_583,N_29468,N_29953);
or UO_584 (O_584,N_29246,N_29822);
nand UO_585 (O_585,N_28927,N_28937);
or UO_586 (O_586,N_28548,N_29273);
nor UO_587 (O_587,N_28698,N_29775);
or UO_588 (O_588,N_29496,N_29050);
nand UO_589 (O_589,N_29096,N_29831);
nor UO_590 (O_590,N_29062,N_29607);
nor UO_591 (O_591,N_29563,N_29205);
nor UO_592 (O_592,N_28973,N_29090);
xor UO_593 (O_593,N_29621,N_29484);
nand UO_594 (O_594,N_29136,N_28615);
and UO_595 (O_595,N_29985,N_29786);
nor UO_596 (O_596,N_29517,N_29291);
xor UO_597 (O_597,N_28989,N_28843);
nor UO_598 (O_598,N_28979,N_29756);
nand UO_599 (O_599,N_29661,N_29883);
xnor UO_600 (O_600,N_29404,N_28769);
and UO_601 (O_601,N_29841,N_28810);
nand UO_602 (O_602,N_28685,N_28697);
or UO_603 (O_603,N_29244,N_28910);
nand UO_604 (O_604,N_29959,N_29727);
nor UO_605 (O_605,N_29387,N_29310);
nand UO_606 (O_606,N_28896,N_28585);
or UO_607 (O_607,N_28629,N_29949);
or UO_608 (O_608,N_28632,N_29505);
or UO_609 (O_609,N_29359,N_28558);
xor UO_610 (O_610,N_29520,N_29316);
and UO_611 (O_611,N_28543,N_28881);
xnor UO_612 (O_612,N_29249,N_29019);
and UO_613 (O_613,N_29884,N_29181);
or UO_614 (O_614,N_29564,N_29994);
nor UO_615 (O_615,N_29514,N_29318);
xnor UO_616 (O_616,N_28830,N_29217);
xnor UO_617 (O_617,N_28878,N_28751);
or UO_618 (O_618,N_28637,N_29865);
and UO_619 (O_619,N_29245,N_28631);
or UO_620 (O_620,N_29729,N_29592);
xor UO_621 (O_621,N_28938,N_29840);
xor UO_622 (O_622,N_29306,N_29761);
xnor UO_623 (O_623,N_29114,N_29760);
nor UO_624 (O_624,N_29375,N_29386);
and UO_625 (O_625,N_29674,N_29513);
nor UO_626 (O_626,N_29882,N_29452);
and UO_627 (O_627,N_29974,N_28855);
or UO_628 (O_628,N_29139,N_29167);
xor UO_629 (O_629,N_28694,N_29971);
nor UO_630 (O_630,N_29943,N_29477);
xnor UO_631 (O_631,N_28958,N_29708);
or UO_632 (O_632,N_29268,N_29868);
nor UO_633 (O_633,N_29173,N_28565);
or UO_634 (O_634,N_29603,N_29628);
nand UO_635 (O_635,N_28858,N_29317);
nor UO_636 (O_636,N_28960,N_29889);
xor UO_637 (O_637,N_28965,N_29846);
and UO_638 (O_638,N_28747,N_29029);
nand UO_639 (O_639,N_29269,N_29958);
and UO_640 (O_640,N_28760,N_29336);
xor UO_641 (O_641,N_29113,N_28547);
nand UO_642 (O_642,N_28702,N_29279);
xnor UO_643 (O_643,N_28523,N_29465);
nor UO_644 (O_644,N_28854,N_29487);
or UO_645 (O_645,N_28775,N_28803);
xnor UO_646 (O_646,N_29837,N_29875);
xnor UO_647 (O_647,N_28579,N_28942);
nand UO_648 (O_648,N_29833,N_28806);
or UO_649 (O_649,N_28975,N_29368);
xor UO_650 (O_650,N_29640,N_28961);
or UO_651 (O_651,N_29703,N_28886);
or UO_652 (O_652,N_29600,N_29556);
nor UO_653 (O_653,N_28643,N_29165);
or UO_654 (O_654,N_29963,N_29726);
nor UO_655 (O_655,N_29645,N_29962);
xnor UO_656 (O_656,N_29467,N_28825);
nor UO_657 (O_657,N_29585,N_28719);
and UO_658 (O_658,N_29864,N_29232);
nor UO_659 (O_659,N_28550,N_29303);
xnor UO_660 (O_660,N_29596,N_28949);
or UO_661 (O_661,N_29507,N_29064);
and UO_662 (O_662,N_29552,N_28617);
or UO_663 (O_663,N_29827,N_29509);
nor UO_664 (O_664,N_29942,N_28892);
and UO_665 (O_665,N_29817,N_29735);
nand UO_666 (O_666,N_28573,N_29400);
xor UO_667 (O_667,N_29582,N_29497);
or UO_668 (O_668,N_29783,N_29767);
nor UO_669 (O_669,N_29402,N_28690);
nand UO_670 (O_670,N_29951,N_28954);
nand UO_671 (O_671,N_29122,N_29390);
nand UO_672 (O_672,N_29765,N_28636);
and UO_673 (O_673,N_29713,N_29599);
nand UO_674 (O_674,N_28734,N_29376);
nand UO_675 (O_675,N_28640,N_29618);
or UO_676 (O_676,N_29913,N_29787);
nand UO_677 (O_677,N_28933,N_28831);
nor UO_678 (O_678,N_29162,N_28997);
or UO_679 (O_679,N_29835,N_28990);
and UO_680 (O_680,N_29972,N_29185);
and UO_681 (O_681,N_28560,N_29194);
xor UO_682 (O_682,N_29975,N_28767);
or UO_683 (O_683,N_29789,N_28852);
or UO_684 (O_684,N_28761,N_29263);
xnor UO_685 (O_685,N_28786,N_28799);
nor UO_686 (O_686,N_29952,N_29180);
or UO_687 (O_687,N_29880,N_29188);
xor UO_688 (O_688,N_28660,N_29226);
and UO_689 (O_689,N_29998,N_29017);
or UO_690 (O_690,N_28738,N_29516);
nor UO_691 (O_691,N_28669,N_29753);
nor UO_692 (O_692,N_28981,N_29914);
nor UO_693 (O_693,N_28838,N_29190);
nand UO_694 (O_694,N_29711,N_28553);
xor UO_695 (O_695,N_28928,N_28705);
or UO_696 (O_696,N_29208,N_29383);
and UO_697 (O_697,N_29633,N_29511);
xnor UO_698 (O_698,N_28514,N_28948);
nand UO_699 (O_699,N_28554,N_29415);
or UO_700 (O_700,N_29702,N_29622);
and UO_701 (O_701,N_28946,N_29529);
nand UO_702 (O_702,N_28611,N_28695);
nor UO_703 (O_703,N_28586,N_29106);
and UO_704 (O_704,N_29284,N_29077);
or UO_705 (O_705,N_29102,N_29543);
xnor UO_706 (O_706,N_29473,N_29796);
nand UO_707 (O_707,N_29945,N_28541);
or UO_708 (O_708,N_28650,N_29097);
nand UO_709 (O_709,N_29899,N_28530);
nor UO_710 (O_710,N_29069,N_29037);
and UO_711 (O_711,N_29991,N_29931);
xnor UO_712 (O_712,N_29271,N_29736);
and UO_713 (O_713,N_29393,N_28621);
xnor UO_714 (O_714,N_29844,N_29426);
xnor UO_715 (O_715,N_29748,N_29430);
nor UO_716 (O_716,N_28723,N_29872);
nor UO_717 (O_717,N_29675,N_29987);
nand UO_718 (O_718,N_29219,N_29839);
xor UO_719 (O_719,N_28890,N_29903);
nand UO_720 (O_720,N_28904,N_28728);
and UO_721 (O_721,N_29850,N_29967);
nor UO_722 (O_722,N_28992,N_29734);
xor UO_723 (O_723,N_28789,N_29326);
nand UO_724 (O_724,N_28563,N_28795);
and UO_725 (O_725,N_29524,N_29879);
nor UO_726 (O_726,N_28720,N_29752);
and UO_727 (O_727,N_28962,N_29478);
nor UO_728 (O_728,N_29032,N_29928);
nor UO_729 (O_729,N_28624,N_29927);
or UO_730 (O_730,N_29347,N_28872);
and UO_731 (O_731,N_29695,N_29634);
nor UO_732 (O_732,N_29411,N_29590);
and UO_733 (O_733,N_29274,N_29294);
and UO_734 (O_734,N_29932,N_29187);
and UO_735 (O_735,N_29608,N_29610);
xor UO_736 (O_736,N_29626,N_28729);
nand UO_737 (O_737,N_29848,N_28524);
nand UO_738 (O_738,N_28638,N_29826);
or UO_739 (O_739,N_28564,N_28644);
and UO_740 (O_740,N_29785,N_28966);
or UO_741 (O_741,N_29399,N_28882);
nand UO_742 (O_742,N_29311,N_29065);
xor UO_743 (O_743,N_28584,N_29489);
and UO_744 (O_744,N_29223,N_29892);
nand UO_745 (O_745,N_28885,N_29152);
and UO_746 (O_746,N_29369,N_29016);
nor UO_747 (O_747,N_29676,N_29704);
nor UO_748 (O_748,N_29169,N_28630);
xor UO_749 (O_749,N_28676,N_29222);
nor UO_750 (O_750,N_28877,N_28583);
and UO_751 (O_751,N_29926,N_29930);
and UO_752 (O_752,N_28861,N_29975);
or UO_753 (O_753,N_29099,N_29341);
and UO_754 (O_754,N_29587,N_29164);
or UO_755 (O_755,N_28721,N_29325);
nor UO_756 (O_756,N_29985,N_29288);
and UO_757 (O_757,N_28536,N_28715);
nor UO_758 (O_758,N_29585,N_29068);
and UO_759 (O_759,N_29272,N_29316);
nor UO_760 (O_760,N_29224,N_29813);
xor UO_761 (O_761,N_29261,N_29917);
nand UO_762 (O_762,N_29768,N_29880);
nand UO_763 (O_763,N_29318,N_29126);
nor UO_764 (O_764,N_28726,N_28504);
or UO_765 (O_765,N_29108,N_28673);
nor UO_766 (O_766,N_29908,N_28575);
or UO_767 (O_767,N_28841,N_28710);
nor UO_768 (O_768,N_29799,N_29948);
and UO_769 (O_769,N_29025,N_29829);
xnor UO_770 (O_770,N_29979,N_28831);
and UO_771 (O_771,N_29468,N_29485);
nor UO_772 (O_772,N_28579,N_29279);
xnor UO_773 (O_773,N_28907,N_28979);
nand UO_774 (O_774,N_29273,N_29675);
nand UO_775 (O_775,N_29212,N_29855);
and UO_776 (O_776,N_29513,N_29888);
nor UO_777 (O_777,N_29311,N_28696);
nand UO_778 (O_778,N_29079,N_28672);
nand UO_779 (O_779,N_28646,N_29381);
nor UO_780 (O_780,N_29850,N_29844);
nor UO_781 (O_781,N_29934,N_29585);
and UO_782 (O_782,N_29702,N_28931);
and UO_783 (O_783,N_29972,N_29117);
and UO_784 (O_784,N_29654,N_28838);
xor UO_785 (O_785,N_29359,N_29631);
or UO_786 (O_786,N_28955,N_29722);
and UO_787 (O_787,N_29027,N_29469);
and UO_788 (O_788,N_28872,N_29885);
xnor UO_789 (O_789,N_29906,N_29046);
and UO_790 (O_790,N_28694,N_29435);
or UO_791 (O_791,N_28898,N_29948);
or UO_792 (O_792,N_29218,N_28555);
xor UO_793 (O_793,N_29001,N_29095);
nand UO_794 (O_794,N_29554,N_29796);
nor UO_795 (O_795,N_29475,N_29495);
and UO_796 (O_796,N_29166,N_28984);
nor UO_797 (O_797,N_29014,N_28535);
xor UO_798 (O_798,N_29270,N_29650);
and UO_799 (O_799,N_29618,N_28876);
xor UO_800 (O_800,N_29369,N_28646);
nand UO_801 (O_801,N_28923,N_29477);
nand UO_802 (O_802,N_29796,N_29835);
or UO_803 (O_803,N_29952,N_28827);
and UO_804 (O_804,N_29206,N_28839);
or UO_805 (O_805,N_28766,N_29643);
or UO_806 (O_806,N_28860,N_29613);
and UO_807 (O_807,N_29970,N_29082);
nor UO_808 (O_808,N_29571,N_29849);
and UO_809 (O_809,N_29172,N_29704);
nor UO_810 (O_810,N_29310,N_29225);
and UO_811 (O_811,N_29277,N_28536);
or UO_812 (O_812,N_29876,N_29503);
nor UO_813 (O_813,N_29097,N_28639);
and UO_814 (O_814,N_28893,N_28591);
nand UO_815 (O_815,N_29869,N_29029);
nand UO_816 (O_816,N_29957,N_29557);
nand UO_817 (O_817,N_29141,N_29888);
xnor UO_818 (O_818,N_29586,N_29433);
nand UO_819 (O_819,N_28944,N_29771);
or UO_820 (O_820,N_28577,N_28685);
nand UO_821 (O_821,N_29146,N_29193);
nand UO_822 (O_822,N_29071,N_28720);
nor UO_823 (O_823,N_28874,N_29298);
nor UO_824 (O_824,N_29358,N_29009);
nor UO_825 (O_825,N_28774,N_28972);
nand UO_826 (O_826,N_29993,N_28606);
nand UO_827 (O_827,N_29835,N_29343);
and UO_828 (O_828,N_29295,N_28817);
nand UO_829 (O_829,N_28781,N_28909);
xor UO_830 (O_830,N_29912,N_29136);
nor UO_831 (O_831,N_29295,N_29640);
nand UO_832 (O_832,N_29048,N_29705);
nand UO_833 (O_833,N_29481,N_29812);
or UO_834 (O_834,N_28646,N_29038);
nor UO_835 (O_835,N_28563,N_28732);
nor UO_836 (O_836,N_29719,N_28527);
nor UO_837 (O_837,N_29735,N_29698);
nand UO_838 (O_838,N_29930,N_29304);
and UO_839 (O_839,N_29374,N_29590);
or UO_840 (O_840,N_29504,N_29036);
and UO_841 (O_841,N_29010,N_29154);
and UO_842 (O_842,N_29542,N_29367);
nand UO_843 (O_843,N_28688,N_29747);
and UO_844 (O_844,N_28543,N_29318);
nand UO_845 (O_845,N_28546,N_29742);
nor UO_846 (O_846,N_28679,N_29261);
and UO_847 (O_847,N_28769,N_29688);
nand UO_848 (O_848,N_29918,N_29313);
and UO_849 (O_849,N_29724,N_29209);
xnor UO_850 (O_850,N_29173,N_29065);
xnor UO_851 (O_851,N_29973,N_29909);
or UO_852 (O_852,N_29956,N_29543);
and UO_853 (O_853,N_29450,N_29948);
nand UO_854 (O_854,N_29118,N_28814);
xor UO_855 (O_855,N_28676,N_29214);
and UO_856 (O_856,N_29552,N_29845);
nand UO_857 (O_857,N_28705,N_29520);
and UO_858 (O_858,N_29467,N_29952);
nand UO_859 (O_859,N_29618,N_28678);
nand UO_860 (O_860,N_28999,N_29933);
nand UO_861 (O_861,N_29463,N_29823);
and UO_862 (O_862,N_28860,N_29702);
xor UO_863 (O_863,N_28748,N_29566);
nor UO_864 (O_864,N_29500,N_28839);
nor UO_865 (O_865,N_29968,N_28603);
and UO_866 (O_866,N_29295,N_28612);
xnor UO_867 (O_867,N_29288,N_29757);
or UO_868 (O_868,N_29339,N_29075);
nor UO_869 (O_869,N_29344,N_28695);
nand UO_870 (O_870,N_29255,N_29119);
and UO_871 (O_871,N_28575,N_28903);
or UO_872 (O_872,N_29088,N_29129);
or UO_873 (O_873,N_29799,N_29291);
and UO_874 (O_874,N_29659,N_29706);
or UO_875 (O_875,N_29103,N_28734);
or UO_876 (O_876,N_28811,N_29806);
nand UO_877 (O_877,N_28792,N_29042);
xnor UO_878 (O_878,N_29455,N_28948);
nor UO_879 (O_879,N_29190,N_28890);
nor UO_880 (O_880,N_29679,N_29358);
nand UO_881 (O_881,N_29871,N_28963);
and UO_882 (O_882,N_29910,N_28855);
nand UO_883 (O_883,N_29445,N_28592);
nand UO_884 (O_884,N_29469,N_29096);
nor UO_885 (O_885,N_29084,N_29231);
and UO_886 (O_886,N_29891,N_28814);
nor UO_887 (O_887,N_29056,N_28794);
xor UO_888 (O_888,N_29809,N_28554);
nand UO_889 (O_889,N_29643,N_29529);
nand UO_890 (O_890,N_29550,N_29502);
nand UO_891 (O_891,N_29055,N_29565);
and UO_892 (O_892,N_29909,N_29360);
and UO_893 (O_893,N_28732,N_28875);
xnor UO_894 (O_894,N_29821,N_29675);
or UO_895 (O_895,N_29314,N_29302);
and UO_896 (O_896,N_29415,N_28958);
nand UO_897 (O_897,N_29881,N_29163);
and UO_898 (O_898,N_29770,N_29060);
or UO_899 (O_899,N_29804,N_29182);
and UO_900 (O_900,N_28945,N_29515);
nand UO_901 (O_901,N_29949,N_28796);
or UO_902 (O_902,N_29274,N_29907);
xnor UO_903 (O_903,N_29775,N_29846);
nor UO_904 (O_904,N_29006,N_29118);
nand UO_905 (O_905,N_29188,N_29995);
nor UO_906 (O_906,N_28926,N_28563);
or UO_907 (O_907,N_29916,N_29863);
nand UO_908 (O_908,N_28729,N_29095);
xnor UO_909 (O_909,N_29711,N_28688);
or UO_910 (O_910,N_29139,N_28692);
xor UO_911 (O_911,N_28810,N_29365);
or UO_912 (O_912,N_29085,N_29464);
nand UO_913 (O_913,N_29553,N_29510);
xor UO_914 (O_914,N_28637,N_29783);
nand UO_915 (O_915,N_29883,N_29040);
or UO_916 (O_916,N_29451,N_29917);
nor UO_917 (O_917,N_28801,N_28951);
nor UO_918 (O_918,N_29127,N_28697);
xor UO_919 (O_919,N_29247,N_29284);
nand UO_920 (O_920,N_29130,N_28684);
xor UO_921 (O_921,N_28656,N_29591);
and UO_922 (O_922,N_29357,N_29267);
nor UO_923 (O_923,N_29808,N_29570);
nor UO_924 (O_924,N_29955,N_28545);
or UO_925 (O_925,N_29142,N_28975);
nor UO_926 (O_926,N_29950,N_28995);
nor UO_927 (O_927,N_29973,N_29994);
nor UO_928 (O_928,N_29298,N_28616);
or UO_929 (O_929,N_28800,N_28681);
nor UO_930 (O_930,N_28919,N_29660);
and UO_931 (O_931,N_29443,N_29915);
nor UO_932 (O_932,N_29032,N_28554);
nand UO_933 (O_933,N_29083,N_29273);
or UO_934 (O_934,N_29864,N_28945);
xor UO_935 (O_935,N_29958,N_29432);
nor UO_936 (O_936,N_29800,N_29114);
nand UO_937 (O_937,N_29276,N_29238);
nand UO_938 (O_938,N_29513,N_28775);
nand UO_939 (O_939,N_28746,N_29691);
nand UO_940 (O_940,N_29354,N_29898);
nor UO_941 (O_941,N_29214,N_28771);
nand UO_942 (O_942,N_29717,N_29194);
and UO_943 (O_943,N_29003,N_29716);
or UO_944 (O_944,N_29795,N_28504);
and UO_945 (O_945,N_29758,N_29145);
nand UO_946 (O_946,N_29210,N_29111);
xnor UO_947 (O_947,N_28672,N_28730);
nor UO_948 (O_948,N_29043,N_28608);
nand UO_949 (O_949,N_28858,N_29583);
xnor UO_950 (O_950,N_29495,N_29648);
and UO_951 (O_951,N_28829,N_28915);
xor UO_952 (O_952,N_29986,N_29114);
nor UO_953 (O_953,N_29924,N_29998);
and UO_954 (O_954,N_28732,N_28958);
or UO_955 (O_955,N_29383,N_29518);
or UO_956 (O_956,N_29151,N_28552);
xor UO_957 (O_957,N_28689,N_29776);
nor UO_958 (O_958,N_28948,N_28570);
or UO_959 (O_959,N_28859,N_28745);
or UO_960 (O_960,N_29246,N_28703);
nor UO_961 (O_961,N_28634,N_28829);
nor UO_962 (O_962,N_29285,N_29602);
and UO_963 (O_963,N_29482,N_29142);
nand UO_964 (O_964,N_29475,N_29904);
xor UO_965 (O_965,N_29856,N_29755);
or UO_966 (O_966,N_28740,N_29388);
and UO_967 (O_967,N_29745,N_29192);
nor UO_968 (O_968,N_29511,N_29120);
nor UO_969 (O_969,N_29239,N_29192);
or UO_970 (O_970,N_29696,N_29020);
or UO_971 (O_971,N_28774,N_29680);
xnor UO_972 (O_972,N_29458,N_28910);
xor UO_973 (O_973,N_29121,N_29096);
nor UO_974 (O_974,N_28960,N_28809);
or UO_975 (O_975,N_29255,N_29072);
nor UO_976 (O_976,N_29866,N_29590);
and UO_977 (O_977,N_29511,N_28589);
xnor UO_978 (O_978,N_29448,N_28887);
nor UO_979 (O_979,N_29618,N_28722);
or UO_980 (O_980,N_29033,N_29911);
nor UO_981 (O_981,N_29941,N_29870);
nand UO_982 (O_982,N_28617,N_29974);
nand UO_983 (O_983,N_28704,N_28751);
nand UO_984 (O_984,N_29948,N_28651);
nor UO_985 (O_985,N_29892,N_28731);
nor UO_986 (O_986,N_29945,N_28597);
xor UO_987 (O_987,N_29756,N_29740);
and UO_988 (O_988,N_29251,N_29693);
or UO_989 (O_989,N_28848,N_29268);
and UO_990 (O_990,N_29278,N_29272);
and UO_991 (O_991,N_28782,N_29295);
xnor UO_992 (O_992,N_28503,N_29568);
and UO_993 (O_993,N_29860,N_29225);
nor UO_994 (O_994,N_29030,N_28521);
xnor UO_995 (O_995,N_28858,N_29148);
or UO_996 (O_996,N_28671,N_28681);
xnor UO_997 (O_997,N_29265,N_29723);
xnor UO_998 (O_998,N_29537,N_29145);
nor UO_999 (O_999,N_29724,N_29328);
nand UO_1000 (O_1000,N_29989,N_28992);
nand UO_1001 (O_1001,N_29485,N_29743);
xor UO_1002 (O_1002,N_29249,N_28810);
nor UO_1003 (O_1003,N_29080,N_29092);
and UO_1004 (O_1004,N_28852,N_29161);
nand UO_1005 (O_1005,N_29396,N_28639);
nand UO_1006 (O_1006,N_29587,N_29751);
and UO_1007 (O_1007,N_29066,N_28715);
nand UO_1008 (O_1008,N_28831,N_29804);
xnor UO_1009 (O_1009,N_29564,N_29053);
nand UO_1010 (O_1010,N_29018,N_29381);
and UO_1011 (O_1011,N_29139,N_29928);
nand UO_1012 (O_1012,N_29598,N_29127);
and UO_1013 (O_1013,N_29977,N_29144);
and UO_1014 (O_1014,N_29637,N_29434);
nor UO_1015 (O_1015,N_29382,N_29915);
nor UO_1016 (O_1016,N_28783,N_29206);
xnor UO_1017 (O_1017,N_28708,N_29046);
or UO_1018 (O_1018,N_29280,N_29554);
nor UO_1019 (O_1019,N_29003,N_28516);
xor UO_1020 (O_1020,N_29714,N_28725);
nor UO_1021 (O_1021,N_29198,N_29967);
xor UO_1022 (O_1022,N_28561,N_29646);
nor UO_1023 (O_1023,N_29287,N_29397);
xor UO_1024 (O_1024,N_29671,N_29440);
and UO_1025 (O_1025,N_28892,N_29802);
or UO_1026 (O_1026,N_29204,N_29186);
and UO_1027 (O_1027,N_28872,N_29795);
nand UO_1028 (O_1028,N_29693,N_28961);
and UO_1029 (O_1029,N_28732,N_28821);
xor UO_1030 (O_1030,N_29975,N_29139);
and UO_1031 (O_1031,N_28963,N_29726);
or UO_1032 (O_1032,N_28672,N_29295);
or UO_1033 (O_1033,N_29877,N_29970);
nand UO_1034 (O_1034,N_28642,N_29887);
xnor UO_1035 (O_1035,N_29400,N_29382);
or UO_1036 (O_1036,N_29755,N_28678);
xor UO_1037 (O_1037,N_29615,N_29830);
nor UO_1038 (O_1038,N_29291,N_29682);
xnor UO_1039 (O_1039,N_28544,N_28795);
or UO_1040 (O_1040,N_28759,N_29081);
xnor UO_1041 (O_1041,N_28691,N_29066);
and UO_1042 (O_1042,N_29058,N_29707);
nand UO_1043 (O_1043,N_29091,N_28850);
or UO_1044 (O_1044,N_29219,N_29593);
nor UO_1045 (O_1045,N_29489,N_28982);
and UO_1046 (O_1046,N_28529,N_29272);
or UO_1047 (O_1047,N_29768,N_29521);
xor UO_1048 (O_1048,N_29904,N_29497);
nor UO_1049 (O_1049,N_28671,N_29353);
nand UO_1050 (O_1050,N_29057,N_29616);
nor UO_1051 (O_1051,N_29243,N_29026);
and UO_1052 (O_1052,N_29289,N_28683);
or UO_1053 (O_1053,N_29898,N_29840);
and UO_1054 (O_1054,N_29194,N_29078);
xnor UO_1055 (O_1055,N_28903,N_29568);
or UO_1056 (O_1056,N_29128,N_28712);
and UO_1057 (O_1057,N_29087,N_29427);
xor UO_1058 (O_1058,N_29009,N_29898);
xnor UO_1059 (O_1059,N_29586,N_29399);
and UO_1060 (O_1060,N_28849,N_29805);
nand UO_1061 (O_1061,N_28553,N_29898);
nor UO_1062 (O_1062,N_28984,N_29606);
and UO_1063 (O_1063,N_28970,N_28670);
nand UO_1064 (O_1064,N_29261,N_29882);
nor UO_1065 (O_1065,N_29613,N_29507);
nand UO_1066 (O_1066,N_29190,N_29949);
and UO_1067 (O_1067,N_28936,N_28531);
or UO_1068 (O_1068,N_29368,N_28861);
and UO_1069 (O_1069,N_29260,N_29563);
nand UO_1070 (O_1070,N_29403,N_29079);
or UO_1071 (O_1071,N_29314,N_28940);
or UO_1072 (O_1072,N_29693,N_28811);
and UO_1073 (O_1073,N_29548,N_28545);
and UO_1074 (O_1074,N_29963,N_29553);
and UO_1075 (O_1075,N_29854,N_28866);
nand UO_1076 (O_1076,N_29170,N_29629);
xnor UO_1077 (O_1077,N_29623,N_29149);
and UO_1078 (O_1078,N_29516,N_28526);
or UO_1079 (O_1079,N_28713,N_29892);
nor UO_1080 (O_1080,N_28550,N_29653);
nor UO_1081 (O_1081,N_29043,N_29288);
nand UO_1082 (O_1082,N_28752,N_28611);
nor UO_1083 (O_1083,N_28558,N_29643);
and UO_1084 (O_1084,N_29701,N_28617);
nand UO_1085 (O_1085,N_29179,N_29077);
nor UO_1086 (O_1086,N_28543,N_29043);
and UO_1087 (O_1087,N_28739,N_29200);
nor UO_1088 (O_1088,N_29741,N_29540);
and UO_1089 (O_1089,N_29641,N_29253);
nand UO_1090 (O_1090,N_28937,N_29922);
nor UO_1091 (O_1091,N_28985,N_29263);
and UO_1092 (O_1092,N_28669,N_29142);
nor UO_1093 (O_1093,N_29311,N_28892);
or UO_1094 (O_1094,N_28564,N_28723);
and UO_1095 (O_1095,N_28572,N_28869);
or UO_1096 (O_1096,N_29288,N_28977);
and UO_1097 (O_1097,N_29690,N_29914);
nor UO_1098 (O_1098,N_28771,N_29360);
xor UO_1099 (O_1099,N_28916,N_29738);
or UO_1100 (O_1100,N_29795,N_28969);
nor UO_1101 (O_1101,N_28716,N_28725);
nor UO_1102 (O_1102,N_29607,N_29369);
and UO_1103 (O_1103,N_28930,N_29092);
and UO_1104 (O_1104,N_28518,N_28840);
nor UO_1105 (O_1105,N_29291,N_29950);
nor UO_1106 (O_1106,N_29959,N_29806);
xnor UO_1107 (O_1107,N_29335,N_29563);
or UO_1108 (O_1108,N_28684,N_29823);
or UO_1109 (O_1109,N_29866,N_29941);
or UO_1110 (O_1110,N_28628,N_29859);
nand UO_1111 (O_1111,N_29088,N_29782);
or UO_1112 (O_1112,N_28646,N_28690);
nand UO_1113 (O_1113,N_29905,N_28938);
or UO_1114 (O_1114,N_29374,N_28832);
nor UO_1115 (O_1115,N_28799,N_29352);
or UO_1116 (O_1116,N_29085,N_28954);
nand UO_1117 (O_1117,N_28939,N_28631);
and UO_1118 (O_1118,N_29710,N_29258);
and UO_1119 (O_1119,N_29485,N_29875);
and UO_1120 (O_1120,N_28835,N_29304);
or UO_1121 (O_1121,N_29011,N_29492);
nand UO_1122 (O_1122,N_29495,N_29816);
xor UO_1123 (O_1123,N_29436,N_29551);
and UO_1124 (O_1124,N_29163,N_29461);
xnor UO_1125 (O_1125,N_28593,N_29534);
and UO_1126 (O_1126,N_29098,N_28995);
nand UO_1127 (O_1127,N_29377,N_28731);
or UO_1128 (O_1128,N_29791,N_29132);
and UO_1129 (O_1129,N_28806,N_29245);
or UO_1130 (O_1130,N_29059,N_29552);
or UO_1131 (O_1131,N_29390,N_28820);
and UO_1132 (O_1132,N_28779,N_28930);
nand UO_1133 (O_1133,N_29347,N_29002);
and UO_1134 (O_1134,N_29847,N_28560);
nor UO_1135 (O_1135,N_29250,N_29049);
nor UO_1136 (O_1136,N_28873,N_28932);
and UO_1137 (O_1137,N_29057,N_28627);
xor UO_1138 (O_1138,N_28625,N_29843);
nor UO_1139 (O_1139,N_28764,N_28547);
xnor UO_1140 (O_1140,N_29398,N_29570);
nor UO_1141 (O_1141,N_29572,N_29215);
nor UO_1142 (O_1142,N_29475,N_28988);
and UO_1143 (O_1143,N_29409,N_29986);
or UO_1144 (O_1144,N_29562,N_28684);
nor UO_1145 (O_1145,N_29733,N_28775);
xor UO_1146 (O_1146,N_29340,N_29653);
nand UO_1147 (O_1147,N_29318,N_28755);
nand UO_1148 (O_1148,N_28836,N_29559);
nand UO_1149 (O_1149,N_29841,N_29358);
or UO_1150 (O_1150,N_28882,N_29338);
nor UO_1151 (O_1151,N_29056,N_29176);
and UO_1152 (O_1152,N_29858,N_28566);
nor UO_1153 (O_1153,N_28704,N_29096);
or UO_1154 (O_1154,N_28544,N_29926);
or UO_1155 (O_1155,N_29689,N_29278);
nand UO_1156 (O_1156,N_28564,N_29114);
or UO_1157 (O_1157,N_28615,N_28852);
xor UO_1158 (O_1158,N_29847,N_29100);
nand UO_1159 (O_1159,N_28871,N_29308);
and UO_1160 (O_1160,N_29366,N_29666);
nor UO_1161 (O_1161,N_29444,N_29016);
and UO_1162 (O_1162,N_28832,N_28531);
and UO_1163 (O_1163,N_29069,N_28863);
nor UO_1164 (O_1164,N_28590,N_29360);
nor UO_1165 (O_1165,N_28823,N_29701);
nand UO_1166 (O_1166,N_29710,N_29403);
nor UO_1167 (O_1167,N_29550,N_29387);
nor UO_1168 (O_1168,N_29520,N_28612);
xnor UO_1169 (O_1169,N_29346,N_28658);
xor UO_1170 (O_1170,N_29446,N_29582);
nand UO_1171 (O_1171,N_29704,N_29376);
or UO_1172 (O_1172,N_29784,N_29918);
nor UO_1173 (O_1173,N_28653,N_29630);
nor UO_1174 (O_1174,N_29255,N_29149);
nor UO_1175 (O_1175,N_28799,N_29456);
nor UO_1176 (O_1176,N_29618,N_29072);
nor UO_1177 (O_1177,N_29484,N_29513);
and UO_1178 (O_1178,N_28801,N_28853);
xnor UO_1179 (O_1179,N_29261,N_29806);
and UO_1180 (O_1180,N_29313,N_29554);
and UO_1181 (O_1181,N_29681,N_29427);
or UO_1182 (O_1182,N_29896,N_29238);
and UO_1183 (O_1183,N_29549,N_29989);
nand UO_1184 (O_1184,N_29408,N_28955);
and UO_1185 (O_1185,N_28563,N_29307);
nor UO_1186 (O_1186,N_28605,N_29859);
or UO_1187 (O_1187,N_29479,N_29889);
nor UO_1188 (O_1188,N_29090,N_29782);
xor UO_1189 (O_1189,N_29368,N_28531);
nor UO_1190 (O_1190,N_29595,N_28661);
xor UO_1191 (O_1191,N_29146,N_29539);
and UO_1192 (O_1192,N_29008,N_28548);
xor UO_1193 (O_1193,N_28670,N_29634);
and UO_1194 (O_1194,N_29822,N_29995);
or UO_1195 (O_1195,N_29036,N_29919);
or UO_1196 (O_1196,N_28836,N_29340);
xnor UO_1197 (O_1197,N_29886,N_29280);
xor UO_1198 (O_1198,N_29695,N_29910);
nand UO_1199 (O_1199,N_29763,N_29753);
xnor UO_1200 (O_1200,N_29343,N_29597);
and UO_1201 (O_1201,N_29788,N_29121);
or UO_1202 (O_1202,N_28565,N_29490);
and UO_1203 (O_1203,N_28509,N_28744);
nor UO_1204 (O_1204,N_29925,N_28908);
nand UO_1205 (O_1205,N_28784,N_29046);
xor UO_1206 (O_1206,N_29622,N_29595);
or UO_1207 (O_1207,N_29691,N_29345);
nor UO_1208 (O_1208,N_29271,N_28756);
nor UO_1209 (O_1209,N_29945,N_29213);
xnor UO_1210 (O_1210,N_29410,N_29711);
xnor UO_1211 (O_1211,N_29024,N_29358);
xor UO_1212 (O_1212,N_29116,N_28931);
nand UO_1213 (O_1213,N_29401,N_29854);
nor UO_1214 (O_1214,N_28630,N_29545);
nand UO_1215 (O_1215,N_29205,N_29946);
or UO_1216 (O_1216,N_29112,N_29632);
nor UO_1217 (O_1217,N_28842,N_29206);
xnor UO_1218 (O_1218,N_29439,N_29911);
nand UO_1219 (O_1219,N_29713,N_28858);
nand UO_1220 (O_1220,N_29123,N_28552);
and UO_1221 (O_1221,N_29684,N_29917);
nor UO_1222 (O_1222,N_29398,N_29055);
xor UO_1223 (O_1223,N_29199,N_28890);
and UO_1224 (O_1224,N_29228,N_29361);
or UO_1225 (O_1225,N_28841,N_28929);
and UO_1226 (O_1226,N_29447,N_29911);
and UO_1227 (O_1227,N_29088,N_28937);
nand UO_1228 (O_1228,N_28777,N_28903);
nand UO_1229 (O_1229,N_29171,N_28907);
or UO_1230 (O_1230,N_29485,N_29184);
and UO_1231 (O_1231,N_28822,N_29327);
nand UO_1232 (O_1232,N_28902,N_29516);
and UO_1233 (O_1233,N_28884,N_28830);
or UO_1234 (O_1234,N_29149,N_29494);
nor UO_1235 (O_1235,N_29118,N_28676);
or UO_1236 (O_1236,N_29230,N_29900);
xor UO_1237 (O_1237,N_29262,N_29168);
or UO_1238 (O_1238,N_29903,N_28749);
or UO_1239 (O_1239,N_29986,N_29988);
xor UO_1240 (O_1240,N_29214,N_29174);
xnor UO_1241 (O_1241,N_28870,N_29468);
and UO_1242 (O_1242,N_29594,N_29714);
or UO_1243 (O_1243,N_28655,N_28789);
nand UO_1244 (O_1244,N_29086,N_29037);
or UO_1245 (O_1245,N_29773,N_28663);
or UO_1246 (O_1246,N_29907,N_29695);
xnor UO_1247 (O_1247,N_29901,N_29779);
and UO_1248 (O_1248,N_28733,N_29674);
nor UO_1249 (O_1249,N_29314,N_29049);
nand UO_1250 (O_1250,N_29664,N_28902);
and UO_1251 (O_1251,N_29199,N_29789);
xnor UO_1252 (O_1252,N_28590,N_29299);
xor UO_1253 (O_1253,N_28748,N_29143);
nand UO_1254 (O_1254,N_28531,N_29067);
nor UO_1255 (O_1255,N_29140,N_29832);
nand UO_1256 (O_1256,N_29434,N_28942);
xor UO_1257 (O_1257,N_29508,N_29670);
and UO_1258 (O_1258,N_29044,N_29363);
xor UO_1259 (O_1259,N_29542,N_28723);
xnor UO_1260 (O_1260,N_29665,N_29907);
or UO_1261 (O_1261,N_29387,N_29428);
xnor UO_1262 (O_1262,N_29396,N_29527);
nand UO_1263 (O_1263,N_29239,N_29855);
or UO_1264 (O_1264,N_28940,N_29077);
xnor UO_1265 (O_1265,N_29792,N_29289);
and UO_1266 (O_1266,N_28937,N_29427);
xor UO_1267 (O_1267,N_29277,N_29000);
nand UO_1268 (O_1268,N_29329,N_29859);
xnor UO_1269 (O_1269,N_29447,N_29782);
or UO_1270 (O_1270,N_29260,N_28558);
nand UO_1271 (O_1271,N_28945,N_28572);
or UO_1272 (O_1272,N_28866,N_28992);
and UO_1273 (O_1273,N_29890,N_29215);
and UO_1274 (O_1274,N_29479,N_28552);
nor UO_1275 (O_1275,N_28540,N_29175);
or UO_1276 (O_1276,N_29756,N_28778);
xor UO_1277 (O_1277,N_29781,N_28717);
and UO_1278 (O_1278,N_29776,N_28553);
or UO_1279 (O_1279,N_29951,N_28839);
or UO_1280 (O_1280,N_29104,N_28806);
xnor UO_1281 (O_1281,N_29196,N_28621);
nor UO_1282 (O_1282,N_29498,N_28616);
and UO_1283 (O_1283,N_29483,N_28946);
nor UO_1284 (O_1284,N_29893,N_28806);
nor UO_1285 (O_1285,N_29550,N_29965);
and UO_1286 (O_1286,N_29952,N_29406);
or UO_1287 (O_1287,N_28833,N_28589);
or UO_1288 (O_1288,N_28940,N_29742);
or UO_1289 (O_1289,N_29701,N_29029);
and UO_1290 (O_1290,N_29128,N_29452);
nand UO_1291 (O_1291,N_29810,N_29469);
xor UO_1292 (O_1292,N_29808,N_28836);
or UO_1293 (O_1293,N_28565,N_29025);
and UO_1294 (O_1294,N_29814,N_29889);
and UO_1295 (O_1295,N_29528,N_29524);
xnor UO_1296 (O_1296,N_29214,N_28864);
nor UO_1297 (O_1297,N_28958,N_29030);
and UO_1298 (O_1298,N_29928,N_28544);
and UO_1299 (O_1299,N_29322,N_28534);
xor UO_1300 (O_1300,N_29424,N_28901);
nor UO_1301 (O_1301,N_29019,N_28905);
nor UO_1302 (O_1302,N_29999,N_29940);
nand UO_1303 (O_1303,N_28735,N_29807);
or UO_1304 (O_1304,N_29770,N_29077);
and UO_1305 (O_1305,N_29019,N_29068);
and UO_1306 (O_1306,N_28871,N_29913);
nor UO_1307 (O_1307,N_28807,N_28518);
or UO_1308 (O_1308,N_29930,N_29139);
xor UO_1309 (O_1309,N_29176,N_28746);
xor UO_1310 (O_1310,N_28598,N_28808);
or UO_1311 (O_1311,N_29201,N_29825);
xor UO_1312 (O_1312,N_29238,N_28810);
xor UO_1313 (O_1313,N_28653,N_29281);
or UO_1314 (O_1314,N_28723,N_28669);
nor UO_1315 (O_1315,N_29332,N_28500);
nor UO_1316 (O_1316,N_28785,N_29515);
and UO_1317 (O_1317,N_29338,N_29722);
xor UO_1318 (O_1318,N_28728,N_29131);
xnor UO_1319 (O_1319,N_29167,N_29203);
nand UO_1320 (O_1320,N_29757,N_29369);
and UO_1321 (O_1321,N_29332,N_29006);
and UO_1322 (O_1322,N_28772,N_29487);
xor UO_1323 (O_1323,N_29693,N_29118);
nand UO_1324 (O_1324,N_28535,N_28626);
or UO_1325 (O_1325,N_29719,N_29226);
nand UO_1326 (O_1326,N_29071,N_29750);
and UO_1327 (O_1327,N_28838,N_28529);
and UO_1328 (O_1328,N_29207,N_28668);
nand UO_1329 (O_1329,N_29805,N_29908);
xnor UO_1330 (O_1330,N_29664,N_29746);
nand UO_1331 (O_1331,N_29336,N_28851);
nand UO_1332 (O_1332,N_28815,N_28986);
nand UO_1333 (O_1333,N_29837,N_28931);
nand UO_1334 (O_1334,N_28888,N_29670);
or UO_1335 (O_1335,N_28881,N_28712);
nand UO_1336 (O_1336,N_29049,N_28680);
and UO_1337 (O_1337,N_28665,N_29650);
xnor UO_1338 (O_1338,N_29832,N_29464);
xnor UO_1339 (O_1339,N_29568,N_28599);
nand UO_1340 (O_1340,N_28614,N_28602);
nor UO_1341 (O_1341,N_29263,N_28931);
xor UO_1342 (O_1342,N_29459,N_29082);
or UO_1343 (O_1343,N_28901,N_29996);
or UO_1344 (O_1344,N_28522,N_28662);
xor UO_1345 (O_1345,N_29930,N_29048);
and UO_1346 (O_1346,N_29761,N_29836);
and UO_1347 (O_1347,N_28569,N_28997);
nand UO_1348 (O_1348,N_29988,N_29502);
nand UO_1349 (O_1349,N_29051,N_28953);
or UO_1350 (O_1350,N_29320,N_29768);
nand UO_1351 (O_1351,N_29889,N_28879);
and UO_1352 (O_1352,N_28550,N_29876);
nand UO_1353 (O_1353,N_28974,N_29998);
and UO_1354 (O_1354,N_28632,N_29200);
xor UO_1355 (O_1355,N_29856,N_29557);
nand UO_1356 (O_1356,N_28794,N_29044);
nand UO_1357 (O_1357,N_28934,N_29030);
xnor UO_1358 (O_1358,N_28518,N_28789);
or UO_1359 (O_1359,N_29149,N_28856);
and UO_1360 (O_1360,N_28912,N_29761);
xor UO_1361 (O_1361,N_29558,N_29638);
or UO_1362 (O_1362,N_29020,N_29328);
xnor UO_1363 (O_1363,N_29531,N_29513);
and UO_1364 (O_1364,N_29366,N_28639);
or UO_1365 (O_1365,N_29175,N_29806);
xnor UO_1366 (O_1366,N_29023,N_28860);
xnor UO_1367 (O_1367,N_29455,N_28612);
xor UO_1368 (O_1368,N_28503,N_29091);
or UO_1369 (O_1369,N_29820,N_28646);
or UO_1370 (O_1370,N_28574,N_29569);
xnor UO_1371 (O_1371,N_29797,N_29372);
nor UO_1372 (O_1372,N_29792,N_29840);
or UO_1373 (O_1373,N_29984,N_29749);
or UO_1374 (O_1374,N_28902,N_28569);
nor UO_1375 (O_1375,N_28598,N_29031);
and UO_1376 (O_1376,N_29700,N_28914);
nor UO_1377 (O_1377,N_28702,N_29333);
nor UO_1378 (O_1378,N_29491,N_29670);
nor UO_1379 (O_1379,N_29255,N_29237);
xor UO_1380 (O_1380,N_29279,N_29061);
xor UO_1381 (O_1381,N_29737,N_29110);
xor UO_1382 (O_1382,N_28764,N_29661);
nand UO_1383 (O_1383,N_29616,N_28874);
xnor UO_1384 (O_1384,N_29387,N_28922);
or UO_1385 (O_1385,N_28672,N_28555);
nor UO_1386 (O_1386,N_28780,N_29653);
and UO_1387 (O_1387,N_29743,N_29506);
nor UO_1388 (O_1388,N_29235,N_29223);
or UO_1389 (O_1389,N_29268,N_29664);
nand UO_1390 (O_1390,N_29036,N_29615);
nand UO_1391 (O_1391,N_28648,N_29579);
and UO_1392 (O_1392,N_28829,N_29460);
xor UO_1393 (O_1393,N_29441,N_28720);
xor UO_1394 (O_1394,N_29197,N_29219);
or UO_1395 (O_1395,N_28928,N_29226);
xor UO_1396 (O_1396,N_29013,N_28816);
or UO_1397 (O_1397,N_29809,N_29040);
nand UO_1398 (O_1398,N_29415,N_28957);
nand UO_1399 (O_1399,N_29733,N_28836);
nand UO_1400 (O_1400,N_29715,N_29931);
and UO_1401 (O_1401,N_29112,N_29232);
nor UO_1402 (O_1402,N_29961,N_29265);
or UO_1403 (O_1403,N_28686,N_29668);
nand UO_1404 (O_1404,N_29652,N_28611);
nor UO_1405 (O_1405,N_29593,N_29611);
and UO_1406 (O_1406,N_29142,N_29875);
and UO_1407 (O_1407,N_29222,N_29929);
and UO_1408 (O_1408,N_29391,N_29739);
or UO_1409 (O_1409,N_29024,N_28706);
or UO_1410 (O_1410,N_29310,N_29578);
nor UO_1411 (O_1411,N_29494,N_28712);
nor UO_1412 (O_1412,N_29935,N_28757);
nor UO_1413 (O_1413,N_29891,N_29199);
nand UO_1414 (O_1414,N_28813,N_29473);
xnor UO_1415 (O_1415,N_29720,N_29505);
nor UO_1416 (O_1416,N_29093,N_29835);
nor UO_1417 (O_1417,N_29883,N_29525);
and UO_1418 (O_1418,N_29549,N_29640);
and UO_1419 (O_1419,N_29160,N_29200);
and UO_1420 (O_1420,N_29678,N_28540);
or UO_1421 (O_1421,N_29164,N_28679);
xnor UO_1422 (O_1422,N_28661,N_28664);
nor UO_1423 (O_1423,N_28512,N_29948);
xnor UO_1424 (O_1424,N_28974,N_28876);
nor UO_1425 (O_1425,N_29196,N_29024);
xnor UO_1426 (O_1426,N_29882,N_28901);
and UO_1427 (O_1427,N_29350,N_29695);
nor UO_1428 (O_1428,N_29824,N_29565);
nor UO_1429 (O_1429,N_28914,N_28669);
nand UO_1430 (O_1430,N_28920,N_28903);
xor UO_1431 (O_1431,N_29169,N_29420);
and UO_1432 (O_1432,N_29672,N_29234);
or UO_1433 (O_1433,N_29829,N_29811);
nand UO_1434 (O_1434,N_28555,N_29809);
nor UO_1435 (O_1435,N_28970,N_28572);
xor UO_1436 (O_1436,N_29820,N_29221);
nand UO_1437 (O_1437,N_29169,N_29409);
nand UO_1438 (O_1438,N_28752,N_29376);
or UO_1439 (O_1439,N_29254,N_29638);
and UO_1440 (O_1440,N_29135,N_29432);
and UO_1441 (O_1441,N_29622,N_29407);
and UO_1442 (O_1442,N_28702,N_29631);
nor UO_1443 (O_1443,N_29613,N_29190);
nor UO_1444 (O_1444,N_28824,N_29217);
nand UO_1445 (O_1445,N_28900,N_29161);
or UO_1446 (O_1446,N_29101,N_29760);
nand UO_1447 (O_1447,N_29458,N_29024);
nand UO_1448 (O_1448,N_29310,N_29065);
xor UO_1449 (O_1449,N_28798,N_28962);
xnor UO_1450 (O_1450,N_29943,N_29260);
and UO_1451 (O_1451,N_29058,N_29514);
nand UO_1452 (O_1452,N_29601,N_29715);
and UO_1453 (O_1453,N_29225,N_29918);
xor UO_1454 (O_1454,N_28911,N_29963);
nor UO_1455 (O_1455,N_28978,N_29376);
and UO_1456 (O_1456,N_29003,N_29673);
nand UO_1457 (O_1457,N_29157,N_28965);
xnor UO_1458 (O_1458,N_28679,N_28680);
nand UO_1459 (O_1459,N_28712,N_28918);
nand UO_1460 (O_1460,N_28854,N_29094);
nand UO_1461 (O_1461,N_29081,N_28558);
or UO_1462 (O_1462,N_28626,N_29735);
and UO_1463 (O_1463,N_29069,N_29398);
and UO_1464 (O_1464,N_29375,N_28944);
xor UO_1465 (O_1465,N_28936,N_28995);
and UO_1466 (O_1466,N_28953,N_28933);
or UO_1467 (O_1467,N_28947,N_29022);
xnor UO_1468 (O_1468,N_29530,N_29692);
and UO_1469 (O_1469,N_29242,N_28668);
nand UO_1470 (O_1470,N_29156,N_28701);
nand UO_1471 (O_1471,N_28610,N_29393);
xor UO_1472 (O_1472,N_29754,N_29968);
nor UO_1473 (O_1473,N_28775,N_28503);
xnor UO_1474 (O_1474,N_29350,N_29148);
nand UO_1475 (O_1475,N_28704,N_28837);
nor UO_1476 (O_1476,N_28651,N_29420);
xor UO_1477 (O_1477,N_29109,N_29639);
nor UO_1478 (O_1478,N_29758,N_28604);
nor UO_1479 (O_1479,N_29362,N_28561);
and UO_1480 (O_1480,N_29685,N_28752);
and UO_1481 (O_1481,N_29046,N_29650);
nor UO_1482 (O_1482,N_29737,N_29234);
or UO_1483 (O_1483,N_29814,N_29715);
or UO_1484 (O_1484,N_29609,N_29657);
and UO_1485 (O_1485,N_28693,N_28937);
or UO_1486 (O_1486,N_29828,N_29302);
nand UO_1487 (O_1487,N_29045,N_29620);
nor UO_1488 (O_1488,N_28856,N_29175);
nand UO_1489 (O_1489,N_29349,N_29889);
nand UO_1490 (O_1490,N_28864,N_28546);
xnor UO_1491 (O_1491,N_29068,N_28868);
or UO_1492 (O_1492,N_29835,N_29185);
nor UO_1493 (O_1493,N_29339,N_28783);
and UO_1494 (O_1494,N_28766,N_28676);
or UO_1495 (O_1495,N_29801,N_28754);
nor UO_1496 (O_1496,N_29473,N_28578);
nand UO_1497 (O_1497,N_28815,N_28712);
nand UO_1498 (O_1498,N_28768,N_28651);
xor UO_1499 (O_1499,N_29668,N_29297);
xnor UO_1500 (O_1500,N_29823,N_29165);
or UO_1501 (O_1501,N_29044,N_29268);
or UO_1502 (O_1502,N_29312,N_29279);
nand UO_1503 (O_1503,N_28595,N_28857);
and UO_1504 (O_1504,N_28965,N_29035);
and UO_1505 (O_1505,N_29738,N_28537);
and UO_1506 (O_1506,N_29348,N_28965);
and UO_1507 (O_1507,N_29411,N_29127);
nand UO_1508 (O_1508,N_28916,N_29389);
nand UO_1509 (O_1509,N_29249,N_29865);
nor UO_1510 (O_1510,N_29371,N_28673);
xor UO_1511 (O_1511,N_29869,N_29023);
nor UO_1512 (O_1512,N_28540,N_29665);
nand UO_1513 (O_1513,N_29889,N_29514);
or UO_1514 (O_1514,N_28620,N_28855);
and UO_1515 (O_1515,N_29313,N_29178);
and UO_1516 (O_1516,N_29936,N_29229);
and UO_1517 (O_1517,N_28663,N_29415);
nor UO_1518 (O_1518,N_29352,N_28781);
and UO_1519 (O_1519,N_29426,N_29422);
xor UO_1520 (O_1520,N_29978,N_28761);
xnor UO_1521 (O_1521,N_29391,N_28917);
and UO_1522 (O_1522,N_29306,N_28520);
nor UO_1523 (O_1523,N_29334,N_28752);
or UO_1524 (O_1524,N_28603,N_28755);
nand UO_1525 (O_1525,N_29503,N_28788);
xnor UO_1526 (O_1526,N_28826,N_28691);
nor UO_1527 (O_1527,N_29837,N_29690);
nand UO_1528 (O_1528,N_29390,N_29958);
nand UO_1529 (O_1529,N_29740,N_29372);
and UO_1530 (O_1530,N_28748,N_29201);
or UO_1531 (O_1531,N_28888,N_29471);
xor UO_1532 (O_1532,N_29954,N_28884);
and UO_1533 (O_1533,N_29745,N_28776);
nor UO_1534 (O_1534,N_29351,N_29078);
or UO_1535 (O_1535,N_28629,N_29657);
or UO_1536 (O_1536,N_29731,N_29559);
xor UO_1537 (O_1537,N_28766,N_29524);
nor UO_1538 (O_1538,N_28652,N_29407);
nor UO_1539 (O_1539,N_29294,N_29301);
xnor UO_1540 (O_1540,N_28679,N_29968);
xnor UO_1541 (O_1541,N_29803,N_29208);
and UO_1542 (O_1542,N_29299,N_29357);
nor UO_1543 (O_1543,N_28782,N_29712);
and UO_1544 (O_1544,N_29068,N_29881);
xnor UO_1545 (O_1545,N_29537,N_29183);
xnor UO_1546 (O_1546,N_29247,N_29278);
or UO_1547 (O_1547,N_28654,N_28754);
or UO_1548 (O_1548,N_28994,N_29289);
or UO_1549 (O_1549,N_28653,N_29798);
nand UO_1550 (O_1550,N_28936,N_29208);
nand UO_1551 (O_1551,N_28640,N_28582);
or UO_1552 (O_1552,N_29140,N_28821);
or UO_1553 (O_1553,N_28779,N_29607);
nand UO_1554 (O_1554,N_28723,N_29210);
or UO_1555 (O_1555,N_28864,N_28507);
nor UO_1556 (O_1556,N_29219,N_29494);
nand UO_1557 (O_1557,N_28847,N_29712);
and UO_1558 (O_1558,N_28766,N_28532);
xor UO_1559 (O_1559,N_29380,N_28631);
xor UO_1560 (O_1560,N_28732,N_29785);
nor UO_1561 (O_1561,N_28948,N_28793);
nand UO_1562 (O_1562,N_28555,N_29881);
or UO_1563 (O_1563,N_29689,N_28612);
nor UO_1564 (O_1564,N_29298,N_29192);
nand UO_1565 (O_1565,N_28630,N_28800);
xor UO_1566 (O_1566,N_29308,N_28948);
nand UO_1567 (O_1567,N_29942,N_29581);
nand UO_1568 (O_1568,N_29462,N_29209);
or UO_1569 (O_1569,N_28973,N_29505);
nand UO_1570 (O_1570,N_29777,N_28951);
xor UO_1571 (O_1571,N_29016,N_29366);
nor UO_1572 (O_1572,N_29866,N_29912);
or UO_1573 (O_1573,N_29346,N_28544);
nor UO_1574 (O_1574,N_29971,N_29537);
and UO_1575 (O_1575,N_29318,N_29702);
nor UO_1576 (O_1576,N_29570,N_29569);
or UO_1577 (O_1577,N_29050,N_29540);
nor UO_1578 (O_1578,N_29648,N_29783);
nor UO_1579 (O_1579,N_29945,N_29724);
and UO_1580 (O_1580,N_29518,N_29672);
nor UO_1581 (O_1581,N_28717,N_29909);
nor UO_1582 (O_1582,N_29705,N_29454);
and UO_1583 (O_1583,N_29396,N_29801);
nand UO_1584 (O_1584,N_28688,N_29852);
nor UO_1585 (O_1585,N_29381,N_29665);
xor UO_1586 (O_1586,N_28512,N_28896);
and UO_1587 (O_1587,N_29313,N_29088);
xor UO_1588 (O_1588,N_28848,N_28663);
nand UO_1589 (O_1589,N_28731,N_28886);
or UO_1590 (O_1590,N_29032,N_29780);
xnor UO_1591 (O_1591,N_28972,N_28645);
nor UO_1592 (O_1592,N_28778,N_28589);
and UO_1593 (O_1593,N_29411,N_28502);
nor UO_1594 (O_1594,N_29748,N_29564);
nor UO_1595 (O_1595,N_28545,N_29697);
or UO_1596 (O_1596,N_28685,N_28715);
and UO_1597 (O_1597,N_29870,N_28903);
nand UO_1598 (O_1598,N_29948,N_29708);
and UO_1599 (O_1599,N_29024,N_29333);
or UO_1600 (O_1600,N_29923,N_28732);
and UO_1601 (O_1601,N_28587,N_28534);
or UO_1602 (O_1602,N_29904,N_28865);
or UO_1603 (O_1603,N_29678,N_29633);
or UO_1604 (O_1604,N_28776,N_29060);
or UO_1605 (O_1605,N_28961,N_28864);
or UO_1606 (O_1606,N_29781,N_29123);
nor UO_1607 (O_1607,N_28934,N_29576);
or UO_1608 (O_1608,N_28827,N_29925);
xnor UO_1609 (O_1609,N_29118,N_29099);
or UO_1610 (O_1610,N_29537,N_29615);
nand UO_1611 (O_1611,N_28972,N_29201);
and UO_1612 (O_1612,N_28897,N_29345);
or UO_1613 (O_1613,N_28529,N_28650);
or UO_1614 (O_1614,N_28653,N_29523);
xnor UO_1615 (O_1615,N_29583,N_29967);
nor UO_1616 (O_1616,N_29805,N_29872);
or UO_1617 (O_1617,N_28530,N_28876);
nor UO_1618 (O_1618,N_28770,N_28973);
or UO_1619 (O_1619,N_28629,N_29176);
xor UO_1620 (O_1620,N_28501,N_29826);
xor UO_1621 (O_1621,N_29358,N_29205);
or UO_1622 (O_1622,N_29070,N_29094);
or UO_1623 (O_1623,N_29520,N_28808);
or UO_1624 (O_1624,N_29374,N_29229);
or UO_1625 (O_1625,N_28528,N_28504);
and UO_1626 (O_1626,N_28723,N_28817);
nor UO_1627 (O_1627,N_29703,N_29903);
nor UO_1628 (O_1628,N_29811,N_28610);
nor UO_1629 (O_1629,N_29034,N_29391);
xor UO_1630 (O_1630,N_29988,N_29545);
nor UO_1631 (O_1631,N_29057,N_29801);
nor UO_1632 (O_1632,N_29423,N_28549);
nor UO_1633 (O_1633,N_29268,N_28938);
nand UO_1634 (O_1634,N_29487,N_28799);
and UO_1635 (O_1635,N_29868,N_29381);
and UO_1636 (O_1636,N_29588,N_29355);
nor UO_1637 (O_1637,N_29484,N_29315);
or UO_1638 (O_1638,N_29954,N_28824);
xor UO_1639 (O_1639,N_28891,N_28832);
and UO_1640 (O_1640,N_28799,N_29672);
or UO_1641 (O_1641,N_29817,N_28579);
xor UO_1642 (O_1642,N_28891,N_29747);
or UO_1643 (O_1643,N_29811,N_29791);
xor UO_1644 (O_1644,N_29891,N_29023);
xnor UO_1645 (O_1645,N_28602,N_29279);
and UO_1646 (O_1646,N_29014,N_28775);
xnor UO_1647 (O_1647,N_28590,N_28696);
and UO_1648 (O_1648,N_29969,N_29375);
or UO_1649 (O_1649,N_29055,N_28713);
or UO_1650 (O_1650,N_28569,N_29391);
xnor UO_1651 (O_1651,N_29651,N_29326);
xnor UO_1652 (O_1652,N_29580,N_29936);
and UO_1653 (O_1653,N_28674,N_28609);
nand UO_1654 (O_1654,N_29986,N_29442);
and UO_1655 (O_1655,N_29554,N_28845);
and UO_1656 (O_1656,N_28514,N_28767);
and UO_1657 (O_1657,N_28976,N_28793);
nor UO_1658 (O_1658,N_28923,N_29611);
and UO_1659 (O_1659,N_29131,N_29043);
nand UO_1660 (O_1660,N_28841,N_29442);
xnor UO_1661 (O_1661,N_28829,N_29298);
nor UO_1662 (O_1662,N_29746,N_28880);
or UO_1663 (O_1663,N_29794,N_28931);
nor UO_1664 (O_1664,N_29953,N_28975);
and UO_1665 (O_1665,N_29545,N_28624);
xnor UO_1666 (O_1666,N_28913,N_29341);
nand UO_1667 (O_1667,N_29457,N_29423);
nand UO_1668 (O_1668,N_29728,N_28779);
or UO_1669 (O_1669,N_28989,N_29061);
nor UO_1670 (O_1670,N_29113,N_29519);
nor UO_1671 (O_1671,N_29713,N_29042);
and UO_1672 (O_1672,N_28868,N_28772);
and UO_1673 (O_1673,N_29521,N_28554);
nand UO_1674 (O_1674,N_29731,N_29306);
nand UO_1675 (O_1675,N_29597,N_29767);
xnor UO_1676 (O_1676,N_29720,N_29923);
xor UO_1677 (O_1677,N_29773,N_28675);
and UO_1678 (O_1678,N_29408,N_28799);
nor UO_1679 (O_1679,N_29924,N_28567);
or UO_1680 (O_1680,N_29700,N_28639);
nor UO_1681 (O_1681,N_29554,N_29696);
xnor UO_1682 (O_1682,N_29950,N_29369);
or UO_1683 (O_1683,N_29471,N_28796);
xor UO_1684 (O_1684,N_29397,N_29295);
or UO_1685 (O_1685,N_29971,N_29820);
and UO_1686 (O_1686,N_29458,N_28663);
nand UO_1687 (O_1687,N_28579,N_28632);
xor UO_1688 (O_1688,N_28557,N_29973);
and UO_1689 (O_1689,N_28914,N_29807);
xnor UO_1690 (O_1690,N_28948,N_29681);
nand UO_1691 (O_1691,N_29487,N_29930);
and UO_1692 (O_1692,N_29023,N_29888);
nand UO_1693 (O_1693,N_29120,N_29110);
and UO_1694 (O_1694,N_29419,N_29888);
nand UO_1695 (O_1695,N_28736,N_28881);
nand UO_1696 (O_1696,N_29045,N_28754);
xor UO_1697 (O_1697,N_29908,N_29575);
or UO_1698 (O_1698,N_29633,N_28556);
nand UO_1699 (O_1699,N_28934,N_29254);
xnor UO_1700 (O_1700,N_29749,N_29882);
xor UO_1701 (O_1701,N_28744,N_29083);
and UO_1702 (O_1702,N_29117,N_29094);
and UO_1703 (O_1703,N_29806,N_28953);
xor UO_1704 (O_1704,N_28509,N_28655);
or UO_1705 (O_1705,N_29824,N_29009);
nand UO_1706 (O_1706,N_29060,N_29890);
or UO_1707 (O_1707,N_28694,N_29207);
xnor UO_1708 (O_1708,N_28535,N_29100);
or UO_1709 (O_1709,N_28731,N_28923);
nand UO_1710 (O_1710,N_28841,N_29083);
and UO_1711 (O_1711,N_29237,N_29431);
xnor UO_1712 (O_1712,N_29057,N_29163);
xnor UO_1713 (O_1713,N_28695,N_29148);
nand UO_1714 (O_1714,N_28723,N_29992);
or UO_1715 (O_1715,N_28711,N_29714);
or UO_1716 (O_1716,N_28710,N_29191);
and UO_1717 (O_1717,N_29976,N_29066);
or UO_1718 (O_1718,N_28695,N_29444);
nand UO_1719 (O_1719,N_29441,N_28955);
or UO_1720 (O_1720,N_29356,N_29808);
nand UO_1721 (O_1721,N_29025,N_29628);
nand UO_1722 (O_1722,N_29771,N_28778);
nand UO_1723 (O_1723,N_29925,N_29404);
xor UO_1724 (O_1724,N_29426,N_28728);
nand UO_1725 (O_1725,N_29626,N_28985);
and UO_1726 (O_1726,N_29588,N_28937);
and UO_1727 (O_1727,N_28748,N_28788);
or UO_1728 (O_1728,N_28523,N_29369);
nand UO_1729 (O_1729,N_28522,N_29476);
xnor UO_1730 (O_1730,N_29765,N_29114);
xor UO_1731 (O_1731,N_28910,N_28859);
nand UO_1732 (O_1732,N_29328,N_29408);
or UO_1733 (O_1733,N_28880,N_29928);
nor UO_1734 (O_1734,N_29795,N_28780);
and UO_1735 (O_1735,N_29628,N_28512);
nand UO_1736 (O_1736,N_28699,N_28525);
nand UO_1737 (O_1737,N_28553,N_29022);
nor UO_1738 (O_1738,N_28722,N_29156);
or UO_1739 (O_1739,N_29658,N_29614);
or UO_1740 (O_1740,N_28630,N_29497);
xnor UO_1741 (O_1741,N_29672,N_29184);
nor UO_1742 (O_1742,N_29921,N_29058);
nand UO_1743 (O_1743,N_29023,N_29315);
and UO_1744 (O_1744,N_29346,N_29791);
xnor UO_1745 (O_1745,N_28786,N_29588);
or UO_1746 (O_1746,N_29319,N_28812);
xor UO_1747 (O_1747,N_29049,N_28852);
xnor UO_1748 (O_1748,N_29994,N_28915);
and UO_1749 (O_1749,N_29202,N_28549);
and UO_1750 (O_1750,N_29244,N_29527);
nor UO_1751 (O_1751,N_29672,N_29131);
and UO_1752 (O_1752,N_29578,N_28810);
nor UO_1753 (O_1753,N_28951,N_28505);
or UO_1754 (O_1754,N_29736,N_28609);
nor UO_1755 (O_1755,N_29642,N_29237);
nand UO_1756 (O_1756,N_29509,N_29466);
or UO_1757 (O_1757,N_29256,N_28902);
or UO_1758 (O_1758,N_29902,N_29101);
or UO_1759 (O_1759,N_28790,N_29983);
xnor UO_1760 (O_1760,N_28903,N_28884);
nor UO_1761 (O_1761,N_29440,N_29002);
nor UO_1762 (O_1762,N_28927,N_29526);
xor UO_1763 (O_1763,N_29674,N_29974);
and UO_1764 (O_1764,N_29442,N_29213);
and UO_1765 (O_1765,N_29042,N_28746);
nor UO_1766 (O_1766,N_28704,N_28805);
nand UO_1767 (O_1767,N_29754,N_29214);
and UO_1768 (O_1768,N_29595,N_28906);
xor UO_1769 (O_1769,N_29707,N_28939);
xnor UO_1770 (O_1770,N_28744,N_28794);
or UO_1771 (O_1771,N_29949,N_29533);
and UO_1772 (O_1772,N_29298,N_28522);
and UO_1773 (O_1773,N_29807,N_29089);
nor UO_1774 (O_1774,N_29920,N_28902);
nor UO_1775 (O_1775,N_29576,N_29835);
nor UO_1776 (O_1776,N_29444,N_29098);
xnor UO_1777 (O_1777,N_29835,N_29304);
nor UO_1778 (O_1778,N_28835,N_29822);
nand UO_1779 (O_1779,N_29597,N_29106);
and UO_1780 (O_1780,N_29932,N_28654);
and UO_1781 (O_1781,N_29456,N_29534);
nor UO_1782 (O_1782,N_29551,N_29411);
or UO_1783 (O_1783,N_29581,N_28598);
nor UO_1784 (O_1784,N_29861,N_29055);
or UO_1785 (O_1785,N_29113,N_29135);
nor UO_1786 (O_1786,N_29833,N_29602);
nand UO_1787 (O_1787,N_29727,N_29984);
nand UO_1788 (O_1788,N_29567,N_28856);
xnor UO_1789 (O_1789,N_29745,N_29568);
or UO_1790 (O_1790,N_28642,N_29553);
nor UO_1791 (O_1791,N_28543,N_29096);
xnor UO_1792 (O_1792,N_28522,N_29643);
or UO_1793 (O_1793,N_29624,N_29763);
or UO_1794 (O_1794,N_29674,N_29131);
xor UO_1795 (O_1795,N_29672,N_28517);
nor UO_1796 (O_1796,N_29442,N_29733);
nor UO_1797 (O_1797,N_28530,N_28846);
nand UO_1798 (O_1798,N_29701,N_28717);
xor UO_1799 (O_1799,N_29610,N_28897);
and UO_1800 (O_1800,N_29648,N_29291);
nor UO_1801 (O_1801,N_29355,N_28628);
nand UO_1802 (O_1802,N_28979,N_28563);
nor UO_1803 (O_1803,N_29889,N_29661);
xnor UO_1804 (O_1804,N_28707,N_29967);
nand UO_1805 (O_1805,N_28829,N_29776);
or UO_1806 (O_1806,N_29479,N_28691);
nand UO_1807 (O_1807,N_29144,N_29629);
nor UO_1808 (O_1808,N_29236,N_29778);
nand UO_1809 (O_1809,N_29359,N_29311);
nor UO_1810 (O_1810,N_29576,N_29587);
nand UO_1811 (O_1811,N_28833,N_29793);
and UO_1812 (O_1812,N_28612,N_29917);
nor UO_1813 (O_1813,N_29669,N_29703);
xor UO_1814 (O_1814,N_29900,N_29478);
or UO_1815 (O_1815,N_29172,N_29529);
xnor UO_1816 (O_1816,N_29786,N_28851);
and UO_1817 (O_1817,N_29308,N_29213);
and UO_1818 (O_1818,N_28956,N_28651);
and UO_1819 (O_1819,N_29749,N_29139);
or UO_1820 (O_1820,N_28628,N_28646);
and UO_1821 (O_1821,N_29367,N_29608);
or UO_1822 (O_1822,N_29100,N_29782);
or UO_1823 (O_1823,N_29505,N_29730);
or UO_1824 (O_1824,N_29849,N_29761);
nor UO_1825 (O_1825,N_28950,N_29964);
xor UO_1826 (O_1826,N_28504,N_29320);
xnor UO_1827 (O_1827,N_29355,N_29530);
xor UO_1828 (O_1828,N_29637,N_29048);
or UO_1829 (O_1829,N_29476,N_29130);
nand UO_1830 (O_1830,N_29071,N_29053);
nor UO_1831 (O_1831,N_29026,N_28731);
or UO_1832 (O_1832,N_28944,N_28637);
and UO_1833 (O_1833,N_28874,N_29142);
or UO_1834 (O_1834,N_29571,N_28708);
xor UO_1835 (O_1835,N_28516,N_29123);
nor UO_1836 (O_1836,N_28651,N_28815);
xor UO_1837 (O_1837,N_28550,N_29823);
xor UO_1838 (O_1838,N_29463,N_29887);
and UO_1839 (O_1839,N_29862,N_28646);
nand UO_1840 (O_1840,N_28828,N_28500);
xnor UO_1841 (O_1841,N_28789,N_29062);
nand UO_1842 (O_1842,N_29458,N_29716);
nand UO_1843 (O_1843,N_29302,N_29566);
xnor UO_1844 (O_1844,N_28934,N_28886);
or UO_1845 (O_1845,N_29682,N_29542);
and UO_1846 (O_1846,N_28782,N_29786);
xnor UO_1847 (O_1847,N_29498,N_29295);
and UO_1848 (O_1848,N_29537,N_29692);
nand UO_1849 (O_1849,N_28792,N_29133);
nand UO_1850 (O_1850,N_29004,N_29454);
or UO_1851 (O_1851,N_29078,N_29371);
xnor UO_1852 (O_1852,N_29042,N_29869);
nor UO_1853 (O_1853,N_28654,N_29100);
nor UO_1854 (O_1854,N_29380,N_29680);
or UO_1855 (O_1855,N_29812,N_28622);
nor UO_1856 (O_1856,N_29809,N_29546);
nor UO_1857 (O_1857,N_28600,N_28756);
nand UO_1858 (O_1858,N_29674,N_29391);
nand UO_1859 (O_1859,N_28631,N_29686);
nand UO_1860 (O_1860,N_29794,N_29057);
nor UO_1861 (O_1861,N_29198,N_29253);
xnor UO_1862 (O_1862,N_29677,N_29578);
nand UO_1863 (O_1863,N_29308,N_28666);
or UO_1864 (O_1864,N_28983,N_29811);
nor UO_1865 (O_1865,N_29789,N_29876);
nor UO_1866 (O_1866,N_29906,N_28680);
xnor UO_1867 (O_1867,N_29586,N_28656);
nor UO_1868 (O_1868,N_28629,N_29719);
nor UO_1869 (O_1869,N_28737,N_29337);
nor UO_1870 (O_1870,N_29166,N_29838);
and UO_1871 (O_1871,N_29770,N_28951);
xor UO_1872 (O_1872,N_29797,N_29560);
and UO_1873 (O_1873,N_29368,N_29344);
and UO_1874 (O_1874,N_28863,N_28733);
nand UO_1875 (O_1875,N_29147,N_29123);
xor UO_1876 (O_1876,N_28802,N_29801);
xnor UO_1877 (O_1877,N_28901,N_29708);
nand UO_1878 (O_1878,N_28542,N_28994);
xnor UO_1879 (O_1879,N_29798,N_29700);
nand UO_1880 (O_1880,N_29724,N_28769);
nor UO_1881 (O_1881,N_28834,N_28935);
nor UO_1882 (O_1882,N_29192,N_29180);
or UO_1883 (O_1883,N_29323,N_29576);
nor UO_1884 (O_1884,N_29571,N_28815);
nor UO_1885 (O_1885,N_29828,N_29095);
and UO_1886 (O_1886,N_29843,N_29847);
xor UO_1887 (O_1887,N_28973,N_28602);
xor UO_1888 (O_1888,N_28959,N_29719);
and UO_1889 (O_1889,N_29987,N_29197);
nand UO_1890 (O_1890,N_29210,N_28879);
nor UO_1891 (O_1891,N_29075,N_28555);
xnor UO_1892 (O_1892,N_29160,N_28657);
nor UO_1893 (O_1893,N_28706,N_29262);
or UO_1894 (O_1894,N_29056,N_29732);
or UO_1895 (O_1895,N_29132,N_29122);
xor UO_1896 (O_1896,N_29377,N_29828);
xnor UO_1897 (O_1897,N_28852,N_29863);
or UO_1898 (O_1898,N_29899,N_29420);
xnor UO_1899 (O_1899,N_28610,N_29651);
or UO_1900 (O_1900,N_29191,N_28609);
and UO_1901 (O_1901,N_28763,N_29479);
nor UO_1902 (O_1902,N_29445,N_29224);
nor UO_1903 (O_1903,N_29583,N_29577);
or UO_1904 (O_1904,N_28658,N_29497);
and UO_1905 (O_1905,N_29343,N_29135);
and UO_1906 (O_1906,N_29331,N_29854);
nand UO_1907 (O_1907,N_29278,N_29630);
nand UO_1908 (O_1908,N_29754,N_29632);
nor UO_1909 (O_1909,N_29394,N_29038);
nor UO_1910 (O_1910,N_29091,N_29463);
or UO_1911 (O_1911,N_29995,N_29555);
nor UO_1912 (O_1912,N_29267,N_29080);
xnor UO_1913 (O_1913,N_29961,N_28690);
and UO_1914 (O_1914,N_29500,N_28774);
xor UO_1915 (O_1915,N_29961,N_29038);
nor UO_1916 (O_1916,N_28815,N_29207);
xor UO_1917 (O_1917,N_29001,N_29209);
nor UO_1918 (O_1918,N_29055,N_29920);
or UO_1919 (O_1919,N_29737,N_28632);
or UO_1920 (O_1920,N_28606,N_29785);
or UO_1921 (O_1921,N_28687,N_28923);
or UO_1922 (O_1922,N_29383,N_29531);
and UO_1923 (O_1923,N_29865,N_29742);
xor UO_1924 (O_1924,N_29890,N_29415);
nor UO_1925 (O_1925,N_28748,N_28887);
or UO_1926 (O_1926,N_28655,N_28562);
nand UO_1927 (O_1927,N_29680,N_29240);
xor UO_1928 (O_1928,N_28541,N_29075);
nor UO_1929 (O_1929,N_29541,N_29737);
xor UO_1930 (O_1930,N_29451,N_29213);
nand UO_1931 (O_1931,N_29942,N_29924);
nand UO_1932 (O_1932,N_28892,N_29242);
nor UO_1933 (O_1933,N_29578,N_29251);
nor UO_1934 (O_1934,N_29243,N_29234);
xnor UO_1935 (O_1935,N_28944,N_29890);
nand UO_1936 (O_1936,N_29793,N_28525);
nand UO_1937 (O_1937,N_29861,N_28664);
or UO_1938 (O_1938,N_29730,N_29477);
nand UO_1939 (O_1939,N_29134,N_29125);
xor UO_1940 (O_1940,N_28738,N_29166);
nor UO_1941 (O_1941,N_28983,N_29321);
or UO_1942 (O_1942,N_29301,N_29456);
or UO_1943 (O_1943,N_29751,N_29058);
or UO_1944 (O_1944,N_29393,N_29656);
and UO_1945 (O_1945,N_29388,N_29826);
xor UO_1946 (O_1946,N_28711,N_28895);
nor UO_1947 (O_1947,N_28591,N_28680);
and UO_1948 (O_1948,N_29064,N_29970);
xnor UO_1949 (O_1949,N_29316,N_29048);
nand UO_1950 (O_1950,N_29107,N_28808);
nor UO_1951 (O_1951,N_29781,N_29440);
nor UO_1952 (O_1952,N_29242,N_28952);
nand UO_1953 (O_1953,N_29091,N_29936);
nor UO_1954 (O_1954,N_29998,N_29824);
or UO_1955 (O_1955,N_29413,N_28632);
or UO_1956 (O_1956,N_28505,N_29069);
xor UO_1957 (O_1957,N_29919,N_29727);
nand UO_1958 (O_1958,N_29465,N_28921);
and UO_1959 (O_1959,N_28938,N_29473);
xor UO_1960 (O_1960,N_29814,N_29838);
nor UO_1961 (O_1961,N_29078,N_29798);
xor UO_1962 (O_1962,N_28637,N_29515);
nor UO_1963 (O_1963,N_28860,N_29201);
nor UO_1964 (O_1964,N_28755,N_28733);
and UO_1965 (O_1965,N_28706,N_29357);
nor UO_1966 (O_1966,N_29371,N_29275);
and UO_1967 (O_1967,N_28660,N_29338);
and UO_1968 (O_1968,N_28516,N_28770);
and UO_1969 (O_1969,N_29370,N_28959);
and UO_1970 (O_1970,N_29268,N_28940);
xnor UO_1971 (O_1971,N_29236,N_29561);
xor UO_1972 (O_1972,N_29500,N_29162);
and UO_1973 (O_1973,N_28683,N_29216);
nor UO_1974 (O_1974,N_29481,N_28888);
xor UO_1975 (O_1975,N_29534,N_28991);
nand UO_1976 (O_1976,N_29164,N_28645);
and UO_1977 (O_1977,N_28939,N_29345);
nor UO_1978 (O_1978,N_29437,N_28803);
xor UO_1979 (O_1979,N_28711,N_28532);
nor UO_1980 (O_1980,N_28992,N_29742);
and UO_1981 (O_1981,N_29183,N_29280);
and UO_1982 (O_1982,N_28623,N_29295);
nor UO_1983 (O_1983,N_29233,N_29325);
xnor UO_1984 (O_1984,N_29363,N_29297);
nand UO_1985 (O_1985,N_29642,N_28608);
nor UO_1986 (O_1986,N_29344,N_28807);
and UO_1987 (O_1987,N_29099,N_29234);
nor UO_1988 (O_1988,N_29659,N_29058);
nand UO_1989 (O_1989,N_29320,N_29152);
nor UO_1990 (O_1990,N_29016,N_29394);
or UO_1991 (O_1991,N_29940,N_29084);
and UO_1992 (O_1992,N_29514,N_28531);
nor UO_1993 (O_1993,N_28759,N_29808);
nor UO_1994 (O_1994,N_29060,N_29789);
or UO_1995 (O_1995,N_28707,N_29249);
and UO_1996 (O_1996,N_28589,N_28726);
nand UO_1997 (O_1997,N_28877,N_29539);
or UO_1998 (O_1998,N_29665,N_29982);
and UO_1999 (O_1999,N_29330,N_28619);
nor UO_2000 (O_2000,N_28706,N_28758);
nor UO_2001 (O_2001,N_29677,N_28522);
xor UO_2002 (O_2002,N_29899,N_29104);
nand UO_2003 (O_2003,N_28819,N_29788);
or UO_2004 (O_2004,N_28641,N_29277);
or UO_2005 (O_2005,N_29959,N_29970);
nor UO_2006 (O_2006,N_29227,N_28891);
and UO_2007 (O_2007,N_29417,N_29420);
nand UO_2008 (O_2008,N_29014,N_29926);
nor UO_2009 (O_2009,N_28667,N_29514);
xor UO_2010 (O_2010,N_29910,N_29160);
or UO_2011 (O_2011,N_29792,N_28750);
or UO_2012 (O_2012,N_29894,N_29951);
nor UO_2013 (O_2013,N_28875,N_28973);
and UO_2014 (O_2014,N_28765,N_29136);
xnor UO_2015 (O_2015,N_28602,N_29761);
xor UO_2016 (O_2016,N_29863,N_28662);
xor UO_2017 (O_2017,N_28664,N_29873);
xnor UO_2018 (O_2018,N_28848,N_29221);
nand UO_2019 (O_2019,N_29514,N_29364);
and UO_2020 (O_2020,N_28892,N_29834);
and UO_2021 (O_2021,N_28934,N_29739);
and UO_2022 (O_2022,N_28799,N_29067);
and UO_2023 (O_2023,N_29163,N_29819);
nand UO_2024 (O_2024,N_29231,N_29095);
nand UO_2025 (O_2025,N_28563,N_29871);
nand UO_2026 (O_2026,N_29858,N_28501);
xor UO_2027 (O_2027,N_29411,N_28588);
nor UO_2028 (O_2028,N_28649,N_29583);
nand UO_2029 (O_2029,N_28514,N_29990);
and UO_2030 (O_2030,N_29860,N_29303);
xor UO_2031 (O_2031,N_28775,N_29346);
or UO_2032 (O_2032,N_28702,N_28627);
nand UO_2033 (O_2033,N_29096,N_29316);
or UO_2034 (O_2034,N_29326,N_29433);
nand UO_2035 (O_2035,N_29823,N_29211);
nand UO_2036 (O_2036,N_29338,N_29253);
nor UO_2037 (O_2037,N_29247,N_28861);
xor UO_2038 (O_2038,N_29849,N_29064);
nand UO_2039 (O_2039,N_29566,N_29763);
nor UO_2040 (O_2040,N_29673,N_29767);
and UO_2041 (O_2041,N_29840,N_29339);
nand UO_2042 (O_2042,N_28769,N_29254);
xor UO_2043 (O_2043,N_28686,N_28673);
nand UO_2044 (O_2044,N_29307,N_28655);
and UO_2045 (O_2045,N_29878,N_28934);
nand UO_2046 (O_2046,N_29290,N_29118);
or UO_2047 (O_2047,N_29110,N_28627);
nand UO_2048 (O_2048,N_29209,N_29396);
and UO_2049 (O_2049,N_29856,N_28814);
and UO_2050 (O_2050,N_29848,N_28518);
and UO_2051 (O_2051,N_29256,N_29137);
and UO_2052 (O_2052,N_28597,N_29589);
and UO_2053 (O_2053,N_28799,N_28787);
nand UO_2054 (O_2054,N_29683,N_29217);
or UO_2055 (O_2055,N_29946,N_29992);
nand UO_2056 (O_2056,N_29534,N_29763);
nor UO_2057 (O_2057,N_29502,N_28618);
and UO_2058 (O_2058,N_29353,N_28616);
nor UO_2059 (O_2059,N_29219,N_29372);
or UO_2060 (O_2060,N_29892,N_28714);
and UO_2061 (O_2061,N_29098,N_28785);
and UO_2062 (O_2062,N_29044,N_29892);
nand UO_2063 (O_2063,N_28648,N_29305);
and UO_2064 (O_2064,N_29174,N_29142);
nand UO_2065 (O_2065,N_29664,N_29196);
and UO_2066 (O_2066,N_29847,N_29475);
and UO_2067 (O_2067,N_29345,N_28898);
nor UO_2068 (O_2068,N_28872,N_28554);
nor UO_2069 (O_2069,N_29680,N_29650);
nor UO_2070 (O_2070,N_29227,N_29029);
and UO_2071 (O_2071,N_29521,N_29018);
nand UO_2072 (O_2072,N_29220,N_28530);
nand UO_2073 (O_2073,N_28650,N_29636);
or UO_2074 (O_2074,N_28596,N_29215);
nand UO_2075 (O_2075,N_29905,N_29377);
nor UO_2076 (O_2076,N_28730,N_29829);
and UO_2077 (O_2077,N_29978,N_29240);
nor UO_2078 (O_2078,N_29909,N_29384);
nand UO_2079 (O_2079,N_28651,N_29025);
and UO_2080 (O_2080,N_28843,N_29436);
nand UO_2081 (O_2081,N_29799,N_29140);
xnor UO_2082 (O_2082,N_29959,N_29201);
and UO_2083 (O_2083,N_28856,N_29606);
and UO_2084 (O_2084,N_29576,N_29252);
nand UO_2085 (O_2085,N_29534,N_29518);
and UO_2086 (O_2086,N_29447,N_28926);
nand UO_2087 (O_2087,N_29727,N_28617);
nor UO_2088 (O_2088,N_28740,N_29897);
xor UO_2089 (O_2089,N_28731,N_28548);
xor UO_2090 (O_2090,N_29379,N_29308);
nand UO_2091 (O_2091,N_28578,N_28575);
or UO_2092 (O_2092,N_28865,N_29186);
and UO_2093 (O_2093,N_29497,N_29853);
or UO_2094 (O_2094,N_29267,N_28791);
or UO_2095 (O_2095,N_29573,N_29299);
and UO_2096 (O_2096,N_28791,N_29026);
xor UO_2097 (O_2097,N_29652,N_29991);
xor UO_2098 (O_2098,N_28544,N_29658);
nor UO_2099 (O_2099,N_29409,N_29868);
nor UO_2100 (O_2100,N_29299,N_29979);
xnor UO_2101 (O_2101,N_28614,N_29849);
nor UO_2102 (O_2102,N_29636,N_29886);
and UO_2103 (O_2103,N_29606,N_28712);
nor UO_2104 (O_2104,N_29388,N_29373);
or UO_2105 (O_2105,N_28801,N_29112);
xor UO_2106 (O_2106,N_28601,N_29522);
or UO_2107 (O_2107,N_29300,N_29916);
xnor UO_2108 (O_2108,N_29785,N_28728);
or UO_2109 (O_2109,N_29259,N_29734);
or UO_2110 (O_2110,N_29471,N_29388);
nor UO_2111 (O_2111,N_29361,N_29625);
nand UO_2112 (O_2112,N_29147,N_29587);
nand UO_2113 (O_2113,N_28762,N_29081);
xor UO_2114 (O_2114,N_29800,N_29933);
nor UO_2115 (O_2115,N_29230,N_28696);
xor UO_2116 (O_2116,N_29218,N_28676);
xnor UO_2117 (O_2117,N_28742,N_29147);
nand UO_2118 (O_2118,N_29205,N_28996);
and UO_2119 (O_2119,N_29918,N_28612);
and UO_2120 (O_2120,N_29832,N_28816);
and UO_2121 (O_2121,N_28523,N_29703);
xor UO_2122 (O_2122,N_29635,N_29796);
or UO_2123 (O_2123,N_29410,N_29980);
nand UO_2124 (O_2124,N_29764,N_29814);
and UO_2125 (O_2125,N_29296,N_29319);
nor UO_2126 (O_2126,N_29255,N_28515);
nor UO_2127 (O_2127,N_28914,N_28565);
nor UO_2128 (O_2128,N_29830,N_29346);
nand UO_2129 (O_2129,N_29538,N_29671);
nand UO_2130 (O_2130,N_29975,N_29700);
or UO_2131 (O_2131,N_28998,N_29025);
and UO_2132 (O_2132,N_28880,N_28859);
nand UO_2133 (O_2133,N_28948,N_29679);
and UO_2134 (O_2134,N_28774,N_29750);
xor UO_2135 (O_2135,N_29719,N_28598);
nor UO_2136 (O_2136,N_29283,N_28677);
nand UO_2137 (O_2137,N_28765,N_29341);
xnor UO_2138 (O_2138,N_29816,N_29273);
xor UO_2139 (O_2139,N_29137,N_28503);
xor UO_2140 (O_2140,N_28729,N_29656);
xnor UO_2141 (O_2141,N_29690,N_29438);
and UO_2142 (O_2142,N_28578,N_29769);
nand UO_2143 (O_2143,N_29889,N_28937);
nand UO_2144 (O_2144,N_29990,N_29588);
xor UO_2145 (O_2145,N_29720,N_29969);
and UO_2146 (O_2146,N_29637,N_29003);
or UO_2147 (O_2147,N_29633,N_29536);
xor UO_2148 (O_2148,N_29201,N_29044);
nor UO_2149 (O_2149,N_28515,N_28926);
nor UO_2150 (O_2150,N_29976,N_29458);
or UO_2151 (O_2151,N_28690,N_29729);
nand UO_2152 (O_2152,N_29683,N_29493);
and UO_2153 (O_2153,N_29887,N_28684);
xor UO_2154 (O_2154,N_29804,N_29033);
nand UO_2155 (O_2155,N_28979,N_29051);
nand UO_2156 (O_2156,N_29825,N_28969);
and UO_2157 (O_2157,N_29213,N_29335);
nor UO_2158 (O_2158,N_28727,N_28689);
or UO_2159 (O_2159,N_28884,N_29293);
xnor UO_2160 (O_2160,N_29081,N_28931);
nor UO_2161 (O_2161,N_29368,N_28895);
nand UO_2162 (O_2162,N_28730,N_28911);
and UO_2163 (O_2163,N_29228,N_29431);
or UO_2164 (O_2164,N_28996,N_29917);
nand UO_2165 (O_2165,N_29104,N_29865);
nor UO_2166 (O_2166,N_29545,N_28787);
nor UO_2167 (O_2167,N_29702,N_29258);
and UO_2168 (O_2168,N_28811,N_29555);
nand UO_2169 (O_2169,N_29847,N_29408);
xor UO_2170 (O_2170,N_28663,N_29148);
xor UO_2171 (O_2171,N_28747,N_28676);
nand UO_2172 (O_2172,N_29833,N_28922);
nor UO_2173 (O_2173,N_29837,N_28853);
and UO_2174 (O_2174,N_29938,N_29103);
xor UO_2175 (O_2175,N_29449,N_28908);
or UO_2176 (O_2176,N_28939,N_28571);
nor UO_2177 (O_2177,N_29585,N_29061);
nor UO_2178 (O_2178,N_29422,N_29420);
nand UO_2179 (O_2179,N_29583,N_29391);
and UO_2180 (O_2180,N_29522,N_29067);
xor UO_2181 (O_2181,N_29505,N_29122);
nor UO_2182 (O_2182,N_29086,N_29439);
and UO_2183 (O_2183,N_29780,N_29432);
or UO_2184 (O_2184,N_29365,N_29236);
nand UO_2185 (O_2185,N_28856,N_29069);
nand UO_2186 (O_2186,N_29199,N_28632);
nand UO_2187 (O_2187,N_28571,N_28757);
nand UO_2188 (O_2188,N_29814,N_29147);
nand UO_2189 (O_2189,N_29712,N_29407);
and UO_2190 (O_2190,N_28693,N_29949);
nand UO_2191 (O_2191,N_28654,N_29421);
and UO_2192 (O_2192,N_29938,N_29963);
and UO_2193 (O_2193,N_29569,N_28921);
and UO_2194 (O_2194,N_28577,N_29674);
and UO_2195 (O_2195,N_29150,N_29325);
or UO_2196 (O_2196,N_28689,N_28657);
or UO_2197 (O_2197,N_29511,N_29020);
or UO_2198 (O_2198,N_28542,N_29557);
or UO_2199 (O_2199,N_28563,N_28855);
nor UO_2200 (O_2200,N_28778,N_29894);
and UO_2201 (O_2201,N_29251,N_29046);
xnor UO_2202 (O_2202,N_29297,N_29094);
nor UO_2203 (O_2203,N_28785,N_29708);
xor UO_2204 (O_2204,N_28649,N_29725);
xnor UO_2205 (O_2205,N_29486,N_29123);
and UO_2206 (O_2206,N_29375,N_29222);
or UO_2207 (O_2207,N_29631,N_29196);
and UO_2208 (O_2208,N_29052,N_29806);
and UO_2209 (O_2209,N_29141,N_29850);
or UO_2210 (O_2210,N_28995,N_29471);
nand UO_2211 (O_2211,N_28547,N_28896);
or UO_2212 (O_2212,N_28638,N_28985);
or UO_2213 (O_2213,N_29062,N_29633);
nand UO_2214 (O_2214,N_28683,N_29983);
nor UO_2215 (O_2215,N_28703,N_29859);
nand UO_2216 (O_2216,N_29660,N_29040);
or UO_2217 (O_2217,N_29300,N_29114);
xor UO_2218 (O_2218,N_29900,N_28552);
nand UO_2219 (O_2219,N_28520,N_29425);
and UO_2220 (O_2220,N_28771,N_29553);
nor UO_2221 (O_2221,N_29802,N_28938);
or UO_2222 (O_2222,N_29270,N_29041);
or UO_2223 (O_2223,N_28825,N_29390);
xor UO_2224 (O_2224,N_29743,N_29826);
nor UO_2225 (O_2225,N_28717,N_29051);
nand UO_2226 (O_2226,N_29424,N_29750);
and UO_2227 (O_2227,N_29653,N_29224);
xor UO_2228 (O_2228,N_29483,N_29934);
and UO_2229 (O_2229,N_29109,N_29008);
nor UO_2230 (O_2230,N_28627,N_29046);
nand UO_2231 (O_2231,N_29973,N_28876);
nor UO_2232 (O_2232,N_28851,N_28821);
or UO_2233 (O_2233,N_28744,N_29789);
nor UO_2234 (O_2234,N_29337,N_28645);
or UO_2235 (O_2235,N_28653,N_29221);
or UO_2236 (O_2236,N_29286,N_28661);
or UO_2237 (O_2237,N_29848,N_29314);
nor UO_2238 (O_2238,N_28711,N_29865);
nor UO_2239 (O_2239,N_29372,N_29936);
nor UO_2240 (O_2240,N_28681,N_29836);
and UO_2241 (O_2241,N_29287,N_29903);
or UO_2242 (O_2242,N_29954,N_29512);
nor UO_2243 (O_2243,N_29767,N_29748);
or UO_2244 (O_2244,N_29485,N_29128);
xor UO_2245 (O_2245,N_28937,N_28903);
xor UO_2246 (O_2246,N_28944,N_28917);
or UO_2247 (O_2247,N_29568,N_29507);
nand UO_2248 (O_2248,N_29513,N_29577);
xnor UO_2249 (O_2249,N_28759,N_29040);
xor UO_2250 (O_2250,N_29404,N_29602);
and UO_2251 (O_2251,N_28663,N_29965);
nand UO_2252 (O_2252,N_28566,N_29034);
nand UO_2253 (O_2253,N_29341,N_28520);
or UO_2254 (O_2254,N_29922,N_29681);
and UO_2255 (O_2255,N_29351,N_29397);
nand UO_2256 (O_2256,N_29138,N_28657);
and UO_2257 (O_2257,N_29613,N_28941);
xnor UO_2258 (O_2258,N_29895,N_29734);
xnor UO_2259 (O_2259,N_29079,N_28623);
or UO_2260 (O_2260,N_29357,N_29342);
nand UO_2261 (O_2261,N_28740,N_29468);
and UO_2262 (O_2262,N_29365,N_29339);
nor UO_2263 (O_2263,N_29165,N_28604);
and UO_2264 (O_2264,N_29232,N_29758);
nor UO_2265 (O_2265,N_28897,N_29153);
nor UO_2266 (O_2266,N_29287,N_28941);
or UO_2267 (O_2267,N_29504,N_29675);
nor UO_2268 (O_2268,N_28979,N_28687);
or UO_2269 (O_2269,N_29985,N_29790);
xor UO_2270 (O_2270,N_29397,N_29806);
or UO_2271 (O_2271,N_29298,N_28559);
or UO_2272 (O_2272,N_29086,N_29923);
and UO_2273 (O_2273,N_29505,N_29746);
nor UO_2274 (O_2274,N_29632,N_29598);
xnor UO_2275 (O_2275,N_29700,N_29457);
or UO_2276 (O_2276,N_28801,N_28685);
nand UO_2277 (O_2277,N_28698,N_29669);
or UO_2278 (O_2278,N_29698,N_29263);
xor UO_2279 (O_2279,N_29456,N_28709);
nand UO_2280 (O_2280,N_29126,N_29138);
or UO_2281 (O_2281,N_29685,N_28599);
xnor UO_2282 (O_2282,N_28529,N_29099);
and UO_2283 (O_2283,N_28939,N_28875);
and UO_2284 (O_2284,N_29837,N_29435);
and UO_2285 (O_2285,N_28592,N_28710);
or UO_2286 (O_2286,N_28640,N_28865);
nand UO_2287 (O_2287,N_28991,N_28893);
xor UO_2288 (O_2288,N_29520,N_28872);
nor UO_2289 (O_2289,N_29441,N_28862);
or UO_2290 (O_2290,N_28766,N_28572);
nor UO_2291 (O_2291,N_28917,N_29497);
nand UO_2292 (O_2292,N_29107,N_29013);
xnor UO_2293 (O_2293,N_28743,N_28573);
or UO_2294 (O_2294,N_28968,N_29793);
nand UO_2295 (O_2295,N_28614,N_29826);
or UO_2296 (O_2296,N_28966,N_28589);
nor UO_2297 (O_2297,N_28790,N_28928);
or UO_2298 (O_2298,N_29731,N_29027);
nor UO_2299 (O_2299,N_29614,N_29154);
or UO_2300 (O_2300,N_28932,N_29722);
nand UO_2301 (O_2301,N_29814,N_28847);
nor UO_2302 (O_2302,N_29368,N_29817);
or UO_2303 (O_2303,N_29450,N_29006);
nor UO_2304 (O_2304,N_29674,N_28989);
nand UO_2305 (O_2305,N_29990,N_29402);
and UO_2306 (O_2306,N_28516,N_28956);
nand UO_2307 (O_2307,N_28985,N_28684);
or UO_2308 (O_2308,N_28546,N_29945);
nand UO_2309 (O_2309,N_28995,N_29655);
xor UO_2310 (O_2310,N_29337,N_29382);
nor UO_2311 (O_2311,N_28899,N_29968);
and UO_2312 (O_2312,N_29597,N_29019);
xor UO_2313 (O_2313,N_29454,N_28726);
xnor UO_2314 (O_2314,N_28764,N_29827);
nor UO_2315 (O_2315,N_29814,N_29903);
nand UO_2316 (O_2316,N_29618,N_29677);
and UO_2317 (O_2317,N_29885,N_29151);
or UO_2318 (O_2318,N_28970,N_28555);
nor UO_2319 (O_2319,N_29461,N_29054);
nor UO_2320 (O_2320,N_29191,N_29274);
nor UO_2321 (O_2321,N_29461,N_28929);
nand UO_2322 (O_2322,N_28832,N_29841);
nand UO_2323 (O_2323,N_29840,N_28948);
nand UO_2324 (O_2324,N_29719,N_28967);
xor UO_2325 (O_2325,N_29216,N_29728);
or UO_2326 (O_2326,N_28573,N_29554);
nor UO_2327 (O_2327,N_29470,N_28859);
or UO_2328 (O_2328,N_28859,N_29014);
nor UO_2329 (O_2329,N_29605,N_29808);
or UO_2330 (O_2330,N_29684,N_29794);
and UO_2331 (O_2331,N_29349,N_29884);
nor UO_2332 (O_2332,N_29471,N_29702);
or UO_2333 (O_2333,N_29912,N_29680);
xnor UO_2334 (O_2334,N_28838,N_29382);
nor UO_2335 (O_2335,N_28703,N_28788);
nand UO_2336 (O_2336,N_29473,N_28928);
xnor UO_2337 (O_2337,N_29111,N_29828);
nor UO_2338 (O_2338,N_29813,N_28885);
xnor UO_2339 (O_2339,N_29300,N_29202);
xor UO_2340 (O_2340,N_28860,N_29890);
xor UO_2341 (O_2341,N_29783,N_28727);
nor UO_2342 (O_2342,N_28922,N_28662);
or UO_2343 (O_2343,N_29726,N_28529);
nor UO_2344 (O_2344,N_28732,N_28730);
nor UO_2345 (O_2345,N_28965,N_28994);
xor UO_2346 (O_2346,N_28774,N_29944);
xnor UO_2347 (O_2347,N_29865,N_28877);
and UO_2348 (O_2348,N_29440,N_29600);
nor UO_2349 (O_2349,N_28717,N_28954);
nand UO_2350 (O_2350,N_29057,N_28821);
nor UO_2351 (O_2351,N_29801,N_28700);
and UO_2352 (O_2352,N_29030,N_28944);
and UO_2353 (O_2353,N_29006,N_29065);
xnor UO_2354 (O_2354,N_29527,N_28987);
and UO_2355 (O_2355,N_29144,N_28877);
nand UO_2356 (O_2356,N_29415,N_29868);
and UO_2357 (O_2357,N_29109,N_29537);
or UO_2358 (O_2358,N_28579,N_28916);
nor UO_2359 (O_2359,N_29228,N_28716);
nor UO_2360 (O_2360,N_29088,N_29321);
and UO_2361 (O_2361,N_29583,N_29332);
nor UO_2362 (O_2362,N_29672,N_29271);
xor UO_2363 (O_2363,N_28573,N_29473);
and UO_2364 (O_2364,N_29579,N_29855);
nor UO_2365 (O_2365,N_29184,N_28671);
xor UO_2366 (O_2366,N_29652,N_28893);
xnor UO_2367 (O_2367,N_28954,N_28688);
nand UO_2368 (O_2368,N_28535,N_29902);
xor UO_2369 (O_2369,N_29162,N_29456);
or UO_2370 (O_2370,N_29689,N_28857);
xor UO_2371 (O_2371,N_29328,N_29348);
and UO_2372 (O_2372,N_29250,N_28965);
and UO_2373 (O_2373,N_29952,N_28838);
and UO_2374 (O_2374,N_29806,N_29950);
nand UO_2375 (O_2375,N_28629,N_29236);
nor UO_2376 (O_2376,N_29277,N_28686);
or UO_2377 (O_2377,N_29522,N_29136);
xnor UO_2378 (O_2378,N_29675,N_29404);
and UO_2379 (O_2379,N_28899,N_29102);
and UO_2380 (O_2380,N_28798,N_28816);
and UO_2381 (O_2381,N_29546,N_29128);
nand UO_2382 (O_2382,N_29169,N_28625);
or UO_2383 (O_2383,N_29560,N_28994);
nor UO_2384 (O_2384,N_29060,N_29601);
or UO_2385 (O_2385,N_29779,N_29464);
nand UO_2386 (O_2386,N_29211,N_29862);
or UO_2387 (O_2387,N_29332,N_29097);
nor UO_2388 (O_2388,N_28690,N_29468);
xnor UO_2389 (O_2389,N_29766,N_28530);
xor UO_2390 (O_2390,N_28726,N_28752);
and UO_2391 (O_2391,N_29509,N_29621);
nor UO_2392 (O_2392,N_29487,N_28743);
nand UO_2393 (O_2393,N_29194,N_29529);
or UO_2394 (O_2394,N_28927,N_28608);
xor UO_2395 (O_2395,N_28538,N_28828);
or UO_2396 (O_2396,N_29638,N_29362);
or UO_2397 (O_2397,N_29139,N_29925);
nor UO_2398 (O_2398,N_29080,N_29960);
xor UO_2399 (O_2399,N_29580,N_28876);
nand UO_2400 (O_2400,N_29154,N_29508);
nand UO_2401 (O_2401,N_29282,N_29807);
and UO_2402 (O_2402,N_29056,N_28950);
xnor UO_2403 (O_2403,N_29091,N_28540);
nand UO_2404 (O_2404,N_29833,N_29702);
nor UO_2405 (O_2405,N_29937,N_29236);
xnor UO_2406 (O_2406,N_28679,N_29208);
or UO_2407 (O_2407,N_29544,N_29439);
xnor UO_2408 (O_2408,N_29732,N_29358);
xnor UO_2409 (O_2409,N_28622,N_29884);
nor UO_2410 (O_2410,N_28697,N_29449);
nor UO_2411 (O_2411,N_29621,N_29628);
or UO_2412 (O_2412,N_29538,N_29718);
nand UO_2413 (O_2413,N_29193,N_29424);
nand UO_2414 (O_2414,N_28673,N_28508);
xnor UO_2415 (O_2415,N_29393,N_28691);
or UO_2416 (O_2416,N_28801,N_29994);
nand UO_2417 (O_2417,N_29403,N_28511);
and UO_2418 (O_2418,N_29097,N_29189);
nor UO_2419 (O_2419,N_29185,N_29338);
or UO_2420 (O_2420,N_29650,N_29445);
xnor UO_2421 (O_2421,N_28809,N_29950);
or UO_2422 (O_2422,N_29975,N_29963);
nand UO_2423 (O_2423,N_29590,N_29664);
and UO_2424 (O_2424,N_28641,N_29902);
nor UO_2425 (O_2425,N_29759,N_29573);
or UO_2426 (O_2426,N_28750,N_28756);
nor UO_2427 (O_2427,N_29350,N_29562);
and UO_2428 (O_2428,N_29996,N_29276);
xor UO_2429 (O_2429,N_29888,N_29826);
or UO_2430 (O_2430,N_29921,N_29720);
or UO_2431 (O_2431,N_29488,N_29955);
nand UO_2432 (O_2432,N_29591,N_29325);
and UO_2433 (O_2433,N_29287,N_29657);
nor UO_2434 (O_2434,N_28661,N_29649);
or UO_2435 (O_2435,N_28992,N_29699);
xnor UO_2436 (O_2436,N_29069,N_29304);
nor UO_2437 (O_2437,N_29353,N_29633);
or UO_2438 (O_2438,N_29379,N_29313);
nor UO_2439 (O_2439,N_29042,N_29584);
or UO_2440 (O_2440,N_29904,N_28540);
and UO_2441 (O_2441,N_29832,N_28883);
or UO_2442 (O_2442,N_29156,N_29698);
or UO_2443 (O_2443,N_28596,N_28667);
xor UO_2444 (O_2444,N_29964,N_28925);
and UO_2445 (O_2445,N_29610,N_29141);
and UO_2446 (O_2446,N_29687,N_28584);
xor UO_2447 (O_2447,N_29697,N_28953);
nand UO_2448 (O_2448,N_29747,N_29508);
xor UO_2449 (O_2449,N_29491,N_28891);
and UO_2450 (O_2450,N_28656,N_28969);
or UO_2451 (O_2451,N_29379,N_28503);
nor UO_2452 (O_2452,N_28874,N_28589);
or UO_2453 (O_2453,N_29429,N_28840);
or UO_2454 (O_2454,N_29898,N_29008);
or UO_2455 (O_2455,N_28586,N_28810);
nor UO_2456 (O_2456,N_29072,N_28680);
and UO_2457 (O_2457,N_29477,N_28611);
xnor UO_2458 (O_2458,N_29184,N_29912);
nor UO_2459 (O_2459,N_29078,N_28656);
and UO_2460 (O_2460,N_28563,N_28653);
or UO_2461 (O_2461,N_29731,N_29522);
or UO_2462 (O_2462,N_28630,N_29874);
or UO_2463 (O_2463,N_29494,N_29890);
or UO_2464 (O_2464,N_29295,N_28974);
and UO_2465 (O_2465,N_29788,N_29630);
or UO_2466 (O_2466,N_28904,N_29678);
xnor UO_2467 (O_2467,N_28942,N_29536);
xor UO_2468 (O_2468,N_29582,N_29991);
nand UO_2469 (O_2469,N_29519,N_29377);
or UO_2470 (O_2470,N_28901,N_28717);
xor UO_2471 (O_2471,N_29051,N_29433);
nand UO_2472 (O_2472,N_29475,N_29287);
nor UO_2473 (O_2473,N_29402,N_28963);
nand UO_2474 (O_2474,N_29244,N_29143);
and UO_2475 (O_2475,N_28829,N_29008);
nor UO_2476 (O_2476,N_29609,N_29582);
or UO_2477 (O_2477,N_28698,N_29834);
and UO_2478 (O_2478,N_28506,N_29243);
nand UO_2479 (O_2479,N_29985,N_29205);
and UO_2480 (O_2480,N_29046,N_28755);
and UO_2481 (O_2481,N_29121,N_29760);
and UO_2482 (O_2482,N_28551,N_29172);
and UO_2483 (O_2483,N_28780,N_29200);
and UO_2484 (O_2484,N_28898,N_29363);
and UO_2485 (O_2485,N_29294,N_29797);
nor UO_2486 (O_2486,N_29634,N_28741);
and UO_2487 (O_2487,N_28684,N_28672);
nor UO_2488 (O_2488,N_29936,N_29296);
nand UO_2489 (O_2489,N_29413,N_28948);
nand UO_2490 (O_2490,N_29090,N_29086);
or UO_2491 (O_2491,N_28606,N_28568);
xor UO_2492 (O_2492,N_28554,N_28860);
nor UO_2493 (O_2493,N_29975,N_29741);
xor UO_2494 (O_2494,N_29218,N_29109);
or UO_2495 (O_2495,N_29189,N_28766);
and UO_2496 (O_2496,N_29841,N_28554);
nor UO_2497 (O_2497,N_29725,N_29920);
nor UO_2498 (O_2498,N_29029,N_29672);
xnor UO_2499 (O_2499,N_29306,N_28839);
xor UO_2500 (O_2500,N_28714,N_28966);
xnor UO_2501 (O_2501,N_29445,N_29077);
nand UO_2502 (O_2502,N_28810,N_29097);
and UO_2503 (O_2503,N_29554,N_29716);
xnor UO_2504 (O_2504,N_28815,N_28697);
and UO_2505 (O_2505,N_29749,N_28899);
nand UO_2506 (O_2506,N_28841,N_28759);
nor UO_2507 (O_2507,N_29739,N_29410);
nand UO_2508 (O_2508,N_29559,N_29855);
nor UO_2509 (O_2509,N_29744,N_29986);
and UO_2510 (O_2510,N_29946,N_28742);
and UO_2511 (O_2511,N_28604,N_29361);
xor UO_2512 (O_2512,N_29248,N_29812);
nor UO_2513 (O_2513,N_29124,N_29489);
nand UO_2514 (O_2514,N_28898,N_28921);
and UO_2515 (O_2515,N_28608,N_29941);
and UO_2516 (O_2516,N_28948,N_28745);
nor UO_2517 (O_2517,N_29168,N_29111);
and UO_2518 (O_2518,N_29402,N_29167);
nand UO_2519 (O_2519,N_28798,N_29130);
and UO_2520 (O_2520,N_29104,N_28618);
nand UO_2521 (O_2521,N_28553,N_29236);
and UO_2522 (O_2522,N_29085,N_29322);
xor UO_2523 (O_2523,N_29472,N_29916);
nor UO_2524 (O_2524,N_29859,N_29243);
and UO_2525 (O_2525,N_29515,N_29862);
and UO_2526 (O_2526,N_28901,N_28638);
and UO_2527 (O_2527,N_28554,N_29800);
nor UO_2528 (O_2528,N_29508,N_29373);
and UO_2529 (O_2529,N_28991,N_29082);
and UO_2530 (O_2530,N_29004,N_28626);
xor UO_2531 (O_2531,N_28537,N_29390);
nor UO_2532 (O_2532,N_28560,N_29409);
or UO_2533 (O_2533,N_28824,N_29894);
nand UO_2534 (O_2534,N_29194,N_29556);
nor UO_2535 (O_2535,N_29035,N_28829);
nor UO_2536 (O_2536,N_28808,N_29112);
xnor UO_2537 (O_2537,N_28732,N_28781);
nor UO_2538 (O_2538,N_29722,N_29907);
nor UO_2539 (O_2539,N_29889,N_29820);
xnor UO_2540 (O_2540,N_29589,N_29977);
xor UO_2541 (O_2541,N_29743,N_28531);
and UO_2542 (O_2542,N_28622,N_28741);
nand UO_2543 (O_2543,N_28883,N_29615);
and UO_2544 (O_2544,N_28575,N_29363);
xor UO_2545 (O_2545,N_29919,N_29168);
nand UO_2546 (O_2546,N_29184,N_29466);
or UO_2547 (O_2547,N_29713,N_28689);
nand UO_2548 (O_2548,N_28697,N_28633);
nand UO_2549 (O_2549,N_29427,N_28651);
xnor UO_2550 (O_2550,N_29184,N_29327);
xnor UO_2551 (O_2551,N_29884,N_28916);
or UO_2552 (O_2552,N_29068,N_29318);
nor UO_2553 (O_2553,N_29398,N_29377);
xor UO_2554 (O_2554,N_28934,N_28973);
and UO_2555 (O_2555,N_29681,N_29758);
xnor UO_2556 (O_2556,N_29829,N_29839);
and UO_2557 (O_2557,N_29407,N_29459);
nor UO_2558 (O_2558,N_29096,N_29127);
and UO_2559 (O_2559,N_28686,N_28880);
and UO_2560 (O_2560,N_29981,N_29942);
or UO_2561 (O_2561,N_28734,N_28737);
or UO_2562 (O_2562,N_28878,N_29803);
nor UO_2563 (O_2563,N_28670,N_29289);
nor UO_2564 (O_2564,N_28977,N_29816);
nor UO_2565 (O_2565,N_29773,N_29328);
nor UO_2566 (O_2566,N_29702,N_28735);
nand UO_2567 (O_2567,N_29047,N_28867);
and UO_2568 (O_2568,N_29243,N_28534);
nor UO_2569 (O_2569,N_28943,N_28725);
nor UO_2570 (O_2570,N_29741,N_29289);
nand UO_2571 (O_2571,N_28610,N_28854);
nand UO_2572 (O_2572,N_28759,N_28564);
nand UO_2573 (O_2573,N_29995,N_28748);
or UO_2574 (O_2574,N_29645,N_29649);
xor UO_2575 (O_2575,N_28702,N_28846);
nand UO_2576 (O_2576,N_28519,N_29364);
nor UO_2577 (O_2577,N_29315,N_28880);
and UO_2578 (O_2578,N_29060,N_29140);
or UO_2579 (O_2579,N_29096,N_29800);
and UO_2580 (O_2580,N_29164,N_29217);
or UO_2581 (O_2581,N_29722,N_29819);
and UO_2582 (O_2582,N_29952,N_29256);
and UO_2583 (O_2583,N_28985,N_28566);
and UO_2584 (O_2584,N_29916,N_29926);
or UO_2585 (O_2585,N_28922,N_28671);
nor UO_2586 (O_2586,N_28554,N_29649);
nand UO_2587 (O_2587,N_29110,N_29454);
xor UO_2588 (O_2588,N_29923,N_29939);
xor UO_2589 (O_2589,N_29931,N_29817);
xor UO_2590 (O_2590,N_28800,N_29546);
or UO_2591 (O_2591,N_29701,N_29813);
xor UO_2592 (O_2592,N_29842,N_28758);
and UO_2593 (O_2593,N_29365,N_29968);
and UO_2594 (O_2594,N_29890,N_28712);
nor UO_2595 (O_2595,N_29624,N_29157);
xor UO_2596 (O_2596,N_29831,N_29967);
nand UO_2597 (O_2597,N_28996,N_29995);
nor UO_2598 (O_2598,N_29824,N_28605);
nand UO_2599 (O_2599,N_28619,N_28736);
xnor UO_2600 (O_2600,N_29559,N_29999);
nor UO_2601 (O_2601,N_29722,N_29653);
nor UO_2602 (O_2602,N_29567,N_29553);
nand UO_2603 (O_2603,N_29776,N_29011);
or UO_2604 (O_2604,N_29864,N_28716);
and UO_2605 (O_2605,N_29594,N_29981);
and UO_2606 (O_2606,N_28906,N_29561);
nor UO_2607 (O_2607,N_28943,N_28607);
xnor UO_2608 (O_2608,N_28824,N_29462);
nand UO_2609 (O_2609,N_28904,N_29348);
and UO_2610 (O_2610,N_28672,N_29183);
and UO_2611 (O_2611,N_28837,N_29870);
or UO_2612 (O_2612,N_29784,N_29613);
xor UO_2613 (O_2613,N_29973,N_29970);
and UO_2614 (O_2614,N_29657,N_29455);
nor UO_2615 (O_2615,N_29637,N_29448);
nor UO_2616 (O_2616,N_29381,N_28935);
and UO_2617 (O_2617,N_29893,N_29957);
nand UO_2618 (O_2618,N_28976,N_29315);
xor UO_2619 (O_2619,N_29864,N_29444);
and UO_2620 (O_2620,N_29316,N_29500);
nand UO_2621 (O_2621,N_28622,N_29810);
nand UO_2622 (O_2622,N_29230,N_29075);
and UO_2623 (O_2623,N_29941,N_29175);
and UO_2624 (O_2624,N_29538,N_29131);
nand UO_2625 (O_2625,N_29420,N_28725);
or UO_2626 (O_2626,N_28691,N_28847);
or UO_2627 (O_2627,N_29998,N_28660);
nand UO_2628 (O_2628,N_28513,N_29471);
nor UO_2629 (O_2629,N_28718,N_28858);
or UO_2630 (O_2630,N_29424,N_29203);
nand UO_2631 (O_2631,N_29601,N_28954);
nor UO_2632 (O_2632,N_29415,N_28665);
nand UO_2633 (O_2633,N_28624,N_28906);
or UO_2634 (O_2634,N_29527,N_29764);
nor UO_2635 (O_2635,N_28649,N_29130);
nor UO_2636 (O_2636,N_29035,N_29045);
xnor UO_2637 (O_2637,N_29114,N_28679);
and UO_2638 (O_2638,N_29030,N_28765);
xor UO_2639 (O_2639,N_28710,N_29991);
and UO_2640 (O_2640,N_29821,N_29035);
nor UO_2641 (O_2641,N_29542,N_29264);
and UO_2642 (O_2642,N_29077,N_29682);
and UO_2643 (O_2643,N_29574,N_29777);
xor UO_2644 (O_2644,N_29586,N_29291);
xnor UO_2645 (O_2645,N_29622,N_28799);
nand UO_2646 (O_2646,N_29072,N_29725);
and UO_2647 (O_2647,N_28514,N_29035);
xnor UO_2648 (O_2648,N_29948,N_29320);
and UO_2649 (O_2649,N_29797,N_29109);
and UO_2650 (O_2650,N_29663,N_28979);
or UO_2651 (O_2651,N_29390,N_29215);
or UO_2652 (O_2652,N_29472,N_29717);
or UO_2653 (O_2653,N_29681,N_28524);
nand UO_2654 (O_2654,N_29123,N_29225);
nand UO_2655 (O_2655,N_28919,N_28672);
and UO_2656 (O_2656,N_29936,N_28719);
nand UO_2657 (O_2657,N_29011,N_29563);
and UO_2658 (O_2658,N_28957,N_29773);
and UO_2659 (O_2659,N_28977,N_29442);
nor UO_2660 (O_2660,N_28586,N_29049);
nor UO_2661 (O_2661,N_29662,N_29426);
xnor UO_2662 (O_2662,N_29476,N_28850);
xor UO_2663 (O_2663,N_29966,N_28613);
nand UO_2664 (O_2664,N_29604,N_29702);
nor UO_2665 (O_2665,N_29834,N_29619);
nor UO_2666 (O_2666,N_29858,N_29476);
nand UO_2667 (O_2667,N_29060,N_29632);
xor UO_2668 (O_2668,N_28905,N_29250);
and UO_2669 (O_2669,N_28939,N_28704);
xor UO_2670 (O_2670,N_29958,N_28907);
nand UO_2671 (O_2671,N_29036,N_29100);
xnor UO_2672 (O_2672,N_28581,N_29378);
xnor UO_2673 (O_2673,N_28631,N_29252);
or UO_2674 (O_2674,N_28846,N_28844);
xnor UO_2675 (O_2675,N_29044,N_29217);
nand UO_2676 (O_2676,N_29672,N_29099);
xor UO_2677 (O_2677,N_29440,N_29676);
xnor UO_2678 (O_2678,N_29395,N_28551);
nor UO_2679 (O_2679,N_29013,N_29387);
xor UO_2680 (O_2680,N_29392,N_29580);
and UO_2681 (O_2681,N_29800,N_29959);
and UO_2682 (O_2682,N_29840,N_29594);
nand UO_2683 (O_2683,N_29154,N_29661);
nand UO_2684 (O_2684,N_28726,N_29323);
or UO_2685 (O_2685,N_29549,N_28822);
and UO_2686 (O_2686,N_28914,N_28887);
nor UO_2687 (O_2687,N_29706,N_28989);
or UO_2688 (O_2688,N_28590,N_29524);
nor UO_2689 (O_2689,N_28888,N_29724);
nor UO_2690 (O_2690,N_28627,N_29290);
nor UO_2691 (O_2691,N_29925,N_28724);
and UO_2692 (O_2692,N_29532,N_29169);
and UO_2693 (O_2693,N_29801,N_29473);
nor UO_2694 (O_2694,N_29720,N_29483);
or UO_2695 (O_2695,N_29674,N_29593);
xnor UO_2696 (O_2696,N_29750,N_29246);
and UO_2697 (O_2697,N_29830,N_28527);
and UO_2698 (O_2698,N_28630,N_29767);
nand UO_2699 (O_2699,N_29713,N_28894);
xor UO_2700 (O_2700,N_29315,N_29557);
xor UO_2701 (O_2701,N_29567,N_29287);
nor UO_2702 (O_2702,N_29099,N_28890);
or UO_2703 (O_2703,N_29884,N_29421);
and UO_2704 (O_2704,N_29512,N_29770);
and UO_2705 (O_2705,N_29427,N_29805);
xor UO_2706 (O_2706,N_29484,N_29390);
or UO_2707 (O_2707,N_29622,N_29597);
nor UO_2708 (O_2708,N_28902,N_29063);
or UO_2709 (O_2709,N_28675,N_29742);
nor UO_2710 (O_2710,N_28832,N_28850);
nor UO_2711 (O_2711,N_29907,N_29535);
xor UO_2712 (O_2712,N_29321,N_28908);
or UO_2713 (O_2713,N_29817,N_29272);
and UO_2714 (O_2714,N_29637,N_28905);
and UO_2715 (O_2715,N_29217,N_28607);
nor UO_2716 (O_2716,N_28774,N_28501);
nand UO_2717 (O_2717,N_29868,N_29678);
nor UO_2718 (O_2718,N_28658,N_29524);
nand UO_2719 (O_2719,N_28881,N_28561);
nor UO_2720 (O_2720,N_29475,N_29376);
xnor UO_2721 (O_2721,N_29046,N_29604);
or UO_2722 (O_2722,N_28684,N_28910);
and UO_2723 (O_2723,N_28895,N_29506);
xor UO_2724 (O_2724,N_29483,N_29601);
nand UO_2725 (O_2725,N_29675,N_29173);
nor UO_2726 (O_2726,N_28853,N_29170);
nand UO_2727 (O_2727,N_29651,N_28639);
xnor UO_2728 (O_2728,N_29938,N_29309);
nand UO_2729 (O_2729,N_28935,N_29677);
nor UO_2730 (O_2730,N_28723,N_28699);
and UO_2731 (O_2731,N_29359,N_28662);
nand UO_2732 (O_2732,N_29552,N_28907);
xnor UO_2733 (O_2733,N_29064,N_29463);
and UO_2734 (O_2734,N_29511,N_29161);
xor UO_2735 (O_2735,N_29169,N_28948);
nand UO_2736 (O_2736,N_29979,N_29499);
and UO_2737 (O_2737,N_29404,N_29695);
xnor UO_2738 (O_2738,N_28906,N_28813);
and UO_2739 (O_2739,N_29431,N_29938);
or UO_2740 (O_2740,N_28649,N_28962);
or UO_2741 (O_2741,N_29792,N_29467);
nor UO_2742 (O_2742,N_29073,N_29169);
or UO_2743 (O_2743,N_29983,N_29132);
nor UO_2744 (O_2744,N_29117,N_28593);
nor UO_2745 (O_2745,N_29780,N_28822);
or UO_2746 (O_2746,N_29461,N_29519);
or UO_2747 (O_2747,N_28606,N_29570);
and UO_2748 (O_2748,N_28511,N_28980);
nor UO_2749 (O_2749,N_29870,N_29927);
or UO_2750 (O_2750,N_29222,N_28819);
or UO_2751 (O_2751,N_29043,N_28713);
nand UO_2752 (O_2752,N_29988,N_29028);
xnor UO_2753 (O_2753,N_28667,N_28793);
and UO_2754 (O_2754,N_29242,N_28665);
nor UO_2755 (O_2755,N_28783,N_28918);
or UO_2756 (O_2756,N_29311,N_28819);
nor UO_2757 (O_2757,N_28733,N_28518);
xor UO_2758 (O_2758,N_28944,N_29511);
nor UO_2759 (O_2759,N_29349,N_28709);
or UO_2760 (O_2760,N_29002,N_28581);
nand UO_2761 (O_2761,N_29791,N_28597);
nand UO_2762 (O_2762,N_29298,N_29735);
xnor UO_2763 (O_2763,N_28792,N_28594);
and UO_2764 (O_2764,N_28917,N_29037);
nor UO_2765 (O_2765,N_29798,N_28772);
xnor UO_2766 (O_2766,N_28515,N_29898);
and UO_2767 (O_2767,N_29701,N_29829);
and UO_2768 (O_2768,N_28874,N_28894);
and UO_2769 (O_2769,N_29093,N_29876);
nand UO_2770 (O_2770,N_28689,N_28683);
nand UO_2771 (O_2771,N_29461,N_29186);
nor UO_2772 (O_2772,N_29108,N_28572);
and UO_2773 (O_2773,N_29998,N_29612);
or UO_2774 (O_2774,N_28544,N_29690);
and UO_2775 (O_2775,N_28998,N_29618);
or UO_2776 (O_2776,N_29084,N_29238);
and UO_2777 (O_2777,N_29804,N_28807);
xor UO_2778 (O_2778,N_29122,N_29191);
xnor UO_2779 (O_2779,N_28810,N_29807);
and UO_2780 (O_2780,N_28789,N_29006);
and UO_2781 (O_2781,N_29244,N_28856);
xor UO_2782 (O_2782,N_29737,N_29586);
xnor UO_2783 (O_2783,N_29233,N_28951);
nand UO_2784 (O_2784,N_29896,N_29350);
nand UO_2785 (O_2785,N_29653,N_28720);
nor UO_2786 (O_2786,N_29326,N_29590);
nand UO_2787 (O_2787,N_28539,N_29150);
xor UO_2788 (O_2788,N_29598,N_28985);
or UO_2789 (O_2789,N_29600,N_29974);
xor UO_2790 (O_2790,N_29346,N_29988);
nand UO_2791 (O_2791,N_29656,N_29453);
and UO_2792 (O_2792,N_28509,N_28566);
xnor UO_2793 (O_2793,N_29103,N_28672);
nor UO_2794 (O_2794,N_29632,N_29897);
nor UO_2795 (O_2795,N_29587,N_28879);
nand UO_2796 (O_2796,N_29269,N_29369);
or UO_2797 (O_2797,N_29348,N_29861);
nor UO_2798 (O_2798,N_29790,N_29901);
and UO_2799 (O_2799,N_29649,N_28953);
xnor UO_2800 (O_2800,N_28526,N_29651);
and UO_2801 (O_2801,N_29446,N_28642);
nor UO_2802 (O_2802,N_29699,N_29707);
xnor UO_2803 (O_2803,N_28978,N_29952);
nor UO_2804 (O_2804,N_29369,N_29232);
and UO_2805 (O_2805,N_28878,N_29595);
nor UO_2806 (O_2806,N_29356,N_28748);
xor UO_2807 (O_2807,N_29215,N_29886);
nand UO_2808 (O_2808,N_29799,N_28562);
nor UO_2809 (O_2809,N_29140,N_29178);
nand UO_2810 (O_2810,N_29769,N_29855);
nor UO_2811 (O_2811,N_28625,N_29082);
and UO_2812 (O_2812,N_29880,N_28801);
or UO_2813 (O_2813,N_28962,N_29186);
or UO_2814 (O_2814,N_29357,N_29946);
nor UO_2815 (O_2815,N_29148,N_28818);
xnor UO_2816 (O_2816,N_29427,N_28870);
and UO_2817 (O_2817,N_29112,N_29346);
or UO_2818 (O_2818,N_29837,N_29982);
nor UO_2819 (O_2819,N_29164,N_29404);
and UO_2820 (O_2820,N_29003,N_29157);
and UO_2821 (O_2821,N_29867,N_29499);
nand UO_2822 (O_2822,N_29515,N_28711);
nand UO_2823 (O_2823,N_29298,N_29974);
or UO_2824 (O_2824,N_29689,N_29771);
or UO_2825 (O_2825,N_29716,N_28578);
and UO_2826 (O_2826,N_29128,N_28763);
and UO_2827 (O_2827,N_29351,N_29502);
nand UO_2828 (O_2828,N_28974,N_29032);
or UO_2829 (O_2829,N_29296,N_29881);
nor UO_2830 (O_2830,N_28715,N_29233);
nor UO_2831 (O_2831,N_29555,N_29874);
xor UO_2832 (O_2832,N_29139,N_28762);
nor UO_2833 (O_2833,N_28579,N_29665);
nand UO_2834 (O_2834,N_29766,N_29389);
or UO_2835 (O_2835,N_28976,N_29740);
nand UO_2836 (O_2836,N_29195,N_29586);
and UO_2837 (O_2837,N_28524,N_29075);
and UO_2838 (O_2838,N_29581,N_29248);
xnor UO_2839 (O_2839,N_28886,N_28670);
nor UO_2840 (O_2840,N_29642,N_28966);
xor UO_2841 (O_2841,N_28626,N_29774);
nor UO_2842 (O_2842,N_28571,N_28530);
xor UO_2843 (O_2843,N_28724,N_29881);
and UO_2844 (O_2844,N_28860,N_28657);
xnor UO_2845 (O_2845,N_28775,N_29949);
or UO_2846 (O_2846,N_29665,N_29227);
nor UO_2847 (O_2847,N_29657,N_28666);
nor UO_2848 (O_2848,N_29742,N_29198);
or UO_2849 (O_2849,N_28964,N_29762);
nand UO_2850 (O_2850,N_29121,N_28689);
and UO_2851 (O_2851,N_29781,N_29882);
nand UO_2852 (O_2852,N_28836,N_28915);
xor UO_2853 (O_2853,N_29755,N_29757);
or UO_2854 (O_2854,N_28539,N_28555);
or UO_2855 (O_2855,N_29024,N_28510);
nand UO_2856 (O_2856,N_29207,N_29192);
nand UO_2857 (O_2857,N_29155,N_29481);
xnor UO_2858 (O_2858,N_29458,N_29826);
or UO_2859 (O_2859,N_28512,N_28515);
nand UO_2860 (O_2860,N_29759,N_29001);
or UO_2861 (O_2861,N_29314,N_29459);
xnor UO_2862 (O_2862,N_29031,N_29420);
xor UO_2863 (O_2863,N_29060,N_29918);
nor UO_2864 (O_2864,N_29812,N_29786);
or UO_2865 (O_2865,N_29905,N_28952);
or UO_2866 (O_2866,N_28507,N_28681);
nand UO_2867 (O_2867,N_29020,N_28782);
and UO_2868 (O_2868,N_28646,N_28776);
and UO_2869 (O_2869,N_29205,N_29976);
nand UO_2870 (O_2870,N_28742,N_29376);
nand UO_2871 (O_2871,N_28614,N_29312);
or UO_2872 (O_2872,N_29027,N_28731);
nor UO_2873 (O_2873,N_28913,N_29012);
nand UO_2874 (O_2874,N_29080,N_29382);
nor UO_2875 (O_2875,N_29013,N_29881);
or UO_2876 (O_2876,N_28570,N_28562);
or UO_2877 (O_2877,N_28956,N_29065);
nor UO_2878 (O_2878,N_28609,N_28625);
and UO_2879 (O_2879,N_28657,N_29588);
nor UO_2880 (O_2880,N_29795,N_28722);
nand UO_2881 (O_2881,N_29958,N_29783);
xnor UO_2882 (O_2882,N_29249,N_29645);
or UO_2883 (O_2883,N_28925,N_29483);
xor UO_2884 (O_2884,N_28996,N_29901);
nand UO_2885 (O_2885,N_28853,N_29024);
xnor UO_2886 (O_2886,N_29477,N_29628);
and UO_2887 (O_2887,N_29771,N_28897);
nand UO_2888 (O_2888,N_28793,N_29661);
nor UO_2889 (O_2889,N_29586,N_28581);
nand UO_2890 (O_2890,N_29528,N_29855);
or UO_2891 (O_2891,N_29785,N_29684);
xor UO_2892 (O_2892,N_29044,N_28950);
and UO_2893 (O_2893,N_28892,N_28797);
nand UO_2894 (O_2894,N_28787,N_29989);
and UO_2895 (O_2895,N_28701,N_29963);
or UO_2896 (O_2896,N_29452,N_29099);
or UO_2897 (O_2897,N_29999,N_28856);
or UO_2898 (O_2898,N_29338,N_29234);
xor UO_2899 (O_2899,N_29787,N_29793);
nor UO_2900 (O_2900,N_29106,N_29472);
and UO_2901 (O_2901,N_29926,N_29671);
xnor UO_2902 (O_2902,N_29896,N_29314);
nand UO_2903 (O_2903,N_29173,N_28747);
nor UO_2904 (O_2904,N_29898,N_28765);
and UO_2905 (O_2905,N_29968,N_28954);
or UO_2906 (O_2906,N_28813,N_29763);
and UO_2907 (O_2907,N_29724,N_29593);
xor UO_2908 (O_2908,N_29908,N_29532);
xor UO_2909 (O_2909,N_29987,N_28592);
nor UO_2910 (O_2910,N_29209,N_29897);
xor UO_2911 (O_2911,N_29068,N_28763);
and UO_2912 (O_2912,N_29061,N_28901);
and UO_2913 (O_2913,N_29767,N_29965);
xor UO_2914 (O_2914,N_29350,N_29448);
or UO_2915 (O_2915,N_29211,N_28843);
or UO_2916 (O_2916,N_29130,N_29781);
and UO_2917 (O_2917,N_29284,N_29803);
xor UO_2918 (O_2918,N_29898,N_28979);
xor UO_2919 (O_2919,N_29505,N_29395);
nor UO_2920 (O_2920,N_29648,N_29564);
and UO_2921 (O_2921,N_28926,N_29846);
or UO_2922 (O_2922,N_29579,N_28956);
and UO_2923 (O_2923,N_29894,N_29140);
or UO_2924 (O_2924,N_29488,N_29724);
xor UO_2925 (O_2925,N_28663,N_28850);
xnor UO_2926 (O_2926,N_29356,N_29404);
xor UO_2927 (O_2927,N_29673,N_29458);
nor UO_2928 (O_2928,N_29697,N_28927);
or UO_2929 (O_2929,N_29874,N_28994);
xnor UO_2930 (O_2930,N_28771,N_29836);
nand UO_2931 (O_2931,N_29513,N_29428);
or UO_2932 (O_2932,N_28986,N_28747);
and UO_2933 (O_2933,N_29990,N_28954);
nor UO_2934 (O_2934,N_28826,N_29717);
nor UO_2935 (O_2935,N_28773,N_29540);
xor UO_2936 (O_2936,N_28513,N_28880);
nand UO_2937 (O_2937,N_29160,N_28588);
xnor UO_2938 (O_2938,N_29055,N_29135);
nand UO_2939 (O_2939,N_28550,N_29158);
xnor UO_2940 (O_2940,N_29999,N_28931);
nand UO_2941 (O_2941,N_29101,N_28617);
nor UO_2942 (O_2942,N_28656,N_29876);
xor UO_2943 (O_2943,N_29511,N_29010);
nor UO_2944 (O_2944,N_29752,N_29392);
or UO_2945 (O_2945,N_28983,N_29652);
or UO_2946 (O_2946,N_29274,N_29614);
xnor UO_2947 (O_2947,N_29078,N_29254);
xor UO_2948 (O_2948,N_29163,N_28551);
xor UO_2949 (O_2949,N_29684,N_28598);
and UO_2950 (O_2950,N_29431,N_28906);
or UO_2951 (O_2951,N_29626,N_28622);
nand UO_2952 (O_2952,N_28846,N_29439);
xnor UO_2953 (O_2953,N_29193,N_28752);
or UO_2954 (O_2954,N_29503,N_28894);
or UO_2955 (O_2955,N_29958,N_29281);
or UO_2956 (O_2956,N_29921,N_29346);
nor UO_2957 (O_2957,N_29177,N_28740);
or UO_2958 (O_2958,N_29147,N_28726);
nor UO_2959 (O_2959,N_29932,N_29306);
nor UO_2960 (O_2960,N_29059,N_29580);
xnor UO_2961 (O_2961,N_29869,N_29943);
or UO_2962 (O_2962,N_29241,N_28968);
or UO_2963 (O_2963,N_28880,N_29798);
nand UO_2964 (O_2964,N_28988,N_29816);
nand UO_2965 (O_2965,N_29823,N_29220);
xnor UO_2966 (O_2966,N_28827,N_28965);
xor UO_2967 (O_2967,N_29260,N_28700);
xnor UO_2968 (O_2968,N_29690,N_28712);
nand UO_2969 (O_2969,N_29241,N_28804);
nor UO_2970 (O_2970,N_29728,N_29850);
and UO_2971 (O_2971,N_28809,N_28507);
nand UO_2972 (O_2972,N_29142,N_29657);
or UO_2973 (O_2973,N_29427,N_29042);
nand UO_2974 (O_2974,N_29485,N_29388);
xnor UO_2975 (O_2975,N_28573,N_29979);
or UO_2976 (O_2976,N_29151,N_29749);
nand UO_2977 (O_2977,N_28537,N_29157);
nor UO_2978 (O_2978,N_29129,N_29626);
nor UO_2979 (O_2979,N_28641,N_29241);
xor UO_2980 (O_2980,N_28549,N_28694);
nand UO_2981 (O_2981,N_28717,N_28639);
nor UO_2982 (O_2982,N_29403,N_29459);
and UO_2983 (O_2983,N_29234,N_29880);
xnor UO_2984 (O_2984,N_29541,N_28891);
xor UO_2985 (O_2985,N_29615,N_29099);
and UO_2986 (O_2986,N_28507,N_28501);
or UO_2987 (O_2987,N_29970,N_29074);
xnor UO_2988 (O_2988,N_28662,N_28565);
nand UO_2989 (O_2989,N_28514,N_29596);
or UO_2990 (O_2990,N_28802,N_29384);
nand UO_2991 (O_2991,N_29863,N_29387);
nand UO_2992 (O_2992,N_29554,N_29854);
nand UO_2993 (O_2993,N_29215,N_28641);
nand UO_2994 (O_2994,N_28787,N_28547);
nand UO_2995 (O_2995,N_29828,N_29321);
and UO_2996 (O_2996,N_28570,N_29385);
or UO_2997 (O_2997,N_28851,N_29457);
nand UO_2998 (O_2998,N_29220,N_29747);
nand UO_2999 (O_2999,N_29237,N_29571);
or UO_3000 (O_3000,N_29168,N_29467);
or UO_3001 (O_3001,N_29700,N_29777);
nand UO_3002 (O_3002,N_29677,N_29430);
xnor UO_3003 (O_3003,N_28989,N_28793);
nand UO_3004 (O_3004,N_28806,N_29006);
nand UO_3005 (O_3005,N_28849,N_29889);
or UO_3006 (O_3006,N_29338,N_28905);
xor UO_3007 (O_3007,N_29919,N_28775);
nand UO_3008 (O_3008,N_29959,N_29407);
nor UO_3009 (O_3009,N_29180,N_29728);
nor UO_3010 (O_3010,N_29425,N_29364);
or UO_3011 (O_3011,N_29011,N_28681);
nand UO_3012 (O_3012,N_28804,N_29963);
or UO_3013 (O_3013,N_28996,N_29434);
or UO_3014 (O_3014,N_29157,N_29136);
or UO_3015 (O_3015,N_28912,N_29926);
xnor UO_3016 (O_3016,N_29223,N_28867);
nand UO_3017 (O_3017,N_28836,N_28549);
nand UO_3018 (O_3018,N_29717,N_29324);
nand UO_3019 (O_3019,N_29296,N_29605);
xor UO_3020 (O_3020,N_29715,N_29911);
xor UO_3021 (O_3021,N_29412,N_28695);
nor UO_3022 (O_3022,N_29162,N_29455);
nand UO_3023 (O_3023,N_28784,N_29915);
nor UO_3024 (O_3024,N_29394,N_29415);
nand UO_3025 (O_3025,N_29430,N_28539);
or UO_3026 (O_3026,N_28696,N_28786);
and UO_3027 (O_3027,N_28794,N_29931);
or UO_3028 (O_3028,N_28654,N_29588);
and UO_3029 (O_3029,N_29432,N_29469);
or UO_3030 (O_3030,N_28987,N_29546);
and UO_3031 (O_3031,N_28535,N_29307);
and UO_3032 (O_3032,N_29268,N_29558);
xnor UO_3033 (O_3033,N_29116,N_28918);
nand UO_3034 (O_3034,N_28929,N_29466);
xnor UO_3035 (O_3035,N_29025,N_29118);
nor UO_3036 (O_3036,N_29070,N_29061);
nand UO_3037 (O_3037,N_29653,N_29901);
and UO_3038 (O_3038,N_29173,N_29538);
or UO_3039 (O_3039,N_28636,N_29197);
nand UO_3040 (O_3040,N_28522,N_28854);
xnor UO_3041 (O_3041,N_29923,N_29916);
nor UO_3042 (O_3042,N_29700,N_29913);
xor UO_3043 (O_3043,N_29299,N_29243);
nor UO_3044 (O_3044,N_29733,N_28876);
or UO_3045 (O_3045,N_28614,N_29059);
xnor UO_3046 (O_3046,N_29573,N_29231);
nor UO_3047 (O_3047,N_29085,N_29359);
nor UO_3048 (O_3048,N_29999,N_28967);
xor UO_3049 (O_3049,N_28891,N_28821);
nand UO_3050 (O_3050,N_29552,N_28910);
or UO_3051 (O_3051,N_29537,N_29152);
nand UO_3052 (O_3052,N_29784,N_29975);
or UO_3053 (O_3053,N_28894,N_29516);
xor UO_3054 (O_3054,N_29710,N_29337);
nand UO_3055 (O_3055,N_29033,N_28859);
or UO_3056 (O_3056,N_28961,N_28927);
nand UO_3057 (O_3057,N_29296,N_29018);
xor UO_3058 (O_3058,N_29530,N_29381);
nor UO_3059 (O_3059,N_29735,N_29687);
nand UO_3060 (O_3060,N_29361,N_28664);
nand UO_3061 (O_3061,N_28564,N_29113);
xor UO_3062 (O_3062,N_29302,N_29603);
nor UO_3063 (O_3063,N_29054,N_29251);
and UO_3064 (O_3064,N_29599,N_28759);
nor UO_3065 (O_3065,N_29258,N_29519);
and UO_3066 (O_3066,N_29966,N_29538);
nor UO_3067 (O_3067,N_29307,N_28923);
xor UO_3068 (O_3068,N_29579,N_28583);
or UO_3069 (O_3069,N_29049,N_29343);
and UO_3070 (O_3070,N_28733,N_29536);
nor UO_3071 (O_3071,N_28540,N_29401);
nor UO_3072 (O_3072,N_29274,N_29163);
nor UO_3073 (O_3073,N_28716,N_28949);
or UO_3074 (O_3074,N_29125,N_28993);
or UO_3075 (O_3075,N_29300,N_29729);
xnor UO_3076 (O_3076,N_29261,N_29388);
xnor UO_3077 (O_3077,N_29866,N_28507);
xnor UO_3078 (O_3078,N_29267,N_29749);
xnor UO_3079 (O_3079,N_29545,N_29976);
and UO_3080 (O_3080,N_28514,N_29586);
and UO_3081 (O_3081,N_29312,N_29652);
nand UO_3082 (O_3082,N_28517,N_28996);
xor UO_3083 (O_3083,N_28768,N_28895);
and UO_3084 (O_3084,N_28672,N_29477);
or UO_3085 (O_3085,N_29234,N_29156);
or UO_3086 (O_3086,N_29067,N_29901);
xnor UO_3087 (O_3087,N_29975,N_29427);
and UO_3088 (O_3088,N_29756,N_29281);
xnor UO_3089 (O_3089,N_28955,N_29278);
or UO_3090 (O_3090,N_29882,N_29213);
xnor UO_3091 (O_3091,N_28828,N_29671);
xnor UO_3092 (O_3092,N_29596,N_29431);
or UO_3093 (O_3093,N_29010,N_29618);
nor UO_3094 (O_3094,N_28677,N_28534);
and UO_3095 (O_3095,N_29340,N_29352);
or UO_3096 (O_3096,N_29797,N_29220);
and UO_3097 (O_3097,N_29869,N_29279);
xor UO_3098 (O_3098,N_29602,N_28991);
or UO_3099 (O_3099,N_28567,N_29208);
nand UO_3100 (O_3100,N_29356,N_29246);
and UO_3101 (O_3101,N_29061,N_28957);
nand UO_3102 (O_3102,N_28964,N_29848);
and UO_3103 (O_3103,N_28868,N_29736);
or UO_3104 (O_3104,N_28938,N_28575);
and UO_3105 (O_3105,N_29702,N_29067);
nand UO_3106 (O_3106,N_29865,N_28995);
or UO_3107 (O_3107,N_29726,N_28623);
nand UO_3108 (O_3108,N_28913,N_29220);
nor UO_3109 (O_3109,N_29318,N_28687);
xor UO_3110 (O_3110,N_29226,N_28507);
nor UO_3111 (O_3111,N_29823,N_28810);
and UO_3112 (O_3112,N_29124,N_29673);
and UO_3113 (O_3113,N_29669,N_29235);
or UO_3114 (O_3114,N_28788,N_29478);
or UO_3115 (O_3115,N_28784,N_28559);
and UO_3116 (O_3116,N_29550,N_28774);
and UO_3117 (O_3117,N_29099,N_28638);
nor UO_3118 (O_3118,N_29761,N_28959);
nor UO_3119 (O_3119,N_28776,N_29050);
or UO_3120 (O_3120,N_28538,N_29671);
nor UO_3121 (O_3121,N_28798,N_29853);
xnor UO_3122 (O_3122,N_29491,N_29727);
xnor UO_3123 (O_3123,N_29542,N_28668);
xor UO_3124 (O_3124,N_29962,N_29277);
and UO_3125 (O_3125,N_28796,N_29355);
or UO_3126 (O_3126,N_29159,N_28978);
nand UO_3127 (O_3127,N_28983,N_28798);
and UO_3128 (O_3128,N_28802,N_29589);
xor UO_3129 (O_3129,N_28807,N_29385);
and UO_3130 (O_3130,N_29333,N_28846);
and UO_3131 (O_3131,N_29293,N_28509);
or UO_3132 (O_3132,N_29829,N_28808);
xor UO_3133 (O_3133,N_28960,N_29035);
or UO_3134 (O_3134,N_28848,N_29611);
or UO_3135 (O_3135,N_29297,N_29739);
nor UO_3136 (O_3136,N_28836,N_28738);
or UO_3137 (O_3137,N_29466,N_28931);
and UO_3138 (O_3138,N_29766,N_28736);
xor UO_3139 (O_3139,N_28623,N_29265);
nor UO_3140 (O_3140,N_29594,N_28895);
nor UO_3141 (O_3141,N_29581,N_28501);
xor UO_3142 (O_3142,N_29031,N_29116);
or UO_3143 (O_3143,N_29241,N_29143);
and UO_3144 (O_3144,N_29364,N_28503);
nor UO_3145 (O_3145,N_29039,N_29609);
xor UO_3146 (O_3146,N_28550,N_29393);
and UO_3147 (O_3147,N_28847,N_29502);
or UO_3148 (O_3148,N_28704,N_29312);
or UO_3149 (O_3149,N_28696,N_29582);
nand UO_3150 (O_3150,N_29971,N_29412);
nand UO_3151 (O_3151,N_29386,N_29018);
nor UO_3152 (O_3152,N_29855,N_29693);
nand UO_3153 (O_3153,N_29349,N_29522);
or UO_3154 (O_3154,N_29748,N_29995);
xor UO_3155 (O_3155,N_29710,N_29920);
xnor UO_3156 (O_3156,N_29249,N_29936);
xnor UO_3157 (O_3157,N_29834,N_29511);
or UO_3158 (O_3158,N_29019,N_28826);
xor UO_3159 (O_3159,N_29222,N_28617);
nand UO_3160 (O_3160,N_28658,N_29197);
xor UO_3161 (O_3161,N_28878,N_29550);
nand UO_3162 (O_3162,N_29196,N_28559);
nand UO_3163 (O_3163,N_29634,N_28537);
xnor UO_3164 (O_3164,N_28665,N_28857);
xor UO_3165 (O_3165,N_29186,N_29439);
nand UO_3166 (O_3166,N_28896,N_28600);
nor UO_3167 (O_3167,N_28619,N_29461);
nand UO_3168 (O_3168,N_29607,N_29307);
nor UO_3169 (O_3169,N_28961,N_29120);
or UO_3170 (O_3170,N_29623,N_29735);
and UO_3171 (O_3171,N_29702,N_28889);
or UO_3172 (O_3172,N_28569,N_28832);
nand UO_3173 (O_3173,N_28633,N_28878);
or UO_3174 (O_3174,N_29580,N_29411);
or UO_3175 (O_3175,N_28732,N_29563);
or UO_3176 (O_3176,N_29708,N_29996);
or UO_3177 (O_3177,N_28668,N_28976);
xor UO_3178 (O_3178,N_29231,N_29023);
or UO_3179 (O_3179,N_29130,N_29394);
xnor UO_3180 (O_3180,N_28542,N_29618);
nor UO_3181 (O_3181,N_29465,N_29594);
and UO_3182 (O_3182,N_29520,N_28863);
nand UO_3183 (O_3183,N_29555,N_28988);
and UO_3184 (O_3184,N_29551,N_29973);
and UO_3185 (O_3185,N_29218,N_28865);
or UO_3186 (O_3186,N_29207,N_29440);
and UO_3187 (O_3187,N_29695,N_29060);
and UO_3188 (O_3188,N_28973,N_29393);
and UO_3189 (O_3189,N_29447,N_29560);
or UO_3190 (O_3190,N_29983,N_29882);
and UO_3191 (O_3191,N_29500,N_28503);
nand UO_3192 (O_3192,N_28611,N_28873);
nand UO_3193 (O_3193,N_29995,N_28765);
and UO_3194 (O_3194,N_29747,N_29746);
and UO_3195 (O_3195,N_29737,N_28738);
or UO_3196 (O_3196,N_29803,N_28983);
nor UO_3197 (O_3197,N_29057,N_29258);
or UO_3198 (O_3198,N_29851,N_29092);
nor UO_3199 (O_3199,N_29135,N_29151);
or UO_3200 (O_3200,N_29585,N_29793);
xor UO_3201 (O_3201,N_29247,N_28986);
nor UO_3202 (O_3202,N_28612,N_28797);
nor UO_3203 (O_3203,N_29387,N_29276);
or UO_3204 (O_3204,N_29811,N_28860);
nor UO_3205 (O_3205,N_28791,N_28872);
or UO_3206 (O_3206,N_29738,N_29922);
or UO_3207 (O_3207,N_28519,N_28762);
xnor UO_3208 (O_3208,N_29412,N_29947);
or UO_3209 (O_3209,N_28774,N_29483);
and UO_3210 (O_3210,N_29629,N_29015);
nand UO_3211 (O_3211,N_29822,N_29766);
nor UO_3212 (O_3212,N_29714,N_28590);
or UO_3213 (O_3213,N_29137,N_29299);
xor UO_3214 (O_3214,N_28534,N_29004);
or UO_3215 (O_3215,N_29061,N_28625);
nand UO_3216 (O_3216,N_28678,N_29312);
xnor UO_3217 (O_3217,N_29137,N_29158);
or UO_3218 (O_3218,N_29276,N_29954);
nand UO_3219 (O_3219,N_29500,N_29566);
or UO_3220 (O_3220,N_29083,N_29145);
xnor UO_3221 (O_3221,N_29766,N_29048);
and UO_3222 (O_3222,N_29620,N_29187);
xnor UO_3223 (O_3223,N_29844,N_29926);
xnor UO_3224 (O_3224,N_29479,N_29322);
xor UO_3225 (O_3225,N_29583,N_28877);
nor UO_3226 (O_3226,N_29802,N_29970);
nand UO_3227 (O_3227,N_28667,N_29382);
and UO_3228 (O_3228,N_28625,N_29411);
xor UO_3229 (O_3229,N_29222,N_29878);
nand UO_3230 (O_3230,N_29281,N_29336);
or UO_3231 (O_3231,N_29777,N_29116);
nor UO_3232 (O_3232,N_29440,N_28884);
xnor UO_3233 (O_3233,N_28759,N_28796);
xnor UO_3234 (O_3234,N_29296,N_28672);
and UO_3235 (O_3235,N_28856,N_29942);
and UO_3236 (O_3236,N_29098,N_29994);
and UO_3237 (O_3237,N_28531,N_29715);
or UO_3238 (O_3238,N_28626,N_29464);
or UO_3239 (O_3239,N_28622,N_29687);
and UO_3240 (O_3240,N_29723,N_28885);
xnor UO_3241 (O_3241,N_28800,N_29832);
or UO_3242 (O_3242,N_28870,N_29006);
or UO_3243 (O_3243,N_28567,N_29579);
or UO_3244 (O_3244,N_29303,N_28776);
and UO_3245 (O_3245,N_29173,N_29483);
and UO_3246 (O_3246,N_29840,N_28935);
or UO_3247 (O_3247,N_29042,N_28775);
or UO_3248 (O_3248,N_29548,N_28698);
and UO_3249 (O_3249,N_29820,N_28663);
xnor UO_3250 (O_3250,N_28866,N_29007);
xor UO_3251 (O_3251,N_29410,N_28906);
nand UO_3252 (O_3252,N_28845,N_28607);
nand UO_3253 (O_3253,N_29948,N_29973);
and UO_3254 (O_3254,N_29675,N_29535);
nor UO_3255 (O_3255,N_28697,N_28671);
nand UO_3256 (O_3256,N_29043,N_29966);
nor UO_3257 (O_3257,N_28868,N_29396);
nor UO_3258 (O_3258,N_28681,N_29377);
nor UO_3259 (O_3259,N_29593,N_28851);
and UO_3260 (O_3260,N_29827,N_29709);
nor UO_3261 (O_3261,N_29348,N_29178);
and UO_3262 (O_3262,N_28738,N_28859);
or UO_3263 (O_3263,N_29153,N_29828);
xor UO_3264 (O_3264,N_29438,N_28566);
xor UO_3265 (O_3265,N_28700,N_29736);
or UO_3266 (O_3266,N_29031,N_29319);
nor UO_3267 (O_3267,N_29808,N_28659);
or UO_3268 (O_3268,N_29750,N_29998);
and UO_3269 (O_3269,N_29745,N_29550);
and UO_3270 (O_3270,N_29672,N_29252);
nor UO_3271 (O_3271,N_29873,N_29591);
and UO_3272 (O_3272,N_29249,N_29479);
nor UO_3273 (O_3273,N_28958,N_29650);
or UO_3274 (O_3274,N_29327,N_28910);
nor UO_3275 (O_3275,N_28640,N_29731);
nor UO_3276 (O_3276,N_29750,N_29603);
nor UO_3277 (O_3277,N_28993,N_28714);
xnor UO_3278 (O_3278,N_29293,N_29579);
xnor UO_3279 (O_3279,N_29221,N_29715);
nor UO_3280 (O_3280,N_28857,N_28828);
xor UO_3281 (O_3281,N_28682,N_29710);
nor UO_3282 (O_3282,N_28989,N_28788);
xnor UO_3283 (O_3283,N_29261,N_29219);
nand UO_3284 (O_3284,N_29284,N_29175);
or UO_3285 (O_3285,N_29915,N_29852);
xor UO_3286 (O_3286,N_29862,N_28931);
nand UO_3287 (O_3287,N_29642,N_29137);
xor UO_3288 (O_3288,N_29815,N_29458);
or UO_3289 (O_3289,N_28626,N_29368);
nor UO_3290 (O_3290,N_28522,N_29683);
nor UO_3291 (O_3291,N_29563,N_28955);
nor UO_3292 (O_3292,N_29625,N_29460);
or UO_3293 (O_3293,N_29774,N_29766);
and UO_3294 (O_3294,N_28955,N_29684);
nor UO_3295 (O_3295,N_28884,N_29868);
nand UO_3296 (O_3296,N_28541,N_28689);
and UO_3297 (O_3297,N_29065,N_29817);
nand UO_3298 (O_3298,N_29958,N_29156);
and UO_3299 (O_3299,N_28589,N_28974);
and UO_3300 (O_3300,N_28674,N_28615);
and UO_3301 (O_3301,N_28706,N_29987);
nor UO_3302 (O_3302,N_28594,N_28505);
nand UO_3303 (O_3303,N_29826,N_29309);
nor UO_3304 (O_3304,N_29347,N_28781);
nor UO_3305 (O_3305,N_28509,N_29585);
xor UO_3306 (O_3306,N_29417,N_28724);
and UO_3307 (O_3307,N_29795,N_29225);
or UO_3308 (O_3308,N_29853,N_29487);
and UO_3309 (O_3309,N_29596,N_28709);
nor UO_3310 (O_3310,N_29281,N_29876);
and UO_3311 (O_3311,N_28544,N_29130);
xor UO_3312 (O_3312,N_29073,N_28720);
or UO_3313 (O_3313,N_29911,N_29747);
nand UO_3314 (O_3314,N_28752,N_29476);
nor UO_3315 (O_3315,N_29480,N_29092);
or UO_3316 (O_3316,N_29002,N_29096);
nand UO_3317 (O_3317,N_29137,N_28729);
and UO_3318 (O_3318,N_29810,N_28664);
xor UO_3319 (O_3319,N_29567,N_29562);
or UO_3320 (O_3320,N_29117,N_29939);
or UO_3321 (O_3321,N_29230,N_29225);
nor UO_3322 (O_3322,N_29210,N_29114);
nor UO_3323 (O_3323,N_29798,N_29204);
nor UO_3324 (O_3324,N_29880,N_28710);
or UO_3325 (O_3325,N_28631,N_29536);
nor UO_3326 (O_3326,N_29672,N_29946);
nor UO_3327 (O_3327,N_28547,N_28833);
and UO_3328 (O_3328,N_29974,N_29018);
or UO_3329 (O_3329,N_29103,N_29999);
xnor UO_3330 (O_3330,N_28935,N_29366);
or UO_3331 (O_3331,N_29807,N_28862);
or UO_3332 (O_3332,N_29374,N_29269);
nand UO_3333 (O_3333,N_29967,N_29655);
nand UO_3334 (O_3334,N_29404,N_28892);
nor UO_3335 (O_3335,N_29605,N_28594);
and UO_3336 (O_3336,N_29147,N_28689);
and UO_3337 (O_3337,N_29240,N_29575);
nor UO_3338 (O_3338,N_28969,N_29584);
and UO_3339 (O_3339,N_28991,N_28929);
or UO_3340 (O_3340,N_29601,N_29002);
and UO_3341 (O_3341,N_29364,N_28687);
nand UO_3342 (O_3342,N_29522,N_29157);
or UO_3343 (O_3343,N_29147,N_29108);
nor UO_3344 (O_3344,N_29319,N_29539);
or UO_3345 (O_3345,N_28538,N_29199);
or UO_3346 (O_3346,N_28941,N_29691);
nand UO_3347 (O_3347,N_28872,N_28895);
or UO_3348 (O_3348,N_28856,N_29032);
or UO_3349 (O_3349,N_28686,N_29965);
or UO_3350 (O_3350,N_29122,N_29239);
nor UO_3351 (O_3351,N_28785,N_29912);
or UO_3352 (O_3352,N_29588,N_29802);
xnor UO_3353 (O_3353,N_29135,N_29738);
xor UO_3354 (O_3354,N_28550,N_28662);
nor UO_3355 (O_3355,N_28536,N_29409);
nand UO_3356 (O_3356,N_28598,N_29537);
or UO_3357 (O_3357,N_29742,N_29756);
and UO_3358 (O_3358,N_28816,N_28802);
and UO_3359 (O_3359,N_28963,N_29337);
and UO_3360 (O_3360,N_28952,N_28613);
nand UO_3361 (O_3361,N_29448,N_29220);
or UO_3362 (O_3362,N_28732,N_28562);
nor UO_3363 (O_3363,N_29782,N_29699);
nand UO_3364 (O_3364,N_29770,N_28904);
or UO_3365 (O_3365,N_29227,N_28959);
or UO_3366 (O_3366,N_28536,N_29594);
nand UO_3367 (O_3367,N_29575,N_29536);
or UO_3368 (O_3368,N_28869,N_28523);
and UO_3369 (O_3369,N_29762,N_29431);
nor UO_3370 (O_3370,N_29738,N_29277);
or UO_3371 (O_3371,N_29702,N_29560);
nand UO_3372 (O_3372,N_28531,N_29159);
or UO_3373 (O_3373,N_29908,N_28716);
and UO_3374 (O_3374,N_28545,N_28546);
and UO_3375 (O_3375,N_28673,N_29640);
or UO_3376 (O_3376,N_29448,N_29263);
xnor UO_3377 (O_3377,N_29659,N_28674);
nand UO_3378 (O_3378,N_29390,N_28883);
nand UO_3379 (O_3379,N_29357,N_28563);
xor UO_3380 (O_3380,N_29082,N_29891);
or UO_3381 (O_3381,N_29513,N_29341);
nand UO_3382 (O_3382,N_29866,N_29519);
xor UO_3383 (O_3383,N_29285,N_28758);
and UO_3384 (O_3384,N_28505,N_28871);
nand UO_3385 (O_3385,N_29443,N_29942);
or UO_3386 (O_3386,N_28962,N_28539);
or UO_3387 (O_3387,N_29386,N_28831);
nand UO_3388 (O_3388,N_28947,N_29171);
or UO_3389 (O_3389,N_29878,N_28677);
nor UO_3390 (O_3390,N_29138,N_28771);
nor UO_3391 (O_3391,N_29981,N_29405);
xnor UO_3392 (O_3392,N_29871,N_29372);
and UO_3393 (O_3393,N_29396,N_29960);
and UO_3394 (O_3394,N_29886,N_28933);
xnor UO_3395 (O_3395,N_28875,N_28502);
or UO_3396 (O_3396,N_29191,N_29150);
and UO_3397 (O_3397,N_29737,N_28582);
nor UO_3398 (O_3398,N_29178,N_29134);
nor UO_3399 (O_3399,N_29073,N_29257);
or UO_3400 (O_3400,N_29304,N_28624);
nor UO_3401 (O_3401,N_28567,N_28535);
nand UO_3402 (O_3402,N_29968,N_29066);
nor UO_3403 (O_3403,N_29734,N_29614);
nor UO_3404 (O_3404,N_28848,N_28774);
xor UO_3405 (O_3405,N_29024,N_28680);
nor UO_3406 (O_3406,N_29519,N_28788);
nor UO_3407 (O_3407,N_29747,N_29129);
and UO_3408 (O_3408,N_29220,N_29922);
nand UO_3409 (O_3409,N_29408,N_29459);
xnor UO_3410 (O_3410,N_29734,N_29398);
xor UO_3411 (O_3411,N_29126,N_29793);
or UO_3412 (O_3412,N_29084,N_28554);
nand UO_3413 (O_3413,N_29809,N_28989);
and UO_3414 (O_3414,N_29499,N_28533);
and UO_3415 (O_3415,N_29172,N_29957);
nand UO_3416 (O_3416,N_29366,N_28844);
xnor UO_3417 (O_3417,N_29910,N_29547);
nor UO_3418 (O_3418,N_29104,N_28646);
nor UO_3419 (O_3419,N_29265,N_28548);
nor UO_3420 (O_3420,N_29960,N_29931);
nor UO_3421 (O_3421,N_28865,N_29009);
and UO_3422 (O_3422,N_29703,N_29679);
xnor UO_3423 (O_3423,N_28547,N_28729);
nand UO_3424 (O_3424,N_29254,N_29163);
and UO_3425 (O_3425,N_29491,N_28828);
and UO_3426 (O_3426,N_29749,N_29651);
and UO_3427 (O_3427,N_28930,N_29228);
or UO_3428 (O_3428,N_29244,N_29992);
nor UO_3429 (O_3429,N_29180,N_29220);
nand UO_3430 (O_3430,N_28602,N_29874);
and UO_3431 (O_3431,N_29467,N_29103);
and UO_3432 (O_3432,N_28833,N_29517);
and UO_3433 (O_3433,N_29647,N_28611);
and UO_3434 (O_3434,N_29738,N_29980);
nand UO_3435 (O_3435,N_28789,N_29511);
or UO_3436 (O_3436,N_28553,N_29671);
nor UO_3437 (O_3437,N_29460,N_28561);
and UO_3438 (O_3438,N_29575,N_29713);
xor UO_3439 (O_3439,N_29827,N_29998);
or UO_3440 (O_3440,N_28606,N_29750);
nand UO_3441 (O_3441,N_28955,N_29704);
xnor UO_3442 (O_3442,N_29787,N_29022);
nor UO_3443 (O_3443,N_28532,N_29333);
xnor UO_3444 (O_3444,N_29105,N_28676);
and UO_3445 (O_3445,N_29932,N_29972);
or UO_3446 (O_3446,N_29400,N_29262);
or UO_3447 (O_3447,N_28750,N_29860);
xnor UO_3448 (O_3448,N_29506,N_29969);
xor UO_3449 (O_3449,N_29137,N_28900);
and UO_3450 (O_3450,N_28648,N_29038);
nand UO_3451 (O_3451,N_29386,N_29498);
xnor UO_3452 (O_3452,N_29735,N_28832);
and UO_3453 (O_3453,N_29125,N_28989);
xor UO_3454 (O_3454,N_29759,N_29243);
and UO_3455 (O_3455,N_28976,N_29278);
xnor UO_3456 (O_3456,N_29324,N_28982);
nor UO_3457 (O_3457,N_28785,N_29308);
and UO_3458 (O_3458,N_28929,N_28619);
nand UO_3459 (O_3459,N_29237,N_29039);
and UO_3460 (O_3460,N_29753,N_29985);
xnor UO_3461 (O_3461,N_28501,N_29632);
xnor UO_3462 (O_3462,N_29820,N_29291);
xor UO_3463 (O_3463,N_29240,N_29712);
nor UO_3464 (O_3464,N_29283,N_29793);
nor UO_3465 (O_3465,N_28532,N_28832);
nor UO_3466 (O_3466,N_28615,N_29156);
nand UO_3467 (O_3467,N_29801,N_28681);
xnor UO_3468 (O_3468,N_29017,N_29682);
nand UO_3469 (O_3469,N_29554,N_29368);
or UO_3470 (O_3470,N_28695,N_28867);
xor UO_3471 (O_3471,N_29669,N_29314);
or UO_3472 (O_3472,N_29088,N_29130);
or UO_3473 (O_3473,N_29174,N_29334);
or UO_3474 (O_3474,N_29411,N_29124);
or UO_3475 (O_3475,N_29940,N_29777);
xor UO_3476 (O_3476,N_29240,N_29817);
nand UO_3477 (O_3477,N_29963,N_29081);
xnor UO_3478 (O_3478,N_29675,N_29068);
nor UO_3479 (O_3479,N_29249,N_29375);
or UO_3480 (O_3480,N_29192,N_29166);
nand UO_3481 (O_3481,N_29189,N_28727);
nor UO_3482 (O_3482,N_29607,N_29466);
or UO_3483 (O_3483,N_29034,N_29327);
nor UO_3484 (O_3484,N_29830,N_29448);
xor UO_3485 (O_3485,N_29050,N_29094);
or UO_3486 (O_3486,N_29742,N_29768);
nor UO_3487 (O_3487,N_28706,N_28606);
nand UO_3488 (O_3488,N_29039,N_29427);
and UO_3489 (O_3489,N_28941,N_29012);
nand UO_3490 (O_3490,N_29740,N_28602);
nor UO_3491 (O_3491,N_28814,N_29016);
nor UO_3492 (O_3492,N_29906,N_29398);
nor UO_3493 (O_3493,N_28524,N_28620);
or UO_3494 (O_3494,N_29930,N_29717);
and UO_3495 (O_3495,N_29362,N_28945);
and UO_3496 (O_3496,N_29677,N_29326);
xnor UO_3497 (O_3497,N_28638,N_29195);
nand UO_3498 (O_3498,N_29938,N_28704);
or UO_3499 (O_3499,N_29594,N_29223);
endmodule