module basic_1000_10000_1500_2_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5005,N_5007,N_5008,N_5011,N_5014,N_5017,N_5019,N_5020,N_5021,N_5022,N_5024,N_5025,N_5026,N_5030,N_5032,N_5034,N_5036,N_5038,N_5041,N_5042,N_5044,N_5047,N_5048,N_5050,N_5056,N_5057,N_5058,N_5060,N_5063,N_5064,N_5065,N_5067,N_5068,N_5069,N_5073,N_5074,N_5076,N_5078,N_5081,N_5082,N_5083,N_5085,N_5087,N_5088,N_5094,N_5096,N_5097,N_5098,N_5099,N_5102,N_5104,N_5109,N_5111,N_5114,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5123,N_5124,N_5125,N_5128,N_5129,N_5135,N_5136,N_5137,N_5139,N_5140,N_5142,N_5145,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5154,N_5155,N_5156,N_5157,N_5158,N_5160,N_5161,N_5162,N_5163,N_5165,N_5166,N_5167,N_5168,N_5169,N_5171,N_5172,N_5174,N_5175,N_5176,N_5177,N_5178,N_5180,N_5182,N_5183,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5193,N_5194,N_5196,N_5197,N_5199,N_5200,N_5201,N_5202,N_5203,N_5205,N_5206,N_5207,N_5210,N_5211,N_5212,N_5213,N_5215,N_5216,N_5218,N_5220,N_5221,N_5223,N_5224,N_5225,N_5227,N_5229,N_5231,N_5234,N_5235,N_5236,N_5239,N_5241,N_5242,N_5243,N_5246,N_5248,N_5249,N_5252,N_5253,N_5255,N_5258,N_5259,N_5261,N_5262,N_5263,N_5265,N_5266,N_5267,N_5269,N_5272,N_5273,N_5274,N_5275,N_5278,N_5282,N_5283,N_5284,N_5285,N_5286,N_5288,N_5289,N_5290,N_5292,N_5293,N_5294,N_5295,N_5296,N_5299,N_5300,N_5302,N_5303,N_5304,N_5305,N_5307,N_5309,N_5310,N_5311,N_5312,N_5314,N_5315,N_5325,N_5326,N_5327,N_5329,N_5331,N_5332,N_5334,N_5335,N_5336,N_5339,N_5340,N_5343,N_5344,N_5345,N_5348,N_5350,N_5352,N_5353,N_5354,N_5357,N_5358,N_5359,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5370,N_5372,N_5373,N_5374,N_5376,N_5377,N_5380,N_5382,N_5383,N_5384,N_5385,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5398,N_5399,N_5400,N_5402,N_5403,N_5404,N_5406,N_5407,N_5410,N_5411,N_5412,N_5413,N_5416,N_5417,N_5418,N_5419,N_5420,N_5423,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5438,N_5439,N_5440,N_5441,N_5443,N_5445,N_5447,N_5448,N_5449,N_5450,N_5451,N_5454,N_5455,N_5458,N_5460,N_5461,N_5465,N_5466,N_5467,N_5468,N_5470,N_5475,N_5476,N_5478,N_5479,N_5480,N_5481,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5493,N_5494,N_5498,N_5499,N_5500,N_5501,N_5504,N_5506,N_5507,N_5509,N_5510,N_5511,N_5513,N_5514,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5526,N_5527,N_5528,N_5530,N_5532,N_5533,N_5536,N_5537,N_5540,N_5542,N_5543,N_5544,N_5545,N_5546,N_5548,N_5551,N_5552,N_5553,N_5554,N_5555,N_5557,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5568,N_5569,N_5570,N_5571,N_5573,N_5574,N_5577,N_5578,N_5581,N_5582,N_5583,N_5584,N_5585,N_5588,N_5589,N_5591,N_5594,N_5595,N_5596,N_5597,N_5601,N_5604,N_5605,N_5611,N_5612,N_5617,N_5618,N_5620,N_5622,N_5623,N_5624,N_5625,N_5629,N_5630,N_5631,N_5633,N_5634,N_5636,N_5637,N_5638,N_5643,N_5645,N_5647,N_5648,N_5649,N_5651,N_5653,N_5656,N_5659,N_5660,N_5661,N_5664,N_5665,N_5668,N_5669,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5679,N_5680,N_5684,N_5687,N_5688,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5700,N_5701,N_5702,N_5705,N_5706,N_5710,N_5711,N_5714,N_5718,N_5719,N_5721,N_5724,N_5727,N_5728,N_5729,N_5730,N_5734,N_5735,N_5736,N_5737,N_5741,N_5743,N_5744,N_5746,N_5748,N_5749,N_5751,N_5752,N_5755,N_5756,N_5757,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5769,N_5770,N_5772,N_5773,N_5774,N_5775,N_5776,N_5779,N_5781,N_5783,N_5785,N_5786,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5800,N_5802,N_5803,N_5811,N_5812,N_5815,N_5817,N_5818,N_5819,N_5820,N_5823,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5834,N_5836,N_5840,N_5841,N_5842,N_5844,N_5845,N_5848,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5860,N_5862,N_5864,N_5865,N_5869,N_5870,N_5871,N_5873,N_5874,N_5876,N_5877,N_5879,N_5881,N_5882,N_5883,N_5884,N_5888,N_5889,N_5890,N_5891,N_5894,N_5895,N_5899,N_5901,N_5903,N_5904,N_5905,N_5906,N_5908,N_5909,N_5910,N_5914,N_5915,N_5917,N_5918,N_5920,N_5924,N_5926,N_5927,N_5928,N_5930,N_5931,N_5932,N_5934,N_5935,N_5936,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5950,N_5951,N_5953,N_5956,N_5960,N_5962,N_5963,N_5964,N_5965,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5976,N_5978,N_5981,N_5982,N_5983,N_5984,N_5988,N_5990,N_5992,N_5994,N_5995,N_5996,N_5998,N_6001,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6011,N_6012,N_6014,N_6016,N_6017,N_6019,N_6024,N_6025,N_6027,N_6029,N_6030,N_6032,N_6034,N_6036,N_6037,N_6039,N_6040,N_6042,N_6044,N_6045,N_6049,N_6050,N_6051,N_6052,N_6054,N_6057,N_6058,N_6060,N_6062,N_6065,N_6066,N_6067,N_6070,N_6071,N_6074,N_6076,N_6077,N_6079,N_6082,N_6083,N_6087,N_6088,N_6089,N_6092,N_6093,N_6094,N_6099,N_6101,N_6102,N_6103,N_6104,N_6106,N_6107,N_6108,N_6109,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6119,N_6120,N_6121,N_6122,N_6124,N_6125,N_6128,N_6130,N_6132,N_6135,N_6139,N_6140,N_6142,N_6143,N_6144,N_6145,N_6150,N_6151,N_6152,N_6154,N_6155,N_6156,N_6157,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6171,N_6172,N_6179,N_6182,N_6183,N_6184,N_6185,N_6187,N_6189,N_6194,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6205,N_6206,N_6209,N_6210,N_6211,N_6212,N_6216,N_6218,N_6220,N_6224,N_6225,N_6226,N_6227,N_6229,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6241,N_6242,N_6243,N_6244,N_6245,N_6248,N_6250,N_6251,N_6252,N_6253,N_6255,N_6256,N_6257,N_6259,N_6260,N_6261,N_6262,N_6264,N_6269,N_6270,N_6271,N_6272,N_6274,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6296,N_6297,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6317,N_6318,N_6319,N_6320,N_6322,N_6323,N_6325,N_6326,N_6330,N_6331,N_6332,N_6333,N_6335,N_6337,N_6341,N_6343,N_6344,N_6348,N_6349,N_6350,N_6351,N_6354,N_6357,N_6362,N_6364,N_6367,N_6369,N_6371,N_6372,N_6375,N_6376,N_6379,N_6380,N_6382,N_6385,N_6386,N_6390,N_6391,N_6392,N_6395,N_6396,N_6400,N_6401,N_6402,N_6403,N_6405,N_6406,N_6407,N_6409,N_6410,N_6411,N_6414,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6427,N_6429,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6447,N_6448,N_6449,N_6451,N_6456,N_6459,N_6461,N_6462,N_6465,N_6466,N_6467,N_6468,N_6470,N_6471,N_6473,N_6474,N_6475,N_6476,N_6477,N_6480,N_6482,N_6484,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6497,N_6501,N_6502,N_6503,N_6504,N_6507,N_6509,N_6511,N_6512,N_6513,N_6516,N_6517,N_6519,N_6520,N_6523,N_6524,N_6526,N_6527,N_6528,N_6530,N_6531,N_6532,N_6533,N_6534,N_6536,N_6537,N_6538,N_6542,N_6543,N_6546,N_6549,N_6550,N_6551,N_6555,N_6556,N_6560,N_6561,N_6563,N_6565,N_6569,N_6570,N_6571,N_6572,N_6573,N_6575,N_6577,N_6578,N_6579,N_6582,N_6584,N_6586,N_6587,N_6589,N_6592,N_6594,N_6597,N_6598,N_6599,N_6601,N_6605,N_6606,N_6607,N_6608,N_6610,N_6613,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6626,N_6627,N_6629,N_6632,N_6633,N_6634,N_6636,N_6637,N_6640,N_6641,N_6642,N_6644,N_6645,N_6647,N_6650,N_6651,N_6652,N_6654,N_6655,N_6656,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6665,N_6666,N_6667,N_6669,N_6670,N_6673,N_6675,N_6676,N_6677,N_6678,N_6679,N_6681,N_6682,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6693,N_6694,N_6695,N_6696,N_6697,N_6699,N_6702,N_6703,N_6704,N_6707,N_6708,N_6710,N_6711,N_6714,N_6716,N_6717,N_6724,N_6729,N_6730,N_6731,N_6732,N_6733,N_6739,N_6740,N_6741,N_6742,N_6744,N_6745,N_6746,N_6748,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6759,N_6767,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6778,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6790,N_6793,N_6794,N_6797,N_6798,N_6799,N_6801,N_6802,N_6805,N_6807,N_6808,N_6811,N_6814,N_6817,N_6818,N_6820,N_6824,N_6826,N_6827,N_6829,N_6834,N_6835,N_6836,N_6839,N_6841,N_6844,N_6846,N_6847,N_6848,N_6849,N_6850,N_6853,N_6854,N_6855,N_6856,N_6858,N_6859,N_6860,N_6863,N_6867,N_6868,N_6869,N_6871,N_6873,N_6875,N_6878,N_6880,N_6881,N_6882,N_6884,N_6886,N_6887,N_6888,N_6889,N_6890,N_6892,N_6893,N_6895,N_6896,N_6897,N_6899,N_6901,N_6904,N_6906,N_6908,N_6911,N_6915,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6926,N_6927,N_6928,N_6929,N_6931,N_6932,N_6933,N_6934,N_6936,N_6937,N_6938,N_6939,N_6943,N_6944,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6957,N_6959,N_6960,N_6963,N_6966,N_6967,N_6968,N_6970,N_6973,N_6974,N_6979,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6988,N_6991,N_6993,N_6994,N_6995,N_6997,N_6999,N_7000,N_7001,N_7003,N_7004,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7016,N_7017,N_7019,N_7022,N_7024,N_7025,N_7026,N_7028,N_7030,N_7031,N_7032,N_7034,N_7037,N_7038,N_7040,N_7041,N_7042,N_7043,N_7045,N_7046,N_7047,N_7048,N_7049,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7058,N_7059,N_7060,N_7061,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7070,N_7071,N_7073,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7084,N_7086,N_7088,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7105,N_7106,N_7107,N_7110,N_7114,N_7115,N_7117,N_7119,N_7120,N_7121,N_7123,N_7124,N_7125,N_7127,N_7128,N_7129,N_7130,N_7131,N_7133,N_7137,N_7139,N_7140,N_7141,N_7142,N_7143,N_7145,N_7146,N_7148,N_7152,N_7154,N_7155,N_7156,N_7157,N_7160,N_7162,N_7163,N_7164,N_7165,N_7171,N_7173,N_7174,N_7175,N_7176,N_7177,N_7183,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7196,N_7197,N_7198,N_7201,N_7203,N_7204,N_7206,N_7207,N_7208,N_7209,N_7210,N_7212,N_7213,N_7214,N_7217,N_7218,N_7220,N_7221,N_7222,N_7223,N_7225,N_7227,N_7228,N_7229,N_7230,N_7233,N_7235,N_7236,N_7237,N_7239,N_7242,N_7243,N_7245,N_7248,N_7250,N_7251,N_7253,N_7254,N_7255,N_7256,N_7258,N_7259,N_7260,N_7261,N_7262,N_7264,N_7265,N_7268,N_7269,N_7270,N_7271,N_7272,N_7274,N_7276,N_7277,N_7279,N_7280,N_7282,N_7283,N_7284,N_7285,N_7286,N_7289,N_7290,N_7293,N_7294,N_7295,N_7296,N_7298,N_7300,N_7303,N_7304,N_7305,N_7307,N_7308,N_7309,N_7310,N_7311,N_7313,N_7315,N_7316,N_7318,N_7319,N_7322,N_7324,N_7326,N_7327,N_7328,N_7329,N_7330,N_7334,N_7335,N_7336,N_7337,N_7338,N_7341,N_7343,N_7344,N_7345,N_7346,N_7348,N_7349,N_7351,N_7352,N_7354,N_7356,N_7357,N_7363,N_7365,N_7366,N_7367,N_7368,N_7373,N_7375,N_7376,N_7378,N_7379,N_7381,N_7382,N_7383,N_7385,N_7386,N_7387,N_7388,N_7389,N_7393,N_7394,N_7397,N_7399,N_7402,N_7403,N_7404,N_7408,N_7409,N_7412,N_7414,N_7419,N_7421,N_7425,N_7426,N_7427,N_7429,N_7434,N_7436,N_7438,N_7439,N_7443,N_7444,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7455,N_7456,N_7461,N_7462,N_7463,N_7465,N_7466,N_7467,N_7469,N_7470,N_7471,N_7472,N_7473,N_7475,N_7476,N_7479,N_7480,N_7483,N_7484,N_7485,N_7486,N_7487,N_7489,N_7492,N_7493,N_7496,N_7498,N_7499,N_7500,N_7502,N_7503,N_7504,N_7507,N_7508,N_7510,N_7513,N_7514,N_7516,N_7517,N_7520,N_7521,N_7522,N_7523,N_7526,N_7527,N_7529,N_7531,N_7533,N_7534,N_7536,N_7537,N_7538,N_7540,N_7542,N_7544,N_7545,N_7546,N_7547,N_7548,N_7553,N_7554,N_7556,N_7558,N_7559,N_7567,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7580,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7590,N_7592,N_7593,N_7594,N_7595,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7605,N_7607,N_7608,N_7609,N_7610,N_7614,N_7615,N_7618,N_7620,N_7623,N_7624,N_7627,N_7629,N_7630,N_7632,N_7634,N_7635,N_7636,N_7638,N_7641,N_7642,N_7643,N_7645,N_7646,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7660,N_7661,N_7666,N_7668,N_7669,N_7670,N_7671,N_7672,N_7675,N_7676,N_7677,N_7678,N_7679,N_7681,N_7682,N_7683,N_7684,N_7687,N_7689,N_7699,N_7700,N_7701,N_7704,N_7705,N_7706,N_7709,N_7710,N_7712,N_7713,N_7715,N_7716,N_7717,N_7718,N_7719,N_7722,N_7723,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7734,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7745,N_7748,N_7751,N_7752,N_7754,N_7755,N_7756,N_7759,N_7760,N_7761,N_7762,N_7764,N_7765,N_7768,N_7771,N_7773,N_7775,N_7777,N_7778,N_7781,N_7783,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7795,N_7796,N_7798,N_7799,N_7801,N_7803,N_7806,N_7809,N_7811,N_7815,N_7817,N_7818,N_7819,N_7820,N_7821,N_7823,N_7824,N_7826,N_7827,N_7828,N_7831,N_7832,N_7834,N_7835,N_7837,N_7838,N_7840,N_7841,N_7844,N_7846,N_7847,N_7849,N_7852,N_7853,N_7854,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7872,N_7873,N_7876,N_7877,N_7878,N_7879,N_7880,N_7883,N_7885,N_7887,N_7889,N_7891,N_7893,N_7894,N_7895,N_7896,N_7898,N_7899,N_7900,N_7901,N_7902,N_7904,N_7910,N_7911,N_7912,N_7913,N_7914,N_7916,N_7917,N_7923,N_7925,N_7926,N_7929,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7940,N_7944,N_7945,N_7947,N_7949,N_7951,N_7955,N_7956,N_7957,N_7958,N_7960,N_7961,N_7964,N_7965,N_7966,N_7968,N_7972,N_7974,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7986,N_7987,N_7995,N_7999,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8010,N_8011,N_8012,N_8015,N_8016,N_8020,N_8025,N_8026,N_8027,N_8028,N_8029,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8042,N_8045,N_8047,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8061,N_8064,N_8065,N_8067,N_8068,N_8069,N_8070,N_8073,N_8074,N_8075,N_8077,N_8078,N_8080,N_8081,N_8082,N_8083,N_8085,N_8086,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8099,N_8101,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8112,N_8113,N_8114,N_8119,N_8120,N_8125,N_8128,N_8129,N_8130,N_8133,N_8136,N_8137,N_8138,N_8141,N_8144,N_8145,N_8147,N_8148,N_8150,N_8151,N_8152,N_8154,N_8156,N_8157,N_8158,N_8161,N_8162,N_8163,N_8164,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8176,N_8177,N_8179,N_8180,N_8182,N_8183,N_8184,N_8185,N_8186,N_8189,N_8190,N_8192,N_8194,N_8196,N_8197,N_8200,N_8202,N_8204,N_8205,N_8206,N_8208,N_8209,N_8211,N_8213,N_8214,N_8221,N_8222,N_8225,N_8226,N_8227,N_8229,N_8233,N_8234,N_8235,N_8236,N_8239,N_8240,N_8241,N_8242,N_8244,N_8250,N_8251,N_8253,N_8255,N_8256,N_8257,N_8258,N_8260,N_8262,N_8265,N_8268,N_8270,N_8272,N_8273,N_8277,N_8278,N_8279,N_8280,N_8281,N_8283,N_8284,N_8285,N_8286,N_8287,N_8290,N_8291,N_8293,N_8294,N_8296,N_8297,N_8299,N_8301,N_8303,N_8304,N_8305,N_8306,N_8308,N_8309,N_8310,N_8311,N_8312,N_8314,N_8318,N_8320,N_8321,N_8323,N_8325,N_8327,N_8328,N_8329,N_8330,N_8332,N_8333,N_8335,N_8337,N_8340,N_8341,N_8342,N_8343,N_8344,N_8348,N_8349,N_8350,N_8351,N_8352,N_8354,N_8355,N_8357,N_8358,N_8361,N_8362,N_8363,N_8366,N_8367,N_8371,N_8372,N_8373,N_8374,N_8377,N_8378,N_8379,N_8382,N_8384,N_8386,N_8387,N_8390,N_8392,N_8393,N_8394,N_8395,N_8397,N_8399,N_8401,N_8402,N_8404,N_8405,N_8407,N_8410,N_8412,N_8413,N_8414,N_8416,N_8417,N_8419,N_8424,N_8425,N_8428,N_8430,N_8431,N_8433,N_8434,N_8436,N_8437,N_8438,N_8439,N_8440,N_8442,N_8445,N_8447,N_8448,N_8449,N_8450,N_8452,N_8454,N_8457,N_8460,N_8463,N_8464,N_8465,N_8468,N_8469,N_8471,N_8472,N_8474,N_8478,N_8480,N_8481,N_8482,N_8483,N_8487,N_8488,N_8489,N_8491,N_8493,N_8494,N_8495,N_8496,N_8498,N_8499,N_8500,N_8501,N_8504,N_8506,N_8507,N_8508,N_8510,N_8513,N_8514,N_8515,N_8516,N_8519,N_8520,N_8521,N_8522,N_8523,N_8529,N_8531,N_8533,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8546,N_8548,N_8549,N_8552,N_8554,N_8558,N_8563,N_8564,N_8566,N_8571,N_8573,N_8574,N_8575,N_8578,N_8579,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8589,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8605,N_8606,N_8609,N_8615,N_8616,N_8618,N_8620,N_8621,N_8623,N_8624,N_8625,N_8626,N_8629,N_8630,N_8632,N_8633,N_8635,N_8636,N_8640,N_8642,N_8643,N_8644,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8655,N_8656,N_8659,N_8660,N_8661,N_8663,N_8664,N_8665,N_8667,N_8668,N_8669,N_8671,N_8674,N_8676,N_8681,N_8683,N_8685,N_8686,N_8689,N_8690,N_8692,N_8694,N_8696,N_8698,N_8699,N_8700,N_8702,N_8703,N_8704,N_8705,N_8706,N_8709,N_8710,N_8712,N_8716,N_8717,N_8718,N_8720,N_8721,N_8722,N_8729,N_8730,N_8731,N_8732,N_8733,N_8735,N_8736,N_8739,N_8741,N_8742,N_8743,N_8745,N_8746,N_8747,N_8749,N_8751,N_8752,N_8755,N_8756,N_8758,N_8760,N_8762,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8773,N_8774,N_8775,N_8776,N_8779,N_8780,N_8781,N_8782,N_8784,N_8786,N_8787,N_8788,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8797,N_8798,N_8800,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8816,N_8817,N_8819,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8832,N_8834,N_8836,N_8838,N_8840,N_8841,N_8842,N_8843,N_8844,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8855,N_8856,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8865,N_8867,N_8868,N_8869,N_8870,N_8873,N_8874,N_8875,N_8876,N_8878,N_8883,N_8886,N_8888,N_8890,N_8891,N_8892,N_8893,N_8895,N_8898,N_8899,N_8900,N_8901,N_8905,N_8907,N_8908,N_8909,N_8912,N_8915,N_8916,N_8917,N_8920,N_8921,N_8922,N_8924,N_8925,N_8926,N_8928,N_8929,N_8931,N_8933,N_8935,N_8936,N_8937,N_8942,N_8943,N_8944,N_8947,N_8948,N_8952,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8965,N_8968,N_8972,N_8973,N_8976,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8986,N_8987,N_8989,N_8993,N_8996,N_8997,N_8999,N_9001,N_9002,N_9003,N_9004,N_9005,N_9008,N_9010,N_9012,N_9014,N_9016,N_9017,N_9019,N_9021,N_9022,N_9023,N_9028,N_9029,N_9030,N_9031,N_9036,N_9037,N_9038,N_9039,N_9040,N_9042,N_9043,N_9044,N_9046,N_9047,N_9048,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9062,N_9063,N_9066,N_9067,N_9069,N_9070,N_9072,N_9074,N_9075,N_9076,N_9077,N_9079,N_9080,N_9081,N_9083,N_9084,N_9085,N_9088,N_9089,N_9093,N_9095,N_9096,N_9098,N_9103,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9115,N_9116,N_9117,N_9118,N_9120,N_9121,N_9122,N_9123,N_9126,N_9129,N_9130,N_9131,N_9132,N_9133,N_9135,N_9137,N_9138,N_9140,N_9141,N_9143,N_9144,N_9147,N_9149,N_9150,N_9151,N_9152,N_9153,N_9156,N_9157,N_9160,N_9162,N_9163,N_9164,N_9165,N_9168,N_9169,N_9170,N_9173,N_9174,N_9175,N_9176,N_9180,N_9181,N_9182,N_9183,N_9186,N_9190,N_9191,N_9192,N_9193,N_9194,N_9196,N_9197,N_9199,N_9201,N_9202,N_9203,N_9204,N_9206,N_9208,N_9210,N_9211,N_9213,N_9215,N_9217,N_9222,N_9224,N_9225,N_9228,N_9229,N_9231,N_9232,N_9233,N_9234,N_9235,N_9237,N_9239,N_9240,N_9241,N_9243,N_9248,N_9250,N_9251,N_9252,N_9253,N_9254,N_9256,N_9258,N_9260,N_9261,N_9265,N_9266,N_9267,N_9269,N_9270,N_9273,N_9277,N_9279,N_9280,N_9282,N_9283,N_9284,N_9287,N_9288,N_9289,N_9290,N_9292,N_9293,N_9296,N_9297,N_9300,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9311,N_9313,N_9314,N_9315,N_9317,N_9318,N_9320,N_9321,N_9322,N_9326,N_9333,N_9335,N_9336,N_9338,N_9339,N_9340,N_9342,N_9343,N_9346,N_9348,N_9349,N_9350,N_9351,N_9354,N_9355,N_9356,N_9357,N_9361,N_9364,N_9365,N_9366,N_9369,N_9370,N_9373,N_9375,N_9379,N_9380,N_9383,N_9384,N_9385,N_9388,N_9389,N_9390,N_9393,N_9394,N_9396,N_9398,N_9400,N_9401,N_9402,N_9405,N_9406,N_9407,N_9408,N_9410,N_9411,N_9412,N_9414,N_9416,N_9418,N_9419,N_9420,N_9422,N_9425,N_9426,N_9427,N_9428,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9438,N_9439,N_9440,N_9441,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9451,N_9453,N_9455,N_9457,N_9458,N_9459,N_9460,N_9462,N_9463,N_9464,N_9465,N_9466,N_9468,N_9470,N_9471,N_9472,N_9473,N_9476,N_9477,N_9480,N_9481,N_9483,N_9484,N_9486,N_9487,N_9488,N_9489,N_9491,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9504,N_9505,N_9506,N_9508,N_9509,N_9510,N_9512,N_9514,N_9516,N_9521,N_9523,N_9524,N_9525,N_9526,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9537,N_9541,N_9547,N_9548,N_9551,N_9553,N_9554,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9566,N_9567,N_9571,N_9572,N_9575,N_9576,N_9577,N_9578,N_9580,N_9581,N_9582,N_9588,N_9589,N_9590,N_9592,N_9593,N_9595,N_9596,N_9597,N_9599,N_9600,N_9602,N_9604,N_9607,N_9609,N_9613,N_9614,N_9618,N_9619,N_9624,N_9625,N_9627,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9639,N_9647,N_9648,N_9654,N_9656,N_9659,N_9661,N_9665,N_9666,N_9667,N_9669,N_9670,N_9671,N_9673,N_9674,N_9676,N_9677,N_9679,N_9680,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9696,N_9697,N_9699,N_9700,N_9703,N_9704,N_9705,N_9706,N_9707,N_9709,N_9710,N_9713,N_9714,N_9715,N_9716,N_9717,N_9722,N_9723,N_9726,N_9728,N_9730,N_9731,N_9732,N_9734,N_9735,N_9736,N_9740,N_9742,N_9745,N_9747,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9757,N_9759,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9772,N_9774,N_9776,N_9777,N_9779,N_9781,N_9782,N_9783,N_9785,N_9787,N_9789,N_9791,N_9794,N_9795,N_9796,N_9797,N_9799,N_9800,N_9801,N_9802,N_9803,N_9810,N_9811,N_9814,N_9815,N_9816,N_9818,N_9819,N_9820,N_9821,N_9822,N_9825,N_9826,N_9827,N_9828,N_9832,N_9834,N_9835,N_9838,N_9839,N_9840,N_9841,N_9842,N_9844,N_9845,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9854,N_9855,N_9856,N_9858,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9872,N_9873,N_9875,N_9876,N_9877,N_9878,N_9882,N_9883,N_9885,N_9887,N_9888,N_9890,N_9891,N_9892,N_9894,N_9895,N_9896,N_9897,N_9899,N_9900,N_9902,N_9903,N_9907,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9916,N_9919,N_9920,N_9923,N_9924,N_9925,N_9926,N_9928,N_9930,N_9932,N_9935,N_9936,N_9937,N_9939,N_9943,N_9944,N_9947,N_9948,N_9950,N_9951,N_9955,N_9956,N_9958,N_9961,N_9965,N_9966,N_9967,N_9969,N_9970,N_9972,N_9973,N_9977,N_9979,N_9980,N_9982,N_9983,N_9985,N_9986,N_9988,N_9992,N_9995,N_9996,N_9997,N_9998;
nor U0 (N_0,In_27,In_511);
nor U1 (N_1,In_41,In_802);
and U2 (N_2,In_73,In_357);
nand U3 (N_3,In_633,In_827);
and U4 (N_4,In_236,In_735);
nor U5 (N_5,In_274,In_321);
nand U6 (N_6,In_222,In_749);
or U7 (N_7,In_255,In_868);
nor U8 (N_8,In_576,In_798);
or U9 (N_9,In_591,In_743);
nor U10 (N_10,In_266,In_111);
and U11 (N_11,In_97,In_597);
nor U12 (N_12,In_230,In_855);
and U13 (N_13,In_930,In_549);
or U14 (N_14,In_962,In_218);
nor U15 (N_15,In_937,In_895);
nor U16 (N_16,In_717,In_156);
nand U17 (N_17,In_692,In_562);
or U18 (N_18,In_420,In_63);
or U19 (N_19,In_838,In_852);
nand U20 (N_20,In_145,In_526);
nor U21 (N_21,In_303,In_793);
nand U22 (N_22,In_744,In_242);
nor U23 (N_23,In_513,In_983);
xor U24 (N_24,In_929,In_415);
and U25 (N_25,In_905,In_517);
xnor U26 (N_26,In_657,In_469);
xnor U27 (N_27,In_699,In_470);
nand U28 (N_28,In_371,In_521);
nor U29 (N_29,In_75,In_882);
or U30 (N_30,In_495,In_378);
nand U31 (N_31,In_965,In_38);
nor U32 (N_32,In_402,In_724);
nor U33 (N_33,In_853,In_836);
or U34 (N_34,In_959,In_751);
nand U35 (N_35,In_279,In_989);
nand U36 (N_36,In_306,In_92);
xnor U37 (N_37,In_880,In_122);
nand U38 (N_38,In_168,In_430);
xnor U39 (N_39,In_36,In_98);
nand U40 (N_40,In_834,In_795);
nand U41 (N_41,In_133,In_747);
nor U42 (N_42,In_803,In_756);
xnor U43 (N_43,In_332,In_897);
nand U44 (N_44,In_90,In_709);
nor U45 (N_45,In_314,In_736);
nand U46 (N_46,In_93,In_734);
or U47 (N_47,In_687,In_450);
xnor U48 (N_48,In_501,In_785);
nor U49 (N_49,In_351,In_523);
or U50 (N_50,In_954,In_758);
nand U51 (N_51,In_577,In_926);
nor U52 (N_52,In_537,In_137);
nor U53 (N_53,In_528,In_10);
nand U54 (N_54,In_573,In_176);
and U55 (N_55,In_559,In_851);
or U56 (N_56,In_14,In_428);
nor U57 (N_57,In_726,In_718);
nand U58 (N_58,In_896,In_197);
or U59 (N_59,In_37,In_149);
nor U60 (N_60,In_147,In_109);
and U61 (N_61,In_201,In_878);
nand U62 (N_62,In_45,In_932);
xor U63 (N_63,In_273,In_369);
nand U64 (N_64,In_150,In_323);
nor U65 (N_65,In_384,In_640);
nor U66 (N_66,In_732,In_984);
and U67 (N_67,In_207,In_655);
and U68 (N_68,In_94,In_365);
and U69 (N_69,In_313,In_460);
nor U70 (N_70,In_858,In_923);
xnor U71 (N_71,In_911,In_754);
nand U72 (N_72,In_432,In_808);
nor U73 (N_73,In_47,In_261);
and U74 (N_74,In_26,In_307);
nor U75 (N_75,In_441,In_114);
and U76 (N_76,In_167,In_978);
xnor U77 (N_77,In_794,In_17);
nor U78 (N_78,In_603,In_714);
nor U79 (N_79,In_115,In_373);
nand U80 (N_80,In_716,In_945);
and U81 (N_81,In_776,In_381);
nor U82 (N_82,In_507,In_278);
nor U83 (N_83,In_52,In_967);
or U84 (N_84,In_998,In_957);
and U85 (N_85,In_169,In_894);
nor U86 (N_86,In_904,In_682);
nor U87 (N_87,In_525,In_812);
nand U88 (N_88,In_686,In_341);
nor U89 (N_89,In_500,In_696);
xor U90 (N_90,In_128,In_366);
or U91 (N_91,In_542,In_473);
nand U92 (N_92,In_489,In_879);
and U93 (N_93,In_418,In_229);
xor U94 (N_94,In_966,In_175);
and U95 (N_95,In_558,In_841);
or U96 (N_96,In_877,In_264);
and U97 (N_97,In_445,In_520);
and U98 (N_98,In_710,In_43);
xor U99 (N_99,In_370,In_297);
and U100 (N_100,In_312,In_654);
or U101 (N_101,In_555,In_24);
and U102 (N_102,In_706,In_829);
and U103 (N_103,In_857,In_202);
nor U104 (N_104,In_474,In_865);
xnor U105 (N_105,In_504,In_497);
or U106 (N_106,In_281,In_826);
nor U107 (N_107,In_112,In_408);
or U108 (N_108,In_590,In_358);
and U109 (N_109,In_985,In_621);
nand U110 (N_110,In_641,In_755);
or U111 (N_111,In_892,In_225);
and U112 (N_112,In_740,In_660);
nand U113 (N_113,In_162,In_205);
and U114 (N_114,In_854,In_174);
nand U115 (N_115,In_126,In_848);
nor U116 (N_116,In_825,In_410);
or U117 (N_117,In_424,In_545);
and U118 (N_118,In_54,In_579);
and U119 (N_119,In_350,In_818);
or U120 (N_120,In_413,In_20);
nor U121 (N_121,In_431,In_448);
and U122 (N_122,In_887,In_153);
xnor U123 (N_123,In_624,In_427);
and U124 (N_124,In_232,In_565);
or U125 (N_125,In_703,In_614);
nor U126 (N_126,In_239,In_914);
nand U127 (N_127,In_846,In_256);
nor U128 (N_128,In_867,In_189);
or U129 (N_129,In_209,In_300);
and U130 (N_130,In_581,In_416);
and U131 (N_131,In_801,In_146);
nand U132 (N_132,In_933,In_570);
and U133 (N_133,In_605,In_425);
xnor U134 (N_134,In_360,In_49);
and U135 (N_135,In_695,In_942);
nor U136 (N_136,In_889,In_117);
nand U137 (N_137,In_646,In_386);
or U138 (N_138,In_301,In_494);
and U139 (N_139,In_505,In_935);
or U140 (N_140,In_287,In_672);
or U141 (N_141,In_739,In_362);
nor U142 (N_142,In_569,In_257);
and U143 (N_143,In_275,In_198);
and U144 (N_144,In_130,In_429);
or U145 (N_145,In_364,In_131);
nor U146 (N_146,In_652,In_951);
nand U147 (N_147,In_804,In_688);
or U148 (N_148,In_401,In_771);
and U149 (N_149,In_102,In_79);
nand U150 (N_150,In_250,In_631);
or U151 (N_151,In_380,In_252);
nand U152 (N_152,In_452,In_200);
or U153 (N_153,In_941,In_188);
and U154 (N_154,In_680,In_639);
xor U155 (N_155,In_553,In_969);
nor U156 (N_156,In_265,In_78);
nand U157 (N_157,In_866,In_757);
nand U158 (N_158,In_763,In_705);
xnor U159 (N_159,In_394,In_293);
and U160 (N_160,In_268,In_220);
nor U161 (N_161,In_439,In_689);
or U162 (N_162,In_21,In_347);
or U163 (N_163,In_320,In_151);
and U164 (N_164,In_18,In_407);
or U165 (N_165,In_701,In_863);
nor U166 (N_166,In_159,In_601);
or U167 (N_167,In_971,In_95);
or U168 (N_168,In_673,In_15);
or U169 (N_169,In_647,In_568);
nand U170 (N_170,In_271,In_847);
nor U171 (N_171,In_694,In_119);
nand U172 (N_172,In_913,In_800);
or U173 (N_173,In_23,In_616);
xnor U174 (N_174,In_330,In_698);
nand U175 (N_175,In_13,In_561);
nor U176 (N_176,In_368,In_564);
and U177 (N_177,In_819,In_515);
or U178 (N_178,In_843,In_25);
nand U179 (N_179,In_886,In_96);
nand U180 (N_180,In_272,In_766);
xnor U181 (N_181,In_912,In_86);
nand U182 (N_182,In_183,In_361);
xor U183 (N_183,In_231,In_872);
xnor U184 (N_184,In_178,In_669);
and U185 (N_185,In_512,In_228);
xor U186 (N_186,In_849,In_830);
nor U187 (N_187,In_638,In_240);
nand U188 (N_188,In_806,In_772);
and U189 (N_189,In_157,In_805);
or U190 (N_190,In_580,In_88);
or U191 (N_191,In_524,In_331);
nand U192 (N_192,In_529,In_124);
nor U193 (N_193,In_491,In_583);
or U194 (N_194,In_9,In_179);
nor U195 (N_195,In_234,In_817);
or U196 (N_196,In_540,In_65);
or U197 (N_197,In_376,In_53);
nor U198 (N_198,In_77,In_963);
xor U199 (N_199,In_636,In_502);
nand U200 (N_200,In_514,In_977);
nor U201 (N_201,In_527,In_767);
nor U202 (N_202,In_574,In_161);
nand U203 (N_203,In_733,In_700);
and U204 (N_204,In_936,In_404);
nand U205 (N_205,In_107,In_283);
nand U206 (N_206,In_51,In_80);
nand U207 (N_207,In_393,In_437);
nor U208 (N_208,In_304,In_685);
xor U209 (N_209,In_241,In_215);
xor U210 (N_210,In_436,In_343);
nand U211 (N_211,In_35,In_349);
and U212 (N_212,In_392,In_869);
xor U213 (N_213,In_728,In_282);
nand U214 (N_214,In_129,In_958);
nand U215 (N_215,In_449,In_876);
and U216 (N_216,In_650,In_5);
nor U217 (N_217,In_503,In_833);
xor U218 (N_218,In_158,In_831);
nor U219 (N_219,In_70,In_213);
nor U220 (N_220,In_651,In_196);
nor U221 (N_221,In_592,In_839);
or U222 (N_222,In_481,In_315);
and U223 (N_223,In_254,In_319);
nor U224 (N_224,In_480,In_888);
and U225 (N_225,In_644,In_656);
nand U226 (N_226,In_943,In_184);
or U227 (N_227,In_377,In_290);
or U228 (N_228,In_375,In_934);
or U229 (N_229,In_248,In_796);
or U230 (N_230,In_308,In_625);
nor U231 (N_231,In_760,In_7);
and U232 (N_232,In_192,In_916);
or U233 (N_233,In_548,In_783);
nor U234 (N_234,In_551,In_970);
nor U235 (N_235,In_211,In_604);
or U236 (N_236,In_132,In_342);
nand U237 (N_237,In_820,In_269);
nand U238 (N_238,In_285,In_779);
or U239 (N_239,In_403,In_901);
xnor U240 (N_240,In_333,In_438);
nand U241 (N_241,In_258,In_510);
nor U242 (N_242,In_60,In_46);
or U243 (N_243,In_856,In_753);
and U244 (N_244,In_667,In_774);
nand U245 (N_245,In_991,In_676);
or U246 (N_246,In_83,In_31);
nor U247 (N_247,In_1,In_367);
xnor U248 (N_248,In_881,In_533);
xnor U249 (N_249,In_2,In_642);
nand U250 (N_250,In_39,In_571);
nor U251 (N_251,In_670,In_987);
or U252 (N_252,In_68,In_467);
nor U253 (N_253,In_340,In_875);
nand U254 (N_254,In_534,In_165);
nor U255 (N_255,In_572,In_873);
and U256 (N_256,In_16,In_884);
nand U257 (N_257,In_182,In_89);
nor U258 (N_258,In_627,In_535);
or U259 (N_259,In_722,In_203);
or U260 (N_260,In_50,In_485);
nand U261 (N_261,In_786,In_994);
nor U262 (N_262,In_457,In_288);
or U263 (N_263,In_900,In_447);
nand U264 (N_264,In_547,In_472);
nor U265 (N_265,In_405,In_488);
or U266 (N_266,In_738,In_406);
xnor U267 (N_267,In_906,In_620);
and U268 (N_268,In_552,In_66);
and U269 (N_269,In_337,In_484);
xnor U270 (N_270,In_219,In_768);
xor U271 (N_271,In_379,In_423);
nand U272 (N_272,In_299,In_560);
nor U273 (N_273,In_166,In_944);
nor U274 (N_274,In_103,In_186);
and U275 (N_275,In_414,In_871);
or U276 (N_276,In_594,In_563);
nand U277 (N_277,In_606,In_910);
nor U278 (N_278,In_458,In_554);
nor U279 (N_279,In_118,In_440);
nor U280 (N_280,In_821,In_359);
or U281 (N_281,In_339,In_216);
nand U282 (N_282,In_777,In_33);
nor U283 (N_283,In_395,In_899);
nand U284 (N_284,In_148,In_160);
and U285 (N_285,In_530,In_61);
or U286 (N_286,In_451,In_674);
or U287 (N_287,In_702,In_536);
nor U288 (N_288,In_354,In_653);
nor U289 (N_289,In_531,In_298);
and U290 (N_290,In_71,In_861);
xnor U291 (N_291,In_557,In_649);
or U292 (N_292,In_6,In_435);
nand U293 (N_293,In_433,In_626);
or U294 (N_294,In_277,In_355);
and U295 (N_295,In_729,In_630);
and U296 (N_296,In_336,In_519);
or U297 (N_297,In_538,In_55);
nand U298 (N_298,In_120,In_338);
or U299 (N_299,In_398,In_328);
nor U300 (N_300,In_302,In_221);
nand U301 (N_301,In_832,In_939);
xor U302 (N_302,In_999,In_543);
nor U303 (N_303,In_334,In_976);
nor U304 (N_304,In_74,In_286);
and U305 (N_305,In_422,In_681);
nand U306 (N_306,In_745,In_32);
xor U307 (N_307,In_292,In_920);
nand U308 (N_308,In_479,In_842);
nor U309 (N_309,In_390,In_609);
and U310 (N_310,In_742,In_922);
nor U311 (N_311,In_588,In_723);
nand U312 (N_312,In_721,In_247);
nor U313 (N_313,In_975,In_586);
xnor U314 (N_314,In_475,In_125);
nor U315 (N_315,In_267,In_731);
xnor U316 (N_316,In_155,In_532);
nor U317 (N_317,In_823,In_665);
xnor U318 (N_318,In_797,In_82);
and U319 (N_319,In_72,In_87);
nor U320 (N_320,In_850,In_693);
nand U321 (N_321,In_311,In_172);
or U322 (N_322,In_421,In_938);
or U323 (N_323,In_496,In_417);
nor U324 (N_324,In_249,In_666);
or U325 (N_325,In_411,In_506);
or U326 (N_326,In_909,In_59);
nand U327 (N_327,In_675,In_11);
or U328 (N_328,In_964,In_468);
and U329 (N_329,In_979,In_101);
nor U330 (N_330,In_612,In_990);
nand U331 (N_331,In_578,In_305);
or U332 (N_332,In_140,In_643);
and U333 (N_333,In_903,In_318);
or U334 (N_334,In_289,In_845);
and U335 (N_335,In_623,In_874);
nand U336 (N_336,In_116,In_3);
and U337 (N_337,In_245,In_815);
nand U338 (N_338,In_566,In_34);
or U339 (N_339,In_142,In_187);
nand U340 (N_340,In_397,In_69);
nor U341 (N_341,In_446,In_509);
nor U342 (N_342,In_382,In_890);
nor U343 (N_343,In_762,In_353);
nor U344 (N_344,In_595,In_141);
nand U345 (N_345,In_658,In_988);
nor U346 (N_346,In_372,In_466);
nand U347 (N_347,In_622,In_345);
nand U348 (N_348,In_860,In_787);
and U349 (N_349,In_199,In_584);
nor U350 (N_350,In_915,In_809);
nand U351 (N_351,In_194,In_493);
nor U352 (N_352,In_346,In_712);
nand U353 (N_353,In_750,In_711);
nor U354 (N_354,In_589,In_948);
and U355 (N_355,In_765,In_206);
nor U356 (N_356,In_918,In_253);
nor U357 (N_357,In_629,In_280);
nor U358 (N_358,In_859,In_173);
and U359 (N_359,In_487,In_177);
and U360 (N_360,In_541,In_727);
and U361 (N_361,In_181,In_329);
nor U362 (N_362,In_764,In_344);
and U363 (N_363,In_953,In_251);
or U364 (N_364,In_262,In_136);
or U365 (N_365,In_81,In_637);
xnor U366 (N_366,In_471,In_409);
and U367 (N_367,In_664,In_388);
or U368 (N_368,In_104,In_227);
or U369 (N_369,In_807,In_518);
nor U370 (N_370,In_224,In_719);
or U371 (N_371,In_974,In_400);
nor U372 (N_372,In_310,In_661);
and U373 (N_373,In_814,In_662);
or U374 (N_374,In_972,In_443);
and U375 (N_375,In_697,In_968);
xnor U376 (N_376,In_725,In_645);
and U377 (N_377,In_214,In_84);
xnor U378 (N_378,In_171,In_309);
and U379 (N_379,In_840,In_508);
or U380 (N_380,In_243,In_907);
nor U381 (N_381,In_789,In_30);
or U382 (N_382,In_356,In_781);
nand U383 (N_383,In_946,In_29);
and U384 (N_384,In_608,In_459);
nor U385 (N_385,In_387,In_539);
nand U386 (N_386,In_134,In_486);
xnor U387 (N_387,In_947,In_891);
xnor U388 (N_388,In_477,In_600);
or U389 (N_389,In_374,In_138);
nor U390 (N_390,In_782,In_960);
or U391 (N_391,In_127,In_811);
nand U392 (N_392,In_788,In_973);
or U393 (N_393,In_810,In_263);
nor U394 (N_394,In_123,In_648);
and U395 (N_395,In_108,In_139);
xnor U396 (N_396,In_226,In_322);
nor U397 (N_397,In_522,In_544);
xnor U398 (N_398,In_659,In_799);
or U399 (N_399,In_291,In_483);
or U400 (N_400,In_883,In_615);
and U401 (N_401,In_844,In_931);
or U402 (N_402,In_980,In_316);
and U403 (N_403,In_56,In_956);
nand U404 (N_404,In_135,In_663);
nand U405 (N_405,In_121,In_412);
nor U406 (N_406,In_992,In_193);
nand U407 (N_407,In_259,In_57);
nand U408 (N_408,In_816,In_498);
nor U409 (N_409,In_940,In_363);
and U410 (N_410,In_22,In_492);
or U411 (N_411,In_949,In_164);
nand U412 (N_412,In_67,In_113);
or U413 (N_413,In_0,In_317);
or U414 (N_414,In_296,In_191);
xor U415 (N_415,In_180,In_596);
or U416 (N_416,In_775,In_585);
nor U417 (N_417,In_628,In_769);
and U418 (N_418,In_204,In_837);
or U419 (N_419,In_454,In_708);
or U420 (N_420,In_598,In_704);
nor U421 (N_421,In_163,In_737);
or U422 (N_422,In_324,In_870);
nand U423 (N_423,In_635,In_678);
nand U424 (N_424,In_143,In_599);
xor U425 (N_425,In_668,In_952);
nor U426 (N_426,In_476,In_752);
nand U427 (N_427,In_270,In_748);
and U428 (N_428,In_679,In_335);
nor U429 (N_429,In_835,In_58);
nor U430 (N_430,In_691,In_284);
nand U431 (N_431,In_741,In_327);
or U432 (N_432,In_210,In_419);
or U433 (N_433,In_455,In_683);
xor U434 (N_434,In_465,In_556);
and U435 (N_435,In_617,In_997);
and U436 (N_436,In_391,In_217);
nand U437 (N_437,In_784,In_813);
and U438 (N_438,In_961,In_864);
nor U439 (N_439,In_383,In_919);
or U440 (N_440,In_294,In_246);
nand U441 (N_441,In_607,In_713);
nor U442 (N_442,In_478,In_238);
nand U443 (N_443,In_778,In_917);
or U444 (N_444,In_276,In_352);
and U445 (N_445,In_195,In_19);
nor U446 (N_446,In_62,In_48);
nor U447 (N_447,In_925,In_634);
nand U448 (N_448,In_100,In_619);
nand U449 (N_449,In_385,In_770);
or U450 (N_450,In_85,In_893);
nand U451 (N_451,In_456,In_223);
nor U452 (N_452,In_862,In_593);
nand U453 (N_453,In_464,In_490);
and U454 (N_454,In_677,In_921);
or U455 (N_455,In_233,In_761);
and U456 (N_456,In_602,In_212);
and U457 (N_457,In_389,In_42);
nand U458 (N_458,In_244,In_618);
or U459 (N_459,In_325,In_707);
and U460 (N_460,In_8,In_190);
nor U461 (N_461,In_791,In_924);
and U462 (N_462,In_986,In_235);
and U463 (N_463,In_690,In_462);
and U464 (N_464,In_898,In_295);
nand U465 (N_465,In_773,In_996);
nand U466 (N_466,In_611,In_824);
nand U467 (N_467,In_780,In_185);
or U468 (N_468,In_575,In_790);
nand U469 (N_469,In_950,In_567);
and U470 (N_470,In_482,In_28);
and U471 (N_471,In_715,In_444);
nor U472 (N_472,In_759,In_106);
nor U473 (N_473,In_152,In_671);
nor U474 (N_474,In_399,In_91);
or U475 (N_475,In_99,In_587);
and U476 (N_476,In_792,In_105);
nor U477 (N_477,In_908,In_64);
or U478 (N_478,In_396,In_546);
nor U479 (N_479,In_76,In_463);
and U480 (N_480,In_4,In_822);
xnor U481 (N_481,In_550,In_981);
or U482 (N_482,In_144,In_746);
nand U483 (N_483,In_434,In_516);
and U484 (N_484,In_499,In_955);
nand U485 (N_485,In_684,In_613);
nor U486 (N_486,In_828,In_170);
xnor U487 (N_487,In_995,In_348);
nand U488 (N_488,In_632,In_885);
nor U489 (N_489,In_154,In_40);
and U490 (N_490,In_927,In_44);
or U491 (N_491,In_582,In_12);
xor U492 (N_492,In_730,In_610);
xnor U493 (N_493,In_461,In_110);
nor U494 (N_494,In_260,In_902);
or U495 (N_495,In_237,In_442);
xnor U496 (N_496,In_453,In_928);
nand U497 (N_497,In_426,In_326);
and U498 (N_498,In_208,In_720);
nand U499 (N_499,In_993,In_982);
and U500 (N_500,In_19,In_80);
nor U501 (N_501,In_715,In_676);
nand U502 (N_502,In_762,In_411);
nand U503 (N_503,In_695,In_877);
nor U504 (N_504,In_938,In_413);
nand U505 (N_505,In_475,In_805);
and U506 (N_506,In_548,In_249);
and U507 (N_507,In_157,In_818);
and U508 (N_508,In_268,In_34);
nor U509 (N_509,In_328,In_613);
and U510 (N_510,In_51,In_553);
nand U511 (N_511,In_213,In_75);
nor U512 (N_512,In_822,In_927);
nor U513 (N_513,In_726,In_141);
nand U514 (N_514,In_792,In_395);
nor U515 (N_515,In_883,In_205);
nand U516 (N_516,In_578,In_294);
xor U517 (N_517,In_507,In_959);
xor U518 (N_518,In_927,In_184);
xnor U519 (N_519,In_474,In_564);
nand U520 (N_520,In_337,In_439);
and U521 (N_521,In_463,In_949);
or U522 (N_522,In_571,In_895);
or U523 (N_523,In_934,In_862);
or U524 (N_524,In_980,In_480);
and U525 (N_525,In_509,In_338);
xnor U526 (N_526,In_748,In_369);
nand U527 (N_527,In_364,In_773);
and U528 (N_528,In_184,In_68);
and U529 (N_529,In_539,In_413);
or U530 (N_530,In_37,In_64);
nand U531 (N_531,In_942,In_820);
or U532 (N_532,In_555,In_511);
nor U533 (N_533,In_168,In_217);
or U534 (N_534,In_798,In_536);
nor U535 (N_535,In_431,In_158);
nor U536 (N_536,In_365,In_870);
or U537 (N_537,In_923,In_365);
and U538 (N_538,In_669,In_239);
or U539 (N_539,In_786,In_296);
and U540 (N_540,In_857,In_311);
and U541 (N_541,In_305,In_611);
nor U542 (N_542,In_945,In_23);
or U543 (N_543,In_657,In_278);
or U544 (N_544,In_585,In_468);
nand U545 (N_545,In_14,In_433);
nand U546 (N_546,In_748,In_914);
xnor U547 (N_547,In_581,In_401);
nand U548 (N_548,In_404,In_711);
nor U549 (N_549,In_263,In_704);
nor U550 (N_550,In_305,In_252);
xor U551 (N_551,In_934,In_785);
nor U552 (N_552,In_717,In_909);
nand U553 (N_553,In_144,In_904);
xor U554 (N_554,In_398,In_221);
and U555 (N_555,In_987,In_807);
nand U556 (N_556,In_39,In_81);
or U557 (N_557,In_96,In_190);
xnor U558 (N_558,In_596,In_452);
nor U559 (N_559,In_372,In_632);
or U560 (N_560,In_8,In_992);
xnor U561 (N_561,In_163,In_510);
nand U562 (N_562,In_987,In_82);
or U563 (N_563,In_84,In_662);
and U564 (N_564,In_65,In_277);
and U565 (N_565,In_30,In_574);
nand U566 (N_566,In_31,In_436);
nand U567 (N_567,In_275,In_836);
xor U568 (N_568,In_957,In_122);
or U569 (N_569,In_797,In_753);
nand U570 (N_570,In_208,In_584);
and U571 (N_571,In_563,In_161);
nor U572 (N_572,In_362,In_186);
and U573 (N_573,In_947,In_982);
nor U574 (N_574,In_59,In_118);
or U575 (N_575,In_936,In_457);
or U576 (N_576,In_117,In_727);
and U577 (N_577,In_37,In_583);
and U578 (N_578,In_181,In_840);
and U579 (N_579,In_421,In_900);
or U580 (N_580,In_779,In_140);
nand U581 (N_581,In_116,In_263);
xor U582 (N_582,In_881,In_345);
nor U583 (N_583,In_799,In_200);
nor U584 (N_584,In_201,In_293);
nand U585 (N_585,In_762,In_332);
and U586 (N_586,In_848,In_411);
or U587 (N_587,In_804,In_733);
and U588 (N_588,In_243,In_263);
or U589 (N_589,In_272,In_572);
and U590 (N_590,In_316,In_658);
nor U591 (N_591,In_28,In_646);
or U592 (N_592,In_750,In_752);
nor U593 (N_593,In_981,In_359);
nand U594 (N_594,In_699,In_702);
and U595 (N_595,In_600,In_28);
nor U596 (N_596,In_7,In_298);
nor U597 (N_597,In_678,In_704);
or U598 (N_598,In_413,In_849);
and U599 (N_599,In_192,In_231);
or U600 (N_600,In_66,In_797);
and U601 (N_601,In_196,In_569);
or U602 (N_602,In_299,In_452);
or U603 (N_603,In_656,In_731);
and U604 (N_604,In_97,In_884);
or U605 (N_605,In_835,In_287);
or U606 (N_606,In_656,In_505);
nand U607 (N_607,In_83,In_30);
and U608 (N_608,In_321,In_997);
nand U609 (N_609,In_371,In_235);
and U610 (N_610,In_950,In_811);
or U611 (N_611,In_597,In_670);
and U612 (N_612,In_822,In_421);
nand U613 (N_613,In_494,In_6);
nor U614 (N_614,In_322,In_146);
nand U615 (N_615,In_604,In_623);
or U616 (N_616,In_93,In_794);
and U617 (N_617,In_561,In_597);
or U618 (N_618,In_916,In_142);
or U619 (N_619,In_798,In_591);
or U620 (N_620,In_860,In_459);
nand U621 (N_621,In_497,In_131);
and U622 (N_622,In_929,In_268);
and U623 (N_623,In_463,In_83);
and U624 (N_624,In_344,In_185);
or U625 (N_625,In_6,In_277);
or U626 (N_626,In_808,In_36);
or U627 (N_627,In_280,In_726);
nand U628 (N_628,In_1,In_254);
or U629 (N_629,In_629,In_661);
and U630 (N_630,In_460,In_146);
and U631 (N_631,In_963,In_858);
nand U632 (N_632,In_920,In_714);
or U633 (N_633,In_925,In_794);
nor U634 (N_634,In_523,In_516);
or U635 (N_635,In_495,In_965);
and U636 (N_636,In_53,In_313);
nor U637 (N_637,In_673,In_815);
xor U638 (N_638,In_13,In_77);
and U639 (N_639,In_583,In_656);
and U640 (N_640,In_489,In_94);
nor U641 (N_641,In_797,In_963);
nand U642 (N_642,In_436,In_965);
nand U643 (N_643,In_220,In_513);
nand U644 (N_644,In_634,In_216);
nor U645 (N_645,In_916,In_56);
or U646 (N_646,In_532,In_432);
nand U647 (N_647,In_103,In_867);
nor U648 (N_648,In_831,In_369);
and U649 (N_649,In_300,In_467);
xnor U650 (N_650,In_465,In_464);
or U651 (N_651,In_103,In_382);
nor U652 (N_652,In_507,In_478);
nand U653 (N_653,In_129,In_493);
nand U654 (N_654,In_424,In_558);
nand U655 (N_655,In_94,In_839);
nand U656 (N_656,In_773,In_50);
or U657 (N_657,In_159,In_709);
or U658 (N_658,In_182,In_351);
or U659 (N_659,In_986,In_459);
or U660 (N_660,In_900,In_101);
or U661 (N_661,In_501,In_399);
and U662 (N_662,In_750,In_959);
xnor U663 (N_663,In_790,In_894);
nor U664 (N_664,In_96,In_683);
and U665 (N_665,In_697,In_484);
nand U666 (N_666,In_877,In_854);
nand U667 (N_667,In_403,In_950);
xor U668 (N_668,In_864,In_639);
or U669 (N_669,In_931,In_286);
nor U670 (N_670,In_952,In_971);
nand U671 (N_671,In_869,In_344);
nor U672 (N_672,In_656,In_12);
and U673 (N_673,In_525,In_106);
nand U674 (N_674,In_606,In_153);
xnor U675 (N_675,In_843,In_489);
and U676 (N_676,In_174,In_146);
and U677 (N_677,In_14,In_688);
nand U678 (N_678,In_97,In_843);
or U679 (N_679,In_939,In_622);
xnor U680 (N_680,In_565,In_498);
nor U681 (N_681,In_370,In_221);
or U682 (N_682,In_648,In_404);
nor U683 (N_683,In_372,In_825);
and U684 (N_684,In_890,In_803);
or U685 (N_685,In_399,In_583);
xor U686 (N_686,In_552,In_192);
or U687 (N_687,In_614,In_510);
or U688 (N_688,In_555,In_331);
nor U689 (N_689,In_214,In_340);
nor U690 (N_690,In_200,In_252);
nor U691 (N_691,In_351,In_957);
and U692 (N_692,In_458,In_929);
or U693 (N_693,In_20,In_571);
or U694 (N_694,In_986,In_103);
nor U695 (N_695,In_73,In_453);
nand U696 (N_696,In_76,In_630);
nor U697 (N_697,In_970,In_174);
nor U698 (N_698,In_683,In_788);
nand U699 (N_699,In_141,In_84);
and U700 (N_700,In_135,In_436);
nor U701 (N_701,In_463,In_437);
or U702 (N_702,In_224,In_344);
xnor U703 (N_703,In_481,In_739);
and U704 (N_704,In_517,In_908);
or U705 (N_705,In_873,In_988);
or U706 (N_706,In_971,In_685);
nor U707 (N_707,In_781,In_842);
or U708 (N_708,In_354,In_681);
or U709 (N_709,In_831,In_345);
and U710 (N_710,In_655,In_953);
xor U711 (N_711,In_119,In_438);
xnor U712 (N_712,In_755,In_220);
xor U713 (N_713,In_194,In_68);
xnor U714 (N_714,In_945,In_655);
or U715 (N_715,In_758,In_237);
nand U716 (N_716,In_494,In_769);
nor U717 (N_717,In_447,In_21);
or U718 (N_718,In_186,In_346);
nand U719 (N_719,In_856,In_548);
nand U720 (N_720,In_19,In_527);
and U721 (N_721,In_135,In_8);
nor U722 (N_722,In_350,In_541);
and U723 (N_723,In_801,In_332);
or U724 (N_724,In_493,In_806);
or U725 (N_725,In_161,In_160);
nand U726 (N_726,In_969,In_775);
nand U727 (N_727,In_360,In_617);
nand U728 (N_728,In_380,In_568);
nor U729 (N_729,In_838,In_82);
and U730 (N_730,In_957,In_402);
nor U731 (N_731,In_895,In_673);
or U732 (N_732,In_369,In_861);
and U733 (N_733,In_320,In_905);
nand U734 (N_734,In_982,In_724);
nand U735 (N_735,In_181,In_120);
and U736 (N_736,In_401,In_881);
nor U737 (N_737,In_109,In_407);
nand U738 (N_738,In_990,In_746);
xnor U739 (N_739,In_172,In_283);
and U740 (N_740,In_838,In_815);
or U741 (N_741,In_681,In_472);
nand U742 (N_742,In_289,In_933);
xnor U743 (N_743,In_958,In_671);
or U744 (N_744,In_216,In_952);
and U745 (N_745,In_23,In_394);
or U746 (N_746,In_190,In_995);
or U747 (N_747,In_943,In_31);
and U748 (N_748,In_887,In_901);
nand U749 (N_749,In_967,In_547);
or U750 (N_750,In_948,In_607);
nand U751 (N_751,In_776,In_410);
nor U752 (N_752,In_385,In_826);
or U753 (N_753,In_52,In_11);
and U754 (N_754,In_252,In_638);
nor U755 (N_755,In_291,In_154);
nor U756 (N_756,In_654,In_343);
nand U757 (N_757,In_305,In_466);
nand U758 (N_758,In_6,In_896);
nor U759 (N_759,In_201,In_50);
nand U760 (N_760,In_673,In_211);
and U761 (N_761,In_667,In_760);
or U762 (N_762,In_751,In_25);
nand U763 (N_763,In_14,In_24);
and U764 (N_764,In_94,In_254);
and U765 (N_765,In_167,In_808);
nor U766 (N_766,In_39,In_304);
and U767 (N_767,In_396,In_264);
nand U768 (N_768,In_605,In_919);
or U769 (N_769,In_162,In_474);
and U770 (N_770,In_689,In_959);
or U771 (N_771,In_408,In_41);
xnor U772 (N_772,In_798,In_190);
nand U773 (N_773,In_181,In_980);
and U774 (N_774,In_843,In_13);
or U775 (N_775,In_910,In_8);
and U776 (N_776,In_472,In_136);
nor U777 (N_777,In_425,In_932);
and U778 (N_778,In_878,In_296);
or U779 (N_779,In_298,In_609);
nor U780 (N_780,In_652,In_933);
and U781 (N_781,In_336,In_345);
and U782 (N_782,In_932,In_79);
or U783 (N_783,In_905,In_271);
and U784 (N_784,In_900,In_912);
nand U785 (N_785,In_284,In_654);
xor U786 (N_786,In_69,In_157);
or U787 (N_787,In_943,In_746);
and U788 (N_788,In_137,In_281);
nand U789 (N_789,In_373,In_825);
xor U790 (N_790,In_408,In_201);
or U791 (N_791,In_381,In_663);
nand U792 (N_792,In_375,In_683);
nand U793 (N_793,In_537,In_396);
and U794 (N_794,In_174,In_788);
xnor U795 (N_795,In_135,In_304);
nor U796 (N_796,In_0,In_306);
nor U797 (N_797,In_301,In_284);
nor U798 (N_798,In_97,In_20);
nand U799 (N_799,In_91,In_396);
nor U800 (N_800,In_124,In_924);
nand U801 (N_801,In_993,In_857);
and U802 (N_802,In_276,In_308);
and U803 (N_803,In_249,In_493);
nand U804 (N_804,In_497,In_511);
nand U805 (N_805,In_205,In_985);
nor U806 (N_806,In_795,In_219);
and U807 (N_807,In_57,In_2);
and U808 (N_808,In_684,In_708);
and U809 (N_809,In_586,In_103);
nor U810 (N_810,In_234,In_559);
and U811 (N_811,In_362,In_20);
and U812 (N_812,In_777,In_916);
or U813 (N_813,In_358,In_100);
xor U814 (N_814,In_370,In_793);
nor U815 (N_815,In_717,In_219);
or U816 (N_816,In_925,In_948);
or U817 (N_817,In_711,In_827);
nor U818 (N_818,In_851,In_965);
or U819 (N_819,In_668,In_542);
nor U820 (N_820,In_88,In_422);
or U821 (N_821,In_560,In_122);
nor U822 (N_822,In_755,In_711);
and U823 (N_823,In_931,In_605);
nand U824 (N_824,In_570,In_21);
and U825 (N_825,In_341,In_515);
and U826 (N_826,In_106,In_449);
and U827 (N_827,In_701,In_914);
nor U828 (N_828,In_175,In_68);
and U829 (N_829,In_323,In_762);
nand U830 (N_830,In_601,In_235);
nand U831 (N_831,In_286,In_864);
nand U832 (N_832,In_35,In_754);
nor U833 (N_833,In_760,In_764);
nor U834 (N_834,In_246,In_633);
nand U835 (N_835,In_750,In_765);
nor U836 (N_836,In_468,In_341);
or U837 (N_837,In_522,In_230);
and U838 (N_838,In_577,In_515);
nand U839 (N_839,In_245,In_163);
xnor U840 (N_840,In_584,In_7);
and U841 (N_841,In_53,In_488);
and U842 (N_842,In_437,In_661);
nor U843 (N_843,In_767,In_50);
nor U844 (N_844,In_25,In_653);
or U845 (N_845,In_369,In_483);
xor U846 (N_846,In_766,In_702);
and U847 (N_847,In_849,In_25);
nor U848 (N_848,In_129,In_193);
nand U849 (N_849,In_960,In_812);
or U850 (N_850,In_743,In_50);
and U851 (N_851,In_199,In_699);
or U852 (N_852,In_286,In_355);
nand U853 (N_853,In_206,In_132);
or U854 (N_854,In_16,In_201);
xnor U855 (N_855,In_574,In_899);
nor U856 (N_856,In_759,In_932);
nor U857 (N_857,In_93,In_471);
or U858 (N_858,In_425,In_575);
nor U859 (N_859,In_209,In_68);
nor U860 (N_860,In_453,In_894);
or U861 (N_861,In_625,In_648);
nand U862 (N_862,In_604,In_194);
nand U863 (N_863,In_673,In_526);
and U864 (N_864,In_159,In_833);
or U865 (N_865,In_799,In_868);
xnor U866 (N_866,In_216,In_104);
nand U867 (N_867,In_382,In_671);
or U868 (N_868,In_949,In_379);
nand U869 (N_869,In_312,In_333);
nand U870 (N_870,In_547,In_667);
nand U871 (N_871,In_823,In_119);
or U872 (N_872,In_806,In_979);
xor U873 (N_873,In_417,In_657);
nand U874 (N_874,In_32,In_664);
or U875 (N_875,In_928,In_707);
and U876 (N_876,In_241,In_835);
and U877 (N_877,In_478,In_502);
and U878 (N_878,In_989,In_376);
nor U879 (N_879,In_952,In_767);
xnor U880 (N_880,In_666,In_346);
or U881 (N_881,In_346,In_912);
and U882 (N_882,In_443,In_995);
nand U883 (N_883,In_141,In_871);
nor U884 (N_884,In_218,In_729);
or U885 (N_885,In_437,In_780);
nand U886 (N_886,In_641,In_700);
or U887 (N_887,In_303,In_782);
nor U888 (N_888,In_872,In_321);
and U889 (N_889,In_21,In_230);
nor U890 (N_890,In_165,In_374);
or U891 (N_891,In_95,In_375);
nor U892 (N_892,In_103,In_159);
nor U893 (N_893,In_916,In_486);
or U894 (N_894,In_276,In_235);
nand U895 (N_895,In_553,In_991);
nor U896 (N_896,In_529,In_68);
or U897 (N_897,In_741,In_155);
and U898 (N_898,In_981,In_748);
nand U899 (N_899,In_207,In_826);
nor U900 (N_900,In_153,In_166);
nand U901 (N_901,In_389,In_718);
and U902 (N_902,In_851,In_617);
and U903 (N_903,In_273,In_810);
or U904 (N_904,In_762,In_407);
and U905 (N_905,In_878,In_567);
and U906 (N_906,In_521,In_24);
nor U907 (N_907,In_775,In_295);
and U908 (N_908,In_491,In_798);
xnor U909 (N_909,In_691,In_412);
nand U910 (N_910,In_650,In_961);
xnor U911 (N_911,In_306,In_957);
and U912 (N_912,In_628,In_367);
xor U913 (N_913,In_370,In_208);
nor U914 (N_914,In_963,In_548);
nor U915 (N_915,In_910,In_31);
nor U916 (N_916,In_169,In_297);
and U917 (N_917,In_3,In_606);
or U918 (N_918,In_220,In_153);
or U919 (N_919,In_543,In_660);
nand U920 (N_920,In_18,In_803);
xnor U921 (N_921,In_88,In_940);
nor U922 (N_922,In_930,In_815);
nand U923 (N_923,In_486,In_309);
nand U924 (N_924,In_462,In_387);
nor U925 (N_925,In_965,In_870);
or U926 (N_926,In_733,In_428);
and U927 (N_927,In_671,In_361);
or U928 (N_928,In_134,In_86);
nor U929 (N_929,In_274,In_392);
and U930 (N_930,In_41,In_128);
and U931 (N_931,In_801,In_779);
or U932 (N_932,In_102,In_830);
nand U933 (N_933,In_974,In_415);
nor U934 (N_934,In_239,In_528);
and U935 (N_935,In_847,In_323);
or U936 (N_936,In_512,In_765);
nand U937 (N_937,In_232,In_428);
xnor U938 (N_938,In_209,In_398);
nand U939 (N_939,In_975,In_694);
nand U940 (N_940,In_991,In_871);
and U941 (N_941,In_189,In_991);
nor U942 (N_942,In_23,In_111);
and U943 (N_943,In_605,In_193);
or U944 (N_944,In_936,In_19);
or U945 (N_945,In_961,In_353);
nor U946 (N_946,In_721,In_929);
nand U947 (N_947,In_829,In_478);
nand U948 (N_948,In_572,In_823);
and U949 (N_949,In_174,In_965);
xnor U950 (N_950,In_805,In_552);
and U951 (N_951,In_437,In_223);
xor U952 (N_952,In_270,In_425);
nor U953 (N_953,In_336,In_663);
nand U954 (N_954,In_313,In_178);
nor U955 (N_955,In_964,In_811);
or U956 (N_956,In_721,In_887);
nor U957 (N_957,In_761,In_591);
and U958 (N_958,In_813,In_649);
nor U959 (N_959,In_952,In_934);
or U960 (N_960,In_249,In_189);
nand U961 (N_961,In_267,In_673);
xnor U962 (N_962,In_522,In_276);
and U963 (N_963,In_505,In_267);
or U964 (N_964,In_477,In_474);
or U965 (N_965,In_988,In_264);
and U966 (N_966,In_686,In_1);
nor U967 (N_967,In_151,In_236);
or U968 (N_968,In_631,In_378);
nor U969 (N_969,In_437,In_206);
nor U970 (N_970,In_836,In_107);
and U971 (N_971,In_400,In_218);
nor U972 (N_972,In_755,In_531);
xor U973 (N_973,In_518,In_634);
and U974 (N_974,In_860,In_494);
nand U975 (N_975,In_515,In_258);
nor U976 (N_976,In_382,In_983);
nand U977 (N_977,In_693,In_125);
and U978 (N_978,In_696,In_426);
nand U979 (N_979,In_740,In_475);
nand U980 (N_980,In_493,In_934);
nand U981 (N_981,In_142,In_930);
or U982 (N_982,In_638,In_73);
and U983 (N_983,In_108,In_429);
xor U984 (N_984,In_357,In_482);
and U985 (N_985,In_549,In_271);
and U986 (N_986,In_288,In_330);
or U987 (N_987,In_517,In_394);
or U988 (N_988,In_954,In_392);
and U989 (N_989,In_828,In_842);
xnor U990 (N_990,In_927,In_319);
nand U991 (N_991,In_426,In_421);
nand U992 (N_992,In_422,In_599);
nand U993 (N_993,In_486,In_109);
and U994 (N_994,In_409,In_136);
xnor U995 (N_995,In_829,In_750);
nand U996 (N_996,In_777,In_330);
xor U997 (N_997,In_756,In_1);
or U998 (N_998,In_875,In_418);
nor U999 (N_999,In_534,In_888);
or U1000 (N_1000,In_754,In_935);
and U1001 (N_1001,In_308,In_714);
nand U1002 (N_1002,In_192,In_140);
and U1003 (N_1003,In_901,In_497);
nor U1004 (N_1004,In_572,In_25);
nand U1005 (N_1005,In_572,In_643);
nand U1006 (N_1006,In_442,In_114);
nand U1007 (N_1007,In_479,In_874);
or U1008 (N_1008,In_586,In_347);
or U1009 (N_1009,In_727,In_671);
or U1010 (N_1010,In_753,In_279);
or U1011 (N_1011,In_103,In_995);
nor U1012 (N_1012,In_587,In_157);
or U1013 (N_1013,In_412,In_103);
or U1014 (N_1014,In_993,In_874);
nand U1015 (N_1015,In_829,In_98);
nor U1016 (N_1016,In_149,In_733);
xnor U1017 (N_1017,In_451,In_890);
and U1018 (N_1018,In_913,In_517);
xnor U1019 (N_1019,In_251,In_779);
nor U1020 (N_1020,In_549,In_84);
and U1021 (N_1021,In_229,In_904);
nand U1022 (N_1022,In_678,In_953);
nor U1023 (N_1023,In_689,In_144);
nand U1024 (N_1024,In_511,In_542);
nor U1025 (N_1025,In_490,In_37);
nor U1026 (N_1026,In_473,In_670);
and U1027 (N_1027,In_203,In_168);
nor U1028 (N_1028,In_760,In_116);
xnor U1029 (N_1029,In_293,In_163);
and U1030 (N_1030,In_615,In_830);
or U1031 (N_1031,In_745,In_67);
and U1032 (N_1032,In_440,In_288);
nor U1033 (N_1033,In_39,In_62);
or U1034 (N_1034,In_548,In_717);
and U1035 (N_1035,In_731,In_276);
or U1036 (N_1036,In_413,In_401);
or U1037 (N_1037,In_408,In_407);
nand U1038 (N_1038,In_271,In_990);
nand U1039 (N_1039,In_782,In_230);
or U1040 (N_1040,In_705,In_222);
xnor U1041 (N_1041,In_942,In_201);
or U1042 (N_1042,In_174,In_736);
nand U1043 (N_1043,In_352,In_856);
or U1044 (N_1044,In_1,In_381);
and U1045 (N_1045,In_213,In_194);
and U1046 (N_1046,In_354,In_778);
nor U1047 (N_1047,In_529,In_495);
or U1048 (N_1048,In_389,In_527);
nand U1049 (N_1049,In_385,In_545);
and U1050 (N_1050,In_549,In_565);
nor U1051 (N_1051,In_888,In_881);
nand U1052 (N_1052,In_57,In_716);
nor U1053 (N_1053,In_782,In_461);
or U1054 (N_1054,In_652,In_82);
or U1055 (N_1055,In_437,In_875);
nand U1056 (N_1056,In_248,In_387);
nand U1057 (N_1057,In_149,In_242);
nand U1058 (N_1058,In_650,In_921);
xnor U1059 (N_1059,In_638,In_776);
nor U1060 (N_1060,In_793,In_258);
nand U1061 (N_1061,In_594,In_716);
nor U1062 (N_1062,In_396,In_605);
or U1063 (N_1063,In_561,In_576);
nand U1064 (N_1064,In_502,In_338);
xor U1065 (N_1065,In_433,In_113);
nor U1066 (N_1066,In_391,In_724);
xor U1067 (N_1067,In_906,In_329);
nor U1068 (N_1068,In_795,In_766);
nor U1069 (N_1069,In_933,In_59);
nand U1070 (N_1070,In_838,In_358);
and U1071 (N_1071,In_391,In_604);
nand U1072 (N_1072,In_475,In_250);
and U1073 (N_1073,In_667,In_874);
xnor U1074 (N_1074,In_893,In_113);
nand U1075 (N_1075,In_587,In_327);
xnor U1076 (N_1076,In_220,In_924);
or U1077 (N_1077,In_180,In_90);
nand U1078 (N_1078,In_355,In_936);
nor U1079 (N_1079,In_350,In_721);
nor U1080 (N_1080,In_194,In_953);
nor U1081 (N_1081,In_30,In_373);
nand U1082 (N_1082,In_623,In_356);
or U1083 (N_1083,In_416,In_712);
or U1084 (N_1084,In_390,In_953);
xor U1085 (N_1085,In_655,In_335);
nand U1086 (N_1086,In_949,In_441);
or U1087 (N_1087,In_196,In_827);
nand U1088 (N_1088,In_692,In_580);
nand U1089 (N_1089,In_564,In_781);
nand U1090 (N_1090,In_474,In_57);
and U1091 (N_1091,In_945,In_661);
nand U1092 (N_1092,In_242,In_127);
or U1093 (N_1093,In_498,In_562);
or U1094 (N_1094,In_53,In_249);
xor U1095 (N_1095,In_283,In_862);
or U1096 (N_1096,In_229,In_79);
and U1097 (N_1097,In_231,In_3);
and U1098 (N_1098,In_557,In_979);
or U1099 (N_1099,In_301,In_183);
or U1100 (N_1100,In_173,In_581);
nand U1101 (N_1101,In_10,In_9);
nor U1102 (N_1102,In_608,In_907);
nor U1103 (N_1103,In_282,In_924);
nand U1104 (N_1104,In_417,In_820);
or U1105 (N_1105,In_780,In_363);
and U1106 (N_1106,In_837,In_103);
xor U1107 (N_1107,In_200,In_260);
or U1108 (N_1108,In_194,In_677);
nand U1109 (N_1109,In_409,In_807);
or U1110 (N_1110,In_426,In_816);
nand U1111 (N_1111,In_600,In_376);
nand U1112 (N_1112,In_186,In_974);
nor U1113 (N_1113,In_313,In_167);
and U1114 (N_1114,In_977,In_70);
nand U1115 (N_1115,In_72,In_712);
nand U1116 (N_1116,In_988,In_747);
nor U1117 (N_1117,In_552,In_194);
or U1118 (N_1118,In_311,In_295);
nor U1119 (N_1119,In_405,In_436);
nor U1120 (N_1120,In_275,In_814);
nor U1121 (N_1121,In_135,In_197);
xor U1122 (N_1122,In_242,In_451);
or U1123 (N_1123,In_435,In_693);
or U1124 (N_1124,In_976,In_486);
or U1125 (N_1125,In_109,In_360);
xnor U1126 (N_1126,In_840,In_220);
and U1127 (N_1127,In_985,In_518);
or U1128 (N_1128,In_529,In_84);
nor U1129 (N_1129,In_691,In_900);
nand U1130 (N_1130,In_754,In_822);
and U1131 (N_1131,In_446,In_673);
nor U1132 (N_1132,In_36,In_863);
nor U1133 (N_1133,In_538,In_785);
or U1134 (N_1134,In_975,In_424);
nand U1135 (N_1135,In_169,In_560);
and U1136 (N_1136,In_356,In_483);
and U1137 (N_1137,In_173,In_520);
or U1138 (N_1138,In_83,In_722);
xnor U1139 (N_1139,In_501,In_7);
nor U1140 (N_1140,In_111,In_347);
and U1141 (N_1141,In_863,In_508);
nor U1142 (N_1142,In_418,In_313);
or U1143 (N_1143,In_393,In_671);
nand U1144 (N_1144,In_94,In_108);
and U1145 (N_1145,In_493,In_739);
or U1146 (N_1146,In_748,In_84);
nor U1147 (N_1147,In_845,In_284);
and U1148 (N_1148,In_967,In_308);
nor U1149 (N_1149,In_196,In_693);
nand U1150 (N_1150,In_385,In_723);
nor U1151 (N_1151,In_451,In_751);
and U1152 (N_1152,In_813,In_580);
nor U1153 (N_1153,In_910,In_975);
nand U1154 (N_1154,In_966,In_419);
and U1155 (N_1155,In_296,In_134);
nor U1156 (N_1156,In_894,In_216);
or U1157 (N_1157,In_87,In_651);
or U1158 (N_1158,In_262,In_527);
and U1159 (N_1159,In_459,In_209);
nand U1160 (N_1160,In_89,In_479);
or U1161 (N_1161,In_207,In_910);
or U1162 (N_1162,In_244,In_908);
nor U1163 (N_1163,In_474,In_75);
and U1164 (N_1164,In_328,In_277);
and U1165 (N_1165,In_975,In_92);
nor U1166 (N_1166,In_528,In_857);
xnor U1167 (N_1167,In_614,In_885);
or U1168 (N_1168,In_571,In_68);
xnor U1169 (N_1169,In_495,In_341);
nand U1170 (N_1170,In_443,In_825);
nand U1171 (N_1171,In_229,In_889);
or U1172 (N_1172,In_877,In_298);
or U1173 (N_1173,In_526,In_442);
nand U1174 (N_1174,In_679,In_471);
or U1175 (N_1175,In_945,In_51);
nand U1176 (N_1176,In_366,In_838);
xor U1177 (N_1177,In_460,In_413);
nand U1178 (N_1178,In_699,In_168);
and U1179 (N_1179,In_440,In_968);
and U1180 (N_1180,In_420,In_674);
nand U1181 (N_1181,In_173,In_572);
nand U1182 (N_1182,In_451,In_196);
or U1183 (N_1183,In_529,In_916);
nand U1184 (N_1184,In_376,In_335);
nor U1185 (N_1185,In_780,In_309);
nor U1186 (N_1186,In_216,In_744);
nand U1187 (N_1187,In_339,In_160);
nand U1188 (N_1188,In_186,In_991);
or U1189 (N_1189,In_83,In_614);
and U1190 (N_1190,In_59,In_199);
or U1191 (N_1191,In_930,In_648);
or U1192 (N_1192,In_283,In_92);
xnor U1193 (N_1193,In_23,In_570);
and U1194 (N_1194,In_696,In_167);
nand U1195 (N_1195,In_665,In_520);
nand U1196 (N_1196,In_907,In_622);
and U1197 (N_1197,In_158,In_675);
nor U1198 (N_1198,In_27,In_421);
and U1199 (N_1199,In_310,In_889);
nor U1200 (N_1200,In_600,In_355);
nor U1201 (N_1201,In_261,In_320);
and U1202 (N_1202,In_742,In_534);
or U1203 (N_1203,In_649,In_969);
nor U1204 (N_1204,In_238,In_68);
and U1205 (N_1205,In_405,In_611);
nand U1206 (N_1206,In_19,In_830);
and U1207 (N_1207,In_133,In_244);
nor U1208 (N_1208,In_140,In_443);
nand U1209 (N_1209,In_96,In_645);
and U1210 (N_1210,In_638,In_701);
xnor U1211 (N_1211,In_824,In_468);
and U1212 (N_1212,In_422,In_81);
and U1213 (N_1213,In_506,In_88);
nand U1214 (N_1214,In_926,In_919);
xnor U1215 (N_1215,In_876,In_5);
or U1216 (N_1216,In_794,In_881);
nand U1217 (N_1217,In_235,In_163);
and U1218 (N_1218,In_715,In_362);
nand U1219 (N_1219,In_994,In_224);
nand U1220 (N_1220,In_594,In_938);
nor U1221 (N_1221,In_967,In_386);
or U1222 (N_1222,In_346,In_766);
or U1223 (N_1223,In_364,In_847);
and U1224 (N_1224,In_932,In_541);
nand U1225 (N_1225,In_648,In_447);
xor U1226 (N_1226,In_167,In_109);
nor U1227 (N_1227,In_702,In_634);
and U1228 (N_1228,In_388,In_447);
or U1229 (N_1229,In_290,In_169);
and U1230 (N_1230,In_556,In_584);
nand U1231 (N_1231,In_125,In_715);
nor U1232 (N_1232,In_989,In_832);
and U1233 (N_1233,In_840,In_376);
nand U1234 (N_1234,In_780,In_95);
nand U1235 (N_1235,In_874,In_141);
xnor U1236 (N_1236,In_676,In_344);
or U1237 (N_1237,In_942,In_508);
nor U1238 (N_1238,In_175,In_207);
nand U1239 (N_1239,In_864,In_108);
or U1240 (N_1240,In_506,In_438);
or U1241 (N_1241,In_163,In_275);
and U1242 (N_1242,In_287,In_301);
nand U1243 (N_1243,In_132,In_283);
nor U1244 (N_1244,In_43,In_263);
and U1245 (N_1245,In_970,In_663);
or U1246 (N_1246,In_471,In_203);
and U1247 (N_1247,In_484,In_561);
and U1248 (N_1248,In_478,In_467);
nor U1249 (N_1249,In_659,In_9);
nand U1250 (N_1250,In_512,In_706);
nor U1251 (N_1251,In_288,In_578);
nand U1252 (N_1252,In_646,In_165);
and U1253 (N_1253,In_859,In_306);
or U1254 (N_1254,In_82,In_526);
nand U1255 (N_1255,In_229,In_9);
nand U1256 (N_1256,In_615,In_652);
and U1257 (N_1257,In_443,In_361);
or U1258 (N_1258,In_824,In_528);
xnor U1259 (N_1259,In_328,In_275);
nor U1260 (N_1260,In_368,In_411);
nor U1261 (N_1261,In_865,In_345);
nand U1262 (N_1262,In_771,In_570);
nand U1263 (N_1263,In_58,In_981);
nor U1264 (N_1264,In_196,In_279);
nor U1265 (N_1265,In_622,In_744);
nor U1266 (N_1266,In_896,In_452);
or U1267 (N_1267,In_179,In_52);
or U1268 (N_1268,In_578,In_574);
nand U1269 (N_1269,In_941,In_698);
nand U1270 (N_1270,In_251,In_501);
and U1271 (N_1271,In_698,In_194);
nand U1272 (N_1272,In_805,In_135);
nand U1273 (N_1273,In_928,In_680);
nor U1274 (N_1274,In_351,In_941);
xnor U1275 (N_1275,In_837,In_248);
and U1276 (N_1276,In_424,In_777);
xnor U1277 (N_1277,In_997,In_462);
nor U1278 (N_1278,In_249,In_875);
or U1279 (N_1279,In_381,In_62);
xor U1280 (N_1280,In_578,In_752);
and U1281 (N_1281,In_725,In_38);
nand U1282 (N_1282,In_701,In_822);
xor U1283 (N_1283,In_153,In_348);
and U1284 (N_1284,In_571,In_954);
nand U1285 (N_1285,In_920,In_466);
nor U1286 (N_1286,In_965,In_96);
nand U1287 (N_1287,In_446,In_71);
and U1288 (N_1288,In_423,In_477);
nand U1289 (N_1289,In_558,In_153);
or U1290 (N_1290,In_302,In_688);
and U1291 (N_1291,In_156,In_410);
and U1292 (N_1292,In_190,In_745);
or U1293 (N_1293,In_796,In_241);
nand U1294 (N_1294,In_415,In_497);
nor U1295 (N_1295,In_732,In_731);
nor U1296 (N_1296,In_122,In_923);
and U1297 (N_1297,In_493,In_902);
and U1298 (N_1298,In_474,In_951);
nand U1299 (N_1299,In_420,In_329);
nand U1300 (N_1300,In_689,In_217);
nand U1301 (N_1301,In_7,In_317);
nor U1302 (N_1302,In_966,In_449);
xor U1303 (N_1303,In_154,In_580);
and U1304 (N_1304,In_634,In_574);
and U1305 (N_1305,In_542,In_759);
and U1306 (N_1306,In_157,In_824);
nand U1307 (N_1307,In_440,In_364);
nor U1308 (N_1308,In_82,In_168);
or U1309 (N_1309,In_880,In_63);
xor U1310 (N_1310,In_96,In_501);
xnor U1311 (N_1311,In_562,In_647);
xor U1312 (N_1312,In_827,In_453);
nand U1313 (N_1313,In_0,In_548);
nor U1314 (N_1314,In_786,In_246);
nand U1315 (N_1315,In_714,In_25);
or U1316 (N_1316,In_393,In_92);
nor U1317 (N_1317,In_252,In_176);
and U1318 (N_1318,In_271,In_176);
or U1319 (N_1319,In_403,In_520);
xnor U1320 (N_1320,In_457,In_322);
nand U1321 (N_1321,In_487,In_763);
or U1322 (N_1322,In_561,In_672);
and U1323 (N_1323,In_911,In_905);
and U1324 (N_1324,In_243,In_275);
and U1325 (N_1325,In_729,In_180);
or U1326 (N_1326,In_570,In_343);
xnor U1327 (N_1327,In_993,In_624);
nand U1328 (N_1328,In_366,In_471);
nor U1329 (N_1329,In_353,In_296);
nand U1330 (N_1330,In_25,In_124);
or U1331 (N_1331,In_904,In_178);
nor U1332 (N_1332,In_971,In_944);
or U1333 (N_1333,In_869,In_377);
xor U1334 (N_1334,In_859,In_475);
and U1335 (N_1335,In_932,In_303);
nor U1336 (N_1336,In_466,In_875);
nor U1337 (N_1337,In_151,In_447);
or U1338 (N_1338,In_177,In_139);
xnor U1339 (N_1339,In_973,In_270);
or U1340 (N_1340,In_754,In_968);
or U1341 (N_1341,In_307,In_656);
or U1342 (N_1342,In_610,In_211);
xnor U1343 (N_1343,In_771,In_467);
xnor U1344 (N_1344,In_383,In_688);
nand U1345 (N_1345,In_157,In_607);
or U1346 (N_1346,In_265,In_310);
and U1347 (N_1347,In_230,In_501);
nor U1348 (N_1348,In_539,In_289);
nand U1349 (N_1349,In_707,In_520);
nor U1350 (N_1350,In_180,In_67);
nor U1351 (N_1351,In_33,In_801);
nor U1352 (N_1352,In_690,In_715);
nor U1353 (N_1353,In_109,In_216);
xor U1354 (N_1354,In_187,In_805);
nor U1355 (N_1355,In_727,In_218);
nand U1356 (N_1356,In_172,In_552);
nor U1357 (N_1357,In_577,In_383);
xor U1358 (N_1358,In_142,In_51);
and U1359 (N_1359,In_608,In_67);
and U1360 (N_1360,In_874,In_577);
nor U1361 (N_1361,In_101,In_595);
and U1362 (N_1362,In_118,In_747);
xor U1363 (N_1363,In_910,In_996);
nand U1364 (N_1364,In_929,In_561);
nand U1365 (N_1365,In_845,In_917);
or U1366 (N_1366,In_912,In_325);
nor U1367 (N_1367,In_149,In_765);
or U1368 (N_1368,In_870,In_343);
or U1369 (N_1369,In_394,In_273);
nor U1370 (N_1370,In_316,In_556);
nor U1371 (N_1371,In_835,In_403);
nand U1372 (N_1372,In_915,In_52);
nor U1373 (N_1373,In_354,In_903);
nand U1374 (N_1374,In_884,In_278);
or U1375 (N_1375,In_480,In_392);
or U1376 (N_1376,In_724,In_475);
nor U1377 (N_1377,In_346,In_308);
nand U1378 (N_1378,In_768,In_939);
and U1379 (N_1379,In_143,In_365);
nand U1380 (N_1380,In_570,In_358);
and U1381 (N_1381,In_130,In_526);
and U1382 (N_1382,In_291,In_854);
or U1383 (N_1383,In_877,In_881);
nand U1384 (N_1384,In_351,In_733);
or U1385 (N_1385,In_791,In_20);
or U1386 (N_1386,In_596,In_347);
and U1387 (N_1387,In_448,In_340);
nor U1388 (N_1388,In_535,In_51);
nor U1389 (N_1389,In_289,In_172);
nor U1390 (N_1390,In_559,In_293);
nor U1391 (N_1391,In_158,In_136);
or U1392 (N_1392,In_532,In_437);
and U1393 (N_1393,In_509,In_407);
nand U1394 (N_1394,In_9,In_755);
or U1395 (N_1395,In_853,In_205);
and U1396 (N_1396,In_478,In_20);
xor U1397 (N_1397,In_536,In_561);
or U1398 (N_1398,In_986,In_410);
and U1399 (N_1399,In_544,In_849);
and U1400 (N_1400,In_115,In_73);
and U1401 (N_1401,In_1,In_517);
nand U1402 (N_1402,In_834,In_761);
nor U1403 (N_1403,In_537,In_202);
or U1404 (N_1404,In_616,In_973);
and U1405 (N_1405,In_814,In_269);
xor U1406 (N_1406,In_440,In_305);
nand U1407 (N_1407,In_292,In_685);
nand U1408 (N_1408,In_424,In_161);
or U1409 (N_1409,In_568,In_444);
nor U1410 (N_1410,In_794,In_724);
nand U1411 (N_1411,In_137,In_412);
or U1412 (N_1412,In_250,In_0);
or U1413 (N_1413,In_596,In_503);
xnor U1414 (N_1414,In_578,In_57);
and U1415 (N_1415,In_306,In_329);
nor U1416 (N_1416,In_906,In_240);
and U1417 (N_1417,In_470,In_531);
nor U1418 (N_1418,In_296,In_954);
xnor U1419 (N_1419,In_745,In_382);
or U1420 (N_1420,In_480,In_306);
xnor U1421 (N_1421,In_849,In_930);
and U1422 (N_1422,In_140,In_101);
xor U1423 (N_1423,In_782,In_264);
nand U1424 (N_1424,In_512,In_986);
xnor U1425 (N_1425,In_623,In_865);
or U1426 (N_1426,In_581,In_751);
and U1427 (N_1427,In_198,In_713);
nand U1428 (N_1428,In_682,In_70);
or U1429 (N_1429,In_50,In_493);
and U1430 (N_1430,In_807,In_728);
nand U1431 (N_1431,In_803,In_592);
nand U1432 (N_1432,In_44,In_468);
nand U1433 (N_1433,In_771,In_752);
xor U1434 (N_1434,In_991,In_148);
nor U1435 (N_1435,In_773,In_524);
or U1436 (N_1436,In_523,In_800);
and U1437 (N_1437,In_593,In_390);
and U1438 (N_1438,In_572,In_347);
nand U1439 (N_1439,In_216,In_781);
and U1440 (N_1440,In_423,In_365);
or U1441 (N_1441,In_22,In_925);
nor U1442 (N_1442,In_54,In_280);
nand U1443 (N_1443,In_284,In_935);
nor U1444 (N_1444,In_846,In_530);
nor U1445 (N_1445,In_23,In_805);
xor U1446 (N_1446,In_30,In_705);
nand U1447 (N_1447,In_563,In_769);
nor U1448 (N_1448,In_887,In_243);
and U1449 (N_1449,In_763,In_25);
nand U1450 (N_1450,In_370,In_417);
and U1451 (N_1451,In_142,In_150);
or U1452 (N_1452,In_350,In_611);
nand U1453 (N_1453,In_129,In_286);
or U1454 (N_1454,In_845,In_43);
nand U1455 (N_1455,In_560,In_958);
nand U1456 (N_1456,In_715,In_420);
and U1457 (N_1457,In_998,In_98);
or U1458 (N_1458,In_927,In_829);
xor U1459 (N_1459,In_388,In_997);
and U1460 (N_1460,In_417,In_137);
nand U1461 (N_1461,In_430,In_328);
xor U1462 (N_1462,In_231,In_182);
and U1463 (N_1463,In_182,In_222);
and U1464 (N_1464,In_965,In_115);
nand U1465 (N_1465,In_99,In_287);
or U1466 (N_1466,In_224,In_737);
nor U1467 (N_1467,In_756,In_552);
nor U1468 (N_1468,In_670,In_136);
xor U1469 (N_1469,In_770,In_363);
or U1470 (N_1470,In_173,In_889);
nand U1471 (N_1471,In_879,In_641);
nor U1472 (N_1472,In_441,In_246);
or U1473 (N_1473,In_768,In_251);
and U1474 (N_1474,In_710,In_750);
xor U1475 (N_1475,In_378,In_739);
nor U1476 (N_1476,In_571,In_677);
nand U1477 (N_1477,In_983,In_759);
or U1478 (N_1478,In_468,In_689);
and U1479 (N_1479,In_512,In_369);
xor U1480 (N_1480,In_976,In_947);
or U1481 (N_1481,In_461,In_109);
nand U1482 (N_1482,In_602,In_310);
or U1483 (N_1483,In_363,In_721);
and U1484 (N_1484,In_371,In_116);
nor U1485 (N_1485,In_217,In_242);
nor U1486 (N_1486,In_813,In_943);
nor U1487 (N_1487,In_408,In_172);
or U1488 (N_1488,In_529,In_254);
and U1489 (N_1489,In_409,In_676);
xnor U1490 (N_1490,In_198,In_845);
or U1491 (N_1491,In_677,In_167);
nor U1492 (N_1492,In_223,In_588);
xor U1493 (N_1493,In_201,In_156);
and U1494 (N_1494,In_957,In_65);
nand U1495 (N_1495,In_859,In_786);
or U1496 (N_1496,In_865,In_695);
and U1497 (N_1497,In_973,In_357);
and U1498 (N_1498,In_469,In_311);
and U1499 (N_1499,In_41,In_327);
nand U1500 (N_1500,In_208,In_191);
xnor U1501 (N_1501,In_145,In_22);
nor U1502 (N_1502,In_980,In_539);
nand U1503 (N_1503,In_178,In_937);
nand U1504 (N_1504,In_745,In_915);
and U1505 (N_1505,In_452,In_486);
nand U1506 (N_1506,In_280,In_563);
and U1507 (N_1507,In_692,In_225);
and U1508 (N_1508,In_200,In_362);
or U1509 (N_1509,In_583,In_22);
or U1510 (N_1510,In_295,In_83);
or U1511 (N_1511,In_407,In_991);
or U1512 (N_1512,In_666,In_676);
and U1513 (N_1513,In_638,In_736);
or U1514 (N_1514,In_718,In_422);
xnor U1515 (N_1515,In_665,In_796);
or U1516 (N_1516,In_414,In_706);
nor U1517 (N_1517,In_579,In_633);
or U1518 (N_1518,In_820,In_633);
nand U1519 (N_1519,In_286,In_669);
nand U1520 (N_1520,In_626,In_17);
and U1521 (N_1521,In_905,In_921);
xnor U1522 (N_1522,In_790,In_992);
xor U1523 (N_1523,In_341,In_427);
nand U1524 (N_1524,In_270,In_927);
or U1525 (N_1525,In_357,In_852);
nand U1526 (N_1526,In_216,In_512);
nand U1527 (N_1527,In_151,In_5);
nor U1528 (N_1528,In_889,In_562);
and U1529 (N_1529,In_342,In_952);
nor U1530 (N_1530,In_336,In_555);
or U1531 (N_1531,In_135,In_945);
or U1532 (N_1532,In_823,In_323);
or U1533 (N_1533,In_96,In_224);
and U1534 (N_1534,In_295,In_16);
and U1535 (N_1535,In_58,In_815);
or U1536 (N_1536,In_647,In_227);
and U1537 (N_1537,In_116,In_81);
nor U1538 (N_1538,In_491,In_309);
nor U1539 (N_1539,In_914,In_800);
nor U1540 (N_1540,In_930,In_927);
nor U1541 (N_1541,In_492,In_3);
or U1542 (N_1542,In_31,In_799);
nor U1543 (N_1543,In_86,In_725);
nand U1544 (N_1544,In_499,In_931);
nand U1545 (N_1545,In_167,In_127);
nor U1546 (N_1546,In_2,In_699);
nand U1547 (N_1547,In_52,In_658);
nand U1548 (N_1548,In_115,In_738);
nand U1549 (N_1549,In_21,In_440);
or U1550 (N_1550,In_931,In_488);
xnor U1551 (N_1551,In_892,In_645);
nand U1552 (N_1552,In_247,In_483);
and U1553 (N_1553,In_324,In_771);
nor U1554 (N_1554,In_456,In_644);
or U1555 (N_1555,In_134,In_154);
and U1556 (N_1556,In_700,In_965);
and U1557 (N_1557,In_673,In_239);
and U1558 (N_1558,In_548,In_792);
or U1559 (N_1559,In_266,In_494);
nor U1560 (N_1560,In_51,In_946);
or U1561 (N_1561,In_663,In_975);
or U1562 (N_1562,In_899,In_724);
or U1563 (N_1563,In_186,In_850);
or U1564 (N_1564,In_71,In_311);
or U1565 (N_1565,In_126,In_363);
and U1566 (N_1566,In_944,In_937);
nor U1567 (N_1567,In_205,In_517);
nor U1568 (N_1568,In_271,In_875);
nand U1569 (N_1569,In_380,In_511);
or U1570 (N_1570,In_819,In_3);
or U1571 (N_1571,In_842,In_92);
and U1572 (N_1572,In_796,In_908);
nor U1573 (N_1573,In_875,In_393);
nor U1574 (N_1574,In_540,In_641);
or U1575 (N_1575,In_32,In_205);
and U1576 (N_1576,In_730,In_374);
and U1577 (N_1577,In_680,In_996);
xor U1578 (N_1578,In_247,In_2);
nand U1579 (N_1579,In_328,In_138);
nand U1580 (N_1580,In_704,In_408);
nor U1581 (N_1581,In_548,In_466);
nand U1582 (N_1582,In_448,In_770);
nand U1583 (N_1583,In_932,In_670);
or U1584 (N_1584,In_430,In_471);
and U1585 (N_1585,In_483,In_375);
nand U1586 (N_1586,In_370,In_412);
xor U1587 (N_1587,In_105,In_756);
and U1588 (N_1588,In_364,In_179);
xor U1589 (N_1589,In_67,In_293);
xor U1590 (N_1590,In_457,In_965);
or U1591 (N_1591,In_595,In_289);
nand U1592 (N_1592,In_511,In_282);
nor U1593 (N_1593,In_792,In_760);
or U1594 (N_1594,In_812,In_106);
nor U1595 (N_1595,In_19,In_675);
xor U1596 (N_1596,In_371,In_255);
xnor U1597 (N_1597,In_874,In_867);
or U1598 (N_1598,In_710,In_517);
xor U1599 (N_1599,In_504,In_984);
xnor U1600 (N_1600,In_630,In_757);
and U1601 (N_1601,In_733,In_145);
nand U1602 (N_1602,In_503,In_779);
nor U1603 (N_1603,In_332,In_178);
nor U1604 (N_1604,In_176,In_548);
and U1605 (N_1605,In_923,In_507);
nor U1606 (N_1606,In_631,In_679);
and U1607 (N_1607,In_742,In_255);
and U1608 (N_1608,In_331,In_934);
or U1609 (N_1609,In_196,In_836);
xor U1610 (N_1610,In_108,In_323);
nor U1611 (N_1611,In_714,In_193);
or U1612 (N_1612,In_491,In_697);
nor U1613 (N_1613,In_593,In_305);
and U1614 (N_1614,In_792,In_557);
nand U1615 (N_1615,In_640,In_411);
nand U1616 (N_1616,In_548,In_854);
nor U1617 (N_1617,In_679,In_822);
nand U1618 (N_1618,In_971,In_961);
and U1619 (N_1619,In_451,In_730);
nor U1620 (N_1620,In_678,In_319);
nor U1621 (N_1621,In_622,In_512);
nor U1622 (N_1622,In_711,In_431);
or U1623 (N_1623,In_877,In_266);
or U1624 (N_1624,In_370,In_480);
and U1625 (N_1625,In_801,In_867);
or U1626 (N_1626,In_272,In_865);
and U1627 (N_1627,In_529,In_387);
nand U1628 (N_1628,In_62,In_764);
and U1629 (N_1629,In_45,In_658);
nand U1630 (N_1630,In_731,In_508);
nor U1631 (N_1631,In_422,In_325);
xor U1632 (N_1632,In_69,In_151);
nand U1633 (N_1633,In_268,In_333);
or U1634 (N_1634,In_415,In_856);
or U1635 (N_1635,In_284,In_157);
or U1636 (N_1636,In_204,In_714);
xnor U1637 (N_1637,In_541,In_721);
nand U1638 (N_1638,In_960,In_270);
nand U1639 (N_1639,In_524,In_489);
or U1640 (N_1640,In_597,In_777);
nor U1641 (N_1641,In_223,In_18);
nor U1642 (N_1642,In_277,In_257);
nor U1643 (N_1643,In_173,In_41);
nor U1644 (N_1644,In_528,In_947);
nor U1645 (N_1645,In_711,In_977);
nand U1646 (N_1646,In_309,In_11);
nand U1647 (N_1647,In_733,In_824);
xor U1648 (N_1648,In_709,In_780);
nand U1649 (N_1649,In_127,In_790);
nand U1650 (N_1650,In_269,In_939);
or U1651 (N_1651,In_558,In_422);
nand U1652 (N_1652,In_826,In_163);
nand U1653 (N_1653,In_316,In_685);
or U1654 (N_1654,In_442,In_262);
xnor U1655 (N_1655,In_447,In_669);
nor U1656 (N_1656,In_712,In_588);
nand U1657 (N_1657,In_66,In_968);
nand U1658 (N_1658,In_664,In_74);
or U1659 (N_1659,In_231,In_517);
nor U1660 (N_1660,In_18,In_267);
nor U1661 (N_1661,In_270,In_307);
or U1662 (N_1662,In_166,In_280);
nand U1663 (N_1663,In_960,In_203);
nand U1664 (N_1664,In_521,In_504);
nand U1665 (N_1665,In_78,In_902);
nor U1666 (N_1666,In_656,In_676);
nor U1667 (N_1667,In_325,In_21);
or U1668 (N_1668,In_727,In_143);
nand U1669 (N_1669,In_291,In_872);
nor U1670 (N_1670,In_438,In_971);
nor U1671 (N_1671,In_742,In_363);
or U1672 (N_1672,In_213,In_61);
and U1673 (N_1673,In_73,In_384);
or U1674 (N_1674,In_959,In_401);
or U1675 (N_1675,In_623,In_302);
and U1676 (N_1676,In_597,In_657);
nand U1677 (N_1677,In_239,In_778);
xor U1678 (N_1678,In_911,In_770);
nor U1679 (N_1679,In_478,In_490);
and U1680 (N_1680,In_935,In_447);
or U1681 (N_1681,In_750,In_61);
or U1682 (N_1682,In_675,In_128);
or U1683 (N_1683,In_810,In_269);
or U1684 (N_1684,In_376,In_578);
and U1685 (N_1685,In_615,In_51);
or U1686 (N_1686,In_482,In_314);
or U1687 (N_1687,In_353,In_473);
and U1688 (N_1688,In_111,In_865);
and U1689 (N_1689,In_348,In_511);
or U1690 (N_1690,In_89,In_611);
and U1691 (N_1691,In_691,In_865);
and U1692 (N_1692,In_443,In_200);
and U1693 (N_1693,In_630,In_427);
or U1694 (N_1694,In_687,In_43);
and U1695 (N_1695,In_970,In_703);
or U1696 (N_1696,In_56,In_324);
or U1697 (N_1697,In_100,In_522);
nand U1698 (N_1698,In_323,In_43);
nand U1699 (N_1699,In_989,In_243);
xnor U1700 (N_1700,In_452,In_932);
nor U1701 (N_1701,In_614,In_670);
nor U1702 (N_1702,In_5,In_611);
and U1703 (N_1703,In_199,In_66);
xnor U1704 (N_1704,In_79,In_227);
or U1705 (N_1705,In_263,In_154);
nor U1706 (N_1706,In_654,In_35);
nand U1707 (N_1707,In_832,In_439);
or U1708 (N_1708,In_269,In_178);
nor U1709 (N_1709,In_891,In_628);
nand U1710 (N_1710,In_663,In_229);
or U1711 (N_1711,In_587,In_541);
and U1712 (N_1712,In_711,In_481);
and U1713 (N_1713,In_982,In_894);
or U1714 (N_1714,In_368,In_499);
nand U1715 (N_1715,In_301,In_134);
nor U1716 (N_1716,In_938,In_574);
or U1717 (N_1717,In_999,In_328);
and U1718 (N_1718,In_417,In_933);
and U1719 (N_1719,In_747,In_990);
nor U1720 (N_1720,In_295,In_530);
and U1721 (N_1721,In_328,In_570);
nor U1722 (N_1722,In_980,In_617);
and U1723 (N_1723,In_294,In_53);
nor U1724 (N_1724,In_903,In_785);
nor U1725 (N_1725,In_979,In_639);
nand U1726 (N_1726,In_720,In_292);
and U1727 (N_1727,In_995,In_275);
and U1728 (N_1728,In_755,In_423);
nand U1729 (N_1729,In_70,In_823);
and U1730 (N_1730,In_973,In_384);
and U1731 (N_1731,In_100,In_933);
nand U1732 (N_1732,In_207,In_509);
nor U1733 (N_1733,In_584,In_815);
and U1734 (N_1734,In_739,In_455);
and U1735 (N_1735,In_111,In_532);
or U1736 (N_1736,In_205,In_455);
xor U1737 (N_1737,In_154,In_107);
xor U1738 (N_1738,In_854,In_678);
xnor U1739 (N_1739,In_242,In_58);
and U1740 (N_1740,In_388,In_225);
nor U1741 (N_1741,In_481,In_749);
nor U1742 (N_1742,In_12,In_120);
nand U1743 (N_1743,In_423,In_735);
nand U1744 (N_1744,In_146,In_114);
or U1745 (N_1745,In_694,In_638);
nor U1746 (N_1746,In_476,In_83);
xnor U1747 (N_1747,In_27,In_704);
or U1748 (N_1748,In_56,In_429);
nor U1749 (N_1749,In_592,In_961);
nor U1750 (N_1750,In_6,In_657);
and U1751 (N_1751,In_662,In_386);
nor U1752 (N_1752,In_602,In_163);
nor U1753 (N_1753,In_192,In_704);
nor U1754 (N_1754,In_885,In_233);
and U1755 (N_1755,In_616,In_805);
and U1756 (N_1756,In_568,In_797);
nand U1757 (N_1757,In_855,In_41);
nand U1758 (N_1758,In_730,In_731);
and U1759 (N_1759,In_986,In_706);
xnor U1760 (N_1760,In_766,In_598);
or U1761 (N_1761,In_932,In_994);
xnor U1762 (N_1762,In_340,In_878);
nor U1763 (N_1763,In_69,In_427);
nor U1764 (N_1764,In_201,In_664);
and U1765 (N_1765,In_858,In_302);
or U1766 (N_1766,In_840,In_349);
and U1767 (N_1767,In_855,In_102);
nand U1768 (N_1768,In_458,In_50);
and U1769 (N_1769,In_628,In_60);
or U1770 (N_1770,In_604,In_267);
nand U1771 (N_1771,In_754,In_780);
nand U1772 (N_1772,In_43,In_16);
nand U1773 (N_1773,In_550,In_579);
nor U1774 (N_1774,In_825,In_587);
nand U1775 (N_1775,In_341,In_238);
and U1776 (N_1776,In_41,In_874);
nor U1777 (N_1777,In_506,In_499);
and U1778 (N_1778,In_253,In_201);
or U1779 (N_1779,In_190,In_517);
xor U1780 (N_1780,In_202,In_953);
nand U1781 (N_1781,In_36,In_474);
or U1782 (N_1782,In_666,In_248);
xor U1783 (N_1783,In_303,In_415);
or U1784 (N_1784,In_418,In_512);
and U1785 (N_1785,In_693,In_351);
and U1786 (N_1786,In_619,In_905);
nor U1787 (N_1787,In_312,In_975);
nand U1788 (N_1788,In_612,In_616);
or U1789 (N_1789,In_625,In_793);
nand U1790 (N_1790,In_870,In_970);
nand U1791 (N_1791,In_992,In_880);
or U1792 (N_1792,In_750,In_521);
nor U1793 (N_1793,In_539,In_190);
or U1794 (N_1794,In_552,In_9);
and U1795 (N_1795,In_799,In_275);
and U1796 (N_1796,In_499,In_50);
nand U1797 (N_1797,In_139,In_290);
or U1798 (N_1798,In_649,In_365);
and U1799 (N_1799,In_644,In_364);
and U1800 (N_1800,In_150,In_421);
xnor U1801 (N_1801,In_333,In_873);
or U1802 (N_1802,In_832,In_758);
and U1803 (N_1803,In_360,In_560);
nand U1804 (N_1804,In_924,In_241);
nor U1805 (N_1805,In_948,In_310);
and U1806 (N_1806,In_283,In_118);
or U1807 (N_1807,In_117,In_404);
nand U1808 (N_1808,In_162,In_831);
or U1809 (N_1809,In_232,In_214);
nand U1810 (N_1810,In_341,In_823);
nand U1811 (N_1811,In_626,In_723);
nand U1812 (N_1812,In_643,In_155);
and U1813 (N_1813,In_925,In_754);
nand U1814 (N_1814,In_99,In_317);
and U1815 (N_1815,In_523,In_187);
nand U1816 (N_1816,In_652,In_804);
and U1817 (N_1817,In_195,In_0);
and U1818 (N_1818,In_437,In_246);
or U1819 (N_1819,In_885,In_513);
and U1820 (N_1820,In_48,In_126);
or U1821 (N_1821,In_363,In_113);
nand U1822 (N_1822,In_404,In_164);
nor U1823 (N_1823,In_59,In_133);
nand U1824 (N_1824,In_208,In_249);
and U1825 (N_1825,In_271,In_959);
and U1826 (N_1826,In_266,In_758);
and U1827 (N_1827,In_859,In_571);
xor U1828 (N_1828,In_150,In_895);
xnor U1829 (N_1829,In_11,In_637);
nor U1830 (N_1830,In_462,In_877);
nand U1831 (N_1831,In_651,In_710);
and U1832 (N_1832,In_404,In_90);
nand U1833 (N_1833,In_594,In_493);
nor U1834 (N_1834,In_195,In_201);
nand U1835 (N_1835,In_470,In_317);
or U1836 (N_1836,In_905,In_662);
and U1837 (N_1837,In_785,In_463);
or U1838 (N_1838,In_828,In_727);
nand U1839 (N_1839,In_431,In_445);
or U1840 (N_1840,In_946,In_93);
xnor U1841 (N_1841,In_316,In_77);
and U1842 (N_1842,In_547,In_94);
or U1843 (N_1843,In_474,In_774);
xor U1844 (N_1844,In_695,In_772);
or U1845 (N_1845,In_177,In_464);
nor U1846 (N_1846,In_416,In_322);
nand U1847 (N_1847,In_777,In_828);
nand U1848 (N_1848,In_352,In_27);
or U1849 (N_1849,In_805,In_631);
or U1850 (N_1850,In_598,In_63);
and U1851 (N_1851,In_439,In_90);
and U1852 (N_1852,In_818,In_4);
and U1853 (N_1853,In_763,In_501);
nand U1854 (N_1854,In_815,In_254);
nor U1855 (N_1855,In_436,In_246);
or U1856 (N_1856,In_665,In_991);
or U1857 (N_1857,In_137,In_47);
nand U1858 (N_1858,In_66,In_735);
nor U1859 (N_1859,In_438,In_585);
nor U1860 (N_1860,In_44,In_527);
and U1861 (N_1861,In_756,In_441);
xnor U1862 (N_1862,In_955,In_753);
or U1863 (N_1863,In_169,In_546);
nand U1864 (N_1864,In_89,In_764);
nor U1865 (N_1865,In_269,In_908);
or U1866 (N_1866,In_302,In_214);
or U1867 (N_1867,In_4,In_800);
nor U1868 (N_1868,In_419,In_682);
nor U1869 (N_1869,In_542,In_837);
nand U1870 (N_1870,In_729,In_621);
nor U1871 (N_1871,In_558,In_479);
nand U1872 (N_1872,In_286,In_906);
and U1873 (N_1873,In_298,In_492);
and U1874 (N_1874,In_243,In_488);
nand U1875 (N_1875,In_191,In_156);
nand U1876 (N_1876,In_899,In_382);
xnor U1877 (N_1877,In_655,In_309);
nor U1878 (N_1878,In_818,In_490);
xnor U1879 (N_1879,In_13,In_353);
nor U1880 (N_1880,In_94,In_292);
nor U1881 (N_1881,In_44,In_582);
or U1882 (N_1882,In_555,In_719);
or U1883 (N_1883,In_312,In_307);
nand U1884 (N_1884,In_535,In_592);
or U1885 (N_1885,In_475,In_537);
nor U1886 (N_1886,In_968,In_466);
nand U1887 (N_1887,In_790,In_734);
or U1888 (N_1888,In_481,In_637);
nor U1889 (N_1889,In_918,In_512);
and U1890 (N_1890,In_913,In_509);
and U1891 (N_1891,In_72,In_347);
nor U1892 (N_1892,In_269,In_572);
nand U1893 (N_1893,In_648,In_170);
nor U1894 (N_1894,In_499,In_844);
nor U1895 (N_1895,In_54,In_245);
and U1896 (N_1896,In_21,In_936);
xnor U1897 (N_1897,In_426,In_860);
nand U1898 (N_1898,In_785,In_969);
nand U1899 (N_1899,In_382,In_274);
nor U1900 (N_1900,In_731,In_372);
nor U1901 (N_1901,In_824,In_593);
nand U1902 (N_1902,In_854,In_661);
nand U1903 (N_1903,In_16,In_163);
or U1904 (N_1904,In_385,In_318);
nor U1905 (N_1905,In_671,In_40);
xnor U1906 (N_1906,In_529,In_206);
nor U1907 (N_1907,In_733,In_608);
nor U1908 (N_1908,In_664,In_738);
nor U1909 (N_1909,In_619,In_743);
and U1910 (N_1910,In_497,In_327);
or U1911 (N_1911,In_54,In_357);
or U1912 (N_1912,In_802,In_760);
and U1913 (N_1913,In_26,In_419);
or U1914 (N_1914,In_445,In_542);
nand U1915 (N_1915,In_275,In_448);
xor U1916 (N_1916,In_772,In_277);
or U1917 (N_1917,In_636,In_592);
nand U1918 (N_1918,In_824,In_608);
and U1919 (N_1919,In_823,In_360);
and U1920 (N_1920,In_507,In_568);
nand U1921 (N_1921,In_496,In_342);
nand U1922 (N_1922,In_921,In_909);
or U1923 (N_1923,In_520,In_269);
or U1924 (N_1924,In_800,In_243);
nor U1925 (N_1925,In_202,In_534);
or U1926 (N_1926,In_934,In_282);
and U1927 (N_1927,In_307,In_282);
or U1928 (N_1928,In_43,In_343);
nand U1929 (N_1929,In_120,In_858);
or U1930 (N_1930,In_787,In_290);
or U1931 (N_1931,In_339,In_156);
nor U1932 (N_1932,In_530,In_307);
and U1933 (N_1933,In_491,In_515);
or U1934 (N_1934,In_328,In_880);
or U1935 (N_1935,In_947,In_267);
xor U1936 (N_1936,In_591,In_733);
and U1937 (N_1937,In_621,In_326);
or U1938 (N_1938,In_923,In_780);
nand U1939 (N_1939,In_539,In_717);
nor U1940 (N_1940,In_72,In_703);
and U1941 (N_1941,In_660,In_754);
nor U1942 (N_1942,In_816,In_864);
nand U1943 (N_1943,In_246,In_157);
and U1944 (N_1944,In_701,In_472);
and U1945 (N_1945,In_792,In_820);
or U1946 (N_1946,In_197,In_214);
xnor U1947 (N_1947,In_436,In_883);
and U1948 (N_1948,In_704,In_733);
nor U1949 (N_1949,In_676,In_274);
or U1950 (N_1950,In_184,In_997);
xor U1951 (N_1951,In_109,In_27);
nor U1952 (N_1952,In_347,In_675);
and U1953 (N_1953,In_621,In_874);
and U1954 (N_1954,In_574,In_205);
xnor U1955 (N_1955,In_54,In_562);
nor U1956 (N_1956,In_356,In_366);
nand U1957 (N_1957,In_16,In_896);
nand U1958 (N_1958,In_582,In_236);
nand U1959 (N_1959,In_160,In_666);
nand U1960 (N_1960,In_396,In_61);
xor U1961 (N_1961,In_100,In_762);
nand U1962 (N_1962,In_655,In_82);
xor U1963 (N_1963,In_435,In_449);
nor U1964 (N_1964,In_151,In_314);
xor U1965 (N_1965,In_31,In_333);
xnor U1966 (N_1966,In_457,In_139);
and U1967 (N_1967,In_116,In_208);
or U1968 (N_1968,In_949,In_205);
and U1969 (N_1969,In_162,In_378);
xor U1970 (N_1970,In_640,In_811);
nand U1971 (N_1971,In_488,In_60);
or U1972 (N_1972,In_41,In_150);
nand U1973 (N_1973,In_463,In_207);
nor U1974 (N_1974,In_531,In_578);
or U1975 (N_1975,In_849,In_426);
nand U1976 (N_1976,In_185,In_273);
nor U1977 (N_1977,In_458,In_126);
nand U1978 (N_1978,In_204,In_523);
xor U1979 (N_1979,In_552,In_38);
nand U1980 (N_1980,In_457,In_268);
xor U1981 (N_1981,In_696,In_710);
or U1982 (N_1982,In_440,In_798);
nor U1983 (N_1983,In_206,In_290);
nand U1984 (N_1984,In_536,In_443);
nand U1985 (N_1985,In_524,In_657);
and U1986 (N_1986,In_687,In_622);
nand U1987 (N_1987,In_469,In_135);
xor U1988 (N_1988,In_609,In_453);
nor U1989 (N_1989,In_681,In_120);
nand U1990 (N_1990,In_820,In_671);
nand U1991 (N_1991,In_204,In_944);
or U1992 (N_1992,In_983,In_397);
and U1993 (N_1993,In_160,In_390);
xnor U1994 (N_1994,In_279,In_451);
nor U1995 (N_1995,In_617,In_691);
xnor U1996 (N_1996,In_398,In_566);
and U1997 (N_1997,In_516,In_107);
and U1998 (N_1998,In_281,In_470);
and U1999 (N_1999,In_31,In_82);
nor U2000 (N_2000,In_112,In_62);
nand U2001 (N_2001,In_627,In_590);
and U2002 (N_2002,In_734,In_881);
nor U2003 (N_2003,In_256,In_637);
nor U2004 (N_2004,In_209,In_307);
and U2005 (N_2005,In_599,In_369);
nand U2006 (N_2006,In_79,In_290);
and U2007 (N_2007,In_213,In_68);
or U2008 (N_2008,In_388,In_223);
nand U2009 (N_2009,In_517,In_425);
nor U2010 (N_2010,In_495,In_989);
nand U2011 (N_2011,In_17,In_259);
nand U2012 (N_2012,In_198,In_847);
nand U2013 (N_2013,In_884,In_933);
or U2014 (N_2014,In_813,In_705);
or U2015 (N_2015,In_698,In_294);
or U2016 (N_2016,In_774,In_280);
nor U2017 (N_2017,In_372,In_816);
or U2018 (N_2018,In_467,In_116);
or U2019 (N_2019,In_891,In_190);
and U2020 (N_2020,In_72,In_99);
or U2021 (N_2021,In_971,In_514);
or U2022 (N_2022,In_12,In_596);
and U2023 (N_2023,In_139,In_322);
nand U2024 (N_2024,In_905,In_573);
nand U2025 (N_2025,In_2,In_738);
and U2026 (N_2026,In_447,In_449);
nand U2027 (N_2027,In_244,In_567);
and U2028 (N_2028,In_339,In_486);
or U2029 (N_2029,In_797,In_700);
and U2030 (N_2030,In_500,In_438);
or U2031 (N_2031,In_678,In_600);
nor U2032 (N_2032,In_651,In_619);
or U2033 (N_2033,In_614,In_997);
nor U2034 (N_2034,In_392,In_224);
or U2035 (N_2035,In_609,In_683);
nand U2036 (N_2036,In_956,In_296);
and U2037 (N_2037,In_414,In_849);
xor U2038 (N_2038,In_196,In_187);
nor U2039 (N_2039,In_521,In_732);
or U2040 (N_2040,In_779,In_349);
and U2041 (N_2041,In_15,In_217);
or U2042 (N_2042,In_448,In_103);
or U2043 (N_2043,In_712,In_414);
and U2044 (N_2044,In_617,In_34);
xor U2045 (N_2045,In_93,In_679);
nand U2046 (N_2046,In_175,In_132);
or U2047 (N_2047,In_617,In_442);
nand U2048 (N_2048,In_874,In_555);
and U2049 (N_2049,In_768,In_431);
nand U2050 (N_2050,In_971,In_506);
or U2051 (N_2051,In_821,In_997);
nor U2052 (N_2052,In_107,In_248);
nand U2053 (N_2053,In_819,In_684);
or U2054 (N_2054,In_201,In_521);
nor U2055 (N_2055,In_503,In_679);
nor U2056 (N_2056,In_565,In_918);
or U2057 (N_2057,In_836,In_400);
or U2058 (N_2058,In_827,In_4);
xor U2059 (N_2059,In_747,In_731);
nand U2060 (N_2060,In_158,In_8);
or U2061 (N_2061,In_314,In_476);
nor U2062 (N_2062,In_603,In_598);
nor U2063 (N_2063,In_501,In_370);
nand U2064 (N_2064,In_535,In_65);
or U2065 (N_2065,In_110,In_937);
nand U2066 (N_2066,In_696,In_240);
nor U2067 (N_2067,In_440,In_212);
nor U2068 (N_2068,In_384,In_758);
nor U2069 (N_2069,In_211,In_328);
nor U2070 (N_2070,In_931,In_742);
nor U2071 (N_2071,In_789,In_923);
nand U2072 (N_2072,In_835,In_893);
nand U2073 (N_2073,In_732,In_773);
and U2074 (N_2074,In_946,In_650);
or U2075 (N_2075,In_345,In_844);
nor U2076 (N_2076,In_794,In_497);
nand U2077 (N_2077,In_544,In_728);
nor U2078 (N_2078,In_392,In_912);
and U2079 (N_2079,In_676,In_608);
nor U2080 (N_2080,In_276,In_135);
nor U2081 (N_2081,In_921,In_487);
or U2082 (N_2082,In_356,In_699);
or U2083 (N_2083,In_443,In_267);
and U2084 (N_2084,In_501,In_280);
nor U2085 (N_2085,In_340,In_207);
or U2086 (N_2086,In_540,In_416);
nand U2087 (N_2087,In_515,In_628);
nor U2088 (N_2088,In_757,In_487);
nand U2089 (N_2089,In_343,In_491);
or U2090 (N_2090,In_126,In_481);
nor U2091 (N_2091,In_778,In_972);
or U2092 (N_2092,In_24,In_437);
or U2093 (N_2093,In_953,In_375);
nor U2094 (N_2094,In_999,In_194);
or U2095 (N_2095,In_139,In_683);
nand U2096 (N_2096,In_218,In_281);
xor U2097 (N_2097,In_664,In_973);
xnor U2098 (N_2098,In_354,In_299);
nor U2099 (N_2099,In_641,In_22);
nor U2100 (N_2100,In_390,In_852);
and U2101 (N_2101,In_876,In_601);
xor U2102 (N_2102,In_187,In_732);
or U2103 (N_2103,In_415,In_808);
nand U2104 (N_2104,In_350,In_599);
nor U2105 (N_2105,In_685,In_590);
nor U2106 (N_2106,In_809,In_277);
nand U2107 (N_2107,In_997,In_272);
nand U2108 (N_2108,In_931,In_282);
nand U2109 (N_2109,In_751,In_566);
nand U2110 (N_2110,In_165,In_898);
nor U2111 (N_2111,In_838,In_730);
nor U2112 (N_2112,In_163,In_772);
or U2113 (N_2113,In_353,In_917);
xor U2114 (N_2114,In_525,In_608);
nor U2115 (N_2115,In_995,In_318);
nand U2116 (N_2116,In_127,In_953);
xor U2117 (N_2117,In_388,In_759);
nand U2118 (N_2118,In_279,In_359);
nand U2119 (N_2119,In_689,In_210);
and U2120 (N_2120,In_130,In_55);
nor U2121 (N_2121,In_325,In_626);
nand U2122 (N_2122,In_259,In_582);
and U2123 (N_2123,In_169,In_446);
nand U2124 (N_2124,In_434,In_903);
nand U2125 (N_2125,In_929,In_820);
nor U2126 (N_2126,In_843,In_142);
and U2127 (N_2127,In_207,In_534);
xnor U2128 (N_2128,In_788,In_274);
and U2129 (N_2129,In_507,In_248);
and U2130 (N_2130,In_251,In_209);
nor U2131 (N_2131,In_465,In_155);
xnor U2132 (N_2132,In_809,In_285);
nor U2133 (N_2133,In_339,In_607);
or U2134 (N_2134,In_616,In_30);
xnor U2135 (N_2135,In_184,In_279);
nand U2136 (N_2136,In_34,In_290);
nand U2137 (N_2137,In_630,In_249);
nand U2138 (N_2138,In_505,In_871);
or U2139 (N_2139,In_466,In_253);
nor U2140 (N_2140,In_953,In_92);
nand U2141 (N_2141,In_200,In_211);
and U2142 (N_2142,In_601,In_97);
or U2143 (N_2143,In_824,In_661);
nand U2144 (N_2144,In_258,In_809);
or U2145 (N_2145,In_68,In_786);
nand U2146 (N_2146,In_753,In_558);
nor U2147 (N_2147,In_499,In_518);
nand U2148 (N_2148,In_103,In_126);
nor U2149 (N_2149,In_63,In_232);
and U2150 (N_2150,In_502,In_161);
nand U2151 (N_2151,In_556,In_638);
or U2152 (N_2152,In_269,In_324);
and U2153 (N_2153,In_84,In_511);
nor U2154 (N_2154,In_133,In_546);
nand U2155 (N_2155,In_818,In_291);
or U2156 (N_2156,In_88,In_171);
nor U2157 (N_2157,In_956,In_193);
and U2158 (N_2158,In_21,In_453);
and U2159 (N_2159,In_694,In_827);
nor U2160 (N_2160,In_55,In_788);
nand U2161 (N_2161,In_470,In_981);
and U2162 (N_2162,In_627,In_198);
and U2163 (N_2163,In_141,In_778);
xnor U2164 (N_2164,In_531,In_887);
nand U2165 (N_2165,In_271,In_728);
nor U2166 (N_2166,In_373,In_678);
or U2167 (N_2167,In_79,In_695);
nand U2168 (N_2168,In_289,In_268);
nand U2169 (N_2169,In_387,In_606);
xnor U2170 (N_2170,In_913,In_215);
nor U2171 (N_2171,In_675,In_367);
nand U2172 (N_2172,In_785,In_884);
nand U2173 (N_2173,In_379,In_957);
nand U2174 (N_2174,In_103,In_226);
and U2175 (N_2175,In_400,In_795);
or U2176 (N_2176,In_598,In_664);
nor U2177 (N_2177,In_971,In_570);
or U2178 (N_2178,In_422,In_864);
or U2179 (N_2179,In_697,In_879);
and U2180 (N_2180,In_761,In_676);
and U2181 (N_2181,In_20,In_593);
or U2182 (N_2182,In_749,In_156);
nand U2183 (N_2183,In_658,In_345);
nand U2184 (N_2184,In_231,In_366);
nand U2185 (N_2185,In_379,In_863);
nand U2186 (N_2186,In_356,In_480);
or U2187 (N_2187,In_574,In_885);
xor U2188 (N_2188,In_119,In_453);
or U2189 (N_2189,In_451,In_447);
nand U2190 (N_2190,In_717,In_294);
and U2191 (N_2191,In_892,In_547);
and U2192 (N_2192,In_753,In_272);
xnor U2193 (N_2193,In_909,In_691);
xnor U2194 (N_2194,In_978,In_934);
or U2195 (N_2195,In_264,In_231);
nand U2196 (N_2196,In_164,In_706);
nand U2197 (N_2197,In_37,In_263);
nor U2198 (N_2198,In_655,In_319);
nand U2199 (N_2199,In_754,In_215);
or U2200 (N_2200,In_994,In_188);
nand U2201 (N_2201,In_249,In_570);
nor U2202 (N_2202,In_952,In_851);
or U2203 (N_2203,In_592,In_149);
nand U2204 (N_2204,In_225,In_624);
and U2205 (N_2205,In_176,In_448);
xnor U2206 (N_2206,In_186,In_344);
nand U2207 (N_2207,In_698,In_183);
nand U2208 (N_2208,In_180,In_284);
nand U2209 (N_2209,In_519,In_281);
nand U2210 (N_2210,In_557,In_909);
or U2211 (N_2211,In_101,In_549);
or U2212 (N_2212,In_915,In_526);
or U2213 (N_2213,In_304,In_489);
or U2214 (N_2214,In_478,In_593);
and U2215 (N_2215,In_533,In_70);
nand U2216 (N_2216,In_380,In_706);
nor U2217 (N_2217,In_701,In_492);
xnor U2218 (N_2218,In_730,In_773);
and U2219 (N_2219,In_733,In_537);
and U2220 (N_2220,In_168,In_145);
nand U2221 (N_2221,In_111,In_770);
nor U2222 (N_2222,In_182,In_191);
and U2223 (N_2223,In_926,In_341);
nand U2224 (N_2224,In_281,In_929);
or U2225 (N_2225,In_15,In_147);
nor U2226 (N_2226,In_74,In_321);
nand U2227 (N_2227,In_929,In_523);
or U2228 (N_2228,In_542,In_181);
or U2229 (N_2229,In_980,In_30);
or U2230 (N_2230,In_609,In_375);
or U2231 (N_2231,In_568,In_755);
and U2232 (N_2232,In_613,In_979);
and U2233 (N_2233,In_829,In_100);
and U2234 (N_2234,In_774,In_277);
xor U2235 (N_2235,In_47,In_781);
xor U2236 (N_2236,In_742,In_81);
nor U2237 (N_2237,In_740,In_546);
nand U2238 (N_2238,In_445,In_699);
and U2239 (N_2239,In_452,In_519);
or U2240 (N_2240,In_718,In_217);
nand U2241 (N_2241,In_994,In_778);
or U2242 (N_2242,In_199,In_353);
or U2243 (N_2243,In_118,In_31);
xor U2244 (N_2244,In_854,In_743);
and U2245 (N_2245,In_556,In_534);
or U2246 (N_2246,In_403,In_562);
or U2247 (N_2247,In_177,In_262);
xor U2248 (N_2248,In_678,In_540);
or U2249 (N_2249,In_970,In_93);
and U2250 (N_2250,In_104,In_684);
xnor U2251 (N_2251,In_715,In_702);
nor U2252 (N_2252,In_379,In_843);
nor U2253 (N_2253,In_161,In_885);
or U2254 (N_2254,In_508,In_49);
or U2255 (N_2255,In_582,In_470);
nor U2256 (N_2256,In_71,In_300);
and U2257 (N_2257,In_122,In_551);
nor U2258 (N_2258,In_634,In_877);
nand U2259 (N_2259,In_648,In_984);
nor U2260 (N_2260,In_724,In_347);
and U2261 (N_2261,In_879,In_944);
nand U2262 (N_2262,In_875,In_828);
nand U2263 (N_2263,In_113,In_528);
nand U2264 (N_2264,In_815,In_574);
nand U2265 (N_2265,In_207,In_164);
nor U2266 (N_2266,In_207,In_122);
nor U2267 (N_2267,In_796,In_217);
and U2268 (N_2268,In_706,In_282);
or U2269 (N_2269,In_481,In_586);
and U2270 (N_2270,In_569,In_803);
nand U2271 (N_2271,In_98,In_361);
and U2272 (N_2272,In_656,In_867);
nor U2273 (N_2273,In_159,In_157);
nand U2274 (N_2274,In_700,In_130);
xnor U2275 (N_2275,In_322,In_123);
xor U2276 (N_2276,In_318,In_0);
or U2277 (N_2277,In_768,In_709);
nor U2278 (N_2278,In_777,In_264);
nand U2279 (N_2279,In_6,In_859);
or U2280 (N_2280,In_856,In_232);
or U2281 (N_2281,In_395,In_542);
and U2282 (N_2282,In_964,In_672);
nor U2283 (N_2283,In_739,In_759);
nor U2284 (N_2284,In_388,In_939);
nor U2285 (N_2285,In_818,In_688);
nand U2286 (N_2286,In_75,In_868);
nand U2287 (N_2287,In_921,In_822);
or U2288 (N_2288,In_828,In_854);
and U2289 (N_2289,In_246,In_56);
nand U2290 (N_2290,In_952,In_783);
and U2291 (N_2291,In_800,In_857);
and U2292 (N_2292,In_291,In_735);
nor U2293 (N_2293,In_682,In_193);
or U2294 (N_2294,In_825,In_134);
nand U2295 (N_2295,In_937,In_768);
nand U2296 (N_2296,In_156,In_190);
nor U2297 (N_2297,In_551,In_284);
nor U2298 (N_2298,In_587,In_471);
xor U2299 (N_2299,In_186,In_755);
nor U2300 (N_2300,In_597,In_630);
and U2301 (N_2301,In_725,In_931);
nor U2302 (N_2302,In_593,In_843);
and U2303 (N_2303,In_84,In_845);
and U2304 (N_2304,In_750,In_643);
nor U2305 (N_2305,In_273,In_193);
or U2306 (N_2306,In_925,In_738);
and U2307 (N_2307,In_696,In_843);
xnor U2308 (N_2308,In_523,In_202);
nand U2309 (N_2309,In_81,In_703);
or U2310 (N_2310,In_640,In_718);
and U2311 (N_2311,In_248,In_920);
nor U2312 (N_2312,In_242,In_760);
xor U2313 (N_2313,In_100,In_858);
nor U2314 (N_2314,In_181,In_58);
xnor U2315 (N_2315,In_403,In_610);
or U2316 (N_2316,In_24,In_782);
nand U2317 (N_2317,In_285,In_27);
nor U2318 (N_2318,In_227,In_766);
and U2319 (N_2319,In_603,In_909);
nand U2320 (N_2320,In_438,In_381);
and U2321 (N_2321,In_768,In_76);
nor U2322 (N_2322,In_796,In_521);
or U2323 (N_2323,In_426,In_806);
nand U2324 (N_2324,In_605,In_701);
nand U2325 (N_2325,In_677,In_245);
and U2326 (N_2326,In_864,In_766);
nand U2327 (N_2327,In_524,In_45);
and U2328 (N_2328,In_850,In_996);
or U2329 (N_2329,In_538,In_571);
and U2330 (N_2330,In_726,In_600);
or U2331 (N_2331,In_556,In_551);
nand U2332 (N_2332,In_717,In_638);
nor U2333 (N_2333,In_185,In_569);
xor U2334 (N_2334,In_917,In_696);
xor U2335 (N_2335,In_844,In_409);
and U2336 (N_2336,In_181,In_66);
nand U2337 (N_2337,In_95,In_667);
or U2338 (N_2338,In_341,In_405);
nor U2339 (N_2339,In_780,In_830);
nor U2340 (N_2340,In_971,In_177);
and U2341 (N_2341,In_352,In_821);
nand U2342 (N_2342,In_160,In_491);
nor U2343 (N_2343,In_783,In_977);
and U2344 (N_2344,In_31,In_78);
and U2345 (N_2345,In_18,In_937);
or U2346 (N_2346,In_962,In_235);
and U2347 (N_2347,In_920,In_376);
or U2348 (N_2348,In_654,In_326);
nand U2349 (N_2349,In_449,In_173);
or U2350 (N_2350,In_893,In_187);
or U2351 (N_2351,In_174,In_97);
nor U2352 (N_2352,In_769,In_677);
nor U2353 (N_2353,In_256,In_300);
or U2354 (N_2354,In_808,In_526);
or U2355 (N_2355,In_675,In_681);
and U2356 (N_2356,In_685,In_771);
xor U2357 (N_2357,In_270,In_988);
nor U2358 (N_2358,In_46,In_159);
nand U2359 (N_2359,In_979,In_342);
nor U2360 (N_2360,In_1,In_967);
and U2361 (N_2361,In_463,In_794);
and U2362 (N_2362,In_730,In_335);
nand U2363 (N_2363,In_620,In_5);
nand U2364 (N_2364,In_496,In_580);
and U2365 (N_2365,In_310,In_172);
and U2366 (N_2366,In_283,In_934);
nand U2367 (N_2367,In_166,In_183);
nor U2368 (N_2368,In_680,In_0);
and U2369 (N_2369,In_701,In_859);
nor U2370 (N_2370,In_173,In_688);
and U2371 (N_2371,In_593,In_502);
nor U2372 (N_2372,In_463,In_948);
and U2373 (N_2373,In_636,In_910);
or U2374 (N_2374,In_338,In_4);
nor U2375 (N_2375,In_930,In_15);
or U2376 (N_2376,In_13,In_919);
and U2377 (N_2377,In_171,In_528);
or U2378 (N_2378,In_101,In_829);
nor U2379 (N_2379,In_630,In_272);
and U2380 (N_2380,In_847,In_320);
and U2381 (N_2381,In_824,In_290);
nand U2382 (N_2382,In_460,In_674);
nor U2383 (N_2383,In_0,In_763);
or U2384 (N_2384,In_442,In_3);
or U2385 (N_2385,In_372,In_6);
nand U2386 (N_2386,In_206,In_181);
and U2387 (N_2387,In_646,In_838);
and U2388 (N_2388,In_308,In_526);
or U2389 (N_2389,In_462,In_6);
and U2390 (N_2390,In_15,In_880);
nand U2391 (N_2391,In_391,In_463);
nand U2392 (N_2392,In_768,In_964);
and U2393 (N_2393,In_72,In_926);
nor U2394 (N_2394,In_266,In_258);
nor U2395 (N_2395,In_383,In_698);
or U2396 (N_2396,In_700,In_976);
and U2397 (N_2397,In_107,In_378);
nand U2398 (N_2398,In_981,In_352);
and U2399 (N_2399,In_571,In_175);
nor U2400 (N_2400,In_989,In_82);
nand U2401 (N_2401,In_122,In_429);
and U2402 (N_2402,In_671,In_953);
nand U2403 (N_2403,In_711,In_553);
and U2404 (N_2404,In_648,In_908);
or U2405 (N_2405,In_168,In_965);
nor U2406 (N_2406,In_108,In_624);
and U2407 (N_2407,In_257,In_740);
nor U2408 (N_2408,In_485,In_940);
or U2409 (N_2409,In_968,In_536);
xnor U2410 (N_2410,In_485,In_83);
nand U2411 (N_2411,In_288,In_242);
nand U2412 (N_2412,In_337,In_325);
nor U2413 (N_2413,In_58,In_127);
and U2414 (N_2414,In_490,In_672);
xnor U2415 (N_2415,In_515,In_970);
and U2416 (N_2416,In_513,In_538);
xnor U2417 (N_2417,In_743,In_1);
or U2418 (N_2418,In_917,In_507);
nand U2419 (N_2419,In_139,In_537);
nand U2420 (N_2420,In_818,In_640);
xnor U2421 (N_2421,In_208,In_509);
xnor U2422 (N_2422,In_51,In_976);
nand U2423 (N_2423,In_285,In_317);
xor U2424 (N_2424,In_908,In_92);
nand U2425 (N_2425,In_17,In_218);
nand U2426 (N_2426,In_160,In_14);
nor U2427 (N_2427,In_133,In_659);
or U2428 (N_2428,In_229,In_960);
nor U2429 (N_2429,In_772,In_955);
or U2430 (N_2430,In_215,In_59);
or U2431 (N_2431,In_123,In_138);
and U2432 (N_2432,In_682,In_199);
nand U2433 (N_2433,In_423,In_917);
and U2434 (N_2434,In_664,In_799);
and U2435 (N_2435,In_905,In_542);
or U2436 (N_2436,In_919,In_32);
nor U2437 (N_2437,In_281,In_531);
or U2438 (N_2438,In_707,In_581);
nand U2439 (N_2439,In_163,In_612);
nor U2440 (N_2440,In_758,In_69);
nor U2441 (N_2441,In_26,In_989);
and U2442 (N_2442,In_475,In_396);
nand U2443 (N_2443,In_163,In_704);
nand U2444 (N_2444,In_831,In_586);
and U2445 (N_2445,In_500,In_393);
or U2446 (N_2446,In_754,In_668);
or U2447 (N_2447,In_494,In_798);
nand U2448 (N_2448,In_154,In_255);
and U2449 (N_2449,In_438,In_191);
nand U2450 (N_2450,In_716,In_700);
nand U2451 (N_2451,In_802,In_682);
nor U2452 (N_2452,In_161,In_904);
and U2453 (N_2453,In_854,In_26);
nand U2454 (N_2454,In_430,In_755);
or U2455 (N_2455,In_5,In_726);
nand U2456 (N_2456,In_106,In_76);
and U2457 (N_2457,In_912,In_924);
and U2458 (N_2458,In_190,In_881);
or U2459 (N_2459,In_36,In_769);
or U2460 (N_2460,In_307,In_139);
nor U2461 (N_2461,In_186,In_61);
nand U2462 (N_2462,In_404,In_568);
or U2463 (N_2463,In_543,In_710);
nand U2464 (N_2464,In_964,In_532);
and U2465 (N_2465,In_132,In_49);
or U2466 (N_2466,In_480,In_849);
nor U2467 (N_2467,In_920,In_84);
and U2468 (N_2468,In_379,In_425);
or U2469 (N_2469,In_945,In_320);
xnor U2470 (N_2470,In_229,In_313);
and U2471 (N_2471,In_737,In_67);
nand U2472 (N_2472,In_138,In_41);
and U2473 (N_2473,In_336,In_254);
nand U2474 (N_2474,In_850,In_491);
nand U2475 (N_2475,In_672,In_926);
or U2476 (N_2476,In_67,In_292);
or U2477 (N_2477,In_996,In_144);
and U2478 (N_2478,In_577,In_590);
and U2479 (N_2479,In_22,In_454);
nor U2480 (N_2480,In_157,In_547);
or U2481 (N_2481,In_218,In_302);
and U2482 (N_2482,In_943,In_789);
and U2483 (N_2483,In_95,In_680);
nand U2484 (N_2484,In_460,In_504);
or U2485 (N_2485,In_367,In_973);
nand U2486 (N_2486,In_246,In_629);
or U2487 (N_2487,In_688,In_41);
nor U2488 (N_2488,In_222,In_854);
nand U2489 (N_2489,In_728,In_962);
or U2490 (N_2490,In_409,In_830);
nand U2491 (N_2491,In_155,In_342);
and U2492 (N_2492,In_114,In_588);
or U2493 (N_2493,In_171,In_871);
or U2494 (N_2494,In_714,In_872);
and U2495 (N_2495,In_766,In_553);
nor U2496 (N_2496,In_151,In_581);
nand U2497 (N_2497,In_476,In_31);
or U2498 (N_2498,In_738,In_537);
nor U2499 (N_2499,In_994,In_380);
nand U2500 (N_2500,In_701,In_49);
and U2501 (N_2501,In_712,In_466);
and U2502 (N_2502,In_658,In_352);
or U2503 (N_2503,In_166,In_710);
xnor U2504 (N_2504,In_568,In_573);
or U2505 (N_2505,In_556,In_236);
nor U2506 (N_2506,In_107,In_430);
and U2507 (N_2507,In_693,In_177);
and U2508 (N_2508,In_23,In_975);
or U2509 (N_2509,In_442,In_878);
or U2510 (N_2510,In_409,In_936);
nand U2511 (N_2511,In_756,In_796);
or U2512 (N_2512,In_17,In_235);
or U2513 (N_2513,In_644,In_734);
and U2514 (N_2514,In_246,In_678);
nand U2515 (N_2515,In_819,In_554);
and U2516 (N_2516,In_756,In_986);
xor U2517 (N_2517,In_695,In_665);
and U2518 (N_2518,In_807,In_706);
xnor U2519 (N_2519,In_288,In_895);
nor U2520 (N_2520,In_518,In_910);
xnor U2521 (N_2521,In_480,In_685);
nand U2522 (N_2522,In_336,In_979);
nand U2523 (N_2523,In_579,In_938);
and U2524 (N_2524,In_290,In_800);
nand U2525 (N_2525,In_845,In_567);
xor U2526 (N_2526,In_187,In_539);
nor U2527 (N_2527,In_587,In_28);
nor U2528 (N_2528,In_281,In_142);
or U2529 (N_2529,In_98,In_124);
and U2530 (N_2530,In_65,In_178);
and U2531 (N_2531,In_458,In_211);
or U2532 (N_2532,In_186,In_339);
and U2533 (N_2533,In_108,In_610);
and U2534 (N_2534,In_823,In_255);
nor U2535 (N_2535,In_277,In_139);
and U2536 (N_2536,In_340,In_981);
xnor U2537 (N_2537,In_981,In_155);
and U2538 (N_2538,In_565,In_479);
and U2539 (N_2539,In_773,In_203);
nand U2540 (N_2540,In_833,In_402);
nor U2541 (N_2541,In_332,In_104);
or U2542 (N_2542,In_954,In_108);
or U2543 (N_2543,In_564,In_826);
or U2544 (N_2544,In_402,In_434);
xor U2545 (N_2545,In_154,In_779);
xor U2546 (N_2546,In_272,In_685);
nand U2547 (N_2547,In_116,In_262);
and U2548 (N_2548,In_78,In_982);
nand U2549 (N_2549,In_229,In_866);
nand U2550 (N_2550,In_199,In_639);
or U2551 (N_2551,In_90,In_791);
or U2552 (N_2552,In_434,In_520);
nor U2553 (N_2553,In_569,In_525);
nor U2554 (N_2554,In_897,In_809);
or U2555 (N_2555,In_55,In_992);
or U2556 (N_2556,In_992,In_891);
and U2557 (N_2557,In_919,In_378);
or U2558 (N_2558,In_684,In_814);
and U2559 (N_2559,In_737,In_125);
and U2560 (N_2560,In_70,In_839);
nor U2561 (N_2561,In_355,In_863);
nor U2562 (N_2562,In_781,In_811);
nor U2563 (N_2563,In_390,In_176);
nand U2564 (N_2564,In_80,In_917);
nor U2565 (N_2565,In_143,In_356);
or U2566 (N_2566,In_735,In_57);
xnor U2567 (N_2567,In_440,In_49);
nor U2568 (N_2568,In_293,In_333);
nand U2569 (N_2569,In_178,In_445);
nor U2570 (N_2570,In_971,In_716);
and U2571 (N_2571,In_792,In_904);
or U2572 (N_2572,In_317,In_620);
and U2573 (N_2573,In_342,In_385);
nor U2574 (N_2574,In_39,In_40);
or U2575 (N_2575,In_420,In_188);
or U2576 (N_2576,In_895,In_849);
xor U2577 (N_2577,In_171,In_569);
nor U2578 (N_2578,In_119,In_376);
or U2579 (N_2579,In_115,In_277);
xnor U2580 (N_2580,In_184,In_251);
and U2581 (N_2581,In_208,In_286);
or U2582 (N_2582,In_445,In_48);
nand U2583 (N_2583,In_977,In_803);
and U2584 (N_2584,In_894,In_743);
or U2585 (N_2585,In_777,In_193);
nand U2586 (N_2586,In_110,In_306);
xnor U2587 (N_2587,In_394,In_380);
and U2588 (N_2588,In_673,In_677);
nand U2589 (N_2589,In_219,In_404);
nand U2590 (N_2590,In_344,In_779);
or U2591 (N_2591,In_188,In_594);
nor U2592 (N_2592,In_456,In_745);
nor U2593 (N_2593,In_575,In_323);
nand U2594 (N_2594,In_450,In_621);
xor U2595 (N_2595,In_966,In_184);
and U2596 (N_2596,In_824,In_899);
or U2597 (N_2597,In_5,In_250);
and U2598 (N_2598,In_888,In_659);
nor U2599 (N_2599,In_647,In_904);
nor U2600 (N_2600,In_180,In_512);
xor U2601 (N_2601,In_349,In_112);
nand U2602 (N_2602,In_321,In_758);
nand U2603 (N_2603,In_410,In_838);
or U2604 (N_2604,In_739,In_546);
nand U2605 (N_2605,In_493,In_846);
nand U2606 (N_2606,In_641,In_363);
and U2607 (N_2607,In_178,In_707);
xor U2608 (N_2608,In_912,In_259);
nand U2609 (N_2609,In_65,In_508);
xnor U2610 (N_2610,In_471,In_314);
and U2611 (N_2611,In_492,In_190);
xor U2612 (N_2612,In_690,In_802);
nor U2613 (N_2613,In_826,In_129);
xor U2614 (N_2614,In_425,In_856);
nand U2615 (N_2615,In_589,In_222);
xnor U2616 (N_2616,In_461,In_21);
or U2617 (N_2617,In_312,In_544);
nand U2618 (N_2618,In_537,In_944);
nor U2619 (N_2619,In_431,In_735);
or U2620 (N_2620,In_816,In_231);
nor U2621 (N_2621,In_273,In_652);
nand U2622 (N_2622,In_576,In_607);
or U2623 (N_2623,In_761,In_35);
and U2624 (N_2624,In_218,In_182);
nor U2625 (N_2625,In_12,In_444);
and U2626 (N_2626,In_519,In_526);
or U2627 (N_2627,In_449,In_704);
nor U2628 (N_2628,In_846,In_368);
or U2629 (N_2629,In_169,In_943);
or U2630 (N_2630,In_677,In_33);
and U2631 (N_2631,In_410,In_861);
and U2632 (N_2632,In_770,In_564);
nor U2633 (N_2633,In_759,In_988);
xor U2634 (N_2634,In_393,In_442);
nand U2635 (N_2635,In_722,In_377);
or U2636 (N_2636,In_337,In_219);
or U2637 (N_2637,In_994,In_661);
or U2638 (N_2638,In_204,In_71);
nand U2639 (N_2639,In_53,In_182);
nand U2640 (N_2640,In_874,In_970);
or U2641 (N_2641,In_822,In_671);
and U2642 (N_2642,In_293,In_753);
nand U2643 (N_2643,In_202,In_98);
nand U2644 (N_2644,In_466,In_179);
nor U2645 (N_2645,In_9,In_152);
nor U2646 (N_2646,In_136,In_693);
nor U2647 (N_2647,In_221,In_179);
and U2648 (N_2648,In_988,In_607);
and U2649 (N_2649,In_886,In_902);
nor U2650 (N_2650,In_67,In_137);
and U2651 (N_2651,In_390,In_356);
nor U2652 (N_2652,In_822,In_372);
nor U2653 (N_2653,In_429,In_576);
and U2654 (N_2654,In_76,In_404);
or U2655 (N_2655,In_501,In_596);
nand U2656 (N_2656,In_365,In_469);
and U2657 (N_2657,In_492,In_990);
nor U2658 (N_2658,In_584,In_127);
nand U2659 (N_2659,In_883,In_52);
nor U2660 (N_2660,In_272,In_566);
nand U2661 (N_2661,In_576,In_679);
and U2662 (N_2662,In_704,In_295);
nand U2663 (N_2663,In_138,In_31);
nor U2664 (N_2664,In_115,In_339);
and U2665 (N_2665,In_314,In_609);
nand U2666 (N_2666,In_143,In_67);
nor U2667 (N_2667,In_836,In_510);
or U2668 (N_2668,In_524,In_281);
nor U2669 (N_2669,In_357,In_476);
or U2670 (N_2670,In_864,In_889);
nor U2671 (N_2671,In_242,In_60);
nand U2672 (N_2672,In_271,In_612);
and U2673 (N_2673,In_238,In_549);
and U2674 (N_2674,In_112,In_433);
nor U2675 (N_2675,In_475,In_37);
nand U2676 (N_2676,In_79,In_882);
nand U2677 (N_2677,In_779,In_642);
or U2678 (N_2678,In_673,In_898);
and U2679 (N_2679,In_59,In_610);
nand U2680 (N_2680,In_248,In_538);
or U2681 (N_2681,In_69,In_351);
nand U2682 (N_2682,In_541,In_57);
nand U2683 (N_2683,In_825,In_908);
nand U2684 (N_2684,In_117,In_119);
or U2685 (N_2685,In_502,In_343);
or U2686 (N_2686,In_795,In_971);
and U2687 (N_2687,In_909,In_499);
or U2688 (N_2688,In_665,In_9);
nor U2689 (N_2689,In_664,In_116);
and U2690 (N_2690,In_534,In_172);
and U2691 (N_2691,In_889,In_167);
and U2692 (N_2692,In_77,In_22);
nor U2693 (N_2693,In_549,In_858);
nor U2694 (N_2694,In_990,In_428);
and U2695 (N_2695,In_762,In_800);
or U2696 (N_2696,In_771,In_578);
or U2697 (N_2697,In_759,In_154);
nor U2698 (N_2698,In_893,In_816);
and U2699 (N_2699,In_742,In_581);
nand U2700 (N_2700,In_450,In_179);
xnor U2701 (N_2701,In_140,In_826);
and U2702 (N_2702,In_507,In_933);
or U2703 (N_2703,In_445,In_571);
and U2704 (N_2704,In_923,In_735);
nor U2705 (N_2705,In_186,In_161);
or U2706 (N_2706,In_827,In_534);
or U2707 (N_2707,In_364,In_52);
nor U2708 (N_2708,In_688,In_249);
and U2709 (N_2709,In_83,In_662);
nor U2710 (N_2710,In_563,In_87);
and U2711 (N_2711,In_908,In_594);
or U2712 (N_2712,In_267,In_174);
and U2713 (N_2713,In_442,In_555);
nor U2714 (N_2714,In_680,In_973);
nand U2715 (N_2715,In_283,In_895);
nand U2716 (N_2716,In_822,In_306);
nor U2717 (N_2717,In_983,In_926);
or U2718 (N_2718,In_229,In_514);
or U2719 (N_2719,In_734,In_739);
nand U2720 (N_2720,In_220,In_135);
or U2721 (N_2721,In_377,In_830);
nor U2722 (N_2722,In_22,In_105);
or U2723 (N_2723,In_554,In_300);
and U2724 (N_2724,In_451,In_28);
nand U2725 (N_2725,In_410,In_279);
nand U2726 (N_2726,In_705,In_787);
and U2727 (N_2727,In_469,In_218);
nor U2728 (N_2728,In_912,In_759);
or U2729 (N_2729,In_444,In_165);
nand U2730 (N_2730,In_10,In_437);
or U2731 (N_2731,In_418,In_562);
and U2732 (N_2732,In_264,In_9);
or U2733 (N_2733,In_245,In_633);
and U2734 (N_2734,In_24,In_411);
nor U2735 (N_2735,In_641,In_913);
nand U2736 (N_2736,In_602,In_200);
nand U2737 (N_2737,In_846,In_441);
nor U2738 (N_2738,In_851,In_459);
xor U2739 (N_2739,In_159,In_113);
and U2740 (N_2740,In_697,In_506);
and U2741 (N_2741,In_931,In_138);
nand U2742 (N_2742,In_697,In_488);
xor U2743 (N_2743,In_365,In_786);
nor U2744 (N_2744,In_965,In_868);
and U2745 (N_2745,In_895,In_906);
or U2746 (N_2746,In_657,In_639);
nor U2747 (N_2747,In_403,In_762);
nand U2748 (N_2748,In_224,In_100);
and U2749 (N_2749,In_170,In_69);
nand U2750 (N_2750,In_398,In_410);
nand U2751 (N_2751,In_6,In_547);
or U2752 (N_2752,In_730,In_122);
nor U2753 (N_2753,In_850,In_767);
and U2754 (N_2754,In_518,In_996);
nand U2755 (N_2755,In_183,In_930);
nor U2756 (N_2756,In_152,In_893);
and U2757 (N_2757,In_340,In_675);
or U2758 (N_2758,In_1,In_261);
or U2759 (N_2759,In_612,In_238);
or U2760 (N_2760,In_224,In_608);
or U2761 (N_2761,In_127,In_951);
nand U2762 (N_2762,In_285,In_562);
xor U2763 (N_2763,In_51,In_751);
xnor U2764 (N_2764,In_540,In_156);
and U2765 (N_2765,In_849,In_850);
or U2766 (N_2766,In_661,In_210);
nor U2767 (N_2767,In_942,In_612);
nor U2768 (N_2768,In_177,In_536);
nor U2769 (N_2769,In_424,In_706);
and U2770 (N_2770,In_612,In_941);
nand U2771 (N_2771,In_803,In_709);
nand U2772 (N_2772,In_382,In_179);
nand U2773 (N_2773,In_57,In_161);
and U2774 (N_2774,In_371,In_527);
and U2775 (N_2775,In_345,In_643);
nand U2776 (N_2776,In_423,In_551);
nand U2777 (N_2777,In_639,In_125);
and U2778 (N_2778,In_898,In_111);
or U2779 (N_2779,In_953,In_927);
nor U2780 (N_2780,In_545,In_301);
or U2781 (N_2781,In_266,In_651);
nor U2782 (N_2782,In_320,In_914);
or U2783 (N_2783,In_78,In_828);
nand U2784 (N_2784,In_740,In_942);
and U2785 (N_2785,In_205,In_170);
or U2786 (N_2786,In_510,In_944);
nand U2787 (N_2787,In_38,In_690);
xor U2788 (N_2788,In_556,In_172);
and U2789 (N_2789,In_955,In_568);
nand U2790 (N_2790,In_166,In_464);
nand U2791 (N_2791,In_443,In_95);
nand U2792 (N_2792,In_261,In_657);
nand U2793 (N_2793,In_514,In_529);
or U2794 (N_2794,In_96,In_659);
or U2795 (N_2795,In_323,In_689);
or U2796 (N_2796,In_163,In_156);
or U2797 (N_2797,In_266,In_81);
xor U2798 (N_2798,In_973,In_815);
nand U2799 (N_2799,In_103,In_601);
xnor U2800 (N_2800,In_727,In_456);
or U2801 (N_2801,In_782,In_470);
and U2802 (N_2802,In_827,In_92);
nor U2803 (N_2803,In_269,In_31);
or U2804 (N_2804,In_533,In_699);
and U2805 (N_2805,In_917,In_737);
xnor U2806 (N_2806,In_28,In_464);
nor U2807 (N_2807,In_560,In_559);
nand U2808 (N_2808,In_519,In_35);
or U2809 (N_2809,In_62,In_358);
or U2810 (N_2810,In_278,In_490);
and U2811 (N_2811,In_659,In_501);
nand U2812 (N_2812,In_914,In_416);
nor U2813 (N_2813,In_521,In_944);
nor U2814 (N_2814,In_936,In_741);
or U2815 (N_2815,In_582,In_52);
nand U2816 (N_2816,In_158,In_313);
or U2817 (N_2817,In_946,In_318);
and U2818 (N_2818,In_388,In_859);
and U2819 (N_2819,In_975,In_619);
or U2820 (N_2820,In_312,In_140);
and U2821 (N_2821,In_165,In_917);
nand U2822 (N_2822,In_129,In_720);
nor U2823 (N_2823,In_28,In_348);
nand U2824 (N_2824,In_663,In_555);
nand U2825 (N_2825,In_570,In_801);
and U2826 (N_2826,In_648,In_132);
and U2827 (N_2827,In_458,In_681);
nor U2828 (N_2828,In_999,In_953);
and U2829 (N_2829,In_212,In_239);
and U2830 (N_2830,In_841,In_236);
nor U2831 (N_2831,In_372,In_423);
and U2832 (N_2832,In_162,In_969);
nor U2833 (N_2833,In_477,In_449);
nor U2834 (N_2834,In_591,In_23);
xor U2835 (N_2835,In_854,In_241);
and U2836 (N_2836,In_247,In_421);
xnor U2837 (N_2837,In_853,In_721);
and U2838 (N_2838,In_836,In_829);
and U2839 (N_2839,In_744,In_317);
nor U2840 (N_2840,In_708,In_372);
xnor U2841 (N_2841,In_703,In_248);
and U2842 (N_2842,In_362,In_961);
xnor U2843 (N_2843,In_745,In_639);
nand U2844 (N_2844,In_413,In_403);
xnor U2845 (N_2845,In_201,In_888);
or U2846 (N_2846,In_643,In_114);
or U2847 (N_2847,In_915,In_769);
or U2848 (N_2848,In_824,In_737);
nand U2849 (N_2849,In_419,In_177);
and U2850 (N_2850,In_542,In_58);
or U2851 (N_2851,In_984,In_651);
xor U2852 (N_2852,In_409,In_832);
or U2853 (N_2853,In_13,In_391);
and U2854 (N_2854,In_657,In_222);
or U2855 (N_2855,In_437,In_322);
nor U2856 (N_2856,In_432,In_310);
or U2857 (N_2857,In_110,In_279);
or U2858 (N_2858,In_70,In_614);
nor U2859 (N_2859,In_668,In_593);
and U2860 (N_2860,In_951,In_958);
nor U2861 (N_2861,In_196,In_647);
and U2862 (N_2862,In_917,In_896);
nor U2863 (N_2863,In_177,In_106);
nor U2864 (N_2864,In_313,In_430);
and U2865 (N_2865,In_497,In_473);
or U2866 (N_2866,In_366,In_991);
nor U2867 (N_2867,In_428,In_761);
or U2868 (N_2868,In_302,In_821);
nand U2869 (N_2869,In_761,In_816);
and U2870 (N_2870,In_158,In_931);
xor U2871 (N_2871,In_85,In_928);
nand U2872 (N_2872,In_613,In_417);
nand U2873 (N_2873,In_312,In_44);
nand U2874 (N_2874,In_787,In_452);
xor U2875 (N_2875,In_272,In_798);
and U2876 (N_2876,In_434,In_720);
and U2877 (N_2877,In_842,In_957);
nand U2878 (N_2878,In_347,In_194);
and U2879 (N_2879,In_813,In_433);
nand U2880 (N_2880,In_55,In_267);
or U2881 (N_2881,In_86,In_146);
or U2882 (N_2882,In_672,In_552);
and U2883 (N_2883,In_284,In_711);
or U2884 (N_2884,In_513,In_16);
and U2885 (N_2885,In_812,In_117);
and U2886 (N_2886,In_323,In_208);
and U2887 (N_2887,In_532,In_160);
and U2888 (N_2888,In_83,In_341);
nor U2889 (N_2889,In_366,In_823);
and U2890 (N_2890,In_387,In_741);
and U2891 (N_2891,In_941,In_316);
nor U2892 (N_2892,In_10,In_664);
nand U2893 (N_2893,In_832,In_646);
and U2894 (N_2894,In_371,In_529);
and U2895 (N_2895,In_734,In_797);
nand U2896 (N_2896,In_478,In_678);
nand U2897 (N_2897,In_372,In_645);
and U2898 (N_2898,In_564,In_746);
nand U2899 (N_2899,In_101,In_180);
or U2900 (N_2900,In_86,In_693);
or U2901 (N_2901,In_161,In_975);
nand U2902 (N_2902,In_302,In_533);
or U2903 (N_2903,In_727,In_324);
and U2904 (N_2904,In_670,In_246);
and U2905 (N_2905,In_280,In_881);
or U2906 (N_2906,In_309,In_389);
nor U2907 (N_2907,In_209,In_69);
xor U2908 (N_2908,In_724,In_250);
nand U2909 (N_2909,In_371,In_283);
nor U2910 (N_2910,In_331,In_345);
or U2911 (N_2911,In_465,In_229);
or U2912 (N_2912,In_826,In_211);
or U2913 (N_2913,In_143,In_885);
or U2914 (N_2914,In_474,In_308);
or U2915 (N_2915,In_599,In_639);
or U2916 (N_2916,In_117,In_589);
xnor U2917 (N_2917,In_336,In_483);
xnor U2918 (N_2918,In_353,In_432);
and U2919 (N_2919,In_901,In_116);
and U2920 (N_2920,In_375,In_842);
nor U2921 (N_2921,In_245,In_959);
or U2922 (N_2922,In_810,In_767);
nand U2923 (N_2923,In_684,In_434);
nor U2924 (N_2924,In_900,In_315);
and U2925 (N_2925,In_746,In_824);
and U2926 (N_2926,In_359,In_582);
nor U2927 (N_2927,In_830,In_850);
or U2928 (N_2928,In_915,In_982);
xnor U2929 (N_2929,In_847,In_250);
nor U2930 (N_2930,In_475,In_720);
nor U2931 (N_2931,In_622,In_895);
nor U2932 (N_2932,In_700,In_212);
or U2933 (N_2933,In_305,In_633);
and U2934 (N_2934,In_8,In_751);
nand U2935 (N_2935,In_204,In_505);
nor U2936 (N_2936,In_800,In_212);
xnor U2937 (N_2937,In_678,In_684);
and U2938 (N_2938,In_54,In_968);
and U2939 (N_2939,In_316,In_214);
nand U2940 (N_2940,In_839,In_386);
and U2941 (N_2941,In_583,In_636);
xnor U2942 (N_2942,In_166,In_252);
and U2943 (N_2943,In_284,In_916);
nor U2944 (N_2944,In_237,In_464);
or U2945 (N_2945,In_306,In_111);
or U2946 (N_2946,In_454,In_947);
or U2947 (N_2947,In_174,In_322);
or U2948 (N_2948,In_11,In_268);
or U2949 (N_2949,In_10,In_379);
or U2950 (N_2950,In_786,In_222);
or U2951 (N_2951,In_744,In_83);
xnor U2952 (N_2952,In_270,In_658);
or U2953 (N_2953,In_248,In_793);
and U2954 (N_2954,In_477,In_620);
nor U2955 (N_2955,In_287,In_611);
nor U2956 (N_2956,In_324,In_275);
nor U2957 (N_2957,In_419,In_473);
nor U2958 (N_2958,In_620,In_432);
nand U2959 (N_2959,In_762,In_448);
nor U2960 (N_2960,In_332,In_307);
nand U2961 (N_2961,In_356,In_808);
and U2962 (N_2962,In_816,In_129);
nand U2963 (N_2963,In_165,In_641);
or U2964 (N_2964,In_112,In_197);
nor U2965 (N_2965,In_332,In_324);
or U2966 (N_2966,In_913,In_41);
nor U2967 (N_2967,In_349,In_287);
and U2968 (N_2968,In_916,In_870);
and U2969 (N_2969,In_820,In_978);
xor U2970 (N_2970,In_883,In_490);
nand U2971 (N_2971,In_27,In_603);
or U2972 (N_2972,In_110,In_176);
and U2973 (N_2973,In_867,In_393);
nand U2974 (N_2974,In_577,In_988);
and U2975 (N_2975,In_857,In_361);
nor U2976 (N_2976,In_936,In_397);
nand U2977 (N_2977,In_775,In_310);
nor U2978 (N_2978,In_324,In_488);
xor U2979 (N_2979,In_596,In_356);
xnor U2980 (N_2980,In_705,In_100);
or U2981 (N_2981,In_583,In_777);
and U2982 (N_2982,In_439,In_580);
nor U2983 (N_2983,In_806,In_640);
xnor U2984 (N_2984,In_754,In_941);
nand U2985 (N_2985,In_165,In_957);
or U2986 (N_2986,In_462,In_492);
or U2987 (N_2987,In_952,In_275);
xor U2988 (N_2988,In_535,In_343);
nand U2989 (N_2989,In_920,In_932);
or U2990 (N_2990,In_444,In_589);
nand U2991 (N_2991,In_586,In_283);
and U2992 (N_2992,In_806,In_167);
nor U2993 (N_2993,In_984,In_377);
and U2994 (N_2994,In_247,In_570);
nor U2995 (N_2995,In_594,In_606);
or U2996 (N_2996,In_488,In_925);
nor U2997 (N_2997,In_366,In_736);
or U2998 (N_2998,In_667,In_246);
nand U2999 (N_2999,In_398,In_415);
and U3000 (N_3000,In_938,In_548);
and U3001 (N_3001,In_415,In_430);
and U3002 (N_3002,In_632,In_167);
nand U3003 (N_3003,In_649,In_335);
or U3004 (N_3004,In_837,In_625);
nor U3005 (N_3005,In_273,In_787);
nor U3006 (N_3006,In_316,In_657);
xor U3007 (N_3007,In_361,In_124);
nor U3008 (N_3008,In_132,In_706);
and U3009 (N_3009,In_925,In_844);
nand U3010 (N_3010,In_280,In_130);
and U3011 (N_3011,In_954,In_766);
and U3012 (N_3012,In_262,In_650);
xnor U3013 (N_3013,In_833,In_114);
nor U3014 (N_3014,In_981,In_71);
and U3015 (N_3015,In_798,In_296);
and U3016 (N_3016,In_111,In_720);
or U3017 (N_3017,In_520,In_958);
or U3018 (N_3018,In_182,In_593);
and U3019 (N_3019,In_118,In_236);
or U3020 (N_3020,In_692,In_718);
xnor U3021 (N_3021,In_304,In_329);
nand U3022 (N_3022,In_637,In_539);
nor U3023 (N_3023,In_215,In_689);
nand U3024 (N_3024,In_884,In_793);
and U3025 (N_3025,In_503,In_894);
nor U3026 (N_3026,In_444,In_333);
nor U3027 (N_3027,In_389,In_233);
nor U3028 (N_3028,In_498,In_318);
xnor U3029 (N_3029,In_174,In_713);
nor U3030 (N_3030,In_49,In_793);
and U3031 (N_3031,In_409,In_458);
xnor U3032 (N_3032,In_503,In_410);
nor U3033 (N_3033,In_761,In_869);
xnor U3034 (N_3034,In_920,In_440);
and U3035 (N_3035,In_101,In_686);
xnor U3036 (N_3036,In_890,In_775);
xnor U3037 (N_3037,In_820,In_78);
nor U3038 (N_3038,In_495,In_521);
xnor U3039 (N_3039,In_724,In_94);
and U3040 (N_3040,In_948,In_372);
nor U3041 (N_3041,In_179,In_320);
nor U3042 (N_3042,In_142,In_98);
xor U3043 (N_3043,In_434,In_86);
nor U3044 (N_3044,In_643,In_134);
nor U3045 (N_3045,In_41,In_703);
or U3046 (N_3046,In_991,In_795);
or U3047 (N_3047,In_595,In_912);
and U3048 (N_3048,In_302,In_733);
nand U3049 (N_3049,In_840,In_564);
or U3050 (N_3050,In_192,In_889);
and U3051 (N_3051,In_940,In_499);
and U3052 (N_3052,In_822,In_153);
nand U3053 (N_3053,In_688,In_395);
nand U3054 (N_3054,In_533,In_745);
or U3055 (N_3055,In_176,In_996);
and U3056 (N_3056,In_957,In_327);
or U3057 (N_3057,In_135,In_42);
nor U3058 (N_3058,In_219,In_192);
or U3059 (N_3059,In_18,In_301);
nor U3060 (N_3060,In_131,In_755);
nand U3061 (N_3061,In_237,In_889);
and U3062 (N_3062,In_401,In_147);
and U3063 (N_3063,In_780,In_837);
xnor U3064 (N_3064,In_762,In_663);
and U3065 (N_3065,In_585,In_616);
and U3066 (N_3066,In_164,In_797);
or U3067 (N_3067,In_209,In_887);
nand U3068 (N_3068,In_671,In_7);
nor U3069 (N_3069,In_399,In_774);
nor U3070 (N_3070,In_711,In_589);
nand U3071 (N_3071,In_178,In_802);
or U3072 (N_3072,In_618,In_552);
nand U3073 (N_3073,In_655,In_892);
nor U3074 (N_3074,In_640,In_133);
nor U3075 (N_3075,In_376,In_589);
and U3076 (N_3076,In_469,In_282);
or U3077 (N_3077,In_268,In_828);
or U3078 (N_3078,In_675,In_92);
or U3079 (N_3079,In_435,In_684);
xnor U3080 (N_3080,In_882,In_210);
xor U3081 (N_3081,In_628,In_830);
and U3082 (N_3082,In_811,In_401);
and U3083 (N_3083,In_77,In_530);
nand U3084 (N_3084,In_525,In_825);
or U3085 (N_3085,In_329,In_928);
nor U3086 (N_3086,In_958,In_327);
or U3087 (N_3087,In_294,In_580);
nor U3088 (N_3088,In_600,In_896);
nor U3089 (N_3089,In_534,In_355);
xnor U3090 (N_3090,In_885,In_379);
nor U3091 (N_3091,In_694,In_594);
nand U3092 (N_3092,In_507,In_934);
xnor U3093 (N_3093,In_684,In_716);
nand U3094 (N_3094,In_212,In_457);
and U3095 (N_3095,In_553,In_549);
or U3096 (N_3096,In_773,In_479);
nand U3097 (N_3097,In_432,In_14);
or U3098 (N_3098,In_901,In_809);
or U3099 (N_3099,In_332,In_932);
nand U3100 (N_3100,In_985,In_289);
and U3101 (N_3101,In_912,In_863);
or U3102 (N_3102,In_481,In_404);
or U3103 (N_3103,In_952,In_57);
or U3104 (N_3104,In_220,In_986);
or U3105 (N_3105,In_910,In_221);
nand U3106 (N_3106,In_121,In_345);
nor U3107 (N_3107,In_994,In_628);
or U3108 (N_3108,In_512,In_743);
nor U3109 (N_3109,In_368,In_117);
or U3110 (N_3110,In_17,In_448);
or U3111 (N_3111,In_520,In_787);
nor U3112 (N_3112,In_701,In_719);
nand U3113 (N_3113,In_230,In_726);
or U3114 (N_3114,In_695,In_39);
or U3115 (N_3115,In_99,In_350);
nand U3116 (N_3116,In_942,In_101);
nand U3117 (N_3117,In_169,In_330);
xnor U3118 (N_3118,In_121,In_196);
nor U3119 (N_3119,In_434,In_626);
and U3120 (N_3120,In_80,In_623);
or U3121 (N_3121,In_2,In_215);
or U3122 (N_3122,In_80,In_457);
nor U3123 (N_3123,In_512,In_219);
nand U3124 (N_3124,In_456,In_652);
nor U3125 (N_3125,In_267,In_294);
nand U3126 (N_3126,In_308,In_609);
or U3127 (N_3127,In_851,In_351);
nand U3128 (N_3128,In_466,In_615);
nand U3129 (N_3129,In_55,In_409);
xor U3130 (N_3130,In_438,In_366);
or U3131 (N_3131,In_695,In_129);
nor U3132 (N_3132,In_963,In_37);
nand U3133 (N_3133,In_790,In_537);
xor U3134 (N_3134,In_328,In_978);
and U3135 (N_3135,In_308,In_725);
or U3136 (N_3136,In_68,In_787);
and U3137 (N_3137,In_120,In_323);
nor U3138 (N_3138,In_543,In_752);
and U3139 (N_3139,In_487,In_494);
and U3140 (N_3140,In_939,In_558);
and U3141 (N_3141,In_547,In_889);
nor U3142 (N_3142,In_942,In_711);
or U3143 (N_3143,In_603,In_345);
or U3144 (N_3144,In_300,In_58);
nand U3145 (N_3145,In_343,In_756);
nand U3146 (N_3146,In_390,In_512);
nand U3147 (N_3147,In_223,In_623);
nand U3148 (N_3148,In_509,In_454);
or U3149 (N_3149,In_140,In_41);
and U3150 (N_3150,In_276,In_851);
nand U3151 (N_3151,In_342,In_302);
and U3152 (N_3152,In_966,In_197);
and U3153 (N_3153,In_685,In_421);
or U3154 (N_3154,In_393,In_884);
or U3155 (N_3155,In_727,In_18);
and U3156 (N_3156,In_149,In_270);
xor U3157 (N_3157,In_784,In_380);
nor U3158 (N_3158,In_142,In_633);
nand U3159 (N_3159,In_444,In_673);
nor U3160 (N_3160,In_302,In_457);
or U3161 (N_3161,In_83,In_597);
nand U3162 (N_3162,In_788,In_235);
xnor U3163 (N_3163,In_877,In_160);
and U3164 (N_3164,In_217,In_943);
nor U3165 (N_3165,In_812,In_777);
nand U3166 (N_3166,In_762,In_300);
and U3167 (N_3167,In_938,In_821);
nor U3168 (N_3168,In_724,In_360);
nand U3169 (N_3169,In_787,In_420);
or U3170 (N_3170,In_70,In_120);
nand U3171 (N_3171,In_459,In_398);
nand U3172 (N_3172,In_629,In_745);
and U3173 (N_3173,In_693,In_464);
xnor U3174 (N_3174,In_4,In_652);
nand U3175 (N_3175,In_595,In_31);
nand U3176 (N_3176,In_438,In_698);
and U3177 (N_3177,In_181,In_871);
nor U3178 (N_3178,In_709,In_648);
nor U3179 (N_3179,In_907,In_758);
xnor U3180 (N_3180,In_201,In_291);
and U3181 (N_3181,In_371,In_942);
and U3182 (N_3182,In_771,In_633);
and U3183 (N_3183,In_778,In_410);
or U3184 (N_3184,In_236,In_308);
and U3185 (N_3185,In_123,In_1);
nor U3186 (N_3186,In_477,In_833);
or U3187 (N_3187,In_806,In_172);
xor U3188 (N_3188,In_343,In_406);
nor U3189 (N_3189,In_198,In_884);
nand U3190 (N_3190,In_325,In_747);
nand U3191 (N_3191,In_45,In_577);
and U3192 (N_3192,In_998,In_2);
nand U3193 (N_3193,In_158,In_439);
nand U3194 (N_3194,In_498,In_645);
and U3195 (N_3195,In_357,In_600);
nor U3196 (N_3196,In_252,In_427);
xnor U3197 (N_3197,In_922,In_918);
nor U3198 (N_3198,In_541,In_395);
nand U3199 (N_3199,In_603,In_53);
and U3200 (N_3200,In_95,In_741);
and U3201 (N_3201,In_431,In_538);
and U3202 (N_3202,In_780,In_498);
nand U3203 (N_3203,In_72,In_901);
or U3204 (N_3204,In_247,In_130);
or U3205 (N_3205,In_415,In_560);
or U3206 (N_3206,In_930,In_451);
or U3207 (N_3207,In_160,In_567);
nand U3208 (N_3208,In_917,In_253);
or U3209 (N_3209,In_174,In_894);
or U3210 (N_3210,In_733,In_112);
xnor U3211 (N_3211,In_463,In_328);
xnor U3212 (N_3212,In_121,In_641);
xnor U3213 (N_3213,In_362,In_275);
nor U3214 (N_3214,In_586,In_85);
nand U3215 (N_3215,In_817,In_285);
nor U3216 (N_3216,In_627,In_63);
nand U3217 (N_3217,In_6,In_82);
or U3218 (N_3218,In_812,In_836);
and U3219 (N_3219,In_741,In_128);
nor U3220 (N_3220,In_881,In_394);
nor U3221 (N_3221,In_251,In_539);
or U3222 (N_3222,In_201,In_712);
xor U3223 (N_3223,In_413,In_222);
nor U3224 (N_3224,In_626,In_396);
or U3225 (N_3225,In_722,In_380);
nand U3226 (N_3226,In_34,In_740);
and U3227 (N_3227,In_973,In_755);
and U3228 (N_3228,In_457,In_300);
nand U3229 (N_3229,In_273,In_216);
and U3230 (N_3230,In_290,In_505);
or U3231 (N_3231,In_6,In_57);
nand U3232 (N_3232,In_126,In_699);
and U3233 (N_3233,In_578,In_124);
or U3234 (N_3234,In_106,In_919);
nand U3235 (N_3235,In_995,In_687);
nand U3236 (N_3236,In_115,In_451);
or U3237 (N_3237,In_101,In_853);
nor U3238 (N_3238,In_432,In_59);
nor U3239 (N_3239,In_21,In_528);
xnor U3240 (N_3240,In_439,In_938);
and U3241 (N_3241,In_849,In_673);
or U3242 (N_3242,In_30,In_708);
and U3243 (N_3243,In_841,In_94);
nor U3244 (N_3244,In_414,In_125);
nor U3245 (N_3245,In_307,In_994);
and U3246 (N_3246,In_845,In_873);
or U3247 (N_3247,In_920,In_502);
nor U3248 (N_3248,In_311,In_265);
nor U3249 (N_3249,In_887,In_498);
and U3250 (N_3250,In_321,In_759);
and U3251 (N_3251,In_177,In_92);
or U3252 (N_3252,In_586,In_587);
nor U3253 (N_3253,In_382,In_545);
nor U3254 (N_3254,In_671,In_69);
xnor U3255 (N_3255,In_692,In_662);
nor U3256 (N_3256,In_363,In_373);
or U3257 (N_3257,In_562,In_155);
nor U3258 (N_3258,In_95,In_61);
and U3259 (N_3259,In_288,In_733);
xnor U3260 (N_3260,In_737,In_145);
nand U3261 (N_3261,In_85,In_718);
and U3262 (N_3262,In_941,In_783);
xor U3263 (N_3263,In_130,In_431);
and U3264 (N_3264,In_450,In_564);
nor U3265 (N_3265,In_879,In_375);
nand U3266 (N_3266,In_26,In_916);
or U3267 (N_3267,In_755,In_229);
or U3268 (N_3268,In_958,In_18);
nor U3269 (N_3269,In_20,In_984);
nor U3270 (N_3270,In_57,In_846);
nor U3271 (N_3271,In_169,In_615);
xnor U3272 (N_3272,In_829,In_37);
nor U3273 (N_3273,In_665,In_481);
nand U3274 (N_3274,In_250,In_220);
nand U3275 (N_3275,In_986,In_847);
and U3276 (N_3276,In_772,In_204);
xnor U3277 (N_3277,In_44,In_553);
nand U3278 (N_3278,In_192,In_943);
or U3279 (N_3279,In_145,In_743);
xor U3280 (N_3280,In_779,In_905);
and U3281 (N_3281,In_129,In_781);
nor U3282 (N_3282,In_583,In_516);
nand U3283 (N_3283,In_866,In_712);
nand U3284 (N_3284,In_223,In_312);
and U3285 (N_3285,In_822,In_201);
nand U3286 (N_3286,In_210,In_119);
nor U3287 (N_3287,In_415,In_328);
nor U3288 (N_3288,In_154,In_327);
and U3289 (N_3289,In_521,In_331);
or U3290 (N_3290,In_61,In_514);
or U3291 (N_3291,In_164,In_312);
and U3292 (N_3292,In_565,In_344);
or U3293 (N_3293,In_833,In_589);
nand U3294 (N_3294,In_965,In_337);
nand U3295 (N_3295,In_671,In_776);
nor U3296 (N_3296,In_445,In_777);
nand U3297 (N_3297,In_770,In_609);
nand U3298 (N_3298,In_720,In_342);
nand U3299 (N_3299,In_497,In_806);
nor U3300 (N_3300,In_800,In_309);
or U3301 (N_3301,In_726,In_785);
and U3302 (N_3302,In_728,In_172);
or U3303 (N_3303,In_320,In_276);
nand U3304 (N_3304,In_236,In_878);
and U3305 (N_3305,In_978,In_847);
and U3306 (N_3306,In_216,In_935);
and U3307 (N_3307,In_305,In_895);
xor U3308 (N_3308,In_669,In_155);
nor U3309 (N_3309,In_726,In_481);
or U3310 (N_3310,In_9,In_353);
and U3311 (N_3311,In_833,In_117);
nand U3312 (N_3312,In_863,In_792);
nand U3313 (N_3313,In_837,In_672);
and U3314 (N_3314,In_389,In_765);
and U3315 (N_3315,In_632,In_316);
nor U3316 (N_3316,In_358,In_892);
nand U3317 (N_3317,In_889,In_56);
or U3318 (N_3318,In_365,In_350);
or U3319 (N_3319,In_273,In_138);
or U3320 (N_3320,In_709,In_720);
nor U3321 (N_3321,In_629,In_407);
or U3322 (N_3322,In_823,In_280);
nor U3323 (N_3323,In_652,In_761);
and U3324 (N_3324,In_17,In_579);
nor U3325 (N_3325,In_395,In_897);
and U3326 (N_3326,In_845,In_841);
nor U3327 (N_3327,In_656,In_943);
nor U3328 (N_3328,In_932,In_653);
nand U3329 (N_3329,In_561,In_292);
nand U3330 (N_3330,In_50,In_60);
or U3331 (N_3331,In_971,In_917);
or U3332 (N_3332,In_100,In_35);
nand U3333 (N_3333,In_699,In_712);
nor U3334 (N_3334,In_790,In_125);
or U3335 (N_3335,In_556,In_872);
nand U3336 (N_3336,In_914,In_357);
or U3337 (N_3337,In_274,In_496);
nand U3338 (N_3338,In_60,In_123);
and U3339 (N_3339,In_218,In_408);
or U3340 (N_3340,In_988,In_618);
nand U3341 (N_3341,In_837,In_176);
and U3342 (N_3342,In_709,In_479);
or U3343 (N_3343,In_752,In_250);
nand U3344 (N_3344,In_384,In_394);
xnor U3345 (N_3345,In_842,In_205);
nor U3346 (N_3346,In_75,In_428);
nand U3347 (N_3347,In_782,In_592);
nor U3348 (N_3348,In_522,In_49);
or U3349 (N_3349,In_420,In_530);
nand U3350 (N_3350,In_521,In_861);
or U3351 (N_3351,In_641,In_797);
or U3352 (N_3352,In_533,In_671);
nand U3353 (N_3353,In_230,In_844);
nor U3354 (N_3354,In_100,In_173);
nand U3355 (N_3355,In_440,In_766);
or U3356 (N_3356,In_183,In_99);
nand U3357 (N_3357,In_587,In_786);
nand U3358 (N_3358,In_987,In_418);
or U3359 (N_3359,In_740,In_499);
nand U3360 (N_3360,In_535,In_514);
nand U3361 (N_3361,In_727,In_135);
or U3362 (N_3362,In_953,In_982);
nand U3363 (N_3363,In_490,In_254);
nand U3364 (N_3364,In_872,In_419);
and U3365 (N_3365,In_88,In_149);
xnor U3366 (N_3366,In_425,In_287);
nand U3367 (N_3367,In_280,In_727);
nand U3368 (N_3368,In_460,In_786);
nand U3369 (N_3369,In_327,In_577);
or U3370 (N_3370,In_242,In_117);
or U3371 (N_3371,In_353,In_864);
nor U3372 (N_3372,In_788,In_918);
nand U3373 (N_3373,In_10,In_94);
or U3374 (N_3374,In_265,In_167);
xnor U3375 (N_3375,In_417,In_28);
or U3376 (N_3376,In_577,In_371);
nand U3377 (N_3377,In_704,In_838);
nor U3378 (N_3378,In_721,In_345);
or U3379 (N_3379,In_697,In_689);
and U3380 (N_3380,In_121,In_398);
nand U3381 (N_3381,In_343,In_149);
nand U3382 (N_3382,In_421,In_227);
nand U3383 (N_3383,In_763,In_684);
nand U3384 (N_3384,In_953,In_187);
or U3385 (N_3385,In_265,In_643);
xor U3386 (N_3386,In_204,In_181);
and U3387 (N_3387,In_90,In_422);
nor U3388 (N_3388,In_408,In_428);
or U3389 (N_3389,In_293,In_840);
or U3390 (N_3390,In_109,In_490);
and U3391 (N_3391,In_619,In_890);
or U3392 (N_3392,In_613,In_215);
nand U3393 (N_3393,In_396,In_659);
nand U3394 (N_3394,In_750,In_365);
xnor U3395 (N_3395,In_832,In_559);
or U3396 (N_3396,In_181,In_602);
xnor U3397 (N_3397,In_189,In_219);
nand U3398 (N_3398,In_776,In_382);
nor U3399 (N_3399,In_912,In_579);
or U3400 (N_3400,In_396,In_857);
and U3401 (N_3401,In_217,In_846);
nand U3402 (N_3402,In_865,In_670);
or U3403 (N_3403,In_386,In_618);
xnor U3404 (N_3404,In_623,In_633);
or U3405 (N_3405,In_635,In_974);
or U3406 (N_3406,In_105,In_639);
nor U3407 (N_3407,In_80,In_548);
nor U3408 (N_3408,In_997,In_815);
nand U3409 (N_3409,In_575,In_874);
xnor U3410 (N_3410,In_664,In_662);
or U3411 (N_3411,In_934,In_273);
or U3412 (N_3412,In_936,In_406);
or U3413 (N_3413,In_252,In_259);
or U3414 (N_3414,In_594,In_501);
or U3415 (N_3415,In_432,In_316);
nor U3416 (N_3416,In_700,In_724);
nand U3417 (N_3417,In_305,In_181);
and U3418 (N_3418,In_151,In_741);
nor U3419 (N_3419,In_655,In_345);
nor U3420 (N_3420,In_102,In_389);
xnor U3421 (N_3421,In_126,In_300);
nor U3422 (N_3422,In_337,In_304);
nor U3423 (N_3423,In_391,In_966);
or U3424 (N_3424,In_695,In_383);
nor U3425 (N_3425,In_353,In_241);
or U3426 (N_3426,In_112,In_852);
nand U3427 (N_3427,In_53,In_687);
nor U3428 (N_3428,In_341,In_329);
nor U3429 (N_3429,In_25,In_240);
nor U3430 (N_3430,In_994,In_910);
nand U3431 (N_3431,In_890,In_105);
nand U3432 (N_3432,In_685,In_280);
and U3433 (N_3433,In_523,In_694);
xor U3434 (N_3434,In_701,In_574);
and U3435 (N_3435,In_308,In_643);
nor U3436 (N_3436,In_427,In_993);
or U3437 (N_3437,In_181,In_733);
nor U3438 (N_3438,In_284,In_532);
nor U3439 (N_3439,In_76,In_455);
or U3440 (N_3440,In_251,In_176);
xor U3441 (N_3441,In_386,In_794);
or U3442 (N_3442,In_15,In_413);
or U3443 (N_3443,In_191,In_47);
or U3444 (N_3444,In_696,In_923);
and U3445 (N_3445,In_922,In_485);
and U3446 (N_3446,In_825,In_866);
or U3447 (N_3447,In_836,In_611);
and U3448 (N_3448,In_43,In_638);
nand U3449 (N_3449,In_880,In_182);
and U3450 (N_3450,In_256,In_271);
or U3451 (N_3451,In_924,In_505);
xnor U3452 (N_3452,In_774,In_111);
nor U3453 (N_3453,In_380,In_418);
and U3454 (N_3454,In_878,In_237);
or U3455 (N_3455,In_391,In_335);
nand U3456 (N_3456,In_200,In_643);
and U3457 (N_3457,In_234,In_456);
nor U3458 (N_3458,In_167,In_694);
nand U3459 (N_3459,In_279,In_614);
and U3460 (N_3460,In_799,In_85);
and U3461 (N_3461,In_759,In_415);
nand U3462 (N_3462,In_762,In_935);
or U3463 (N_3463,In_205,In_958);
and U3464 (N_3464,In_47,In_838);
nor U3465 (N_3465,In_949,In_613);
and U3466 (N_3466,In_380,In_493);
or U3467 (N_3467,In_52,In_169);
nand U3468 (N_3468,In_790,In_400);
xor U3469 (N_3469,In_971,In_72);
nor U3470 (N_3470,In_623,In_555);
or U3471 (N_3471,In_695,In_408);
nor U3472 (N_3472,In_75,In_39);
or U3473 (N_3473,In_529,In_474);
nor U3474 (N_3474,In_984,In_100);
nor U3475 (N_3475,In_672,In_524);
nand U3476 (N_3476,In_90,In_805);
nor U3477 (N_3477,In_892,In_467);
nand U3478 (N_3478,In_880,In_515);
and U3479 (N_3479,In_619,In_21);
and U3480 (N_3480,In_731,In_988);
nor U3481 (N_3481,In_205,In_968);
nor U3482 (N_3482,In_836,In_528);
nor U3483 (N_3483,In_163,In_180);
or U3484 (N_3484,In_509,In_442);
nand U3485 (N_3485,In_777,In_354);
and U3486 (N_3486,In_476,In_431);
nor U3487 (N_3487,In_27,In_877);
xor U3488 (N_3488,In_840,In_669);
nand U3489 (N_3489,In_512,In_88);
or U3490 (N_3490,In_465,In_190);
nand U3491 (N_3491,In_695,In_972);
or U3492 (N_3492,In_479,In_978);
nand U3493 (N_3493,In_885,In_935);
nor U3494 (N_3494,In_949,In_850);
or U3495 (N_3495,In_818,In_17);
nand U3496 (N_3496,In_966,In_292);
nor U3497 (N_3497,In_134,In_535);
nand U3498 (N_3498,In_130,In_229);
nor U3499 (N_3499,In_33,In_980);
and U3500 (N_3500,In_199,In_944);
nand U3501 (N_3501,In_437,In_216);
nand U3502 (N_3502,In_411,In_570);
or U3503 (N_3503,In_935,In_472);
and U3504 (N_3504,In_360,In_587);
nand U3505 (N_3505,In_662,In_381);
nand U3506 (N_3506,In_719,In_885);
or U3507 (N_3507,In_266,In_708);
or U3508 (N_3508,In_123,In_371);
and U3509 (N_3509,In_505,In_408);
nand U3510 (N_3510,In_466,In_748);
xnor U3511 (N_3511,In_535,In_788);
nand U3512 (N_3512,In_252,In_990);
xor U3513 (N_3513,In_139,In_915);
and U3514 (N_3514,In_981,In_549);
xor U3515 (N_3515,In_52,In_759);
nor U3516 (N_3516,In_784,In_55);
and U3517 (N_3517,In_255,In_383);
nor U3518 (N_3518,In_983,In_246);
nand U3519 (N_3519,In_617,In_148);
and U3520 (N_3520,In_808,In_573);
nand U3521 (N_3521,In_90,In_339);
nor U3522 (N_3522,In_109,In_516);
nor U3523 (N_3523,In_726,In_756);
nor U3524 (N_3524,In_729,In_175);
nand U3525 (N_3525,In_795,In_295);
xnor U3526 (N_3526,In_838,In_368);
nor U3527 (N_3527,In_733,In_599);
or U3528 (N_3528,In_123,In_132);
nand U3529 (N_3529,In_208,In_926);
xor U3530 (N_3530,In_724,In_319);
nand U3531 (N_3531,In_288,In_567);
and U3532 (N_3532,In_630,In_870);
and U3533 (N_3533,In_187,In_796);
and U3534 (N_3534,In_115,In_441);
and U3535 (N_3535,In_167,In_569);
nor U3536 (N_3536,In_965,In_940);
nand U3537 (N_3537,In_931,In_963);
nor U3538 (N_3538,In_410,In_379);
nand U3539 (N_3539,In_231,In_284);
nand U3540 (N_3540,In_361,In_924);
nand U3541 (N_3541,In_351,In_894);
nand U3542 (N_3542,In_319,In_72);
and U3543 (N_3543,In_67,In_834);
nand U3544 (N_3544,In_5,In_148);
nor U3545 (N_3545,In_795,In_349);
nor U3546 (N_3546,In_239,In_605);
nor U3547 (N_3547,In_718,In_847);
and U3548 (N_3548,In_93,In_592);
nor U3549 (N_3549,In_643,In_433);
or U3550 (N_3550,In_366,In_163);
xor U3551 (N_3551,In_718,In_39);
xor U3552 (N_3552,In_757,In_242);
or U3553 (N_3553,In_524,In_804);
nor U3554 (N_3554,In_507,In_771);
nand U3555 (N_3555,In_630,In_736);
and U3556 (N_3556,In_917,In_666);
and U3557 (N_3557,In_825,In_303);
nor U3558 (N_3558,In_589,In_427);
or U3559 (N_3559,In_997,In_675);
xor U3560 (N_3560,In_829,In_366);
and U3561 (N_3561,In_747,In_332);
or U3562 (N_3562,In_254,In_18);
nor U3563 (N_3563,In_277,In_980);
or U3564 (N_3564,In_596,In_943);
nand U3565 (N_3565,In_538,In_531);
or U3566 (N_3566,In_379,In_505);
nand U3567 (N_3567,In_392,In_265);
or U3568 (N_3568,In_361,In_609);
or U3569 (N_3569,In_439,In_825);
or U3570 (N_3570,In_180,In_806);
or U3571 (N_3571,In_864,In_471);
nand U3572 (N_3572,In_761,In_162);
nand U3573 (N_3573,In_937,In_523);
and U3574 (N_3574,In_290,In_888);
or U3575 (N_3575,In_125,In_196);
and U3576 (N_3576,In_601,In_986);
nand U3577 (N_3577,In_295,In_275);
nand U3578 (N_3578,In_122,In_649);
nor U3579 (N_3579,In_85,In_406);
and U3580 (N_3580,In_440,In_261);
nand U3581 (N_3581,In_62,In_443);
nor U3582 (N_3582,In_830,In_81);
nor U3583 (N_3583,In_363,In_225);
or U3584 (N_3584,In_391,In_218);
and U3585 (N_3585,In_464,In_85);
nand U3586 (N_3586,In_330,In_971);
or U3587 (N_3587,In_67,In_785);
or U3588 (N_3588,In_978,In_507);
and U3589 (N_3589,In_860,In_979);
nor U3590 (N_3590,In_107,In_316);
nor U3591 (N_3591,In_580,In_281);
nand U3592 (N_3592,In_426,In_836);
nor U3593 (N_3593,In_460,In_739);
nor U3594 (N_3594,In_834,In_974);
or U3595 (N_3595,In_663,In_491);
or U3596 (N_3596,In_912,In_706);
nand U3597 (N_3597,In_818,In_973);
nand U3598 (N_3598,In_82,In_665);
or U3599 (N_3599,In_799,In_748);
nor U3600 (N_3600,In_174,In_286);
or U3601 (N_3601,In_950,In_641);
and U3602 (N_3602,In_273,In_635);
or U3603 (N_3603,In_38,In_966);
xor U3604 (N_3604,In_199,In_98);
and U3605 (N_3605,In_882,In_814);
and U3606 (N_3606,In_537,In_876);
and U3607 (N_3607,In_289,In_779);
nor U3608 (N_3608,In_880,In_695);
or U3609 (N_3609,In_150,In_978);
or U3610 (N_3610,In_903,In_79);
and U3611 (N_3611,In_854,In_60);
or U3612 (N_3612,In_284,In_31);
or U3613 (N_3613,In_916,In_744);
nand U3614 (N_3614,In_195,In_13);
nor U3615 (N_3615,In_192,In_850);
nand U3616 (N_3616,In_7,In_980);
and U3617 (N_3617,In_973,In_884);
or U3618 (N_3618,In_964,In_276);
and U3619 (N_3619,In_274,In_528);
and U3620 (N_3620,In_13,In_574);
xnor U3621 (N_3621,In_666,In_660);
or U3622 (N_3622,In_193,In_160);
xor U3623 (N_3623,In_700,In_517);
nand U3624 (N_3624,In_827,In_953);
nand U3625 (N_3625,In_88,In_152);
nor U3626 (N_3626,In_921,In_464);
nand U3627 (N_3627,In_315,In_638);
nand U3628 (N_3628,In_360,In_0);
xor U3629 (N_3629,In_115,In_476);
or U3630 (N_3630,In_498,In_940);
nand U3631 (N_3631,In_532,In_441);
and U3632 (N_3632,In_191,In_967);
or U3633 (N_3633,In_824,In_974);
and U3634 (N_3634,In_609,In_147);
nand U3635 (N_3635,In_215,In_33);
and U3636 (N_3636,In_117,In_414);
nand U3637 (N_3637,In_624,In_10);
and U3638 (N_3638,In_205,In_326);
or U3639 (N_3639,In_771,In_346);
and U3640 (N_3640,In_452,In_400);
and U3641 (N_3641,In_384,In_141);
and U3642 (N_3642,In_169,In_877);
or U3643 (N_3643,In_8,In_866);
nor U3644 (N_3644,In_164,In_364);
nor U3645 (N_3645,In_665,In_169);
and U3646 (N_3646,In_224,In_752);
and U3647 (N_3647,In_877,In_521);
or U3648 (N_3648,In_911,In_357);
and U3649 (N_3649,In_906,In_691);
or U3650 (N_3650,In_190,In_972);
and U3651 (N_3651,In_51,In_613);
or U3652 (N_3652,In_253,In_661);
and U3653 (N_3653,In_520,In_856);
nand U3654 (N_3654,In_904,In_401);
nor U3655 (N_3655,In_469,In_647);
or U3656 (N_3656,In_834,In_822);
nor U3657 (N_3657,In_958,In_277);
and U3658 (N_3658,In_70,In_962);
and U3659 (N_3659,In_465,In_274);
xnor U3660 (N_3660,In_374,In_663);
nor U3661 (N_3661,In_242,In_545);
nand U3662 (N_3662,In_163,In_286);
nor U3663 (N_3663,In_355,In_599);
and U3664 (N_3664,In_932,In_784);
or U3665 (N_3665,In_288,In_121);
and U3666 (N_3666,In_66,In_274);
or U3667 (N_3667,In_295,In_87);
nor U3668 (N_3668,In_222,In_565);
nor U3669 (N_3669,In_805,In_747);
and U3670 (N_3670,In_523,In_940);
nand U3671 (N_3671,In_657,In_232);
nand U3672 (N_3672,In_157,In_768);
nand U3673 (N_3673,In_71,In_0);
xor U3674 (N_3674,In_462,In_275);
or U3675 (N_3675,In_960,In_9);
and U3676 (N_3676,In_200,In_67);
or U3677 (N_3677,In_620,In_869);
nor U3678 (N_3678,In_464,In_319);
nand U3679 (N_3679,In_852,In_973);
xor U3680 (N_3680,In_248,In_185);
nand U3681 (N_3681,In_455,In_848);
nand U3682 (N_3682,In_637,In_786);
and U3683 (N_3683,In_784,In_94);
nor U3684 (N_3684,In_76,In_642);
or U3685 (N_3685,In_729,In_889);
nor U3686 (N_3686,In_504,In_874);
nor U3687 (N_3687,In_896,In_887);
xor U3688 (N_3688,In_803,In_457);
and U3689 (N_3689,In_719,In_570);
xnor U3690 (N_3690,In_86,In_751);
nor U3691 (N_3691,In_346,In_420);
nor U3692 (N_3692,In_882,In_122);
or U3693 (N_3693,In_211,In_223);
nand U3694 (N_3694,In_363,In_195);
xnor U3695 (N_3695,In_389,In_224);
nand U3696 (N_3696,In_39,In_292);
nand U3697 (N_3697,In_578,In_978);
nand U3698 (N_3698,In_923,In_163);
and U3699 (N_3699,In_766,In_852);
nor U3700 (N_3700,In_527,In_788);
nand U3701 (N_3701,In_400,In_20);
nor U3702 (N_3702,In_290,In_254);
and U3703 (N_3703,In_618,In_172);
nor U3704 (N_3704,In_50,In_138);
or U3705 (N_3705,In_24,In_213);
nor U3706 (N_3706,In_383,In_17);
nand U3707 (N_3707,In_311,In_772);
nand U3708 (N_3708,In_125,In_50);
xor U3709 (N_3709,In_758,In_85);
nand U3710 (N_3710,In_84,In_815);
nand U3711 (N_3711,In_553,In_719);
nor U3712 (N_3712,In_343,In_562);
and U3713 (N_3713,In_561,In_65);
and U3714 (N_3714,In_330,In_230);
or U3715 (N_3715,In_825,In_928);
or U3716 (N_3716,In_442,In_527);
nand U3717 (N_3717,In_259,In_387);
nor U3718 (N_3718,In_826,In_678);
and U3719 (N_3719,In_440,In_227);
or U3720 (N_3720,In_182,In_40);
nor U3721 (N_3721,In_524,In_58);
or U3722 (N_3722,In_518,In_345);
or U3723 (N_3723,In_626,In_198);
or U3724 (N_3724,In_126,In_191);
and U3725 (N_3725,In_870,In_819);
xnor U3726 (N_3726,In_256,In_59);
and U3727 (N_3727,In_434,In_354);
or U3728 (N_3728,In_813,In_489);
and U3729 (N_3729,In_318,In_66);
or U3730 (N_3730,In_168,In_763);
nand U3731 (N_3731,In_429,In_774);
or U3732 (N_3732,In_108,In_459);
nand U3733 (N_3733,In_208,In_693);
nor U3734 (N_3734,In_831,In_225);
nor U3735 (N_3735,In_408,In_839);
and U3736 (N_3736,In_779,In_531);
or U3737 (N_3737,In_351,In_927);
and U3738 (N_3738,In_497,In_192);
or U3739 (N_3739,In_943,In_524);
nor U3740 (N_3740,In_414,In_923);
and U3741 (N_3741,In_785,In_269);
or U3742 (N_3742,In_868,In_668);
and U3743 (N_3743,In_339,In_913);
or U3744 (N_3744,In_902,In_776);
nor U3745 (N_3745,In_222,In_274);
or U3746 (N_3746,In_364,In_459);
nor U3747 (N_3747,In_679,In_377);
xor U3748 (N_3748,In_794,In_282);
nor U3749 (N_3749,In_810,In_617);
nand U3750 (N_3750,In_933,In_996);
or U3751 (N_3751,In_310,In_30);
and U3752 (N_3752,In_917,In_166);
or U3753 (N_3753,In_626,In_140);
nor U3754 (N_3754,In_170,In_418);
nand U3755 (N_3755,In_808,In_728);
and U3756 (N_3756,In_255,In_289);
xor U3757 (N_3757,In_570,In_280);
nor U3758 (N_3758,In_447,In_642);
nor U3759 (N_3759,In_381,In_676);
nand U3760 (N_3760,In_936,In_679);
nand U3761 (N_3761,In_476,In_701);
or U3762 (N_3762,In_244,In_534);
and U3763 (N_3763,In_589,In_153);
or U3764 (N_3764,In_162,In_257);
nor U3765 (N_3765,In_49,In_759);
nor U3766 (N_3766,In_437,In_815);
nand U3767 (N_3767,In_810,In_700);
nand U3768 (N_3768,In_948,In_577);
or U3769 (N_3769,In_176,In_511);
nor U3770 (N_3770,In_463,In_527);
or U3771 (N_3771,In_0,In_103);
and U3772 (N_3772,In_761,In_888);
nor U3773 (N_3773,In_26,In_37);
nand U3774 (N_3774,In_372,In_366);
or U3775 (N_3775,In_54,In_565);
or U3776 (N_3776,In_950,In_364);
and U3777 (N_3777,In_597,In_458);
or U3778 (N_3778,In_950,In_149);
nor U3779 (N_3779,In_589,In_425);
nand U3780 (N_3780,In_595,In_275);
nor U3781 (N_3781,In_757,In_97);
or U3782 (N_3782,In_593,In_347);
xor U3783 (N_3783,In_371,In_370);
nand U3784 (N_3784,In_885,In_438);
nor U3785 (N_3785,In_214,In_764);
and U3786 (N_3786,In_339,In_365);
xor U3787 (N_3787,In_123,In_919);
and U3788 (N_3788,In_37,In_769);
nand U3789 (N_3789,In_588,In_678);
or U3790 (N_3790,In_855,In_164);
or U3791 (N_3791,In_384,In_661);
or U3792 (N_3792,In_990,In_145);
or U3793 (N_3793,In_779,In_168);
xor U3794 (N_3794,In_899,In_705);
nor U3795 (N_3795,In_121,In_532);
nand U3796 (N_3796,In_153,In_793);
or U3797 (N_3797,In_454,In_760);
xnor U3798 (N_3798,In_791,In_362);
or U3799 (N_3799,In_344,In_155);
xnor U3800 (N_3800,In_855,In_761);
nand U3801 (N_3801,In_667,In_751);
or U3802 (N_3802,In_142,In_12);
and U3803 (N_3803,In_977,In_520);
nand U3804 (N_3804,In_413,In_914);
and U3805 (N_3805,In_781,In_66);
or U3806 (N_3806,In_690,In_844);
or U3807 (N_3807,In_776,In_795);
nor U3808 (N_3808,In_774,In_43);
nand U3809 (N_3809,In_270,In_134);
and U3810 (N_3810,In_988,In_723);
and U3811 (N_3811,In_174,In_14);
or U3812 (N_3812,In_654,In_247);
and U3813 (N_3813,In_696,In_37);
or U3814 (N_3814,In_319,In_749);
and U3815 (N_3815,In_400,In_49);
nand U3816 (N_3816,In_385,In_905);
and U3817 (N_3817,In_226,In_768);
nor U3818 (N_3818,In_241,In_338);
nor U3819 (N_3819,In_846,In_126);
or U3820 (N_3820,In_397,In_706);
nand U3821 (N_3821,In_234,In_398);
nor U3822 (N_3822,In_777,In_513);
xor U3823 (N_3823,In_797,In_511);
and U3824 (N_3824,In_952,In_505);
nand U3825 (N_3825,In_355,In_443);
nand U3826 (N_3826,In_947,In_184);
and U3827 (N_3827,In_483,In_344);
nand U3828 (N_3828,In_418,In_177);
xnor U3829 (N_3829,In_776,In_310);
and U3830 (N_3830,In_41,In_153);
xor U3831 (N_3831,In_22,In_660);
and U3832 (N_3832,In_697,In_809);
nand U3833 (N_3833,In_914,In_955);
nor U3834 (N_3834,In_128,In_337);
or U3835 (N_3835,In_414,In_634);
nand U3836 (N_3836,In_317,In_152);
nor U3837 (N_3837,In_881,In_577);
and U3838 (N_3838,In_244,In_935);
xor U3839 (N_3839,In_912,In_425);
or U3840 (N_3840,In_905,In_295);
and U3841 (N_3841,In_26,In_218);
or U3842 (N_3842,In_940,In_553);
nand U3843 (N_3843,In_860,In_862);
and U3844 (N_3844,In_593,In_443);
or U3845 (N_3845,In_578,In_820);
nand U3846 (N_3846,In_373,In_39);
nor U3847 (N_3847,In_822,In_114);
or U3848 (N_3848,In_169,In_913);
or U3849 (N_3849,In_174,In_527);
and U3850 (N_3850,In_969,In_357);
nor U3851 (N_3851,In_609,In_169);
nand U3852 (N_3852,In_785,In_350);
nor U3853 (N_3853,In_204,In_155);
and U3854 (N_3854,In_954,In_570);
and U3855 (N_3855,In_561,In_70);
and U3856 (N_3856,In_938,In_550);
nor U3857 (N_3857,In_448,In_234);
nand U3858 (N_3858,In_305,In_3);
nand U3859 (N_3859,In_754,In_360);
nand U3860 (N_3860,In_65,In_183);
and U3861 (N_3861,In_418,In_73);
nand U3862 (N_3862,In_110,In_183);
and U3863 (N_3863,In_745,In_323);
nand U3864 (N_3864,In_641,In_758);
or U3865 (N_3865,In_571,In_726);
or U3866 (N_3866,In_516,In_779);
or U3867 (N_3867,In_125,In_529);
xnor U3868 (N_3868,In_523,In_885);
nor U3869 (N_3869,In_516,In_437);
nand U3870 (N_3870,In_579,In_840);
nand U3871 (N_3871,In_974,In_310);
nand U3872 (N_3872,In_734,In_725);
and U3873 (N_3873,In_252,In_317);
nor U3874 (N_3874,In_99,In_648);
and U3875 (N_3875,In_589,In_323);
nor U3876 (N_3876,In_454,In_237);
nand U3877 (N_3877,In_236,In_111);
xnor U3878 (N_3878,In_939,In_386);
and U3879 (N_3879,In_651,In_529);
and U3880 (N_3880,In_652,In_685);
or U3881 (N_3881,In_357,In_845);
and U3882 (N_3882,In_102,In_666);
nand U3883 (N_3883,In_702,In_690);
and U3884 (N_3884,In_619,In_613);
nand U3885 (N_3885,In_474,In_626);
xor U3886 (N_3886,In_962,In_285);
nand U3887 (N_3887,In_641,In_841);
and U3888 (N_3888,In_273,In_760);
or U3889 (N_3889,In_67,In_98);
nand U3890 (N_3890,In_614,In_790);
xor U3891 (N_3891,In_69,In_454);
xnor U3892 (N_3892,In_450,In_577);
nand U3893 (N_3893,In_893,In_758);
nand U3894 (N_3894,In_328,In_93);
nor U3895 (N_3895,In_358,In_72);
and U3896 (N_3896,In_136,In_936);
nor U3897 (N_3897,In_834,In_516);
or U3898 (N_3898,In_323,In_376);
nor U3899 (N_3899,In_879,In_803);
or U3900 (N_3900,In_568,In_228);
nand U3901 (N_3901,In_872,In_632);
xor U3902 (N_3902,In_547,In_849);
or U3903 (N_3903,In_319,In_965);
nor U3904 (N_3904,In_985,In_909);
and U3905 (N_3905,In_935,In_941);
and U3906 (N_3906,In_807,In_4);
xnor U3907 (N_3907,In_286,In_722);
and U3908 (N_3908,In_200,In_993);
or U3909 (N_3909,In_473,In_984);
or U3910 (N_3910,In_357,In_875);
nor U3911 (N_3911,In_796,In_527);
and U3912 (N_3912,In_690,In_659);
or U3913 (N_3913,In_835,In_997);
nand U3914 (N_3914,In_138,In_987);
or U3915 (N_3915,In_629,In_275);
nand U3916 (N_3916,In_937,In_722);
nor U3917 (N_3917,In_159,In_477);
or U3918 (N_3918,In_874,In_89);
nor U3919 (N_3919,In_20,In_906);
and U3920 (N_3920,In_624,In_972);
or U3921 (N_3921,In_925,In_879);
and U3922 (N_3922,In_294,In_619);
nor U3923 (N_3923,In_480,In_712);
xor U3924 (N_3924,In_71,In_597);
nand U3925 (N_3925,In_652,In_803);
nor U3926 (N_3926,In_843,In_342);
or U3927 (N_3927,In_43,In_644);
or U3928 (N_3928,In_226,In_535);
and U3929 (N_3929,In_250,In_15);
nand U3930 (N_3930,In_622,In_859);
nor U3931 (N_3931,In_946,In_543);
xor U3932 (N_3932,In_656,In_811);
nand U3933 (N_3933,In_107,In_544);
and U3934 (N_3934,In_613,In_179);
or U3935 (N_3935,In_335,In_895);
nand U3936 (N_3936,In_983,In_280);
nor U3937 (N_3937,In_37,In_556);
xnor U3938 (N_3938,In_724,In_230);
and U3939 (N_3939,In_541,In_693);
and U3940 (N_3940,In_863,In_42);
and U3941 (N_3941,In_560,In_676);
xnor U3942 (N_3942,In_692,In_369);
nor U3943 (N_3943,In_247,In_927);
or U3944 (N_3944,In_110,In_469);
nand U3945 (N_3945,In_430,In_943);
nand U3946 (N_3946,In_745,In_172);
or U3947 (N_3947,In_323,In_215);
or U3948 (N_3948,In_464,In_363);
nor U3949 (N_3949,In_242,In_191);
and U3950 (N_3950,In_335,In_326);
or U3951 (N_3951,In_488,In_853);
or U3952 (N_3952,In_181,In_923);
nor U3953 (N_3953,In_847,In_555);
xnor U3954 (N_3954,In_632,In_971);
nand U3955 (N_3955,In_851,In_674);
and U3956 (N_3956,In_134,In_808);
and U3957 (N_3957,In_995,In_886);
or U3958 (N_3958,In_336,In_782);
nand U3959 (N_3959,In_362,In_998);
or U3960 (N_3960,In_370,In_192);
nor U3961 (N_3961,In_24,In_583);
nor U3962 (N_3962,In_525,In_919);
and U3963 (N_3963,In_568,In_660);
and U3964 (N_3964,In_203,In_215);
xor U3965 (N_3965,In_668,In_507);
and U3966 (N_3966,In_404,In_338);
and U3967 (N_3967,In_245,In_745);
nand U3968 (N_3968,In_845,In_388);
or U3969 (N_3969,In_302,In_901);
and U3970 (N_3970,In_903,In_390);
or U3971 (N_3971,In_580,In_490);
nand U3972 (N_3972,In_143,In_52);
nor U3973 (N_3973,In_577,In_105);
or U3974 (N_3974,In_996,In_467);
xor U3975 (N_3975,In_62,In_212);
nand U3976 (N_3976,In_840,In_949);
nand U3977 (N_3977,In_861,In_77);
nand U3978 (N_3978,In_5,In_263);
or U3979 (N_3979,In_660,In_411);
or U3980 (N_3980,In_659,In_200);
nand U3981 (N_3981,In_270,In_716);
xor U3982 (N_3982,In_810,In_806);
or U3983 (N_3983,In_820,In_707);
nand U3984 (N_3984,In_55,In_852);
or U3985 (N_3985,In_924,In_42);
or U3986 (N_3986,In_173,In_734);
or U3987 (N_3987,In_517,In_145);
xnor U3988 (N_3988,In_731,In_502);
and U3989 (N_3989,In_347,In_574);
nor U3990 (N_3990,In_806,In_191);
xnor U3991 (N_3991,In_344,In_663);
nand U3992 (N_3992,In_227,In_945);
nor U3993 (N_3993,In_413,In_877);
and U3994 (N_3994,In_303,In_377);
or U3995 (N_3995,In_968,In_33);
and U3996 (N_3996,In_933,In_848);
nand U3997 (N_3997,In_494,In_828);
nor U3998 (N_3998,In_841,In_260);
nand U3999 (N_3999,In_935,In_384);
xor U4000 (N_4000,In_20,In_747);
xnor U4001 (N_4001,In_665,In_525);
nor U4002 (N_4002,In_277,In_825);
or U4003 (N_4003,In_188,In_300);
and U4004 (N_4004,In_186,In_125);
nand U4005 (N_4005,In_198,In_771);
nor U4006 (N_4006,In_110,In_845);
or U4007 (N_4007,In_511,In_316);
nor U4008 (N_4008,In_13,In_270);
and U4009 (N_4009,In_92,In_30);
nand U4010 (N_4010,In_49,In_914);
or U4011 (N_4011,In_699,In_558);
nand U4012 (N_4012,In_962,In_242);
and U4013 (N_4013,In_658,In_412);
and U4014 (N_4014,In_817,In_992);
nor U4015 (N_4015,In_107,In_695);
nor U4016 (N_4016,In_758,In_599);
or U4017 (N_4017,In_472,In_809);
nand U4018 (N_4018,In_886,In_882);
nand U4019 (N_4019,In_850,In_534);
or U4020 (N_4020,In_319,In_986);
or U4021 (N_4021,In_383,In_441);
xor U4022 (N_4022,In_879,In_713);
nor U4023 (N_4023,In_727,In_691);
or U4024 (N_4024,In_717,In_577);
nor U4025 (N_4025,In_253,In_618);
or U4026 (N_4026,In_643,In_459);
nor U4027 (N_4027,In_381,In_553);
and U4028 (N_4028,In_58,In_228);
nor U4029 (N_4029,In_304,In_992);
or U4030 (N_4030,In_872,In_839);
nand U4031 (N_4031,In_55,In_309);
nand U4032 (N_4032,In_336,In_996);
nand U4033 (N_4033,In_298,In_684);
and U4034 (N_4034,In_787,In_43);
xnor U4035 (N_4035,In_816,In_215);
xor U4036 (N_4036,In_423,In_349);
nand U4037 (N_4037,In_858,In_380);
xor U4038 (N_4038,In_860,In_967);
nor U4039 (N_4039,In_885,In_711);
or U4040 (N_4040,In_610,In_477);
nor U4041 (N_4041,In_396,In_460);
nor U4042 (N_4042,In_281,In_709);
or U4043 (N_4043,In_981,In_119);
and U4044 (N_4044,In_805,In_367);
nand U4045 (N_4045,In_935,In_727);
nand U4046 (N_4046,In_157,In_9);
nor U4047 (N_4047,In_401,In_373);
and U4048 (N_4048,In_244,In_308);
or U4049 (N_4049,In_997,In_968);
and U4050 (N_4050,In_637,In_392);
nor U4051 (N_4051,In_13,In_878);
or U4052 (N_4052,In_239,In_934);
xnor U4053 (N_4053,In_27,In_314);
and U4054 (N_4054,In_192,In_85);
and U4055 (N_4055,In_700,In_358);
nor U4056 (N_4056,In_599,In_835);
nor U4057 (N_4057,In_448,In_812);
nor U4058 (N_4058,In_826,In_150);
nor U4059 (N_4059,In_989,In_285);
nand U4060 (N_4060,In_918,In_869);
nor U4061 (N_4061,In_604,In_329);
nor U4062 (N_4062,In_576,In_274);
or U4063 (N_4063,In_304,In_312);
or U4064 (N_4064,In_903,In_157);
and U4065 (N_4065,In_705,In_296);
or U4066 (N_4066,In_396,In_652);
or U4067 (N_4067,In_632,In_581);
nand U4068 (N_4068,In_300,In_200);
nand U4069 (N_4069,In_340,In_261);
and U4070 (N_4070,In_391,In_807);
or U4071 (N_4071,In_246,In_262);
and U4072 (N_4072,In_146,In_239);
and U4073 (N_4073,In_502,In_779);
xnor U4074 (N_4074,In_16,In_533);
or U4075 (N_4075,In_775,In_27);
nand U4076 (N_4076,In_789,In_655);
and U4077 (N_4077,In_715,In_83);
nor U4078 (N_4078,In_746,In_806);
and U4079 (N_4079,In_308,In_458);
nor U4080 (N_4080,In_862,In_707);
xnor U4081 (N_4081,In_690,In_196);
nor U4082 (N_4082,In_728,In_419);
and U4083 (N_4083,In_587,In_954);
nor U4084 (N_4084,In_134,In_972);
and U4085 (N_4085,In_114,In_925);
nor U4086 (N_4086,In_658,In_953);
xor U4087 (N_4087,In_809,In_446);
xor U4088 (N_4088,In_200,In_796);
nor U4089 (N_4089,In_411,In_645);
or U4090 (N_4090,In_607,In_67);
or U4091 (N_4091,In_64,In_22);
and U4092 (N_4092,In_446,In_584);
or U4093 (N_4093,In_599,In_271);
and U4094 (N_4094,In_445,In_930);
nor U4095 (N_4095,In_403,In_645);
nand U4096 (N_4096,In_792,In_859);
and U4097 (N_4097,In_964,In_499);
nand U4098 (N_4098,In_638,In_875);
nor U4099 (N_4099,In_431,In_864);
and U4100 (N_4100,In_82,In_996);
nor U4101 (N_4101,In_599,In_759);
nand U4102 (N_4102,In_677,In_343);
and U4103 (N_4103,In_671,In_935);
and U4104 (N_4104,In_462,In_632);
nand U4105 (N_4105,In_295,In_274);
nand U4106 (N_4106,In_351,In_269);
nand U4107 (N_4107,In_642,In_637);
nor U4108 (N_4108,In_21,In_176);
or U4109 (N_4109,In_580,In_182);
and U4110 (N_4110,In_111,In_201);
and U4111 (N_4111,In_724,In_923);
nor U4112 (N_4112,In_847,In_523);
or U4113 (N_4113,In_640,In_317);
or U4114 (N_4114,In_33,In_40);
or U4115 (N_4115,In_862,In_940);
and U4116 (N_4116,In_369,In_759);
nand U4117 (N_4117,In_749,In_173);
nor U4118 (N_4118,In_621,In_147);
and U4119 (N_4119,In_869,In_339);
and U4120 (N_4120,In_685,In_9);
xnor U4121 (N_4121,In_644,In_673);
or U4122 (N_4122,In_457,In_886);
nor U4123 (N_4123,In_267,In_571);
nor U4124 (N_4124,In_866,In_117);
nor U4125 (N_4125,In_288,In_898);
nand U4126 (N_4126,In_774,In_40);
and U4127 (N_4127,In_338,In_385);
or U4128 (N_4128,In_516,In_559);
nor U4129 (N_4129,In_50,In_334);
nor U4130 (N_4130,In_919,In_853);
and U4131 (N_4131,In_751,In_588);
or U4132 (N_4132,In_858,In_418);
nand U4133 (N_4133,In_332,In_713);
and U4134 (N_4134,In_584,In_36);
nor U4135 (N_4135,In_831,In_623);
nor U4136 (N_4136,In_557,In_314);
nor U4137 (N_4137,In_873,In_316);
or U4138 (N_4138,In_679,In_353);
or U4139 (N_4139,In_311,In_334);
or U4140 (N_4140,In_706,In_564);
and U4141 (N_4141,In_260,In_903);
and U4142 (N_4142,In_732,In_846);
or U4143 (N_4143,In_829,In_850);
nand U4144 (N_4144,In_882,In_831);
nand U4145 (N_4145,In_93,In_345);
xnor U4146 (N_4146,In_232,In_662);
nand U4147 (N_4147,In_124,In_93);
or U4148 (N_4148,In_405,In_886);
or U4149 (N_4149,In_27,In_583);
nand U4150 (N_4150,In_607,In_539);
and U4151 (N_4151,In_308,In_935);
or U4152 (N_4152,In_508,In_833);
or U4153 (N_4153,In_388,In_550);
and U4154 (N_4154,In_715,In_565);
and U4155 (N_4155,In_233,In_540);
nand U4156 (N_4156,In_583,In_870);
nor U4157 (N_4157,In_154,In_932);
nor U4158 (N_4158,In_265,In_475);
and U4159 (N_4159,In_469,In_126);
or U4160 (N_4160,In_178,In_489);
nand U4161 (N_4161,In_935,In_403);
nand U4162 (N_4162,In_259,In_257);
xor U4163 (N_4163,In_664,In_960);
nand U4164 (N_4164,In_596,In_861);
or U4165 (N_4165,In_989,In_232);
and U4166 (N_4166,In_328,In_426);
and U4167 (N_4167,In_828,In_570);
or U4168 (N_4168,In_564,In_68);
or U4169 (N_4169,In_482,In_324);
nand U4170 (N_4170,In_341,In_843);
nand U4171 (N_4171,In_152,In_878);
or U4172 (N_4172,In_979,In_881);
or U4173 (N_4173,In_829,In_965);
and U4174 (N_4174,In_481,In_157);
and U4175 (N_4175,In_445,In_515);
or U4176 (N_4176,In_561,In_496);
or U4177 (N_4177,In_689,In_989);
or U4178 (N_4178,In_627,In_301);
or U4179 (N_4179,In_385,In_373);
xnor U4180 (N_4180,In_8,In_195);
nor U4181 (N_4181,In_338,In_439);
nand U4182 (N_4182,In_836,In_59);
or U4183 (N_4183,In_866,In_721);
or U4184 (N_4184,In_215,In_805);
and U4185 (N_4185,In_453,In_986);
and U4186 (N_4186,In_396,In_380);
and U4187 (N_4187,In_867,In_37);
and U4188 (N_4188,In_116,In_819);
nor U4189 (N_4189,In_96,In_452);
or U4190 (N_4190,In_43,In_765);
or U4191 (N_4191,In_831,In_936);
nand U4192 (N_4192,In_451,In_830);
or U4193 (N_4193,In_95,In_34);
or U4194 (N_4194,In_961,In_783);
or U4195 (N_4195,In_893,In_498);
nand U4196 (N_4196,In_382,In_325);
and U4197 (N_4197,In_251,In_214);
nor U4198 (N_4198,In_757,In_786);
or U4199 (N_4199,In_474,In_868);
and U4200 (N_4200,In_487,In_715);
or U4201 (N_4201,In_638,In_132);
or U4202 (N_4202,In_677,In_728);
nand U4203 (N_4203,In_545,In_648);
and U4204 (N_4204,In_605,In_957);
nand U4205 (N_4205,In_890,In_957);
nand U4206 (N_4206,In_542,In_783);
and U4207 (N_4207,In_578,In_576);
or U4208 (N_4208,In_335,In_163);
or U4209 (N_4209,In_525,In_358);
or U4210 (N_4210,In_768,In_490);
and U4211 (N_4211,In_394,In_56);
nand U4212 (N_4212,In_764,In_229);
nand U4213 (N_4213,In_628,In_498);
nand U4214 (N_4214,In_56,In_632);
and U4215 (N_4215,In_65,In_171);
nor U4216 (N_4216,In_587,In_882);
nor U4217 (N_4217,In_638,In_700);
nor U4218 (N_4218,In_769,In_114);
nor U4219 (N_4219,In_859,In_756);
nor U4220 (N_4220,In_58,In_171);
and U4221 (N_4221,In_926,In_773);
and U4222 (N_4222,In_536,In_415);
and U4223 (N_4223,In_238,In_271);
nand U4224 (N_4224,In_12,In_524);
nand U4225 (N_4225,In_901,In_961);
or U4226 (N_4226,In_470,In_206);
and U4227 (N_4227,In_331,In_124);
nor U4228 (N_4228,In_722,In_315);
and U4229 (N_4229,In_603,In_804);
nand U4230 (N_4230,In_150,In_258);
nor U4231 (N_4231,In_665,In_500);
or U4232 (N_4232,In_463,In_120);
nand U4233 (N_4233,In_124,In_89);
nor U4234 (N_4234,In_940,In_646);
nand U4235 (N_4235,In_214,In_526);
nor U4236 (N_4236,In_977,In_497);
or U4237 (N_4237,In_64,In_683);
or U4238 (N_4238,In_313,In_78);
nand U4239 (N_4239,In_177,In_665);
xnor U4240 (N_4240,In_884,In_983);
xor U4241 (N_4241,In_185,In_653);
nor U4242 (N_4242,In_277,In_424);
nor U4243 (N_4243,In_829,In_757);
xnor U4244 (N_4244,In_351,In_116);
or U4245 (N_4245,In_584,In_891);
or U4246 (N_4246,In_463,In_365);
or U4247 (N_4247,In_376,In_38);
xor U4248 (N_4248,In_165,In_683);
nand U4249 (N_4249,In_404,In_750);
nand U4250 (N_4250,In_655,In_450);
and U4251 (N_4251,In_18,In_208);
and U4252 (N_4252,In_856,In_413);
nor U4253 (N_4253,In_159,In_208);
or U4254 (N_4254,In_689,In_186);
and U4255 (N_4255,In_599,In_365);
or U4256 (N_4256,In_477,In_310);
or U4257 (N_4257,In_673,In_350);
or U4258 (N_4258,In_127,In_536);
and U4259 (N_4259,In_999,In_187);
and U4260 (N_4260,In_450,In_745);
nor U4261 (N_4261,In_784,In_110);
nand U4262 (N_4262,In_26,In_265);
or U4263 (N_4263,In_867,In_869);
nor U4264 (N_4264,In_406,In_627);
nor U4265 (N_4265,In_459,In_811);
and U4266 (N_4266,In_261,In_68);
nor U4267 (N_4267,In_784,In_681);
or U4268 (N_4268,In_384,In_32);
nor U4269 (N_4269,In_54,In_438);
nor U4270 (N_4270,In_383,In_195);
or U4271 (N_4271,In_246,In_417);
or U4272 (N_4272,In_95,In_929);
and U4273 (N_4273,In_303,In_587);
and U4274 (N_4274,In_450,In_638);
nor U4275 (N_4275,In_339,In_305);
nor U4276 (N_4276,In_551,In_858);
nor U4277 (N_4277,In_324,In_550);
and U4278 (N_4278,In_504,In_402);
nand U4279 (N_4279,In_698,In_819);
or U4280 (N_4280,In_857,In_119);
or U4281 (N_4281,In_429,In_687);
and U4282 (N_4282,In_313,In_153);
or U4283 (N_4283,In_72,In_963);
nand U4284 (N_4284,In_41,In_634);
nand U4285 (N_4285,In_888,In_800);
nand U4286 (N_4286,In_440,In_772);
nand U4287 (N_4287,In_562,In_500);
or U4288 (N_4288,In_822,In_423);
xnor U4289 (N_4289,In_207,In_407);
or U4290 (N_4290,In_381,In_406);
nand U4291 (N_4291,In_367,In_113);
or U4292 (N_4292,In_29,In_238);
and U4293 (N_4293,In_25,In_481);
and U4294 (N_4294,In_597,In_61);
or U4295 (N_4295,In_321,In_220);
or U4296 (N_4296,In_77,In_822);
and U4297 (N_4297,In_245,In_661);
or U4298 (N_4298,In_405,In_762);
or U4299 (N_4299,In_723,In_692);
or U4300 (N_4300,In_722,In_497);
nor U4301 (N_4301,In_728,In_57);
nor U4302 (N_4302,In_119,In_691);
and U4303 (N_4303,In_188,In_908);
and U4304 (N_4304,In_983,In_913);
and U4305 (N_4305,In_166,In_879);
and U4306 (N_4306,In_647,In_247);
xor U4307 (N_4307,In_619,In_636);
xor U4308 (N_4308,In_679,In_629);
nor U4309 (N_4309,In_805,In_919);
nor U4310 (N_4310,In_764,In_608);
or U4311 (N_4311,In_484,In_920);
nor U4312 (N_4312,In_996,In_759);
nor U4313 (N_4313,In_229,In_183);
nand U4314 (N_4314,In_882,In_163);
or U4315 (N_4315,In_232,In_262);
xor U4316 (N_4316,In_544,In_44);
and U4317 (N_4317,In_74,In_800);
nor U4318 (N_4318,In_11,In_332);
nand U4319 (N_4319,In_831,In_333);
nor U4320 (N_4320,In_632,In_359);
and U4321 (N_4321,In_560,In_345);
nor U4322 (N_4322,In_973,In_261);
and U4323 (N_4323,In_427,In_638);
nor U4324 (N_4324,In_327,In_36);
nand U4325 (N_4325,In_455,In_387);
or U4326 (N_4326,In_633,In_852);
nor U4327 (N_4327,In_67,In_473);
or U4328 (N_4328,In_308,In_32);
and U4329 (N_4329,In_167,In_766);
xnor U4330 (N_4330,In_136,In_811);
xor U4331 (N_4331,In_900,In_266);
or U4332 (N_4332,In_117,In_694);
nand U4333 (N_4333,In_52,In_80);
and U4334 (N_4334,In_158,In_92);
nand U4335 (N_4335,In_213,In_442);
or U4336 (N_4336,In_291,In_420);
nand U4337 (N_4337,In_233,In_45);
nand U4338 (N_4338,In_517,In_692);
or U4339 (N_4339,In_275,In_550);
xnor U4340 (N_4340,In_589,In_274);
and U4341 (N_4341,In_832,In_272);
nand U4342 (N_4342,In_610,In_226);
and U4343 (N_4343,In_384,In_569);
and U4344 (N_4344,In_451,In_207);
and U4345 (N_4345,In_361,In_767);
nand U4346 (N_4346,In_654,In_945);
nor U4347 (N_4347,In_354,In_270);
or U4348 (N_4348,In_220,In_336);
xnor U4349 (N_4349,In_602,In_731);
nand U4350 (N_4350,In_333,In_336);
nor U4351 (N_4351,In_863,In_590);
or U4352 (N_4352,In_652,In_490);
nand U4353 (N_4353,In_717,In_422);
nor U4354 (N_4354,In_393,In_581);
nor U4355 (N_4355,In_322,In_419);
nor U4356 (N_4356,In_587,In_341);
or U4357 (N_4357,In_943,In_314);
nor U4358 (N_4358,In_565,In_783);
nand U4359 (N_4359,In_205,In_939);
xnor U4360 (N_4360,In_54,In_829);
nand U4361 (N_4361,In_321,In_398);
nand U4362 (N_4362,In_19,In_98);
or U4363 (N_4363,In_174,In_974);
xor U4364 (N_4364,In_872,In_772);
and U4365 (N_4365,In_596,In_710);
and U4366 (N_4366,In_982,In_170);
nand U4367 (N_4367,In_427,In_48);
or U4368 (N_4368,In_610,In_9);
xnor U4369 (N_4369,In_148,In_187);
nand U4370 (N_4370,In_251,In_572);
and U4371 (N_4371,In_956,In_896);
and U4372 (N_4372,In_94,In_471);
or U4373 (N_4373,In_456,In_294);
nand U4374 (N_4374,In_104,In_19);
nor U4375 (N_4375,In_902,In_981);
or U4376 (N_4376,In_460,In_1);
and U4377 (N_4377,In_201,In_910);
and U4378 (N_4378,In_46,In_977);
nand U4379 (N_4379,In_218,In_516);
nand U4380 (N_4380,In_927,In_216);
or U4381 (N_4381,In_769,In_130);
or U4382 (N_4382,In_546,In_697);
or U4383 (N_4383,In_771,In_178);
or U4384 (N_4384,In_497,In_845);
and U4385 (N_4385,In_216,In_830);
xnor U4386 (N_4386,In_220,In_233);
nand U4387 (N_4387,In_959,In_541);
or U4388 (N_4388,In_739,In_913);
nand U4389 (N_4389,In_202,In_949);
nand U4390 (N_4390,In_381,In_499);
nor U4391 (N_4391,In_17,In_878);
or U4392 (N_4392,In_944,In_744);
or U4393 (N_4393,In_979,In_963);
and U4394 (N_4394,In_919,In_79);
or U4395 (N_4395,In_18,In_953);
nor U4396 (N_4396,In_986,In_458);
and U4397 (N_4397,In_866,In_528);
and U4398 (N_4398,In_489,In_597);
nand U4399 (N_4399,In_467,In_596);
xnor U4400 (N_4400,In_449,In_662);
nor U4401 (N_4401,In_669,In_725);
nor U4402 (N_4402,In_899,In_944);
nor U4403 (N_4403,In_966,In_893);
or U4404 (N_4404,In_728,In_494);
nor U4405 (N_4405,In_936,In_309);
and U4406 (N_4406,In_257,In_332);
nand U4407 (N_4407,In_760,In_963);
nand U4408 (N_4408,In_44,In_549);
nand U4409 (N_4409,In_713,In_327);
nand U4410 (N_4410,In_927,In_190);
nand U4411 (N_4411,In_611,In_110);
nor U4412 (N_4412,In_591,In_663);
nand U4413 (N_4413,In_413,In_625);
nand U4414 (N_4414,In_127,In_177);
or U4415 (N_4415,In_30,In_629);
or U4416 (N_4416,In_490,In_696);
nor U4417 (N_4417,In_727,In_53);
or U4418 (N_4418,In_18,In_363);
nor U4419 (N_4419,In_681,In_553);
and U4420 (N_4420,In_69,In_663);
and U4421 (N_4421,In_148,In_585);
nand U4422 (N_4422,In_689,In_695);
or U4423 (N_4423,In_139,In_121);
nand U4424 (N_4424,In_478,In_384);
nor U4425 (N_4425,In_870,In_169);
and U4426 (N_4426,In_527,In_319);
xnor U4427 (N_4427,In_262,In_629);
or U4428 (N_4428,In_937,In_943);
and U4429 (N_4429,In_512,In_58);
nand U4430 (N_4430,In_397,In_820);
and U4431 (N_4431,In_169,In_438);
nand U4432 (N_4432,In_874,In_423);
and U4433 (N_4433,In_801,In_78);
or U4434 (N_4434,In_141,In_23);
and U4435 (N_4435,In_111,In_652);
or U4436 (N_4436,In_817,In_250);
xnor U4437 (N_4437,In_447,In_46);
nand U4438 (N_4438,In_312,In_791);
nor U4439 (N_4439,In_113,In_52);
and U4440 (N_4440,In_951,In_396);
and U4441 (N_4441,In_698,In_586);
nor U4442 (N_4442,In_124,In_817);
nor U4443 (N_4443,In_808,In_621);
and U4444 (N_4444,In_341,In_412);
nor U4445 (N_4445,In_776,In_452);
nand U4446 (N_4446,In_367,In_771);
or U4447 (N_4447,In_226,In_624);
or U4448 (N_4448,In_574,In_685);
or U4449 (N_4449,In_531,In_203);
xor U4450 (N_4450,In_24,In_407);
and U4451 (N_4451,In_455,In_746);
xor U4452 (N_4452,In_657,In_988);
xnor U4453 (N_4453,In_33,In_812);
and U4454 (N_4454,In_163,In_348);
nor U4455 (N_4455,In_751,In_884);
or U4456 (N_4456,In_70,In_973);
xnor U4457 (N_4457,In_400,In_14);
or U4458 (N_4458,In_808,In_704);
nand U4459 (N_4459,In_361,In_377);
nand U4460 (N_4460,In_599,In_112);
xor U4461 (N_4461,In_260,In_213);
nor U4462 (N_4462,In_299,In_30);
or U4463 (N_4463,In_127,In_45);
and U4464 (N_4464,In_706,In_89);
nand U4465 (N_4465,In_958,In_269);
and U4466 (N_4466,In_353,In_682);
or U4467 (N_4467,In_84,In_586);
nand U4468 (N_4468,In_347,In_241);
xor U4469 (N_4469,In_245,In_914);
nor U4470 (N_4470,In_337,In_610);
and U4471 (N_4471,In_222,In_75);
or U4472 (N_4472,In_812,In_128);
nand U4473 (N_4473,In_516,In_951);
nor U4474 (N_4474,In_214,In_512);
or U4475 (N_4475,In_893,In_969);
nor U4476 (N_4476,In_690,In_62);
nand U4477 (N_4477,In_740,In_571);
or U4478 (N_4478,In_87,In_320);
nand U4479 (N_4479,In_142,In_22);
nand U4480 (N_4480,In_71,In_92);
nand U4481 (N_4481,In_957,In_34);
xnor U4482 (N_4482,In_149,In_653);
nor U4483 (N_4483,In_921,In_708);
xor U4484 (N_4484,In_340,In_579);
or U4485 (N_4485,In_458,In_330);
nor U4486 (N_4486,In_678,In_218);
xnor U4487 (N_4487,In_307,In_104);
nand U4488 (N_4488,In_525,In_442);
nand U4489 (N_4489,In_839,In_873);
nor U4490 (N_4490,In_944,In_333);
or U4491 (N_4491,In_789,In_692);
nand U4492 (N_4492,In_89,In_137);
xor U4493 (N_4493,In_950,In_653);
or U4494 (N_4494,In_254,In_28);
or U4495 (N_4495,In_926,In_30);
or U4496 (N_4496,In_223,In_238);
and U4497 (N_4497,In_615,In_55);
or U4498 (N_4498,In_85,In_820);
nor U4499 (N_4499,In_534,In_616);
xnor U4500 (N_4500,In_338,In_656);
or U4501 (N_4501,In_465,In_652);
and U4502 (N_4502,In_349,In_276);
nand U4503 (N_4503,In_814,In_906);
nor U4504 (N_4504,In_425,In_269);
and U4505 (N_4505,In_120,In_614);
or U4506 (N_4506,In_667,In_418);
or U4507 (N_4507,In_577,In_282);
nor U4508 (N_4508,In_860,In_777);
nor U4509 (N_4509,In_212,In_64);
or U4510 (N_4510,In_300,In_747);
and U4511 (N_4511,In_657,In_226);
nor U4512 (N_4512,In_729,In_150);
or U4513 (N_4513,In_946,In_425);
or U4514 (N_4514,In_927,In_573);
nand U4515 (N_4515,In_758,In_329);
xor U4516 (N_4516,In_589,In_364);
and U4517 (N_4517,In_435,In_644);
xor U4518 (N_4518,In_795,In_983);
and U4519 (N_4519,In_522,In_354);
and U4520 (N_4520,In_594,In_861);
nor U4521 (N_4521,In_345,In_738);
nor U4522 (N_4522,In_459,In_395);
or U4523 (N_4523,In_167,In_184);
or U4524 (N_4524,In_69,In_851);
nand U4525 (N_4525,In_601,In_185);
nand U4526 (N_4526,In_716,In_911);
or U4527 (N_4527,In_104,In_701);
nor U4528 (N_4528,In_24,In_224);
or U4529 (N_4529,In_502,In_202);
nand U4530 (N_4530,In_254,In_163);
nand U4531 (N_4531,In_273,In_495);
or U4532 (N_4532,In_219,In_529);
and U4533 (N_4533,In_270,In_670);
and U4534 (N_4534,In_10,In_888);
xor U4535 (N_4535,In_148,In_691);
and U4536 (N_4536,In_77,In_882);
or U4537 (N_4537,In_514,In_616);
or U4538 (N_4538,In_247,In_153);
nor U4539 (N_4539,In_68,In_483);
or U4540 (N_4540,In_414,In_104);
nor U4541 (N_4541,In_418,In_488);
nor U4542 (N_4542,In_965,In_418);
or U4543 (N_4543,In_736,In_135);
nand U4544 (N_4544,In_63,In_841);
nand U4545 (N_4545,In_472,In_984);
or U4546 (N_4546,In_455,In_331);
nor U4547 (N_4547,In_711,In_285);
xnor U4548 (N_4548,In_943,In_381);
and U4549 (N_4549,In_619,In_879);
nand U4550 (N_4550,In_777,In_468);
nor U4551 (N_4551,In_474,In_747);
nor U4552 (N_4552,In_3,In_133);
nor U4553 (N_4553,In_260,In_608);
nor U4554 (N_4554,In_323,In_227);
nand U4555 (N_4555,In_295,In_38);
nor U4556 (N_4556,In_655,In_750);
nor U4557 (N_4557,In_788,In_629);
or U4558 (N_4558,In_41,In_586);
nor U4559 (N_4559,In_585,In_231);
or U4560 (N_4560,In_529,In_232);
nor U4561 (N_4561,In_319,In_362);
or U4562 (N_4562,In_192,In_933);
nor U4563 (N_4563,In_984,In_593);
and U4564 (N_4564,In_912,In_809);
nand U4565 (N_4565,In_6,In_761);
nand U4566 (N_4566,In_360,In_175);
and U4567 (N_4567,In_945,In_64);
nand U4568 (N_4568,In_598,In_286);
xnor U4569 (N_4569,In_833,In_577);
nor U4570 (N_4570,In_430,In_440);
or U4571 (N_4571,In_127,In_636);
nand U4572 (N_4572,In_505,In_595);
nand U4573 (N_4573,In_385,In_139);
or U4574 (N_4574,In_752,In_717);
or U4575 (N_4575,In_88,In_81);
xnor U4576 (N_4576,In_938,In_429);
and U4577 (N_4577,In_510,In_608);
xnor U4578 (N_4578,In_896,In_167);
nor U4579 (N_4579,In_895,In_265);
or U4580 (N_4580,In_904,In_383);
and U4581 (N_4581,In_690,In_397);
nor U4582 (N_4582,In_417,In_858);
nor U4583 (N_4583,In_58,In_284);
or U4584 (N_4584,In_696,In_484);
nor U4585 (N_4585,In_978,In_749);
or U4586 (N_4586,In_299,In_438);
nand U4587 (N_4587,In_240,In_634);
nand U4588 (N_4588,In_893,In_876);
and U4589 (N_4589,In_484,In_471);
or U4590 (N_4590,In_597,In_912);
nand U4591 (N_4591,In_814,In_838);
nand U4592 (N_4592,In_488,In_763);
or U4593 (N_4593,In_779,In_734);
nor U4594 (N_4594,In_397,In_481);
nand U4595 (N_4595,In_362,In_639);
nand U4596 (N_4596,In_565,In_503);
and U4597 (N_4597,In_655,In_588);
and U4598 (N_4598,In_829,In_980);
xnor U4599 (N_4599,In_799,In_63);
nand U4600 (N_4600,In_939,In_369);
and U4601 (N_4601,In_421,In_707);
and U4602 (N_4602,In_432,In_781);
or U4603 (N_4603,In_291,In_764);
and U4604 (N_4604,In_275,In_612);
or U4605 (N_4605,In_172,In_593);
or U4606 (N_4606,In_861,In_17);
nor U4607 (N_4607,In_794,In_795);
nor U4608 (N_4608,In_330,In_375);
nand U4609 (N_4609,In_547,In_459);
nand U4610 (N_4610,In_781,In_614);
or U4611 (N_4611,In_243,In_291);
nor U4612 (N_4612,In_465,In_412);
nand U4613 (N_4613,In_500,In_913);
or U4614 (N_4614,In_795,In_113);
and U4615 (N_4615,In_186,In_260);
nand U4616 (N_4616,In_230,In_132);
nand U4617 (N_4617,In_649,In_641);
xnor U4618 (N_4618,In_573,In_727);
nand U4619 (N_4619,In_353,In_793);
and U4620 (N_4620,In_576,In_998);
and U4621 (N_4621,In_540,In_223);
nand U4622 (N_4622,In_800,In_418);
and U4623 (N_4623,In_593,In_96);
or U4624 (N_4624,In_411,In_682);
xor U4625 (N_4625,In_793,In_592);
nand U4626 (N_4626,In_273,In_537);
nand U4627 (N_4627,In_786,In_634);
nand U4628 (N_4628,In_158,In_861);
xor U4629 (N_4629,In_299,In_420);
nand U4630 (N_4630,In_455,In_69);
nor U4631 (N_4631,In_16,In_587);
nor U4632 (N_4632,In_365,In_79);
or U4633 (N_4633,In_738,In_25);
nand U4634 (N_4634,In_539,In_257);
or U4635 (N_4635,In_567,In_380);
nor U4636 (N_4636,In_249,In_311);
nor U4637 (N_4637,In_623,In_475);
xor U4638 (N_4638,In_986,In_709);
nand U4639 (N_4639,In_722,In_744);
nor U4640 (N_4640,In_637,In_482);
or U4641 (N_4641,In_869,In_118);
nand U4642 (N_4642,In_218,In_390);
nand U4643 (N_4643,In_61,In_783);
or U4644 (N_4644,In_830,In_921);
and U4645 (N_4645,In_512,In_648);
nor U4646 (N_4646,In_8,In_283);
nor U4647 (N_4647,In_583,In_814);
or U4648 (N_4648,In_242,In_996);
nand U4649 (N_4649,In_722,In_469);
nand U4650 (N_4650,In_510,In_428);
nor U4651 (N_4651,In_749,In_158);
nor U4652 (N_4652,In_858,In_446);
and U4653 (N_4653,In_161,In_958);
nand U4654 (N_4654,In_745,In_287);
and U4655 (N_4655,In_179,In_483);
and U4656 (N_4656,In_703,In_276);
and U4657 (N_4657,In_67,In_35);
nand U4658 (N_4658,In_251,In_380);
or U4659 (N_4659,In_819,In_589);
and U4660 (N_4660,In_665,In_178);
nor U4661 (N_4661,In_146,In_150);
and U4662 (N_4662,In_493,In_267);
nand U4663 (N_4663,In_163,In_684);
and U4664 (N_4664,In_657,In_624);
and U4665 (N_4665,In_758,In_474);
nor U4666 (N_4666,In_163,In_502);
nand U4667 (N_4667,In_533,In_406);
nand U4668 (N_4668,In_397,In_612);
nor U4669 (N_4669,In_320,In_339);
nand U4670 (N_4670,In_808,In_166);
xor U4671 (N_4671,In_934,In_303);
or U4672 (N_4672,In_964,In_98);
and U4673 (N_4673,In_385,In_31);
or U4674 (N_4674,In_680,In_667);
xor U4675 (N_4675,In_840,In_675);
and U4676 (N_4676,In_153,In_107);
and U4677 (N_4677,In_173,In_754);
nand U4678 (N_4678,In_568,In_391);
and U4679 (N_4679,In_717,In_656);
nand U4680 (N_4680,In_107,In_559);
xnor U4681 (N_4681,In_740,In_791);
or U4682 (N_4682,In_203,In_526);
nor U4683 (N_4683,In_494,In_772);
or U4684 (N_4684,In_889,In_497);
or U4685 (N_4685,In_731,In_373);
or U4686 (N_4686,In_712,In_197);
nor U4687 (N_4687,In_168,In_153);
and U4688 (N_4688,In_287,In_176);
and U4689 (N_4689,In_476,In_557);
nand U4690 (N_4690,In_482,In_790);
and U4691 (N_4691,In_47,In_719);
nor U4692 (N_4692,In_714,In_333);
or U4693 (N_4693,In_49,In_590);
xnor U4694 (N_4694,In_353,In_739);
or U4695 (N_4695,In_92,In_414);
or U4696 (N_4696,In_165,In_928);
or U4697 (N_4697,In_490,In_882);
nor U4698 (N_4698,In_863,In_536);
or U4699 (N_4699,In_179,In_139);
xor U4700 (N_4700,In_504,In_939);
and U4701 (N_4701,In_812,In_214);
nand U4702 (N_4702,In_139,In_433);
nand U4703 (N_4703,In_950,In_962);
nor U4704 (N_4704,In_342,In_8);
or U4705 (N_4705,In_79,In_185);
or U4706 (N_4706,In_98,In_63);
xor U4707 (N_4707,In_276,In_430);
and U4708 (N_4708,In_179,In_877);
and U4709 (N_4709,In_331,In_645);
or U4710 (N_4710,In_185,In_313);
xnor U4711 (N_4711,In_206,In_358);
nor U4712 (N_4712,In_337,In_274);
nor U4713 (N_4713,In_892,In_359);
nand U4714 (N_4714,In_851,In_284);
nand U4715 (N_4715,In_548,In_959);
and U4716 (N_4716,In_226,In_906);
and U4717 (N_4717,In_311,In_888);
nand U4718 (N_4718,In_779,In_330);
and U4719 (N_4719,In_468,In_377);
xnor U4720 (N_4720,In_665,In_441);
and U4721 (N_4721,In_145,In_11);
and U4722 (N_4722,In_558,In_574);
or U4723 (N_4723,In_845,In_728);
nand U4724 (N_4724,In_136,In_930);
and U4725 (N_4725,In_72,In_775);
nor U4726 (N_4726,In_305,In_574);
and U4727 (N_4727,In_263,In_229);
nor U4728 (N_4728,In_391,In_286);
nor U4729 (N_4729,In_870,In_932);
nand U4730 (N_4730,In_289,In_296);
nor U4731 (N_4731,In_335,In_707);
nor U4732 (N_4732,In_273,In_681);
nand U4733 (N_4733,In_916,In_651);
or U4734 (N_4734,In_956,In_612);
nand U4735 (N_4735,In_382,In_945);
or U4736 (N_4736,In_845,In_803);
nand U4737 (N_4737,In_888,In_234);
and U4738 (N_4738,In_93,In_947);
and U4739 (N_4739,In_17,In_415);
nor U4740 (N_4740,In_569,In_362);
nand U4741 (N_4741,In_82,In_938);
and U4742 (N_4742,In_718,In_390);
or U4743 (N_4743,In_851,In_71);
and U4744 (N_4744,In_286,In_262);
and U4745 (N_4745,In_489,In_974);
nand U4746 (N_4746,In_544,In_758);
nor U4747 (N_4747,In_372,In_374);
xor U4748 (N_4748,In_22,In_179);
xnor U4749 (N_4749,In_974,In_816);
nor U4750 (N_4750,In_232,In_834);
xor U4751 (N_4751,In_922,In_373);
and U4752 (N_4752,In_351,In_496);
xor U4753 (N_4753,In_584,In_200);
nand U4754 (N_4754,In_676,In_756);
and U4755 (N_4755,In_39,In_633);
nor U4756 (N_4756,In_436,In_635);
or U4757 (N_4757,In_268,In_899);
nor U4758 (N_4758,In_725,In_814);
xnor U4759 (N_4759,In_986,In_476);
or U4760 (N_4760,In_0,In_214);
xor U4761 (N_4761,In_119,In_942);
nor U4762 (N_4762,In_242,In_431);
xor U4763 (N_4763,In_695,In_349);
and U4764 (N_4764,In_220,In_575);
nor U4765 (N_4765,In_523,In_542);
nand U4766 (N_4766,In_581,In_272);
and U4767 (N_4767,In_736,In_555);
nand U4768 (N_4768,In_243,In_264);
and U4769 (N_4769,In_156,In_120);
or U4770 (N_4770,In_237,In_287);
and U4771 (N_4771,In_291,In_501);
nand U4772 (N_4772,In_551,In_791);
and U4773 (N_4773,In_630,In_627);
or U4774 (N_4774,In_938,In_968);
or U4775 (N_4775,In_817,In_941);
and U4776 (N_4776,In_962,In_80);
and U4777 (N_4777,In_917,In_151);
xnor U4778 (N_4778,In_214,In_998);
nor U4779 (N_4779,In_763,In_852);
and U4780 (N_4780,In_600,In_674);
nand U4781 (N_4781,In_133,In_42);
nor U4782 (N_4782,In_699,In_192);
nor U4783 (N_4783,In_313,In_544);
xor U4784 (N_4784,In_804,In_143);
nand U4785 (N_4785,In_594,In_936);
nand U4786 (N_4786,In_217,In_941);
and U4787 (N_4787,In_526,In_311);
or U4788 (N_4788,In_249,In_262);
xnor U4789 (N_4789,In_90,In_906);
nor U4790 (N_4790,In_579,In_106);
or U4791 (N_4791,In_67,In_880);
nand U4792 (N_4792,In_708,In_661);
nand U4793 (N_4793,In_673,In_484);
or U4794 (N_4794,In_842,In_290);
and U4795 (N_4795,In_68,In_842);
or U4796 (N_4796,In_562,In_192);
nor U4797 (N_4797,In_733,In_442);
and U4798 (N_4798,In_76,In_253);
and U4799 (N_4799,In_71,In_326);
nand U4800 (N_4800,In_783,In_390);
and U4801 (N_4801,In_843,In_564);
or U4802 (N_4802,In_649,In_939);
or U4803 (N_4803,In_912,In_693);
xnor U4804 (N_4804,In_690,In_211);
and U4805 (N_4805,In_383,In_869);
nand U4806 (N_4806,In_416,In_415);
nor U4807 (N_4807,In_106,In_983);
nand U4808 (N_4808,In_611,In_605);
nand U4809 (N_4809,In_707,In_624);
xor U4810 (N_4810,In_882,In_815);
nor U4811 (N_4811,In_35,In_759);
and U4812 (N_4812,In_20,In_479);
xnor U4813 (N_4813,In_10,In_679);
nand U4814 (N_4814,In_358,In_659);
or U4815 (N_4815,In_989,In_193);
nor U4816 (N_4816,In_341,In_367);
xnor U4817 (N_4817,In_637,In_139);
or U4818 (N_4818,In_688,In_68);
and U4819 (N_4819,In_566,In_704);
or U4820 (N_4820,In_14,In_821);
or U4821 (N_4821,In_771,In_217);
or U4822 (N_4822,In_355,In_621);
nand U4823 (N_4823,In_704,In_54);
and U4824 (N_4824,In_894,In_842);
nand U4825 (N_4825,In_146,In_246);
and U4826 (N_4826,In_703,In_503);
or U4827 (N_4827,In_27,In_565);
xor U4828 (N_4828,In_793,In_608);
nand U4829 (N_4829,In_199,In_56);
xor U4830 (N_4830,In_88,In_51);
or U4831 (N_4831,In_663,In_961);
and U4832 (N_4832,In_229,In_420);
or U4833 (N_4833,In_168,In_90);
or U4834 (N_4834,In_17,In_991);
or U4835 (N_4835,In_723,In_25);
and U4836 (N_4836,In_532,In_340);
and U4837 (N_4837,In_430,In_298);
nand U4838 (N_4838,In_754,In_262);
xor U4839 (N_4839,In_785,In_465);
nand U4840 (N_4840,In_467,In_182);
xnor U4841 (N_4841,In_676,In_63);
nand U4842 (N_4842,In_288,In_700);
nor U4843 (N_4843,In_626,In_525);
xnor U4844 (N_4844,In_490,In_504);
and U4845 (N_4845,In_75,In_975);
nor U4846 (N_4846,In_270,In_689);
and U4847 (N_4847,In_340,In_624);
or U4848 (N_4848,In_412,In_834);
nor U4849 (N_4849,In_328,In_707);
xor U4850 (N_4850,In_726,In_396);
and U4851 (N_4851,In_88,In_90);
nand U4852 (N_4852,In_191,In_756);
and U4853 (N_4853,In_266,In_237);
or U4854 (N_4854,In_448,In_262);
and U4855 (N_4855,In_881,In_976);
nor U4856 (N_4856,In_528,In_768);
and U4857 (N_4857,In_206,In_98);
nor U4858 (N_4858,In_485,In_212);
nand U4859 (N_4859,In_469,In_268);
and U4860 (N_4860,In_555,In_152);
or U4861 (N_4861,In_126,In_905);
and U4862 (N_4862,In_132,In_253);
nand U4863 (N_4863,In_358,In_273);
or U4864 (N_4864,In_71,In_408);
and U4865 (N_4865,In_277,In_81);
and U4866 (N_4866,In_972,In_899);
nand U4867 (N_4867,In_877,In_137);
nor U4868 (N_4868,In_617,In_308);
nand U4869 (N_4869,In_736,In_548);
nor U4870 (N_4870,In_43,In_634);
or U4871 (N_4871,In_581,In_244);
nor U4872 (N_4872,In_595,In_521);
nand U4873 (N_4873,In_738,In_284);
or U4874 (N_4874,In_791,In_126);
and U4875 (N_4875,In_900,In_713);
nor U4876 (N_4876,In_225,In_707);
nand U4877 (N_4877,In_239,In_725);
nor U4878 (N_4878,In_876,In_985);
or U4879 (N_4879,In_870,In_536);
xnor U4880 (N_4880,In_857,In_580);
or U4881 (N_4881,In_213,In_829);
xor U4882 (N_4882,In_62,In_416);
nand U4883 (N_4883,In_929,In_429);
xor U4884 (N_4884,In_473,In_289);
nor U4885 (N_4885,In_142,In_399);
and U4886 (N_4886,In_298,In_526);
or U4887 (N_4887,In_610,In_440);
nor U4888 (N_4888,In_24,In_633);
and U4889 (N_4889,In_713,In_375);
nor U4890 (N_4890,In_224,In_592);
or U4891 (N_4891,In_938,In_279);
nand U4892 (N_4892,In_123,In_249);
and U4893 (N_4893,In_722,In_726);
nor U4894 (N_4894,In_166,In_180);
nor U4895 (N_4895,In_531,In_72);
and U4896 (N_4896,In_401,In_232);
xnor U4897 (N_4897,In_341,In_373);
or U4898 (N_4898,In_401,In_414);
or U4899 (N_4899,In_433,In_674);
or U4900 (N_4900,In_377,In_524);
or U4901 (N_4901,In_722,In_932);
xnor U4902 (N_4902,In_108,In_24);
nand U4903 (N_4903,In_701,In_806);
xor U4904 (N_4904,In_901,In_456);
nor U4905 (N_4905,In_804,In_120);
nor U4906 (N_4906,In_80,In_68);
or U4907 (N_4907,In_340,In_217);
nand U4908 (N_4908,In_457,In_357);
and U4909 (N_4909,In_75,In_218);
xnor U4910 (N_4910,In_676,In_287);
or U4911 (N_4911,In_273,In_675);
and U4912 (N_4912,In_607,In_473);
nand U4913 (N_4913,In_70,In_236);
nor U4914 (N_4914,In_376,In_795);
or U4915 (N_4915,In_903,In_96);
xor U4916 (N_4916,In_427,In_914);
or U4917 (N_4917,In_906,In_821);
and U4918 (N_4918,In_944,In_245);
xor U4919 (N_4919,In_304,In_960);
and U4920 (N_4920,In_320,In_737);
and U4921 (N_4921,In_606,In_536);
xnor U4922 (N_4922,In_52,In_140);
nor U4923 (N_4923,In_514,In_111);
nand U4924 (N_4924,In_768,In_15);
nand U4925 (N_4925,In_223,In_721);
nor U4926 (N_4926,In_177,In_977);
and U4927 (N_4927,In_515,In_74);
and U4928 (N_4928,In_777,In_527);
nor U4929 (N_4929,In_583,In_138);
and U4930 (N_4930,In_142,In_60);
or U4931 (N_4931,In_120,In_190);
xor U4932 (N_4932,In_117,In_353);
xor U4933 (N_4933,In_21,In_968);
and U4934 (N_4934,In_768,In_109);
nor U4935 (N_4935,In_38,In_168);
and U4936 (N_4936,In_271,In_863);
nor U4937 (N_4937,In_162,In_927);
and U4938 (N_4938,In_46,In_642);
and U4939 (N_4939,In_601,In_813);
and U4940 (N_4940,In_211,In_159);
xor U4941 (N_4941,In_788,In_525);
nor U4942 (N_4942,In_523,In_456);
nor U4943 (N_4943,In_313,In_428);
nor U4944 (N_4944,In_365,In_491);
nand U4945 (N_4945,In_754,In_824);
nand U4946 (N_4946,In_238,In_814);
and U4947 (N_4947,In_690,In_954);
nand U4948 (N_4948,In_949,In_781);
or U4949 (N_4949,In_2,In_866);
or U4950 (N_4950,In_520,In_206);
nand U4951 (N_4951,In_702,In_434);
nand U4952 (N_4952,In_543,In_750);
nor U4953 (N_4953,In_326,In_145);
and U4954 (N_4954,In_247,In_518);
xnor U4955 (N_4955,In_936,In_995);
nor U4956 (N_4956,In_253,In_223);
nor U4957 (N_4957,In_132,In_616);
or U4958 (N_4958,In_135,In_840);
xnor U4959 (N_4959,In_965,In_469);
nand U4960 (N_4960,In_755,In_846);
nand U4961 (N_4961,In_575,In_314);
and U4962 (N_4962,In_838,In_708);
nor U4963 (N_4963,In_535,In_641);
nand U4964 (N_4964,In_781,In_976);
nand U4965 (N_4965,In_158,In_459);
and U4966 (N_4966,In_667,In_376);
and U4967 (N_4967,In_437,In_839);
nand U4968 (N_4968,In_804,In_437);
or U4969 (N_4969,In_957,In_137);
nor U4970 (N_4970,In_371,In_403);
nand U4971 (N_4971,In_747,In_924);
nor U4972 (N_4972,In_130,In_859);
or U4973 (N_4973,In_194,In_310);
nand U4974 (N_4974,In_166,In_76);
nand U4975 (N_4975,In_341,In_382);
and U4976 (N_4976,In_896,In_40);
or U4977 (N_4977,In_546,In_202);
nor U4978 (N_4978,In_746,In_122);
nand U4979 (N_4979,In_763,In_547);
nor U4980 (N_4980,In_812,In_674);
or U4981 (N_4981,In_22,In_200);
nor U4982 (N_4982,In_388,In_167);
xor U4983 (N_4983,In_960,In_455);
nor U4984 (N_4984,In_70,In_394);
nand U4985 (N_4985,In_771,In_383);
and U4986 (N_4986,In_390,In_159);
and U4987 (N_4987,In_77,In_559);
nor U4988 (N_4988,In_932,In_214);
or U4989 (N_4989,In_754,In_165);
nor U4990 (N_4990,In_698,In_893);
nor U4991 (N_4991,In_285,In_448);
nand U4992 (N_4992,In_154,In_193);
and U4993 (N_4993,In_297,In_884);
nand U4994 (N_4994,In_21,In_465);
nand U4995 (N_4995,In_899,In_618);
and U4996 (N_4996,In_7,In_244);
or U4997 (N_4997,In_24,In_32);
or U4998 (N_4998,In_26,In_277);
xnor U4999 (N_4999,In_338,In_162);
nand U5000 (N_5000,N_3307,N_4144);
and U5001 (N_5001,N_154,N_887);
nor U5002 (N_5002,N_4378,N_1061);
and U5003 (N_5003,N_2316,N_3439);
and U5004 (N_5004,N_3776,N_4138);
nor U5005 (N_5005,N_4872,N_3441);
nand U5006 (N_5006,N_3453,N_14);
and U5007 (N_5007,N_1843,N_3855);
nor U5008 (N_5008,N_805,N_442);
and U5009 (N_5009,N_1840,N_1466);
nand U5010 (N_5010,N_594,N_2324);
xor U5011 (N_5011,N_3949,N_4371);
nor U5012 (N_5012,N_2006,N_3127);
nor U5013 (N_5013,N_2587,N_4042);
nor U5014 (N_5014,N_2075,N_3030);
and U5015 (N_5015,N_3994,N_770);
xor U5016 (N_5016,N_3344,N_4635);
nor U5017 (N_5017,N_4999,N_3697);
or U5018 (N_5018,N_60,N_4172);
and U5019 (N_5019,N_823,N_437);
nand U5020 (N_5020,N_3639,N_1679);
and U5021 (N_5021,N_406,N_2588);
nor U5022 (N_5022,N_32,N_3885);
nor U5023 (N_5023,N_683,N_1251);
or U5024 (N_5024,N_767,N_2394);
or U5025 (N_5025,N_4672,N_1726);
nand U5026 (N_5026,N_2156,N_620);
or U5027 (N_5027,N_636,N_4163);
nand U5028 (N_5028,N_2379,N_1921);
or U5029 (N_5029,N_2054,N_28);
or U5030 (N_5030,N_4058,N_1282);
and U5031 (N_5031,N_1980,N_4469);
and U5032 (N_5032,N_1108,N_1393);
and U5033 (N_5033,N_1274,N_3930);
or U5034 (N_5034,N_1511,N_4847);
or U5035 (N_5035,N_3286,N_3736);
nand U5036 (N_5036,N_3141,N_3998);
xor U5037 (N_5037,N_1874,N_3982);
nand U5038 (N_5038,N_13,N_666);
nand U5039 (N_5039,N_1261,N_2363);
or U5040 (N_5040,N_1837,N_2844);
nor U5041 (N_5041,N_1468,N_734);
nand U5042 (N_5042,N_3508,N_4094);
and U5043 (N_5043,N_1407,N_1971);
and U5044 (N_5044,N_170,N_1758);
nor U5045 (N_5045,N_2958,N_963);
or U5046 (N_5046,N_2777,N_1250);
nor U5047 (N_5047,N_3381,N_3246);
and U5048 (N_5048,N_3212,N_3694);
or U5049 (N_5049,N_644,N_4742);
or U5050 (N_5050,N_567,N_3415);
nand U5051 (N_5051,N_4297,N_3470);
and U5052 (N_5052,N_2366,N_648);
and U5053 (N_5053,N_2430,N_4400);
and U5054 (N_5054,N_744,N_305);
nor U5055 (N_5055,N_3714,N_3443);
xnor U5056 (N_5056,N_3020,N_545);
or U5057 (N_5057,N_1849,N_3856);
nor U5058 (N_5058,N_565,N_1053);
and U5059 (N_5059,N_1464,N_586);
or U5060 (N_5060,N_2954,N_2769);
and U5061 (N_5061,N_2544,N_3250);
xor U5062 (N_5062,N_921,N_4521);
and U5063 (N_5063,N_2778,N_1986);
nor U5064 (N_5064,N_1516,N_1804);
nand U5065 (N_5065,N_2765,N_3922);
or U5066 (N_5066,N_1982,N_2618);
nor U5067 (N_5067,N_896,N_317);
nor U5068 (N_5068,N_4804,N_4468);
and U5069 (N_5069,N_1071,N_2716);
nor U5070 (N_5070,N_819,N_3379);
or U5071 (N_5071,N_3341,N_1336);
xnor U5072 (N_5072,N_4370,N_917);
nor U5073 (N_5073,N_3901,N_2894);
nor U5074 (N_5074,N_2758,N_2371);
and U5075 (N_5075,N_2627,N_2891);
nor U5076 (N_5076,N_4159,N_3013);
or U5077 (N_5077,N_112,N_1182);
xnor U5078 (N_5078,N_109,N_4887);
xnor U5079 (N_5079,N_414,N_3108);
or U5080 (N_5080,N_272,N_4553);
nor U5081 (N_5081,N_3870,N_3647);
or U5082 (N_5082,N_4272,N_1345);
nor U5083 (N_5083,N_4942,N_3792);
nand U5084 (N_5084,N_1825,N_4634);
nand U5085 (N_5085,N_2550,N_4682);
and U5086 (N_5086,N_3198,N_1927);
or U5087 (N_5087,N_144,N_621);
nand U5088 (N_5088,N_3176,N_3819);
or U5089 (N_5089,N_4707,N_4274);
and U5090 (N_5090,N_2412,N_4994);
nand U5091 (N_5091,N_2672,N_1458);
nor U5092 (N_5092,N_1646,N_4062);
nor U5093 (N_5093,N_4348,N_1950);
or U5094 (N_5094,N_4245,N_4109);
or U5095 (N_5095,N_4552,N_2142);
and U5096 (N_5096,N_3906,N_3703);
and U5097 (N_5097,N_438,N_39);
or U5098 (N_5098,N_2434,N_1203);
nand U5099 (N_5099,N_2116,N_1710);
nor U5100 (N_5100,N_1248,N_3527);
or U5101 (N_5101,N_3000,N_2056);
nor U5102 (N_5102,N_3388,N_2942);
nand U5103 (N_5103,N_1272,N_3285);
or U5104 (N_5104,N_4064,N_88);
or U5105 (N_5105,N_1830,N_4656);
xnor U5106 (N_5106,N_4751,N_1500);
xor U5107 (N_5107,N_390,N_1519);
xor U5108 (N_5108,N_2915,N_2922);
nor U5109 (N_5109,N_418,N_4915);
or U5110 (N_5110,N_2904,N_2433);
or U5111 (N_5111,N_167,N_709);
nor U5112 (N_5112,N_2037,N_4797);
nor U5113 (N_5113,N_3546,N_1300);
xor U5114 (N_5114,N_435,N_3917);
and U5115 (N_5115,N_1976,N_1910);
nor U5116 (N_5116,N_153,N_123);
xor U5117 (N_5117,N_2735,N_1659);
nand U5118 (N_5118,N_2086,N_1795);
nor U5119 (N_5119,N_1010,N_1496);
xnor U5120 (N_5120,N_451,N_925);
and U5121 (N_5121,N_3366,N_4228);
nor U5122 (N_5122,N_331,N_4305);
and U5123 (N_5123,N_445,N_219);
and U5124 (N_5124,N_2516,N_2873);
xor U5125 (N_5125,N_1836,N_1457);
nor U5126 (N_5126,N_2034,N_1227);
nand U5127 (N_5127,N_4281,N_3663);
nor U5128 (N_5128,N_1286,N_25);
and U5129 (N_5129,N_537,N_1588);
nand U5130 (N_5130,N_1509,N_473);
xor U5131 (N_5131,N_3566,N_3825);
xor U5132 (N_5132,N_4466,N_4736);
and U5133 (N_5133,N_2595,N_3710);
nor U5134 (N_5134,N_3996,N_1696);
nand U5135 (N_5135,N_4750,N_2444);
nor U5136 (N_5136,N_1740,N_4752);
nand U5137 (N_5137,N_3808,N_2380);
or U5138 (N_5138,N_212,N_2402);
and U5139 (N_5139,N_1481,N_2918);
nand U5140 (N_5140,N_1290,N_4203);
nand U5141 (N_5141,N_4963,N_4002);
nor U5142 (N_5142,N_2538,N_2440);
or U5143 (N_5143,N_3383,N_2274);
or U5144 (N_5144,N_4168,N_1433);
nand U5145 (N_5145,N_1903,N_183);
nor U5146 (N_5146,N_4800,N_3175);
nor U5147 (N_5147,N_141,N_4410);
or U5148 (N_5148,N_2928,N_1949);
or U5149 (N_5149,N_3425,N_4354);
xor U5150 (N_5150,N_3724,N_3923);
nor U5151 (N_5151,N_3753,N_3993);
and U5152 (N_5152,N_3267,N_2344);
nand U5153 (N_5153,N_4366,N_3317);
nand U5154 (N_5154,N_814,N_3665);
and U5155 (N_5155,N_3177,N_2685);
nor U5156 (N_5156,N_3274,N_3877);
and U5157 (N_5157,N_3931,N_4383);
and U5158 (N_5158,N_4584,N_1121);
or U5159 (N_5159,N_511,N_2136);
or U5160 (N_5160,N_4987,N_1177);
xor U5161 (N_5161,N_42,N_4143);
nor U5162 (N_5162,N_3880,N_1224);
nand U5163 (N_5163,N_1213,N_3801);
or U5164 (N_5164,N_1576,N_3152);
or U5165 (N_5165,N_4500,N_3109);
and U5166 (N_5166,N_249,N_4294);
xor U5167 (N_5167,N_4273,N_1629);
and U5168 (N_5168,N_3651,N_1941);
nand U5169 (N_5169,N_4463,N_3363);
or U5170 (N_5170,N_1233,N_427);
or U5171 (N_5171,N_2794,N_951);
nand U5172 (N_5172,N_3131,N_3616);
nand U5173 (N_5173,N_613,N_580);
nor U5174 (N_5174,N_577,N_4063);
xor U5175 (N_5175,N_3833,N_4097);
or U5176 (N_5176,N_4701,N_3796);
nand U5177 (N_5177,N_865,N_3688);
nor U5178 (N_5178,N_3079,N_987);
and U5179 (N_5179,N_3253,N_2214);
and U5180 (N_5180,N_2376,N_1166);
and U5181 (N_5181,N_3056,N_992);
or U5182 (N_5182,N_4379,N_3842);
nand U5183 (N_5183,N_3029,N_3895);
or U5184 (N_5184,N_1819,N_1926);
or U5185 (N_5185,N_4661,N_4067);
or U5186 (N_5186,N_1195,N_206);
nand U5187 (N_5187,N_1403,N_2682);
nand U5188 (N_5188,N_352,N_999);
nor U5189 (N_5189,N_3794,N_2955);
nand U5190 (N_5190,N_2767,N_888);
and U5191 (N_5191,N_1953,N_1373);
xor U5192 (N_5192,N_4938,N_4928);
and U5193 (N_5193,N_1120,N_4591);
or U5194 (N_5194,N_4706,N_713);
nand U5195 (N_5195,N_1262,N_3186);
nand U5196 (N_5196,N_924,N_407);
nand U5197 (N_5197,N_4194,N_3843);
or U5198 (N_5198,N_3898,N_2077);
nand U5199 (N_5199,N_1367,N_3699);
nor U5200 (N_5200,N_561,N_812);
and U5201 (N_5201,N_4319,N_4766);
nor U5202 (N_5202,N_2471,N_3164);
nand U5203 (N_5203,N_2935,N_1324);
nand U5204 (N_5204,N_4489,N_936);
nor U5205 (N_5205,N_4747,N_3723);
nor U5206 (N_5206,N_3101,N_4032);
and U5207 (N_5207,N_4996,N_1967);
nor U5208 (N_5208,N_3720,N_4108);
nor U5209 (N_5209,N_3437,N_3064);
or U5210 (N_5210,N_3584,N_1278);
nand U5211 (N_5211,N_3272,N_747);
nand U5212 (N_5212,N_1868,N_2177);
xnor U5213 (N_5213,N_2602,N_2429);
nand U5214 (N_5214,N_4516,N_3838);
or U5215 (N_5215,N_609,N_2045);
and U5216 (N_5216,N_794,N_1800);
nand U5217 (N_5217,N_993,N_4445);
xnor U5218 (N_5218,N_1236,N_4806);
xor U5219 (N_5219,N_3042,N_3811);
and U5220 (N_5220,N_487,N_4594);
or U5221 (N_5221,N_4288,N_33);
and U5222 (N_5222,N_4531,N_1561);
xor U5223 (N_5223,N_4761,N_2872);
and U5224 (N_5224,N_3468,N_23);
nand U5225 (N_5225,N_2104,N_3913);
xnor U5226 (N_5226,N_4517,N_4611);
or U5227 (N_5227,N_984,N_470);
and U5228 (N_5228,N_505,N_2293);
or U5229 (N_5229,N_4035,N_2534);
nor U5230 (N_5230,N_3802,N_1332);
and U5231 (N_5231,N_825,N_3849);
and U5232 (N_5232,N_755,N_3134);
nand U5233 (N_5233,N_308,N_4432);
or U5234 (N_5234,N_4171,N_3247);
and U5235 (N_5235,N_4221,N_1657);
and U5236 (N_5236,N_2666,N_1304);
nand U5237 (N_5237,N_52,N_4433);
xor U5238 (N_5238,N_3325,N_253);
nand U5239 (N_5239,N_4808,N_824);
or U5240 (N_5240,N_4323,N_4258);
nand U5241 (N_5241,N_616,N_119);
nand U5242 (N_5242,N_4382,N_240);
or U5243 (N_5243,N_2524,N_903);
or U5244 (N_5244,N_3786,N_2657);
and U5245 (N_5245,N_4496,N_355);
nor U5246 (N_5246,N_1467,N_3268);
and U5247 (N_5247,N_4413,N_2360);
nand U5248 (N_5248,N_1655,N_3878);
nand U5249 (N_5249,N_2438,N_1906);
nor U5250 (N_5250,N_2493,N_3479);
nand U5251 (N_5251,N_997,N_3512);
nand U5252 (N_5252,N_877,N_945);
nand U5253 (N_5253,N_3826,N_4932);
xnor U5254 (N_5254,N_2292,N_2317);
or U5255 (N_5255,N_2604,N_4003);
or U5256 (N_5256,N_2377,N_4353);
nor U5257 (N_5257,N_1489,N_3306);
nand U5258 (N_5258,N_1198,N_676);
and U5259 (N_5259,N_3561,N_3912);
nor U5260 (N_5260,N_3160,N_1720);
xnor U5261 (N_5261,N_2178,N_1199);
nand U5262 (N_5262,N_3916,N_8);
or U5263 (N_5263,N_4230,N_3464);
and U5264 (N_5264,N_1383,N_3220);
and U5265 (N_5265,N_4749,N_2101);
nand U5266 (N_5266,N_497,N_1423);
xor U5267 (N_5267,N_920,N_3988);
nor U5268 (N_5268,N_185,N_1070);
nor U5269 (N_5269,N_4135,N_3618);
nor U5270 (N_5270,N_659,N_288);
nor U5271 (N_5271,N_3296,N_3503);
or U5272 (N_5272,N_353,N_4638);
nor U5273 (N_5273,N_4375,N_3195);
nor U5274 (N_5274,N_1578,N_2067);
or U5275 (N_5275,N_575,N_2082);
xnor U5276 (N_5276,N_283,N_2611);
nand U5277 (N_5277,N_907,N_2837);
nor U5278 (N_5278,N_4670,N_2912);
xnor U5279 (N_5279,N_3172,N_3829);
or U5280 (N_5280,N_1246,N_1252);
and U5281 (N_5281,N_4271,N_973);
nand U5282 (N_5282,N_83,N_2109);
xor U5283 (N_5283,N_2365,N_306);
xor U5284 (N_5284,N_1447,N_2966);
or U5285 (N_5285,N_4267,N_4420);
nor U5286 (N_5286,N_2031,N_341);
nor U5287 (N_5287,N_4089,N_981);
and U5288 (N_5288,N_3129,N_3444);
nor U5289 (N_5289,N_3867,N_3487);
nor U5290 (N_5290,N_496,N_886);
nand U5291 (N_5291,N_1875,N_1529);
nand U5292 (N_5292,N_4199,N_4033);
and U5293 (N_5293,N_4099,N_892);
nor U5294 (N_5294,N_939,N_2535);
and U5295 (N_5295,N_4438,N_2830);
or U5296 (N_5296,N_3461,N_3036);
nor U5297 (N_5297,N_2924,N_1148);
and U5298 (N_5298,N_560,N_4373);
and U5299 (N_5299,N_2449,N_4845);
nor U5300 (N_5300,N_1994,N_737);
xor U5301 (N_5301,N_1890,N_4139);
and U5302 (N_5302,N_1594,N_2882);
and U5303 (N_5303,N_1226,N_1190);
nand U5304 (N_5304,N_2736,N_1975);
or U5305 (N_5305,N_3427,N_2845);
and U5306 (N_5306,N_4912,N_1216);
xor U5307 (N_5307,N_3257,N_2683);
nor U5308 (N_5308,N_231,N_535);
or U5309 (N_5309,N_1015,N_1707);
nor U5310 (N_5310,N_328,N_4975);
nand U5311 (N_5311,N_2481,N_4494);
or U5312 (N_5312,N_1023,N_4873);
nand U5313 (N_5313,N_55,N_374);
and U5314 (N_5314,N_4302,N_3019);
and U5315 (N_5315,N_2393,N_1674);
xnor U5316 (N_5316,N_1438,N_2164);
and U5317 (N_5317,N_2373,N_4180);
and U5318 (N_5318,N_1682,N_4614);
nand U5319 (N_5319,N_2636,N_855);
and U5320 (N_5320,N_2853,N_2842);
or U5321 (N_5321,N_4493,N_938);
nor U5322 (N_5322,N_1144,N_2840);
or U5323 (N_5323,N_749,N_2585);
or U5324 (N_5324,N_1530,N_3100);
nand U5325 (N_5325,N_464,N_3418);
nand U5326 (N_5326,N_2149,N_3865);
or U5327 (N_5327,N_1970,N_3936);
or U5328 (N_5328,N_3778,N_4697);
and U5329 (N_5329,N_608,N_357);
and U5330 (N_5330,N_1220,N_434);
xor U5331 (N_5331,N_4709,N_1063);
nand U5332 (N_5332,N_1491,N_1887);
nor U5333 (N_5333,N_3386,N_3282);
and U5334 (N_5334,N_4911,N_398);
or U5335 (N_5335,N_3436,N_628);
nor U5336 (N_5336,N_841,N_1479);
or U5337 (N_5337,N_361,N_147);
and U5338 (N_5338,N_1571,N_489);
or U5339 (N_5339,N_4619,N_3679);
xnor U5340 (N_5340,N_4418,N_4934);
nand U5341 (N_5341,N_1384,N_289);
or U5342 (N_5342,N_3517,N_1968);
or U5343 (N_5343,N_3026,N_1590);
nor U5344 (N_5344,N_3634,N_2617);
or U5345 (N_5345,N_4939,N_1934);
xor U5346 (N_5346,N_964,N_932);
nand U5347 (N_5347,N_889,N_3368);
or U5348 (N_5348,N_576,N_3645);
or U5349 (N_5349,N_612,N_4023);
nand U5350 (N_5350,N_3822,N_2804);
or U5351 (N_5351,N_2515,N_1753);
nor U5352 (N_5352,N_4976,N_3223);
and U5353 (N_5353,N_4653,N_4000);
nor U5354 (N_5354,N_3620,N_4811);
nor U5355 (N_5355,N_2755,N_3623);
and U5356 (N_5356,N_867,N_2404);
nor U5357 (N_5357,N_1222,N_2332);
xnor U5358 (N_5358,N_453,N_956);
nor U5359 (N_5359,N_2581,N_3446);
or U5360 (N_5360,N_4728,N_1490);
xor U5361 (N_5361,N_2879,N_1852);
or U5362 (N_5362,N_3169,N_1204);
nor U5363 (N_5363,N_522,N_3067);
and U5364 (N_5364,N_3393,N_4457);
or U5365 (N_5365,N_2629,N_1879);
and U5366 (N_5366,N_4234,N_2382);
nand U5367 (N_5367,N_2841,N_2695);
nor U5368 (N_5368,N_2829,N_764);
nand U5369 (N_5369,N_4897,N_942);
xnor U5370 (N_5370,N_1784,N_1902);
and U5371 (N_5371,N_961,N_3312);
and U5372 (N_5372,N_670,N_1528);
nand U5373 (N_5373,N_2257,N_3509);
and U5374 (N_5374,N_4395,N_4151);
xor U5375 (N_5375,N_1164,N_379);
nand U5376 (N_5376,N_1087,N_4291);
and U5377 (N_5377,N_3583,N_1265);
nand U5378 (N_5378,N_4372,N_778);
or U5379 (N_5379,N_2354,N_2398);
nor U5380 (N_5380,N_2210,N_4338);
nor U5381 (N_5381,N_3330,N_4224);
nor U5382 (N_5382,N_2194,N_1109);
or U5383 (N_5383,N_4188,N_432);
or U5384 (N_5384,N_1340,N_2175);
or U5385 (N_5385,N_1572,N_1047);
and U5386 (N_5386,N_2776,N_4773);
xor U5387 (N_5387,N_2009,N_915);
or U5388 (N_5388,N_2172,N_4905);
and U5389 (N_5389,N_3073,N_108);
nor U5390 (N_5390,N_383,N_1983);
nor U5391 (N_5391,N_4166,N_2489);
or U5392 (N_5392,N_3232,N_3408);
and U5393 (N_5393,N_2941,N_1929);
nor U5394 (N_5394,N_2750,N_507);
and U5395 (N_5395,N_4001,N_772);
nand U5396 (N_5396,N_2472,N_935);
and U5397 (N_5397,N_4536,N_2867);
nand U5398 (N_5398,N_1469,N_251);
and U5399 (N_5399,N_1494,N_155);
nor U5400 (N_5400,N_2634,N_4786);
or U5401 (N_5401,N_2239,N_2367);
nor U5402 (N_5402,N_1106,N_4828);
nor U5403 (N_5403,N_4557,N_4982);
and U5404 (N_5404,N_2329,N_1689);
nor U5405 (N_5405,N_1142,N_1292);
nand U5406 (N_5406,N_4787,N_2105);
nor U5407 (N_5407,N_3119,N_2482);
nand U5408 (N_5408,N_3767,N_4237);
or U5409 (N_5409,N_3587,N_4152);
xnor U5410 (N_5410,N_2852,N_3151);
nand U5411 (N_5411,N_2410,N_4376);
nand U5412 (N_5412,N_2361,N_3486);
or U5413 (N_5413,N_4704,N_2388);
or U5414 (N_5414,N_2170,N_3200);
nand U5415 (N_5415,N_3277,N_640);
nand U5416 (N_5416,N_4121,N_2923);
xor U5417 (N_5417,N_160,N_4694);
nand U5418 (N_5418,N_3760,N_4101);
or U5419 (N_5419,N_330,N_4231);
and U5420 (N_5420,N_3084,N_2509);
and U5421 (N_5421,N_584,N_1211);
xnor U5422 (N_5422,N_4599,N_2222);
or U5423 (N_5423,N_4385,N_2181);
xnor U5424 (N_5424,N_4538,N_4443);
nor U5425 (N_5425,N_2927,N_4793);
nor U5426 (N_5426,N_752,N_4232);
and U5427 (N_5427,N_2754,N_806);
or U5428 (N_5428,N_1610,N_699);
nor U5429 (N_5429,N_3451,N_2994);
nand U5430 (N_5430,N_3422,N_1596);
and U5431 (N_5431,N_1193,N_1611);
nor U5432 (N_5432,N_856,N_3866);
or U5433 (N_5433,N_3733,N_3953);
xnor U5434 (N_5434,N_2235,N_3090);
nor U5435 (N_5435,N_3255,N_2058);
or U5436 (N_5436,N_4660,N_4763);
xnor U5437 (N_5437,N_1764,N_1427);
nor U5438 (N_5438,N_4542,N_2443);
or U5439 (N_5439,N_2151,N_1418);
and U5440 (N_5440,N_50,N_277);
and U5441 (N_5441,N_1169,N_2816);
and U5442 (N_5442,N_657,N_2134);
nand U5443 (N_5443,N_1456,N_2810);
xor U5444 (N_5444,N_1000,N_1998);
nand U5445 (N_5445,N_3372,N_4907);
and U5446 (N_5446,N_3832,N_2036);
or U5447 (N_5447,N_694,N_3705);
and U5448 (N_5448,N_4040,N_2176);
nand U5449 (N_5449,N_2702,N_2762);
or U5450 (N_5450,N_3555,N_264);
nand U5451 (N_5451,N_40,N_669);
nor U5452 (N_5452,N_73,N_3224);
xor U5453 (N_5453,N_4822,N_3681);
nor U5454 (N_5454,N_501,N_1854);
or U5455 (N_5455,N_2578,N_4947);
nor U5456 (N_5456,N_1989,N_3984);
or U5457 (N_5457,N_692,N_2661);
or U5458 (N_5458,N_4504,N_2589);
or U5459 (N_5459,N_269,N_3745);
nor U5460 (N_5460,N_4283,N_16);
or U5461 (N_5461,N_3412,N_2798);
and U5462 (N_5462,N_547,N_2263);
and U5463 (N_5463,N_928,N_2949);
and U5464 (N_5464,N_1221,N_1280);
or U5465 (N_5465,N_1358,N_3511);
nand U5466 (N_5466,N_930,N_93);
nand U5467 (N_5467,N_549,N_603);
xnor U5468 (N_5468,N_1871,N_1425);
or U5469 (N_5469,N_1586,N_4765);
nor U5470 (N_5470,N_1894,N_1513);
and U5471 (N_5471,N_4598,N_1256);
and U5472 (N_5472,N_3294,N_4544);
nand U5473 (N_5473,N_4859,N_1567);
or U5474 (N_5474,N_1125,N_2183);
or U5475 (N_5475,N_2158,N_2061);
and U5476 (N_5476,N_3331,N_661);
or U5477 (N_5477,N_4356,N_4080);
nor U5478 (N_5478,N_4241,N_1492);
or U5479 (N_5479,N_1102,N_4309);
xor U5480 (N_5480,N_879,N_1900);
and U5481 (N_5481,N_2732,N_1766);
xor U5482 (N_5482,N_1618,N_708);
nor U5483 (N_5483,N_3899,N_1090);
xor U5484 (N_5484,N_2824,N_465);
and U5485 (N_5485,N_3513,N_4970);
and U5486 (N_5486,N_3932,N_3962);
nor U5487 (N_5487,N_1913,N_1330);
nand U5488 (N_5488,N_4861,N_1709);
nand U5489 (N_5489,N_1035,N_509);
nor U5490 (N_5490,N_3083,N_3840);
nor U5491 (N_5491,N_3188,N_732);
and U5492 (N_5492,N_1229,N_989);
or U5493 (N_5493,N_583,N_4325);
xnor U5494 (N_5494,N_2473,N_2261);
and U5495 (N_5495,N_1756,N_4113);
nor U5496 (N_5496,N_2582,N_1381);
nand U5497 (N_5497,N_1559,N_3295);
nand U5498 (N_5498,N_1680,N_4729);
xnor U5499 (N_5499,N_38,N_2890);
nor U5500 (N_5500,N_2335,N_385);
xnor U5501 (N_5501,N_3991,N_2610);
xor U5502 (N_5502,N_788,N_3148);
or U5503 (N_5503,N_4546,N_4406);
nor U5504 (N_5504,N_3092,N_1692);
xor U5505 (N_5505,N_4147,N_4190);
nor U5506 (N_5506,N_2147,N_2499);
nor U5507 (N_5507,N_3967,N_4702);
nor U5508 (N_5508,N_349,N_3920);
and U5509 (N_5509,N_3270,N_4606);
and U5510 (N_5510,N_368,N_4346);
nand U5511 (N_5511,N_3021,N_562);
nor U5512 (N_5512,N_3828,N_191);
and U5513 (N_5513,N_4005,N_4512);
nand U5514 (N_5514,N_161,N_2281);
nor U5515 (N_5515,N_2246,N_4387);
nand U5516 (N_5516,N_2770,N_2011);
and U5517 (N_5517,N_4242,N_417);
and U5518 (N_5518,N_3287,N_4290);
and U5519 (N_5519,N_4876,N_2139);
or U5520 (N_5520,N_1557,N_1257);
or U5521 (N_5521,N_2032,N_492);
or U5522 (N_5522,N_1593,N_1137);
xnor U5523 (N_5523,N_1553,N_3876);
and U5524 (N_5524,N_1454,N_701);
nor U5525 (N_5525,N_3156,N_4936);
nand U5526 (N_5526,N_4015,N_3574);
and U5527 (N_5527,N_1311,N_2639);
xor U5528 (N_5528,N_4472,N_1534);
or U5529 (N_5529,N_4452,N_1249);
or U5530 (N_5530,N_2635,N_4110);
and U5531 (N_5531,N_4365,N_3735);
xnor U5532 (N_5532,N_4096,N_1757);
nor U5533 (N_5533,N_1329,N_4017);
or U5534 (N_5534,N_1339,N_3674);
or U5535 (N_5535,N_801,N_2742);
nand U5536 (N_5536,N_3426,N_138);
nor U5537 (N_5537,N_4501,N_1560);
nand U5538 (N_5538,N_2125,N_2740);
nand U5539 (N_5539,N_1622,N_3995);
xnor U5540 (N_5540,N_190,N_654);
and U5541 (N_5541,N_3279,N_2046);
nand U5542 (N_5542,N_3219,N_4078);
nand U5543 (N_5543,N_1397,N_2013);
nand U5544 (N_5544,N_3406,N_213);
nand U5545 (N_5545,N_1714,N_2463);
and U5546 (N_5546,N_1880,N_1793);
nand U5547 (N_5547,N_67,N_4451);
nor U5548 (N_5548,N_1940,N_949);
and U5549 (N_5549,N_4102,N_4439);
nand U5550 (N_5550,N_4481,N_1573);
nand U5551 (N_5551,N_181,N_4367);
or U5552 (N_5552,N_4721,N_908);
nand U5553 (N_5553,N_4627,N_1991);
nand U5554 (N_5554,N_578,N_2939);
xnor U5555 (N_5555,N_2518,N_2656);
nand U5556 (N_5556,N_486,N_4154);
or U5557 (N_5557,N_672,N_1029);
nand U5558 (N_5558,N_3118,N_2899);
nor U5559 (N_5559,N_1535,N_1021);
nand U5560 (N_5560,N_1092,N_598);
or U5561 (N_5561,N_2039,N_839);
xnor U5562 (N_5562,N_4571,N_335);
or U5563 (N_5563,N_1574,N_4559);
xnor U5564 (N_5564,N_3396,N_3480);
nand U5565 (N_5565,N_4940,N_1732);
and U5566 (N_5566,N_1592,N_128);
nor U5567 (N_5567,N_292,N_2505);
or U5568 (N_5568,N_627,N_2179);
nand U5569 (N_5569,N_4588,N_4465);
nand U5570 (N_5570,N_479,N_2290);
or U5571 (N_5571,N_455,N_2352);
and U5572 (N_5572,N_1037,N_3027);
or U5573 (N_5573,N_4795,N_2648);
nand U5574 (N_5574,N_4509,N_2881);
nand U5575 (N_5575,N_4448,N_765);
nor U5576 (N_5576,N_1052,N_974);
and U5577 (N_5577,N_3040,N_2469);
nor U5578 (N_5578,N_2917,N_1270);
or U5579 (N_5579,N_4260,N_2312);
nand U5580 (N_5580,N_1392,N_3554);
nor U5581 (N_5581,N_3732,N_4201);
or U5582 (N_5582,N_2231,N_4415);
or U5583 (N_5583,N_44,N_1380);
or U5584 (N_5584,N_295,N_484);
nand U5585 (N_5585,N_2229,N_3891);
and U5586 (N_5586,N_1684,N_1542);
or U5587 (N_5587,N_2334,N_3248);
nand U5588 (N_5588,N_775,N_4657);
and U5589 (N_5589,N_4009,N_2734);
or U5590 (N_5590,N_1738,N_3947);
xnor U5591 (N_5591,N_1355,N_3283);
nand U5592 (N_5592,N_3450,N_4025);
nand U5593 (N_5593,N_4184,N_3698);
or U5594 (N_5594,N_3756,N_2240);
or U5595 (N_5595,N_3628,N_3273);
or U5596 (N_5596,N_4674,N_140);
xnor U5597 (N_5597,N_2987,N_2284);
or U5598 (N_5598,N_3249,N_4885);
xnor U5599 (N_5599,N_168,N_4671);
xnor U5600 (N_5600,N_78,N_4727);
or U5601 (N_5601,N_397,N_4175);
and U5602 (N_5602,N_3636,N_2028);
and U5603 (N_5603,N_934,N_1116);
nand U5604 (N_5604,N_3552,N_2159);
nor U5605 (N_5605,N_3977,N_568);
and U5606 (N_5606,N_2145,N_3711);
nand U5607 (N_5607,N_3975,N_1315);
and U5608 (N_5608,N_103,N_4212);
nand U5609 (N_5609,N_4183,N_1059);
and U5610 (N_5610,N_122,N_3338);
nor U5611 (N_5611,N_202,N_4510);
or U5612 (N_5612,N_2189,N_2849);
nor U5613 (N_5613,N_3667,N_847);
nand U5614 (N_5614,N_2706,N_4879);
nand U5615 (N_5615,N_1883,N_836);
and U5616 (N_5616,N_3890,N_3238);
and U5617 (N_5617,N_3664,N_2791);
and U5618 (N_5618,N_553,N_914);
and U5619 (N_5619,N_395,N_1742);
or U5620 (N_5620,N_3918,N_3942);
and U5621 (N_5621,N_679,N_2403);
nor U5622 (N_5622,N_439,N_1178);
xnor U5623 (N_5623,N_1154,N_3231);
and U5624 (N_5624,N_3979,N_2549);
or U5625 (N_5625,N_1207,N_651);
or U5626 (N_5626,N_2932,N_1767);
or U5627 (N_5627,N_475,N_1214);
nand U5628 (N_5628,N_4105,N_2305);
nand U5629 (N_5629,N_1253,N_3434);
nor U5630 (N_5630,N_2820,N_401);
nor U5631 (N_5631,N_2323,N_63);
and U5632 (N_5632,N_3862,N_145);
nand U5633 (N_5633,N_51,N_2594);
nor U5634 (N_5634,N_4589,N_2282);
xnor U5635 (N_5635,N_9,N_2536);
or U5636 (N_5636,N_1939,N_4084);
and U5637 (N_5637,N_596,N_1094);
and U5638 (N_5638,N_3501,N_4208);
or U5639 (N_5639,N_3680,N_4579);
or U5640 (N_5640,N_129,N_286);
and U5641 (N_5641,N_791,N_808);
and U5642 (N_5642,N_2992,N_3058);
or U5643 (N_5643,N_91,N_4675);
nand U5644 (N_5644,N_4809,N_4477);
nand U5645 (N_5645,N_194,N_2828);
xor U5646 (N_5646,N_4525,N_3215);
and U5647 (N_5647,N_4658,N_1708);
nand U5648 (N_5648,N_1275,N_2783);
and U5649 (N_5649,N_4286,N_287);
nand U5650 (N_5650,N_1930,N_2593);
nor U5651 (N_5651,N_1920,N_4296);
or U5652 (N_5652,N_4174,N_3959);
xor U5653 (N_5653,N_1683,N_224);
or U5654 (N_5654,N_1243,N_2021);
and U5655 (N_5655,N_4044,N_197);
and U5656 (N_5656,N_4743,N_3668);
nor U5657 (N_5657,N_4558,N_2268);
or U5658 (N_5658,N_1587,N_503);
xnor U5659 (N_5659,N_4287,N_3500);
nor U5660 (N_5660,N_2107,N_4490);
and U5661 (N_5661,N_301,N_148);
nand U5662 (N_5662,N_4858,N_2501);
and U5663 (N_5663,N_1310,N_3173);
xor U5664 (N_5664,N_2863,N_102);
or U5665 (N_5665,N_2539,N_4303);
and U5666 (N_5666,N_3162,N_4050);
or U5667 (N_5667,N_2678,N_2108);
xor U5668 (N_5668,N_2040,N_3060);
or U5669 (N_5669,N_1984,N_2756);
nand U5670 (N_5670,N_1729,N_2553);
nor U5671 (N_5671,N_3696,N_599);
and U5672 (N_5672,N_2609,N_3646);
and U5673 (N_5673,N_4846,N_4550);
and U5674 (N_5674,N_2739,N_1394);
nand U5675 (N_5675,N_3097,N_211);
or U5676 (N_5676,N_2168,N_4083);
and U5677 (N_5677,N_1161,N_205);
nand U5678 (N_5678,N_2823,N_3834);
nand U5679 (N_5679,N_2573,N_4430);
xor U5680 (N_5680,N_459,N_2626);
and U5681 (N_5681,N_2960,N_382);
nor U5682 (N_5682,N_2174,N_250);
nor U5683 (N_5683,N_4548,N_3218);
nand U5684 (N_5684,N_4864,N_1273);
and U5685 (N_5685,N_4259,N_3689);
nor U5686 (N_5686,N_279,N_2864);
and U5687 (N_5687,N_3709,N_4106);
nor U5688 (N_5688,N_2401,N_3447);
or U5689 (N_5689,N_4350,N_4349);
or U5690 (N_5690,N_2300,N_1321);
or U5691 (N_5691,N_2461,N_4953);
and U5692 (N_5692,N_719,N_2192);
nor U5693 (N_5693,N_3271,N_840);
and U5694 (N_5694,N_828,N_4345);
and U5695 (N_5695,N_142,N_702);
nand U5696 (N_5696,N_4758,N_4875);
and U5697 (N_5697,N_2291,N_3375);
nand U5698 (N_5698,N_3612,N_4256);
and U5699 (N_5699,N_821,N_1602);
or U5700 (N_5700,N_1077,N_4043);
or U5701 (N_5701,N_2537,N_3204);
nor U5702 (N_5702,N_2940,N_911);
or U5703 (N_5703,N_3599,N_2605);
nand U5704 (N_5704,N_2936,N_1086);
nor U5705 (N_5705,N_2081,N_36);
or U5706 (N_5706,N_3194,N_4791);
or U5707 (N_5707,N_1728,N_1350);
nand U5708 (N_5708,N_1434,N_893);
nand U5709 (N_5709,N_4798,N_1685);
and U5710 (N_5710,N_3759,N_4262);
nand U5711 (N_5711,N_4275,N_1671);
and U5712 (N_5712,N_2933,N_4825);
nand U5713 (N_5713,N_1140,N_954);
and U5714 (N_5714,N_1378,N_1391);
and U5715 (N_5715,N_3768,N_3661);
or U5716 (N_5716,N_717,N_3600);
and U5717 (N_5717,N_4498,N_3577);
nor U5718 (N_5718,N_3506,N_1111);
nor U5719 (N_5719,N_4951,N_3637);
and U5720 (N_5720,N_4813,N_230);
nand U5721 (N_5721,N_508,N_860);
xnor U5722 (N_5722,N_389,N_1595);
and U5723 (N_5723,N_1565,N_995);
xnor U5724 (N_5724,N_4978,N_4645);
or U5725 (N_5725,N_4789,N_4980);
and U5726 (N_5726,N_3591,N_3262);
nor U5727 (N_5727,N_1523,N_554);
and U5728 (N_5728,N_3174,N_3990);
xor U5729 (N_5729,N_4524,N_4414);
xor U5730 (N_5730,N_3281,N_4254);
nor U5731 (N_5731,N_3763,N_4399);
xor U5732 (N_5732,N_273,N_3941);
and U5733 (N_5733,N_4577,N_3448);
or U5734 (N_5734,N_1325,N_1797);
or U5735 (N_5735,N_3254,N_884);
nand U5736 (N_5736,N_2171,N_4683);
or U5737 (N_5737,N_2838,N_298);
and U5738 (N_5738,N_4126,N_4479);
or U5739 (N_5739,N_215,N_3691);
or U5740 (N_5740,N_421,N_1642);
nand U5741 (N_5741,N_902,N_2567);
nor U5742 (N_5742,N_2447,N_4893);
nor U5743 (N_5743,N_506,N_1711);
nand U5744 (N_5744,N_158,N_2862);
nor U5745 (N_5745,N_990,N_871);
nand U5746 (N_5746,N_1677,N_4146);
nor U5747 (N_5747,N_2907,N_1548);
xor U5748 (N_5748,N_493,N_2066);
or U5749 (N_5749,N_4625,N_1580);
nor U5750 (N_5750,N_4329,N_3362);
nand U5751 (N_5751,N_2019,N_4013);
and U5752 (N_5752,N_4107,N_3851);
nor U5753 (N_5753,N_164,N_3364);
nand U5754 (N_5754,N_2720,N_4903);
nand U5755 (N_5755,N_766,N_3061);
and U5756 (N_5756,N_4666,N_3754);
nand U5757 (N_5757,N_1189,N_4985);
nand U5758 (N_5758,N_1319,N_1068);
and U5759 (N_5759,N_4347,N_2114);
or U5760 (N_5760,N_136,N_233);
and U5761 (N_5761,N_315,N_4223);
xnor U5762 (N_5762,N_3111,N_3044);
nand U5763 (N_5763,N_2267,N_1547);
nand U5764 (N_5764,N_2091,N_3730);
nand U5765 (N_5765,N_1351,N_2253);
or U5766 (N_5766,N_3106,N_3588);
nand U5767 (N_5767,N_1072,N_4407);
and U5768 (N_5768,N_3065,N_3033);
nor U5769 (N_5769,N_721,N_21);
nor U5770 (N_5770,N_232,N_3971);
nand U5771 (N_5771,N_3496,N_2999);
nand U5772 (N_5772,N_1312,N_3069);
or U5773 (N_5773,N_1223,N_4663);
and U5774 (N_5774,N_2556,N_1091);
nor U5775 (N_5775,N_4837,N_4604);
and U5776 (N_5776,N_81,N_3835);
xnor U5777 (N_5777,N_2254,N_607);
xnor U5778 (N_5778,N_2647,N_574);
or U5779 (N_5779,N_3844,N_4087);
nand U5780 (N_5780,N_722,N_4);
xor U5781 (N_5781,N_3476,N_834);
nand U5782 (N_5782,N_3521,N_2963);
nor U5783 (N_5783,N_4495,N_4768);
and U5784 (N_5784,N_420,N_3999);
and U5785 (N_5785,N_872,N_838);
nand U5786 (N_5786,N_1598,N_1406);
or U5787 (N_5787,N_1855,N_975);
and U5788 (N_5788,N_2586,N_1891);
or U5789 (N_5789,N_2191,N_3442);
or U5790 (N_5790,N_4198,N_1196);
nand U5791 (N_5791,N_54,N_3046);
nor U5792 (N_5792,N_4642,N_853);
nand U5793 (N_5793,N_3823,N_2005);
and U5794 (N_5794,N_4028,N_4610);
or U5795 (N_5795,N_3209,N_4251);
nand U5796 (N_5796,N_2485,N_3657);
or U5797 (N_5797,N_753,N_89);
xnor U5798 (N_5798,N_1483,N_4079);
nor U5799 (N_5799,N_241,N_1577);
and U5800 (N_5800,N_2413,N_874);
nor U5801 (N_5801,N_901,N_1947);
nor U5802 (N_5802,N_1518,N_3551);
or U5803 (N_5803,N_1656,N_1905);
and U5804 (N_5804,N_2646,N_290);
nand U5805 (N_5805,N_491,N_2700);
and U5806 (N_5806,N_1563,N_2458);
nand U5807 (N_5807,N_4778,N_2638);
and U5808 (N_5808,N_1556,N_110);
or U5809 (N_5809,N_4944,N_499);
and U5810 (N_5810,N_696,N_1485);
and U5811 (N_5811,N_582,N_4162);
nand U5812 (N_5812,N_754,N_1877);
or U5813 (N_5813,N_3731,N_1401);
and U5814 (N_5814,N_1143,N_3686);
nor U5815 (N_5815,N_2785,N_2523);
nand U5816 (N_5816,N_463,N_1873);
nand U5817 (N_5817,N_2022,N_4026);
or U5818 (N_5818,N_2351,N_1631);
nor U5819 (N_5819,N_2285,N_75);
nand U5820 (N_5820,N_1727,N_2896);
or U5821 (N_5821,N_156,N_4889);
nor U5822 (N_5822,N_3499,N_4781);
nor U5823 (N_5823,N_1411,N_4997);
and U5824 (N_5824,N_4217,N_3430);
or U5825 (N_5825,N_4070,N_873);
nand U5826 (N_5826,N_2569,N_3197);
nand U5827 (N_5827,N_3677,N_2527);
nand U5828 (N_5828,N_2321,N_3650);
nand U5829 (N_5829,N_4990,N_3649);
nor U5830 (N_5830,N_1022,N_422);
nand U5831 (N_5831,N_4404,N_2336);
and U5832 (N_5832,N_4870,N_2146);
nor U5833 (N_5833,N_3087,N_1997);
or U5834 (N_5834,N_4590,N_3653);
nor U5835 (N_5835,N_1859,N_3099);
xor U5836 (N_5836,N_3354,N_2921);
or U5837 (N_5837,N_706,N_1626);
nor U5838 (N_5838,N_366,N_4722);
nand U5839 (N_5839,N_65,N_4735);
and U5840 (N_5840,N_113,N_329);
or U5841 (N_5841,N_1990,N_1388);
or U5842 (N_5842,N_3739,N_3171);
or U5843 (N_5843,N_3007,N_1952);
nand U5844 (N_5844,N_4030,N_2141);
and U5845 (N_5845,N_829,N_3278);
or U5846 (N_5846,N_1649,N_3568);
or U5847 (N_5847,N_2744,N_4782);
or U5848 (N_5848,N_1958,N_4744);
nand U5849 (N_5849,N_2358,N_1041);
nand U5850 (N_5850,N_2007,N_4233);
nand U5851 (N_5851,N_4193,N_6);
nand U5852 (N_5852,N_3259,N_2866);
and U5853 (N_5853,N_2885,N_4012);
nand U5854 (N_5854,N_2399,N_1385);
xor U5855 (N_5855,N_4336,N_3516);
nand U5856 (N_5856,N_413,N_1546);
nor U5857 (N_5857,N_2089,N_3750);
and U5858 (N_5858,N_105,N_3035);
or U5859 (N_5859,N_1165,N_408);
nand U5860 (N_5860,N_2956,N_2484);
nand U5861 (N_5861,N_2825,N_2381);
nor U5862 (N_5862,N_96,N_4422);
nand U5863 (N_5863,N_2016,N_2123);
and U5864 (N_5864,N_1759,N_246);
nand U5865 (N_5865,N_2834,N_4453);
or U5866 (N_5866,N_2592,N_4711);
xor U5867 (N_5867,N_454,N_1503);
and U5868 (N_5868,N_3562,N_1167);
and U5869 (N_5869,N_1141,N_3817);
nor U5870 (N_5870,N_4318,N_4626);
or U5871 (N_5871,N_1507,N_2737);
xnor U5872 (N_5872,N_3384,N_3718);
or U5873 (N_5873,N_3903,N_4377);
or U5874 (N_5874,N_2884,N_4880);
or U5875 (N_5875,N_2161,N_4431);
or U5876 (N_5876,N_45,N_1453);
or U5877 (N_5877,N_1153,N_4118);
nor U5878 (N_5878,N_2185,N_4899);
and U5879 (N_5879,N_1181,N_2901);
nor U5880 (N_5880,N_2318,N_2888);
nand U5881 (N_5881,N_4476,N_4686);
and U5882 (N_5882,N_180,N_2460);
or U5883 (N_5883,N_2049,N_485);
or U5884 (N_5884,N_912,N_1609);
nand U5885 (N_5885,N_1426,N_3514);
nor U5886 (N_5886,N_3687,N_4441);
nor U5887 (N_5887,N_3701,N_4330);
and U5888 (N_5888,N_3859,N_1404);
or U5889 (N_5889,N_3497,N_3672);
xor U5890 (N_5890,N_1735,N_4908);
nor U5891 (N_5891,N_803,N_458);
xor U5892 (N_5892,N_2003,N_4851);
nor U5893 (N_5893,N_1841,N_1117);
nor U5894 (N_5894,N_3445,N_3598);
nor U5895 (N_5895,N_1835,N_371);
xnor U5896 (N_5896,N_1600,N_529);
and U5897 (N_5897,N_2980,N_3524);
nand U5898 (N_5898,N_2997,N_1667);
and U5899 (N_5899,N_2584,N_1884);
nand U5900 (N_5900,N_4182,N_3845);
and U5901 (N_5901,N_1459,N_786);
and U5902 (N_5902,N_3181,N_2269);
or U5903 (N_5903,N_1695,N_3103);
nand U5904 (N_5904,N_1865,N_2406);
nand U5905 (N_5905,N_2790,N_3006);
and U5906 (N_5906,N_256,N_736);
xor U5907 (N_5907,N_3590,N_3413);
nor U5908 (N_5908,N_700,N_4358);
nor U5909 (N_5909,N_440,N_813);
or U5910 (N_5910,N_2397,N_3606);
and U5911 (N_5911,N_2200,N_4142);
and U5912 (N_5912,N_2247,N_143);
and U5913 (N_5913,N_1156,N_2805);
or U5914 (N_5914,N_1612,N_163);
and U5915 (N_5915,N_3682,N_4529);
or U5916 (N_5916,N_2715,N_4351);
and U5917 (N_5917,N_1653,N_1691);
nor U5918 (N_5918,N_4304,N_1123);
or U5919 (N_5919,N_988,N_2779);
or U5920 (N_5920,N_4470,N_4461);
or U5921 (N_5921,N_1614,N_4613);
nand U5922 (N_5922,N_1132,N_1042);
or U5923 (N_5923,N_4902,N_4519);
nand U5924 (N_5924,N_234,N_2787);
nor U5925 (N_5925,N_1549,N_80);
xnor U5926 (N_5926,N_24,N_2616);
xnor U5927 (N_5927,N_2971,N_1361);
and U5928 (N_5928,N_3909,N_216);
or U5929 (N_5929,N_1780,N_4723);
and U5930 (N_5930,N_2688,N_4282);
nand U5931 (N_5931,N_2378,N_4278);
and U5932 (N_5932,N_1943,N_4849);
or U5933 (N_5933,N_3530,N_319);
nand U5934 (N_5934,N_3288,N_1792);
or U5935 (N_5935,N_4200,N_1749);
and U5936 (N_5936,N_3203,N_4165);
nor U5937 (N_5937,N_729,N_2494);
nand U5938 (N_5938,N_3660,N_3531);
and U5939 (N_5939,N_3615,N_3907);
nand U5940 (N_5940,N_4238,N_2224);
xor U5941 (N_5941,N_3704,N_2152);
xor U5942 (N_5942,N_4615,N_1540);
nor U5943 (N_5943,N_2920,N_566);
nand U5944 (N_5944,N_4580,N_4995);
nand U5945 (N_5945,N_771,N_2244);
nand U5946 (N_5946,N_1700,N_1338);
nand U5947 (N_5947,N_3793,N_2835);
and U5948 (N_5948,N_1044,N_468);
or U5949 (N_5949,N_1828,N_1809);
nor U5950 (N_5950,N_2711,N_1013);
xor U5951 (N_5951,N_3575,N_3673);
and U5952 (N_5952,N_1488,N_1755);
and U5953 (N_5953,N_1285,N_3915);
nand U5954 (N_5954,N_46,N_4037);
nand U5955 (N_5955,N_2652,N_4311);
xnor U5956 (N_5956,N_3863,N_4393);
and U5957 (N_5957,N_2807,N_3569);
nand U5958 (N_5958,N_3370,N_4300);
and U5959 (N_5959,N_1966,N_4636);
and U5960 (N_5960,N_1948,N_2342);
nand U5961 (N_5961,N_733,N_3121);
or U5962 (N_5962,N_2079,N_1375);
and U5963 (N_5963,N_4488,N_3762);
and U5964 (N_5964,N_918,N_478);
nor U5965 (N_5965,N_490,N_2659);
nand U5966 (N_5966,N_2069,N_3349);
nor U5967 (N_5967,N_4540,N_3452);
nor U5968 (N_5968,N_3960,N_4826);
and U5969 (N_5969,N_135,N_1045);
nor U5970 (N_5970,N_263,N_4655);
and U5971 (N_5971,N_4192,N_894);
nand U5972 (N_5972,N_3091,N_664);
nor U5973 (N_5973,N_2680,N_391);
nor U5974 (N_5974,N_4181,N_655);
nand U5975 (N_5975,N_4317,N_3130);
nand U5976 (N_5976,N_127,N_2327);
nand U5977 (N_5977,N_2000,N_1647);
or U5978 (N_5978,N_4444,N_2658);
nor U5979 (N_5979,N_2050,N_1002);
or U5980 (N_5980,N_1616,N_940);
xor U5981 (N_5981,N_2157,N_543);
and U5982 (N_5982,N_3082,N_605);
or U5983 (N_5983,N_1308,N_2119);
or U5984 (N_5984,N_2699,N_3078);
and U5985 (N_5985,N_3123,N_595);
and U5986 (N_5986,N_4137,N_4913);
or U5987 (N_5987,N_4396,N_3199);
nor U5988 (N_5988,N_483,N_4016);
or U5989 (N_5989,N_3904,N_4021);
nor U5990 (N_5990,N_2208,N_3128);
and U5991 (N_5991,N_4343,N_4714);
or U5992 (N_5992,N_3032,N_3095);
and U5993 (N_5993,N_1279,N_2615);
nand U5994 (N_5994,N_633,N_1944);
and U5995 (N_5995,N_3928,N_2969);
or U5996 (N_5996,N_2072,N_3308);
or U5997 (N_5997,N_3788,N_4266);
nand U5998 (N_5998,N_2287,N_587);
and U5999 (N_5999,N_1625,N_510);
xnor U6000 (N_6000,N_1703,N_4755);
nand U6001 (N_6001,N_3343,N_375);
and U6002 (N_6002,N_4881,N_686);
or U6003 (N_6003,N_2709,N_653);
or U6004 (N_6004,N_3265,N_2590);
and U6005 (N_6005,N_1909,N_960);
nor U6006 (N_6006,N_682,N_2938);
or U6007 (N_6007,N_1964,N_817);
xor U6008 (N_6008,N_1313,N_3038);
nand U6009 (N_6009,N_3609,N_2124);
or U6010 (N_6010,N_4261,N_43);
nand U6011 (N_6011,N_416,N_71);
nand U6012 (N_6012,N_3233,N_87);
nor U6013 (N_6013,N_3469,N_1185);
and U6014 (N_6014,N_3938,N_2106);
and U6015 (N_6015,N_4600,N_4560);
or U6016 (N_6016,N_1963,N_3039);
nor U6017 (N_6017,N_176,N_1621);
and U6018 (N_6018,N_4884,N_730);
and U6019 (N_6019,N_2621,N_4374);
and U6020 (N_6020,N_2059,N_3812);
nand U6021 (N_6021,N_4895,N_1788);
or U6022 (N_6022,N_2775,N_2510);
xnor U6023 (N_6023,N_3570,N_1619);
or U6024 (N_6024,N_1615,N_4119);
or U6025 (N_6025,N_3871,N_1295);
and U6026 (N_6026,N_523,N_2813);
or U6027 (N_6027,N_1267,N_2726);
nor U6028 (N_6028,N_3827,N_2727);
and U6029 (N_6029,N_426,N_1263);
nor U6030 (N_6030,N_4547,N_3488);
or U6031 (N_6031,N_1765,N_1377);
or U6032 (N_6032,N_4342,N_1098);
nand U6033 (N_6033,N_3954,N_4719);
and U6034 (N_6034,N_4041,N_300);
and U6035 (N_6035,N_2353,N_4740);
nor U6036 (N_6036,N_2641,N_3809);
and U6037 (N_6037,N_1133,N_635);
nand U6038 (N_6038,N_3429,N_1264);
and U6039 (N_6039,N_3815,N_3459);
nor U6040 (N_6040,N_2796,N_3230);
nor U6041 (N_6041,N_4992,N_3269);
nor U6042 (N_6042,N_2309,N_4677);
or U6043 (N_6043,N_4341,N_1477);
or U6044 (N_6044,N_1620,N_1520);
nand U6045 (N_6045,N_4528,N_4862);
and U6046 (N_6046,N_861,N_4700);
nand U6047 (N_6047,N_735,N_3721);
and U6048 (N_6048,N_780,N_3945);
nand U6049 (N_6049,N_1493,N_198);
or U6050 (N_6050,N_4447,N_4421);
nand U6051 (N_6051,N_3260,N_3601);
nor U6052 (N_6052,N_1155,N_3068);
and U6053 (N_6053,N_2547,N_528);
and U6054 (N_6054,N_367,N_1782);
nor U6055 (N_6055,N_1551,N_3063);
and U6056 (N_6056,N_1333,N_4386);
nor U6057 (N_6057,N_2654,N_3401);
or U6058 (N_6058,N_4603,N_2418);
nor U6059 (N_6059,N_1768,N_2743);
xor U6060 (N_6060,N_1400,N_3652);
nand U6061 (N_6061,N_3158,N_641);
and U6062 (N_6062,N_1552,N_2572);
nor U6063 (N_6063,N_688,N_3392);
xor U6064 (N_6064,N_41,N_1217);
nor U6065 (N_6065,N_111,N_178);
or U6066 (N_6066,N_3934,N_1173);
xor U6067 (N_6067,N_3391,N_4020);
nor U6068 (N_6068,N_76,N_1031);
xor U6069 (N_6069,N_1845,N_4648);
nor U6070 (N_6070,N_1305,N_2780);
nor U6071 (N_6071,N_4214,N_3328);
or U6072 (N_6072,N_2206,N_3545);
or U6073 (N_6073,N_323,N_986);
xnor U6074 (N_6074,N_1923,N_1698);
and U6075 (N_6075,N_1769,N_1569);
nor U6076 (N_6076,N_1135,N_2645);
xnor U6077 (N_6077,N_1369,N_4036);
and U6078 (N_6078,N_387,N_4715);
and U6079 (N_6079,N_2042,N_1694);
xor U6080 (N_6080,N_1277,N_3400);
and U6081 (N_6081,N_1776,N_2902);
and U6082 (N_6082,N_2925,N_441);
nand U6083 (N_6083,N_59,N_3234);
and U6084 (N_6084,N_637,N_4051);
xor U6085 (N_6085,N_3293,N_1247);
nand U6086 (N_6086,N_4039,N_3310);
or U6087 (N_6087,N_4480,N_2868);
or U6088 (N_6088,N_4955,N_2357);
xnor U6089 (N_6089,N_3345,N_4066);
xnor U6090 (N_6090,N_3520,N_4024);
or U6091 (N_6091,N_851,N_978);
and U6092 (N_6092,N_4446,N_3473);
nor U6093 (N_6093,N_3116,N_2369);
xor U6094 (N_6094,N_4436,N_4586);
nor U6095 (N_6095,N_3905,N_1107);
xor U6096 (N_6096,N_1420,N_2631);
and U6097 (N_6097,N_3104,N_3882);
or U6098 (N_6098,N_4601,N_2944);
and U6099 (N_6099,N_2764,N_4085);
and U6100 (N_6100,N_4757,N_2875);
and U6101 (N_6101,N_4801,N_1942);
xnor U6102 (N_6102,N_631,N_3432);
and U6103 (N_6103,N_4115,N_943);
nor U6104 (N_6104,N_1084,N_969);
or U6105 (N_6105,N_1824,N_685);
or U6106 (N_6106,N_2577,N_3410);
and U6107 (N_6107,N_2315,N_4384);
or U6108 (N_6108,N_1171,N_1007);
and U6109 (N_6109,N_533,N_394);
or U6110 (N_6110,N_2298,N_3752);
or U6111 (N_6111,N_2409,N_2910);
nand U6112 (N_6112,N_693,N_2977);
nor U6113 (N_6113,N_3883,N_1288);
nor U6114 (N_6114,N_2632,N_2026);
and U6115 (N_6115,N_3770,N_1575);
and U6116 (N_6116,N_4483,N_2018);
and U6117 (N_6117,N_3155,N_130);
xor U6118 (N_6118,N_1861,N_3892);
and U6119 (N_6119,N_570,N_3557);
or U6120 (N_6120,N_3676,N_1147);
nand U6121 (N_6121,N_3780,N_4127);
nor U6122 (N_6122,N_4098,N_321);
or U6123 (N_6123,N_3538,N_796);
nand U6124 (N_6124,N_695,N_3847);
nand U6125 (N_6125,N_4022,N_184);
nand U6126 (N_6126,N_1352,N_2306);
and U6127 (N_6127,N_476,N_1675);
and U6128 (N_6128,N_186,N_1139);
nand U6129 (N_6129,N_2098,N_4437);
and U6130 (N_6130,N_1818,N_4008);
nor U6131 (N_6131,N_3542,N_2025);
or U6132 (N_6132,N_3154,N_4090);
nor U6133 (N_6133,N_3435,N_3884);
nand U6134 (N_6134,N_1543,N_3205);
nand U6135 (N_6135,N_2554,N_4930);
or U6136 (N_6136,N_2717,N_1514);
or U6137 (N_6137,N_1613,N_3358);
or U6138 (N_6138,N_1882,N_4830);
and U6139 (N_6139,N_1110,N_2568);
and U6140 (N_6140,N_2978,N_2846);
nand U6141 (N_6141,N_904,N_2988);
nand U6142 (N_6142,N_1362,N_2128);
nand U6143 (N_6143,N_3096,N_419);
nor U6144 (N_6144,N_4247,N_2897);
or U6145 (N_6145,N_3182,N_98);
and U6146 (N_6146,N_2076,N_259);
or U6147 (N_6147,N_3983,N_4061);
nand U6148 (N_6148,N_2964,N_3023);
or U6149 (N_6149,N_3357,N_1717);
or U6150 (N_6150,N_450,N_1527);
nand U6151 (N_6151,N_4696,N_56);
or U6152 (N_6152,N_4817,N_1497);
xnor U6153 (N_6153,N_1395,N_1417);
xnor U6154 (N_6154,N_2623,N_322);
or U6155 (N_6155,N_2328,N_3654);
and U6156 (N_6156,N_727,N_1638);
nor U6157 (N_6157,N_2526,N_3564);
and U6158 (N_6158,N_2217,N_1713);
and U6159 (N_6159,N_2043,N_3009);
nand U6160 (N_6160,N_1778,N_1405);
nand U6161 (N_6161,N_1131,N_3115);
or U6162 (N_6162,N_743,N_4459);
and U6163 (N_6163,N_2965,N_2325);
nor U6164 (N_6164,N_3414,N_1472);
nor U6165 (N_6165,N_763,N_2252);
or U6166 (N_6166,N_2385,N_3957);
and U6167 (N_6167,N_3785,N_1328);
xor U6168 (N_6168,N_2340,N_2929);
xor U6169 (N_6169,N_2219,N_3539);
nor U6170 (N_6170,N_781,N_1723);
nor U6171 (N_6171,N_1057,N_2710);
nor U6172 (N_6172,N_2733,N_1349);
nand U6173 (N_6173,N_4010,N_2390);
nand U6174 (N_6174,N_645,N_2596);
nor U6175 (N_6175,N_3908,N_2117);
nor U6176 (N_6176,N_4900,N_1550);
nor U6177 (N_6177,N_2350,N_2533);
and U6178 (N_6178,N_2486,N_2546);
nor U6179 (N_6179,N_1919,N_2431);
xnor U6180 (N_6180,N_1322,N_1159);
nor U6181 (N_6181,N_2302,N_4597);
or U6182 (N_6182,N_3886,N_1743);
or U6183 (N_6183,N_2930,N_2679);
nand U6184 (N_6184,N_22,N_1074);
or U6185 (N_6185,N_2197,N_1995);
or U6186 (N_6186,N_4417,N_223);
or U6187 (N_6187,N_2644,N_423);
nand U6188 (N_6188,N_3360,N_660);
and U6189 (N_6189,N_4563,N_2249);
nand U6190 (N_6190,N_3625,N_4654);
or U6191 (N_6191,N_1815,N_49);
nand U6192 (N_6192,N_1897,N_1628);
nor U6193 (N_6193,N_4935,N_3301);
and U6194 (N_6194,N_1113,N_718);
nor U6195 (N_6195,N_1666,N_2564);
nand U6196 (N_6196,N_1386,N_1915);
nor U6197 (N_6197,N_3191,N_274);
nor U6198 (N_6198,N_3771,N_4738);
or U6199 (N_6199,N_1763,N_3187);
nor U6200 (N_6200,N_4326,N_4769);
nand U6201 (N_6201,N_3565,N_1302);
and U6202 (N_6202,N_1151,N_4842);
nor U6203 (N_6203,N_2722,N_217);
nand U6204 (N_6204,N_4539,N_4429);
nand U6205 (N_6205,N_3327,N_3081);
or U6206 (N_6206,N_1408,N_37);
nand U6207 (N_6207,N_376,N_4888);
nand U6208 (N_6208,N_2407,N_2651);
and U6209 (N_6209,N_3854,N_2479);
xor U6210 (N_6210,N_48,N_447);
nand U6211 (N_6211,N_2694,N_1733);
and U6212 (N_6212,N_2184,N_1289);
nand U6213 (N_6213,N_4585,N_1512);
and U6214 (N_6214,N_1931,N_3782);
xnor U6215 (N_6215,N_2600,N_2848);
and U6216 (N_6216,N_4556,N_4454);
nor U6217 (N_6217,N_1643,N_467);
or U6218 (N_6218,N_712,N_4731);
nor U6219 (N_6219,N_4790,N_4530);
or U6220 (N_6220,N_3075,N_1499);
nor U6221 (N_6221,N_1149,N_1981);
and U6222 (N_6222,N_2719,N_297);
or U6223 (N_6223,N_1060,N_3800);
nand U6224 (N_6224,N_3526,N_1005);
nand U6225 (N_6225,N_3603,N_3872);
nand U6226 (N_6226,N_53,N_3532);
and U6227 (N_6227,N_2020,N_2575);
xnor U6228 (N_6228,N_199,N_4321);
nand U6229 (N_6229,N_991,N_4762);
nand U6230 (N_6230,N_2560,N_2876);
xor U6231 (N_6231,N_1201,N_513);
xor U6232 (N_6232,N_2664,N_1241);
nor U6233 (N_6233,N_4057,N_3631);
nand U6234 (N_6234,N_4235,N_4896);
and U6235 (N_6235,N_2256,N_728);
and U6236 (N_6236,N_4574,N_2511);
or U6237 (N_6237,N_2836,N_2432);
nor U6238 (N_6238,N_601,N_3420);
and U6239 (N_6239,N_4576,N_3868);
xnor U6240 (N_6240,N_3244,N_2299);
nor U6241 (N_6241,N_4503,N_1389);
nor U6242 (N_6242,N_2911,N_1937);
or U6243 (N_6243,N_396,N_3300);
or U6244 (N_6244,N_4878,N_1371);
nor U6245 (N_6245,N_798,N_1049);
nor U6246 (N_6246,N_2008,N_579);
nor U6247 (N_6247,N_2650,N_3684);
and U6248 (N_6248,N_27,N_2288);
nor U6249 (N_6249,N_4746,N_4917);
or U6250 (N_6250,N_844,N_3519);
nor U6251 (N_6251,N_1904,N_555);
xor U6252 (N_6252,N_3740,N_4153);
nor U6253 (N_6253,N_4810,N_1470);
xnor U6254 (N_6254,N_2886,N_698);
xnor U6255 (N_6255,N_4170,N_2400);
nand U6256 (N_6256,N_1012,N_1209);
nor U6257 (N_6257,N_1536,N_4841);
xnor U6258 (N_6258,N_638,N_327);
nand U6259 (N_6259,N_4705,N_2051);
or U6260 (N_6260,N_4741,N_4473);
or U6261 (N_6261,N_386,N_3347);
nor U6262 (N_6262,N_2233,N_4277);
or U6263 (N_6263,N_339,N_1907);
nor U6264 (N_6264,N_4344,N_4460);
or U6265 (N_6265,N_4068,N_2667);
xnor U6266 (N_6266,N_4855,N_3966);
nor U6267 (N_6267,N_4045,N_2462);
nand U6268 (N_6268,N_1985,N_4578);
xor U6269 (N_6269,N_1662,N_162);
nand U6270 (N_6270,N_2993,N_1669);
or U6271 (N_6271,N_95,N_4555);
nand U6272 (N_6272,N_4796,N_2529);
or U6273 (N_6273,N_1024,N_4405);
xnor U6274 (N_6274,N_3860,N_3041);
nor U6275 (N_6275,N_4784,N_4236);
nand U6276 (N_6276,N_3477,N_1838);
nor U6277 (N_6277,N_3986,N_384);
nor U6278 (N_6278,N_3887,N_4991);
xor U6279 (N_6279,N_2236,N_1331);
or U6280 (N_6280,N_1917,N_3371);
nor U6281 (N_6281,N_3225,N_3132);
or U6282 (N_6282,N_3072,N_1654);
and U6283 (N_6283,N_2655,N_494);
nand U6284 (N_6284,N_3113,N_2703);
nand U6285 (N_6285,N_2759,N_472);
nor U6286 (N_6286,N_4293,N_1475);
nor U6287 (N_6287,N_1112,N_4515);
or U6288 (N_6288,N_1851,N_2597);
and U6289 (N_6289,N_3241,N_4695);
or U6290 (N_6290,N_4844,N_3178);
or U6291 (N_6291,N_4592,N_1450);
xor U6292 (N_6292,N_926,N_4581);
and U6293 (N_6293,N_2279,N_4086);
nor U6294 (N_6294,N_4818,N_2675);
and U6295 (N_6295,N_409,N_756);
and U6296 (N_6296,N_1495,N_1416);
nor U6297 (N_6297,N_481,N_746);
and U6298 (N_6298,N_3761,N_3751);
and U6299 (N_6299,N_2689,N_4449);
and U6300 (N_6300,N_3726,N_3580);
xnor U6301 (N_6301,N_1605,N_3791);
nand U6302 (N_6302,N_4310,N_4643);
and U6303 (N_6303,N_1987,N_1762);
nor U6304 (N_6304,N_2839,N_4312);
nor U6305 (N_6305,N_3964,N_4328);
and U6306 (N_6306,N_2199,N_363);
and U6307 (N_6307,N_3292,N_517);
and U6308 (N_6308,N_173,N_2326);
nand U6309 (N_6309,N_1268,N_471);
and U6310 (N_6310,N_207,N_209);
nand U6311 (N_6311,N_3136,N_668);
or U6312 (N_6312,N_2495,N_4734);
or U6313 (N_6313,N_1630,N_3416);
nand U6314 (N_6314,N_90,N_4160);
or U6315 (N_6315,N_4209,N_4487);
or U6316 (N_6316,N_66,N_1081);
and U6317 (N_6317,N_77,N_2612);
or U6318 (N_6318,N_304,N_203);
and U6319 (N_6319,N_2541,N_1188);
nor U6320 (N_6320,N_1260,N_1739);
or U6321 (N_6321,N_3456,N_229);
or U6322 (N_6322,N_933,N_1170);
nor U6323 (N_6323,N_174,N_689);
nand U6324 (N_6324,N_551,N_1508);
and U6325 (N_6325,N_1681,N_4921);
xnor U6326 (N_6326,N_3748,N_1866);
and U6327 (N_6327,N_1933,N_3074);
and U6328 (N_6328,N_4710,N_1237);
xor U6329 (N_6329,N_3837,N_4863);
nor U6330 (N_6330,N_2551,N_2331);
xnor U6331 (N_6331,N_4389,N_3889);
nand U6332 (N_6332,N_2232,N_3334);
nor U6333 (N_6333,N_2065,N_4340);
or U6334 (N_6334,N_3627,N_4960);
nand U6335 (N_6335,N_4754,N_4832);
and U6336 (N_6336,N_2725,N_3963);
xor U6337 (N_6337,N_4668,N_3978);
and U6338 (N_6338,N_344,N_514);
and U6339 (N_6339,N_1745,N_4732);
nor U6340 (N_6340,N_3303,N_680);
and U6341 (N_6341,N_2906,N_3758);
or U6342 (N_6342,N_2456,N_2230);
nand U6343 (N_6343,N_1636,N_2492);
nand U6344 (N_6344,N_2030,N_1399);
nand U6345 (N_6345,N_3528,N_4471);
or U6346 (N_6346,N_931,N_2426);
or U6347 (N_6347,N_3624,N_4708);
or U6348 (N_6348,N_1916,N_238);
or U6349 (N_6349,N_2057,N_134);
nor U6350 (N_6350,N_3712,N_4775);
nor U6351 (N_6351,N_531,N_1435);
and U6352 (N_6352,N_3715,N_4867);
xor U6353 (N_6353,N_2196,N_2103);
or U6354 (N_6354,N_2985,N_1365);
or U6355 (N_6355,N_2856,N_12);
nor U6356 (N_6356,N_1396,N_4055);
nor U6357 (N_6357,N_133,N_3781);
nor U6358 (N_6358,N_600,N_3280);
or U6359 (N_6359,N_2423,N_869);
nand U6360 (N_6360,N_4220,N_2943);
nand U6361 (N_6361,N_842,N_3333);
and U6362 (N_6362,N_1634,N_1473);
xor U6363 (N_6363,N_1570,N_4883);
or U6364 (N_6364,N_1817,N_2566);
nor U6365 (N_6365,N_2599,N_959);
or U6366 (N_6366,N_538,N_4332);
or U6367 (N_6367,N_3161,N_4279);
or U6368 (N_6368,N_1829,N_2757);
xnor U6369 (N_6369,N_4368,N_3992);
or U6370 (N_6370,N_2950,N_4772);
nand U6371 (N_6371,N_3493,N_4073);
nand U6372 (N_6372,N_316,N_4988);
or U6373 (N_6373,N_4725,N_3779);
xnor U6374 (N_6374,N_2974,N_2424);
and U6375 (N_6375,N_927,N_1016);
and U6376 (N_6376,N_4924,N_1781);
or U6377 (N_6377,N_2506,N_3359);
nand U6378 (N_6378,N_17,N_2237);
nand U6379 (N_6379,N_237,N_985);
nor U6380 (N_6380,N_2517,N_1752);
and U6381 (N_6381,N_3563,N_3080);
and U6382 (N_6382,N_204,N_3572);
or U6383 (N_6383,N_629,N_4785);
nor U6384 (N_6384,N_1803,N_3184);
xor U6385 (N_6385,N_4966,N_4593);
nor U6386 (N_6386,N_2914,N_2528);
or U6387 (N_6387,N_1390,N_1040);
or U6388 (N_6388,N_983,N_830);
nor U6389 (N_6389,N_2913,N_4179);
nor U6390 (N_6390,N_449,N_258);
or U6391 (N_6391,N_1754,N_2368);
and U6392 (N_6392,N_4156,N_2277);
nand U6393 (N_6393,N_4952,N_977);
or U6394 (N_6394,N_47,N_1775);
nand U6395 (N_6395,N_4640,N_1925);
and U6396 (N_6396,N_3535,N_526);
and U6397 (N_6397,N_4981,N_1892);
nand U6398 (N_6398,N_512,N_1665);
or U6399 (N_6399,N_2961,N_3533);
and U6400 (N_6400,N_3110,N_4922);
nor U6401 (N_6401,N_3356,N_1650);
and U6402 (N_6402,N_3365,N_3471);
and U6403 (N_6403,N_1554,N_4225);
and U6404 (N_6404,N_2809,N_3378);
or U6405 (N_6405,N_2799,N_1230);
nand U6406 (N_6406,N_2223,N_3135);
nor U6407 (N_6407,N_1446,N_4427);
nor U6408 (N_6408,N_2422,N_4363);
and U6409 (N_6409,N_4680,N_953);
and U6410 (N_6410,N_354,N_979);
or U6411 (N_6411,N_3153,N_1505);
nand U6412 (N_6412,N_4167,N_3494);
nand U6413 (N_6413,N_4331,N_3850);
nand U6414 (N_6414,N_4280,N_3536);
or U6415 (N_6415,N_1066,N_3789);
nor U6416 (N_6416,N_4149,N_4946);
nand U6417 (N_6417,N_469,N_3602);
xor U6418 (N_6418,N_3454,N_2607);
and U6419 (N_6419,N_1704,N_3839);
and U6420 (N_6420,N_1668,N_318);
nand U6421 (N_6421,N_2198,N_2457);
nor U6422 (N_6422,N_2012,N_3747);
nor U6423 (N_6423,N_2213,N_1402);
nand U6424 (N_6424,N_2203,N_359);
xor U6425 (N_6425,N_3814,N_1633);
nor U6426 (N_6426,N_4252,N_550);
and U6427 (N_6427,N_1672,N_4583);
and U6428 (N_6428,N_4216,N_777);
and U6429 (N_6429,N_1303,N_3683);
xnor U6430 (N_6430,N_2092,N_1215);
nor U6431 (N_6431,N_188,N_2314);
xnor U6432 (N_6432,N_4313,N_1969);
nor U6433 (N_6433,N_3398,N_3399);
and U6434 (N_6434,N_118,N_4814);
and U6435 (N_6435,N_3085,N_4411);
and U6436 (N_6436,N_589,N_1522);
or U6437 (N_6437,N_2624,N_2270);
nand U6438 (N_6438,N_3376,N_4687);
nor U6439 (N_6439,N_1918,N_3395);
nand U6440 (N_6440,N_3185,N_4678);
nor U6441 (N_6441,N_4618,N_1162);
xor U6442 (N_6442,N_266,N_3507);
nor U6443 (N_6443,N_1415,N_2608);
and U6444 (N_6444,N_85,N_2015);
nand U6445 (N_6445,N_3505,N_225);
xnor U6446 (N_6446,N_2384,N_4807);
or U6447 (N_6447,N_946,N_2530);
and U6448 (N_6448,N_1062,N_4150);
or U6449 (N_6449,N_3632,N_4360);
nor U6450 (N_6450,N_751,N_2698);
and U6451 (N_6451,N_2242,N_4320);
xnor U6452 (N_6452,N_4699,N_2957);
nand U6453 (N_6453,N_649,N_1899);
nor U6454 (N_6454,N_1712,N_254);
nand U6455 (N_6455,N_2693,N_2519);
or U6456 (N_6456,N_1210,N_3719);
or U6457 (N_6457,N_2417,N_3540);
nand U6458 (N_6458,N_3428,N_1856);
nor U6459 (N_6459,N_2831,N_776);
or U6460 (N_6460,N_3965,N_4852);
xor U6461 (N_6461,N_1568,N_2064);
or U6462 (N_6462,N_4607,N_3336);
nor U6463 (N_6463,N_502,N_2441);
and U6464 (N_6464,N_3206,N_4783);
or U6465 (N_6465,N_2563,N_2286);
nand U6466 (N_6466,N_1244,N_2359);
nor U6467 (N_6467,N_2083,N_3722);
nor U6468 (N_6468,N_3342,N_222);
and U6469 (N_6469,N_3138,N_1225);
and U6470 (N_6470,N_1271,N_760);
nor U6471 (N_6471,N_2278,N_4187);
nand U6472 (N_6472,N_2387,N_4069);
xnor U6473 (N_6473,N_2909,N_4364);
or U6474 (N_6474,N_3629,N_1172);
nor U6475 (N_6475,N_498,N_971);
nor U6476 (N_6476,N_2803,N_3749);
nand U6477 (N_6477,N_3374,N_2508);
and U6478 (N_6478,N_941,N_1979);
xor U6479 (N_6479,N_452,N_1935);
nand U6480 (N_6480,N_2087,N_3502);
nand U6481 (N_6481,N_2099,N_126);
or U6482 (N_6482,N_3235,N_2745);
xor U6483 (N_6483,N_282,N_1462);
and U6484 (N_6484,N_3952,N_1168);
nand U6485 (N_6485,N_955,N_278);
nand U6486 (N_6486,N_4038,N_3217);
and U6487 (N_6487,N_937,N_4052);
or U6488 (N_6488,N_4646,N_652);
nand U6489 (N_6489,N_1584,N_1348);
nand U6490 (N_6490,N_3669,N_1234);
xnor U6491 (N_6491,N_3024,N_1960);
and U6492 (N_6492,N_2148,N_3022);
nand U6493 (N_6493,N_3818,N_1585);
nor U6494 (N_6494,N_2521,N_1640);
nand U6495 (N_6495,N_2370,N_1601);
nand U6496 (N_6496,N_3742,N_4189);
nor U6497 (N_6497,N_1136,N_2696);
nor U6498 (N_6498,N_3644,N_4926);
nor U6499 (N_6499,N_3504,N_3806);
and U6500 (N_6500,N_2120,N_1878);
and U6501 (N_6501,N_3323,N_1526);
or U6502 (N_6502,N_3387,N_411);
nand U6503 (N_6503,N_3582,N_1069);
or U6504 (N_6504,N_3226,N_1823);
or U6505 (N_6505,N_1101,N_4937);
nand U6506 (N_6506,N_2038,N_1912);
or U6507 (N_6507,N_3846,N_4423);
or U6508 (N_6508,N_2576,N_2952);
and U6509 (N_6509,N_1822,N_1820);
xor U6510 (N_6510,N_1476,N_524);
or U6511 (N_6511,N_3438,N_811);
and U6512 (N_6512,N_1287,N_1306);
nor U6513 (N_6513,N_3737,N_4148);
and U6514 (N_6514,N_460,N_381);
nor U6515 (N_6515,N_1075,N_4408);
nand U6516 (N_6516,N_2027,N_1093);
and U6517 (N_6517,N_1078,N_2513);
nand U6518 (N_6518,N_1555,N_1770);
nand U6519 (N_6519,N_2731,N_1445);
nor U6520 (N_6520,N_1335,N_4979);
and U6521 (N_6521,N_3592,N_3655);
xor U6522 (N_6522,N_4011,N_3324);
or U6523 (N_6523,N_2847,N_564);
and U6524 (N_6524,N_4612,N_572);
or U6525 (N_6525,N_3824,N_3914);
nand U6526 (N_6526,N_1959,N_1724);
or U6527 (N_6527,N_3481,N_835);
nand U6528 (N_6528,N_4780,N_101);
and U6529 (N_6529,N_4865,N_2345);
nor U6530 (N_6530,N_1702,N_3813);
and U6531 (N_6531,N_2502,N_4839);
nor U6532 (N_6532,N_1048,N_3201);
xor U6533 (N_6533,N_4886,N_1660);
nor U6534 (N_6534,N_370,N_4250);
and U6535 (N_6535,N_1028,N_3585);
xnor U6536 (N_6536,N_2874,N_3853);
and U6537 (N_6537,N_3946,N_4712);
nor U6538 (N_6538,N_137,N_3086);
and U6539 (N_6539,N_3981,N_4957);
nand U6540 (N_6540,N_1316,N_2215);
and U6541 (N_6541,N_876,N_2391);
nand U6542 (N_6542,N_4685,N_4972);
or U6543 (N_6543,N_2669,N_2583);
and U6544 (N_6544,N_996,N_4335);
and U6545 (N_6545,N_4511,N_4486);
and U6546 (N_6546,N_1307,N_1455);
and U6547 (N_6547,N_724,N_4764);
xnor U6548 (N_6548,N_4779,N_3772);
xnor U6549 (N_6549,N_2995,N_2677);
nand U6550 (N_6550,N_1537,N_2959);
or U6551 (N_6551,N_1790,N_833);
or U6552 (N_6552,N_1992,N_2193);
nor U6553 (N_6553,N_2346,N_1320);
nand U6554 (N_6554,N_346,N_3495);
nor U6555 (N_6555,N_3326,N_878);
nor U6556 (N_6556,N_569,N_4362);
xor U6557 (N_6557,N_159,N_4518);
and U6558 (N_6558,N_3594,N_4688);
nand U6559 (N_6559,N_4506,N_1443);
nand U6560 (N_6560,N_3163,N_2093);
and U6561 (N_6561,N_255,N_1122);
nor U6562 (N_6562,N_1532,N_1104);
nor U6563 (N_6563,N_3893,N_1734);
nor U6564 (N_6564,N_3596,N_2420);
and U6565 (N_6565,N_3980,N_1283);
nor U6566 (N_6566,N_625,N_2333);
nor U6567 (N_6567,N_827,N_536);
or U6568 (N_6568,N_4392,N_1124);
or U6569 (N_6569,N_2746,N_2188);
nand U6570 (N_6570,N_3012,N_3417);
nand U6571 (N_6571,N_2797,N_5);
and U6572 (N_6572,N_592,N_3927);
xor U6573 (N_6573,N_3237,N_1208);
and U6574 (N_6574,N_4462,N_4866);
nand U6575 (N_6575,N_3208,N_1701);
and U6576 (N_6576,N_3298,N_615);
or U6577 (N_6577,N_4623,N_3929);
nor U6578 (N_6578,N_604,N_4301);
or U6579 (N_6579,N_1673,N_4923);
and U6580 (N_6580,N_3544,N_880);
nand U6581 (N_6581,N_558,N_4397);
xnor U6582 (N_6582,N_2090,N_1026);
nand U6583 (N_6583,N_1413,N_3380);
nand U6584 (N_6584,N_4596,N_2211);
nand U6585 (N_6585,N_3943,N_79);
nand U6586 (N_6586,N_1150,N_70);
nor U6587 (N_6587,N_2313,N_456);
and U6588 (N_6588,N_2795,N_2111);
or U6589 (N_6589,N_750,N_4827);
and U6590 (N_6590,N_2532,N_738);
or U6591 (N_6591,N_2395,N_1951);
and U6592 (N_6592,N_4918,N_1850);
or U6593 (N_6593,N_2832,N_151);
or U6594 (N_6594,N_3729,N_152);
nor U6595 (N_6595,N_3728,N_4211);
and U6596 (N_6596,N_4091,N_2396);
nand U6597 (N_6597,N_309,N_2773);
nand U6598 (N_6598,N_3857,N_1050);
and U6599 (N_6599,N_267,N_239);
and U6600 (N_6600,N_1688,N_2857);
and U6601 (N_6601,N_704,N_4176);
nand U6602 (N_6602,N_114,N_758);
nand U6603 (N_6603,N_281,N_1080);
nand U6604 (N_6604,N_1439,N_461);
and U6605 (N_6605,N_4965,N_4474);
and U6606 (N_6606,N_4631,N_1017);
and U6607 (N_6607,N_2893,N_4435);
or U6608 (N_6608,N_1816,N_1011);
and U6609 (N_6609,N_1255,N_715);
nor U6610 (N_6610,N_3263,N_4641);
or U6611 (N_6611,N_2228,N_790);
nor U6612 (N_6612,N_3377,N_1258);
xnor U6613 (N_6613,N_2984,N_1599);
and U6614 (N_6614,N_4359,N_1814);
or U6615 (N_6615,N_3167,N_2154);
or U6616 (N_6616,N_3145,N_1805);
nor U6617 (N_6617,N_2190,N_1105);
nand U6618 (N_6618,N_726,N_1191);
nand U6619 (N_6619,N_1589,N_3933);
nor U6620 (N_6620,N_3166,N_1973);
nor U6621 (N_6621,N_4499,N_1);
nand U6622 (N_6622,N_3873,N_2558);
and U6623 (N_6623,N_546,N_3798);
nor U6624 (N_6624,N_3607,N_3150);
nand U6625 (N_6625,N_3367,N_4428);
and U6626 (N_6626,N_1474,N_3369);
nand U6627 (N_6627,N_4624,N_2238);
nand U6628 (N_6628,N_4532,N_4412);
nand U6629 (N_6629,N_360,N_4161);
xor U6630 (N_6630,N_1444,N_1359);
or U6631 (N_6631,N_3423,N_74);
nand U6632 (N_6632,N_311,N_1839);
or U6633 (N_6633,N_591,N_1465);
nand U6634 (N_6634,N_1239,N_2112);
nor U6635 (N_6635,N_242,N_1678);
xnor U6636 (N_6636,N_2766,N_4249);
nand U6637 (N_6637,N_132,N_3578);
or U6638 (N_6638,N_1487,N_866);
or U6639 (N_6639,N_1988,N_248);
and U6640 (N_6640,N_2768,N_457);
nand U6641 (N_6641,N_4527,N_1751);
and U6642 (N_6642,N_3016,N_4609);
or U6643 (N_6643,N_2801,N_4838);
or U6644 (N_6644,N_3595,N_4948);
or U6645 (N_6645,N_4890,N_94);
and U6646 (N_6646,N_1658,N_1033);
nor U6647 (N_6647,N_4570,N_373);
and U6648 (N_6648,N_1079,N_1774);
xor U6649 (N_6649,N_1025,N_3717);
xor U6650 (N_6650,N_1158,N_2559);
xnor U6651 (N_6651,N_1579,N_2579);
nor U6652 (N_6652,N_2014,N_4651);
nor U6653 (N_6653,N_2459,N_2234);
xor U6654 (N_6654,N_3189,N_1791);
or U6655 (N_6655,N_3935,N_1872);
nor U6656 (N_6656,N_2216,N_740);
or U6657 (N_6657,N_3970,N_2001);
and U6658 (N_6658,N_1846,N_3924);
and U6659 (N_6659,N_976,N_2068);
nor U6660 (N_6660,N_189,N_2916);
and U6661 (N_6661,N_4006,N_966);
or U6662 (N_6662,N_4130,N_2415);
nand U6663 (N_6663,N_2543,N_4164);
nand U6664 (N_6664,N_4075,N_2162);
nand U6665 (N_6665,N_2427,N_1715);
xor U6666 (N_6666,N_4667,N_4424);
and U6667 (N_6667,N_3490,N_4537);
or U6668 (N_6668,N_4246,N_4120);
nor U6669 (N_6669,N_882,N_1100);
nand U6670 (N_6670,N_4145,N_2976);
or U6671 (N_6671,N_4566,N_1965);
or U6672 (N_6672,N_11,N_714);
or U6673 (N_6673,N_4815,N_2701);
nand U6674 (N_6674,N_196,N_4919);
and U6675 (N_6675,N_1157,N_3455);
nor U6676 (N_6676,N_3518,N_826);
nand U6677 (N_6677,N_4270,N_3005);
nor U6678 (N_6678,N_2871,N_466);
and U6679 (N_6679,N_4771,N_4244);
and U6680 (N_6680,N_4894,N_2671);
nor U6681 (N_6681,N_1908,N_4158);
nor U6682 (N_6682,N_622,N_2771);
nor U6683 (N_6683,N_117,N_684);
or U6684 (N_6684,N_2227,N_4829);
nand U6685 (N_6685,N_3925,N_2552);
and U6686 (N_6686,N_2741,N_4777);
or U6687 (N_6687,N_2212,N_3685);
nor U6688 (N_6688,N_4425,N_2356);
nor U6689 (N_6689,N_1911,N_900);
nor U6690 (N_6690,N_3764,N_4522);
and U6691 (N_6691,N_3258,N_542);
or U6692 (N_6692,N_4019,N_3638);
nand U6693 (N_6693,N_1368,N_916);
and U6694 (N_6694,N_1807,N_4523);
nor U6695 (N_6695,N_520,N_3656);
and U6696 (N_6696,N_2557,N_2167);
nand U6697 (N_6697,N_4941,N_4984);
and U6698 (N_6698,N_1309,N_320);
nor U6699 (N_6699,N_2375,N_994);
nor U6700 (N_6700,N_3678,N_500);
nand U6701 (N_6701,N_4048,N_120);
or U6702 (N_6702,N_2446,N_3648);
nand U6703 (N_6703,N_630,N_430);
nand U6704 (N_6704,N_1932,N_2968);
or U6705 (N_6705,N_4679,N_4869);
or U6706 (N_6706,N_3765,N_3558);
nor U6707 (N_6707,N_1460,N_3240);
or U6708 (N_6708,N_3614,N_1184);
or U6709 (N_6709,N_2273,N_4484);
xnor U6710 (N_6710,N_2514,N_4369);
nor U6711 (N_6711,N_2411,N_1936);
or U6712 (N_6712,N_400,N_2218);
or U6713 (N_6713,N_1515,N_4394);
nand U6714 (N_6714,N_307,N_3146);
or U6715 (N_6715,N_4850,N_1773);
nand U6716 (N_6716,N_820,N_4673);
or U6717 (N_6717,N_4693,N_1478);
or U6718 (N_6718,N_3210,N_2565);
and U6719 (N_6719,N_1372,N_4464);
nor U6720 (N_6720,N_2900,N_4440);
and U6721 (N_6721,N_62,N_2947);
nand U6722 (N_6722,N_1896,N_831);
nand U6723 (N_6723,N_2752,N_4195);
nor U6724 (N_6724,N_3553,N_3321);
nand U6725 (N_6725,N_947,N_2774);
nand U6726 (N_6726,N_3617,N_3820);
and U6727 (N_6727,N_982,N_2981);
nor U6728 (N_6728,N_4426,N_4207);
and U6729 (N_6729,N_3304,N_2386);
and U6730 (N_6730,N_244,N_115);
or U6731 (N_6731,N_2439,N_2035);
and U6732 (N_6732,N_593,N_2905);
xnor U6733 (N_6733,N_1194,N_3140);
xnor U6734 (N_6734,N_2094,N_1436);
or U6735 (N_6735,N_4434,N_2483);
or U6736 (N_6736,N_2878,N_3956);
and U6737 (N_6737,N_2138,N_1449);
nor U6738 (N_6738,N_2843,N_816);
or U6739 (N_6739,N_15,N_4669);
and U6740 (N_6740,N_2250,N_2002);
nor U6741 (N_6741,N_1269,N_1799);
nand U6742 (N_6742,N_822,N_1690);
nor U6743 (N_6743,N_3955,N_57);
nor U6744 (N_6744,N_1422,N_3057);
and U6745 (N_6745,N_4968,N_3902);
or U6746 (N_6746,N_1632,N_929);
nor U6747 (N_6747,N_687,N_4074);
or U6748 (N_6748,N_4339,N_3407);
nor U6749 (N_6749,N_2137,N_4284);
and U6750 (N_6750,N_26,N_1956);
and U6751 (N_6751,N_3114,N_1471);
nand U6752 (N_6752,N_2498,N_4018);
nand U6753 (N_6753,N_3864,N_2772);
xnor U6754 (N_6754,N_3593,N_462);
or U6755 (N_6755,N_2265,N_121);
nor U6756 (N_6756,N_1853,N_3483);
and U6757 (N_6757,N_3951,N_3337);
nand U6758 (N_6758,N_1545,N_4659);
or U6759 (N_6759,N_4569,N_810);
or U6760 (N_6760,N_3498,N_1346);
and U6761 (N_6761,N_4191,N_2865);
or U6762 (N_6762,N_20,N_3911);
and U6763 (N_6763,N_858,N_1020);
nand U6764 (N_6764,N_1566,N_2173);
or U6765 (N_6765,N_1705,N_86);
and U6766 (N_6766,N_2926,N_3);
and U6767 (N_6767,N_1200,N_815);
or U6768 (N_6768,N_4698,N_787);
or U6769 (N_6769,N_2163,N_4125);
and U6770 (N_6770,N_4128,N_265);
and U6771 (N_6771,N_4633,N_2522);
and U6772 (N_6772,N_4945,N_2973);
nand U6773 (N_6773,N_677,N_4514);
or U6774 (N_6774,N_563,N_2436);
nor U6775 (N_6775,N_405,N_2129);
nor U6776 (N_6776,N_837,N_2967);
nor U6777 (N_6777,N_1637,N_3894);
and U6778 (N_6778,N_540,N_3179);
and U6779 (N_6779,N_429,N_3221);
or U6780 (N_6780,N_965,N_1323);
nand U6781 (N_6781,N_3989,N_3738);
nor U6782 (N_6782,N_2892,N_3939);
and U6783 (N_6783,N_2468,N_1999);
nor U6784 (N_6784,N_1096,N_3716);
and U6785 (N_6785,N_2713,N_3071);
nand U6786 (N_6786,N_4901,N_2642);
nor U6787 (N_6787,N_2503,N_3746);
nor U6788 (N_6788,N_124,N_4986);
nor U6789 (N_6789,N_3692,N_262);
nor U6790 (N_6790,N_3147,N_2789);
or U6791 (N_6791,N_1089,N_3239);
and U6792 (N_6792,N_4314,N_1801);
nor U6793 (N_6793,N_2435,N_3852);
nand U6794 (N_6794,N_4549,N_236);
nand U6795 (N_6795,N_948,N_4352);
nor U6796 (N_6796,N_4713,N_3836);
and U6797 (N_6797,N_1533,N_4904);
or U6798 (N_6798,N_3409,N_2817);
nand U6799 (N_6799,N_2150,N_61);
nor U6800 (N_6800,N_3159,N_280);
nand U6801 (N_6801,N_1827,N_3662);
and U6802 (N_6802,N_3266,N_1761);
nor U6803 (N_6803,N_4692,N_4269);
and U6804 (N_6804,N_4324,N_2295);
nor U6805 (N_6805,N_4805,N_1145);
nor U6806 (N_6806,N_3541,N_1748);
xor U6807 (N_6807,N_2047,N_1730);
and U6808 (N_6808,N_4046,N_4831);
nand U6809 (N_6809,N_859,N_868);
nand U6810 (N_6810,N_3921,N_2989);
or U6811 (N_6811,N_588,N_3755);
and U6812 (N_6812,N_347,N_624);
nor U6813 (N_6813,N_2808,N_2023);
nor U6814 (N_6814,N_910,N_433);
nand U6815 (N_6815,N_2712,N_4605);
nor U6816 (N_6816,N_1521,N_2272);
nor U6817 (N_6817,N_843,N_2296);
and U6818 (N_6818,N_2155,N_4882);
xnor U6819 (N_6819,N_4961,N_4681);
nand U6820 (N_6820,N_1354,N_3031);
nand U6821 (N_6821,N_369,N_678);
and U6822 (N_6822,N_2470,N_1777);
or U6823 (N_6823,N_2723,N_1299);
or U6824 (N_6824,N_2793,N_646);
nand U6825 (N_6825,N_2017,N_1129);
nor U6826 (N_6826,N_2591,N_2812);
and U6827 (N_6827,N_1558,N_4820);
nor U6828 (N_6828,N_950,N_898);
nand U6829 (N_6829,N_4482,N_3549);
nand U6830 (N_6830,N_3011,N_3543);
or U6831 (N_6831,N_3034,N_518);
and U6832 (N_6832,N_3017,N_4977);
and U6833 (N_6833,N_424,N_2707);
or U6834 (N_6834,N_647,N_3671);
or U6835 (N_6835,N_3102,N_1419);
nor U6836 (N_6836,N_1212,N_3089);
nand U6837 (N_6837,N_1232,N_364);
or U6838 (N_6838,N_2097,N_2811);
xor U6839 (N_6839,N_2934,N_2338);
nand U6840 (N_6840,N_2428,N_1869);
or U6841 (N_6841,N_377,N_1858);
xnor U6842 (N_6842,N_2414,N_1996);
and U6843 (N_6843,N_3202,N_1876);
nand U6844 (N_6844,N_2280,N_3157);
or U6845 (N_6845,N_3340,N_3858);
or U6846 (N_6846,N_3950,N_3948);
or U6847 (N_6847,N_1889,N_899);
nand U6848 (N_6848,N_4491,N_1442);
or U6849 (N_6849,N_1721,N_3659);
or U6850 (N_6850,N_2297,N_3190);
or U6851 (N_6851,N_3054,N_1429);
and U6852 (N_6852,N_1541,N_3621);
nor U6853 (N_6853,N_2945,N_2751);
nand U6854 (N_6854,N_3002,N_4478);
nand U6855 (N_6855,N_2555,N_3335);
and U6856 (N_6856,N_3775,N_1957);
or U6857 (N_6857,N_482,N_1693);
and U6858 (N_6858,N_4027,N_146);
nand U6859 (N_6859,N_3094,N_1746);
or U6860 (N_6860,N_2962,N_1798);
and U6861 (N_6861,N_2220,N_1591);
or U6862 (N_6862,N_3126,N_4628);
nand U6863 (N_6863,N_72,N_1364);
and U6864 (N_6864,N_2870,N_7);
nand U6865 (N_6865,N_4962,N_2542);
or U6866 (N_6866,N_897,N_179);
and U6867 (N_6867,N_2133,N_116);
nor U6868 (N_6868,N_2,N_3708);
nor U6869 (N_6869,N_1779,N_3018);
nor U6870 (N_6870,N_1736,N_4285);
or U6871 (N_6871,N_2580,N_4967);
or U6872 (N_6872,N_3329,N_3028);
and U6873 (N_6873,N_402,N_4910);
nor U6874 (N_6874,N_611,N_723);
or U6875 (N_6875,N_792,N_3969);
nand U6876 (N_6876,N_1771,N_1301);
nor U6877 (N_6877,N_3640,N_2060);
nand U6878 (N_6878,N_2169,N_1914);
nand U6879 (N_6879,N_175,N_245);
nor U6880 (N_6880,N_3482,N_4554);
nand U6881 (N_6881,N_345,N_1664);
and U6882 (N_6882,N_2073,N_1281);
nand U6883 (N_6883,N_3773,N_3690);
nor U6884 (N_6884,N_2869,N_3613);
or U6885 (N_6885,N_104,N_1370);
nor U6886 (N_6886,N_1366,N_1138);
or U6887 (N_6887,N_2684,N_2520);
nor U6888 (N_6888,N_854,N_4973);
nand U6889 (N_6889,N_1254,N_1099);
and U6890 (N_6890,N_4134,N_2310);
nand U6891 (N_6891,N_4974,N_2289);
nor U6892 (N_6892,N_2601,N_585);
nor U6893 (N_6893,N_1810,N_3510);
nand U6894 (N_6894,N_4718,N_2221);
and U6895 (N_6895,N_4909,N_2497);
or U6896 (N_6896,N_1356,N_2078);
nand U6897 (N_6897,N_4116,N_2721);
xnor U6898 (N_6898,N_58,N_3229);
and U6899 (N_6899,N_3315,N_1862);
xor U6900 (N_6900,N_731,N_2630);
nor U6901 (N_6901,N_4218,N_2826);
and U6902 (N_6902,N_1032,N_2153);
nor U6903 (N_6903,N_667,N_905);
nor U6904 (N_6904,N_539,N_4178);
nor U6905 (N_6905,N_4299,N_4649);
nor U6906 (N_6906,N_602,N_710);
and U6907 (N_6907,N_2343,N_2670);
xor U6908 (N_6908,N_4526,N_3142);
or U6909 (N_6909,N_3869,N_1344);
xnor U6910 (N_6910,N_2052,N_1796);
or U6911 (N_6911,N_285,N_4969);
and U6912 (N_6912,N_968,N_4759);
nand U6913 (N_6913,N_2118,N_4315);
nand U6914 (N_6914,N_864,N_2819);
and U6915 (N_6915,N_4840,N_2491);
nor U6916 (N_6916,N_4507,N_4289);
nor U6917 (N_6917,N_3319,N_4416);
nand U6918 (N_6918,N_221,N_4157);
or U6919 (N_6919,N_4587,N_3025);
nor U6920 (N_6920,N_1961,N_3987);
nand U6921 (N_6921,N_3275,N_3419);
nand U6922 (N_6922,N_1718,N_31);
nor U6923 (N_6923,N_3059,N_1451);
nor U6924 (N_6924,N_3610,N_1448);
nor U6925 (N_6925,N_4788,N_2110);
or U6926 (N_6926,N_557,N_4327);
nand U6927 (N_6927,N_1506,N_3385);
xnor U6928 (N_6928,N_2275,N_2728);
nor U6929 (N_6929,N_314,N_2859);
nand U6930 (N_6930,N_3706,N_2243);
and U6931 (N_6931,N_1652,N_2660);
or U6932 (N_6932,N_2643,N_2704);
xnor U6933 (N_6933,N_619,N_1972);
nand U6934 (N_6934,N_4836,N_1786);
or U6935 (N_6935,N_1687,N_1128);
and U6936 (N_6936,N_1095,N_4455);
nand U6937 (N_6937,N_610,N_3227);
and U6938 (N_6938,N_2681,N_2598);
nand U6939 (N_6939,N_2691,N_3314);
or U6940 (N_6940,N_1461,N_4877);
or U6941 (N_6941,N_3290,N_1118);
and U6942 (N_6942,N_243,N_906);
and U6943 (N_6943,N_2761,N_2455);
and U6944 (N_6944,N_909,N_2818);
nor U6945 (N_6945,N_1624,N_3675);
nand U6946 (N_6946,N_1706,N_617);
nor U6947 (N_6947,N_1806,N_3449);
or U6948 (N_6948,N_2466,N_3137);
nor U6949 (N_6949,N_2784,N_404);
or U6950 (N_6950,N_3284,N_4989);
nor U6951 (N_6951,N_3139,N_2490);
xnor U6952 (N_6952,N_4650,N_4475);
and U6953 (N_6953,N_3222,N_762);
or U6954 (N_6954,N_2512,N_2140);
nand U6955 (N_6955,N_1206,N_697);
nand U6956 (N_6956,N_1127,N_1993);
or U6957 (N_6957,N_2800,N_3633);
and U6958 (N_6958,N_2425,N_4205);
or U6959 (N_6959,N_1639,N_228);
or U6960 (N_6960,N_2095,N_2996);
xor U6961 (N_6961,N_2450,N_3537);
and U6962 (N_6962,N_3604,N_34);
nand U6963 (N_6963,N_4776,N_4632);
nand U6964 (N_6964,N_4264,N_2860);
nand U6965 (N_6965,N_556,N_4551);
nand U6966 (N_6966,N_1284,N_1486);
or U6967 (N_6967,N_1641,N_1334);
nand U6968 (N_6968,N_552,N_4561);
and U6969 (N_6969,N_2953,N_4753);
or U6970 (N_6970,N_2121,N_3919);
or U6971 (N_6971,N_3556,N_2127);
nor U6972 (N_6972,N_2201,N_3805);
nand U6973 (N_6973,N_913,N_252);
xor U6974 (N_6974,N_4173,N_2990);
or U6975 (N_6975,N_3774,N_2895);
nor U6976 (N_6976,N_3045,N_748);
and U6977 (N_6977,N_3757,N_1114);
or U6978 (N_6978,N_1955,N_739);
nand U6979 (N_6979,N_3144,N_757);
nand U6980 (N_6980,N_495,N_388);
and U6981 (N_6981,N_2625,N_3861);
nor U6982 (N_6982,N_634,N_343);
nor U6983 (N_6983,N_703,N_1326);
nor U6984 (N_6984,N_1259,N_3311);
nand U6985 (N_6985,N_919,N_4716);
or U6986 (N_6986,N_3807,N_783);
nor U6987 (N_6987,N_303,N_3489);
nor U6988 (N_6988,N_1187,N_3766);
nor U6989 (N_6989,N_3403,N_4802);
xor U6990 (N_6990,N_681,N_4620);
nor U6991 (N_6991,N_1719,N_2437);
xor U6992 (N_6992,N_1870,N_862);
or U6993 (N_6993,N_1834,N_3795);
and U6994 (N_6994,N_2880,N_1186);
or U6995 (N_6995,N_2419,N_4155);
and U6996 (N_6996,N_4206,N_741);
nand U6997 (N_6997,N_3784,N_3213);
nand U6998 (N_6998,N_1430,N_4034);
and U6999 (N_6999,N_4575,N_2815);
nor U7000 (N_7000,N_632,N_650);
nand U7001 (N_7001,N_3727,N_488);
nand U7002 (N_7002,N_399,N_3586);
or U7003 (N_7003,N_626,N_4497);
nand U7004 (N_7004,N_1231,N_431);
nand U7005 (N_7005,N_1848,N_4931);
and U7006 (N_7006,N_998,N_3926);
xnor U7007 (N_7007,N_1103,N_3252);
and U7008 (N_7008,N_4853,N_2301);
or U7009 (N_7009,N_3463,N_1789);
xor U7010 (N_7010,N_29,N_4202);
nor U7011 (N_7011,N_82,N_3831);
xor U7012 (N_7012,N_4140,N_1410);
nand U7013 (N_7013,N_1484,N_534);
nor U7014 (N_7014,N_4691,N_3010);
nand U7015 (N_7015,N_623,N_769);
nand U7016 (N_7016,N_795,N_1648);
or U7017 (N_7017,N_2248,N_2781);
and U7018 (N_7018,N_195,N_261);
or U7019 (N_7019,N_4133,N_2187);
and U7020 (N_7020,N_3297,N_2858);
nor U7021 (N_7021,N_1034,N_2303);
or U7022 (N_7022,N_944,N_2475);
nor U7023 (N_7023,N_2628,N_1003);
nand U7024 (N_7024,N_4419,N_3332);
nor U7025 (N_7025,N_1725,N_2855);
and U7026 (N_7026,N_1027,N_4124);
and U7027 (N_7027,N_2080,N_3276);
or U7028 (N_7028,N_2186,N_3207);
or U7029 (N_7029,N_3117,N_875);
nand U7030 (N_7030,N_891,N_268);
and U7031 (N_7031,N_4239,N_171);
nand U7032 (N_7032,N_3713,N_325);
and U7033 (N_7033,N_1163,N_192);
nand U7034 (N_7034,N_2283,N_2355);
xnor U7035 (N_7035,N_1893,N_1146);
or U7036 (N_7036,N_4823,N_2126);
and U7037 (N_7037,N_4874,N_1670);
nor U7038 (N_7038,N_4630,N_639);
or U7039 (N_7039,N_3168,N_340);
and U7040 (N_7040,N_1176,N_3214);
or U7041 (N_7041,N_275,N_3743);
nor U7042 (N_7042,N_3433,N_1502);
nand U7043 (N_7043,N_1180,N_2668);
nand U7044 (N_7044,N_2070,N_2241);
nand U7045 (N_7045,N_3573,N_2898);
nand U7046 (N_7046,N_850,N_4253);
or U7047 (N_7047,N_100,N_2048);
or U7048 (N_7048,N_4819,N_4622);
nand U7049 (N_7049,N_4054,N_3972);
nand U7050 (N_7050,N_1831,N_4076);
nand U7051 (N_7051,N_2649,N_4136);
or U7052 (N_7052,N_4690,N_4767);
or U7053 (N_7053,N_2266,N_1978);
and U7054 (N_7054,N_1293,N_3841);
nor U7055 (N_7055,N_4568,N_4543);
nand U7056 (N_7056,N_4647,N_2948);
nand U7057 (N_7057,N_980,N_3243);
nor U7058 (N_7058,N_2307,N_4971);
nor U7059 (N_7059,N_2507,N_3534);
nor U7060 (N_7060,N_4007,N_3626);
nor U7061 (N_7061,N_643,N_443);
or U7062 (N_7062,N_3670,N_2478);
or U7063 (N_7063,N_1785,N_3589);
or U7064 (N_7064,N_1046,N_662);
xnor U7065 (N_7065,N_4541,N_890);
and U7066 (N_7066,N_516,N_4737);
nand U7067 (N_7067,N_313,N_2226);
and U7068 (N_7068,N_338,N_257);
and U7069 (N_7069,N_1924,N_1538);
and U7070 (N_7070,N_1627,N_92);
nand U7071 (N_7071,N_1039,N_64);
and U7072 (N_7072,N_4717,N_3567);
or U7073 (N_7073,N_296,N_4665);
nor U7074 (N_7074,N_1115,N_1030);
nor U7075 (N_7075,N_1376,N_797);
and U7076 (N_7076,N_99,N_312);
nand U7077 (N_7077,N_2488,N_1617);
nor U7078 (N_7078,N_4545,N_1962);
nand U7079 (N_7079,N_1065,N_1202);
and U7080 (N_7080,N_1240,N_4306);
xnor U7081 (N_7081,N_333,N_4081);
nor U7082 (N_7082,N_4401,N_68);
nand U7083 (N_7083,N_4129,N_711);
nand U7084 (N_7084,N_3630,N_2970);
and U7085 (N_7085,N_2311,N_3289);
nor U7086 (N_7086,N_218,N_3077);
and U7087 (N_7087,N_2931,N_642);
nand U7088 (N_7088,N_4652,N_881);
nor U7089 (N_7089,N_4502,N_3093);
nand U7090 (N_7090,N_3597,N_1772);
nand U7091 (N_7091,N_356,N_2349);
or U7092 (N_7092,N_1517,N_477);
nor U7093 (N_7093,N_4572,N_412);
or U7094 (N_7094,N_4141,N_380);
xnor U7095 (N_7095,N_885,N_2674);
nor U7096 (N_7096,N_3879,N_4229);
xor U7097 (N_7097,N_3107,N_1886);
xor U7098 (N_7098,N_779,N_3622);
nand U7099 (N_7099,N_1056,N_1480);
nand U7100 (N_7100,N_2504,N_4123);
nor U7101 (N_7101,N_1205,N_1054);
and U7102 (N_7102,N_3491,N_2714);
nand U7103 (N_7103,N_3052,N_3149);
nor U7104 (N_7104,N_1363,N_2883);
or U7105 (N_7105,N_271,N_1564);
or U7106 (N_7106,N_4664,N_3611);
and U7107 (N_7107,N_857,N_1058);
nand U7108 (N_7108,N_235,N_581);
nor U7109 (N_7109,N_2372,N_3465);
nand U7110 (N_7110,N_4219,N_2255);
or U7111 (N_7111,N_3608,N_4582);
and U7112 (N_7112,N_4177,N_883);
or U7113 (N_7113,N_2998,N_4213);
or U7114 (N_7114,N_4533,N_2975);
and U7115 (N_7115,N_2451,N_1387);
nand U7116 (N_7116,N_2143,N_4703);
and U7117 (N_7117,N_970,N_4112);
nor U7118 (N_7118,N_4629,N_4060);
and U7119 (N_7119,N_2180,N_342);
nor U7120 (N_7120,N_4803,N_365);
and U7121 (N_7121,N_2946,N_2570);
or U7122 (N_7122,N_131,N_474);
nand U7123 (N_7123,N_1318,N_962);
and U7124 (N_7124,N_1130,N_1347);
nand U7125 (N_7125,N_671,N_4843);
nor U7126 (N_7126,N_425,N_1440);
nand U7127 (N_7127,N_1844,N_334);
and U7128 (N_7128,N_1623,N_1160);
or U7129 (N_7129,N_2330,N_1847);
nor U7130 (N_7130,N_958,N_541);
or U7131 (N_7131,N_1954,N_2622);
and U7132 (N_7132,N_97,N_519);
xnor U7133 (N_7133,N_4508,N_326);
nand U7134 (N_7134,N_2603,N_1245);
or U7135 (N_7135,N_571,N_1421);
or U7136 (N_7136,N_2833,N_3804);
nand U7137 (N_7137,N_393,N_4458);
xnor U7138 (N_7138,N_2362,N_3472);
nor U7139 (N_7139,N_4914,N_2389);
nand U7140 (N_7140,N_3373,N_3635);
and U7141 (N_7141,N_2245,N_1842);
and U7142 (N_7142,N_4954,N_4292);
or U7143 (N_7143,N_3196,N_3881);
xor U7144 (N_7144,N_1744,N_1661);
nand U7145 (N_7145,N_182,N_1608);
nor U7146 (N_7146,N_3695,N_4276);
or U7147 (N_7147,N_1432,N_1716);
nor U7148 (N_7148,N_800,N_807);
nor U7149 (N_7149,N_4950,N_4916);
nor U7150 (N_7150,N_284,N_2574);
nor U7151 (N_7151,N_3958,N_2792);
and U7152 (N_7152,N_1863,N_3581);
and U7153 (N_7153,N_1437,N_1544);
and U7154 (N_7154,N_3744,N_4920);
or U7155 (N_7155,N_3666,N_1794);
or U7156 (N_7156,N_2718,N_4726);
or U7157 (N_7157,N_4402,N_3397);
nand U7158 (N_7158,N_3125,N_1463);
xor U7159 (N_7159,N_4186,N_2487);
nor U7160 (N_7160,N_789,N_1812);
or U7161 (N_7161,N_521,N_2972);
or U7162 (N_7162,N_3088,N_3707);
nor U7163 (N_7163,N_3803,N_2697);
or U7164 (N_7164,N_1922,N_2548);
and U7165 (N_7165,N_1428,N_606);
nor U7166 (N_7166,N_2320,N_210);
nand U7167 (N_7167,N_4381,N_1296);
or U7168 (N_7168,N_3874,N_4268);
or U7169 (N_7169,N_848,N_2850);
or U7170 (N_7170,N_1291,N_559);
and U7171 (N_7171,N_2903,N_4255);
and U7172 (N_7172,N_2294,N_1977);
and U7173 (N_7173,N_2619,N_3001);
or U7174 (N_7174,N_2877,N_260);
nor U7175 (N_7175,N_3937,N_4248);
nor U7176 (N_7176,N_4095,N_2392);
and U7177 (N_7177,N_1219,N_922);
xnor U7178 (N_7178,N_3900,N_1635);
xor U7179 (N_7179,N_1686,N_1218);
xnor U7180 (N_7180,N_157,N_1097);
nand U7181 (N_7181,N_107,N_1737);
xnor U7182 (N_7182,N_3004,N_3547);
nand U7183 (N_7183,N_428,N_2827);
xnor U7184 (N_7184,N_3318,N_4316);
or U7185 (N_7185,N_2562,N_832);
and U7186 (N_7186,N_3076,N_3405);
nor U7187 (N_7187,N_4132,N_2782);
nor U7188 (N_7188,N_1266,N_3394);
nor U7189 (N_7189,N_4467,N_1412);
nand U7190 (N_7190,N_208,N_3003);
or U7191 (N_7191,N_4014,N_3440);
xnor U7192 (N_7192,N_310,N_2676);
xor U7193 (N_7193,N_1183,N_3910);
nand U7194 (N_7194,N_410,N_4092);
or U7195 (N_7195,N_690,N_2131);
or U7196 (N_7196,N_4103,N_3216);
nor U7197 (N_7197,N_4943,N_1833);
nand U7198 (N_7198,N_895,N_4562);
nand U7199 (N_7199,N_4565,N_2474);
nor U7200 (N_7200,N_247,N_720);
nor U7201 (N_7201,N_675,N_658);
or U7202 (N_7202,N_4684,N_504);
or U7203 (N_7203,N_1175,N_4442);
or U7204 (N_7204,N_4263,N_2802);
nor U7205 (N_7205,N_2088,N_4745);
xnor U7206 (N_7206,N_3313,N_1192);
xor U7207 (N_7207,N_3799,N_849);
and U7208 (N_7208,N_3236,N_4760);
xnor U7209 (N_7209,N_1134,N_106);
nor U7210 (N_7210,N_4122,N_1073);
xor U7211 (N_7211,N_2889,N_2705);
nor U7212 (N_7212,N_4856,N_2753);
nand U7213 (N_7213,N_3165,N_1374);
nand U7214 (N_7214,N_532,N_3264);
or U7215 (N_7215,N_348,N_3133);
and U7216 (N_7216,N_4834,N_1001);
nand U7217 (N_7217,N_35,N_2033);
nand U7218 (N_7218,N_4333,N_1008);
and U7219 (N_7219,N_3810,N_2122);
nor U7220 (N_7220,N_214,N_1501);
nor U7221 (N_7221,N_656,N_573);
and U7222 (N_7222,N_3355,N_1750);
nand U7223 (N_7223,N_4756,N_2748);
or U7224 (N_7224,N_665,N_1431);
nand U7225 (N_7225,N_3529,N_4520);
or U7226 (N_7226,N_392,N_446);
or U7227 (N_7227,N_716,N_4361);
nor U7228 (N_7228,N_1036,N_4226);
and U7229 (N_7229,N_1747,N_1811);
nor U7230 (N_7230,N_3643,N_187);
and U7231 (N_7231,N_1885,N_350);
or U7232 (N_7232,N_1398,N_3783);
nand U7233 (N_7233,N_358,N_149);
or U7234 (N_7234,N_3055,N_4720);
xor U7235 (N_7235,N_3474,N_3560);
and U7236 (N_7236,N_3571,N_3523);
and U7237 (N_7237,N_4956,N_444);
nand U7238 (N_7238,N_1379,N_527);
and U7239 (N_7239,N_3985,N_1409);
xnor U7240 (N_7240,N_2480,N_3658);
nand U7241 (N_7241,N_4053,N_4117);
xnor U7242 (N_7242,N_967,N_324);
or U7243 (N_7243,N_4104,N_3037);
nor U7244 (N_7244,N_759,N_1606);
nand U7245 (N_7245,N_2074,N_3944);
nand U7246 (N_7246,N_3353,N_4456);
nor U7247 (N_7247,N_1019,N_3700);
xor U7248 (N_7248,N_4240,N_525);
or U7249 (N_7249,N_2445,N_2937);
nand U7250 (N_7250,N_1945,N_2442);
nor U7251 (N_7251,N_3940,N_2464);
and U7252 (N_7252,N_4595,N_2951);
nor U7253 (N_7253,N_4029,N_2724);
nor U7254 (N_7254,N_3066,N_4056);
and U7255 (N_7255,N_3389,N_1946);
xor U7256 (N_7256,N_2115,N_2854);
and U7257 (N_7257,N_4513,N_2540);
and U7258 (N_7258,N_3352,N_1238);
nor U7259 (N_7259,N_172,N_2525);
or U7260 (N_7260,N_3478,N_2160);
nor U7261 (N_7261,N_2271,N_4215);
nand U7262 (N_7262,N_226,N_1582);
or U7263 (N_7263,N_2991,N_4998);
or U7264 (N_7264,N_3559,N_515);
or U7265 (N_7265,N_1006,N_4169);
and U7266 (N_7266,N_3576,N_150);
nand U7267 (N_7267,N_177,N_4860);
nor U7268 (N_7268,N_3411,N_3053);
or U7269 (N_7269,N_2405,N_125);
or U7270 (N_7270,N_2251,N_4573);
and U7271 (N_7271,N_3183,N_1064);
and U7272 (N_7272,N_3741,N_4409);
nand U7273 (N_7273,N_852,N_1663);
nor U7274 (N_7274,N_30,N_1731);
nor U7275 (N_7275,N_3460,N_2637);
or U7276 (N_7276,N_1974,N_3047);
and U7277 (N_7277,N_3180,N_2571);
nor U7278 (N_7278,N_1604,N_1813);
nor U7279 (N_7279,N_4204,N_2408);
nand U7280 (N_7280,N_4072,N_1787);
and U7281 (N_7281,N_2453,N_707);
or U7282 (N_7282,N_2822,N_2760);
xor U7283 (N_7283,N_2708,N_773);
or U7284 (N_7284,N_3550,N_1051);
and U7285 (N_7285,N_1414,N_378);
or U7286 (N_7286,N_3346,N_3619);
nor U7287 (N_7287,N_673,N_351);
and U7288 (N_7288,N_4949,N_3848);
nand U7289 (N_7289,N_2204,N_1597);
xor U7290 (N_7290,N_1082,N_745);
nor U7291 (N_7291,N_1382,N_2465);
nand U7292 (N_7292,N_0,N_448);
xor U7293 (N_7293,N_4031,N_2448);
nor U7294 (N_7294,N_4564,N_1928);
xor U7295 (N_7295,N_4059,N_590);
and U7296 (N_7296,N_2814,N_1826);
or U7297 (N_7297,N_3525,N_2085);
and U7298 (N_7298,N_1009,N_3787);
or U7299 (N_7299,N_2786,N_3404);
and U7300 (N_7300,N_3299,N_1525);
and U7301 (N_7301,N_4111,N_1697);
nand U7302 (N_7302,N_4065,N_1888);
xnor U7303 (N_7303,N_1242,N_845);
xor U7304 (N_7304,N_1083,N_1898);
or U7305 (N_7305,N_2044,N_3105);
and U7306 (N_7306,N_2821,N_4100);
nand U7307 (N_7307,N_1938,N_3192);
or U7308 (N_7308,N_3458,N_3642);
nor U7309 (N_7309,N_4689,N_4857);
nor U7310 (N_7310,N_972,N_18);
nor U7311 (N_7311,N_4724,N_1783);
nor U7312 (N_7312,N_2062,N_1076);
and U7313 (N_7313,N_4816,N_1179);
and U7314 (N_7314,N_1881,N_4892);
nand U7315 (N_7315,N_2202,N_2788);
nor U7316 (N_7316,N_1857,N_4388);
xor U7317 (N_7317,N_4617,N_3261);
xnor U7318 (N_7318,N_2053,N_863);
nand U7319 (N_7319,N_4983,N_2545);
nand U7320 (N_7320,N_4792,N_3702);
or U7321 (N_7321,N_2130,N_1531);
or U7322 (N_7322,N_4621,N_291);
nand U7323 (N_7323,N_4774,N_200);
or U7324 (N_7324,N_923,N_2383);
or U7325 (N_7325,N_4833,N_2100);
nor U7326 (N_7326,N_784,N_2982);
nand U7327 (N_7327,N_2347,N_4794);
nor U7328 (N_7328,N_768,N_1085);
nand U7329 (N_7329,N_3390,N_1562);
or U7330 (N_7330,N_2653,N_1152);
nor U7331 (N_7331,N_2861,N_3051);
or U7332 (N_7332,N_2665,N_705);
nand U7333 (N_7333,N_4799,N_1607);
nor U7334 (N_7334,N_1651,N_870);
xnor U7335 (N_7335,N_618,N_1510);
or U7336 (N_7336,N_2135,N_3050);
and U7337 (N_7337,N_2686,N_2374);
or U7338 (N_7338,N_3143,N_3316);
and U7339 (N_7339,N_957,N_3309);
and U7340 (N_7340,N_691,N_84);
or U7341 (N_7341,N_4927,N_2029);
or U7342 (N_7342,N_1337,N_294);
nor U7343 (N_7343,N_4049,N_2260);
nand U7344 (N_7344,N_270,N_1038);
and U7345 (N_7345,N_742,N_3548);
or U7346 (N_7346,N_2144,N_1452);
nor U7347 (N_7347,N_4265,N_2041);
nand U7348 (N_7348,N_1539,N_2640);
or U7349 (N_7349,N_3043,N_3251);
xnor U7350 (N_7350,N_2887,N_4197);
and U7351 (N_7351,N_2763,N_193);
or U7352 (N_7352,N_3424,N_4608);
and U7353 (N_7353,N_3973,N_4824);
and U7354 (N_7354,N_4958,N_4993);
nand U7355 (N_7355,N_3605,N_2496);
and U7356 (N_7356,N_2341,N_597);
and U7357 (N_7357,N_3382,N_2687);
nand U7358 (N_7358,N_4748,N_4959);
or U7359 (N_7359,N_2620,N_2749);
and U7360 (N_7360,N_415,N_3693);
nand U7361 (N_7361,N_3522,N_2738);
nor U7362 (N_7362,N_2613,N_3816);
nor U7363 (N_7363,N_337,N_1441);
nor U7364 (N_7364,N_2010,N_2205);
or U7365 (N_7365,N_3008,N_1317);
nor U7366 (N_7366,N_3122,N_2055);
nand U7367 (N_7367,N_2421,N_2986);
or U7368 (N_7368,N_2851,N_2322);
and U7369 (N_7369,N_3402,N_4933);
nor U7370 (N_7370,N_2165,N_4114);
or U7371 (N_7371,N_362,N_4243);
and U7372 (N_7372,N_2132,N_1043);
nor U7373 (N_7373,N_2730,N_4662);
nor U7374 (N_7374,N_436,N_2339);
or U7375 (N_7375,N_4185,N_2262);
or U7376 (N_7376,N_4821,N_2452);
nor U7377 (N_7377,N_3830,N_725);
and U7378 (N_7378,N_804,N_1722);
and U7379 (N_7379,N_4602,N_2084);
nor U7380 (N_7380,N_3348,N_201);
nor U7381 (N_7381,N_4964,N_4307);
nor U7382 (N_7382,N_663,N_1004);
nand U7383 (N_7383,N_3242,N_166);
or U7384 (N_7384,N_4308,N_4071);
nor U7385 (N_7385,N_3725,N_2690);
nand U7386 (N_7386,N_1583,N_1603);
and U7387 (N_7387,N_1014,N_1482);
nand U7388 (N_7388,N_3968,N_1119);
nor U7389 (N_7389,N_1699,N_4077);
nand U7390 (N_7390,N_4298,N_4848);
xor U7391 (N_7391,N_1821,N_4355);
nand U7392 (N_7392,N_10,N_4257);
nor U7393 (N_7393,N_4733,N_785);
nor U7394 (N_7394,N_4227,N_3734);
and U7395 (N_7395,N_3193,N_4088);
nand U7396 (N_7396,N_1235,N_2729);
nand U7397 (N_7397,N_1644,N_1067);
nand U7398 (N_7398,N_4534,N_1676);
nor U7399 (N_7399,N_2983,N_952);
nor U7400 (N_7400,N_1297,N_4871);
nor U7401 (N_7401,N_793,N_3797);
nand U7402 (N_7402,N_3462,N_2454);
or U7403 (N_7403,N_4004,N_3015);
or U7404 (N_7404,N_4485,N_1808);
and U7405 (N_7405,N_4898,N_1342);
or U7406 (N_7406,N_1360,N_4131);
and U7407 (N_7407,N_3475,N_1298);
nor U7408 (N_7408,N_1357,N_3485);
or U7409 (N_7409,N_4380,N_799);
nand U7410 (N_7410,N_3976,N_1504);
nand U7411 (N_7411,N_3070,N_4295);
and U7412 (N_7412,N_1760,N_3361);
xnor U7413 (N_7413,N_1424,N_3112);
and U7414 (N_7414,N_2195,N_139);
and U7415 (N_7415,N_3322,N_3351);
and U7416 (N_7416,N_2531,N_3897);
or U7417 (N_7417,N_1343,N_2209);
and U7418 (N_7418,N_4637,N_614);
and U7419 (N_7419,N_2467,N_1645);
or U7420 (N_7420,N_2063,N_19);
nor U7421 (N_7421,N_2337,N_4222);
nor U7422 (N_7422,N_4450,N_2561);
xnor U7423 (N_7423,N_3014,N_3211);
and U7424 (N_7424,N_1524,N_818);
and U7425 (N_7425,N_4739,N_809);
nand U7426 (N_7426,N_3641,N_4925);
or U7427 (N_7427,N_4357,N_372);
nor U7428 (N_7428,N_3302,N_4868);
and U7429 (N_7429,N_2476,N_276);
xor U7430 (N_7430,N_4196,N_2606);
nor U7431 (N_7431,N_4391,N_3062);
nor U7432 (N_7432,N_69,N_4390);
nor U7433 (N_7433,N_2633,N_1197);
nor U7434 (N_7434,N_2225,N_4676);
nor U7435 (N_7435,N_2919,N_761);
nor U7436 (N_7436,N_3245,N_3098);
xnor U7437 (N_7437,N_169,N_3467);
nand U7438 (N_7438,N_293,N_2182);
and U7439 (N_7439,N_1341,N_1901);
xnor U7440 (N_7440,N_2096,N_544);
nand U7441 (N_7441,N_2614,N_2102);
or U7442 (N_7442,N_2500,N_4567);
or U7443 (N_7443,N_3769,N_4891);
or U7444 (N_7444,N_1294,N_3049);
nand U7445 (N_7445,N_4730,N_2979);
or U7446 (N_7446,N_4082,N_2258);
or U7447 (N_7447,N_3875,N_1867);
nor U7448 (N_7448,N_1314,N_1055);
nand U7449 (N_7449,N_2908,N_3350);
nand U7450 (N_7450,N_2166,N_2663);
xnor U7451 (N_7451,N_1353,N_2662);
or U7452 (N_7452,N_4929,N_3256);
or U7453 (N_7453,N_530,N_1228);
nand U7454 (N_7454,N_802,N_4505);
or U7455 (N_7455,N_4770,N_4854);
nor U7456 (N_7456,N_4492,N_4047);
or U7457 (N_7457,N_227,N_3305);
nor U7458 (N_7458,N_4093,N_2259);
xor U7459 (N_7459,N_2319,N_3821);
or U7460 (N_7460,N_1895,N_3120);
nor U7461 (N_7461,N_4398,N_2348);
or U7462 (N_7462,N_302,N_674);
nand U7463 (N_7463,N_1832,N_220);
nor U7464 (N_7464,N_3997,N_3291);
nand U7465 (N_7465,N_846,N_1860);
or U7466 (N_7466,N_4835,N_3320);
or U7467 (N_7467,N_1864,N_165);
and U7468 (N_7468,N_2276,N_2113);
xor U7469 (N_7469,N_3777,N_548);
and U7470 (N_7470,N_3790,N_782);
nand U7471 (N_7471,N_4535,N_3466);
or U7472 (N_7472,N_3961,N_1174);
nand U7473 (N_7473,N_3888,N_1018);
and U7474 (N_7474,N_1276,N_4616);
and U7475 (N_7475,N_4322,N_1498);
or U7476 (N_7476,N_3431,N_1741);
nor U7477 (N_7477,N_3492,N_2304);
and U7478 (N_7478,N_2024,N_1802);
nand U7479 (N_7479,N_2673,N_1327);
nor U7480 (N_7480,N_4403,N_4639);
and U7481 (N_7481,N_2477,N_2207);
or U7482 (N_7482,N_2416,N_299);
nand U7483 (N_7483,N_3484,N_336);
or U7484 (N_7484,N_4210,N_2071);
nor U7485 (N_7485,N_3515,N_774);
and U7486 (N_7486,N_3228,N_2308);
and U7487 (N_7487,N_1126,N_4812);
nand U7488 (N_7488,N_2264,N_332);
or U7489 (N_7489,N_3896,N_3974);
and U7490 (N_7490,N_2004,N_1088);
nand U7491 (N_7491,N_480,N_2806);
and U7492 (N_7492,N_4644,N_403);
nand U7493 (N_7493,N_4337,N_2692);
xor U7494 (N_7494,N_3421,N_3048);
and U7495 (N_7495,N_3339,N_1581);
or U7496 (N_7496,N_2747,N_2364);
nor U7497 (N_7497,N_4334,N_4906);
nor U7498 (N_7498,N_3457,N_3170);
nor U7499 (N_7499,N_3124,N_3579);
nor U7500 (N_7500,N_952,N_1406);
xnor U7501 (N_7501,N_218,N_2714);
or U7502 (N_7502,N_4425,N_1900);
nor U7503 (N_7503,N_2756,N_3419);
nor U7504 (N_7504,N_4290,N_3734);
nand U7505 (N_7505,N_4302,N_3160);
nand U7506 (N_7506,N_1274,N_280);
nand U7507 (N_7507,N_1807,N_923);
nand U7508 (N_7508,N_2571,N_4602);
nor U7509 (N_7509,N_2554,N_408);
and U7510 (N_7510,N_683,N_1244);
nor U7511 (N_7511,N_4622,N_46);
and U7512 (N_7512,N_690,N_182);
nor U7513 (N_7513,N_3320,N_3586);
or U7514 (N_7514,N_1218,N_416);
xnor U7515 (N_7515,N_229,N_3829);
nand U7516 (N_7516,N_346,N_3184);
nor U7517 (N_7517,N_4727,N_202);
or U7518 (N_7518,N_1112,N_4326);
and U7519 (N_7519,N_3640,N_1111);
nor U7520 (N_7520,N_996,N_2128);
nand U7521 (N_7521,N_446,N_2007);
and U7522 (N_7522,N_3213,N_4539);
xor U7523 (N_7523,N_1571,N_319);
xnor U7524 (N_7524,N_309,N_4544);
or U7525 (N_7525,N_216,N_1098);
nor U7526 (N_7526,N_4334,N_2345);
nor U7527 (N_7527,N_1296,N_2368);
nor U7528 (N_7528,N_3134,N_4071);
nor U7529 (N_7529,N_2454,N_2897);
xor U7530 (N_7530,N_1649,N_4975);
or U7531 (N_7531,N_1684,N_4259);
nand U7532 (N_7532,N_2046,N_2326);
and U7533 (N_7533,N_3134,N_4081);
nand U7534 (N_7534,N_4686,N_1335);
nand U7535 (N_7535,N_3061,N_698);
or U7536 (N_7536,N_3570,N_1551);
nor U7537 (N_7537,N_3470,N_3285);
or U7538 (N_7538,N_4521,N_1588);
xnor U7539 (N_7539,N_1200,N_1552);
and U7540 (N_7540,N_2485,N_1208);
nand U7541 (N_7541,N_2699,N_1292);
nand U7542 (N_7542,N_1101,N_3808);
nor U7543 (N_7543,N_2705,N_4512);
nor U7544 (N_7544,N_1171,N_299);
and U7545 (N_7545,N_2672,N_2568);
or U7546 (N_7546,N_4961,N_4867);
xor U7547 (N_7547,N_4569,N_4872);
nand U7548 (N_7548,N_87,N_1440);
xor U7549 (N_7549,N_3184,N_4136);
and U7550 (N_7550,N_3842,N_3358);
and U7551 (N_7551,N_4114,N_261);
or U7552 (N_7552,N_4951,N_3043);
nor U7553 (N_7553,N_1119,N_3553);
xnor U7554 (N_7554,N_3065,N_2295);
or U7555 (N_7555,N_2059,N_916);
and U7556 (N_7556,N_3566,N_4862);
and U7557 (N_7557,N_4221,N_1554);
nand U7558 (N_7558,N_4459,N_4491);
or U7559 (N_7559,N_383,N_3501);
nand U7560 (N_7560,N_2011,N_1585);
nand U7561 (N_7561,N_2730,N_874);
nor U7562 (N_7562,N_1761,N_3181);
nand U7563 (N_7563,N_529,N_583);
or U7564 (N_7564,N_300,N_1177);
nor U7565 (N_7565,N_1769,N_191);
and U7566 (N_7566,N_903,N_4257);
xnor U7567 (N_7567,N_2308,N_2563);
nor U7568 (N_7568,N_4250,N_4667);
and U7569 (N_7569,N_70,N_2153);
nor U7570 (N_7570,N_760,N_1608);
and U7571 (N_7571,N_3559,N_2356);
and U7572 (N_7572,N_529,N_4283);
nand U7573 (N_7573,N_592,N_4176);
nand U7574 (N_7574,N_3100,N_3794);
nand U7575 (N_7575,N_2373,N_1652);
and U7576 (N_7576,N_2335,N_2868);
nor U7577 (N_7577,N_4151,N_3571);
nand U7578 (N_7578,N_477,N_4284);
nor U7579 (N_7579,N_1653,N_1437);
nor U7580 (N_7580,N_44,N_257);
nor U7581 (N_7581,N_1328,N_4970);
or U7582 (N_7582,N_1267,N_3129);
or U7583 (N_7583,N_1690,N_2211);
nand U7584 (N_7584,N_1769,N_1860);
and U7585 (N_7585,N_1595,N_324);
nand U7586 (N_7586,N_4097,N_2432);
or U7587 (N_7587,N_1371,N_1552);
or U7588 (N_7588,N_4701,N_2852);
nor U7589 (N_7589,N_3048,N_4586);
and U7590 (N_7590,N_1458,N_3811);
or U7591 (N_7591,N_2070,N_2840);
nand U7592 (N_7592,N_1867,N_2116);
nand U7593 (N_7593,N_586,N_3828);
and U7594 (N_7594,N_1706,N_1528);
nand U7595 (N_7595,N_948,N_4770);
and U7596 (N_7596,N_4238,N_4991);
nand U7597 (N_7597,N_4234,N_4727);
nand U7598 (N_7598,N_1063,N_459);
nor U7599 (N_7599,N_2522,N_1291);
nor U7600 (N_7600,N_927,N_3231);
and U7601 (N_7601,N_3256,N_3057);
and U7602 (N_7602,N_3029,N_4266);
nand U7603 (N_7603,N_1992,N_4687);
or U7604 (N_7604,N_1152,N_749);
and U7605 (N_7605,N_317,N_3482);
or U7606 (N_7606,N_2496,N_2253);
or U7607 (N_7607,N_3181,N_1431);
or U7608 (N_7608,N_1987,N_1738);
and U7609 (N_7609,N_1025,N_806);
xnor U7610 (N_7610,N_229,N_2273);
nor U7611 (N_7611,N_1336,N_4020);
nand U7612 (N_7612,N_535,N_3191);
and U7613 (N_7613,N_3882,N_489);
and U7614 (N_7614,N_3085,N_3224);
and U7615 (N_7615,N_4168,N_2586);
or U7616 (N_7616,N_894,N_1604);
nor U7617 (N_7617,N_89,N_2309);
xor U7618 (N_7618,N_4340,N_607);
or U7619 (N_7619,N_4510,N_4368);
and U7620 (N_7620,N_3768,N_4418);
xnor U7621 (N_7621,N_2205,N_2944);
or U7622 (N_7622,N_3605,N_474);
and U7623 (N_7623,N_379,N_3157);
nand U7624 (N_7624,N_4986,N_4264);
nand U7625 (N_7625,N_1655,N_1635);
or U7626 (N_7626,N_1856,N_4362);
and U7627 (N_7627,N_283,N_2873);
and U7628 (N_7628,N_1795,N_4263);
nand U7629 (N_7629,N_733,N_2705);
or U7630 (N_7630,N_2918,N_1000);
nand U7631 (N_7631,N_4608,N_3161);
nand U7632 (N_7632,N_4962,N_2221);
or U7633 (N_7633,N_4874,N_4530);
or U7634 (N_7634,N_4758,N_1597);
nand U7635 (N_7635,N_1491,N_2113);
or U7636 (N_7636,N_764,N_2582);
nor U7637 (N_7637,N_2200,N_4130);
nand U7638 (N_7638,N_3007,N_4238);
nand U7639 (N_7639,N_4657,N_3447);
and U7640 (N_7640,N_2651,N_951);
or U7641 (N_7641,N_3942,N_157);
xor U7642 (N_7642,N_274,N_289);
and U7643 (N_7643,N_3682,N_999);
xor U7644 (N_7644,N_2483,N_901);
nor U7645 (N_7645,N_4036,N_621);
nand U7646 (N_7646,N_700,N_1635);
nand U7647 (N_7647,N_2,N_2986);
nand U7648 (N_7648,N_771,N_2364);
or U7649 (N_7649,N_4831,N_2256);
and U7650 (N_7650,N_793,N_4275);
nand U7651 (N_7651,N_4598,N_2446);
nand U7652 (N_7652,N_1163,N_486);
or U7653 (N_7653,N_4721,N_575);
and U7654 (N_7654,N_1305,N_934);
nand U7655 (N_7655,N_3006,N_1807);
or U7656 (N_7656,N_3591,N_687);
nor U7657 (N_7657,N_2874,N_180);
nand U7658 (N_7658,N_4636,N_4846);
or U7659 (N_7659,N_2553,N_4373);
nand U7660 (N_7660,N_3483,N_67);
and U7661 (N_7661,N_1357,N_2824);
nor U7662 (N_7662,N_2111,N_4199);
nor U7663 (N_7663,N_1551,N_71);
nor U7664 (N_7664,N_3224,N_3878);
and U7665 (N_7665,N_2178,N_3268);
xnor U7666 (N_7666,N_3930,N_2080);
nor U7667 (N_7667,N_2489,N_2513);
nand U7668 (N_7668,N_1997,N_3678);
nand U7669 (N_7669,N_1186,N_2820);
nor U7670 (N_7670,N_812,N_4006);
and U7671 (N_7671,N_4935,N_408);
nor U7672 (N_7672,N_174,N_4080);
nor U7673 (N_7673,N_941,N_2918);
nor U7674 (N_7674,N_1417,N_4494);
and U7675 (N_7675,N_2776,N_342);
nand U7676 (N_7676,N_842,N_1571);
nor U7677 (N_7677,N_3931,N_2625);
or U7678 (N_7678,N_575,N_4941);
nor U7679 (N_7679,N_1811,N_780);
nand U7680 (N_7680,N_2496,N_4596);
nand U7681 (N_7681,N_3844,N_1973);
and U7682 (N_7682,N_4648,N_3905);
nand U7683 (N_7683,N_2811,N_221);
nor U7684 (N_7684,N_2726,N_4102);
and U7685 (N_7685,N_2317,N_3795);
and U7686 (N_7686,N_544,N_3283);
xnor U7687 (N_7687,N_848,N_4995);
or U7688 (N_7688,N_4053,N_1368);
and U7689 (N_7689,N_2914,N_4175);
nand U7690 (N_7690,N_4317,N_3777);
and U7691 (N_7691,N_2262,N_939);
nand U7692 (N_7692,N_2368,N_915);
and U7693 (N_7693,N_3439,N_2372);
nor U7694 (N_7694,N_420,N_2575);
nand U7695 (N_7695,N_791,N_2131);
nor U7696 (N_7696,N_3813,N_2085);
and U7697 (N_7697,N_469,N_713);
and U7698 (N_7698,N_1034,N_1217);
xor U7699 (N_7699,N_3006,N_2027);
nand U7700 (N_7700,N_3005,N_1176);
and U7701 (N_7701,N_3094,N_2914);
nor U7702 (N_7702,N_2778,N_978);
or U7703 (N_7703,N_3573,N_3489);
xnor U7704 (N_7704,N_3582,N_673);
xor U7705 (N_7705,N_1522,N_2729);
nand U7706 (N_7706,N_2202,N_3798);
nor U7707 (N_7707,N_3726,N_722);
or U7708 (N_7708,N_526,N_3112);
nor U7709 (N_7709,N_1677,N_1900);
and U7710 (N_7710,N_3166,N_267);
or U7711 (N_7711,N_3772,N_3003);
nor U7712 (N_7712,N_2051,N_4918);
nor U7713 (N_7713,N_1556,N_3815);
or U7714 (N_7714,N_83,N_2896);
nand U7715 (N_7715,N_4512,N_4866);
and U7716 (N_7716,N_82,N_3102);
and U7717 (N_7717,N_2979,N_3780);
nand U7718 (N_7718,N_252,N_2682);
or U7719 (N_7719,N_234,N_93);
nor U7720 (N_7720,N_2577,N_1527);
xnor U7721 (N_7721,N_4872,N_4733);
nand U7722 (N_7722,N_1778,N_3164);
nor U7723 (N_7723,N_1514,N_654);
and U7724 (N_7724,N_1088,N_3380);
nor U7725 (N_7725,N_2925,N_4344);
xnor U7726 (N_7726,N_1898,N_2141);
nor U7727 (N_7727,N_4522,N_2107);
and U7728 (N_7728,N_2498,N_1659);
or U7729 (N_7729,N_725,N_1139);
or U7730 (N_7730,N_3421,N_4426);
nor U7731 (N_7731,N_4659,N_925);
and U7732 (N_7732,N_3322,N_4612);
xnor U7733 (N_7733,N_3757,N_4848);
nand U7734 (N_7734,N_2875,N_1637);
nand U7735 (N_7735,N_2741,N_1025);
or U7736 (N_7736,N_339,N_4490);
or U7737 (N_7737,N_865,N_4536);
nand U7738 (N_7738,N_536,N_3383);
or U7739 (N_7739,N_639,N_824);
nor U7740 (N_7740,N_636,N_2811);
or U7741 (N_7741,N_551,N_3314);
xnor U7742 (N_7742,N_2490,N_1307);
nand U7743 (N_7743,N_1537,N_1400);
or U7744 (N_7744,N_1472,N_4684);
xor U7745 (N_7745,N_1426,N_2225);
nor U7746 (N_7746,N_3265,N_4176);
and U7747 (N_7747,N_1129,N_1436);
nand U7748 (N_7748,N_502,N_139);
and U7749 (N_7749,N_1539,N_2157);
nor U7750 (N_7750,N_3919,N_559);
and U7751 (N_7751,N_327,N_3683);
or U7752 (N_7752,N_1878,N_4998);
xnor U7753 (N_7753,N_180,N_914);
and U7754 (N_7754,N_2167,N_67);
nand U7755 (N_7755,N_3818,N_4432);
and U7756 (N_7756,N_3120,N_367);
nand U7757 (N_7757,N_4587,N_2043);
or U7758 (N_7758,N_4835,N_1707);
nor U7759 (N_7759,N_4519,N_2799);
nor U7760 (N_7760,N_2233,N_1479);
xor U7761 (N_7761,N_2962,N_2184);
or U7762 (N_7762,N_2216,N_3766);
nand U7763 (N_7763,N_1371,N_1464);
nand U7764 (N_7764,N_4789,N_2262);
xor U7765 (N_7765,N_287,N_4513);
or U7766 (N_7766,N_2344,N_3437);
nand U7767 (N_7767,N_2526,N_958);
nand U7768 (N_7768,N_770,N_589);
and U7769 (N_7769,N_3172,N_2912);
and U7770 (N_7770,N_3122,N_2857);
and U7771 (N_7771,N_128,N_2194);
and U7772 (N_7772,N_1792,N_973);
nand U7773 (N_7773,N_4730,N_2711);
and U7774 (N_7774,N_573,N_454);
or U7775 (N_7775,N_3526,N_3265);
and U7776 (N_7776,N_2736,N_1596);
or U7777 (N_7777,N_3153,N_2415);
or U7778 (N_7778,N_1736,N_2683);
nor U7779 (N_7779,N_3505,N_4569);
nor U7780 (N_7780,N_1129,N_594);
nor U7781 (N_7781,N_4376,N_1459);
or U7782 (N_7782,N_4862,N_86);
xnor U7783 (N_7783,N_2742,N_1572);
or U7784 (N_7784,N_4273,N_3419);
or U7785 (N_7785,N_3375,N_1115);
or U7786 (N_7786,N_4010,N_624);
or U7787 (N_7787,N_3133,N_2309);
or U7788 (N_7788,N_3741,N_3566);
and U7789 (N_7789,N_3322,N_1596);
nand U7790 (N_7790,N_2040,N_4114);
nor U7791 (N_7791,N_2465,N_3345);
nor U7792 (N_7792,N_1099,N_771);
xnor U7793 (N_7793,N_4964,N_3521);
nor U7794 (N_7794,N_1405,N_880);
nand U7795 (N_7795,N_3270,N_375);
nor U7796 (N_7796,N_1608,N_273);
or U7797 (N_7797,N_1501,N_3968);
xnor U7798 (N_7798,N_1420,N_4727);
nand U7799 (N_7799,N_1952,N_4193);
nor U7800 (N_7800,N_648,N_1469);
or U7801 (N_7801,N_4913,N_958);
or U7802 (N_7802,N_998,N_106);
nor U7803 (N_7803,N_1799,N_2131);
nand U7804 (N_7804,N_838,N_3105);
and U7805 (N_7805,N_988,N_68);
nor U7806 (N_7806,N_2419,N_2641);
nor U7807 (N_7807,N_2756,N_1265);
nor U7808 (N_7808,N_4191,N_2412);
or U7809 (N_7809,N_3464,N_3384);
nor U7810 (N_7810,N_1014,N_3196);
xor U7811 (N_7811,N_712,N_1828);
nor U7812 (N_7812,N_1149,N_4237);
or U7813 (N_7813,N_4797,N_3838);
xnor U7814 (N_7814,N_4048,N_4756);
and U7815 (N_7815,N_2482,N_3627);
or U7816 (N_7816,N_3993,N_1581);
and U7817 (N_7817,N_1669,N_1956);
xor U7818 (N_7818,N_2576,N_3120);
nand U7819 (N_7819,N_4603,N_3235);
nand U7820 (N_7820,N_2530,N_2220);
nand U7821 (N_7821,N_2046,N_3093);
or U7822 (N_7822,N_2977,N_3426);
nand U7823 (N_7823,N_1345,N_4826);
and U7824 (N_7824,N_109,N_827);
or U7825 (N_7825,N_4252,N_4972);
or U7826 (N_7826,N_3609,N_4788);
nand U7827 (N_7827,N_4254,N_1640);
nand U7828 (N_7828,N_495,N_2838);
or U7829 (N_7829,N_3212,N_4994);
or U7830 (N_7830,N_4404,N_102);
and U7831 (N_7831,N_766,N_2034);
or U7832 (N_7832,N_838,N_2885);
or U7833 (N_7833,N_855,N_2525);
or U7834 (N_7834,N_4866,N_3984);
xor U7835 (N_7835,N_4750,N_2327);
nand U7836 (N_7836,N_3533,N_3001);
and U7837 (N_7837,N_4833,N_4618);
nor U7838 (N_7838,N_3626,N_4537);
or U7839 (N_7839,N_4828,N_1105);
or U7840 (N_7840,N_2582,N_1066);
nor U7841 (N_7841,N_3136,N_2484);
nand U7842 (N_7842,N_1033,N_3112);
nand U7843 (N_7843,N_4753,N_79);
or U7844 (N_7844,N_186,N_4174);
or U7845 (N_7845,N_2366,N_1969);
nor U7846 (N_7846,N_1839,N_4200);
and U7847 (N_7847,N_2926,N_2844);
or U7848 (N_7848,N_4725,N_4447);
or U7849 (N_7849,N_3321,N_1400);
nor U7850 (N_7850,N_2465,N_4792);
and U7851 (N_7851,N_4487,N_308);
xor U7852 (N_7852,N_330,N_3097);
nor U7853 (N_7853,N_3681,N_3764);
and U7854 (N_7854,N_3557,N_4466);
or U7855 (N_7855,N_379,N_501);
or U7856 (N_7856,N_4377,N_1510);
and U7857 (N_7857,N_872,N_4036);
nand U7858 (N_7858,N_3173,N_1948);
nor U7859 (N_7859,N_1835,N_746);
or U7860 (N_7860,N_760,N_3296);
nand U7861 (N_7861,N_3565,N_4312);
nand U7862 (N_7862,N_4418,N_2111);
nand U7863 (N_7863,N_4037,N_4203);
or U7864 (N_7864,N_1598,N_3890);
nor U7865 (N_7865,N_479,N_1848);
or U7866 (N_7866,N_4911,N_3801);
or U7867 (N_7867,N_3843,N_2899);
and U7868 (N_7868,N_2850,N_2494);
nand U7869 (N_7869,N_720,N_4950);
nand U7870 (N_7870,N_2086,N_3396);
nand U7871 (N_7871,N_3503,N_475);
and U7872 (N_7872,N_4777,N_2229);
nand U7873 (N_7873,N_1538,N_1366);
xnor U7874 (N_7874,N_2813,N_288);
xor U7875 (N_7875,N_2888,N_319);
nor U7876 (N_7876,N_4981,N_1974);
nand U7877 (N_7877,N_2795,N_3872);
nand U7878 (N_7878,N_207,N_3804);
or U7879 (N_7879,N_845,N_2196);
and U7880 (N_7880,N_2671,N_1283);
and U7881 (N_7881,N_4404,N_3041);
or U7882 (N_7882,N_957,N_486);
or U7883 (N_7883,N_1643,N_917);
or U7884 (N_7884,N_13,N_2289);
or U7885 (N_7885,N_3118,N_205);
nor U7886 (N_7886,N_3735,N_703);
nor U7887 (N_7887,N_3600,N_3770);
nand U7888 (N_7888,N_95,N_2369);
or U7889 (N_7889,N_2936,N_1108);
nor U7890 (N_7890,N_3079,N_2567);
nand U7891 (N_7891,N_3501,N_4522);
and U7892 (N_7892,N_2168,N_1475);
and U7893 (N_7893,N_2919,N_4443);
and U7894 (N_7894,N_740,N_2481);
and U7895 (N_7895,N_4219,N_4687);
nor U7896 (N_7896,N_2184,N_3200);
or U7897 (N_7897,N_200,N_1577);
or U7898 (N_7898,N_1578,N_3440);
or U7899 (N_7899,N_1444,N_2963);
nor U7900 (N_7900,N_4972,N_344);
or U7901 (N_7901,N_908,N_1238);
or U7902 (N_7902,N_4123,N_583);
nand U7903 (N_7903,N_2124,N_4088);
nor U7904 (N_7904,N_168,N_3533);
nand U7905 (N_7905,N_1567,N_3960);
or U7906 (N_7906,N_4355,N_3234);
and U7907 (N_7907,N_3665,N_4255);
and U7908 (N_7908,N_4713,N_1760);
nand U7909 (N_7909,N_2288,N_3162);
xnor U7910 (N_7910,N_4949,N_4328);
nor U7911 (N_7911,N_3096,N_2412);
or U7912 (N_7912,N_4206,N_2065);
nand U7913 (N_7913,N_123,N_705);
and U7914 (N_7914,N_4134,N_1027);
nor U7915 (N_7915,N_4092,N_3023);
and U7916 (N_7916,N_4981,N_23);
and U7917 (N_7917,N_4027,N_4916);
or U7918 (N_7918,N_3641,N_3062);
nor U7919 (N_7919,N_2,N_688);
nand U7920 (N_7920,N_2590,N_1837);
nand U7921 (N_7921,N_4107,N_3709);
xnor U7922 (N_7922,N_2716,N_3033);
nor U7923 (N_7923,N_1223,N_3362);
nand U7924 (N_7924,N_1642,N_4651);
nor U7925 (N_7925,N_4645,N_4493);
nand U7926 (N_7926,N_3649,N_1269);
nand U7927 (N_7927,N_2992,N_2850);
nand U7928 (N_7928,N_792,N_1597);
nand U7929 (N_7929,N_1890,N_4315);
nor U7930 (N_7930,N_3945,N_497);
and U7931 (N_7931,N_2957,N_4589);
nor U7932 (N_7932,N_2024,N_50);
nand U7933 (N_7933,N_709,N_2461);
nand U7934 (N_7934,N_4168,N_772);
nand U7935 (N_7935,N_258,N_885);
or U7936 (N_7936,N_1418,N_2210);
or U7937 (N_7937,N_180,N_4619);
or U7938 (N_7938,N_4913,N_2915);
nor U7939 (N_7939,N_3370,N_4078);
and U7940 (N_7940,N_3387,N_999);
or U7941 (N_7941,N_2421,N_2298);
nand U7942 (N_7942,N_245,N_315);
nand U7943 (N_7943,N_1573,N_2373);
nor U7944 (N_7944,N_4680,N_337);
nand U7945 (N_7945,N_2338,N_391);
and U7946 (N_7946,N_2038,N_2488);
nor U7947 (N_7947,N_3386,N_541);
nor U7948 (N_7948,N_3750,N_3462);
and U7949 (N_7949,N_1758,N_360);
nor U7950 (N_7950,N_303,N_3833);
nand U7951 (N_7951,N_2858,N_2749);
nand U7952 (N_7952,N_4090,N_3134);
xor U7953 (N_7953,N_2182,N_4981);
xor U7954 (N_7954,N_194,N_152);
nor U7955 (N_7955,N_1878,N_406);
nor U7956 (N_7956,N_3958,N_2268);
and U7957 (N_7957,N_2848,N_633);
nor U7958 (N_7958,N_1635,N_4762);
and U7959 (N_7959,N_1789,N_4813);
and U7960 (N_7960,N_2318,N_920);
and U7961 (N_7961,N_348,N_4887);
nor U7962 (N_7962,N_2043,N_4764);
nor U7963 (N_7963,N_2290,N_2667);
nor U7964 (N_7964,N_1025,N_4300);
and U7965 (N_7965,N_2402,N_3321);
and U7966 (N_7966,N_4043,N_4684);
or U7967 (N_7967,N_602,N_84);
and U7968 (N_7968,N_2299,N_4114);
nand U7969 (N_7969,N_3295,N_2487);
xor U7970 (N_7970,N_2543,N_3692);
nor U7971 (N_7971,N_536,N_1183);
or U7972 (N_7972,N_4785,N_1944);
nor U7973 (N_7973,N_2192,N_4711);
nor U7974 (N_7974,N_3388,N_1288);
or U7975 (N_7975,N_4687,N_4434);
nor U7976 (N_7976,N_1243,N_4608);
or U7977 (N_7977,N_1207,N_298);
or U7978 (N_7978,N_4202,N_3901);
nor U7979 (N_7979,N_4665,N_463);
nor U7980 (N_7980,N_1169,N_4132);
nor U7981 (N_7981,N_1497,N_18);
and U7982 (N_7982,N_4608,N_3208);
nor U7983 (N_7983,N_3474,N_545);
nor U7984 (N_7984,N_3561,N_1403);
nand U7985 (N_7985,N_3314,N_1081);
nor U7986 (N_7986,N_2068,N_3001);
nand U7987 (N_7987,N_3074,N_1833);
or U7988 (N_7988,N_2230,N_1777);
xor U7989 (N_7989,N_552,N_2037);
nor U7990 (N_7990,N_1484,N_967);
nand U7991 (N_7991,N_1772,N_2992);
nor U7992 (N_7992,N_2862,N_4437);
and U7993 (N_7993,N_4111,N_335);
xor U7994 (N_7994,N_2552,N_318);
and U7995 (N_7995,N_3257,N_1055);
or U7996 (N_7996,N_3568,N_1501);
nor U7997 (N_7997,N_1211,N_1395);
or U7998 (N_7998,N_4950,N_2197);
xor U7999 (N_7999,N_4214,N_2149);
nand U8000 (N_8000,N_1449,N_4446);
nand U8001 (N_8001,N_3867,N_4333);
nor U8002 (N_8002,N_1251,N_2883);
and U8003 (N_8003,N_3430,N_4994);
nor U8004 (N_8004,N_347,N_1908);
and U8005 (N_8005,N_553,N_1057);
and U8006 (N_8006,N_2342,N_4742);
and U8007 (N_8007,N_649,N_1236);
nor U8008 (N_8008,N_3130,N_3716);
nor U8009 (N_8009,N_4996,N_3783);
xor U8010 (N_8010,N_3703,N_525);
or U8011 (N_8011,N_2768,N_4336);
nand U8012 (N_8012,N_1642,N_2261);
and U8013 (N_8013,N_3771,N_1282);
nor U8014 (N_8014,N_1964,N_839);
nand U8015 (N_8015,N_4921,N_170);
nor U8016 (N_8016,N_628,N_1487);
xor U8017 (N_8017,N_3287,N_4244);
nor U8018 (N_8018,N_3249,N_3925);
or U8019 (N_8019,N_229,N_122);
xor U8020 (N_8020,N_3980,N_637);
or U8021 (N_8021,N_3797,N_3985);
or U8022 (N_8022,N_4634,N_926);
nand U8023 (N_8023,N_3981,N_3826);
and U8024 (N_8024,N_1891,N_2671);
and U8025 (N_8025,N_633,N_4676);
nand U8026 (N_8026,N_2845,N_438);
and U8027 (N_8027,N_4392,N_2536);
nand U8028 (N_8028,N_719,N_1773);
nor U8029 (N_8029,N_4499,N_3142);
and U8030 (N_8030,N_4531,N_3341);
and U8031 (N_8031,N_611,N_4398);
nand U8032 (N_8032,N_4724,N_3530);
nor U8033 (N_8033,N_741,N_3673);
nand U8034 (N_8034,N_382,N_2801);
nor U8035 (N_8035,N_4536,N_1026);
and U8036 (N_8036,N_788,N_760);
and U8037 (N_8037,N_4031,N_2084);
xnor U8038 (N_8038,N_1247,N_2414);
nor U8039 (N_8039,N_375,N_1488);
and U8040 (N_8040,N_1036,N_1169);
and U8041 (N_8041,N_2065,N_171);
nor U8042 (N_8042,N_4115,N_4779);
and U8043 (N_8043,N_370,N_4233);
and U8044 (N_8044,N_175,N_667);
nand U8045 (N_8045,N_1718,N_37);
nor U8046 (N_8046,N_3101,N_3439);
or U8047 (N_8047,N_3419,N_3180);
or U8048 (N_8048,N_1523,N_2718);
nand U8049 (N_8049,N_4946,N_4246);
or U8050 (N_8050,N_780,N_3406);
and U8051 (N_8051,N_1372,N_437);
nor U8052 (N_8052,N_3424,N_147);
nand U8053 (N_8053,N_1645,N_727);
nor U8054 (N_8054,N_4402,N_1146);
or U8055 (N_8055,N_3609,N_2854);
nor U8056 (N_8056,N_4910,N_808);
or U8057 (N_8057,N_2035,N_3884);
and U8058 (N_8058,N_2118,N_1544);
or U8059 (N_8059,N_4293,N_968);
nand U8060 (N_8060,N_3332,N_1586);
or U8061 (N_8061,N_4794,N_3179);
xnor U8062 (N_8062,N_1679,N_4927);
nor U8063 (N_8063,N_4514,N_25);
xnor U8064 (N_8064,N_2039,N_1991);
nor U8065 (N_8065,N_1375,N_1511);
or U8066 (N_8066,N_2850,N_4596);
nand U8067 (N_8067,N_2576,N_4970);
or U8068 (N_8068,N_2515,N_4348);
nor U8069 (N_8069,N_2588,N_4295);
xor U8070 (N_8070,N_2627,N_3907);
nand U8071 (N_8071,N_1619,N_61);
nand U8072 (N_8072,N_3873,N_1627);
nor U8073 (N_8073,N_4593,N_3260);
or U8074 (N_8074,N_2967,N_959);
nand U8075 (N_8075,N_4804,N_2188);
nand U8076 (N_8076,N_1210,N_3823);
nand U8077 (N_8077,N_1227,N_1126);
nand U8078 (N_8078,N_3008,N_2702);
xor U8079 (N_8079,N_1194,N_3808);
nand U8080 (N_8080,N_1190,N_2506);
nand U8081 (N_8081,N_1831,N_2471);
or U8082 (N_8082,N_1415,N_3608);
xor U8083 (N_8083,N_3929,N_4641);
nand U8084 (N_8084,N_4898,N_4381);
nand U8085 (N_8085,N_3986,N_3260);
or U8086 (N_8086,N_1983,N_2226);
nor U8087 (N_8087,N_816,N_1708);
or U8088 (N_8088,N_4639,N_33);
xor U8089 (N_8089,N_1693,N_537);
nor U8090 (N_8090,N_983,N_4351);
or U8091 (N_8091,N_152,N_292);
nor U8092 (N_8092,N_3305,N_395);
or U8093 (N_8093,N_4711,N_1632);
xnor U8094 (N_8094,N_1021,N_2011);
nand U8095 (N_8095,N_860,N_4705);
nor U8096 (N_8096,N_968,N_3655);
xor U8097 (N_8097,N_4101,N_4064);
or U8098 (N_8098,N_925,N_2106);
nor U8099 (N_8099,N_3484,N_720);
or U8100 (N_8100,N_2508,N_2619);
or U8101 (N_8101,N_642,N_1568);
or U8102 (N_8102,N_1835,N_1707);
or U8103 (N_8103,N_2829,N_3495);
and U8104 (N_8104,N_4018,N_3419);
and U8105 (N_8105,N_2953,N_2485);
or U8106 (N_8106,N_2941,N_2580);
or U8107 (N_8107,N_4357,N_666);
and U8108 (N_8108,N_4035,N_3929);
and U8109 (N_8109,N_1139,N_2025);
and U8110 (N_8110,N_3595,N_3983);
and U8111 (N_8111,N_4559,N_978);
nand U8112 (N_8112,N_1442,N_4198);
or U8113 (N_8113,N_4820,N_2570);
and U8114 (N_8114,N_284,N_2089);
or U8115 (N_8115,N_1571,N_1615);
and U8116 (N_8116,N_3879,N_2227);
or U8117 (N_8117,N_1498,N_1393);
nand U8118 (N_8118,N_2063,N_427);
and U8119 (N_8119,N_4900,N_2391);
and U8120 (N_8120,N_200,N_931);
nand U8121 (N_8121,N_4061,N_4226);
and U8122 (N_8122,N_3824,N_2697);
and U8123 (N_8123,N_795,N_3835);
nor U8124 (N_8124,N_2793,N_2322);
nor U8125 (N_8125,N_1494,N_2656);
nor U8126 (N_8126,N_2245,N_4158);
nor U8127 (N_8127,N_3532,N_1634);
and U8128 (N_8128,N_4214,N_3385);
or U8129 (N_8129,N_2581,N_2788);
nor U8130 (N_8130,N_4440,N_1996);
nand U8131 (N_8131,N_461,N_2485);
nor U8132 (N_8132,N_2574,N_3350);
or U8133 (N_8133,N_1153,N_4072);
xor U8134 (N_8134,N_4846,N_4262);
nand U8135 (N_8135,N_1748,N_960);
nand U8136 (N_8136,N_2068,N_4383);
or U8137 (N_8137,N_3403,N_2701);
nand U8138 (N_8138,N_731,N_3018);
and U8139 (N_8139,N_810,N_1565);
nor U8140 (N_8140,N_4375,N_4213);
and U8141 (N_8141,N_3474,N_2537);
xor U8142 (N_8142,N_512,N_1426);
nand U8143 (N_8143,N_126,N_1948);
nor U8144 (N_8144,N_3230,N_837);
and U8145 (N_8145,N_1391,N_1579);
and U8146 (N_8146,N_3887,N_2741);
nand U8147 (N_8147,N_1731,N_2389);
and U8148 (N_8148,N_2520,N_4881);
or U8149 (N_8149,N_3971,N_1976);
nand U8150 (N_8150,N_2687,N_2746);
xnor U8151 (N_8151,N_1456,N_1826);
nor U8152 (N_8152,N_2055,N_2047);
nand U8153 (N_8153,N_4854,N_3466);
nor U8154 (N_8154,N_2294,N_2052);
and U8155 (N_8155,N_1728,N_886);
nor U8156 (N_8156,N_1553,N_2373);
nand U8157 (N_8157,N_3730,N_4622);
nand U8158 (N_8158,N_1602,N_480);
nor U8159 (N_8159,N_1224,N_66);
nand U8160 (N_8160,N_1472,N_4489);
and U8161 (N_8161,N_102,N_3483);
xor U8162 (N_8162,N_4795,N_1142);
nand U8163 (N_8163,N_4234,N_930);
nand U8164 (N_8164,N_1502,N_1034);
nand U8165 (N_8165,N_1711,N_2906);
and U8166 (N_8166,N_692,N_3923);
and U8167 (N_8167,N_4376,N_665);
xnor U8168 (N_8168,N_3080,N_2137);
xor U8169 (N_8169,N_625,N_1900);
and U8170 (N_8170,N_3416,N_4862);
or U8171 (N_8171,N_2568,N_2611);
xnor U8172 (N_8172,N_2901,N_2388);
or U8173 (N_8173,N_240,N_1001);
or U8174 (N_8174,N_243,N_1278);
nor U8175 (N_8175,N_29,N_4022);
nor U8176 (N_8176,N_1998,N_3899);
nand U8177 (N_8177,N_671,N_302);
or U8178 (N_8178,N_4836,N_1387);
nand U8179 (N_8179,N_815,N_1145);
nand U8180 (N_8180,N_1647,N_2555);
or U8181 (N_8181,N_4814,N_2366);
nor U8182 (N_8182,N_2497,N_4802);
and U8183 (N_8183,N_927,N_2366);
nor U8184 (N_8184,N_3403,N_2491);
and U8185 (N_8185,N_2923,N_4077);
nor U8186 (N_8186,N_552,N_4995);
nand U8187 (N_8187,N_4202,N_3371);
nor U8188 (N_8188,N_4465,N_2101);
or U8189 (N_8189,N_575,N_3482);
or U8190 (N_8190,N_3670,N_4639);
nand U8191 (N_8191,N_718,N_4253);
or U8192 (N_8192,N_2862,N_206);
nor U8193 (N_8193,N_3154,N_758);
nand U8194 (N_8194,N_1376,N_101);
nand U8195 (N_8195,N_1761,N_4220);
and U8196 (N_8196,N_897,N_1347);
and U8197 (N_8197,N_1268,N_2922);
nand U8198 (N_8198,N_4438,N_2058);
and U8199 (N_8199,N_2111,N_3746);
or U8200 (N_8200,N_1192,N_988);
xnor U8201 (N_8201,N_3595,N_2938);
and U8202 (N_8202,N_89,N_3070);
nand U8203 (N_8203,N_2777,N_793);
or U8204 (N_8204,N_4747,N_187);
xor U8205 (N_8205,N_2826,N_3320);
nand U8206 (N_8206,N_3290,N_1615);
or U8207 (N_8207,N_1015,N_3111);
and U8208 (N_8208,N_2872,N_3586);
nand U8209 (N_8209,N_1982,N_395);
nor U8210 (N_8210,N_1476,N_4993);
nand U8211 (N_8211,N_4531,N_1338);
nor U8212 (N_8212,N_4260,N_3303);
xnor U8213 (N_8213,N_4134,N_485);
xnor U8214 (N_8214,N_2956,N_321);
nand U8215 (N_8215,N_2882,N_2044);
or U8216 (N_8216,N_119,N_3541);
and U8217 (N_8217,N_3372,N_336);
and U8218 (N_8218,N_559,N_2310);
and U8219 (N_8219,N_4475,N_1448);
nor U8220 (N_8220,N_517,N_4236);
or U8221 (N_8221,N_829,N_4980);
or U8222 (N_8222,N_1025,N_524);
nand U8223 (N_8223,N_332,N_693);
or U8224 (N_8224,N_4483,N_85);
nand U8225 (N_8225,N_4429,N_2773);
xnor U8226 (N_8226,N_4575,N_2423);
nand U8227 (N_8227,N_1485,N_3898);
nand U8228 (N_8228,N_2044,N_741);
nand U8229 (N_8229,N_4807,N_4570);
nor U8230 (N_8230,N_2712,N_1700);
nor U8231 (N_8231,N_4374,N_3890);
nand U8232 (N_8232,N_1203,N_473);
nor U8233 (N_8233,N_1871,N_2149);
nand U8234 (N_8234,N_4842,N_4195);
or U8235 (N_8235,N_2549,N_3);
nand U8236 (N_8236,N_2404,N_2472);
or U8237 (N_8237,N_4684,N_4306);
or U8238 (N_8238,N_4627,N_3200);
nor U8239 (N_8239,N_2090,N_3894);
xnor U8240 (N_8240,N_3264,N_4201);
nor U8241 (N_8241,N_1579,N_1534);
nand U8242 (N_8242,N_4730,N_859);
nand U8243 (N_8243,N_2325,N_37);
nand U8244 (N_8244,N_2648,N_49);
nor U8245 (N_8245,N_13,N_4840);
nand U8246 (N_8246,N_2809,N_4015);
and U8247 (N_8247,N_4219,N_4290);
nand U8248 (N_8248,N_3805,N_82);
nor U8249 (N_8249,N_909,N_37);
and U8250 (N_8250,N_2519,N_1882);
or U8251 (N_8251,N_2101,N_2039);
nor U8252 (N_8252,N_1004,N_263);
nor U8253 (N_8253,N_1516,N_3833);
or U8254 (N_8254,N_2250,N_2645);
nand U8255 (N_8255,N_3468,N_3928);
and U8256 (N_8256,N_355,N_4111);
and U8257 (N_8257,N_24,N_1703);
and U8258 (N_8258,N_2416,N_819);
nor U8259 (N_8259,N_1768,N_3058);
xor U8260 (N_8260,N_2173,N_1950);
nor U8261 (N_8261,N_381,N_2996);
or U8262 (N_8262,N_3547,N_1195);
or U8263 (N_8263,N_1808,N_1159);
nor U8264 (N_8264,N_1424,N_3690);
nand U8265 (N_8265,N_3583,N_1059);
nand U8266 (N_8266,N_2729,N_1190);
nand U8267 (N_8267,N_3067,N_1049);
xor U8268 (N_8268,N_4117,N_3270);
and U8269 (N_8269,N_1823,N_2892);
xnor U8270 (N_8270,N_3088,N_3082);
xnor U8271 (N_8271,N_3327,N_2965);
or U8272 (N_8272,N_3750,N_1209);
or U8273 (N_8273,N_2698,N_306);
or U8274 (N_8274,N_2352,N_3821);
nand U8275 (N_8275,N_665,N_1334);
xnor U8276 (N_8276,N_4388,N_4463);
nand U8277 (N_8277,N_4985,N_4038);
nor U8278 (N_8278,N_54,N_285);
nand U8279 (N_8279,N_3481,N_1028);
nand U8280 (N_8280,N_3994,N_4557);
nor U8281 (N_8281,N_4010,N_2709);
nand U8282 (N_8282,N_85,N_2214);
nand U8283 (N_8283,N_1487,N_173);
nand U8284 (N_8284,N_2767,N_1437);
nand U8285 (N_8285,N_2024,N_1280);
nor U8286 (N_8286,N_495,N_3336);
nand U8287 (N_8287,N_2557,N_1727);
or U8288 (N_8288,N_1587,N_4386);
nand U8289 (N_8289,N_4197,N_938);
and U8290 (N_8290,N_2685,N_4334);
nand U8291 (N_8291,N_4299,N_3877);
or U8292 (N_8292,N_3968,N_1353);
xor U8293 (N_8293,N_3578,N_3184);
or U8294 (N_8294,N_669,N_2383);
nand U8295 (N_8295,N_1842,N_4500);
nand U8296 (N_8296,N_3766,N_3706);
and U8297 (N_8297,N_447,N_1580);
nor U8298 (N_8298,N_4955,N_1970);
or U8299 (N_8299,N_4988,N_3322);
and U8300 (N_8300,N_1553,N_4350);
and U8301 (N_8301,N_4521,N_430);
nand U8302 (N_8302,N_1231,N_197);
nor U8303 (N_8303,N_4282,N_3407);
or U8304 (N_8304,N_4637,N_672);
and U8305 (N_8305,N_2463,N_173);
and U8306 (N_8306,N_2607,N_2068);
nand U8307 (N_8307,N_4232,N_3579);
and U8308 (N_8308,N_835,N_286);
nand U8309 (N_8309,N_3983,N_1660);
nor U8310 (N_8310,N_4409,N_803);
xor U8311 (N_8311,N_2252,N_344);
nor U8312 (N_8312,N_344,N_384);
nor U8313 (N_8313,N_1992,N_1300);
nand U8314 (N_8314,N_4445,N_919);
and U8315 (N_8315,N_4342,N_749);
nand U8316 (N_8316,N_321,N_4380);
and U8317 (N_8317,N_1135,N_2176);
or U8318 (N_8318,N_1523,N_4488);
and U8319 (N_8319,N_1756,N_4506);
nand U8320 (N_8320,N_1103,N_1334);
nor U8321 (N_8321,N_1102,N_755);
nand U8322 (N_8322,N_4602,N_66);
or U8323 (N_8323,N_2934,N_1606);
and U8324 (N_8324,N_305,N_4011);
and U8325 (N_8325,N_3610,N_3506);
and U8326 (N_8326,N_4986,N_4702);
nand U8327 (N_8327,N_4196,N_2668);
or U8328 (N_8328,N_4964,N_1884);
nor U8329 (N_8329,N_3031,N_2891);
nor U8330 (N_8330,N_1504,N_1426);
or U8331 (N_8331,N_2785,N_1264);
nand U8332 (N_8332,N_441,N_4478);
nand U8333 (N_8333,N_35,N_4582);
nand U8334 (N_8334,N_2113,N_4960);
or U8335 (N_8335,N_4365,N_2421);
and U8336 (N_8336,N_1028,N_377);
xnor U8337 (N_8337,N_2361,N_2618);
nor U8338 (N_8338,N_3410,N_4525);
and U8339 (N_8339,N_3292,N_3343);
nand U8340 (N_8340,N_4468,N_3147);
or U8341 (N_8341,N_597,N_4338);
and U8342 (N_8342,N_3395,N_3602);
or U8343 (N_8343,N_1649,N_1982);
xnor U8344 (N_8344,N_4786,N_3214);
nor U8345 (N_8345,N_1818,N_1384);
or U8346 (N_8346,N_1713,N_960);
or U8347 (N_8347,N_207,N_2130);
nor U8348 (N_8348,N_1821,N_3722);
nand U8349 (N_8349,N_3788,N_391);
nor U8350 (N_8350,N_3810,N_3348);
and U8351 (N_8351,N_1845,N_780);
or U8352 (N_8352,N_4751,N_4473);
nor U8353 (N_8353,N_2818,N_2426);
or U8354 (N_8354,N_3432,N_763);
nor U8355 (N_8355,N_1321,N_3976);
or U8356 (N_8356,N_3951,N_1936);
and U8357 (N_8357,N_1272,N_3938);
xnor U8358 (N_8358,N_298,N_2380);
nand U8359 (N_8359,N_652,N_1110);
nor U8360 (N_8360,N_3843,N_900);
and U8361 (N_8361,N_3034,N_1079);
and U8362 (N_8362,N_912,N_4697);
nand U8363 (N_8363,N_3135,N_1834);
nor U8364 (N_8364,N_2654,N_590);
nor U8365 (N_8365,N_2363,N_866);
or U8366 (N_8366,N_4492,N_573);
nor U8367 (N_8367,N_1951,N_163);
and U8368 (N_8368,N_3909,N_3607);
and U8369 (N_8369,N_654,N_2765);
or U8370 (N_8370,N_4648,N_890);
nand U8371 (N_8371,N_774,N_2941);
nor U8372 (N_8372,N_4156,N_3324);
and U8373 (N_8373,N_4379,N_338);
or U8374 (N_8374,N_4898,N_4580);
nor U8375 (N_8375,N_2489,N_4495);
or U8376 (N_8376,N_4117,N_3886);
or U8377 (N_8377,N_81,N_2754);
nor U8378 (N_8378,N_2203,N_1111);
nand U8379 (N_8379,N_530,N_4281);
xor U8380 (N_8380,N_4887,N_3891);
and U8381 (N_8381,N_872,N_4046);
and U8382 (N_8382,N_3642,N_4734);
or U8383 (N_8383,N_656,N_1615);
and U8384 (N_8384,N_3,N_2211);
or U8385 (N_8385,N_1970,N_4172);
and U8386 (N_8386,N_1972,N_2667);
nand U8387 (N_8387,N_4445,N_833);
nor U8388 (N_8388,N_754,N_2199);
or U8389 (N_8389,N_578,N_2387);
xor U8390 (N_8390,N_2017,N_322);
nand U8391 (N_8391,N_2048,N_853);
or U8392 (N_8392,N_4400,N_1763);
xnor U8393 (N_8393,N_3583,N_2521);
and U8394 (N_8394,N_987,N_423);
xor U8395 (N_8395,N_775,N_1185);
nor U8396 (N_8396,N_3820,N_4081);
and U8397 (N_8397,N_842,N_4671);
nand U8398 (N_8398,N_3221,N_3774);
or U8399 (N_8399,N_1614,N_2534);
and U8400 (N_8400,N_4255,N_2333);
or U8401 (N_8401,N_4802,N_1465);
xnor U8402 (N_8402,N_731,N_1549);
nand U8403 (N_8403,N_2083,N_3792);
or U8404 (N_8404,N_1019,N_3553);
nand U8405 (N_8405,N_3613,N_2680);
or U8406 (N_8406,N_3827,N_975);
nand U8407 (N_8407,N_3911,N_1995);
or U8408 (N_8408,N_885,N_505);
nor U8409 (N_8409,N_3425,N_2868);
xor U8410 (N_8410,N_1139,N_3478);
nor U8411 (N_8411,N_4608,N_1010);
xnor U8412 (N_8412,N_4424,N_4378);
nand U8413 (N_8413,N_4858,N_2911);
nand U8414 (N_8414,N_4616,N_2888);
or U8415 (N_8415,N_1475,N_3028);
nor U8416 (N_8416,N_638,N_2362);
and U8417 (N_8417,N_2090,N_841);
or U8418 (N_8418,N_4980,N_3505);
nand U8419 (N_8419,N_624,N_122);
nor U8420 (N_8420,N_2606,N_1280);
and U8421 (N_8421,N_399,N_1756);
and U8422 (N_8422,N_4326,N_2749);
nor U8423 (N_8423,N_2049,N_705);
nor U8424 (N_8424,N_4770,N_3498);
nor U8425 (N_8425,N_4714,N_4019);
or U8426 (N_8426,N_3382,N_4507);
or U8427 (N_8427,N_99,N_834);
or U8428 (N_8428,N_2680,N_649);
and U8429 (N_8429,N_1679,N_1001);
nand U8430 (N_8430,N_1158,N_501);
nor U8431 (N_8431,N_715,N_1676);
and U8432 (N_8432,N_1402,N_98);
and U8433 (N_8433,N_2599,N_4512);
nand U8434 (N_8434,N_816,N_2488);
and U8435 (N_8435,N_2459,N_3303);
nand U8436 (N_8436,N_3893,N_4561);
or U8437 (N_8437,N_477,N_316);
nand U8438 (N_8438,N_4752,N_4211);
nor U8439 (N_8439,N_2983,N_2753);
nand U8440 (N_8440,N_3729,N_4891);
and U8441 (N_8441,N_1002,N_15);
or U8442 (N_8442,N_56,N_4752);
nor U8443 (N_8443,N_3969,N_4498);
nand U8444 (N_8444,N_4909,N_4559);
and U8445 (N_8445,N_2582,N_461);
nand U8446 (N_8446,N_4889,N_3761);
and U8447 (N_8447,N_1829,N_279);
and U8448 (N_8448,N_3308,N_1006);
and U8449 (N_8449,N_3115,N_3611);
nor U8450 (N_8450,N_31,N_2463);
nand U8451 (N_8451,N_4722,N_121);
or U8452 (N_8452,N_4991,N_3401);
and U8453 (N_8453,N_2740,N_2187);
nor U8454 (N_8454,N_2317,N_4763);
and U8455 (N_8455,N_4412,N_2143);
and U8456 (N_8456,N_2020,N_952);
nand U8457 (N_8457,N_532,N_3883);
nand U8458 (N_8458,N_4823,N_386);
or U8459 (N_8459,N_3428,N_3418);
or U8460 (N_8460,N_551,N_4865);
and U8461 (N_8461,N_2292,N_884);
or U8462 (N_8462,N_4039,N_3543);
nand U8463 (N_8463,N_1800,N_2222);
nand U8464 (N_8464,N_1201,N_1888);
nor U8465 (N_8465,N_2876,N_4089);
nand U8466 (N_8466,N_949,N_4960);
and U8467 (N_8467,N_2882,N_525);
nor U8468 (N_8468,N_1239,N_3475);
nor U8469 (N_8469,N_3436,N_3422);
xor U8470 (N_8470,N_2509,N_4169);
or U8471 (N_8471,N_523,N_1199);
nor U8472 (N_8472,N_3553,N_3068);
or U8473 (N_8473,N_191,N_1548);
nor U8474 (N_8474,N_1356,N_2307);
and U8475 (N_8475,N_453,N_2769);
and U8476 (N_8476,N_3869,N_1122);
nor U8477 (N_8477,N_2866,N_2170);
xnor U8478 (N_8478,N_235,N_1669);
and U8479 (N_8479,N_3797,N_4016);
and U8480 (N_8480,N_2785,N_2810);
and U8481 (N_8481,N_4231,N_1125);
or U8482 (N_8482,N_431,N_2795);
nor U8483 (N_8483,N_3375,N_1508);
nand U8484 (N_8484,N_2264,N_2739);
nand U8485 (N_8485,N_4492,N_3668);
nand U8486 (N_8486,N_2975,N_3047);
and U8487 (N_8487,N_3628,N_2776);
and U8488 (N_8488,N_4701,N_2431);
or U8489 (N_8489,N_1372,N_115);
or U8490 (N_8490,N_1038,N_1131);
nor U8491 (N_8491,N_1297,N_1651);
xor U8492 (N_8492,N_2899,N_2857);
or U8493 (N_8493,N_4900,N_884);
or U8494 (N_8494,N_1992,N_2199);
nor U8495 (N_8495,N_3223,N_890);
nand U8496 (N_8496,N_554,N_2924);
or U8497 (N_8497,N_3009,N_2594);
nor U8498 (N_8498,N_2952,N_983);
nand U8499 (N_8499,N_4125,N_1790);
and U8500 (N_8500,N_1600,N_2156);
nand U8501 (N_8501,N_1095,N_2795);
or U8502 (N_8502,N_1120,N_927);
or U8503 (N_8503,N_2610,N_3203);
and U8504 (N_8504,N_3163,N_1570);
or U8505 (N_8505,N_2558,N_3364);
nand U8506 (N_8506,N_1694,N_1573);
or U8507 (N_8507,N_2120,N_4487);
nor U8508 (N_8508,N_1745,N_4004);
nand U8509 (N_8509,N_3430,N_4243);
or U8510 (N_8510,N_1284,N_1809);
or U8511 (N_8511,N_2272,N_4213);
and U8512 (N_8512,N_3244,N_1647);
and U8513 (N_8513,N_3877,N_1382);
nand U8514 (N_8514,N_125,N_1678);
nor U8515 (N_8515,N_2654,N_3765);
nand U8516 (N_8516,N_4989,N_2941);
nand U8517 (N_8517,N_286,N_1370);
nor U8518 (N_8518,N_1826,N_799);
nor U8519 (N_8519,N_3784,N_3519);
nor U8520 (N_8520,N_4908,N_4999);
nand U8521 (N_8521,N_1700,N_2883);
xor U8522 (N_8522,N_3894,N_3223);
nor U8523 (N_8523,N_583,N_3896);
xnor U8524 (N_8524,N_64,N_4494);
or U8525 (N_8525,N_507,N_2040);
nand U8526 (N_8526,N_1013,N_3693);
nor U8527 (N_8527,N_4963,N_149);
nand U8528 (N_8528,N_4924,N_2271);
nor U8529 (N_8529,N_3074,N_2513);
and U8530 (N_8530,N_4425,N_3024);
or U8531 (N_8531,N_3393,N_3095);
and U8532 (N_8532,N_360,N_2313);
or U8533 (N_8533,N_229,N_587);
or U8534 (N_8534,N_426,N_4140);
nor U8535 (N_8535,N_298,N_3724);
nor U8536 (N_8536,N_786,N_1045);
nand U8537 (N_8537,N_1192,N_3371);
nor U8538 (N_8538,N_594,N_1299);
nand U8539 (N_8539,N_2022,N_4380);
nor U8540 (N_8540,N_3795,N_1386);
nor U8541 (N_8541,N_2309,N_647);
nor U8542 (N_8542,N_1089,N_180);
nand U8543 (N_8543,N_1459,N_1569);
nor U8544 (N_8544,N_1624,N_1672);
or U8545 (N_8545,N_1890,N_2772);
nand U8546 (N_8546,N_317,N_261);
nand U8547 (N_8547,N_1705,N_1055);
and U8548 (N_8548,N_2835,N_184);
or U8549 (N_8549,N_3047,N_272);
or U8550 (N_8550,N_3321,N_4643);
nor U8551 (N_8551,N_4206,N_4697);
nand U8552 (N_8552,N_321,N_573);
or U8553 (N_8553,N_1599,N_1874);
nor U8554 (N_8554,N_1092,N_4267);
or U8555 (N_8555,N_2714,N_967);
and U8556 (N_8556,N_747,N_1938);
nand U8557 (N_8557,N_1751,N_449);
nand U8558 (N_8558,N_3823,N_4981);
and U8559 (N_8559,N_475,N_942);
or U8560 (N_8560,N_239,N_2079);
nor U8561 (N_8561,N_3655,N_3118);
nand U8562 (N_8562,N_1683,N_1949);
xor U8563 (N_8563,N_1282,N_4605);
or U8564 (N_8564,N_2649,N_456);
nand U8565 (N_8565,N_1703,N_1639);
nor U8566 (N_8566,N_55,N_3518);
or U8567 (N_8567,N_737,N_2241);
nor U8568 (N_8568,N_1500,N_165);
or U8569 (N_8569,N_1843,N_3431);
and U8570 (N_8570,N_1928,N_2484);
xor U8571 (N_8571,N_1378,N_1439);
or U8572 (N_8572,N_4333,N_131);
nor U8573 (N_8573,N_4400,N_3537);
nand U8574 (N_8574,N_4750,N_3770);
nand U8575 (N_8575,N_2711,N_4417);
nor U8576 (N_8576,N_4994,N_4190);
and U8577 (N_8577,N_2349,N_3120);
xor U8578 (N_8578,N_907,N_4933);
nor U8579 (N_8579,N_3940,N_1024);
and U8580 (N_8580,N_1206,N_3586);
nand U8581 (N_8581,N_1332,N_4216);
nor U8582 (N_8582,N_3081,N_4005);
and U8583 (N_8583,N_1842,N_2632);
nor U8584 (N_8584,N_3,N_2373);
xnor U8585 (N_8585,N_1836,N_2719);
xor U8586 (N_8586,N_332,N_1365);
or U8587 (N_8587,N_4427,N_1888);
nand U8588 (N_8588,N_3573,N_3821);
nand U8589 (N_8589,N_983,N_266);
xnor U8590 (N_8590,N_4960,N_1239);
nand U8591 (N_8591,N_2947,N_2005);
or U8592 (N_8592,N_3526,N_4354);
or U8593 (N_8593,N_4938,N_2259);
nor U8594 (N_8594,N_1129,N_2606);
nand U8595 (N_8595,N_1483,N_3089);
and U8596 (N_8596,N_3775,N_930);
nor U8597 (N_8597,N_1985,N_4155);
nand U8598 (N_8598,N_14,N_3123);
or U8599 (N_8599,N_2809,N_3410);
nor U8600 (N_8600,N_1732,N_87);
nand U8601 (N_8601,N_2740,N_799);
or U8602 (N_8602,N_4696,N_1180);
and U8603 (N_8603,N_4916,N_2712);
and U8604 (N_8604,N_1620,N_2026);
and U8605 (N_8605,N_167,N_415);
nand U8606 (N_8606,N_2146,N_53);
and U8607 (N_8607,N_3632,N_2966);
nor U8608 (N_8608,N_3992,N_3615);
or U8609 (N_8609,N_339,N_1816);
and U8610 (N_8610,N_4449,N_3632);
nand U8611 (N_8611,N_4475,N_588);
xor U8612 (N_8612,N_4918,N_2970);
and U8613 (N_8613,N_4242,N_4812);
nand U8614 (N_8614,N_481,N_211);
nand U8615 (N_8615,N_4442,N_1810);
nor U8616 (N_8616,N_841,N_3325);
nand U8617 (N_8617,N_1655,N_4191);
and U8618 (N_8618,N_3588,N_3026);
xnor U8619 (N_8619,N_2718,N_858);
and U8620 (N_8620,N_2626,N_2927);
nand U8621 (N_8621,N_713,N_4917);
and U8622 (N_8622,N_1190,N_3292);
or U8623 (N_8623,N_1567,N_1744);
or U8624 (N_8624,N_3379,N_640);
nand U8625 (N_8625,N_3567,N_1375);
nor U8626 (N_8626,N_292,N_2172);
nor U8627 (N_8627,N_2771,N_631);
or U8628 (N_8628,N_1943,N_2223);
nand U8629 (N_8629,N_3064,N_2687);
and U8630 (N_8630,N_3975,N_3161);
or U8631 (N_8631,N_656,N_4502);
nand U8632 (N_8632,N_3010,N_3394);
nand U8633 (N_8633,N_2232,N_4190);
nand U8634 (N_8634,N_3437,N_2022);
xor U8635 (N_8635,N_2232,N_357);
or U8636 (N_8636,N_3852,N_3754);
and U8637 (N_8637,N_4823,N_2141);
and U8638 (N_8638,N_4065,N_2136);
nand U8639 (N_8639,N_459,N_4634);
or U8640 (N_8640,N_4583,N_1628);
or U8641 (N_8641,N_4584,N_2134);
nor U8642 (N_8642,N_2094,N_2316);
or U8643 (N_8643,N_3680,N_1049);
and U8644 (N_8644,N_2323,N_565);
nand U8645 (N_8645,N_3177,N_1110);
nor U8646 (N_8646,N_982,N_4064);
or U8647 (N_8647,N_579,N_2888);
nand U8648 (N_8648,N_1169,N_3881);
nand U8649 (N_8649,N_4834,N_4906);
or U8650 (N_8650,N_4381,N_4440);
and U8651 (N_8651,N_1514,N_4023);
or U8652 (N_8652,N_176,N_2386);
nand U8653 (N_8653,N_4581,N_4192);
or U8654 (N_8654,N_2693,N_1316);
and U8655 (N_8655,N_1283,N_310);
or U8656 (N_8656,N_3077,N_4224);
nand U8657 (N_8657,N_3667,N_4054);
or U8658 (N_8658,N_2536,N_1687);
and U8659 (N_8659,N_1627,N_2237);
nand U8660 (N_8660,N_3939,N_204);
and U8661 (N_8661,N_3834,N_2244);
nand U8662 (N_8662,N_3281,N_1903);
nor U8663 (N_8663,N_4341,N_2889);
nand U8664 (N_8664,N_1262,N_2882);
xor U8665 (N_8665,N_4152,N_4647);
nand U8666 (N_8666,N_2417,N_3555);
nand U8667 (N_8667,N_2331,N_1640);
xor U8668 (N_8668,N_3280,N_3825);
and U8669 (N_8669,N_3732,N_592);
nand U8670 (N_8670,N_1141,N_3027);
and U8671 (N_8671,N_4002,N_1272);
nand U8672 (N_8672,N_1442,N_4409);
nor U8673 (N_8673,N_1129,N_4402);
nand U8674 (N_8674,N_3037,N_3548);
xor U8675 (N_8675,N_4902,N_3188);
nor U8676 (N_8676,N_2544,N_4464);
nand U8677 (N_8677,N_1194,N_2875);
or U8678 (N_8678,N_1455,N_1053);
and U8679 (N_8679,N_3152,N_1403);
nor U8680 (N_8680,N_3834,N_3015);
or U8681 (N_8681,N_3434,N_2606);
nor U8682 (N_8682,N_4302,N_960);
nor U8683 (N_8683,N_4993,N_222);
and U8684 (N_8684,N_1667,N_4046);
or U8685 (N_8685,N_13,N_2174);
or U8686 (N_8686,N_2920,N_3434);
nor U8687 (N_8687,N_49,N_2263);
nor U8688 (N_8688,N_1535,N_3949);
or U8689 (N_8689,N_2231,N_286);
xnor U8690 (N_8690,N_2753,N_2473);
and U8691 (N_8691,N_252,N_3686);
or U8692 (N_8692,N_313,N_3093);
and U8693 (N_8693,N_3883,N_483);
or U8694 (N_8694,N_7,N_1965);
nand U8695 (N_8695,N_0,N_3837);
nand U8696 (N_8696,N_4447,N_3718);
and U8697 (N_8697,N_2305,N_2198);
nand U8698 (N_8698,N_933,N_342);
xnor U8699 (N_8699,N_4155,N_1967);
or U8700 (N_8700,N_3391,N_574);
or U8701 (N_8701,N_3408,N_3897);
nand U8702 (N_8702,N_2271,N_2708);
nor U8703 (N_8703,N_3317,N_2105);
or U8704 (N_8704,N_2534,N_4922);
nor U8705 (N_8705,N_4291,N_4725);
or U8706 (N_8706,N_3227,N_2905);
nand U8707 (N_8707,N_502,N_241);
or U8708 (N_8708,N_867,N_3448);
nand U8709 (N_8709,N_644,N_3480);
or U8710 (N_8710,N_3076,N_4562);
nor U8711 (N_8711,N_1051,N_4181);
nor U8712 (N_8712,N_2550,N_1768);
nor U8713 (N_8713,N_355,N_1235);
nor U8714 (N_8714,N_1758,N_3936);
and U8715 (N_8715,N_244,N_3975);
nand U8716 (N_8716,N_306,N_4774);
or U8717 (N_8717,N_1062,N_2877);
and U8718 (N_8718,N_4608,N_4620);
nand U8719 (N_8719,N_2354,N_2088);
nand U8720 (N_8720,N_2053,N_508);
nor U8721 (N_8721,N_4493,N_3993);
nor U8722 (N_8722,N_1987,N_702);
nor U8723 (N_8723,N_2892,N_3603);
nand U8724 (N_8724,N_3844,N_345);
or U8725 (N_8725,N_4778,N_213);
and U8726 (N_8726,N_3762,N_2490);
or U8727 (N_8727,N_625,N_4274);
nor U8728 (N_8728,N_1371,N_4602);
xor U8729 (N_8729,N_1457,N_2316);
nand U8730 (N_8730,N_4330,N_609);
nand U8731 (N_8731,N_2375,N_671);
nand U8732 (N_8732,N_2007,N_840);
and U8733 (N_8733,N_1342,N_737);
or U8734 (N_8734,N_1211,N_2745);
xnor U8735 (N_8735,N_3506,N_4969);
nor U8736 (N_8736,N_2565,N_2446);
or U8737 (N_8737,N_1870,N_3122);
or U8738 (N_8738,N_1177,N_88);
and U8739 (N_8739,N_811,N_2138);
and U8740 (N_8740,N_4900,N_3535);
or U8741 (N_8741,N_430,N_1012);
or U8742 (N_8742,N_4673,N_2028);
nor U8743 (N_8743,N_1469,N_3692);
nor U8744 (N_8744,N_1031,N_4680);
nor U8745 (N_8745,N_4133,N_1880);
nand U8746 (N_8746,N_638,N_4745);
nand U8747 (N_8747,N_559,N_1244);
nand U8748 (N_8748,N_2859,N_3579);
or U8749 (N_8749,N_3078,N_966);
nand U8750 (N_8750,N_1698,N_191);
or U8751 (N_8751,N_3133,N_92);
xor U8752 (N_8752,N_3609,N_3529);
xnor U8753 (N_8753,N_3242,N_4619);
nand U8754 (N_8754,N_767,N_2551);
or U8755 (N_8755,N_3789,N_2444);
or U8756 (N_8756,N_1742,N_41);
or U8757 (N_8757,N_891,N_4266);
nor U8758 (N_8758,N_541,N_4248);
or U8759 (N_8759,N_3468,N_1002);
and U8760 (N_8760,N_2452,N_2461);
nand U8761 (N_8761,N_1528,N_1106);
nor U8762 (N_8762,N_1896,N_1102);
nand U8763 (N_8763,N_917,N_1294);
xnor U8764 (N_8764,N_4522,N_3652);
and U8765 (N_8765,N_3550,N_614);
nand U8766 (N_8766,N_419,N_3261);
or U8767 (N_8767,N_2291,N_3276);
or U8768 (N_8768,N_4373,N_663);
xor U8769 (N_8769,N_1644,N_1933);
nand U8770 (N_8770,N_1014,N_4655);
nand U8771 (N_8771,N_1099,N_2181);
and U8772 (N_8772,N_2846,N_4210);
nand U8773 (N_8773,N_4076,N_2595);
or U8774 (N_8774,N_4888,N_457);
nor U8775 (N_8775,N_446,N_3486);
nor U8776 (N_8776,N_4180,N_431);
and U8777 (N_8777,N_4437,N_1182);
nand U8778 (N_8778,N_482,N_271);
and U8779 (N_8779,N_1146,N_1432);
and U8780 (N_8780,N_1888,N_484);
xor U8781 (N_8781,N_209,N_3015);
nor U8782 (N_8782,N_2896,N_4036);
nand U8783 (N_8783,N_3261,N_2968);
or U8784 (N_8784,N_185,N_4086);
and U8785 (N_8785,N_2209,N_3644);
nor U8786 (N_8786,N_3517,N_4073);
nand U8787 (N_8787,N_391,N_724);
nor U8788 (N_8788,N_4179,N_2068);
and U8789 (N_8789,N_720,N_2033);
or U8790 (N_8790,N_4592,N_2299);
nand U8791 (N_8791,N_1738,N_4379);
and U8792 (N_8792,N_1842,N_4579);
nor U8793 (N_8793,N_1190,N_3669);
and U8794 (N_8794,N_2429,N_2072);
or U8795 (N_8795,N_28,N_3187);
xor U8796 (N_8796,N_631,N_1487);
or U8797 (N_8797,N_905,N_4192);
nor U8798 (N_8798,N_2387,N_3273);
or U8799 (N_8799,N_4889,N_1335);
and U8800 (N_8800,N_4873,N_4933);
or U8801 (N_8801,N_695,N_4442);
nor U8802 (N_8802,N_2788,N_3288);
and U8803 (N_8803,N_3989,N_2288);
nand U8804 (N_8804,N_4501,N_4439);
or U8805 (N_8805,N_2287,N_1947);
or U8806 (N_8806,N_3608,N_4259);
and U8807 (N_8807,N_4570,N_1174);
nor U8808 (N_8808,N_4467,N_4027);
and U8809 (N_8809,N_1433,N_360);
or U8810 (N_8810,N_2009,N_2007);
and U8811 (N_8811,N_3054,N_3684);
nand U8812 (N_8812,N_4213,N_1124);
nor U8813 (N_8813,N_3571,N_2300);
nor U8814 (N_8814,N_2273,N_3088);
and U8815 (N_8815,N_2565,N_3448);
and U8816 (N_8816,N_186,N_2007);
nand U8817 (N_8817,N_4109,N_1127);
and U8818 (N_8818,N_2991,N_2314);
xnor U8819 (N_8819,N_4657,N_2177);
nor U8820 (N_8820,N_464,N_4031);
and U8821 (N_8821,N_3848,N_3809);
nand U8822 (N_8822,N_3933,N_1942);
or U8823 (N_8823,N_490,N_4317);
or U8824 (N_8824,N_3629,N_2424);
and U8825 (N_8825,N_3740,N_4680);
or U8826 (N_8826,N_1834,N_2859);
nand U8827 (N_8827,N_1615,N_4969);
nand U8828 (N_8828,N_901,N_3736);
or U8829 (N_8829,N_3983,N_2218);
and U8830 (N_8830,N_1126,N_4419);
nand U8831 (N_8831,N_2280,N_3759);
or U8832 (N_8832,N_416,N_2417);
xor U8833 (N_8833,N_1523,N_1024);
and U8834 (N_8834,N_3797,N_3022);
or U8835 (N_8835,N_1975,N_2948);
nor U8836 (N_8836,N_2799,N_3963);
xnor U8837 (N_8837,N_4010,N_4059);
or U8838 (N_8838,N_4197,N_1044);
nand U8839 (N_8839,N_4987,N_2700);
nor U8840 (N_8840,N_298,N_2069);
and U8841 (N_8841,N_4377,N_1527);
nor U8842 (N_8842,N_375,N_1178);
or U8843 (N_8843,N_4130,N_1103);
or U8844 (N_8844,N_1620,N_2085);
and U8845 (N_8845,N_3475,N_3774);
or U8846 (N_8846,N_1484,N_4650);
and U8847 (N_8847,N_1198,N_1404);
or U8848 (N_8848,N_137,N_3741);
and U8849 (N_8849,N_3739,N_2633);
nand U8850 (N_8850,N_1254,N_2668);
or U8851 (N_8851,N_1049,N_166);
nand U8852 (N_8852,N_2470,N_3601);
or U8853 (N_8853,N_3033,N_4197);
nand U8854 (N_8854,N_2731,N_3424);
nor U8855 (N_8855,N_2756,N_1396);
nor U8856 (N_8856,N_4853,N_2989);
nand U8857 (N_8857,N_4175,N_4702);
and U8858 (N_8858,N_3532,N_2041);
nor U8859 (N_8859,N_1030,N_3144);
nor U8860 (N_8860,N_2043,N_2633);
or U8861 (N_8861,N_4881,N_3659);
nand U8862 (N_8862,N_3027,N_4330);
nand U8863 (N_8863,N_2625,N_262);
nand U8864 (N_8864,N_1358,N_697);
or U8865 (N_8865,N_428,N_91);
or U8866 (N_8866,N_3561,N_1039);
and U8867 (N_8867,N_861,N_720);
nand U8868 (N_8868,N_4609,N_4675);
or U8869 (N_8869,N_1579,N_1379);
or U8870 (N_8870,N_2072,N_753);
nor U8871 (N_8871,N_1462,N_2145);
nand U8872 (N_8872,N_546,N_1390);
nand U8873 (N_8873,N_4398,N_1827);
xor U8874 (N_8874,N_993,N_443);
nor U8875 (N_8875,N_728,N_2834);
xor U8876 (N_8876,N_3381,N_691);
or U8877 (N_8877,N_3896,N_3772);
nand U8878 (N_8878,N_4936,N_4786);
or U8879 (N_8879,N_3514,N_2974);
nand U8880 (N_8880,N_3908,N_2490);
xnor U8881 (N_8881,N_813,N_1542);
nor U8882 (N_8882,N_2390,N_4988);
xnor U8883 (N_8883,N_4976,N_3087);
nand U8884 (N_8884,N_3784,N_677);
nand U8885 (N_8885,N_3331,N_2979);
or U8886 (N_8886,N_267,N_559);
xor U8887 (N_8887,N_1209,N_1358);
or U8888 (N_8888,N_1112,N_489);
or U8889 (N_8889,N_4554,N_9);
xor U8890 (N_8890,N_4882,N_2073);
and U8891 (N_8891,N_2487,N_2513);
xor U8892 (N_8892,N_3595,N_1525);
xnor U8893 (N_8893,N_185,N_3217);
xor U8894 (N_8894,N_3263,N_4792);
nand U8895 (N_8895,N_1467,N_457);
or U8896 (N_8896,N_4673,N_4983);
nor U8897 (N_8897,N_1705,N_4745);
and U8898 (N_8898,N_293,N_973);
nand U8899 (N_8899,N_3490,N_2494);
and U8900 (N_8900,N_4514,N_4730);
or U8901 (N_8901,N_1337,N_3331);
nor U8902 (N_8902,N_2368,N_4722);
nor U8903 (N_8903,N_3758,N_2714);
nor U8904 (N_8904,N_1017,N_4725);
nor U8905 (N_8905,N_4975,N_2655);
or U8906 (N_8906,N_4687,N_1678);
nor U8907 (N_8907,N_3296,N_3763);
and U8908 (N_8908,N_2054,N_4357);
or U8909 (N_8909,N_4832,N_580);
or U8910 (N_8910,N_4158,N_749);
or U8911 (N_8911,N_3202,N_507);
and U8912 (N_8912,N_2821,N_2246);
or U8913 (N_8913,N_3228,N_984);
and U8914 (N_8914,N_4484,N_798);
or U8915 (N_8915,N_4265,N_453);
and U8916 (N_8916,N_3956,N_1630);
or U8917 (N_8917,N_4481,N_4387);
xor U8918 (N_8918,N_2135,N_3001);
nor U8919 (N_8919,N_2159,N_3685);
nor U8920 (N_8920,N_826,N_1814);
nor U8921 (N_8921,N_2864,N_4587);
nand U8922 (N_8922,N_3512,N_3265);
and U8923 (N_8923,N_4796,N_4774);
or U8924 (N_8924,N_3574,N_1058);
nand U8925 (N_8925,N_3388,N_3866);
nand U8926 (N_8926,N_61,N_349);
and U8927 (N_8927,N_209,N_4246);
nand U8928 (N_8928,N_2922,N_4101);
nor U8929 (N_8929,N_1015,N_4768);
or U8930 (N_8930,N_2188,N_4257);
nor U8931 (N_8931,N_4496,N_4106);
nand U8932 (N_8932,N_903,N_598);
and U8933 (N_8933,N_1591,N_414);
nand U8934 (N_8934,N_23,N_1852);
xnor U8935 (N_8935,N_456,N_2394);
nand U8936 (N_8936,N_4662,N_562);
nand U8937 (N_8937,N_1525,N_3562);
nand U8938 (N_8938,N_1045,N_3045);
nand U8939 (N_8939,N_3910,N_4802);
xnor U8940 (N_8940,N_808,N_286);
or U8941 (N_8941,N_204,N_1513);
xnor U8942 (N_8942,N_4283,N_1633);
nand U8943 (N_8943,N_1530,N_2987);
nor U8944 (N_8944,N_2909,N_2829);
nor U8945 (N_8945,N_1671,N_2229);
nand U8946 (N_8946,N_3974,N_324);
nor U8947 (N_8947,N_4844,N_1306);
nand U8948 (N_8948,N_3080,N_2008);
nor U8949 (N_8949,N_3509,N_2794);
or U8950 (N_8950,N_2585,N_1734);
and U8951 (N_8951,N_618,N_2087);
and U8952 (N_8952,N_4654,N_4726);
nor U8953 (N_8953,N_1619,N_3799);
nand U8954 (N_8954,N_4471,N_598);
and U8955 (N_8955,N_2646,N_1488);
nor U8956 (N_8956,N_2888,N_1141);
nand U8957 (N_8957,N_2366,N_4059);
nor U8958 (N_8958,N_2889,N_845);
or U8959 (N_8959,N_3276,N_2529);
or U8960 (N_8960,N_3736,N_3190);
xnor U8961 (N_8961,N_457,N_968);
nand U8962 (N_8962,N_1791,N_1828);
xnor U8963 (N_8963,N_540,N_4219);
xnor U8964 (N_8964,N_730,N_1168);
nor U8965 (N_8965,N_1633,N_4139);
nand U8966 (N_8966,N_2437,N_1497);
or U8967 (N_8967,N_3450,N_2201);
xnor U8968 (N_8968,N_3092,N_1437);
nand U8969 (N_8969,N_156,N_3560);
or U8970 (N_8970,N_1221,N_4535);
nand U8971 (N_8971,N_859,N_2311);
and U8972 (N_8972,N_3779,N_4807);
nor U8973 (N_8973,N_1982,N_386);
and U8974 (N_8974,N_1144,N_2007);
and U8975 (N_8975,N_756,N_2998);
and U8976 (N_8976,N_3058,N_1262);
xor U8977 (N_8977,N_2489,N_1166);
nor U8978 (N_8978,N_250,N_497);
nand U8979 (N_8979,N_2799,N_3920);
nand U8980 (N_8980,N_1851,N_2958);
and U8981 (N_8981,N_3366,N_1740);
nor U8982 (N_8982,N_497,N_1406);
and U8983 (N_8983,N_3691,N_2387);
nand U8984 (N_8984,N_4915,N_125);
nand U8985 (N_8985,N_3614,N_652);
nand U8986 (N_8986,N_32,N_4785);
nand U8987 (N_8987,N_488,N_526);
and U8988 (N_8988,N_1795,N_3377);
nor U8989 (N_8989,N_4157,N_4903);
and U8990 (N_8990,N_2285,N_3411);
or U8991 (N_8991,N_1929,N_4962);
nand U8992 (N_8992,N_1192,N_908);
and U8993 (N_8993,N_4881,N_478);
nor U8994 (N_8994,N_472,N_2508);
or U8995 (N_8995,N_168,N_4107);
and U8996 (N_8996,N_3911,N_1381);
nand U8997 (N_8997,N_3593,N_3775);
nor U8998 (N_8998,N_460,N_1568);
or U8999 (N_8999,N_1605,N_2812);
or U9000 (N_9000,N_1918,N_2757);
or U9001 (N_9001,N_93,N_1375);
nor U9002 (N_9002,N_2259,N_2029);
and U9003 (N_9003,N_1917,N_187);
or U9004 (N_9004,N_2526,N_3027);
or U9005 (N_9005,N_3071,N_2574);
nand U9006 (N_9006,N_944,N_1699);
or U9007 (N_9007,N_3367,N_2618);
nor U9008 (N_9008,N_4588,N_2970);
and U9009 (N_9009,N_3024,N_4520);
nand U9010 (N_9010,N_4164,N_1526);
and U9011 (N_9011,N_4289,N_3447);
and U9012 (N_9012,N_532,N_3152);
or U9013 (N_9013,N_3924,N_4727);
or U9014 (N_9014,N_1019,N_209);
xor U9015 (N_9015,N_1984,N_3233);
nor U9016 (N_9016,N_2060,N_4142);
nand U9017 (N_9017,N_1765,N_4485);
nand U9018 (N_9018,N_3872,N_3502);
and U9019 (N_9019,N_4427,N_3982);
or U9020 (N_9020,N_1499,N_994);
and U9021 (N_9021,N_61,N_4072);
or U9022 (N_9022,N_3425,N_2553);
nand U9023 (N_9023,N_4524,N_886);
nand U9024 (N_9024,N_1377,N_1438);
nand U9025 (N_9025,N_1319,N_1867);
nand U9026 (N_9026,N_1484,N_261);
or U9027 (N_9027,N_1727,N_375);
or U9028 (N_9028,N_2164,N_1616);
nand U9029 (N_9029,N_2523,N_3397);
nand U9030 (N_9030,N_2365,N_436);
nand U9031 (N_9031,N_4544,N_583);
and U9032 (N_9032,N_3032,N_1008);
and U9033 (N_9033,N_723,N_1267);
nand U9034 (N_9034,N_3235,N_1063);
or U9035 (N_9035,N_509,N_3839);
and U9036 (N_9036,N_723,N_4581);
nor U9037 (N_9037,N_2863,N_3964);
nor U9038 (N_9038,N_24,N_2415);
nor U9039 (N_9039,N_2882,N_1513);
nand U9040 (N_9040,N_2303,N_1255);
or U9041 (N_9041,N_335,N_4991);
nand U9042 (N_9042,N_1078,N_2177);
and U9043 (N_9043,N_2882,N_1588);
and U9044 (N_9044,N_259,N_1916);
nand U9045 (N_9045,N_2270,N_1401);
and U9046 (N_9046,N_1302,N_816);
nand U9047 (N_9047,N_980,N_1485);
and U9048 (N_9048,N_2245,N_2590);
nor U9049 (N_9049,N_439,N_3583);
nor U9050 (N_9050,N_3481,N_402);
or U9051 (N_9051,N_1511,N_4603);
nor U9052 (N_9052,N_3688,N_1402);
and U9053 (N_9053,N_1012,N_757);
nor U9054 (N_9054,N_794,N_34);
xor U9055 (N_9055,N_3232,N_4460);
nor U9056 (N_9056,N_2091,N_4862);
nor U9057 (N_9057,N_562,N_2477);
or U9058 (N_9058,N_4171,N_1572);
nor U9059 (N_9059,N_341,N_2484);
nor U9060 (N_9060,N_1677,N_4520);
xnor U9061 (N_9061,N_4273,N_2155);
nor U9062 (N_9062,N_1749,N_1896);
xnor U9063 (N_9063,N_924,N_1659);
nand U9064 (N_9064,N_4287,N_4035);
nor U9065 (N_9065,N_974,N_4924);
nand U9066 (N_9066,N_1904,N_1500);
nand U9067 (N_9067,N_3599,N_932);
and U9068 (N_9068,N_2308,N_64);
nand U9069 (N_9069,N_4992,N_1919);
nor U9070 (N_9070,N_4758,N_2479);
and U9071 (N_9071,N_3483,N_730);
xnor U9072 (N_9072,N_1670,N_2145);
and U9073 (N_9073,N_658,N_463);
or U9074 (N_9074,N_4412,N_2532);
nand U9075 (N_9075,N_439,N_2671);
and U9076 (N_9076,N_155,N_2724);
or U9077 (N_9077,N_104,N_1103);
nand U9078 (N_9078,N_4760,N_1377);
nor U9079 (N_9079,N_3284,N_18);
and U9080 (N_9080,N_280,N_858);
xnor U9081 (N_9081,N_703,N_2945);
nor U9082 (N_9082,N_4737,N_834);
xor U9083 (N_9083,N_251,N_2288);
and U9084 (N_9084,N_1728,N_1190);
nor U9085 (N_9085,N_3537,N_1821);
nand U9086 (N_9086,N_4571,N_4903);
nand U9087 (N_9087,N_4770,N_3996);
nor U9088 (N_9088,N_4126,N_4434);
nand U9089 (N_9089,N_2477,N_69);
nand U9090 (N_9090,N_2384,N_3717);
nor U9091 (N_9091,N_1534,N_3761);
nand U9092 (N_9092,N_3363,N_1401);
nand U9093 (N_9093,N_2520,N_4294);
xnor U9094 (N_9094,N_4587,N_2538);
xnor U9095 (N_9095,N_1082,N_2847);
or U9096 (N_9096,N_2708,N_2594);
nor U9097 (N_9097,N_2363,N_4560);
nor U9098 (N_9098,N_1978,N_1456);
and U9099 (N_9099,N_188,N_3775);
and U9100 (N_9100,N_2968,N_1616);
nand U9101 (N_9101,N_1632,N_4683);
nand U9102 (N_9102,N_2932,N_901);
nor U9103 (N_9103,N_1469,N_2457);
nor U9104 (N_9104,N_1309,N_3931);
and U9105 (N_9105,N_1674,N_3151);
xor U9106 (N_9106,N_1540,N_4033);
nor U9107 (N_9107,N_3432,N_3100);
or U9108 (N_9108,N_2188,N_1870);
and U9109 (N_9109,N_1483,N_4375);
xnor U9110 (N_9110,N_2362,N_3099);
xnor U9111 (N_9111,N_671,N_652);
or U9112 (N_9112,N_3947,N_1695);
xnor U9113 (N_9113,N_4448,N_1056);
nand U9114 (N_9114,N_4908,N_1557);
or U9115 (N_9115,N_2739,N_3894);
or U9116 (N_9116,N_2810,N_1656);
nand U9117 (N_9117,N_1721,N_595);
nand U9118 (N_9118,N_3988,N_2446);
or U9119 (N_9119,N_1736,N_664);
or U9120 (N_9120,N_795,N_4189);
nand U9121 (N_9121,N_2350,N_1912);
and U9122 (N_9122,N_748,N_3718);
or U9123 (N_9123,N_2495,N_2249);
or U9124 (N_9124,N_2701,N_4927);
nand U9125 (N_9125,N_298,N_430);
xor U9126 (N_9126,N_201,N_3562);
and U9127 (N_9127,N_4055,N_1378);
nor U9128 (N_9128,N_2197,N_1044);
nand U9129 (N_9129,N_4863,N_1940);
xor U9130 (N_9130,N_3145,N_4644);
or U9131 (N_9131,N_2700,N_1335);
nand U9132 (N_9132,N_1668,N_2793);
nor U9133 (N_9133,N_3660,N_2538);
and U9134 (N_9134,N_916,N_4228);
xnor U9135 (N_9135,N_2744,N_1197);
and U9136 (N_9136,N_2881,N_2204);
nand U9137 (N_9137,N_65,N_4050);
nor U9138 (N_9138,N_4743,N_1264);
nor U9139 (N_9139,N_1712,N_2460);
nand U9140 (N_9140,N_2659,N_4480);
nand U9141 (N_9141,N_2683,N_1949);
nand U9142 (N_9142,N_3985,N_1307);
xnor U9143 (N_9143,N_371,N_822);
nor U9144 (N_9144,N_3717,N_1996);
and U9145 (N_9145,N_3017,N_1158);
nand U9146 (N_9146,N_945,N_1111);
nor U9147 (N_9147,N_1227,N_810);
xnor U9148 (N_9148,N_3061,N_1784);
nand U9149 (N_9149,N_1741,N_4470);
or U9150 (N_9150,N_3374,N_4262);
and U9151 (N_9151,N_3936,N_4202);
xnor U9152 (N_9152,N_1495,N_2876);
or U9153 (N_9153,N_2273,N_1221);
or U9154 (N_9154,N_654,N_700);
nor U9155 (N_9155,N_4,N_3018);
or U9156 (N_9156,N_3225,N_1287);
nand U9157 (N_9157,N_1271,N_1015);
or U9158 (N_9158,N_3803,N_4772);
xor U9159 (N_9159,N_1696,N_3392);
and U9160 (N_9160,N_4968,N_593);
or U9161 (N_9161,N_3314,N_4386);
xnor U9162 (N_9162,N_3626,N_4265);
or U9163 (N_9163,N_3054,N_4500);
nor U9164 (N_9164,N_1540,N_2225);
and U9165 (N_9165,N_1325,N_4938);
nor U9166 (N_9166,N_197,N_4408);
and U9167 (N_9167,N_2627,N_1130);
or U9168 (N_9168,N_1926,N_1871);
nand U9169 (N_9169,N_1089,N_1898);
nor U9170 (N_9170,N_4883,N_2639);
or U9171 (N_9171,N_4604,N_1235);
xor U9172 (N_9172,N_4711,N_1284);
or U9173 (N_9173,N_4658,N_4987);
and U9174 (N_9174,N_3832,N_1226);
or U9175 (N_9175,N_2096,N_4457);
xnor U9176 (N_9176,N_3863,N_2069);
or U9177 (N_9177,N_3016,N_4965);
xnor U9178 (N_9178,N_1541,N_3707);
and U9179 (N_9179,N_543,N_2211);
nor U9180 (N_9180,N_3797,N_3573);
nand U9181 (N_9181,N_2235,N_900);
and U9182 (N_9182,N_2855,N_1374);
xor U9183 (N_9183,N_2629,N_4024);
nor U9184 (N_9184,N_2610,N_2357);
and U9185 (N_9185,N_1692,N_3812);
and U9186 (N_9186,N_624,N_760);
or U9187 (N_9187,N_562,N_2848);
nor U9188 (N_9188,N_935,N_1017);
or U9189 (N_9189,N_653,N_2026);
nor U9190 (N_9190,N_709,N_1675);
and U9191 (N_9191,N_3434,N_3292);
and U9192 (N_9192,N_4553,N_3475);
and U9193 (N_9193,N_1499,N_2924);
and U9194 (N_9194,N_1324,N_3532);
or U9195 (N_9195,N_2712,N_4228);
nand U9196 (N_9196,N_2508,N_588);
nand U9197 (N_9197,N_1843,N_2182);
nor U9198 (N_9198,N_1017,N_1563);
and U9199 (N_9199,N_3530,N_674);
nand U9200 (N_9200,N_4335,N_4934);
nor U9201 (N_9201,N_2071,N_4053);
xor U9202 (N_9202,N_781,N_1689);
or U9203 (N_9203,N_2167,N_4102);
nand U9204 (N_9204,N_3742,N_1849);
nor U9205 (N_9205,N_3656,N_632);
xor U9206 (N_9206,N_3672,N_2084);
or U9207 (N_9207,N_1438,N_2135);
nor U9208 (N_9208,N_3245,N_1118);
or U9209 (N_9209,N_716,N_2466);
xnor U9210 (N_9210,N_3051,N_3981);
nand U9211 (N_9211,N_716,N_3170);
and U9212 (N_9212,N_4037,N_3618);
or U9213 (N_9213,N_1954,N_4802);
nand U9214 (N_9214,N_467,N_2385);
and U9215 (N_9215,N_3459,N_1099);
nand U9216 (N_9216,N_2704,N_2076);
or U9217 (N_9217,N_2625,N_914);
or U9218 (N_9218,N_1804,N_3768);
nor U9219 (N_9219,N_1554,N_3632);
and U9220 (N_9220,N_4215,N_1988);
nand U9221 (N_9221,N_490,N_3511);
nand U9222 (N_9222,N_1422,N_4694);
nand U9223 (N_9223,N_4662,N_2484);
nor U9224 (N_9224,N_3827,N_1226);
or U9225 (N_9225,N_726,N_4821);
nor U9226 (N_9226,N_941,N_4546);
and U9227 (N_9227,N_2681,N_3675);
and U9228 (N_9228,N_1968,N_2374);
nand U9229 (N_9229,N_4927,N_2319);
and U9230 (N_9230,N_4520,N_1445);
nand U9231 (N_9231,N_4683,N_455);
and U9232 (N_9232,N_2942,N_2631);
and U9233 (N_9233,N_1551,N_2599);
or U9234 (N_9234,N_2334,N_4408);
nor U9235 (N_9235,N_340,N_3826);
xnor U9236 (N_9236,N_408,N_1911);
nor U9237 (N_9237,N_1094,N_4688);
xnor U9238 (N_9238,N_369,N_2110);
and U9239 (N_9239,N_3307,N_4867);
nand U9240 (N_9240,N_4727,N_2557);
nor U9241 (N_9241,N_1262,N_1941);
xnor U9242 (N_9242,N_4573,N_1660);
and U9243 (N_9243,N_2351,N_3851);
and U9244 (N_9244,N_755,N_2894);
and U9245 (N_9245,N_4047,N_4987);
nor U9246 (N_9246,N_1322,N_378);
and U9247 (N_9247,N_3230,N_224);
xor U9248 (N_9248,N_8,N_3673);
xor U9249 (N_9249,N_1353,N_2346);
nor U9250 (N_9250,N_3594,N_710);
or U9251 (N_9251,N_1083,N_2315);
nand U9252 (N_9252,N_833,N_4032);
nor U9253 (N_9253,N_3849,N_542);
or U9254 (N_9254,N_1575,N_2332);
nor U9255 (N_9255,N_2806,N_726);
nor U9256 (N_9256,N_4165,N_4131);
or U9257 (N_9257,N_3410,N_2359);
nor U9258 (N_9258,N_3333,N_3536);
and U9259 (N_9259,N_758,N_1360);
nand U9260 (N_9260,N_3043,N_2720);
nor U9261 (N_9261,N_1197,N_4751);
or U9262 (N_9262,N_320,N_2286);
xnor U9263 (N_9263,N_4409,N_2802);
and U9264 (N_9264,N_4379,N_1424);
xnor U9265 (N_9265,N_1580,N_1107);
and U9266 (N_9266,N_228,N_4690);
and U9267 (N_9267,N_3903,N_4622);
and U9268 (N_9268,N_3330,N_3784);
nand U9269 (N_9269,N_4929,N_3296);
and U9270 (N_9270,N_3991,N_3167);
nand U9271 (N_9271,N_1017,N_2422);
nor U9272 (N_9272,N_1230,N_4407);
nor U9273 (N_9273,N_2162,N_1113);
xor U9274 (N_9274,N_594,N_3218);
xor U9275 (N_9275,N_1574,N_3184);
nor U9276 (N_9276,N_4194,N_3902);
or U9277 (N_9277,N_3683,N_104);
or U9278 (N_9278,N_3665,N_283);
nand U9279 (N_9279,N_1359,N_4775);
and U9280 (N_9280,N_3546,N_334);
nor U9281 (N_9281,N_2994,N_3662);
and U9282 (N_9282,N_2880,N_4440);
or U9283 (N_9283,N_406,N_1760);
or U9284 (N_9284,N_1499,N_374);
xor U9285 (N_9285,N_268,N_667);
xor U9286 (N_9286,N_3202,N_846);
nor U9287 (N_9287,N_2455,N_2742);
and U9288 (N_9288,N_4868,N_1625);
or U9289 (N_9289,N_3426,N_1854);
xnor U9290 (N_9290,N_3448,N_4870);
nand U9291 (N_9291,N_120,N_4856);
or U9292 (N_9292,N_2493,N_816);
and U9293 (N_9293,N_4261,N_3660);
and U9294 (N_9294,N_1639,N_4267);
nor U9295 (N_9295,N_4125,N_76);
xnor U9296 (N_9296,N_4157,N_3826);
and U9297 (N_9297,N_4610,N_3629);
and U9298 (N_9298,N_4518,N_3983);
and U9299 (N_9299,N_439,N_1675);
or U9300 (N_9300,N_2798,N_1182);
or U9301 (N_9301,N_3855,N_260);
nand U9302 (N_9302,N_1472,N_3036);
or U9303 (N_9303,N_1908,N_3270);
nand U9304 (N_9304,N_4874,N_833);
or U9305 (N_9305,N_1145,N_1568);
nand U9306 (N_9306,N_2819,N_500);
nor U9307 (N_9307,N_4583,N_2228);
and U9308 (N_9308,N_1993,N_2844);
or U9309 (N_9309,N_2424,N_3564);
or U9310 (N_9310,N_2212,N_303);
nor U9311 (N_9311,N_2002,N_2);
and U9312 (N_9312,N_3620,N_3775);
nor U9313 (N_9313,N_2142,N_4727);
nor U9314 (N_9314,N_2458,N_2342);
xor U9315 (N_9315,N_2582,N_976);
and U9316 (N_9316,N_1383,N_4325);
nand U9317 (N_9317,N_4903,N_396);
or U9318 (N_9318,N_2005,N_926);
or U9319 (N_9319,N_246,N_1255);
nor U9320 (N_9320,N_2583,N_1822);
nand U9321 (N_9321,N_3366,N_3610);
nand U9322 (N_9322,N_2837,N_581);
or U9323 (N_9323,N_141,N_3154);
and U9324 (N_9324,N_4287,N_2421);
nand U9325 (N_9325,N_3058,N_4261);
nor U9326 (N_9326,N_3435,N_3036);
nand U9327 (N_9327,N_161,N_703);
nor U9328 (N_9328,N_583,N_2590);
and U9329 (N_9329,N_1592,N_1613);
or U9330 (N_9330,N_4817,N_2620);
or U9331 (N_9331,N_2108,N_2650);
xnor U9332 (N_9332,N_4532,N_561);
xnor U9333 (N_9333,N_3740,N_3090);
and U9334 (N_9334,N_1057,N_1657);
or U9335 (N_9335,N_2818,N_3021);
and U9336 (N_9336,N_1206,N_974);
xor U9337 (N_9337,N_1810,N_484);
or U9338 (N_9338,N_3940,N_1812);
nand U9339 (N_9339,N_2323,N_761);
nand U9340 (N_9340,N_2053,N_4629);
and U9341 (N_9341,N_3809,N_3534);
nor U9342 (N_9342,N_1562,N_4333);
nor U9343 (N_9343,N_3144,N_4590);
and U9344 (N_9344,N_4408,N_3560);
nor U9345 (N_9345,N_1502,N_4929);
xor U9346 (N_9346,N_1547,N_663);
and U9347 (N_9347,N_1741,N_605);
nand U9348 (N_9348,N_778,N_2015);
or U9349 (N_9349,N_4553,N_3412);
and U9350 (N_9350,N_910,N_4253);
or U9351 (N_9351,N_344,N_2974);
and U9352 (N_9352,N_4715,N_1454);
nor U9353 (N_9353,N_1165,N_525);
or U9354 (N_9354,N_328,N_3065);
nand U9355 (N_9355,N_2482,N_3001);
or U9356 (N_9356,N_1693,N_4087);
and U9357 (N_9357,N_296,N_4720);
nor U9358 (N_9358,N_3966,N_3790);
and U9359 (N_9359,N_4967,N_1230);
and U9360 (N_9360,N_2969,N_1754);
or U9361 (N_9361,N_899,N_616);
or U9362 (N_9362,N_812,N_1684);
nand U9363 (N_9363,N_3265,N_3565);
and U9364 (N_9364,N_1639,N_3235);
or U9365 (N_9365,N_1807,N_1036);
xnor U9366 (N_9366,N_1827,N_3011);
and U9367 (N_9367,N_1164,N_2640);
and U9368 (N_9368,N_2094,N_526);
and U9369 (N_9369,N_1750,N_1756);
and U9370 (N_9370,N_4916,N_1174);
nor U9371 (N_9371,N_1706,N_489);
nand U9372 (N_9372,N_4874,N_2385);
or U9373 (N_9373,N_783,N_89);
or U9374 (N_9374,N_437,N_1046);
or U9375 (N_9375,N_3354,N_2608);
nand U9376 (N_9376,N_1930,N_2496);
and U9377 (N_9377,N_1409,N_107);
or U9378 (N_9378,N_4209,N_1716);
and U9379 (N_9379,N_4194,N_1499);
and U9380 (N_9380,N_4989,N_3058);
and U9381 (N_9381,N_295,N_3470);
or U9382 (N_9382,N_3282,N_1568);
or U9383 (N_9383,N_2091,N_458);
nand U9384 (N_9384,N_508,N_1112);
nand U9385 (N_9385,N_3692,N_4603);
and U9386 (N_9386,N_4928,N_1871);
and U9387 (N_9387,N_4264,N_2386);
and U9388 (N_9388,N_1191,N_2253);
xor U9389 (N_9389,N_815,N_1349);
or U9390 (N_9390,N_16,N_335);
nor U9391 (N_9391,N_4452,N_3171);
nand U9392 (N_9392,N_4816,N_3034);
nand U9393 (N_9393,N_685,N_4470);
and U9394 (N_9394,N_4010,N_4661);
xnor U9395 (N_9395,N_1966,N_3283);
nand U9396 (N_9396,N_1580,N_1711);
and U9397 (N_9397,N_426,N_2482);
nor U9398 (N_9398,N_4834,N_1523);
nor U9399 (N_9399,N_1151,N_3136);
or U9400 (N_9400,N_2606,N_2864);
and U9401 (N_9401,N_3892,N_779);
and U9402 (N_9402,N_4940,N_55);
nand U9403 (N_9403,N_3835,N_2297);
or U9404 (N_9404,N_869,N_3887);
or U9405 (N_9405,N_1621,N_2128);
and U9406 (N_9406,N_4248,N_4312);
xor U9407 (N_9407,N_1082,N_4921);
or U9408 (N_9408,N_3238,N_4941);
and U9409 (N_9409,N_3636,N_2896);
nor U9410 (N_9410,N_3046,N_4205);
and U9411 (N_9411,N_3419,N_268);
and U9412 (N_9412,N_295,N_2161);
nor U9413 (N_9413,N_1871,N_3440);
nand U9414 (N_9414,N_949,N_931);
and U9415 (N_9415,N_1684,N_1741);
nand U9416 (N_9416,N_1468,N_3022);
or U9417 (N_9417,N_1435,N_2423);
xnor U9418 (N_9418,N_513,N_3088);
or U9419 (N_9419,N_2894,N_4917);
and U9420 (N_9420,N_2238,N_3183);
nor U9421 (N_9421,N_1389,N_1362);
xnor U9422 (N_9422,N_1604,N_3617);
nand U9423 (N_9423,N_3574,N_1450);
nor U9424 (N_9424,N_166,N_4413);
xnor U9425 (N_9425,N_4509,N_4046);
or U9426 (N_9426,N_3691,N_598);
or U9427 (N_9427,N_1096,N_4238);
and U9428 (N_9428,N_643,N_3609);
nor U9429 (N_9429,N_4851,N_3473);
nand U9430 (N_9430,N_4932,N_618);
nor U9431 (N_9431,N_138,N_1845);
nor U9432 (N_9432,N_171,N_660);
or U9433 (N_9433,N_1720,N_1220);
nand U9434 (N_9434,N_2063,N_2157);
or U9435 (N_9435,N_2500,N_2315);
or U9436 (N_9436,N_4587,N_3350);
or U9437 (N_9437,N_1186,N_720);
or U9438 (N_9438,N_1025,N_738);
or U9439 (N_9439,N_2891,N_2615);
and U9440 (N_9440,N_1046,N_981);
and U9441 (N_9441,N_4593,N_2645);
nor U9442 (N_9442,N_1249,N_2718);
and U9443 (N_9443,N_3459,N_1193);
and U9444 (N_9444,N_1519,N_3764);
and U9445 (N_9445,N_3048,N_2893);
or U9446 (N_9446,N_2798,N_4171);
nor U9447 (N_9447,N_1329,N_2338);
nor U9448 (N_9448,N_1247,N_3719);
nor U9449 (N_9449,N_661,N_3205);
xor U9450 (N_9450,N_496,N_646);
nor U9451 (N_9451,N_3961,N_1288);
and U9452 (N_9452,N_663,N_4323);
or U9453 (N_9453,N_4128,N_4352);
nand U9454 (N_9454,N_4404,N_3616);
nor U9455 (N_9455,N_2680,N_787);
nand U9456 (N_9456,N_3863,N_3489);
nand U9457 (N_9457,N_1030,N_268);
or U9458 (N_9458,N_2174,N_4692);
xnor U9459 (N_9459,N_1531,N_811);
xnor U9460 (N_9460,N_747,N_1053);
nor U9461 (N_9461,N_3294,N_2319);
nor U9462 (N_9462,N_1587,N_4745);
nand U9463 (N_9463,N_4656,N_1573);
or U9464 (N_9464,N_2513,N_696);
and U9465 (N_9465,N_2280,N_4859);
and U9466 (N_9466,N_2320,N_4914);
and U9467 (N_9467,N_2485,N_329);
nand U9468 (N_9468,N_3840,N_246);
nand U9469 (N_9469,N_4428,N_2214);
nor U9470 (N_9470,N_2577,N_184);
nor U9471 (N_9471,N_256,N_1087);
xor U9472 (N_9472,N_731,N_1774);
and U9473 (N_9473,N_214,N_4873);
xnor U9474 (N_9474,N_51,N_2500);
or U9475 (N_9475,N_2212,N_3983);
xnor U9476 (N_9476,N_3354,N_2632);
and U9477 (N_9477,N_4411,N_2705);
nand U9478 (N_9478,N_3876,N_1674);
or U9479 (N_9479,N_1595,N_3763);
nor U9480 (N_9480,N_226,N_2280);
or U9481 (N_9481,N_819,N_3301);
xnor U9482 (N_9482,N_589,N_3190);
or U9483 (N_9483,N_3160,N_3283);
nor U9484 (N_9484,N_334,N_2551);
or U9485 (N_9485,N_3344,N_280);
or U9486 (N_9486,N_836,N_3471);
xnor U9487 (N_9487,N_4337,N_248);
nor U9488 (N_9488,N_4443,N_1782);
and U9489 (N_9489,N_3241,N_2919);
nor U9490 (N_9490,N_680,N_1660);
nand U9491 (N_9491,N_1505,N_4578);
and U9492 (N_9492,N_534,N_3727);
nor U9493 (N_9493,N_836,N_771);
nor U9494 (N_9494,N_3105,N_4107);
nor U9495 (N_9495,N_2722,N_4436);
nor U9496 (N_9496,N_4239,N_3406);
nor U9497 (N_9497,N_2503,N_576);
and U9498 (N_9498,N_941,N_4993);
nor U9499 (N_9499,N_2259,N_1473);
nand U9500 (N_9500,N_2806,N_4381);
or U9501 (N_9501,N_1115,N_873);
and U9502 (N_9502,N_669,N_1577);
nand U9503 (N_9503,N_2627,N_2452);
nand U9504 (N_9504,N_2575,N_4966);
and U9505 (N_9505,N_2343,N_2567);
or U9506 (N_9506,N_4155,N_1266);
and U9507 (N_9507,N_4564,N_3487);
or U9508 (N_9508,N_1648,N_3173);
and U9509 (N_9509,N_4711,N_3412);
and U9510 (N_9510,N_2343,N_1569);
nand U9511 (N_9511,N_2512,N_1225);
nor U9512 (N_9512,N_780,N_3820);
and U9513 (N_9513,N_632,N_3464);
nor U9514 (N_9514,N_158,N_2343);
or U9515 (N_9515,N_3437,N_1445);
nand U9516 (N_9516,N_2234,N_396);
and U9517 (N_9517,N_2378,N_3187);
nand U9518 (N_9518,N_3592,N_4624);
nand U9519 (N_9519,N_1701,N_223);
or U9520 (N_9520,N_115,N_684);
nor U9521 (N_9521,N_4244,N_3452);
nor U9522 (N_9522,N_2352,N_1179);
or U9523 (N_9523,N_1357,N_618);
or U9524 (N_9524,N_3169,N_1562);
or U9525 (N_9525,N_2954,N_2806);
nand U9526 (N_9526,N_4269,N_1057);
nand U9527 (N_9527,N_2185,N_1484);
and U9528 (N_9528,N_4858,N_3661);
nand U9529 (N_9529,N_4953,N_4312);
and U9530 (N_9530,N_1157,N_2504);
and U9531 (N_9531,N_1846,N_1426);
nor U9532 (N_9532,N_120,N_2509);
and U9533 (N_9533,N_4315,N_2958);
and U9534 (N_9534,N_4856,N_1407);
and U9535 (N_9535,N_3044,N_4620);
nand U9536 (N_9536,N_4115,N_3750);
nor U9537 (N_9537,N_3383,N_3282);
or U9538 (N_9538,N_3777,N_2319);
nor U9539 (N_9539,N_4697,N_2668);
nor U9540 (N_9540,N_1902,N_1690);
and U9541 (N_9541,N_2516,N_4461);
or U9542 (N_9542,N_3403,N_697);
and U9543 (N_9543,N_2495,N_714);
nand U9544 (N_9544,N_3930,N_1801);
or U9545 (N_9545,N_978,N_1826);
nor U9546 (N_9546,N_3398,N_3521);
and U9547 (N_9547,N_3303,N_1251);
nor U9548 (N_9548,N_1506,N_4785);
and U9549 (N_9549,N_2279,N_4322);
and U9550 (N_9550,N_3218,N_2952);
nand U9551 (N_9551,N_4337,N_1882);
or U9552 (N_9552,N_152,N_4247);
or U9553 (N_9553,N_211,N_2770);
nor U9554 (N_9554,N_3397,N_2178);
nand U9555 (N_9555,N_597,N_3356);
or U9556 (N_9556,N_4016,N_302);
or U9557 (N_9557,N_2612,N_3579);
or U9558 (N_9558,N_2813,N_3951);
and U9559 (N_9559,N_1421,N_2395);
xor U9560 (N_9560,N_2762,N_4633);
nand U9561 (N_9561,N_4802,N_2924);
nor U9562 (N_9562,N_4895,N_1911);
nand U9563 (N_9563,N_1227,N_3082);
nor U9564 (N_9564,N_1000,N_3043);
and U9565 (N_9565,N_2760,N_264);
nand U9566 (N_9566,N_4863,N_4411);
nor U9567 (N_9567,N_3652,N_4897);
nand U9568 (N_9568,N_4837,N_865);
and U9569 (N_9569,N_173,N_4285);
nand U9570 (N_9570,N_4008,N_1690);
and U9571 (N_9571,N_3135,N_1938);
xnor U9572 (N_9572,N_2109,N_2003);
nand U9573 (N_9573,N_1732,N_4);
nand U9574 (N_9574,N_3943,N_2440);
and U9575 (N_9575,N_4623,N_1045);
xor U9576 (N_9576,N_4375,N_4578);
and U9577 (N_9577,N_1318,N_2199);
xor U9578 (N_9578,N_2208,N_584);
nand U9579 (N_9579,N_816,N_315);
or U9580 (N_9580,N_2154,N_114);
nor U9581 (N_9581,N_171,N_4985);
nand U9582 (N_9582,N_3361,N_1655);
and U9583 (N_9583,N_538,N_3422);
nor U9584 (N_9584,N_2152,N_1247);
xnor U9585 (N_9585,N_4802,N_3537);
nor U9586 (N_9586,N_2829,N_439);
and U9587 (N_9587,N_909,N_3111);
nor U9588 (N_9588,N_4712,N_4789);
nand U9589 (N_9589,N_4121,N_2366);
and U9590 (N_9590,N_117,N_3381);
or U9591 (N_9591,N_798,N_205);
or U9592 (N_9592,N_485,N_2167);
nor U9593 (N_9593,N_1197,N_344);
nand U9594 (N_9594,N_2226,N_1729);
nand U9595 (N_9595,N_3186,N_4586);
or U9596 (N_9596,N_4374,N_2047);
xnor U9597 (N_9597,N_1499,N_79);
nand U9598 (N_9598,N_1176,N_3896);
nand U9599 (N_9599,N_1399,N_921);
and U9600 (N_9600,N_2484,N_4484);
nand U9601 (N_9601,N_3497,N_2751);
or U9602 (N_9602,N_2743,N_3927);
or U9603 (N_9603,N_807,N_2912);
and U9604 (N_9604,N_2396,N_2225);
and U9605 (N_9605,N_1,N_374);
xnor U9606 (N_9606,N_256,N_2799);
nor U9607 (N_9607,N_81,N_4856);
nor U9608 (N_9608,N_3090,N_4814);
and U9609 (N_9609,N_1614,N_1046);
nand U9610 (N_9610,N_1014,N_2655);
nor U9611 (N_9611,N_1735,N_4040);
and U9612 (N_9612,N_3994,N_2313);
or U9613 (N_9613,N_843,N_94);
and U9614 (N_9614,N_1244,N_31);
nor U9615 (N_9615,N_2943,N_949);
nand U9616 (N_9616,N_1152,N_3629);
and U9617 (N_9617,N_4985,N_2947);
nand U9618 (N_9618,N_4820,N_2292);
or U9619 (N_9619,N_3905,N_326);
and U9620 (N_9620,N_3427,N_3357);
and U9621 (N_9621,N_1530,N_4469);
nor U9622 (N_9622,N_29,N_4421);
xor U9623 (N_9623,N_4790,N_3521);
or U9624 (N_9624,N_3455,N_4056);
xnor U9625 (N_9625,N_3724,N_3301);
nor U9626 (N_9626,N_414,N_825);
nand U9627 (N_9627,N_2767,N_148);
and U9628 (N_9628,N_360,N_1330);
nor U9629 (N_9629,N_3415,N_2273);
xnor U9630 (N_9630,N_611,N_2272);
and U9631 (N_9631,N_860,N_3092);
nand U9632 (N_9632,N_2524,N_739);
nand U9633 (N_9633,N_1478,N_3051);
xnor U9634 (N_9634,N_3934,N_2972);
nor U9635 (N_9635,N_3985,N_4104);
nand U9636 (N_9636,N_1834,N_2446);
nor U9637 (N_9637,N_4094,N_3867);
or U9638 (N_9638,N_3298,N_1679);
nor U9639 (N_9639,N_2741,N_580);
and U9640 (N_9640,N_2450,N_1879);
and U9641 (N_9641,N_1147,N_3488);
nand U9642 (N_9642,N_3983,N_470);
or U9643 (N_9643,N_2775,N_4658);
and U9644 (N_9644,N_240,N_1789);
and U9645 (N_9645,N_4081,N_3277);
xor U9646 (N_9646,N_3115,N_4188);
xor U9647 (N_9647,N_4622,N_2076);
xnor U9648 (N_9648,N_3986,N_3283);
xor U9649 (N_9649,N_1015,N_4500);
or U9650 (N_9650,N_1308,N_4624);
nand U9651 (N_9651,N_3371,N_3361);
and U9652 (N_9652,N_487,N_2671);
nand U9653 (N_9653,N_1035,N_145);
and U9654 (N_9654,N_3987,N_2459);
or U9655 (N_9655,N_378,N_111);
xor U9656 (N_9656,N_3901,N_2953);
nor U9657 (N_9657,N_322,N_4016);
nand U9658 (N_9658,N_3370,N_2026);
and U9659 (N_9659,N_2585,N_4227);
nand U9660 (N_9660,N_1819,N_1830);
nor U9661 (N_9661,N_688,N_4350);
or U9662 (N_9662,N_4037,N_1599);
nor U9663 (N_9663,N_1218,N_284);
nor U9664 (N_9664,N_241,N_2460);
nand U9665 (N_9665,N_1933,N_624);
and U9666 (N_9666,N_2172,N_4111);
nor U9667 (N_9667,N_4291,N_747);
nand U9668 (N_9668,N_4815,N_2079);
nor U9669 (N_9669,N_3691,N_2949);
nor U9670 (N_9670,N_2260,N_788);
xnor U9671 (N_9671,N_3717,N_4350);
nor U9672 (N_9672,N_1119,N_2660);
and U9673 (N_9673,N_2912,N_217);
nand U9674 (N_9674,N_1969,N_3482);
nand U9675 (N_9675,N_2815,N_852);
nor U9676 (N_9676,N_167,N_2200);
nand U9677 (N_9677,N_297,N_3781);
nand U9678 (N_9678,N_750,N_3000);
and U9679 (N_9679,N_1364,N_3032);
nor U9680 (N_9680,N_1782,N_3730);
and U9681 (N_9681,N_1961,N_149);
or U9682 (N_9682,N_1973,N_3395);
nor U9683 (N_9683,N_3622,N_2931);
nor U9684 (N_9684,N_3580,N_2624);
or U9685 (N_9685,N_4945,N_1574);
nor U9686 (N_9686,N_4053,N_1113);
or U9687 (N_9687,N_1907,N_4585);
nor U9688 (N_9688,N_3457,N_3196);
nand U9689 (N_9689,N_124,N_3097);
nand U9690 (N_9690,N_2326,N_3141);
or U9691 (N_9691,N_1706,N_905);
and U9692 (N_9692,N_3839,N_123);
nand U9693 (N_9693,N_934,N_1779);
xnor U9694 (N_9694,N_1899,N_1848);
or U9695 (N_9695,N_3705,N_223);
and U9696 (N_9696,N_3911,N_4459);
and U9697 (N_9697,N_4465,N_3287);
and U9698 (N_9698,N_3858,N_3431);
and U9699 (N_9699,N_315,N_1260);
or U9700 (N_9700,N_440,N_2888);
nand U9701 (N_9701,N_547,N_3094);
xnor U9702 (N_9702,N_584,N_1821);
nor U9703 (N_9703,N_2949,N_292);
nor U9704 (N_9704,N_3932,N_538);
nand U9705 (N_9705,N_1737,N_3676);
and U9706 (N_9706,N_2791,N_773);
nand U9707 (N_9707,N_1681,N_2472);
nand U9708 (N_9708,N_1704,N_2225);
or U9709 (N_9709,N_2694,N_4880);
or U9710 (N_9710,N_1672,N_2300);
and U9711 (N_9711,N_4015,N_3981);
nand U9712 (N_9712,N_1679,N_4933);
or U9713 (N_9713,N_3288,N_1841);
nor U9714 (N_9714,N_4776,N_1913);
nand U9715 (N_9715,N_4532,N_4110);
nor U9716 (N_9716,N_4215,N_2347);
xnor U9717 (N_9717,N_3567,N_431);
nor U9718 (N_9718,N_3247,N_1595);
xor U9719 (N_9719,N_286,N_3757);
and U9720 (N_9720,N_2171,N_921);
and U9721 (N_9721,N_4700,N_4416);
xnor U9722 (N_9722,N_1701,N_4159);
nand U9723 (N_9723,N_2712,N_2988);
nand U9724 (N_9724,N_912,N_3223);
and U9725 (N_9725,N_4449,N_3213);
nand U9726 (N_9726,N_4497,N_4375);
nor U9727 (N_9727,N_2421,N_2725);
nand U9728 (N_9728,N_3518,N_4060);
and U9729 (N_9729,N_541,N_749);
nand U9730 (N_9730,N_3232,N_3965);
and U9731 (N_9731,N_3370,N_2342);
and U9732 (N_9732,N_276,N_2655);
xor U9733 (N_9733,N_62,N_2930);
or U9734 (N_9734,N_1316,N_3337);
or U9735 (N_9735,N_4348,N_1671);
or U9736 (N_9736,N_881,N_4706);
or U9737 (N_9737,N_3369,N_26);
nor U9738 (N_9738,N_4355,N_3585);
and U9739 (N_9739,N_47,N_2110);
and U9740 (N_9740,N_1567,N_4287);
nor U9741 (N_9741,N_4690,N_2114);
or U9742 (N_9742,N_3177,N_803);
nor U9743 (N_9743,N_4964,N_2209);
and U9744 (N_9744,N_2937,N_4896);
and U9745 (N_9745,N_140,N_4083);
or U9746 (N_9746,N_706,N_1229);
or U9747 (N_9747,N_1616,N_4598);
nor U9748 (N_9748,N_300,N_4594);
nor U9749 (N_9749,N_2491,N_2577);
and U9750 (N_9750,N_1680,N_2430);
nor U9751 (N_9751,N_3167,N_3939);
xnor U9752 (N_9752,N_2237,N_1238);
nor U9753 (N_9753,N_1013,N_1393);
and U9754 (N_9754,N_1518,N_1764);
nor U9755 (N_9755,N_2347,N_4559);
nand U9756 (N_9756,N_4281,N_146);
nand U9757 (N_9757,N_2016,N_1693);
and U9758 (N_9758,N_2649,N_2368);
nor U9759 (N_9759,N_818,N_3737);
and U9760 (N_9760,N_2203,N_3593);
nand U9761 (N_9761,N_2889,N_3777);
or U9762 (N_9762,N_1289,N_741);
nand U9763 (N_9763,N_20,N_1425);
nand U9764 (N_9764,N_738,N_2881);
or U9765 (N_9765,N_2263,N_3554);
xnor U9766 (N_9766,N_3920,N_1072);
or U9767 (N_9767,N_490,N_1136);
or U9768 (N_9768,N_4019,N_2942);
nor U9769 (N_9769,N_3316,N_947);
nand U9770 (N_9770,N_2064,N_170);
or U9771 (N_9771,N_3922,N_4570);
nand U9772 (N_9772,N_1131,N_1908);
nor U9773 (N_9773,N_1027,N_1933);
nor U9774 (N_9774,N_3477,N_3938);
or U9775 (N_9775,N_4319,N_4927);
xor U9776 (N_9776,N_1851,N_3150);
nor U9777 (N_9777,N_3526,N_3020);
nor U9778 (N_9778,N_1943,N_4919);
and U9779 (N_9779,N_344,N_4000);
nand U9780 (N_9780,N_2219,N_2948);
nor U9781 (N_9781,N_982,N_2789);
and U9782 (N_9782,N_2297,N_1749);
nand U9783 (N_9783,N_4859,N_1136);
or U9784 (N_9784,N_3870,N_66);
nand U9785 (N_9785,N_2305,N_3742);
and U9786 (N_9786,N_439,N_2704);
or U9787 (N_9787,N_2690,N_3422);
xor U9788 (N_9788,N_1653,N_1598);
nor U9789 (N_9789,N_2776,N_418);
and U9790 (N_9790,N_3193,N_3302);
nor U9791 (N_9791,N_1626,N_385);
and U9792 (N_9792,N_2667,N_4099);
and U9793 (N_9793,N_4142,N_1257);
nand U9794 (N_9794,N_1754,N_4641);
nor U9795 (N_9795,N_2653,N_2551);
nand U9796 (N_9796,N_2786,N_606);
or U9797 (N_9797,N_4233,N_4387);
or U9798 (N_9798,N_662,N_3720);
nand U9799 (N_9799,N_2315,N_1774);
and U9800 (N_9800,N_4120,N_3667);
nor U9801 (N_9801,N_3512,N_4953);
nor U9802 (N_9802,N_4436,N_2600);
and U9803 (N_9803,N_3227,N_4276);
nand U9804 (N_9804,N_2903,N_275);
or U9805 (N_9805,N_1682,N_3074);
nor U9806 (N_9806,N_4855,N_1813);
or U9807 (N_9807,N_2063,N_3484);
nor U9808 (N_9808,N_2391,N_1413);
nand U9809 (N_9809,N_179,N_635);
nor U9810 (N_9810,N_1585,N_1564);
nand U9811 (N_9811,N_638,N_82);
xor U9812 (N_9812,N_4486,N_3798);
and U9813 (N_9813,N_559,N_1867);
xnor U9814 (N_9814,N_2753,N_3288);
nor U9815 (N_9815,N_2044,N_3723);
and U9816 (N_9816,N_3306,N_1273);
nor U9817 (N_9817,N_2593,N_1796);
nand U9818 (N_9818,N_4102,N_4821);
or U9819 (N_9819,N_1558,N_3028);
nor U9820 (N_9820,N_4010,N_3576);
and U9821 (N_9821,N_2274,N_2877);
xnor U9822 (N_9822,N_2388,N_3249);
and U9823 (N_9823,N_4488,N_4399);
and U9824 (N_9824,N_4993,N_1054);
nand U9825 (N_9825,N_67,N_1469);
and U9826 (N_9826,N_3745,N_737);
nor U9827 (N_9827,N_2250,N_1733);
nor U9828 (N_9828,N_2921,N_874);
or U9829 (N_9829,N_1631,N_3360);
or U9830 (N_9830,N_2555,N_4008);
nand U9831 (N_9831,N_3217,N_3031);
and U9832 (N_9832,N_1391,N_2043);
nor U9833 (N_9833,N_2973,N_1227);
and U9834 (N_9834,N_623,N_1906);
and U9835 (N_9835,N_3472,N_1671);
and U9836 (N_9836,N_2935,N_4445);
nor U9837 (N_9837,N_2824,N_585);
nand U9838 (N_9838,N_143,N_2613);
nand U9839 (N_9839,N_2200,N_1655);
or U9840 (N_9840,N_2562,N_2324);
or U9841 (N_9841,N_3858,N_4949);
nand U9842 (N_9842,N_4057,N_2327);
and U9843 (N_9843,N_634,N_4168);
or U9844 (N_9844,N_3906,N_4327);
and U9845 (N_9845,N_2025,N_4564);
and U9846 (N_9846,N_3018,N_4324);
and U9847 (N_9847,N_4445,N_3137);
or U9848 (N_9848,N_1615,N_4422);
xnor U9849 (N_9849,N_876,N_4023);
or U9850 (N_9850,N_866,N_4208);
nand U9851 (N_9851,N_2129,N_164);
or U9852 (N_9852,N_1341,N_4551);
or U9853 (N_9853,N_3293,N_140);
nor U9854 (N_9854,N_877,N_646);
nor U9855 (N_9855,N_838,N_424);
or U9856 (N_9856,N_1842,N_4710);
and U9857 (N_9857,N_2937,N_2381);
nand U9858 (N_9858,N_297,N_3156);
nand U9859 (N_9859,N_3204,N_1562);
nor U9860 (N_9860,N_2834,N_1033);
and U9861 (N_9861,N_3976,N_4970);
and U9862 (N_9862,N_3316,N_2982);
nor U9863 (N_9863,N_4741,N_3646);
or U9864 (N_9864,N_1848,N_1966);
nand U9865 (N_9865,N_1095,N_2497);
nor U9866 (N_9866,N_1244,N_2179);
nor U9867 (N_9867,N_630,N_274);
nand U9868 (N_9868,N_4451,N_4195);
nor U9869 (N_9869,N_4071,N_4804);
xor U9870 (N_9870,N_4919,N_1602);
xnor U9871 (N_9871,N_1577,N_32);
or U9872 (N_9872,N_3571,N_1619);
and U9873 (N_9873,N_2917,N_2874);
nor U9874 (N_9874,N_3884,N_1834);
and U9875 (N_9875,N_619,N_1073);
or U9876 (N_9876,N_2963,N_1563);
nand U9877 (N_9877,N_3072,N_376);
and U9878 (N_9878,N_3243,N_4189);
nand U9879 (N_9879,N_2374,N_4956);
nor U9880 (N_9880,N_4743,N_216);
nand U9881 (N_9881,N_4663,N_3079);
and U9882 (N_9882,N_1375,N_2940);
xnor U9883 (N_9883,N_1678,N_1113);
nand U9884 (N_9884,N_4760,N_2777);
nand U9885 (N_9885,N_675,N_1116);
nor U9886 (N_9886,N_4097,N_3951);
nand U9887 (N_9887,N_2898,N_807);
nor U9888 (N_9888,N_1478,N_1841);
nand U9889 (N_9889,N_157,N_1253);
nand U9890 (N_9890,N_213,N_3748);
nor U9891 (N_9891,N_1534,N_4481);
and U9892 (N_9892,N_3914,N_2873);
or U9893 (N_9893,N_2444,N_76);
or U9894 (N_9894,N_1998,N_4506);
xor U9895 (N_9895,N_1952,N_234);
nor U9896 (N_9896,N_3153,N_204);
or U9897 (N_9897,N_746,N_2054);
and U9898 (N_9898,N_4989,N_3270);
and U9899 (N_9899,N_295,N_1745);
nand U9900 (N_9900,N_3150,N_4172);
or U9901 (N_9901,N_3800,N_1832);
or U9902 (N_9902,N_4512,N_309);
and U9903 (N_9903,N_4695,N_268);
nor U9904 (N_9904,N_4971,N_2551);
nand U9905 (N_9905,N_1522,N_3365);
nor U9906 (N_9906,N_3204,N_2103);
and U9907 (N_9907,N_4456,N_2469);
and U9908 (N_9908,N_2126,N_2821);
and U9909 (N_9909,N_199,N_1022);
nor U9910 (N_9910,N_3443,N_3745);
xor U9911 (N_9911,N_213,N_764);
or U9912 (N_9912,N_3120,N_3985);
or U9913 (N_9913,N_3203,N_1736);
or U9914 (N_9914,N_4290,N_3939);
xnor U9915 (N_9915,N_3349,N_506);
nand U9916 (N_9916,N_370,N_3951);
xnor U9917 (N_9917,N_1555,N_4296);
and U9918 (N_9918,N_2680,N_2053);
or U9919 (N_9919,N_3612,N_2331);
nand U9920 (N_9920,N_94,N_1913);
nand U9921 (N_9921,N_555,N_1472);
nor U9922 (N_9922,N_1234,N_2437);
and U9923 (N_9923,N_4228,N_4375);
nand U9924 (N_9924,N_898,N_4110);
nor U9925 (N_9925,N_2139,N_1188);
or U9926 (N_9926,N_2078,N_1015);
nor U9927 (N_9927,N_587,N_37);
or U9928 (N_9928,N_3671,N_3708);
nor U9929 (N_9929,N_4258,N_3723);
or U9930 (N_9930,N_4267,N_2411);
and U9931 (N_9931,N_1905,N_670);
nor U9932 (N_9932,N_2608,N_1713);
nand U9933 (N_9933,N_4497,N_1869);
nor U9934 (N_9934,N_1594,N_3462);
nand U9935 (N_9935,N_1373,N_3222);
nand U9936 (N_9936,N_71,N_3008);
and U9937 (N_9937,N_1570,N_405);
nor U9938 (N_9938,N_919,N_2488);
nand U9939 (N_9939,N_2638,N_931);
nor U9940 (N_9940,N_3644,N_3481);
nand U9941 (N_9941,N_2744,N_4820);
nor U9942 (N_9942,N_3447,N_1999);
nand U9943 (N_9943,N_1836,N_1942);
xnor U9944 (N_9944,N_1634,N_3984);
or U9945 (N_9945,N_3065,N_1630);
nor U9946 (N_9946,N_4580,N_4611);
or U9947 (N_9947,N_317,N_822);
and U9948 (N_9948,N_4987,N_3516);
nor U9949 (N_9949,N_4831,N_3574);
xnor U9950 (N_9950,N_169,N_2803);
nor U9951 (N_9951,N_3612,N_2935);
and U9952 (N_9952,N_2268,N_1145);
nor U9953 (N_9953,N_1776,N_2338);
nand U9954 (N_9954,N_1217,N_1210);
or U9955 (N_9955,N_1033,N_3856);
nor U9956 (N_9956,N_2353,N_4675);
or U9957 (N_9957,N_2666,N_601);
or U9958 (N_9958,N_2897,N_7);
nand U9959 (N_9959,N_1467,N_4680);
and U9960 (N_9960,N_1249,N_251);
nor U9961 (N_9961,N_1918,N_2493);
nand U9962 (N_9962,N_4297,N_3911);
or U9963 (N_9963,N_3934,N_3629);
xnor U9964 (N_9964,N_4470,N_267);
or U9965 (N_9965,N_4515,N_1414);
nor U9966 (N_9966,N_4015,N_865);
and U9967 (N_9967,N_181,N_3940);
or U9968 (N_9968,N_830,N_1335);
and U9969 (N_9969,N_3492,N_1625);
nand U9970 (N_9970,N_4412,N_3952);
xor U9971 (N_9971,N_4499,N_295);
or U9972 (N_9972,N_3571,N_1070);
and U9973 (N_9973,N_4453,N_915);
nand U9974 (N_9974,N_2792,N_3652);
nor U9975 (N_9975,N_199,N_1360);
and U9976 (N_9976,N_108,N_59);
nand U9977 (N_9977,N_651,N_902);
and U9978 (N_9978,N_2624,N_3125);
nand U9979 (N_9979,N_4156,N_4892);
or U9980 (N_9980,N_3751,N_2855);
nand U9981 (N_9981,N_3806,N_4518);
nand U9982 (N_9982,N_2009,N_3279);
nand U9983 (N_9983,N_3393,N_4157);
nor U9984 (N_9984,N_3945,N_846);
nand U9985 (N_9985,N_4349,N_3905);
and U9986 (N_9986,N_793,N_1679);
and U9987 (N_9987,N_1021,N_1281);
and U9988 (N_9988,N_3860,N_4035);
nor U9989 (N_9989,N_1790,N_1515);
and U9990 (N_9990,N_1874,N_1870);
and U9991 (N_9991,N_3710,N_180);
xor U9992 (N_9992,N_2474,N_887);
or U9993 (N_9993,N_3655,N_3903);
nand U9994 (N_9994,N_4615,N_4017);
or U9995 (N_9995,N_1689,N_281);
nor U9996 (N_9996,N_2825,N_2016);
and U9997 (N_9997,N_4430,N_4665);
nand U9998 (N_9998,N_3709,N_4422);
or U9999 (N_9999,N_1267,N_2417);
and UO_0 (O_0,N_6502,N_9656);
or UO_1 (O_1,N_9123,N_5119);
nand UO_2 (O_2,N_8213,N_6690);
nand UO_3 (O_3,N_9835,N_7916);
nor UO_4 (O_4,N_7315,N_8624);
or UO_5 (O_5,N_5894,N_8152);
nor UO_6 (O_6,N_9690,N_7025);
or UO_7 (O_7,N_7650,N_8205);
nand UO_8 (O_8,N_6283,N_7055);
and UO_9 (O_9,N_5570,N_9038);
and UO_10 (O_10,N_7716,N_9039);
nand UO_11 (O_11,N_8869,N_9019);
nand UO_12 (O_12,N_9865,N_8469);
nor UO_13 (O_13,N_8558,N_9618);
nand UO_14 (O_14,N_6011,N_6014);
nor UO_15 (O_15,N_5340,N_5114);
and UO_16 (O_16,N_5231,N_5493);
nand UO_17 (O_17,N_8841,N_8037);
nor UO_18 (O_18,N_8410,N_5776);
nor UO_19 (O_19,N_9716,N_9630);
nand UO_20 (O_20,N_5760,N_5310);
or UO_21 (O_21,N_8982,N_8741);
or UO_22 (O_22,N_9883,N_5984);
and UO_23 (O_23,N_8656,N_5382);
nor UO_24 (O_24,N_9501,N_5679);
or UO_25 (O_25,N_5128,N_7148);
nand UO_26 (O_26,N_9767,N_6811);
and UO_27 (O_27,N_9349,N_8803);
nand UO_28 (O_28,N_6185,N_5741);
and UO_29 (O_29,N_5354,N_6121);
nand UO_30 (O_30,N_5139,N_9706);
nor UO_31 (O_31,N_6106,N_7727);
or UO_32 (O_32,N_9686,N_9156);
or UO_33 (O_33,N_7160,N_7282);
and UO_34 (O_34,N_8640,N_6929);
and UO_35 (O_35,N_7965,N_7860);
nand UO_36 (O_36,N_8540,N_5737);
or UO_37 (O_37,N_5545,N_7381);
xor UO_38 (O_38,N_6926,N_8694);
nor UO_39 (O_39,N_8542,N_7131);
and UO_40 (O_40,N_6751,N_5014);
nor UO_41 (O_41,N_8069,N_8700);
nor UO_42 (O_42,N_8605,N_5288);
xnor UO_43 (O_43,N_5380,N_6209);
and UO_44 (O_44,N_8371,N_5873);
xnor UO_45 (O_45,N_5284,N_7618);
nor UO_46 (O_46,N_9814,N_5186);
nand UO_47 (O_47,N_6272,N_5283);
xor UO_48 (O_48,N_8862,N_6331);
nand UO_49 (O_49,N_9827,N_6732);
nor UO_50 (O_50,N_6369,N_7599);
and UO_51 (O_51,N_7781,N_9774);
and UO_52 (O_52,N_7762,N_7214);
and UO_53 (O_53,N_8137,N_9059);
or UO_54 (O_54,N_9890,N_7324);
or UO_55 (O_55,N_5764,N_6301);
and UO_56 (O_56,N_5488,N_9866);
nor UO_57 (O_57,N_5924,N_9722);
or UO_58 (O_58,N_7022,N_9046);
or UO_59 (O_59,N_8008,N_5278);
or UO_60 (O_60,N_6675,N_9175);
nor UO_61 (O_61,N_6386,N_6229);
xnor UO_62 (O_62,N_8986,N_8330);
and UO_63 (O_63,N_5978,N_9284);
nor UO_64 (O_64,N_8182,N_5026);
or UO_65 (O_65,N_7646,N_7308);
xnor UO_66 (O_66,N_5790,N_6716);
nand UO_67 (O_67,N_6473,N_7597);
xor UO_68 (O_68,N_6536,N_8419);
xnor UO_69 (O_69,N_9447,N_8439);
or UO_70 (O_70,N_5561,N_5677);
nand UO_71 (O_71,N_7546,N_8948);
nand UO_72 (O_72,N_6561,N_7752);
and UO_73 (O_73,N_5357,N_7979);
xnor UO_74 (O_74,N_6578,N_9267);
and UO_75 (O_75,N_9237,N_6029);
or UO_76 (O_76,N_9747,N_9943);
or UO_77 (O_77,N_7510,N_5345);
and UO_78 (O_78,N_8563,N_7127);
nand UO_79 (O_79,N_9083,N_6171);
nor UO_80 (O_80,N_7012,N_7070);
nand UO_81 (O_81,N_7643,N_6443);
nand UO_82 (O_82,N_6162,N_8661);
and UO_83 (O_83,N_9592,N_6784);
or UO_84 (O_84,N_5890,N_6157);
or UO_85 (O_85,N_9430,N_6005);
nor UO_86 (O_86,N_5242,N_9666);
or UO_87 (O_87,N_7483,N_8922);
and UO_88 (O_88,N_9704,N_8141);
or UO_89 (O_89,N_9578,N_8114);
nor UO_90 (O_90,N_8874,N_5848);
or UO_91 (O_91,N_8883,N_6187);
or UO_92 (O_92,N_5210,N_9180);
and UO_93 (O_93,N_8895,N_7385);
or UO_94 (O_94,N_6507,N_5851);
nor UO_95 (O_95,N_8085,N_5951);
nor UO_96 (O_96,N_7641,N_5176);
or UO_97 (O_97,N_6225,N_9266);
or UO_98 (O_98,N_9373,N_5774);
nor UO_99 (O_99,N_5451,N_8523);
nor UO_100 (O_100,N_7318,N_9781);
nor UO_101 (O_101,N_5557,N_7761);
or UO_102 (O_102,N_7427,N_8489);
and UO_103 (O_103,N_5225,N_8003);
xor UO_104 (O_104,N_9877,N_7233);
xor UO_105 (O_105,N_6633,N_6679);
xnor UO_106 (O_106,N_6115,N_5312);
or UO_107 (O_107,N_7718,N_5083);
nor UO_108 (O_108,N_6923,N_5359);
and UO_109 (O_109,N_5842,N_9031);
or UO_110 (O_110,N_9107,N_9422);
and UO_111 (O_111,N_8849,N_6122);
and UO_112 (O_112,N_5480,N_5755);
nor UO_113 (O_113,N_7463,N_6695);
and UO_114 (O_114,N_5930,N_7925);
and UO_115 (O_115,N_5292,N_6437);
nand UO_116 (O_116,N_5030,N_5510);
nand UO_117 (O_117,N_6799,N_8500);
and UO_118 (O_118,N_5019,N_7533);
nor UO_119 (O_119,N_7742,N_5765);
and UO_120 (O_120,N_5917,N_8192);
xor UO_121 (O_121,N_6248,N_9973);
and UO_122 (O_122,N_7656,N_9541);
and UO_123 (O_123,N_8011,N_5908);
or UO_124 (O_124,N_5934,N_9380);
or UO_125 (O_125,N_5901,N_7059);
or UO_126 (O_126,N_9624,N_6391);
xnor UO_127 (O_127,N_5853,N_6656);
nor UO_128 (O_128,N_6859,N_6697);
and UO_129 (O_129,N_5604,N_8712);
nor UO_130 (O_130,N_9869,N_9138);
and UO_131 (O_131,N_9872,N_9389);
or UO_132 (O_132,N_7583,N_6688);
or UO_133 (O_133,N_5950,N_8284);
or UO_134 (O_134,N_6589,N_6983);
or UO_135 (O_135,N_7484,N_6550);
nand UO_136 (O_136,N_7156,N_5259);
nor UO_137 (O_137,N_5174,N_6252);
nor UO_138 (O_138,N_8349,N_9050);
and UO_139 (O_139,N_8308,N_6280);
nand UO_140 (O_140,N_7569,N_9862);
or UO_141 (O_141,N_8253,N_7467);
nand UO_142 (O_142,N_9269,N_7926);
nand UO_143 (O_143,N_5825,N_5454);
or UO_144 (O_144,N_6650,N_8448);
nand UO_145 (O_145,N_5562,N_6532);
nand UO_146 (O_146,N_8083,N_6471);
nor UO_147 (O_147,N_6465,N_9566);
and UO_148 (O_148,N_8888,N_6292);
and UO_149 (O_149,N_5203,N_8739);
xor UO_150 (O_150,N_7283,N_6189);
nand UO_151 (O_151,N_6211,N_8842);
or UO_152 (O_152,N_8262,N_5516);
xor UO_153 (O_153,N_6995,N_5372);
nor UO_154 (O_154,N_9150,N_8742);
and UO_155 (O_155,N_6474,N_5618);
xor UO_156 (O_156,N_5205,N_5500);
or UO_157 (O_157,N_7627,N_7655);
or UO_158 (O_158,N_6717,N_9661);
nand UO_159 (O_159,N_9252,N_7540);
nand UO_160 (O_160,N_5374,N_8794);
or UO_161 (O_161,N_7645,N_6613);
nand UO_162 (O_162,N_5206,N_6462);
xor UO_163 (O_163,N_8549,N_6708);
nor UO_164 (O_164,N_8671,N_8642);
nand UO_165 (O_165,N_6313,N_5385);
nand UO_166 (O_166,N_8290,N_8520);
xnor UO_167 (O_167,N_8186,N_5366);
or UO_168 (O_168,N_7375,N_6523);
nand UO_169 (O_169,N_9412,N_9343);
or UO_170 (O_170,N_9069,N_7654);
nor UO_171 (O_171,N_7937,N_6050);
nor UO_172 (O_172,N_6054,N_7256);
or UO_173 (O_173,N_8957,N_9864);
nor UO_174 (O_174,N_5746,N_5511);
nand UO_175 (O_175,N_7271,N_6623);
and UO_176 (O_176,N_6164,N_9705);
nand UO_177 (O_177,N_7945,N_8394);
or UO_178 (O_178,N_7877,N_5450);
xor UO_179 (O_179,N_5182,N_7601);
or UO_180 (O_180,N_5102,N_7554);
nor UO_181 (O_181,N_8648,N_9001);
and UO_182 (O_182,N_8943,N_8239);
nand UO_183 (O_183,N_7311,N_9418);
nand UO_184 (O_184,N_9789,N_7773);
and UO_185 (O_185,N_5486,N_5255);
nand UO_186 (O_186,N_6264,N_8416);
nand UO_187 (O_187,N_7091,N_7608);
and UO_188 (O_188,N_7913,N_5680);
or UO_189 (O_189,N_9505,N_9845);
nand UO_190 (O_190,N_7259,N_6776);
and UO_191 (O_191,N_7732,N_7394);
and UO_192 (O_192,N_9891,N_9336);
nand UO_193 (O_193,N_9633,N_6348);
nor UO_194 (O_194,N_8270,N_6144);
and UO_195 (O_195,N_5802,N_6707);
or UO_196 (O_196,N_6582,N_5389);
or UO_197 (O_197,N_9625,N_5520);
xor UO_198 (O_198,N_9547,N_8594);
or UO_199 (O_199,N_7389,N_8571);
nand UO_200 (O_200,N_5796,N_9688);
nor UO_201 (O_201,N_8357,N_5140);
xor UO_202 (O_202,N_5969,N_5675);
or UO_203 (O_203,N_6748,N_7740);
nor UO_204 (O_204,N_8465,N_9832);
nand UO_205 (O_205,N_8493,N_9427);
nand UO_206 (O_206,N_8036,N_8731);
and UO_207 (O_207,N_5335,N_6401);
nand UO_208 (O_208,N_5834,N_9730);
nor UO_209 (O_209,N_7966,N_5410);
and UO_210 (O_210,N_5620,N_5935);
nor UO_211 (O_211,N_7472,N_9752);
or UO_212 (O_212,N_7614,N_6130);
nor UO_213 (O_213,N_8325,N_7900);
or UO_214 (O_214,N_7011,N_8578);
nand UO_215 (O_215,N_5564,N_5074);
nor UO_216 (O_216,N_7356,N_8909);
and UO_217 (O_217,N_6538,N_7465);
and UO_218 (O_218,N_6944,N_8052);
xnor UO_219 (O_219,N_7217,N_8335);
xnor UO_220 (O_220,N_6807,N_5364);
or UO_221 (O_221,N_5398,N_5353);
or UO_222 (O_222,N_6008,N_7274);
nor UO_223 (O_223,N_6019,N_5243);
nor UO_224 (O_224,N_7139,N_7558);
nor UO_225 (O_225,N_9939,N_8272);
or UO_226 (O_226,N_5303,N_9215);
nor UO_227 (O_227,N_9571,N_9463);
nor UO_228 (O_228,N_9948,N_5948);
or UO_229 (O_229,N_7499,N_5282);
or UO_230 (O_230,N_9406,N_9590);
nor UO_231 (O_231,N_7671,N_7522);
nand UO_232 (O_232,N_8659,N_7553);
nor UO_233 (O_233,N_7009,N_5336);
xor UO_234 (O_234,N_6953,N_9112);
or UO_235 (O_235,N_5350,N_5734);
xnor UO_236 (O_236,N_7154,N_6948);
and UO_237 (O_237,N_6546,N_8299);
nor UO_238 (O_238,N_9852,N_5285);
or UO_239 (O_239,N_9998,N_7192);
and UO_240 (O_240,N_9365,N_8004);
xor UO_241 (O_241,N_6302,N_7056);
or UO_242 (O_242,N_5491,N_5705);
and UO_243 (O_243,N_5578,N_8858);
and UO_244 (O_244,N_9196,N_7286);
or UO_245 (O_245,N_5418,N_8702);
or UO_246 (O_246,N_5168,N_9466);
or UO_247 (O_247,N_6579,N_5246);
and UO_248 (O_248,N_8810,N_9576);
and UO_249 (O_249,N_6376,N_5309);
or UO_250 (O_250,N_6739,N_8538);
or UO_251 (O_251,N_9410,N_5332);
nand UO_252 (O_252,N_7545,N_6678);
nand UO_253 (O_253,N_8893,N_8176);
or UO_254 (O_254,N_7221,N_6778);
or UO_255 (O_255,N_5905,N_6152);
nand UO_256 (O_256,N_9785,N_7038);
and UO_257 (O_257,N_6960,N_6986);
nor UO_258 (O_258,N_6262,N_6200);
and UO_259 (O_259,N_9441,N_9639);
xnor UO_260 (O_260,N_6093,N_5936);
or UO_261 (O_261,N_8374,N_5982);
or UO_262 (O_262,N_8147,N_8025);
xnor UO_263 (O_263,N_5770,N_8720);
and UO_264 (O_264,N_7493,N_7096);
nor UO_265 (O_265,N_6873,N_9980);
nand UO_266 (O_266,N_7788,N_7088);
or UO_267 (O_267,N_8696,N_6745);
or UO_268 (O_268,N_9489,N_9022);
nor UO_269 (O_269,N_6676,N_6468);
nor UO_270 (O_270,N_9439,N_5038);
or UO_271 (O_271,N_5082,N_7017);
and UO_272 (O_272,N_6082,N_8851);
or UO_273 (O_273,N_8464,N_5191);
or UO_274 (O_274,N_5272,N_9593);
nor UO_275 (O_275,N_7756,N_7713);
nand UO_276 (O_276,N_5120,N_5762);
nand UO_277 (O_277,N_6850,N_6057);
nor UO_278 (O_278,N_6563,N_9428);
xnor UO_279 (O_279,N_5458,N_8120);
xnor UO_280 (O_280,N_9532,N_8363);
nor UO_281 (O_281,N_5022,N_9581);
or UO_282 (O_282,N_9841,N_8414);
nor UO_283 (O_283,N_9670,N_9111);
and UO_284 (O_284,N_5788,N_5548);
nor UO_285 (O_285,N_7751,N_9293);
nand UO_286 (O_286,N_9924,N_6237);
nand UO_287 (O_287,N_9659,N_8440);
or UO_288 (O_288,N_6750,N_7336);
or UO_289 (O_289,N_9619,N_8250);
and UO_290 (O_290,N_6950,N_9265);
nor UO_291 (O_291,N_5773,N_6062);
or UO_292 (O_292,N_9354,N_5196);
nand UO_293 (O_293,N_8166,N_6868);
nor UO_294 (O_294,N_5820,N_9680);
and UO_295 (O_295,N_7120,N_5724);
and UO_296 (O_296,N_7093,N_8522);
and UO_297 (O_297,N_7099,N_9333);
or UO_298 (O_298,N_5207,N_9512);
nor UO_299 (O_299,N_9017,N_8942);
nor UO_300 (O_300,N_7352,N_8055);
nor UO_301 (O_301,N_6774,N_6116);
and UO_302 (O_302,N_9340,N_8993);
or UO_303 (O_303,N_6284,N_9302);
nor UO_304 (O_304,N_8698,N_5714);
nand UO_305 (O_305,N_5659,N_7531);
and UO_306 (O_306,N_8265,N_5147);
nor UO_307 (O_307,N_5388,N_5478);
nand UO_308 (O_308,N_9339,N_9753);
nor UO_309 (O_309,N_9476,N_9596);
and UO_310 (O_310,N_7485,N_8859);
or UO_311 (O_311,N_6981,N_7117);
and UO_312 (O_312,N_9213,N_9074);
nand UO_313 (O_313,N_5142,N_9916);
nand UO_314 (O_314,N_8499,N_6744);
and UO_315 (O_315,N_5965,N_5743);
nor UO_316 (O_316,N_6119,N_8660);
or UO_317 (O_317,N_5800,N_6661);
nand UO_318 (O_318,N_9321,N_5944);
nand UO_319 (O_319,N_9126,N_6344);
nand UO_320 (O_320,N_6927,N_9411);
and UO_321 (O_321,N_8399,N_6781);
or UO_322 (O_322,N_8161,N_6439);
nor UO_323 (O_323,N_6681,N_8506);
nand UO_324 (O_324,N_6531,N_5290);
nor UO_325 (O_325,N_8564,N_9109);
and UO_326 (O_326,N_8980,N_7580);
nand UO_327 (O_327,N_8344,N_9308);
nor UO_328 (O_328,N_8057,N_7669);
nor UO_329 (O_329,N_6037,N_6444);
nand UO_330 (O_330,N_7133,N_5116);
or UO_331 (O_331,N_7125,N_8669);
or UO_332 (O_332,N_7365,N_5673);
and UO_333 (O_333,N_8310,N_9366);
and UO_334 (O_334,N_9499,N_7053);
xnor UO_335 (O_335,N_8769,N_6300);
or UO_336 (O_336,N_8101,N_7097);
and UO_337 (O_337,N_9057,N_9882);
nor UO_338 (O_338,N_9455,N_5202);
or UO_339 (O_339,N_9531,N_7799);
nor UO_340 (O_340,N_8907,N_5730);
and UO_341 (O_341,N_8206,N_6890);
or UO_342 (O_342,N_6087,N_5429);
and UO_343 (O_343,N_7261,N_8601);
nand UO_344 (O_344,N_7887,N_5927);
nand UO_345 (O_345,N_7803,N_7862);
nor UO_346 (O_346,N_9514,N_8743);
and UO_347 (O_347,N_5914,N_8733);
nor UO_348 (O_348,N_9162,N_9740);
or UO_349 (O_349,N_8067,N_8384);
or UO_350 (O_350,N_5327,N_6504);
and UO_351 (O_351,N_6274,N_5968);
or UO_352 (O_352,N_9967,N_5736);
or UO_353 (O_353,N_8925,N_9529);
nor UO_354 (O_354,N_9047,N_9174);
nor UO_355 (O_355,N_9444,N_6573);
or UO_356 (O_356,N_8573,N_6640);
nand UO_357 (O_357,N_6101,N_8482);
or UO_358 (O_358,N_6442,N_7869);
nor UO_359 (O_359,N_7208,N_5213);
or UO_360 (O_360,N_8546,N_8595);
nor UO_361 (O_361,N_6878,N_5852);
nor UO_362 (O_362,N_5293,N_6077);
and UO_363 (O_363,N_6993,N_9679);
or UO_364 (O_364,N_5660,N_5702);
nor UO_365 (O_365,N_5123,N_6492);
and UO_366 (O_366,N_7068,N_5286);
and UO_367 (O_367,N_7206,N_9816);
nand UO_368 (O_368,N_7210,N_5668);
or UO_369 (O_369,N_9152,N_5011);
nand UO_370 (O_370,N_9671,N_6315);
or UO_371 (O_371,N_8710,N_8430);
xor UO_372 (O_372,N_8073,N_7513);
nand UO_373 (O_373,N_9936,N_8471);
nand UO_374 (O_374,N_8480,N_9966);
and UO_375 (O_375,N_8646,N_8593);
nand UO_376 (O_376,N_6400,N_7305);
or UO_377 (O_377,N_5404,N_6931);
nand UO_378 (O_378,N_5509,N_9243);
nor UO_379 (O_379,N_5402,N_8800);
and UO_380 (O_380,N_5329,N_5121);
nor UO_381 (O_381,N_9133,N_5165);
xor UO_382 (O_382,N_6622,N_9648);
and UO_383 (O_383,N_8816,N_6168);
and UO_384 (O_384,N_7258,N_8086);
nand UO_385 (O_385,N_9521,N_7600);
nand UO_386 (O_386,N_5087,N_6520);
or UO_387 (O_387,N_5069,N_7045);
xnor UO_388 (O_388,N_9240,N_9926);
or UO_389 (O_389,N_6755,N_7419);
nand UO_390 (O_390,N_6730,N_7052);
or UO_391 (O_391,N_9609,N_9110);
and UO_392 (O_392,N_6322,N_6773);
xnor UO_393 (O_393,N_7201,N_6449);
or UO_394 (O_394,N_6997,N_9689);
nor UO_395 (O_395,N_8583,N_6421);
or UO_396 (O_396,N_5596,N_8876);
or UO_397 (O_397,N_5068,N_5792);
or UO_398 (O_398,N_6770,N_5882);
nand UO_399 (O_399,N_7827,N_5624);
nand UO_400 (O_400,N_8704,N_7598);
nand UO_401 (O_401,N_9762,N_6296);
and UO_402 (O_402,N_6245,N_6565);
and UO_403 (O_403,N_5099,N_8579);
and UO_404 (O_404,N_7710,N_7351);
nor UO_405 (O_405,N_9600,N_8806);
xnor UO_406 (O_406,N_8050,N_9895);
and UO_407 (O_407,N_6371,N_5972);
or UO_408 (O_408,N_6310,N_5637);
nor UO_409 (O_409,N_6634,N_8387);
or UO_410 (O_410,N_5862,N_9121);
or UO_411 (O_411,N_9726,N_6306);
nor UO_412 (O_412,N_6888,N_6904);
nand UO_413 (O_413,N_7503,N_8474);
or UO_414 (O_414,N_8054,N_6629);
nand UO_415 (O_415,N_8829,N_9408);
nor UO_416 (O_416,N_9440,N_7188);
and UO_417 (O_417,N_7632,N_6255);
nor UO_418 (O_418,N_6801,N_7368);
and UO_419 (O_419,N_9602,N_9280);
or UO_420 (O_420,N_9260,N_8863);
xnor UO_421 (O_421,N_7146,N_9734);
and UO_422 (O_422,N_8225,N_6407);
and UO_423 (O_423,N_9524,N_8144);
and UO_424 (O_424,N_6571,N_5096);
xnor UO_425 (O_425,N_5735,N_5392);
nand UO_426 (O_426,N_5996,N_7584);
nand UO_427 (O_427,N_8297,N_6682);
or UO_428 (O_428,N_8437,N_7143);
nand UO_429 (O_429,N_6259,N_8717);
nand UO_430 (O_430,N_7683,N_9419);
nand UO_431 (O_431,N_6798,N_6089);
xor UO_432 (O_432,N_6420,N_6092);
nor UO_433 (O_433,N_8001,N_5425);
nor UO_434 (O_434,N_9802,N_6509);
or UO_435 (O_435,N_7586,N_6103);
and UO_436 (O_436,N_7574,N_5367);
nor UO_437 (O_437,N_9509,N_7880);
nand UO_438 (O_438,N_6281,N_5412);
nand UO_439 (O_439,N_5532,N_8596);
nand UO_440 (O_440,N_7891,N_9459);
nor UO_441 (O_441,N_5199,N_7452);
or UO_442 (O_442,N_6244,N_8931);
or UO_443 (O_443,N_6406,N_7940);
and UO_444 (O_444,N_7280,N_8047);
xor UO_445 (O_445,N_5428,N_8808);
nand UO_446 (O_446,N_9842,N_9176);
nand UO_447 (O_447,N_9635,N_9935);
and UO_448 (O_448,N_5148,N_5895);
or UO_449 (O_449,N_6642,N_8928);
nor UO_450 (O_450,N_9815,N_8031);
nor UO_451 (O_451,N_5177,N_8867);
xor UO_452 (O_452,N_6261,N_5056);
or UO_453 (O_453,N_7329,N_7129);
nand UO_454 (O_454,N_6911,N_9077);
and UO_455 (O_455,N_5617,N_8600);
and UO_456 (O_456,N_5455,N_8209);
nor UO_457 (O_457,N_9383,N_9575);
nor UO_458 (O_458,N_7157,N_9338);
and UO_459 (O_459,N_8028,N_5431);
nand UO_460 (O_460,N_7679,N_5300);
or UO_461 (O_461,N_9070,N_5048);
nor UO_462 (O_462,N_8107,N_8606);
nand UO_463 (O_463,N_5221,N_6308);
or UO_464 (O_464,N_8537,N_7456);
or UO_465 (O_465,N_7473,N_5178);
nand UO_466 (O_466,N_5163,N_8901);
nor UO_467 (O_467,N_8764,N_6984);
nand UO_468 (O_468,N_8309,N_8956);
and UO_469 (O_469,N_6901,N_7783);
nand UO_470 (O_470,N_6139,N_8119);
nand UO_471 (O_471,N_6769,N_7634);
or UO_472 (O_472,N_7084,N_9251);
and UO_473 (O_473,N_5274,N_9248);
and UO_474 (O_474,N_5024,N_8984);
or UO_475 (O_475,N_8099,N_5910);
nand UO_476 (O_476,N_9390,N_9925);
or UO_477 (O_477,N_7345,N_7947);
xnor UO_478 (O_478,N_9120,N_7290);
or UO_479 (O_479,N_9961,N_6783);
nand UO_480 (O_480,N_9229,N_9130);
and UO_481 (O_481,N_7898,N_6729);
nand UO_482 (O_482,N_9292,N_6405);
nand UO_483 (O_483,N_8745,N_8026);
and UO_484 (O_484,N_5744,N_9674);
or UO_485 (O_485,N_5467,N_5479);
xor UO_486 (O_486,N_9553,N_8976);
and UO_487 (O_487,N_8170,N_6714);
or UO_488 (O_488,N_6108,N_6949);
xor UO_489 (O_489,N_7486,N_5645);
xnor UO_490 (O_490,N_9095,N_5523);
and UO_491 (O_491,N_8826,N_6686);
nor UO_492 (O_492,N_7527,N_9369);
and UO_493 (O_493,N_5883,N_8496);
nor UO_494 (O_494,N_8655,N_5721);
nand UO_495 (O_495,N_8840,N_6232);
or UO_496 (O_496,N_5236,N_8965);
xor UO_497 (O_497,N_9350,N_8779);
and UO_498 (O_498,N_7453,N_7841);
or UO_499 (O_499,N_8449,N_6459);
nor UO_500 (O_500,N_9561,N_6012);
xnor UO_501 (O_501,N_5400,N_7934);
and UO_502 (O_502,N_5193,N_9614);
and UO_503 (O_503,N_6040,N_5158);
nor UO_504 (O_504,N_6549,N_9040);
and UO_505 (O_505,N_9487,N_5994);
xnor UO_506 (O_506,N_5573,N_7046);
or UO_507 (O_507,N_7791,N_6326);
and UO_508 (O_508,N_8681,N_9777);
nor UO_509 (O_509,N_6742,N_7114);
nor UO_510 (O_510,N_8685,N_9342);
nor UO_511 (O_511,N_5568,N_9402);
and UO_512 (O_512,N_7760,N_5470);
and UO_513 (O_513,N_7507,N_8138);
xnor UO_514 (O_514,N_5289,N_8348);
or UO_515 (O_515,N_8690,N_9222);
nor UO_516 (O_516,N_8163,N_6486);
nand UO_517 (O_517,N_7700,N_6482);
and UO_518 (O_518,N_7470,N_9834);
or UO_519 (O_519,N_8327,N_9309);
nand UO_520 (O_520,N_5416,N_6746);
nor UO_521 (O_521,N_7115,N_7652);
and UO_522 (O_522,N_9723,N_9847);
xnor UO_523 (O_523,N_5577,N_5622);
or UO_524 (O_524,N_6867,N_5466);
nor UO_525 (O_525,N_6109,N_8051);
and UO_526 (O_526,N_9700,N_7272);
xnor UO_527 (O_527,N_5945,N_7487);
and UO_528 (O_528,N_6848,N_6058);
and UO_529 (O_529,N_8090,N_9558);
nor UO_530 (O_530,N_9204,N_9765);
nor UO_531 (O_531,N_7026,N_8706);
nor UO_532 (O_532,N_9496,N_5942);
nand UO_533 (O_533,N_7980,N_5552);
xnor UO_534 (O_534,N_7379,N_7348);
and UO_535 (O_535,N_6385,N_5145);
nand UO_536 (O_536,N_7811,N_6317);
nor UO_537 (O_537,N_5507,N_7338);
or UO_538 (O_538,N_8625,N_5727);
and UO_539 (O_539,N_6847,N_9060);
and UO_540 (O_540,N_9497,N_6887);
xnor UO_541 (O_541,N_8457,N_6253);
or UO_542 (O_542,N_7142,N_6488);
and UO_543 (O_543,N_7076,N_5827);
and UO_544 (O_544,N_9500,N_6754);
xnor UO_545 (O_545,N_8766,N_8255);
nor UO_546 (O_546,N_9300,N_8807);
or UO_547 (O_547,N_5763,N_9794);
and UO_548 (O_548,N_8080,N_5940);
nand UO_549 (O_549,N_6829,N_7956);
nor UO_550 (O_550,N_6711,N_9868);
or UO_551 (O_551,N_5368,N_8329);
or UO_552 (O_552,N_8729,N_9537);
nand UO_553 (O_553,N_9885,N_7058);
and UO_554 (O_554,N_6197,N_9937);
or UO_555 (O_555,N_9992,N_5137);
nor UO_556 (O_556,N_7865,N_5756);
or UO_557 (O_557,N_5542,N_6869);
or UO_558 (O_558,N_7255,N_7508);
nor UO_559 (O_559,N_7968,N_6341);
or UO_560 (O_560,N_7222,N_8827);
nand UO_561 (O_561,N_7204,N_9116);
xnor UO_562 (O_562,N_8814,N_7986);
nand UO_563 (O_563,N_9950,N_9914);
or UO_564 (O_564,N_9557,N_6114);
xor UO_565 (O_565,N_6199,N_7984);
nor UO_566 (O_566,N_7414,N_5828);
or UO_567 (O_567,N_7014,N_7778);
nand UO_568 (O_568,N_6988,N_7387);
nor UO_569 (O_569,N_6767,N_7357);
or UO_570 (O_570,N_5269,N_6660);
nand UO_571 (O_571,N_8454,N_5990);
nor UO_572 (O_572,N_8136,N_7624);
nor UO_573 (O_573,N_7443,N_8959);
nor UO_574 (O_574,N_5248,N_6599);
nor UO_575 (O_575,N_9699,N_5926);
nor UO_576 (O_576,N_5817,N_7298);
nand UO_577 (O_577,N_5794,N_7666);
nor UO_578 (O_578,N_8332,N_5481);
or UO_579 (O_579,N_6818,N_9783);
or UO_580 (O_580,N_9528,N_9755);
nor UO_581 (O_581,N_9084,N_5611);
nand UO_582 (O_582,N_5918,N_9048);
and UO_583 (O_583,N_5785,N_7777);
nand UO_584 (O_584,N_6166,N_9892);
nand UO_585 (O_585,N_9153,N_7295);
nor UO_586 (O_586,N_8488,N_8834);
nand UO_587 (O_587,N_5156,N_5266);
or UO_588 (O_588,N_7343,N_8342);
and UO_589 (O_589,N_8804,N_6052);
xnor UO_590 (O_590,N_7615,N_7587);
and UO_591 (O_591,N_5150,N_8110);
nand UO_592 (O_592,N_7585,N_9894);
nand UO_593 (O_593,N_8762,N_7103);
xor UO_594 (O_594,N_7220,N_8498);
nor UO_595 (O_595,N_8491,N_8260);
xnor UO_596 (O_596,N_6045,N_5995);
or UO_597 (O_597,N_6947,N_9995);
nor UO_598 (O_598,N_5860,N_5261);
or UO_599 (O_599,N_9757,N_9970);
or UO_600 (O_600,N_7000,N_5589);
xnor UO_601 (O_601,N_7896,N_7861);
and UO_602 (O_602,N_9559,N_7260);
and UO_603 (O_603,N_9977,N_9654);
nand UO_604 (O_604,N_8664,N_9607);
or UO_605 (O_605,N_6145,N_9201);
nor UO_606 (O_606,N_7675,N_5343);
nor UO_607 (O_607,N_5339,N_5981);
nand UO_608 (O_608,N_6372,N_5931);
or UO_609 (O_609,N_7479,N_9053);
or UO_610 (O_610,N_8039,N_6733);
and UO_611 (O_611,N_8179,N_7300);
or UO_612 (O_612,N_6435,N_6380);
nand UO_613 (O_613,N_8006,N_5085);
or UO_614 (O_614,N_9432,N_7409);
nor UO_615 (O_615,N_6820,N_5889);
or UO_616 (O_616,N_7176,N_8584);
xor UO_617 (O_617,N_5584,N_7595);
or UO_618 (O_618,N_6156,N_6409);
xor UO_619 (O_619,N_6074,N_5447);
nor UO_620 (O_620,N_7450,N_8095);
xnor UO_621 (O_621,N_5194,N_5234);
nand UO_622 (O_622,N_6417,N_5487);
and UO_623 (O_623,N_6620,N_6893);
or UO_624 (O_624,N_6364,N_9364);
nor UO_625 (O_625,N_7653,N_6396);
or UO_626 (O_626,N_9003,N_8091);
nor UO_627 (O_627,N_9029,N_8515);
and UO_628 (O_628,N_9856,N_5021);
or UO_629 (O_629,N_7853,N_7322);
nor UO_630 (O_630,N_7041,N_6985);
nand UO_631 (O_631,N_7873,N_5387);
or UO_632 (O_632,N_9464,N_7548);
nor UO_633 (O_633,N_7207,N_5781);
nand UO_634 (O_634,N_8828,N_5007);
nand UO_635 (O_635,N_7064,N_5494);
nor UO_636 (O_636,N_8273,N_5649);
nand UO_637 (O_637,N_9420,N_6503);
nor UO_638 (O_638,N_5775,N_7517);
or UO_639 (O_639,N_5461,N_9525);
or UO_640 (O_640,N_6143,N_8908);
xor UO_641 (O_641,N_8049,N_8351);
and UO_642 (O_642,N_9801,N_6354);
nand UO_643 (O_643,N_8597,N_8402);
nand UO_644 (O_644,N_7972,N_6349);
nand UO_645 (O_645,N_9965,N_6632);
and UO_646 (O_646,N_7455,N_6120);
and UO_647 (O_647,N_8390,N_5818);
or UO_648 (O_648,N_9304,N_5826);
nor UO_649 (O_649,N_5612,N_6128);
nor UO_650 (O_650,N_7771,N_6936);
nand UO_651 (O_651,N_9170,N_8755);
and UO_652 (O_652,N_8372,N_5215);
nand UO_653 (O_653,N_5050,N_7894);
nor UO_654 (O_654,N_8767,N_8075);
xnor UO_655 (O_655,N_7571,N_7870);
and UO_656 (O_656,N_8652,N_6693);
or UO_657 (O_657,N_8635,N_8033);
and UO_658 (O_658,N_6782,N_5915);
nor UO_659 (O_659,N_7137,N_6854);
nand UO_660 (O_660,N_5761,N_6652);
nor UO_661 (O_661,N_6954,N_9072);
nand UO_662 (O_662,N_6375,N_7951);
xor UO_663 (O_663,N_5819,N_9375);
nand UO_664 (O_664,N_8792,N_8038);
xnor UO_665 (O_665,N_5258,N_7448);
nor UO_666 (O_666,N_8629,N_7094);
or UO_667 (O_667,N_5653,N_5769);
and UO_668 (O_668,N_9443,N_9217);
xnor UO_669 (O_669,N_9850,N_8797);
and UO_670 (O_670,N_6670,N_9232);
or UO_671 (O_671,N_9858,N_9135);
nor UO_672 (O_672,N_6448,N_8367);
nand UO_673 (O_673,N_6466,N_7904);
and UO_674 (O_674,N_9416,N_5426);
nor UO_675 (O_675,N_6938,N_5081);
xor UO_676 (O_676,N_7689,N_8856);
nor UO_677 (O_677,N_6337,N_7130);
nand UO_678 (O_678,N_8268,N_7248);
nand UO_679 (O_679,N_6666,N_8425);
xor UO_680 (O_680,N_7189,N_9480);
nand UO_681 (O_681,N_6163,N_5229);
and UO_682 (O_682,N_7661,N_7876);
nand UO_683 (O_683,N_8929,N_8125);
xnor UO_684 (O_684,N_5672,N_7008);
nand UO_685 (O_685,N_5433,N_7028);
nand UO_686 (O_686,N_5569,N_8846);
nand UO_687 (O_687,N_8598,N_5436);
nand UO_688 (O_688,N_9506,N_5443);
nor UO_689 (O_689,N_6227,N_7337);
and UO_690 (O_690,N_6343,N_7899);
and UO_691 (O_691,N_6456,N_7605);
nand UO_692 (O_692,N_5797,N_9736);
and UO_693 (O_693,N_6881,N_9224);
nand UO_694 (O_694,N_7538,N_5157);
nor UO_695 (O_695,N_8756,N_8626);
or UO_696 (O_696,N_7745,N_8760);
nand UO_697 (O_697,N_5344,N_9043);
nand UO_698 (O_698,N_7294,N_8586);
or UO_699 (O_699,N_9317,N_7209);
nand UO_700 (O_700,N_5117,N_7040);
and UO_701 (O_701,N_9288,N_7858);
or UO_702 (O_702,N_5829,N_9928);
or UO_703 (O_703,N_6293,N_7572);
and UO_704 (O_704,N_9875,N_8401);
nor UO_705 (O_705,N_6184,N_6533);
or UO_706 (O_706,N_6835,N_9052);
nor UO_707 (O_707,N_5729,N_9037);
nor UO_708 (O_708,N_9164,N_6516);
and UO_709 (O_709,N_8197,N_8056);
nand UO_710 (O_710,N_7955,N_6206);
nor UO_711 (O_711,N_5695,N_5953);
or UO_712 (O_712,N_5413,N_5044);
nand UO_713 (O_713,N_9491,N_9398);
and UO_714 (O_714,N_6594,N_8162);
or UO_715 (O_715,N_6226,N_7285);
or UO_716 (O_716,N_8373,N_9468);
and UO_717 (O_717,N_5448,N_6694);
and UO_718 (O_718,N_9407,N_5656);
or UO_719 (O_719,N_6476,N_6526);
xor UO_720 (O_720,N_6974,N_6294);
nor UO_721 (O_721,N_7500,N_8074);
and UO_722 (O_722,N_5498,N_5909);
and UO_723 (O_723,N_5155,N_7367);
nand UO_724 (O_724,N_6410,N_5218);
nor UO_725 (O_725,N_5983,N_8103);
nor UO_726 (O_726,N_5964,N_6973);
and UO_727 (O_727,N_6939,N_8599);
and UO_728 (O_728,N_5314,N_8236);
xor UO_729 (O_729,N_9548,N_8251);
or UO_730 (O_730,N_9750,N_6856);
or UO_731 (O_731,N_5651,N_6318);
xnor UO_732 (O_732,N_7910,N_5630);
nand UO_733 (O_733,N_5094,N_5307);
nor UO_734 (O_734,N_6601,N_7402);
or UO_735 (O_735,N_5522,N_7095);
xor UO_736 (O_736,N_8012,N_6333);
nand UO_737 (O_737,N_8177,N_6357);
nor UO_738 (O_738,N_5544,N_7037);
xnor UO_739 (O_739,N_8184,N_5200);
nand UO_740 (O_740,N_8428,N_8514);
nand UO_741 (O_741,N_7792,N_8002);
and UO_742 (O_742,N_6618,N_6160);
nor UO_743 (O_743,N_8689,N_5789);
and UO_744 (O_744,N_7067,N_7155);
nand UO_745 (O_745,N_8291,N_9014);
and UO_746 (O_746,N_6689,N_5305);
nand UO_747 (O_747,N_9471,N_6009);
or UO_748 (O_748,N_5420,N_5946);
and UO_749 (O_749,N_5869,N_6937);
nand UO_750 (O_750,N_6908,N_9356);
nor UO_751 (O_751,N_8321,N_7049);
nor UO_752 (O_752,N_5299,N_9401);
nor UO_753 (O_753,N_9761,N_9982);
or UO_754 (O_754,N_5876,N_6104);
or UO_755 (O_755,N_5197,N_5694);
or UO_756 (O_756,N_6070,N_9819);
nand UO_757 (O_757,N_9516,N_7066);
or UO_758 (O_758,N_7119,N_9861);
and UO_759 (O_759,N_5879,N_7889);
or UO_760 (O_760,N_6827,N_5377);
or UO_761 (O_761,N_8683,N_8510);
and UO_762 (O_762,N_6513,N_8771);
xor UO_763 (O_763,N_9588,N_9296);
or UO_764 (O_764,N_6669,N_7818);
and UO_765 (O_765,N_5904,N_9434);
and UO_766 (O_766,N_6311,N_7866);
and UO_767 (O_767,N_6752,N_7191);
and UO_768 (O_768,N_8860,N_7878);
and UO_769 (O_769,N_9631,N_7397);
nand UO_770 (O_770,N_6350,N_7736);
and UO_771 (O_771,N_8183,N_5311);
nor UO_772 (O_772,N_6309,N_5434);
nand UO_773 (O_773,N_5665,N_7253);
and UO_774 (O_774,N_8035,N_6875);
xnor UO_775 (O_775,N_5514,N_5419);
nor UO_776 (O_776,N_6527,N_8413);
and UO_777 (O_777,N_8746,N_9754);
and UO_778 (O_778,N_9098,N_6691);
xor UO_779 (O_779,N_8915,N_5171);
or UO_780 (O_780,N_7223,N_9772);
nand UO_781 (O_781,N_5411,N_8105);
nor UO_782 (O_782,N_9796,N_8978);
and UO_783 (O_783,N_9766,N_9563);
and UO_784 (O_784,N_5088,N_8395);
nand UO_785 (O_785,N_8811,N_6970);
and UO_786 (O_786,N_8296,N_5441);
nand UO_787 (O_787,N_8812,N_7334);
nor UO_788 (O_788,N_6113,N_9396);
or UO_789 (O_789,N_8987,N_5932);
or UO_790 (O_790,N_8463,N_9182);
nand UO_791 (O_791,N_5390,N_5235);
nand UO_792 (O_792,N_7885,N_7042);
nand UO_793 (O_793,N_7344,N_7228);
xnor UO_794 (O_794,N_9193,N_6924);
nor UO_795 (O_795,N_9446,N_9956);
xnor UO_796 (O_796,N_5125,N_9250);
or UO_797 (O_797,N_6575,N_8077);
and UO_798 (O_798,N_8843,N_9582);
nor UO_799 (O_799,N_8825,N_6140);
and UO_800 (O_800,N_9088,N_6025);
and UO_801 (O_801,N_9021,N_8200);
and UO_802 (O_802,N_8716,N_6135);
nand UO_803 (O_803,N_7642,N_7917);
and UO_804 (O_804,N_8616,N_8650);
nor UO_805 (O_805,N_8064,N_8350);
xor UO_806 (O_806,N_6390,N_9687);
nor UO_807 (O_807,N_7748,N_8112);
or UO_808 (O_808,N_9683,N_6416);
xnor UO_809 (O_809,N_7516,N_8603);
and UO_810 (O_810,N_9315,N_8092);
nand UO_811 (O_811,N_7559,N_5499);
or UO_812 (O_812,N_5475,N_6621);
or UO_813 (O_813,N_6543,N_9149);
or UO_814 (O_814,N_8786,N_6946);
nor UO_815 (O_815,N_9685,N_5855);
or UO_816 (O_816,N_5601,N_7623);
nor UO_817 (O_817,N_9634,N_5865);
nor UO_818 (O_818,N_6530,N_6951);
or UO_819 (O_819,N_9194,N_5391);
nand UO_820 (O_820,N_6696,N_8539);
nand UO_821 (O_821,N_6703,N_9066);
nand UO_822 (O_822,N_7701,N_9597);
xor UO_823 (O_823,N_8507,N_6605);
or UO_824 (O_824,N_6556,N_9595);
nor UO_825 (O_825,N_8404,N_5468);
xnor UO_826 (O_826,N_9436,N_7001);
and UO_827 (O_827,N_7593,N_8968);
nor UO_828 (O_828,N_7704,N_8774);
and UO_829 (O_829,N_5063,N_9140);
xnor UO_830 (O_830,N_7677,N_7982);
and UO_831 (O_831,N_8311,N_8164);
nand UO_832 (O_832,N_9488,N_7245);
and UO_833 (O_833,N_8651,N_8058);
nor UO_834 (O_834,N_5899,N_6560);
and UO_835 (O_835,N_5521,N_7964);
or UO_836 (O_836,N_8229,N_5844);
and UO_837 (O_837,N_8732,N_7635);
xnor UO_838 (O_838,N_7476,N_7489);
or UO_839 (O_839,N_9348,N_8392);
or UO_840 (O_840,N_5836,N_5795);
nor UO_841 (O_841,N_5383,N_7403);
nand UO_842 (O_842,N_7447,N_5560);
or UO_843 (O_843,N_9709,N_6863);
or UO_844 (O_844,N_7977,N_5160);
and UO_845 (O_845,N_6006,N_7838);
nand UO_846 (O_846,N_6934,N_8442);
nor UO_847 (O_847,N_9810,N_5766);
and UO_848 (O_848,N_6610,N_9715);
and UO_849 (O_849,N_9825,N_7471);
nand UO_850 (O_850,N_7844,N_9460);
nor UO_851 (O_851,N_6534,N_9258);
nor UO_852 (O_852,N_6071,N_9253);
nand UO_853 (O_853,N_9228,N_8378);
nor UO_854 (O_854,N_9997,N_6928);
nand UO_855 (O_855,N_9800,N_7426);
xor UO_856 (O_856,N_6257,N_9567);
nor UO_857 (O_857,N_8089,N_6470);
or UO_858 (O_858,N_9076,N_7834);
or UO_859 (O_859,N_9955,N_7828);
or UO_860 (O_860,N_7265,N_7250);
xor UO_861 (O_861,N_6684,N_8960);
nand UO_862 (O_862,N_8686,N_7251);
nor UO_863 (O_863,N_9779,N_9203);
and UO_864 (O_864,N_5546,N_5854);
nor UO_865 (O_865,N_7107,N_8787);
and UO_866 (O_866,N_6079,N_8999);
and UO_867 (O_867,N_5166,N_8620);
nor UO_868 (O_868,N_8487,N_7712);
or UO_869 (O_869,N_7162,N_6076);
nor UO_870 (O_870,N_5352,N_8615);
nor UO_871 (O_871,N_8997,N_5295);
xor UO_872 (O_872,N_9361,N_8412);
nor UO_873 (O_873,N_8784,N_8106);
and UO_874 (O_874,N_6886,N_5224);
nand UO_875 (O_875,N_8791,N_6994);
or UO_876 (O_876,N_5941,N_7504);
or UO_877 (O_877,N_6494,N_9867);
nand UO_878 (O_878,N_6658,N_5585);
and UO_879 (O_879,N_8438,N_8521);
nor UO_880 (O_880,N_5519,N_8890);
xnor UO_881 (O_881,N_5581,N_8936);
and UO_882 (O_882,N_9560,N_8424);
or UO_883 (O_883,N_7755,N_5183);
and UO_884 (O_884,N_5275,N_5791);
or UO_885 (O_885,N_7289,N_8305);
and UO_886 (O_886,N_6477,N_8306);
nor UO_887 (O_887,N_9131,N_5629);
nor UO_888 (O_888,N_6802,N_7229);
nor UO_889 (O_889,N_6606,N_8362);
and UO_890 (O_890,N_8718,N_6999);
nor UO_891 (O_891,N_7835,N_5728);
or UO_892 (O_892,N_7789,N_5543);
xnor UO_893 (O_893,N_8478,N_5151);
and UO_894 (O_894,N_8768,N_7071);
nand UO_895 (O_895,N_5365,N_9305);
nor UO_896 (O_896,N_8582,N_8312);
nor UO_897 (O_897,N_7279,N_6933);
and UO_898 (O_898,N_9714,N_8234);
nand UO_899 (O_899,N_6659,N_6794);
or UO_900 (O_900,N_8361,N_7868);
nor UO_901 (O_901,N_9822,N_8240);
xnor UO_902 (O_902,N_6155,N_6587);
nand UO_903 (O_903,N_5563,N_9483);
nand UO_904 (O_904,N_5180,N_6151);
or UO_905 (O_905,N_8320,N_5399);
nor UO_906 (O_906,N_7124,N_7408);
or UO_907 (O_907,N_6201,N_6312);
and UO_908 (O_908,N_9400,N_5136);
or UO_909 (O_909,N_8258,N_8552);
nor UO_910 (O_910,N_7326,N_7768);
nand UO_911 (O_911,N_5749,N_8150);
nor UO_912 (O_912,N_5267,N_6959);
and UO_913 (O_913,N_5974,N_6304);
xor UO_914 (O_914,N_6233,N_7739);
nand UO_915 (O_915,N_5172,N_6644);
and UO_916 (O_916,N_8167,N_8798);
nand UO_917 (O_917,N_7090,N_6860);
nor UO_918 (O_918,N_6617,N_8653);
or UO_919 (O_919,N_7944,N_8916);
and UO_920 (O_920,N_5109,N_8328);
nor UO_921 (O_921,N_9848,N_7100);
nor UO_922 (O_922,N_8623,N_7588);
and UO_923 (O_923,N_5537,N_5706);
and UO_924 (O_924,N_6892,N_5190);
or UO_925 (O_925,N_9081,N_9951);
or UO_926 (O_926,N_6179,N_5881);
nand UO_927 (O_927,N_5527,N_6884);
or UO_928 (O_928,N_5973,N_8981);
and UO_929 (O_929,N_7024,N_6537);
nor UO_930 (O_930,N_9669,N_9197);
and UO_931 (O_931,N_6805,N_7765);
nand UO_932 (O_932,N_8104,N_9863);
and UO_933 (O_933,N_9186,N_8996);
or UO_934 (O_934,N_7929,N_5870);
xor UO_935 (O_935,N_8935,N_7235);
nand UO_936 (O_936,N_7687,N_5625);
and UO_937 (O_937,N_9838,N_7310);
nand UO_938 (O_938,N_5373,N_8575);
nor UO_939 (O_939,N_7607,N_9911);
nor UO_940 (O_940,N_8875,N_9191);
or UO_941 (O_941,N_9523,N_8873);
nor UO_942 (O_942,N_8838,N_6853);
and UO_943 (O_943,N_9313,N_5555);
nand UO_944 (O_944,N_7817,N_7475);
or UO_945 (O_945,N_7183,N_6382);
xor UO_946 (O_946,N_7164,N_8665);
and UO_947 (O_947,N_7047,N_6619);
xor UO_948 (O_948,N_8751,N_9599);
and UO_949 (O_949,N_7376,N_6475);
xor UO_950 (O_950,N_6524,N_9289);
nand UO_951 (O_951,N_6269,N_7254);
xnor UO_952 (O_952,N_7386,N_7171);
or UO_953 (O_953,N_7373,N_6290);
nor UO_954 (O_954,N_7186,N_6921);
or UO_955 (O_955,N_8304,N_5058);
nand UO_956 (O_956,N_7212,N_5553);
nand UO_957 (O_957,N_6624,N_5124);
nand UO_958 (O_958,N_8285,N_8899);
or UO_959 (O_959,N_9117,N_6427);
nand UO_960 (O_960,N_8070,N_8180);
nor UO_961 (O_961,N_8947,N_5967);
nor UO_962 (O_962,N_6445,N_7547);
xnor UO_963 (O_963,N_6167,N_8196);
nor UO_964 (O_964,N_8010,N_8920);
or UO_965 (O_965,N_6517,N_7496);
nand UO_966 (O_966,N_8333,N_7079);
and UO_967 (O_967,N_9254,N_7847);
nand UO_968 (O_968,N_6194,N_6030);
or UO_969 (O_969,N_7976,N_7462);
and UO_970 (O_970,N_9728,N_9075);
and UO_971 (O_971,N_6637,N_7461);
and UO_972 (O_972,N_5490,N_7775);
or UO_973 (O_973,N_6198,N_7726);
nor UO_974 (O_974,N_8585,N_6251);
and UO_975 (O_975,N_7187,N_6150);
or UO_976 (O_976,N_6662,N_6667);
and UO_977 (O_977,N_6759,N_8354);
nor UO_978 (O_978,N_7867,N_6871);
nor UO_979 (O_979,N_6636,N_5065);
nor UO_980 (O_980,N_9393,N_8341);
nor UO_981 (O_981,N_5591,N_6236);
nand UO_982 (O_982,N_7194,N_8097);
xor UO_983 (O_983,N_9676,N_8513);
nand UO_984 (O_984,N_8781,N_9457);
nor UO_985 (O_985,N_5710,N_8618);
or UO_986 (O_986,N_6943,N_9944);
xnor UO_987 (O_987,N_8983,N_8844);
xnor UO_988 (O_988,N_8256,N_6651);
nor UO_989 (O_989,N_8736,N_7826);
nand UO_990 (O_990,N_7705,N_9495);
or UO_991 (O_991,N_8544,N_6849);
and UO_992 (O_992,N_5812,N_5020);
nor UO_993 (O_993,N_5700,N_7879);
or UO_994 (O_994,N_5393,N_7152);
or UO_995 (O_995,N_5167,N_8494);
nand UO_996 (O_996,N_7363,N_7421);
nor UO_997 (O_997,N_6279,N_9776);
xor UO_998 (O_998,N_5241,N_6066);
xnor UO_999 (O_999,N_9731,N_7961);
nand UO_1000 (O_1000,N_5430,N_9183);
and UO_1001 (O_1001,N_7722,N_5216);
nor UO_1002 (O_1002,N_9510,N_6702);
or UO_1003 (O_1003,N_5262,N_8157);
and UO_1004 (O_1004,N_6231,N_7140);
xnor UO_1005 (O_1005,N_7230,N_7449);
nand UO_1006 (O_1006,N_8221,N_5135);
nand UO_1007 (O_1007,N_7110,N_7610);
xor UO_1008 (O_1008,N_5161,N_6004);
xnor UO_1009 (O_1009,N_7092,N_9818);
and UO_1010 (O_1010,N_5871,N_9425);
nand UO_1011 (O_1011,N_7717,N_5325);
or UO_1012 (O_1012,N_7101,N_7872);
nand UO_1013 (O_1013,N_9647,N_8504);
nor UO_1014 (O_1014,N_8817,N_8865);
nand UO_1015 (O_1015,N_7319,N_8020);
nand UO_1016 (O_1016,N_8758,N_5384);
or UO_1017 (O_1017,N_9147,N_5823);
nor UO_1018 (O_1018,N_7438,N_9067);
nand UO_1019 (O_1019,N_6963,N_6511);
nor UO_1020 (O_1020,N_7236,N_6367);
nor UO_1021 (O_1021,N_8788,N_8355);
and UO_1022 (O_1022,N_9458,N_8293);
and UO_1023 (O_1023,N_6855,N_8483);
nor UO_1024 (O_1024,N_7854,N_7730);
and UO_1025 (O_1025,N_6319,N_7893);
xor UO_1026 (O_1026,N_5891,N_9208);
or UO_1027 (O_1027,N_6512,N_6165);
or UO_1028 (O_1028,N_5076,N_7003);
or UO_1029 (O_1029,N_6982,N_7859);
nand UO_1030 (O_1030,N_9873,N_9141);
and UO_1031 (O_1031,N_6379,N_6967);
and UO_1032 (O_1032,N_8433,N_5098);
or UO_1033 (O_1033,N_9173,N_8892);
nor UO_1034 (O_1034,N_9002,N_6183);
nand UO_1035 (O_1035,N_8171,N_8516);
nor UO_1036 (O_1036,N_8382,N_8721);
and UO_1037 (O_1037,N_7815,N_6242);
nor UO_1038 (O_1038,N_7738,N_9504);
nand UO_1039 (O_1039,N_7602,N_6899);
or UO_1040 (O_1040,N_6335,N_5988);
or UO_1041 (O_1041,N_8699,N_6814);
nand UO_1042 (O_1042,N_9665,N_6598);
or UO_1043 (O_1043,N_7630,N_8445);
nand UO_1044 (O_1044,N_8337,N_9782);
nand UO_1045 (O_1045,N_8674,N_8647);
or UO_1046 (O_1046,N_6724,N_8168);
nand UO_1047 (O_1047,N_7823,N_7277);
and UO_1048 (O_1048,N_6501,N_9143);
nor UO_1049 (O_1049,N_6051,N_9684);
or UO_1050 (O_1050,N_9307,N_9157);
or UO_1051 (O_1051,N_5697,N_5530);
xor UO_1052 (O_1052,N_9985,N_9453);
nand UO_1053 (O_1053,N_9058,N_8061);
nor UO_1054 (O_1054,N_8830,N_9118);
or UO_1055 (O_1055,N_8782,N_6497);
nor UO_1056 (O_1056,N_6016,N_8955);
or UO_1057 (O_1057,N_8813,N_7754);
nand UO_1058 (O_1058,N_9996,N_9983);
nand UO_1059 (O_1059,N_5485,N_5877);
or UO_1060 (O_1060,N_5067,N_9530);
and UO_1061 (O_1061,N_6979,N_7609);
or UO_1062 (O_1062,N_9357,N_9902);
and UO_1063 (O_1063,N_8468,N_8129);
nand UO_1064 (O_1064,N_8156,N_7723);
nor UO_1065 (O_1065,N_7902,N_7759);
or UO_1066 (O_1066,N_9231,N_5504);
and UO_1067 (O_1067,N_8417,N_5719);
nand UO_1068 (O_1068,N_5751,N_7425);
or UO_1069 (O_1069,N_5249,N_8204);
and UO_1070 (O_1070,N_6577,N_9484);
nand UO_1071 (O_1071,N_8501,N_6570);
and UO_1072 (O_1072,N_9079,N_8280);
nand UO_1073 (O_1073,N_5189,N_8226);
or UO_1074 (O_1074,N_5438,N_8133);
and UO_1075 (O_1075,N_8722,N_7657);
nand UO_1076 (O_1076,N_9063,N_8405);
xnor UO_1077 (O_1077,N_8032,N_9062);
nand UO_1078 (O_1078,N_9004,N_6677);
nand UO_1079 (O_1079,N_7141,N_9044);
nor UO_1080 (O_1080,N_7393,N_6787);
or UO_1081 (O_1081,N_6731,N_9151);
nor UO_1082 (O_1082,N_5798,N_8676);
nor UO_1083 (O_1083,N_9930,N_9448);
nand UO_1084 (O_1084,N_8301,N_8407);
nor UO_1085 (O_1085,N_5078,N_7080);
or UO_1086 (O_1086,N_5302,N_6920);
or UO_1087 (O_1087,N_5363,N_6616);
nor UO_1088 (O_1088,N_8870,N_6088);
nand UO_1089 (O_1089,N_9012,N_7492);
xor UO_1090 (O_1090,N_7883,N_9210);
and UO_1091 (O_1091,N_9797,N_9192);
nand UO_1092 (O_1092,N_6235,N_5169);
nand UO_1093 (O_1093,N_8805,N_7923);
nand UO_1094 (O_1094,N_5643,N_9554);
nand UO_1095 (O_1095,N_9481,N_5669);
nand UO_1096 (O_1096,N_6440,N_7729);
nand UO_1097 (O_1097,N_8034,N_6844);
and UO_1098 (O_1098,N_8961,N_9534);
xnor UO_1099 (O_1099,N_9426,N_6663);
or UO_1100 (O_1100,N_8836,N_7073);
nand UO_1101 (O_1101,N_9030,N_5962);
nor UO_1102 (O_1102,N_9160,N_8495);
and UO_1103 (O_1103,N_6042,N_9335);
nor UO_1104 (O_1104,N_6351,N_7852);
nand UO_1105 (O_1105,N_6858,N_5403);
and UO_1106 (O_1106,N_9008,N_5032);
nor UO_1107 (O_1107,N_5692,N_8029);
or UO_1108 (O_1108,N_7787,N_9896);
or UO_1109 (O_1109,N_5811,N_8529);
and UO_1110 (O_1110,N_7809,N_5476);
nand UO_1111 (O_1111,N_7313,N_6001);
and UO_1112 (O_1112,N_5489,N_7262);
nand UO_1113 (O_1113,N_8222,N_8211);
nor UO_1114 (O_1114,N_6641,N_9840);
nand UO_1115 (O_1115,N_7981,N_8933);
and UO_1116 (O_1116,N_7316,N_5060);
or UO_1117 (O_1117,N_9080,N_8972);
and UO_1118 (O_1118,N_9912,N_5693);
and UO_1119 (O_1119,N_6060,N_8587);
nand UO_1120 (O_1120,N_6673,N_5998);
nor UO_1121 (O_1121,N_7404,N_9311);
and UO_1122 (O_1122,N_5201,N_9132);
and UO_1123 (O_1123,N_5664,N_7529);
nand UO_1124 (O_1124,N_9763,N_9225);
and UO_1125 (O_1125,N_8898,N_9314);
or UO_1126 (O_1126,N_5041,N_8294);
and UO_1127 (O_1127,N_8886,N_5526);
nor UO_1128 (O_1128,N_8283,N_8632);
nor UO_1129 (O_1129,N_5906,N_7846);
nand UO_1130 (O_1130,N_8279,N_8574);
xnor UO_1131 (O_1131,N_8773,N_5864);
nand UO_1132 (O_1132,N_5005,N_5097);
and UO_1133 (O_1133,N_5772,N_5017);
xor UO_1134 (O_1134,N_6282,N_7933);
or UO_1135 (O_1135,N_6655,N_6793);
or UO_1136 (O_1136,N_5884,N_7061);
or UO_1137 (O_1137,N_7048,N_8589);
xor UO_1138 (O_1138,N_6414,N_6528);
or UO_1139 (O_1139,N_5759,N_7895);
nand UO_1140 (O_1140,N_6846,N_6740);
nor UO_1141 (O_1141,N_6411,N_8878);
or UO_1142 (O_1142,N_8227,N_7383);
and UO_1143 (O_1143,N_9562,N_8602);
nand UO_1144 (O_1144,N_9277,N_6645);
nor UO_1145 (O_1145,N_6797,N_9580);
nand UO_1146 (O_1146,N_8848,N_8649);
xor UO_1147 (O_1147,N_9878,N_6896);
and UO_1148 (O_1148,N_8891,N_5767);
and UO_1149 (O_1149,N_9370,N_5518);
xnor UO_1150 (O_1150,N_7660,N_7715);
nand UO_1151 (O_1151,N_7034,N_5595);
nor UO_1152 (O_1152,N_7764,N_7498);
nand UO_1153 (O_1153,N_7521,N_6142);
nor UO_1154 (O_1154,N_6161,N_5803);
and UO_1155 (O_1155,N_8194,N_8190);
nand UO_1156 (O_1156,N_9799,N_7649);
nand UO_1157 (O_1157,N_5920,N_5588);
xor UO_1158 (O_1158,N_5227,N_6403);
or UO_1159 (O_1159,N_9435,N_9564);
nor UO_1160 (O_1160,N_7914,N_7436);
nand UO_1161 (O_1161,N_6826,N_5631);
or UO_1162 (O_1162,N_7502,N_9351);
nor UO_1163 (O_1163,N_7534,N_9355);
and UO_1164 (O_1164,N_9235,N_7366);
nand UO_1165 (O_1165,N_6271,N_8352);
nor UO_1166 (O_1166,N_9900,N_8113);
nor UO_1167 (O_1167,N_7102,N_7514);
or UO_1168 (O_1168,N_7901,N_9677);
and UO_1169 (O_1169,N_5162,N_6362);
xnor UO_1170 (O_1170,N_7480,N_8917);
and UO_1171 (O_1171,N_9279,N_9849);
or UO_1172 (O_1172,N_8481,N_8952);
or UO_1173 (O_1173,N_6569,N_7526);
and UO_1174 (O_1174,N_6542,N_8286);
or UO_1175 (O_1175,N_9759,N_5265);
nor UO_1176 (O_1176,N_9042,N_9979);
xnor UO_1177 (O_1177,N_7523,N_5551);
nand UO_1178 (O_1178,N_7636,N_6699);
nand UO_1179 (O_1179,N_9093,N_7542);
and UO_1180 (O_1180,N_6027,N_7831);
or UO_1181 (O_1181,N_8765,N_6597);
and UO_1182 (O_1182,N_7165,N_8548);
nand UO_1183 (O_1183,N_9282,N_9820);
and UO_1184 (O_1184,N_9322,N_9828);
or UO_1185 (O_1185,N_8042,N_9932);
or UO_1186 (O_1186,N_9270,N_9811);
nor UO_1187 (O_1187,N_6392,N_5633);
or UO_1188 (O_1188,N_6785,N_8065);
or UO_1189 (O_1189,N_7270,N_6325);
nand UO_1190 (O_1190,N_8318,N_8809);
or UO_1191 (O_1191,N_8340,N_6824);
or UO_1192 (O_1192,N_6572,N_7798);
and UO_1193 (O_1193,N_9089,N_8944);
or UO_1194 (O_1194,N_6895,N_8861);
nand UO_1195 (O_1195,N_6647,N_9113);
nor UO_1196 (O_1196,N_9713,N_5154);
xor UO_1197 (O_1197,N_5574,N_7590);
or UO_1198 (O_1198,N_5252,N_8379);
xnor UO_1199 (O_1199,N_9986,N_5025);
and UO_1200 (O_1200,N_9165,N_8850);
or UO_1201 (O_1201,N_6172,N_7911);
nor UO_1202 (O_1202,N_9791,N_5684);
nand UO_1203 (O_1203,N_7796,N_5506);
nand UO_1204 (O_1204,N_9844,N_8130);
nand UO_1205 (O_1205,N_6205,N_5687);
or UO_1206 (O_1206,N_5104,N_5783);
nand UO_1207 (O_1207,N_7243,N_5676);
or UO_1208 (O_1208,N_7668,N_6250);
xor UO_1209 (O_1209,N_8081,N_7444);
nand UO_1210 (O_1210,N_6836,N_7681);
nor UO_1211 (O_1211,N_9256,N_8554);
nand UO_1212 (O_1212,N_6395,N_8730);
nand UO_1213 (O_1213,N_5992,N_6490);
or UO_1214 (O_1214,N_7327,N_7304);
nor UO_1215 (O_1215,N_6132,N_9287);
nand UO_1216 (O_1216,N_5073,N_8108);
nor UO_1217 (O_1217,N_5517,N_6441);
xor UO_1218 (O_1218,N_8278,N_9839);
and UO_1219 (O_1219,N_8703,N_8005);
nand UO_1220 (O_1220,N_7469,N_8855);
and UO_1221 (O_1221,N_5129,N_7995);
or UO_1222 (O_1222,N_7145,N_5273);
nor UO_1223 (O_1223,N_6882,N_5440);
or UO_1224 (O_1224,N_8015,N_6003);
or UO_1225 (O_1225,N_9876,N_8244);
nor UO_1226 (O_1226,N_8900,N_9855);
and UO_1227 (O_1227,N_9384,N_7999);
or UO_1228 (O_1228,N_9462,N_5623);
nand UO_1229 (O_1229,N_9707,N_8790);
nor UO_1230 (O_1230,N_5036,N_6125);
xnor UO_1231 (O_1231,N_7676,N_8776);
and UO_1232 (O_1232,N_6216,N_8027);
nand UO_1233 (O_1233,N_6241,N_5963);
or UO_1234 (O_1234,N_8281,N_9445);
nand UO_1235 (O_1235,N_7293,N_8233);
and UO_1236 (O_1236,N_7412,N_5449);
or UO_1237 (O_1237,N_6919,N_9735);
nand UO_1238 (O_1238,N_9379,N_9920);
nor UO_1239 (O_1239,N_7793,N_8832);
nor UO_1240 (O_1240,N_5605,N_7203);
and UO_1241 (O_1241,N_8868,N_9108);
and UO_1242 (O_1242,N_6196,N_5501);
or UO_1243 (O_1243,N_7592,N_9627);
or UO_1244 (O_1244,N_7670,N_6256);
nor UO_1245 (O_1245,N_9907,N_8169);
or UO_1246 (O_1246,N_6402,N_5559);
and UO_1247 (O_1247,N_7556,N_7349);
and UO_1248 (O_1248,N_9103,N_6017);
nand UO_1249 (O_1249,N_8531,N_6243);
nand UO_1250 (O_1250,N_8621,N_9691);
xnor UO_1251 (O_1251,N_9465,N_7573);
or UO_1252 (O_1252,N_8257,N_9005);
nor UO_1253 (O_1253,N_5970,N_6906);
and UO_1254 (O_1254,N_9306,N_7983);
nor UO_1255 (O_1255,N_9697,N_9414);
nand UO_1256 (O_1256,N_5439,N_5874);
xor UO_1257 (O_1257,N_5358,N_8819);
or UO_1258 (O_1258,N_5636,N_8154);
nand UO_1259 (O_1259,N_5465,N_7075);
and UO_1260 (O_1260,N_6775,N_7570);
and UO_1261 (O_1261,N_5840,N_5212);
and UO_1262 (O_1262,N_7309,N_8434);
or UO_1263 (O_1263,N_6880,N_6889);
nor UO_1264 (O_1264,N_6991,N_9137);
and UO_1265 (O_1265,N_9696,N_9211);
nand UO_1266 (O_1266,N_7086,N_9438);
and UO_1267 (O_1267,N_6067,N_7638);
or UO_1268 (O_1268,N_8989,N_7741);
xnor UO_1269 (O_1269,N_7335,N_5674);
or UO_1270 (O_1270,N_6419,N_9556);
or UO_1271 (O_1271,N_6436,N_6102);
and UO_1272 (O_1272,N_6036,N_8185);
xnor UO_1273 (O_1273,N_6592,N_8158);
nand UO_1274 (O_1274,N_9572,N_8460);
nor UO_1275 (O_1275,N_8780,N_9129);
and UO_1276 (O_1276,N_5263,N_7832);
and UO_1277 (O_1277,N_8533,N_5688);
nor UO_1278 (O_1278,N_7567,N_5304);
and UO_1279 (O_1279,N_5583,N_6034);
or UO_1280 (O_1280,N_9096,N_9851);
nand UO_1281 (O_1281,N_6429,N_9826);
nor UO_1282 (O_1282,N_6555,N_7620);
nand UO_1283 (O_1283,N_6297,N_5718);
or UO_1284 (O_1284,N_8094,N_9115);
xor UO_1285 (O_1285,N_7264,N_9787);
xor UO_1286 (O_1286,N_9888,N_7341);
or UO_1287 (O_1287,N_9742,N_7106);
xnor UO_1288 (O_1288,N_9431,N_9903);
nand UO_1289 (O_1289,N_8793,N_7330);
nand UO_1290 (O_1290,N_8314,N_7594);
nand UO_1291 (O_1291,N_5786,N_9803);
or UO_1292 (O_1292,N_7974,N_6484);
nor UO_1293 (O_1293,N_9233,N_6032);
and UO_1294 (O_1294,N_7672,N_8668);
nor UO_1295 (O_1295,N_9887,N_9710);
nor UO_1296 (O_1296,N_6968,N_9577);
nor UO_1297 (O_1297,N_9051,N_8377);
nor UO_1298 (O_1298,N_9190,N_7837);
or UO_1299 (O_1299,N_8937,N_8566);
nand UO_1300 (O_1300,N_5960,N_9909);
nand UO_1301 (O_1301,N_7706,N_5348);
nor UO_1302 (O_1302,N_8609,N_7239);
or UO_1303 (O_1303,N_9318,N_7957);
or UO_1304 (O_1304,N_7237,N_8747);
and UO_1305 (O_1305,N_5253,N_7121);
and UO_1306 (O_1306,N_6493,N_9636);
and UO_1307 (O_1307,N_7544,N_5513);
nand UO_1308 (O_1308,N_5423,N_8366);
nor UO_1309 (O_1309,N_7225,N_7030);
or UO_1310 (O_1310,N_7098,N_7709);
nand UO_1311 (O_1311,N_8128,N_7719);
xnor UO_1312 (O_1312,N_7284,N_7520);
or UO_1313 (O_1313,N_9016,N_9055);
and UO_1314 (O_1314,N_6808,N_5331);
nor UO_1315 (O_1315,N_6451,N_9667);
nand UO_1316 (O_1316,N_8954,N_6551);
nand UO_1317 (O_1317,N_5793,N_8235);
and UO_1318 (O_1318,N_8358,N_6083);
nor UO_1319 (O_1319,N_6710,N_8508);
and UO_1320 (O_1320,N_6159,N_8644);
nand UO_1321 (O_1321,N_6314,N_6438);
and UO_1322 (O_1322,N_9477,N_6112);
and UO_1323 (O_1323,N_6741,N_5845);
nand UO_1324 (O_1324,N_9673,N_9768);
nand UO_1325 (O_1325,N_5661,N_6461);
nand UO_1326 (O_1326,N_6932,N_5427);
xor UO_1327 (O_1327,N_5976,N_9923);
nor UO_1328 (O_1328,N_9470,N_6107);
nand UO_1329 (O_1329,N_7177,N_8958);
nand UO_1330 (O_1330,N_9433,N_9234);
nand UO_1331 (O_1331,N_7960,N_7536);
or UO_1332 (O_1332,N_6212,N_8303);
nand UO_1333 (O_1333,N_7382,N_7734);
or UO_1334 (O_1334,N_9122,N_7043);
and UO_1335 (O_1335,N_6234,N_9241);
and UO_1336 (O_1336,N_7728,N_9682);
or UO_1337 (O_1337,N_6202,N_8905);
and UO_1338 (O_1338,N_5315,N_9056);
xor UO_1339 (O_1339,N_7163,N_7678);
or UO_1340 (O_1340,N_6897,N_7054);
nor UO_1341 (O_1341,N_6491,N_5711);
nand UO_1342 (O_1342,N_8053,N_5118);
and UO_1343 (O_1343,N_6447,N_7303);
nand UO_1344 (O_1344,N_8979,N_9745);
and UO_1345 (O_1345,N_7276,N_6627);
and UO_1346 (O_1346,N_9717,N_5460);
xor UO_1347 (O_1347,N_7218,N_7737);
nor UO_1348 (O_1348,N_7429,N_5971);
or UO_1349 (O_1349,N_6839,N_8151);
nor UO_1350 (O_1350,N_5850,N_8924);
or UO_1351 (O_1351,N_7065,N_7857);
nor UO_1352 (O_1352,N_5752,N_8007);
xor UO_1353 (O_1353,N_9913,N_6584);
nor UO_1354 (O_1354,N_7268,N_7795);
or UO_1355 (O_1355,N_9206,N_6332);
nor UO_1356 (O_1356,N_8973,N_8202);
and UO_1357 (O_1357,N_7328,N_5187);
and UO_1358 (O_1358,N_5406,N_8795);
and UO_1359 (O_1359,N_7032,N_6685);
or UO_1360 (O_1360,N_6124,N_8735);
nand UO_1361 (O_1361,N_9405,N_6704);
nor UO_1362 (O_1362,N_6039,N_6224);
and UO_1363 (O_1363,N_8667,N_7193);
or UO_1364 (O_1364,N_6467,N_8208);
nand UO_1365 (O_1365,N_8277,N_7227);
xnor UO_1366 (O_1366,N_7819,N_7010);
nand UO_1367 (O_1367,N_5376,N_7466);
xnor UO_1368 (O_1368,N_5638,N_7537);
or UO_1369 (O_1369,N_6841,N_9486);
xor UO_1370 (O_1370,N_6220,N_8636);
and UO_1371 (O_1371,N_6099,N_7399);
or UO_1372 (O_1372,N_9703,N_6834);
nand UO_1373 (O_1373,N_5888,N_7105);
nand UO_1374 (O_1374,N_8519,N_9589);
or UO_1375 (O_1375,N_8543,N_6182);
nor UO_1376 (O_1376,N_9163,N_8343);
xor UO_1377 (O_1377,N_8452,N_6418);
nor UO_1378 (O_1378,N_5294,N_6687);
nor UO_1379 (O_1379,N_8189,N_5296);
or UO_1380 (O_1380,N_5554,N_8705);
and UO_1381 (O_1381,N_8242,N_6487);
or UO_1382 (O_1382,N_5815,N_6753);
nand UO_1383 (O_1383,N_7242,N_9821);
nand UO_1384 (O_1384,N_5540,N_8436);
nor UO_1385 (O_1385,N_8447,N_6320);
xor UO_1386 (O_1386,N_8926,N_9261);
nor UO_1387 (O_1387,N_6615,N_8016);
and UO_1388 (O_1388,N_7451,N_8093);
or UO_1389 (O_1389,N_5149,N_9181);
or UO_1390 (O_1390,N_7949,N_5947);
nand UO_1391 (O_1391,N_7346,N_7932);
and UO_1392 (O_1392,N_8643,N_7824);
xor UO_1393 (O_1393,N_6260,N_8078);
and UO_1394 (O_1394,N_7060,N_9897);
or UO_1395 (O_1395,N_7063,N_6303);
nand UO_1396 (O_1396,N_9508,N_6608);
and UO_1397 (O_1397,N_5696,N_8096);
xnor UO_1398 (O_1398,N_8397,N_7840);
nor UO_1399 (O_1399,N_9385,N_6489);
and UO_1400 (O_1400,N_9988,N_9169);
xor UO_1401 (O_1401,N_5757,N_8241);
or UO_1402 (O_1402,N_7296,N_5034);
nand UO_1403 (O_1403,N_7987,N_6065);
nand UO_1404 (O_1404,N_9795,N_9168);
nand UO_1405 (O_1405,N_8323,N_9526);
nor UO_1406 (O_1406,N_7912,N_9239);
nand UO_1407 (O_1407,N_7175,N_5536);
or UO_1408 (O_1408,N_9972,N_5152);
nand UO_1409 (O_1409,N_7123,N_5334);
xnor UO_1410 (O_1410,N_8287,N_5435);
nor UO_1411 (O_1411,N_9297,N_9451);
or UO_1412 (O_1412,N_6044,N_6790);
nor UO_1413 (O_1413,N_9751,N_7354);
xor UO_1414 (O_1414,N_7684,N_9473);
nand UO_1415 (O_1415,N_8386,N_7077);
nor UO_1416 (O_1416,N_9533,N_9283);
or UO_1417 (O_1417,N_6323,N_9202);
nand UO_1418 (O_1418,N_8752,N_9346);
nand UO_1419 (O_1419,N_8472,N_8393);
nor UO_1420 (O_1420,N_5841,N_7213);
nor UO_1421 (O_1421,N_7682,N_8775);
and UO_1422 (O_1422,N_6049,N_5223);
or UO_1423 (O_1423,N_7173,N_8633);
nor UO_1424 (O_1424,N_6922,N_5943);
xor UO_1425 (O_1425,N_6771,N_6957);
nand UO_1426 (O_1426,N_9958,N_6519);
nand UO_1427 (O_1427,N_5956,N_5047);
and UO_1428 (O_1428,N_7031,N_9604);
nand UO_1429 (O_1429,N_7801,N_7731);
or UO_1430 (O_1430,N_8214,N_8663);
and UO_1431 (O_1431,N_8921,N_7743);
xnor UO_1432 (O_1432,N_7004,N_7699);
or UO_1433 (O_1433,N_7190,N_7197);
and UO_1434 (O_1434,N_5370,N_9010);
or UO_1435 (O_1435,N_9854,N_7935);
and UO_1436 (O_1436,N_9472,N_9144);
or UO_1437 (O_1437,N_6270,N_8068);
nor UO_1438 (O_1438,N_6817,N_6117);
or UO_1439 (O_1439,N_5701,N_9028);
or UO_1440 (O_1440,N_8145,N_9303);
or UO_1441 (O_1441,N_6915,N_5064);
and UO_1442 (O_1442,N_8109,N_9764);
or UO_1443 (O_1443,N_8770,N_6772);
and UO_1444 (O_1444,N_5008,N_5648);
nor UO_1445 (O_1445,N_6330,N_7651);
nor UO_1446 (O_1446,N_6966,N_5188);
nand UO_1447 (O_1447,N_7128,N_5175);
or UO_1448 (O_1448,N_5042,N_5597);
and UO_1449 (O_1449,N_6665,N_5594);
and UO_1450 (O_1450,N_5571,N_7307);
nor UO_1451 (O_1451,N_6210,N_7978);
nor UO_1452 (O_1452,N_5647,N_6007);
nor UO_1453 (O_1453,N_9199,N_9388);
nand UO_1454 (O_1454,N_9732,N_9085);
or UO_1455 (O_1455,N_5220,N_6291);
xnor UO_1456 (O_1456,N_6786,N_8541);
and UO_1457 (O_1457,N_9023,N_5634);
nor UO_1458 (O_1458,N_5445,N_8045);
and UO_1459 (O_1459,N_7378,N_5830);
nand UO_1460 (O_1460,N_9273,N_8082);
nand UO_1461 (O_1461,N_9054,N_5528);
nand UO_1462 (O_1462,N_7439,N_9692);
nand UO_1463 (O_1463,N_8148,N_9919);
nand UO_1464 (O_1464,N_7269,N_8088);
and UO_1465 (O_1465,N_7958,N_7820);
nor UO_1466 (O_1466,N_9899,N_7388);
nand UO_1467 (O_1467,N_5407,N_9969);
or UO_1468 (O_1468,N_9947,N_7019);
nor UO_1469 (O_1469,N_7849,N_5211);
nand UO_1470 (O_1470,N_9036,N_5928);
and UO_1471 (O_1471,N_8749,N_5533);
nor UO_1472 (O_1472,N_9632,N_7629);
and UO_1473 (O_1473,N_6586,N_5524);
or UO_1474 (O_1474,N_5582,N_9910);
nand UO_1475 (O_1475,N_7790,N_6218);
or UO_1476 (O_1476,N_6607,N_8912);
nand UO_1477 (O_1477,N_9320,N_6780);
and UO_1478 (O_1478,N_7806,N_7936);
xor UO_1479 (O_1479,N_5903,N_7821);
or UO_1480 (O_1480,N_5417,N_6952);
nor UO_1481 (O_1481,N_6626,N_5748);
and UO_1482 (O_1482,N_9629,N_7434);
or UO_1483 (O_1483,N_6480,N_7078);
nand UO_1484 (O_1484,N_8630,N_7174);
nor UO_1485 (O_1485,N_6154,N_6305);
or UO_1486 (O_1486,N_5057,N_5326);
and UO_1487 (O_1487,N_9290,N_5484);
xor UO_1488 (O_1488,N_6289,N_5111);
and UO_1489 (O_1489,N_7016,N_5185);
or UO_1490 (O_1490,N_8847,N_7196);
xor UO_1491 (O_1491,N_5432,N_8692);
nor UO_1492 (O_1492,N_9498,N_6094);
nor UO_1493 (O_1493,N_9394,N_8450);
nand UO_1494 (O_1494,N_5239,N_6024);
nand UO_1495 (O_1495,N_6654,N_7013);
nand UO_1496 (O_1496,N_5779,N_7051);
or UO_1497 (O_1497,N_9551,N_7198);
and UO_1498 (O_1498,N_9613,N_8709);
nor UO_1499 (O_1499,N_9326,N_8431);
endmodule