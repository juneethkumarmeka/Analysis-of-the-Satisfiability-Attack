module basic_2000_20000_2500_5_levels_2xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_777,In_955);
or U1 (N_1,In_1453,In_1889);
nor U2 (N_2,In_721,In_175);
nor U3 (N_3,In_57,In_199);
nor U4 (N_4,In_569,In_130);
nand U5 (N_5,In_441,In_1136);
and U6 (N_6,In_36,In_773);
or U7 (N_7,In_1995,In_1823);
nor U8 (N_8,In_1618,In_1779);
or U9 (N_9,In_1123,In_1738);
nor U10 (N_10,In_1298,In_1725);
nor U11 (N_11,In_547,In_58);
or U12 (N_12,In_325,In_949);
or U13 (N_13,In_910,In_1603);
nand U14 (N_14,In_716,In_1800);
or U15 (N_15,In_782,In_585);
nor U16 (N_16,In_1953,In_1081);
nor U17 (N_17,In_1261,In_827);
nand U18 (N_18,In_735,In_848);
nand U19 (N_19,In_855,In_1534);
or U20 (N_20,In_1294,In_1866);
nor U21 (N_21,In_382,In_275);
xor U22 (N_22,In_820,In_1111);
nor U23 (N_23,In_1256,In_1267);
and U24 (N_24,In_1637,In_1323);
or U25 (N_25,In_1705,In_1499);
and U26 (N_26,In_295,In_362);
nand U27 (N_27,In_1372,In_675);
or U28 (N_28,In_1615,In_507);
and U29 (N_29,In_1406,In_231);
nand U30 (N_30,In_673,In_623);
nor U31 (N_31,In_1758,In_1042);
or U32 (N_32,In_845,In_925);
nand U33 (N_33,In_875,In_1908);
nor U34 (N_34,In_23,In_1963);
and U35 (N_35,In_1421,In_907);
or U36 (N_36,In_1225,In_1595);
or U37 (N_37,In_1007,In_884);
and U38 (N_38,In_1792,In_830);
nand U39 (N_39,In_681,In_1934);
or U40 (N_40,In_364,In_248);
nor U41 (N_41,In_1567,In_561);
and U42 (N_42,In_213,In_1229);
or U43 (N_43,In_13,In_1143);
and U44 (N_44,In_885,In_1681);
nor U45 (N_45,In_1396,In_720);
nand U46 (N_46,In_663,In_794);
and U47 (N_47,In_1329,In_968);
or U48 (N_48,In_1080,In_913);
nand U49 (N_49,In_430,In_383);
and U50 (N_50,In_1273,In_698);
nor U51 (N_51,In_128,In_400);
or U52 (N_52,In_262,In_263);
and U53 (N_53,In_1606,In_1194);
nand U54 (N_54,In_82,In_1177);
nor U55 (N_55,In_1634,In_1649);
nor U56 (N_56,In_1068,In_50);
nor U57 (N_57,In_435,In_35);
or U58 (N_58,In_149,In_1895);
or U59 (N_59,In_1633,In_385);
or U60 (N_60,In_305,In_991);
or U61 (N_61,In_388,In_985);
nor U62 (N_62,In_1680,In_683);
nor U63 (N_63,In_1485,In_351);
and U64 (N_64,In_1580,In_670);
and U65 (N_65,In_396,In_1419);
and U66 (N_66,In_78,In_1588);
or U67 (N_67,In_1905,In_967);
nand U68 (N_68,In_1884,In_1906);
and U69 (N_69,In_161,In_265);
nor U70 (N_70,In_1596,In_1556);
nand U71 (N_71,In_1974,In_473);
nor U72 (N_72,In_705,In_1520);
nand U73 (N_73,In_1980,In_646);
nand U74 (N_74,In_142,In_176);
nand U75 (N_75,In_422,In_272);
nor U76 (N_76,In_81,In_210);
and U77 (N_77,In_812,In_1602);
and U78 (N_78,In_702,In_1096);
or U79 (N_79,In_1890,In_1700);
or U80 (N_80,In_1002,In_1166);
nand U81 (N_81,In_1066,In_1063);
nor U82 (N_82,In_497,In_431);
nor U83 (N_83,In_981,In_866);
and U84 (N_84,In_625,In_338);
nand U85 (N_85,In_151,In_116);
and U86 (N_86,In_1959,In_1870);
or U87 (N_87,In_1090,In_674);
or U88 (N_88,In_22,In_1666);
and U89 (N_89,In_584,In_1528);
and U90 (N_90,In_371,In_1262);
or U91 (N_91,In_813,In_1429);
nand U92 (N_92,In_1939,In_559);
nor U93 (N_93,In_294,In_1147);
nand U94 (N_94,In_1028,In_1616);
nor U95 (N_95,In_887,In_434);
nor U96 (N_96,In_924,In_836);
nor U97 (N_97,In_776,In_168);
nand U98 (N_98,In_1020,In_998);
nand U99 (N_99,In_1644,In_620);
nand U100 (N_100,In_150,In_1762);
and U101 (N_101,In_1878,In_1537);
nor U102 (N_102,In_309,In_1141);
or U103 (N_103,In_1629,In_408);
nor U104 (N_104,In_243,In_562);
nor U105 (N_105,In_296,In_277);
nand U106 (N_106,In_297,In_300);
and U107 (N_107,In_958,In_1724);
nand U108 (N_108,In_1348,In_354);
nand U109 (N_109,In_983,In_1051);
nor U110 (N_110,In_1257,In_814);
and U111 (N_111,In_1260,In_235);
and U112 (N_112,In_1555,In_1290);
nor U113 (N_113,In_780,In_1611);
and U114 (N_114,In_1244,In_1103);
nand U115 (N_115,In_443,In_84);
and U116 (N_116,In_117,In_1067);
and U117 (N_117,In_21,In_1820);
nand U118 (N_118,In_344,In_1132);
nor U119 (N_119,In_1749,In_1830);
nand U120 (N_120,In_990,In_881);
nor U121 (N_121,In_1208,In_250);
nand U122 (N_122,In_1516,In_1607);
nor U123 (N_123,In_311,In_64);
nand U124 (N_124,In_221,In_1849);
or U125 (N_125,In_1539,In_1651);
or U126 (N_126,In_629,In_6);
nand U127 (N_127,In_1223,In_1914);
and U128 (N_128,In_1763,In_1947);
nor U129 (N_129,In_342,In_249);
and U130 (N_130,In_650,In_1397);
nand U131 (N_131,In_922,In_904);
or U132 (N_132,In_245,In_741);
and U133 (N_133,In_1722,In_1932);
and U134 (N_134,In_945,In_24);
and U135 (N_135,In_1249,In_1017);
nor U136 (N_136,In_988,In_589);
and U137 (N_137,In_603,In_452);
or U138 (N_138,In_186,In_831);
nor U139 (N_139,In_1466,In_1819);
and U140 (N_140,In_1853,In_1753);
or U141 (N_141,In_1886,In_548);
or U142 (N_142,In_1458,In_1272);
and U143 (N_143,In_1263,In_14);
nor U144 (N_144,In_519,In_736);
and U145 (N_145,In_1535,In_1672);
and U146 (N_146,In_1898,In_510);
and U147 (N_147,In_1719,In_264);
and U148 (N_148,In_1129,In_169);
nand U149 (N_149,In_1969,In_505);
nand U150 (N_150,In_1542,In_1807);
nor U151 (N_151,In_1321,In_1524);
or U152 (N_152,In_484,In_619);
and U153 (N_153,In_1243,In_902);
nand U154 (N_154,In_1676,In_1105);
nor U155 (N_155,In_405,In_1950);
and U156 (N_156,In_1716,In_506);
nor U157 (N_157,In_960,In_786);
and U158 (N_158,In_1825,In_1161);
nor U159 (N_159,In_200,In_899);
and U160 (N_160,In_1482,In_1824);
and U161 (N_161,In_1360,In_304);
nor U162 (N_162,In_1912,In_74);
xnor U163 (N_163,In_1752,In_326);
nand U164 (N_164,In_1018,In_676);
or U165 (N_165,In_1169,In_604);
nand U166 (N_166,In_274,In_428);
nand U167 (N_167,In_891,In_1434);
or U168 (N_168,In_1922,In_89);
nand U169 (N_169,In_1465,In_173);
and U170 (N_170,In_19,In_239);
nor U171 (N_171,In_1411,In_1487);
xor U172 (N_172,In_109,In_933);
nand U173 (N_173,In_826,In_1673);
or U174 (N_174,In_1305,In_1691);
nor U175 (N_175,In_999,In_1173);
nor U176 (N_176,In_1095,In_244);
nor U177 (N_177,In_1627,In_554);
or U178 (N_178,In_324,In_1811);
and U179 (N_179,In_425,In_482);
and U180 (N_180,In_1768,In_890);
or U181 (N_181,In_1423,In_1444);
or U182 (N_182,In_695,In_1435);
xnor U183 (N_183,In_691,In_1571);
nor U184 (N_184,In_872,In_1938);
nand U185 (N_185,In_1944,In_302);
nor U186 (N_186,In_1788,In_1314);
or U187 (N_187,In_1843,In_1238);
nand U188 (N_188,In_1250,In_996);
or U189 (N_189,In_724,In_68);
or U190 (N_190,In_76,In_88);
and U191 (N_191,In_215,In_1858);
nand U192 (N_192,In_1986,In_146);
nor U193 (N_193,In_1341,In_410);
and U194 (N_194,In_1892,In_1041);
nor U195 (N_195,In_556,In_26);
nor U196 (N_196,In_133,In_573);
or U197 (N_197,In_957,In_1258);
and U198 (N_198,In_281,In_163);
nand U199 (N_199,In_1058,In_419);
or U200 (N_200,In_271,In_1027);
nor U201 (N_201,In_1484,In_464);
nand U202 (N_202,In_1349,In_1550);
nor U203 (N_203,In_658,In_1899);
and U204 (N_204,In_1613,In_240);
nand U205 (N_205,In_889,In_1204);
or U206 (N_206,In_1188,In_463);
or U207 (N_207,In_1685,In_591);
or U208 (N_208,In_930,In_1038);
nor U209 (N_209,In_1001,In_105);
nor U210 (N_210,In_896,In_1504);
nand U211 (N_211,In_457,In_1960);
nor U212 (N_212,In_1717,In_1525);
and U213 (N_213,In_1809,In_938);
nor U214 (N_214,In_125,In_1052);
xnor U215 (N_215,In_706,In_112);
nand U216 (N_216,In_1433,In_1375);
and U217 (N_217,In_27,In_1463);
nand U218 (N_218,In_745,In_113);
nand U219 (N_219,In_1108,In_1390);
nand U220 (N_220,In_5,In_404);
nor U221 (N_221,In_937,In_427);
or U222 (N_222,In_723,In_1994);
or U223 (N_223,In_501,In_164);
or U224 (N_224,In_530,In_67);
and U225 (N_225,In_480,In_1954);
nand U226 (N_226,In_1106,In_232);
or U227 (N_227,In_600,In_508);
nor U228 (N_228,In_766,In_550);
nor U229 (N_229,In_71,In_893);
and U230 (N_230,In_16,In_1239);
and U231 (N_231,In_1847,In_1657);
xnor U232 (N_232,In_1765,In_678);
or U233 (N_233,In_883,In_331);
xnor U234 (N_234,In_299,In_1200);
nor U235 (N_235,In_1478,In_1473);
and U236 (N_236,In_1073,In_1569);
nor U237 (N_237,In_0,In_197);
and U238 (N_238,In_1791,In_1436);
nand U239 (N_239,In_1134,In_1382);
xnor U240 (N_240,In_1359,In_1587);
xnor U241 (N_241,In_1923,In_178);
nor U242 (N_242,In_734,In_1842);
nand U243 (N_243,In_788,In_1982);
nand U244 (N_244,In_1011,In_1481);
and U245 (N_245,In_1455,In_316);
nand U246 (N_246,In_1101,In_486);
and U247 (N_247,In_399,In_1220);
nand U248 (N_248,In_1165,In_1167);
nor U249 (N_249,In_1156,In_1623);
and U250 (N_250,In_390,In_516);
xnor U251 (N_251,In_62,In_1075);
nor U252 (N_252,In_1089,In_1352);
xnor U253 (N_253,In_1226,In_312);
nor U254 (N_254,In_1748,In_900);
and U255 (N_255,In_962,In_1171);
or U256 (N_256,In_632,In_141);
and U257 (N_257,In_690,In_1818);
xnor U258 (N_258,In_701,In_1428);
nand U259 (N_259,In_477,In_824);
or U260 (N_260,In_606,In_225);
or U261 (N_261,In_1110,In_1816);
nor U262 (N_262,In_858,In_1495);
nor U263 (N_263,In_223,In_760);
nor U264 (N_264,In_1767,In_1834);
nand U265 (N_265,In_1216,In_122);
nand U266 (N_266,In_1883,In_158);
nor U267 (N_267,In_120,In_461);
or U268 (N_268,In_1660,In_1076);
or U269 (N_269,In_1150,In_1964);
xnor U270 (N_270,In_1726,In_266);
or U271 (N_271,In_187,In_709);
or U272 (N_272,In_1911,In_227);
nor U273 (N_273,In_520,In_1989);
and U274 (N_274,In_1308,In_1064);
or U275 (N_275,In_1747,In_972);
nor U276 (N_276,In_1777,In_1370);
or U277 (N_277,In_1078,In_288);
and U278 (N_278,In_1729,In_7);
and U279 (N_279,In_1284,In_194);
nor U280 (N_280,In_1707,In_1756);
or U281 (N_281,In_1012,In_1692);
or U282 (N_282,In_1868,In_179);
and U283 (N_283,In_689,In_144);
nand U284 (N_284,In_540,In_861);
and U285 (N_285,In_898,In_1712);
nor U286 (N_286,In_166,In_363);
nor U287 (N_287,In_409,In_961);
nand U288 (N_288,In_882,In_353);
nor U289 (N_289,In_1826,In_236);
or U290 (N_290,In_995,In_1355);
or U291 (N_291,In_1835,In_1683);
nor U292 (N_292,In_1293,In_1773);
xnor U293 (N_293,In_515,In_329);
and U294 (N_294,In_1678,In_1715);
or U295 (N_295,In_54,In_340);
and U296 (N_296,In_1965,In_1268);
nor U297 (N_297,In_1379,In_20);
or U298 (N_298,In_1813,In_1449);
or U299 (N_299,In_1316,In_611);
and U300 (N_300,In_320,In_1193);
nor U301 (N_301,In_769,In_1745);
and U302 (N_302,In_842,In_40);
and U303 (N_303,In_1209,In_1266);
and U304 (N_304,In_638,In_586);
nor U305 (N_305,In_1186,In_686);
nor U306 (N_306,In_1276,In_1281);
or U307 (N_307,In_914,In_1462);
and U308 (N_308,In_1903,In_729);
or U309 (N_309,In_867,In_1292);
or U310 (N_310,In_819,In_526);
and U311 (N_311,In_451,In_1227);
or U312 (N_312,In_1415,In_1711);
and U313 (N_313,In_986,In_246);
and U314 (N_314,In_588,In_982);
nand U315 (N_315,In_1560,In_217);
and U316 (N_316,In_1536,In_29);
and U317 (N_317,In_1056,In_1850);
and U318 (N_318,In_37,In_1373);
nand U319 (N_319,In_1006,In_313);
nor U320 (N_320,In_289,In_1205);
nand U321 (N_321,In_1184,In_209);
and U322 (N_322,In_1653,In_1740);
nand U323 (N_323,In_643,In_483);
and U324 (N_324,In_607,In_966);
or U325 (N_325,In_555,In_644);
or U326 (N_326,In_870,In_1398);
or U327 (N_327,In_1581,In_1941);
nand U328 (N_328,In_1174,In_226);
or U329 (N_329,In_596,In_471);
nand U330 (N_330,In_32,In_1840);
nand U331 (N_331,In_139,In_123);
nand U332 (N_332,In_971,In_1918);
nor U333 (N_333,In_1638,In_1195);
nand U334 (N_334,In_825,In_1310);
nand U335 (N_335,In_1985,In_915);
nor U336 (N_336,In_1322,In_1432);
nor U337 (N_337,In_1307,In_370);
nor U338 (N_338,In_1945,In_462);
nor U339 (N_339,In_93,In_946);
and U340 (N_340,In_1927,In_1511);
nor U341 (N_341,In_669,In_534);
or U342 (N_342,In_389,In_1997);
or U343 (N_343,In_1446,In_1877);
or U344 (N_344,In_974,In_594);
or U345 (N_345,In_374,In_1399);
nor U346 (N_346,In_43,In_1741);
xor U347 (N_347,In_1920,In_710);
nand U348 (N_348,In_541,In_1781);
and U349 (N_349,In_579,In_1231);
nand U350 (N_350,In_159,In_1697);
or U351 (N_351,In_613,In_733);
nor U352 (N_352,In_73,In_298);
xnor U353 (N_353,In_648,In_1380);
nor U354 (N_354,In_699,In_1330);
and U355 (N_355,In_1553,In_513);
or U356 (N_356,In_257,In_1916);
nand U357 (N_357,In_259,In_1418);
nand U358 (N_358,In_1326,In_1682);
or U359 (N_359,In_106,In_1211);
or U360 (N_360,In_959,In_1130);
and U361 (N_361,In_228,In_1590);
nand U362 (N_362,In_864,In_684);
nand U363 (N_363,In_795,In_174);
and U364 (N_364,In_254,In_1778);
xnor U365 (N_365,In_1659,In_1494);
or U366 (N_366,In_285,In_1531);
nand U367 (N_367,In_590,In_897);
nand U368 (N_368,In_509,In_1545);
or U369 (N_369,In_916,In_494);
or U370 (N_370,In_479,In_1861);
xor U371 (N_371,In_1182,In_1829);
or U372 (N_372,In_291,In_124);
or U373 (N_373,In_56,In_377);
or U374 (N_374,In_546,In_1732);
or U375 (N_375,In_1139,In_1601);
nand U376 (N_376,In_1277,In_335);
or U377 (N_377,In_1236,In_1029);
and U378 (N_378,In_627,In_977);
nand U379 (N_379,In_207,In_1568);
nor U380 (N_380,In_1207,In_1702);
and U381 (N_381,In_1190,In_70);
nand U382 (N_382,In_1530,In_1955);
and U383 (N_383,In_1241,In_328);
nor U384 (N_384,In_1085,In_160);
nor U385 (N_385,In_1967,In_614);
xor U386 (N_386,In_876,In_52);
or U387 (N_387,In_1839,In_1951);
or U388 (N_388,In_1782,In_514);
or U389 (N_389,In_1652,In_948);
or U390 (N_390,In_1915,In_170);
nand U391 (N_391,In_189,In_844);
xnor U392 (N_392,In_1137,In_1039);
nor U393 (N_393,In_815,In_1586);
nor U394 (N_394,In_1785,In_99);
nor U395 (N_395,In_1460,In_1838);
nand U396 (N_396,In_652,In_1698);
nand U397 (N_397,In_1658,In_181);
and U398 (N_398,In_1030,In_1592);
nand U399 (N_399,In_1439,In_80);
or U400 (N_400,In_1224,In_597);
and U401 (N_401,In_1519,In_905);
nor U402 (N_402,In_1046,In_1936);
or U403 (N_403,In_1252,In_829);
or U404 (N_404,In_1483,In_1114);
nor U405 (N_405,In_970,In_1353);
nor U406 (N_406,In_963,In_94);
nor U407 (N_407,In_475,In_439);
nor U408 (N_408,In_535,In_557);
nand U409 (N_409,In_414,In_1972);
nor U410 (N_410,In_1138,In_1479);
nand U411 (N_411,In_49,In_1891);
or U412 (N_412,In_352,In_1461);
nand U413 (N_413,In_989,In_1392);
or U414 (N_414,In_1160,In_177);
or U415 (N_415,In_637,In_853);
and U416 (N_416,In_1971,In_687);
and U417 (N_417,In_1251,In_145);
or U418 (N_418,In_1509,In_440);
nand U419 (N_419,In_1021,In_315);
nor U420 (N_420,In_233,In_206);
and U421 (N_421,In_1427,In_1100);
and U422 (N_422,In_379,In_1407);
nor U423 (N_423,In_599,In_1597);
and U424 (N_424,In_3,In_247);
or U425 (N_425,In_196,In_1476);
nor U426 (N_426,In_1532,In_86);
nor U427 (N_427,In_1467,In_528);
nor U428 (N_428,In_1146,In_994);
nand U429 (N_429,In_1507,In_919);
nor U430 (N_430,In_656,In_241);
or U431 (N_431,In_1025,In_1946);
nand U432 (N_432,In_577,In_1036);
or U433 (N_433,In_1774,In_69);
nand U434 (N_434,In_47,In_762);
nand U435 (N_435,In_1797,In_877);
and U436 (N_436,In_1966,In_1424);
nand U437 (N_437,In_358,In_224);
nand U438 (N_438,In_807,In_704);
nand U439 (N_439,In_1845,In_672);
nand U440 (N_440,In_1062,In_1014);
nor U441 (N_441,In_242,In_322);
or U442 (N_442,In_1640,In_1733);
nor U443 (N_443,In_975,In_1264);
or U444 (N_444,In_666,In_744);
and U445 (N_445,In_1522,In_1975);
or U446 (N_446,In_1232,In_1503);
nand U447 (N_447,In_135,In_253);
and U448 (N_448,In_268,In_1632);
and U449 (N_449,In_1585,In_886);
nand U450 (N_450,In_15,In_238);
or U451 (N_451,In_759,In_1343);
and U452 (N_452,In_799,In_334);
xnor U453 (N_453,In_485,In_442);
or U454 (N_454,In_849,In_466);
nand U455 (N_455,In_660,In_775);
nor U456 (N_456,In_1621,In_350);
and U457 (N_457,In_51,In_1488);
and U458 (N_458,In_155,In_1514);
nand U459 (N_459,In_127,In_1148);
or U460 (N_460,In_1422,In_517);
and U461 (N_461,In_863,In_46);
nor U462 (N_462,In_1686,In_722);
and U463 (N_463,In_951,In_467);
xor U464 (N_464,In_1269,In_802);
nand U465 (N_465,In_1367,In_1408);
nand U466 (N_466,In_659,In_1766);
nor U467 (N_467,In_1365,In_1901);
and U468 (N_468,In_1882,In_458);
nand U469 (N_469,In_1948,In_688);
or U470 (N_470,In_1356,In_1988);
nand U471 (N_471,In_626,In_406);
xnor U472 (N_472,In_1979,In_993);
nor U473 (N_473,In_1196,In_391);
or U474 (N_474,In_365,In_1486);
nand U475 (N_475,In_1925,In_1197);
nand U476 (N_476,In_1924,In_188);
nand U477 (N_477,In_1142,In_368);
or U478 (N_478,In_1286,In_1783);
and U479 (N_479,In_1704,In_703);
and U480 (N_480,In_793,In_1684);
nor U481 (N_481,In_1098,In_1761);
or U482 (N_482,In_1862,In_39);
and U483 (N_483,In_1278,In_1222);
or U484 (N_484,In_512,In_1902);
and U485 (N_485,In_838,In_908);
and U486 (N_486,In_767,In_470);
or U487 (N_487,In_167,In_888);
or U488 (N_488,In_798,In_746);
nand U489 (N_489,In_1546,In_1589);
nand U490 (N_490,In_1764,In_1949);
and U491 (N_491,In_1500,In_1117);
nor U492 (N_492,In_1646,In_1426);
nand U493 (N_493,In_53,In_859);
nor U494 (N_494,In_911,In_575);
nor U495 (N_495,In_153,In_822);
nor U496 (N_496,In_1641,In_260);
xor U497 (N_497,In_48,In_1931);
nor U498 (N_498,In_1780,In_1475);
nor U499 (N_499,In_347,In_55);
or U500 (N_500,In_621,In_96);
and U501 (N_501,In_634,In_137);
and U502 (N_502,In_18,In_1852);
nand U503 (N_503,In_1430,In_1448);
nor U504 (N_504,In_1794,In_865);
nand U505 (N_505,In_1445,In_172);
or U506 (N_506,In_1389,In_307);
nand U507 (N_507,In_1645,In_796);
nand U508 (N_508,In_1827,In_765);
and U509 (N_509,In_719,In_1315);
nor U510 (N_510,In_1312,In_1416);
and U511 (N_511,In_1973,In_857);
and U512 (N_512,In_1489,In_372);
nand U513 (N_513,In_1234,In_1024);
nand U514 (N_514,In_923,In_339);
xor U515 (N_515,In_1480,In_456);
nand U516 (N_516,In_929,In_1612);
xor U517 (N_517,In_214,In_1559);
nand U518 (N_518,In_1282,In_693);
or U519 (N_519,In_1055,In_789);
and U520 (N_520,In_1378,In_1346);
nor U521 (N_521,In_1736,In_1320);
nand U522 (N_522,In_395,In_1342);
or U523 (N_523,In_792,In_1318);
or U524 (N_524,In_956,In_1071);
and U525 (N_525,In_1087,In_1815);
nand U526 (N_526,In_1677,In_1812);
nand U527 (N_527,In_921,In_503);
nand U528 (N_528,In_661,In_101);
nand U529 (N_529,In_1468,In_59);
nor U530 (N_530,In_944,In_308);
nand U531 (N_531,In_1984,In_801);
and U532 (N_532,In_1998,In_1447);
nor U533 (N_533,In_1414,In_1957);
xor U534 (N_534,In_1162,In_1910);
or U535 (N_535,In_258,In_1218);
or U536 (N_536,In_732,In_803);
nand U537 (N_537,In_498,In_1841);
nor U538 (N_538,In_492,In_1620);
nor U539 (N_539,In_1010,In_208);
nand U540 (N_540,In_751,In_1708);
nor U541 (N_541,In_1793,In_653);
or U542 (N_542,In_1880,In_1942);
or U543 (N_543,In_1650,In_539);
nor U544 (N_544,In_1699,In_805);
nor U545 (N_545,In_360,In_523);
nand U546 (N_546,In_193,In_1893);
or U547 (N_547,In_1319,In_757);
and U548 (N_548,In_1325,In_895);
nand U549 (N_549,In_755,In_455);
nand U550 (N_550,In_785,In_343);
nor U551 (N_551,In_1187,In_34);
nand U552 (N_552,In_500,In_79);
or U553 (N_553,In_1848,In_1317);
nor U554 (N_554,In_715,In_753);
nand U555 (N_555,In_1887,In_287);
nor U556 (N_556,In_1690,In_1155);
xnor U557 (N_557,In_1019,In_1057);
xor U558 (N_558,In_918,In_1576);
nand U559 (N_559,In_1212,In_839);
nor U560 (N_560,In_1737,In_1296);
nand U561 (N_561,In_1863,In_1082);
and U562 (N_562,In_1470,In_44);
or U563 (N_563,In_1119,In_1404);
nand U564 (N_564,In_1798,In_587);
nor U565 (N_565,In_1578,In_685);
nand U566 (N_566,In_1145,In_1151);
and U567 (N_567,In_184,In_1654);
and U568 (N_568,In_469,In_1179);
and U569 (N_569,In_415,In_367);
nor U570 (N_570,In_566,In_1092);
nand U571 (N_571,In_380,In_711);
nor U572 (N_572,In_1043,In_1154);
and U573 (N_573,In_423,In_1127);
nor U574 (N_574,In_204,In_1345);
or U575 (N_575,In_115,In_1832);
or U576 (N_576,In_714,In_1735);
and U577 (N_577,In_327,In_1395);
nand U578 (N_578,In_303,In_1237);
nor U579 (N_579,In_728,In_103);
or U580 (N_580,In_1851,In_381);
or U581 (N_581,In_1566,In_1992);
nor U582 (N_582,In_1583,In_85);
or U583 (N_583,In_903,In_1605);
xnor U584 (N_584,In_1185,In_1926);
or U585 (N_585,In_928,In_1490);
and U586 (N_586,In_293,In_943);
nor U587 (N_587,In_828,In_1561);
nand U588 (N_588,In_880,In_979);
xnor U589 (N_589,In_532,In_529);
and U590 (N_590,In_1958,In_1501);
nor U591 (N_591,In_846,In_121);
xor U592 (N_592,In_191,In_1405);
and U593 (N_593,In_436,In_1180);
nand U594 (N_594,In_1221,In_1450);
and U595 (N_595,In_764,In_333);
or U596 (N_596,In_195,In_1459);
nor U597 (N_597,In_1037,In_1689);
or U598 (N_598,In_927,In_770);
nand U599 (N_599,In_290,In_1135);
nand U600 (N_600,In_1687,In_126);
nand U601 (N_601,In_9,In_1192);
or U602 (N_602,In_108,In_978);
or U603 (N_603,In_493,In_1254);
nor U604 (N_604,In_602,In_1598);
nand U605 (N_605,In_487,In_1584);
or U606 (N_606,In_1437,In_1900);
or U607 (N_607,In_1574,In_1149);
or U608 (N_608,In_657,In_1593);
nand U609 (N_609,In_1909,In_1876);
nand U610 (N_610,In_306,In_279);
nor U611 (N_611,In_1970,In_1077);
and U612 (N_612,In_574,In_616);
and U613 (N_613,In_750,In_1175);
and U614 (N_614,In_592,In_1730);
and U615 (N_615,In_1181,In_1981);
and U616 (N_616,In_1497,In_1);
nor U617 (N_617,In_496,In_878);
and U618 (N_618,In_1344,In_448);
and U619 (N_619,In_459,In_1440);
nand U620 (N_620,In_1074,In_393);
or U621 (N_621,In_1000,In_1183);
nand U622 (N_622,In_1913,In_1990);
nand U623 (N_623,In_1259,In_1210);
nor U624 (N_624,In_1930,In_1701);
nand U625 (N_625,In_154,In_1859);
nand U626 (N_626,In_533,In_1401);
and U627 (N_627,In_1639,In_635);
nand U628 (N_628,In_1993,In_1608);
nand U629 (N_629,In_1943,In_33);
nand U630 (N_630,In_739,In_576);
nor U631 (N_631,In_1512,In_1088);
nand U632 (N_632,In_1956,In_1128);
or U633 (N_633,In_747,In_230);
nor U634 (N_634,In_346,In_1873);
or U635 (N_635,In_1803,In_527);
nor U636 (N_636,In_873,In_114);
or U637 (N_637,In_816,In_931);
or U638 (N_638,In_628,In_1350);
and U639 (N_639,In_1983,In_781);
and U640 (N_640,In_1376,In_373);
and U641 (N_641,In_447,In_1443);
nand U642 (N_642,In_942,In_162);
nor U643 (N_643,In_1810,In_823);
nor U644 (N_644,In_833,In_355);
or U645 (N_645,In_356,In_679);
and U646 (N_646,In_1015,In_1072);
or U647 (N_647,In_1364,In_1648);
nand U648 (N_648,In_1888,In_1517);
nand U649 (N_649,In_1248,In_939);
nor U650 (N_650,In_568,In_840);
nor U651 (N_651,In_1804,In_1802);
or U652 (N_652,In_336,In_438);
nand U653 (N_653,In_595,In_251);
and U654 (N_654,In_1746,In_992);
or U655 (N_655,In_394,In_1358);
or U656 (N_656,In_1049,In_261);
nor U657 (N_657,In_636,In_787);
and U658 (N_658,In_671,In_1496);
nand U659 (N_659,In_1004,In_1933);
or U660 (N_660,In_1340,In_1005);
nor U661 (N_661,In_1591,In_1253);
or U662 (N_662,In_718,In_330);
nor U663 (N_663,In_936,In_98);
or U664 (N_664,In_854,In_947);
or U665 (N_665,In_1026,In_1628);
nor U666 (N_666,In_950,In_713);
nor U667 (N_667,In_45,In_129);
and U668 (N_668,In_1053,In_642);
nand U669 (N_669,In_912,In_1255);
and U670 (N_670,In_1871,In_1083);
nor U671 (N_671,In_645,In_1362);
or U672 (N_672,In_1731,In_1189);
and U673 (N_673,In_633,In_1377);
nand U674 (N_674,In_1045,In_219);
nand U675 (N_675,In_1710,In_1163);
nand U676 (N_676,In_797,In_1033);
nand U677 (N_677,In_1786,In_772);
or U678 (N_678,In_495,In_1662);
and U679 (N_679,In_1327,In_1144);
or U680 (N_680,In_286,In_630);
nor U681 (N_681,In_1297,In_1022);
xnor U682 (N_682,In_1723,In_521);
nor U683 (N_683,In_1991,In_560);
xnor U684 (N_684,In_1454,In_1178);
nand U685 (N_685,In_1604,In_1201);
and U686 (N_686,In_570,In_1573);
or U687 (N_687,In_601,In_1552);
and U688 (N_688,In_1968,In_267);
or U689 (N_689,In_1742,In_1540);
and U690 (N_690,In_1527,In_229);
or U691 (N_691,In_1790,In_522);
and U692 (N_692,In_1881,In_1523);
nand U693 (N_693,In_1642,In_1122);
nor U694 (N_694,In_183,In_1675);
nand U695 (N_695,In_332,In_397);
nor U696 (N_696,In_1713,In_1755);
and U697 (N_697,In_1113,In_774);
nor U698 (N_698,In_1721,In_707);
nor U699 (N_699,In_138,In_1577);
or U700 (N_700,In_1668,In_818);
nor U701 (N_701,In_1565,In_624);
nand U702 (N_702,In_8,In_378);
nand U703 (N_703,In_148,In_847);
nand U704 (N_704,In_1548,In_92);
nand U705 (N_705,In_450,In_835);
nor U706 (N_706,In_77,In_749);
nor U707 (N_707,In_474,In_662);
nor U708 (N_708,In_1291,In_276);
nand U709 (N_709,In_564,In_1003);
xnor U710 (N_710,In_453,In_1775);
nor U711 (N_711,In_1363,In_544);
and U712 (N_712,In_622,In_1357);
nor U713 (N_713,In_449,In_143);
and U714 (N_714,In_869,In_1614);
nor U715 (N_715,In_165,In_270);
or U716 (N_716,In_1158,In_1643);
nand U717 (N_717,In_700,In_1309);
and U718 (N_718,In_1044,In_1714);
and U719 (N_719,In_909,In_768);
or U720 (N_720,In_1728,In_612);
nor U721 (N_721,In_901,In_100);
or U722 (N_722,In_817,In_856);
and U723 (N_723,In_1069,In_1720);
or U724 (N_724,In_1896,In_537);
nor U725 (N_725,In_1772,In_1228);
and U726 (N_726,In_1337,In_1301);
nor U727 (N_727,In_1831,In_1844);
nor U728 (N_728,In_654,In_1594);
nor U729 (N_729,In_580,In_87);
and U730 (N_730,In_1563,In_1787);
nand U731 (N_731,In_1050,In_376);
nor U732 (N_732,In_1904,In_1086);
or U733 (N_733,In_1609,In_1381);
and U734 (N_734,In_369,In_1008);
xnor U735 (N_735,In_1805,In_1394);
and U736 (N_736,In_1289,In_1333);
nand U737 (N_737,In_392,In_578);
and U738 (N_738,In_319,In_476);
or U739 (N_739,In_361,In_743);
or U740 (N_740,In_1894,In_1492);
or U741 (N_741,In_1784,In_1391);
nor U742 (N_742,In_1864,In_610);
or U743 (N_743,In_28,In_926);
nor U744 (N_744,In_843,In_218);
or U745 (N_745,In_871,In_545);
nand U746 (N_746,In_821,In_1734);
or U747 (N_747,In_433,In_572);
nor U748 (N_748,In_1288,In_110);
nand U749 (N_749,In_416,In_756);
nor U750 (N_750,In_491,In_1464);
nor U751 (N_751,In_91,In_941);
nand U752 (N_752,In_424,In_668);
nor U753 (N_753,In_549,In_1176);
and U754 (N_754,In_1107,In_726);
nor U755 (N_755,In_386,In_1600);
and U756 (N_756,In_402,In_1287);
nand U757 (N_757,In_969,In_1799);
nand U758 (N_758,In_278,In_1457);
nand U759 (N_759,In_1907,In_1679);
nand U760 (N_760,In_1295,In_468);
or U761 (N_761,In_1855,In_1328);
or U762 (N_762,In_631,In_667);
nand U763 (N_763,In_1191,In_111);
nor U764 (N_764,In_1121,In_1091);
nor U765 (N_765,In_1199,In_1383);
and U766 (N_766,In_102,In_1562);
or U767 (N_767,In_784,In_1635);
and U768 (N_768,In_976,In_234);
nor U769 (N_769,In_1230,In_1203);
and U770 (N_770,In_1854,In_1727);
nor U771 (N_771,In_60,In_1354);
or U772 (N_772,In_403,In_1403);
nor U773 (N_773,In_964,In_1213);
nor U774 (N_774,In_1366,In_1084);
or U775 (N_775,In_1978,In_708);
nor U776 (N_776,In_314,In_934);
and U777 (N_777,In_478,In_1505);
or U778 (N_778,In_778,In_359);
and U779 (N_779,In_737,In_1977);
or U780 (N_780,In_1198,In_680);
or U781 (N_781,In_738,In_1023);
or U782 (N_782,In_1233,In_252);
nor U783 (N_783,In_1808,In_63);
and U784 (N_784,In_203,In_1079);
or U785 (N_785,In_1451,In_808);
or U786 (N_786,In_1099,In_617);
and U787 (N_787,In_932,In_1617);
and U788 (N_788,In_1929,In_41);
nand U789 (N_789,In_1324,In_997);
nor U790 (N_790,In_1125,In_499);
and U791 (N_791,In_1789,In_502);
and U792 (N_792,In_292,In_1054);
nand U793 (N_793,In_1265,In_134);
nor U794 (N_794,In_1558,In_1335);
nand U795 (N_795,In_1219,In_201);
nor U796 (N_796,In_851,In_345);
or U797 (N_797,In_1417,In_1770);
and U798 (N_798,In_1557,In_525);
and U799 (N_799,In_75,In_273);
and U800 (N_800,In_375,In_581);
or U801 (N_801,In_1070,In_1371);
nor U802 (N_802,In_1526,In_190);
nand U803 (N_803,In_1270,In_1118);
nor U804 (N_804,In_1669,In_1060);
and U805 (N_805,In_140,In_563);
nand U806 (N_806,In_131,In_1471);
or U807 (N_807,In_1857,In_1695);
and U808 (N_808,In_542,In_1283);
and U809 (N_809,In_1009,In_1664);
nand U810 (N_810,In_12,In_558);
and U811 (N_811,In_1332,In_284);
or U812 (N_812,In_790,In_1300);
and U813 (N_813,In_465,In_1303);
nand U814 (N_814,In_1247,In_655);
and U815 (N_815,In_104,In_1215);
nand U816 (N_816,In_543,In_640);
or U817 (N_817,In_1164,In_1102);
nand U818 (N_818,In_283,In_868);
or U819 (N_819,In_834,In_879);
or U820 (N_820,In_748,In_538);
or U821 (N_821,In_198,In_1413);
nor U822 (N_822,In_1874,In_740);
nor U823 (N_823,In_860,In_65);
and U824 (N_824,In_1275,In_804);
nand U825 (N_825,In_1409,In_321);
or U826 (N_826,In_1919,In_30);
and U827 (N_827,In_1334,In_417);
or U828 (N_828,In_730,In_1280);
nor U829 (N_829,In_758,In_1630);
or U830 (N_830,In_212,In_454);
nand U831 (N_831,In_1104,In_437);
or U832 (N_832,In_1172,In_1048);
and U833 (N_833,In_696,In_301);
and U834 (N_834,In_1474,In_1491);
or U835 (N_835,In_1456,In_1061);
or U836 (N_836,In_1837,In_1709);
and U837 (N_837,In_171,In_717);
nor U838 (N_838,In_1533,In_973);
nor U839 (N_839,In_862,In_1647);
nor U840 (N_840,In_1477,In_984);
and U841 (N_841,In_1665,In_1743);
or U842 (N_842,In_504,In_429);
and U843 (N_843,In_1441,In_1109);
or U844 (N_844,In_800,In_1879);
and U845 (N_845,In_1510,In_1836);
nor U846 (N_846,In_1351,In_1897);
or U847 (N_847,In_665,In_1744);
or U848 (N_848,In_1760,In_421);
nand U849 (N_849,In_1452,In_1031);
or U850 (N_850,In_1159,In_387);
nor U851 (N_851,In_1631,In_72);
nand U852 (N_852,In_1544,In_180);
and U853 (N_853,In_1636,In_1610);
or U854 (N_854,In_742,In_1674);
nand U855 (N_855,In_1361,In_446);
and U856 (N_856,In_1387,In_1469);
or U857 (N_857,In_1754,In_1170);
nand U858 (N_858,In_1339,In_524);
nor U859 (N_859,In_892,In_1402);
nor U860 (N_860,In_1521,In_445);
or U861 (N_861,In_1311,In_1869);
nand U862 (N_862,In_1575,In_31);
and U863 (N_863,In_1885,In_472);
nor U864 (N_864,In_980,In_953);
nand U865 (N_865,In_1667,In_1425);
nand U866 (N_866,In_809,In_1817);
or U867 (N_867,In_1828,In_488);
and U868 (N_868,In_754,In_1420);
nor U869 (N_869,In_205,In_1937);
and U870 (N_870,In_1821,In_152);
or U871 (N_871,In_1554,In_97);
nand U872 (N_872,In_1299,In_987);
and U873 (N_873,In_837,In_553);
nor U874 (N_874,In_1140,In_1622);
and U875 (N_875,In_411,In_1624);
or U876 (N_876,In_682,In_783);
and U877 (N_877,In_1168,In_401);
and U878 (N_878,In_185,In_25);
nor U879 (N_879,In_95,In_318);
and U880 (N_880,In_1384,In_202);
or U881 (N_881,In_357,In_1035);
nand U882 (N_882,In_489,In_906);
nand U883 (N_883,In_582,In_639);
and U884 (N_884,In_1718,In_841);
nand U885 (N_885,In_583,In_220);
nand U886 (N_886,In_1769,In_1214);
nor U887 (N_887,In_712,In_806);
nand U888 (N_888,In_1133,In_1860);
and U889 (N_889,In_1619,In_1153);
or U890 (N_890,In_608,In_677);
and U891 (N_891,In_1115,In_1431);
or U892 (N_892,In_567,In_1386);
nor U893 (N_893,In_1917,In_1506);
or U894 (N_894,In_1338,In_1961);
nor U895 (N_895,In_147,In_1549);
and U896 (N_896,In_83,In_1245);
nand U897 (N_897,In_1120,In_1996);
nor U898 (N_898,In_565,In_1385);
nand U899 (N_899,In_647,In_384);
and U900 (N_900,In_651,In_697);
nand U901 (N_901,In_1776,In_1541);
and U902 (N_902,In_1625,In_1157);
or U903 (N_903,In_1759,In_1663);
and U904 (N_904,In_366,In_418);
nand U905 (N_905,In_1040,In_1438);
and U906 (N_906,In_256,In_1570);
and U907 (N_907,In_10,In_1152);
or U908 (N_908,In_107,In_965);
or U909 (N_909,In_763,In_1116);
nor U910 (N_910,In_1757,In_810);
or U911 (N_911,In_952,In_337);
nor U912 (N_912,In_1313,In_920);
and U913 (N_913,In_1626,In_1302);
or U914 (N_914,In_1388,In_157);
nor U915 (N_915,In_407,In_90);
xnor U916 (N_916,In_1962,In_1703);
and U917 (N_917,In_649,In_1306);
nand U918 (N_918,In_1529,In_255);
and U919 (N_919,In_1240,In_42);
and U920 (N_920,In_1833,In_1279);
nand U921 (N_921,In_1935,In_1875);
and U922 (N_922,In_692,In_1661);
or U923 (N_923,In_1059,In_11);
nor U924 (N_924,In_349,In_593);
or U925 (N_925,In_280,In_1750);
and U926 (N_926,In_317,In_1706);
or U927 (N_927,In_1543,In_598);
and U928 (N_928,In_731,In_1034);
nand U929 (N_929,In_132,In_481);
nand U930 (N_930,In_1112,In_694);
nor U931 (N_931,In_1515,In_1551);
nor U932 (N_932,In_874,In_894);
or U933 (N_933,In_531,In_460);
or U934 (N_934,In_211,In_1393);
or U935 (N_935,In_1806,In_1865);
nor U936 (N_936,In_1124,In_1579);
and U937 (N_937,In_1513,In_310);
and U938 (N_938,In_1940,In_1771);
nand U939 (N_939,In_1285,In_1928);
nand U940 (N_940,In_811,In_511);
nand U941 (N_941,In_282,In_1976);
or U942 (N_942,In_1671,In_1582);
and U943 (N_943,In_518,In_1921);
nand U944 (N_944,In_426,In_1412);
nor U945 (N_945,In_1369,In_1271);
and U946 (N_946,In_1822,In_1599);
and U947 (N_947,In_413,In_237);
and U948 (N_948,In_1987,In_1242);
or U949 (N_949,In_4,In_341);
nand U950 (N_950,In_1126,In_771);
nor U951 (N_951,In_727,In_1795);
or U952 (N_952,In_1472,In_192);
nor U953 (N_953,In_348,In_1093);
and U954 (N_954,In_1814,In_935);
xor U955 (N_955,In_1751,In_1999);
nor U956 (N_956,In_1336,In_850);
nand U957 (N_957,In_17,In_222);
nor U958 (N_958,In_269,In_1065);
and U959 (N_959,In_1217,In_1688);
nand U960 (N_960,In_1013,In_156);
or U961 (N_961,In_1016,In_1508);
nor U962 (N_962,In_398,In_761);
nor U963 (N_963,In_571,In_1952);
nor U964 (N_964,In_1655,In_1693);
nor U965 (N_965,In_1872,In_1442);
nand U966 (N_966,In_1047,In_136);
nor U967 (N_967,In_182,In_954);
or U968 (N_968,In_118,In_1304);
nor U969 (N_969,In_1498,In_1400);
and U970 (N_970,In_1518,In_605);
nor U971 (N_971,In_1274,In_1032);
nor U972 (N_972,In_852,In_1801);
nor U973 (N_973,In_1331,In_725);
or U974 (N_974,In_618,In_552);
and U975 (N_975,In_1235,In_412);
nand U976 (N_976,In_420,In_1670);
or U977 (N_977,In_551,In_66);
and U978 (N_978,In_1856,In_216);
nand U979 (N_979,In_940,In_1564);
or U980 (N_980,In_832,In_791);
nand U981 (N_981,In_490,In_1131);
and U982 (N_982,In_119,In_38);
nor U983 (N_983,In_1206,In_1202);
nand U984 (N_984,In_2,In_444);
nand U985 (N_985,In_615,In_1739);
and U986 (N_986,In_1867,In_1097);
nand U987 (N_987,In_1347,In_1796);
nand U988 (N_988,In_1094,In_779);
xor U989 (N_989,In_432,In_1246);
or U990 (N_990,In_61,In_1410);
and U991 (N_991,In_536,In_1572);
nand U992 (N_992,In_664,In_917);
nand U993 (N_993,In_1846,In_609);
nor U994 (N_994,In_1374,In_1502);
or U995 (N_995,In_1696,In_752);
or U996 (N_996,In_641,In_1547);
nor U997 (N_997,In_1656,In_1538);
nand U998 (N_998,In_1368,In_1493);
nand U999 (N_999,In_323,In_1694);
and U1000 (N_1000,In_1568,In_319);
or U1001 (N_1001,In_471,In_96);
nor U1002 (N_1002,In_1102,In_1157);
nor U1003 (N_1003,In_1783,In_1607);
and U1004 (N_1004,In_1884,In_1838);
nand U1005 (N_1005,In_141,In_1220);
or U1006 (N_1006,In_1619,In_735);
and U1007 (N_1007,In_1594,In_1320);
nor U1008 (N_1008,In_101,In_1292);
nor U1009 (N_1009,In_1374,In_1039);
or U1010 (N_1010,In_1944,In_1178);
and U1011 (N_1011,In_1710,In_1297);
and U1012 (N_1012,In_1773,In_300);
or U1013 (N_1013,In_1954,In_1816);
or U1014 (N_1014,In_1873,In_1955);
nor U1015 (N_1015,In_1120,In_1036);
and U1016 (N_1016,In_1997,In_616);
nand U1017 (N_1017,In_1582,In_1928);
nand U1018 (N_1018,In_1838,In_1960);
or U1019 (N_1019,In_801,In_1955);
nand U1020 (N_1020,In_851,In_1245);
and U1021 (N_1021,In_386,In_526);
and U1022 (N_1022,In_1519,In_65);
nand U1023 (N_1023,In_499,In_774);
nand U1024 (N_1024,In_1017,In_1847);
nand U1025 (N_1025,In_1071,In_1150);
or U1026 (N_1026,In_372,In_407);
or U1027 (N_1027,In_1626,In_1422);
or U1028 (N_1028,In_760,In_1224);
or U1029 (N_1029,In_1254,In_1895);
xor U1030 (N_1030,In_5,In_1328);
and U1031 (N_1031,In_1681,In_1491);
and U1032 (N_1032,In_888,In_1236);
nor U1033 (N_1033,In_1945,In_1984);
or U1034 (N_1034,In_257,In_378);
nand U1035 (N_1035,In_101,In_196);
or U1036 (N_1036,In_628,In_1820);
or U1037 (N_1037,In_1868,In_1416);
nor U1038 (N_1038,In_1066,In_596);
or U1039 (N_1039,In_1076,In_92);
nand U1040 (N_1040,In_1930,In_147);
and U1041 (N_1041,In_974,In_54);
nand U1042 (N_1042,In_1611,In_73);
nand U1043 (N_1043,In_1494,In_1119);
and U1044 (N_1044,In_993,In_1356);
and U1045 (N_1045,In_928,In_1404);
nor U1046 (N_1046,In_1282,In_476);
nand U1047 (N_1047,In_712,In_1358);
or U1048 (N_1048,In_1097,In_1751);
nand U1049 (N_1049,In_1926,In_1304);
nand U1050 (N_1050,In_261,In_1159);
nor U1051 (N_1051,In_1244,In_1226);
or U1052 (N_1052,In_773,In_1344);
nand U1053 (N_1053,In_1938,In_1886);
nand U1054 (N_1054,In_764,In_951);
or U1055 (N_1055,In_240,In_1282);
or U1056 (N_1056,In_132,In_1766);
nand U1057 (N_1057,In_1277,In_636);
nor U1058 (N_1058,In_1245,In_1606);
or U1059 (N_1059,In_1256,In_1662);
nor U1060 (N_1060,In_113,In_101);
and U1061 (N_1061,In_1560,In_1542);
and U1062 (N_1062,In_1484,In_320);
nand U1063 (N_1063,In_168,In_869);
nand U1064 (N_1064,In_471,In_1331);
nand U1065 (N_1065,In_1260,In_1349);
xnor U1066 (N_1066,In_437,In_6);
and U1067 (N_1067,In_1936,In_580);
nand U1068 (N_1068,In_830,In_1389);
or U1069 (N_1069,In_1593,In_644);
and U1070 (N_1070,In_1726,In_1920);
nor U1071 (N_1071,In_644,In_1347);
nand U1072 (N_1072,In_350,In_699);
or U1073 (N_1073,In_151,In_355);
nand U1074 (N_1074,In_972,In_1162);
or U1075 (N_1075,In_1207,In_789);
or U1076 (N_1076,In_1946,In_261);
nor U1077 (N_1077,In_536,In_603);
or U1078 (N_1078,In_584,In_1998);
or U1079 (N_1079,In_874,In_537);
nand U1080 (N_1080,In_1505,In_838);
nand U1081 (N_1081,In_1758,In_1207);
or U1082 (N_1082,In_775,In_1107);
and U1083 (N_1083,In_441,In_1126);
nor U1084 (N_1084,In_31,In_1397);
nor U1085 (N_1085,In_627,In_448);
or U1086 (N_1086,In_1127,In_164);
nor U1087 (N_1087,In_430,In_1280);
or U1088 (N_1088,In_1611,In_1811);
and U1089 (N_1089,In_1131,In_241);
and U1090 (N_1090,In_1029,In_858);
or U1091 (N_1091,In_1933,In_124);
nor U1092 (N_1092,In_220,In_1311);
nand U1093 (N_1093,In_1224,In_548);
or U1094 (N_1094,In_208,In_1566);
or U1095 (N_1095,In_1256,In_364);
or U1096 (N_1096,In_257,In_1128);
nor U1097 (N_1097,In_1496,In_1514);
nor U1098 (N_1098,In_157,In_1298);
or U1099 (N_1099,In_1116,In_1411);
nor U1100 (N_1100,In_28,In_1849);
xnor U1101 (N_1101,In_828,In_1393);
and U1102 (N_1102,In_420,In_543);
and U1103 (N_1103,In_616,In_558);
nor U1104 (N_1104,In_1326,In_633);
nor U1105 (N_1105,In_1802,In_1403);
nor U1106 (N_1106,In_595,In_805);
nor U1107 (N_1107,In_261,In_271);
and U1108 (N_1108,In_906,In_21);
or U1109 (N_1109,In_1142,In_99);
and U1110 (N_1110,In_207,In_1328);
and U1111 (N_1111,In_1640,In_70);
nand U1112 (N_1112,In_839,In_864);
nand U1113 (N_1113,In_1711,In_79);
or U1114 (N_1114,In_1724,In_262);
nand U1115 (N_1115,In_610,In_1746);
or U1116 (N_1116,In_1384,In_923);
nand U1117 (N_1117,In_79,In_523);
and U1118 (N_1118,In_242,In_546);
nor U1119 (N_1119,In_735,In_436);
and U1120 (N_1120,In_1343,In_956);
nor U1121 (N_1121,In_544,In_480);
or U1122 (N_1122,In_375,In_20);
nor U1123 (N_1123,In_1380,In_975);
nand U1124 (N_1124,In_452,In_1403);
and U1125 (N_1125,In_364,In_1923);
nand U1126 (N_1126,In_1128,In_1609);
xor U1127 (N_1127,In_1174,In_253);
nand U1128 (N_1128,In_644,In_84);
nand U1129 (N_1129,In_1930,In_1098);
nand U1130 (N_1130,In_474,In_1248);
nor U1131 (N_1131,In_102,In_1180);
nand U1132 (N_1132,In_380,In_13);
nor U1133 (N_1133,In_1458,In_1888);
and U1134 (N_1134,In_1834,In_1398);
nand U1135 (N_1135,In_1544,In_1168);
nor U1136 (N_1136,In_295,In_1006);
and U1137 (N_1137,In_1810,In_155);
or U1138 (N_1138,In_93,In_491);
and U1139 (N_1139,In_166,In_225);
nand U1140 (N_1140,In_576,In_1068);
nand U1141 (N_1141,In_716,In_1707);
or U1142 (N_1142,In_1078,In_806);
nor U1143 (N_1143,In_1849,In_792);
and U1144 (N_1144,In_53,In_710);
nand U1145 (N_1145,In_651,In_1669);
nand U1146 (N_1146,In_164,In_1937);
nor U1147 (N_1147,In_1907,In_1612);
or U1148 (N_1148,In_190,In_235);
nand U1149 (N_1149,In_1464,In_1554);
or U1150 (N_1150,In_1814,In_218);
or U1151 (N_1151,In_1854,In_1303);
nand U1152 (N_1152,In_155,In_376);
nor U1153 (N_1153,In_126,In_1755);
nand U1154 (N_1154,In_1803,In_1091);
nor U1155 (N_1155,In_484,In_1217);
or U1156 (N_1156,In_626,In_852);
and U1157 (N_1157,In_514,In_1429);
and U1158 (N_1158,In_882,In_1583);
nor U1159 (N_1159,In_1537,In_1190);
nor U1160 (N_1160,In_135,In_142);
nor U1161 (N_1161,In_1347,In_1603);
or U1162 (N_1162,In_834,In_1900);
and U1163 (N_1163,In_1023,In_1061);
nand U1164 (N_1164,In_582,In_1807);
nand U1165 (N_1165,In_1635,In_675);
or U1166 (N_1166,In_463,In_1679);
nor U1167 (N_1167,In_806,In_984);
and U1168 (N_1168,In_569,In_199);
and U1169 (N_1169,In_1765,In_734);
nand U1170 (N_1170,In_924,In_1725);
nand U1171 (N_1171,In_1535,In_541);
or U1172 (N_1172,In_995,In_1315);
or U1173 (N_1173,In_1264,In_1203);
and U1174 (N_1174,In_851,In_1623);
nand U1175 (N_1175,In_240,In_1458);
and U1176 (N_1176,In_557,In_1469);
and U1177 (N_1177,In_363,In_1055);
nor U1178 (N_1178,In_102,In_1525);
and U1179 (N_1179,In_1270,In_1356);
nor U1180 (N_1180,In_886,In_1614);
nand U1181 (N_1181,In_211,In_1004);
nand U1182 (N_1182,In_318,In_794);
and U1183 (N_1183,In_1459,In_1375);
nand U1184 (N_1184,In_518,In_1794);
nand U1185 (N_1185,In_130,In_1136);
or U1186 (N_1186,In_791,In_537);
nand U1187 (N_1187,In_592,In_908);
and U1188 (N_1188,In_333,In_1239);
nor U1189 (N_1189,In_900,In_830);
or U1190 (N_1190,In_520,In_528);
or U1191 (N_1191,In_1401,In_1633);
or U1192 (N_1192,In_788,In_740);
nor U1193 (N_1193,In_34,In_310);
and U1194 (N_1194,In_598,In_1885);
nand U1195 (N_1195,In_1285,In_555);
or U1196 (N_1196,In_1327,In_1589);
nand U1197 (N_1197,In_1451,In_571);
nor U1198 (N_1198,In_210,In_567);
and U1199 (N_1199,In_618,In_706);
nor U1200 (N_1200,In_1649,In_645);
and U1201 (N_1201,In_1146,In_783);
nor U1202 (N_1202,In_763,In_371);
nor U1203 (N_1203,In_1203,In_1757);
or U1204 (N_1204,In_116,In_164);
and U1205 (N_1205,In_1847,In_1900);
and U1206 (N_1206,In_1290,In_434);
nand U1207 (N_1207,In_1522,In_608);
nor U1208 (N_1208,In_1419,In_1092);
nor U1209 (N_1209,In_259,In_1238);
or U1210 (N_1210,In_42,In_1953);
and U1211 (N_1211,In_1386,In_750);
and U1212 (N_1212,In_326,In_1161);
or U1213 (N_1213,In_1630,In_858);
nor U1214 (N_1214,In_170,In_468);
nor U1215 (N_1215,In_802,In_1793);
nand U1216 (N_1216,In_947,In_23);
or U1217 (N_1217,In_95,In_1277);
and U1218 (N_1218,In_1967,In_1624);
or U1219 (N_1219,In_633,In_1824);
and U1220 (N_1220,In_1178,In_641);
or U1221 (N_1221,In_1586,In_1070);
nor U1222 (N_1222,In_1255,In_1928);
nor U1223 (N_1223,In_177,In_343);
nor U1224 (N_1224,In_974,In_1937);
and U1225 (N_1225,In_1427,In_582);
nand U1226 (N_1226,In_1284,In_26);
nand U1227 (N_1227,In_601,In_545);
xor U1228 (N_1228,In_542,In_805);
nor U1229 (N_1229,In_1811,In_910);
nor U1230 (N_1230,In_1088,In_951);
xnor U1231 (N_1231,In_580,In_879);
or U1232 (N_1232,In_1812,In_1894);
or U1233 (N_1233,In_606,In_1172);
or U1234 (N_1234,In_133,In_1852);
or U1235 (N_1235,In_1282,In_865);
nor U1236 (N_1236,In_1690,In_1999);
nor U1237 (N_1237,In_1814,In_3);
nand U1238 (N_1238,In_1738,In_502);
nand U1239 (N_1239,In_549,In_1680);
and U1240 (N_1240,In_1982,In_901);
nand U1241 (N_1241,In_1044,In_885);
nor U1242 (N_1242,In_1167,In_1586);
nor U1243 (N_1243,In_1167,In_102);
or U1244 (N_1244,In_649,In_806);
nand U1245 (N_1245,In_1456,In_688);
and U1246 (N_1246,In_384,In_1391);
or U1247 (N_1247,In_1046,In_5);
nand U1248 (N_1248,In_430,In_487);
nor U1249 (N_1249,In_966,In_1678);
nand U1250 (N_1250,In_1424,In_227);
and U1251 (N_1251,In_1090,In_1759);
nor U1252 (N_1252,In_844,In_1127);
and U1253 (N_1253,In_1818,In_1067);
and U1254 (N_1254,In_820,In_1740);
or U1255 (N_1255,In_1296,In_1464);
nand U1256 (N_1256,In_1391,In_1443);
nand U1257 (N_1257,In_295,In_588);
or U1258 (N_1258,In_369,In_1679);
nor U1259 (N_1259,In_1108,In_421);
nand U1260 (N_1260,In_1642,In_1056);
nor U1261 (N_1261,In_928,In_1908);
nand U1262 (N_1262,In_817,In_1346);
nor U1263 (N_1263,In_1861,In_1900);
nand U1264 (N_1264,In_898,In_681);
nand U1265 (N_1265,In_514,In_1724);
and U1266 (N_1266,In_1321,In_422);
and U1267 (N_1267,In_552,In_74);
nor U1268 (N_1268,In_1446,In_1358);
nor U1269 (N_1269,In_342,In_1618);
nand U1270 (N_1270,In_513,In_1516);
and U1271 (N_1271,In_1333,In_117);
nand U1272 (N_1272,In_946,In_1895);
and U1273 (N_1273,In_711,In_918);
and U1274 (N_1274,In_1138,In_1260);
nor U1275 (N_1275,In_103,In_439);
or U1276 (N_1276,In_1838,In_1329);
nor U1277 (N_1277,In_1083,In_1118);
nand U1278 (N_1278,In_280,In_1919);
or U1279 (N_1279,In_509,In_254);
and U1280 (N_1280,In_1452,In_239);
nor U1281 (N_1281,In_232,In_1872);
nand U1282 (N_1282,In_1615,In_90);
nor U1283 (N_1283,In_1274,In_460);
nor U1284 (N_1284,In_1426,In_1959);
nand U1285 (N_1285,In_106,In_746);
or U1286 (N_1286,In_374,In_1004);
nand U1287 (N_1287,In_153,In_991);
nor U1288 (N_1288,In_16,In_1540);
nor U1289 (N_1289,In_281,In_1990);
nand U1290 (N_1290,In_1079,In_1328);
nor U1291 (N_1291,In_459,In_832);
and U1292 (N_1292,In_742,In_705);
and U1293 (N_1293,In_894,In_1272);
nor U1294 (N_1294,In_1397,In_943);
nor U1295 (N_1295,In_488,In_295);
and U1296 (N_1296,In_928,In_803);
and U1297 (N_1297,In_512,In_1897);
nor U1298 (N_1298,In_1366,In_1465);
and U1299 (N_1299,In_1531,In_1907);
and U1300 (N_1300,In_1053,In_1899);
or U1301 (N_1301,In_109,In_1920);
nand U1302 (N_1302,In_247,In_1861);
or U1303 (N_1303,In_658,In_803);
nand U1304 (N_1304,In_1423,In_575);
or U1305 (N_1305,In_888,In_1338);
or U1306 (N_1306,In_577,In_120);
and U1307 (N_1307,In_66,In_1247);
nor U1308 (N_1308,In_743,In_1913);
nand U1309 (N_1309,In_1525,In_541);
nand U1310 (N_1310,In_975,In_1480);
nand U1311 (N_1311,In_355,In_502);
nor U1312 (N_1312,In_1270,In_1313);
and U1313 (N_1313,In_127,In_1800);
nor U1314 (N_1314,In_159,In_1761);
or U1315 (N_1315,In_441,In_754);
or U1316 (N_1316,In_460,In_92);
nor U1317 (N_1317,In_1389,In_624);
and U1318 (N_1318,In_173,In_1093);
and U1319 (N_1319,In_1142,In_51);
nand U1320 (N_1320,In_153,In_82);
and U1321 (N_1321,In_190,In_494);
nand U1322 (N_1322,In_73,In_316);
and U1323 (N_1323,In_1777,In_1942);
and U1324 (N_1324,In_51,In_607);
and U1325 (N_1325,In_564,In_1603);
nand U1326 (N_1326,In_300,In_800);
nand U1327 (N_1327,In_1292,In_94);
and U1328 (N_1328,In_1247,In_1643);
or U1329 (N_1329,In_1427,In_1156);
nor U1330 (N_1330,In_1011,In_39);
or U1331 (N_1331,In_787,In_1307);
and U1332 (N_1332,In_1313,In_1839);
nor U1333 (N_1333,In_1730,In_61);
and U1334 (N_1334,In_485,In_1392);
and U1335 (N_1335,In_1770,In_1353);
nor U1336 (N_1336,In_348,In_621);
nand U1337 (N_1337,In_676,In_1403);
and U1338 (N_1338,In_1053,In_1988);
or U1339 (N_1339,In_1087,In_1268);
nand U1340 (N_1340,In_376,In_638);
nor U1341 (N_1341,In_729,In_99);
nor U1342 (N_1342,In_1995,In_182);
nor U1343 (N_1343,In_1254,In_49);
or U1344 (N_1344,In_108,In_1103);
and U1345 (N_1345,In_796,In_1385);
nand U1346 (N_1346,In_1510,In_624);
xor U1347 (N_1347,In_1674,In_780);
xnor U1348 (N_1348,In_733,In_1408);
nor U1349 (N_1349,In_10,In_1551);
or U1350 (N_1350,In_1224,In_546);
or U1351 (N_1351,In_1341,In_1381);
nand U1352 (N_1352,In_1416,In_1543);
nand U1353 (N_1353,In_233,In_1437);
nand U1354 (N_1354,In_17,In_1978);
nor U1355 (N_1355,In_1240,In_1505);
nor U1356 (N_1356,In_1821,In_1778);
or U1357 (N_1357,In_197,In_462);
or U1358 (N_1358,In_602,In_1546);
and U1359 (N_1359,In_1387,In_1553);
or U1360 (N_1360,In_1702,In_370);
nand U1361 (N_1361,In_1333,In_806);
nand U1362 (N_1362,In_523,In_1215);
nand U1363 (N_1363,In_380,In_135);
or U1364 (N_1364,In_238,In_1546);
and U1365 (N_1365,In_1843,In_1052);
or U1366 (N_1366,In_1989,In_317);
or U1367 (N_1367,In_1721,In_1809);
or U1368 (N_1368,In_808,In_945);
and U1369 (N_1369,In_51,In_1334);
or U1370 (N_1370,In_1956,In_152);
nand U1371 (N_1371,In_875,In_710);
and U1372 (N_1372,In_183,In_99);
nor U1373 (N_1373,In_1241,In_972);
nand U1374 (N_1374,In_1085,In_1020);
or U1375 (N_1375,In_38,In_1585);
nand U1376 (N_1376,In_620,In_574);
nor U1377 (N_1377,In_711,In_686);
nand U1378 (N_1378,In_215,In_1362);
or U1379 (N_1379,In_77,In_1280);
nand U1380 (N_1380,In_257,In_142);
nand U1381 (N_1381,In_1777,In_1353);
and U1382 (N_1382,In_965,In_1660);
or U1383 (N_1383,In_1918,In_811);
or U1384 (N_1384,In_714,In_610);
nor U1385 (N_1385,In_1257,In_731);
nand U1386 (N_1386,In_1629,In_1127);
xnor U1387 (N_1387,In_81,In_1399);
or U1388 (N_1388,In_153,In_874);
and U1389 (N_1389,In_1234,In_1381);
or U1390 (N_1390,In_158,In_1019);
or U1391 (N_1391,In_95,In_211);
nor U1392 (N_1392,In_1601,In_633);
nor U1393 (N_1393,In_1210,In_1645);
nand U1394 (N_1394,In_26,In_162);
or U1395 (N_1395,In_1953,In_216);
or U1396 (N_1396,In_1865,In_1508);
and U1397 (N_1397,In_1769,In_1380);
or U1398 (N_1398,In_555,In_1814);
nand U1399 (N_1399,In_1684,In_762);
nand U1400 (N_1400,In_1430,In_906);
and U1401 (N_1401,In_32,In_612);
nand U1402 (N_1402,In_1056,In_1334);
nor U1403 (N_1403,In_1986,In_1880);
nand U1404 (N_1404,In_1988,In_1377);
and U1405 (N_1405,In_1860,In_1436);
nand U1406 (N_1406,In_250,In_1009);
or U1407 (N_1407,In_1311,In_162);
or U1408 (N_1408,In_60,In_1369);
nor U1409 (N_1409,In_1597,In_1999);
or U1410 (N_1410,In_275,In_1570);
and U1411 (N_1411,In_1170,In_929);
nand U1412 (N_1412,In_916,In_36);
and U1413 (N_1413,In_499,In_1868);
nor U1414 (N_1414,In_958,In_1267);
or U1415 (N_1415,In_64,In_1896);
or U1416 (N_1416,In_1550,In_1424);
and U1417 (N_1417,In_295,In_1129);
nor U1418 (N_1418,In_1754,In_421);
nor U1419 (N_1419,In_1295,In_1018);
nor U1420 (N_1420,In_234,In_970);
and U1421 (N_1421,In_922,In_1462);
nor U1422 (N_1422,In_1549,In_319);
or U1423 (N_1423,In_932,In_1925);
or U1424 (N_1424,In_1448,In_1514);
or U1425 (N_1425,In_685,In_490);
and U1426 (N_1426,In_539,In_265);
xor U1427 (N_1427,In_1621,In_1608);
and U1428 (N_1428,In_106,In_1687);
nand U1429 (N_1429,In_239,In_1340);
or U1430 (N_1430,In_781,In_1017);
or U1431 (N_1431,In_157,In_1453);
or U1432 (N_1432,In_1389,In_850);
or U1433 (N_1433,In_138,In_1911);
or U1434 (N_1434,In_453,In_315);
or U1435 (N_1435,In_1453,In_1894);
or U1436 (N_1436,In_1413,In_1596);
nand U1437 (N_1437,In_489,In_1926);
or U1438 (N_1438,In_1243,In_880);
nor U1439 (N_1439,In_1070,In_926);
and U1440 (N_1440,In_931,In_1737);
nand U1441 (N_1441,In_1935,In_1331);
nand U1442 (N_1442,In_28,In_162);
nand U1443 (N_1443,In_1631,In_1763);
and U1444 (N_1444,In_592,In_1198);
and U1445 (N_1445,In_844,In_1128);
nor U1446 (N_1446,In_271,In_1943);
nand U1447 (N_1447,In_463,In_1913);
and U1448 (N_1448,In_1412,In_649);
nand U1449 (N_1449,In_166,In_1113);
nor U1450 (N_1450,In_794,In_134);
and U1451 (N_1451,In_329,In_1246);
and U1452 (N_1452,In_791,In_843);
and U1453 (N_1453,In_146,In_628);
nand U1454 (N_1454,In_795,In_1897);
nand U1455 (N_1455,In_1905,In_574);
nor U1456 (N_1456,In_345,In_686);
nand U1457 (N_1457,In_1938,In_549);
nor U1458 (N_1458,In_1752,In_1786);
nor U1459 (N_1459,In_225,In_1045);
or U1460 (N_1460,In_866,In_1743);
nand U1461 (N_1461,In_737,In_520);
and U1462 (N_1462,In_136,In_97);
or U1463 (N_1463,In_1082,In_214);
nor U1464 (N_1464,In_665,In_1857);
and U1465 (N_1465,In_1181,In_57);
and U1466 (N_1466,In_689,In_1334);
or U1467 (N_1467,In_257,In_1913);
nand U1468 (N_1468,In_1283,In_1997);
or U1469 (N_1469,In_167,In_1566);
xor U1470 (N_1470,In_790,In_1128);
nand U1471 (N_1471,In_1879,In_1747);
nor U1472 (N_1472,In_402,In_1176);
or U1473 (N_1473,In_749,In_318);
and U1474 (N_1474,In_1390,In_1123);
nor U1475 (N_1475,In_39,In_907);
or U1476 (N_1476,In_363,In_1910);
nor U1477 (N_1477,In_1134,In_1115);
and U1478 (N_1478,In_986,In_315);
or U1479 (N_1479,In_1002,In_113);
or U1480 (N_1480,In_329,In_492);
nand U1481 (N_1481,In_1642,In_1332);
or U1482 (N_1482,In_1810,In_1812);
nor U1483 (N_1483,In_1340,In_337);
or U1484 (N_1484,In_233,In_252);
nand U1485 (N_1485,In_1251,In_1740);
or U1486 (N_1486,In_1889,In_1859);
nor U1487 (N_1487,In_344,In_1966);
and U1488 (N_1488,In_129,In_228);
and U1489 (N_1489,In_1709,In_322);
nor U1490 (N_1490,In_946,In_700);
nand U1491 (N_1491,In_1173,In_32);
and U1492 (N_1492,In_775,In_1031);
or U1493 (N_1493,In_636,In_499);
nand U1494 (N_1494,In_641,In_321);
or U1495 (N_1495,In_1716,In_630);
nand U1496 (N_1496,In_176,In_915);
nand U1497 (N_1497,In_1333,In_1190);
or U1498 (N_1498,In_401,In_371);
and U1499 (N_1499,In_1837,In_896);
nor U1500 (N_1500,In_955,In_976);
or U1501 (N_1501,In_849,In_893);
nand U1502 (N_1502,In_559,In_1217);
nand U1503 (N_1503,In_737,In_108);
or U1504 (N_1504,In_1293,In_468);
and U1505 (N_1505,In_934,In_227);
nor U1506 (N_1506,In_1023,In_526);
nand U1507 (N_1507,In_1077,In_706);
nand U1508 (N_1508,In_1101,In_1804);
nand U1509 (N_1509,In_597,In_1306);
and U1510 (N_1510,In_1260,In_1609);
or U1511 (N_1511,In_1354,In_822);
or U1512 (N_1512,In_875,In_1531);
or U1513 (N_1513,In_939,In_1423);
nand U1514 (N_1514,In_1073,In_370);
nand U1515 (N_1515,In_1919,In_1568);
nor U1516 (N_1516,In_784,In_64);
and U1517 (N_1517,In_575,In_1146);
or U1518 (N_1518,In_35,In_1159);
nand U1519 (N_1519,In_1392,In_265);
or U1520 (N_1520,In_355,In_256);
or U1521 (N_1521,In_227,In_1620);
or U1522 (N_1522,In_761,In_1056);
nor U1523 (N_1523,In_1505,In_1892);
or U1524 (N_1524,In_1871,In_103);
or U1525 (N_1525,In_1224,In_419);
xor U1526 (N_1526,In_1262,In_1930);
nand U1527 (N_1527,In_698,In_884);
or U1528 (N_1528,In_751,In_1350);
and U1529 (N_1529,In_1638,In_1290);
nor U1530 (N_1530,In_908,In_1666);
or U1531 (N_1531,In_1363,In_932);
and U1532 (N_1532,In_803,In_1572);
nand U1533 (N_1533,In_691,In_571);
and U1534 (N_1534,In_442,In_1743);
or U1535 (N_1535,In_1527,In_1423);
or U1536 (N_1536,In_583,In_572);
nand U1537 (N_1537,In_341,In_1642);
nand U1538 (N_1538,In_565,In_1363);
and U1539 (N_1539,In_703,In_1222);
nand U1540 (N_1540,In_240,In_1921);
nand U1541 (N_1541,In_1355,In_304);
nand U1542 (N_1542,In_1978,In_327);
nand U1543 (N_1543,In_292,In_620);
or U1544 (N_1544,In_5,In_1586);
nand U1545 (N_1545,In_1531,In_1676);
nand U1546 (N_1546,In_341,In_496);
nor U1547 (N_1547,In_649,In_1524);
and U1548 (N_1548,In_70,In_137);
and U1549 (N_1549,In_1767,In_1314);
nand U1550 (N_1550,In_1964,In_1621);
nand U1551 (N_1551,In_198,In_1609);
and U1552 (N_1552,In_1908,In_265);
xor U1553 (N_1553,In_1908,In_1051);
xnor U1554 (N_1554,In_1318,In_513);
nand U1555 (N_1555,In_1544,In_1310);
nand U1556 (N_1556,In_1541,In_1460);
xor U1557 (N_1557,In_1345,In_1453);
nand U1558 (N_1558,In_729,In_837);
nand U1559 (N_1559,In_917,In_796);
nor U1560 (N_1560,In_1400,In_1303);
nand U1561 (N_1561,In_24,In_92);
or U1562 (N_1562,In_1078,In_1218);
nor U1563 (N_1563,In_779,In_1436);
nand U1564 (N_1564,In_1404,In_446);
nor U1565 (N_1565,In_1495,In_989);
nor U1566 (N_1566,In_848,In_639);
and U1567 (N_1567,In_274,In_1103);
nand U1568 (N_1568,In_1867,In_989);
nand U1569 (N_1569,In_1745,In_1659);
and U1570 (N_1570,In_1238,In_977);
nor U1571 (N_1571,In_1480,In_1767);
nor U1572 (N_1572,In_1212,In_1744);
nor U1573 (N_1573,In_797,In_274);
or U1574 (N_1574,In_189,In_1329);
and U1575 (N_1575,In_130,In_350);
or U1576 (N_1576,In_1656,In_1110);
nor U1577 (N_1577,In_1783,In_830);
or U1578 (N_1578,In_53,In_1879);
nor U1579 (N_1579,In_140,In_30);
or U1580 (N_1580,In_777,In_226);
or U1581 (N_1581,In_1915,In_1148);
nand U1582 (N_1582,In_1931,In_1848);
nor U1583 (N_1583,In_874,In_1916);
or U1584 (N_1584,In_54,In_379);
and U1585 (N_1585,In_1272,In_42);
or U1586 (N_1586,In_801,In_783);
and U1587 (N_1587,In_1218,In_1454);
and U1588 (N_1588,In_677,In_1749);
and U1589 (N_1589,In_1160,In_983);
nand U1590 (N_1590,In_43,In_1766);
nand U1591 (N_1591,In_676,In_736);
nor U1592 (N_1592,In_1442,In_1077);
and U1593 (N_1593,In_208,In_1044);
xor U1594 (N_1594,In_993,In_169);
and U1595 (N_1595,In_309,In_366);
nor U1596 (N_1596,In_1335,In_787);
or U1597 (N_1597,In_1887,In_421);
nor U1598 (N_1598,In_1548,In_909);
nand U1599 (N_1599,In_868,In_924);
nand U1600 (N_1600,In_1265,In_1538);
and U1601 (N_1601,In_863,In_155);
nor U1602 (N_1602,In_562,In_419);
and U1603 (N_1603,In_542,In_341);
nand U1604 (N_1604,In_1545,In_653);
nor U1605 (N_1605,In_1156,In_1323);
and U1606 (N_1606,In_302,In_1365);
nand U1607 (N_1607,In_952,In_1178);
and U1608 (N_1608,In_1588,In_1943);
or U1609 (N_1609,In_572,In_1896);
nor U1610 (N_1610,In_858,In_62);
nand U1611 (N_1611,In_1922,In_1141);
nor U1612 (N_1612,In_1150,In_748);
xnor U1613 (N_1613,In_520,In_1378);
and U1614 (N_1614,In_868,In_484);
nand U1615 (N_1615,In_511,In_14);
and U1616 (N_1616,In_762,In_1617);
and U1617 (N_1617,In_1799,In_586);
nor U1618 (N_1618,In_809,In_1560);
and U1619 (N_1619,In_1342,In_1149);
and U1620 (N_1620,In_20,In_423);
and U1621 (N_1621,In_409,In_1917);
nand U1622 (N_1622,In_1586,In_73);
or U1623 (N_1623,In_1919,In_1952);
and U1624 (N_1624,In_1207,In_502);
nor U1625 (N_1625,In_610,In_371);
nor U1626 (N_1626,In_1660,In_854);
and U1627 (N_1627,In_490,In_1150);
and U1628 (N_1628,In_1221,In_1728);
nand U1629 (N_1629,In_1434,In_1379);
nor U1630 (N_1630,In_1072,In_1076);
nor U1631 (N_1631,In_1211,In_1306);
and U1632 (N_1632,In_1579,In_1763);
nor U1633 (N_1633,In_1620,In_651);
and U1634 (N_1634,In_1007,In_752);
and U1635 (N_1635,In_1045,In_1451);
nor U1636 (N_1636,In_1537,In_275);
or U1637 (N_1637,In_836,In_1525);
and U1638 (N_1638,In_1873,In_1312);
and U1639 (N_1639,In_1592,In_1927);
nand U1640 (N_1640,In_1033,In_1222);
and U1641 (N_1641,In_1315,In_1760);
and U1642 (N_1642,In_1843,In_322);
or U1643 (N_1643,In_562,In_1017);
nand U1644 (N_1644,In_507,In_1273);
nor U1645 (N_1645,In_1657,In_437);
nand U1646 (N_1646,In_797,In_685);
or U1647 (N_1647,In_1943,In_461);
nand U1648 (N_1648,In_30,In_142);
nor U1649 (N_1649,In_1801,In_610);
nor U1650 (N_1650,In_1946,In_1829);
nor U1651 (N_1651,In_1936,In_982);
nor U1652 (N_1652,In_1736,In_412);
or U1653 (N_1653,In_1831,In_1462);
nand U1654 (N_1654,In_142,In_191);
nand U1655 (N_1655,In_207,In_132);
nor U1656 (N_1656,In_1893,In_980);
nand U1657 (N_1657,In_464,In_720);
and U1658 (N_1658,In_1198,In_1021);
nor U1659 (N_1659,In_472,In_803);
nand U1660 (N_1660,In_275,In_1267);
nand U1661 (N_1661,In_1827,In_1989);
nor U1662 (N_1662,In_1307,In_1444);
and U1663 (N_1663,In_874,In_1352);
and U1664 (N_1664,In_1542,In_597);
and U1665 (N_1665,In_1289,In_1996);
and U1666 (N_1666,In_429,In_1);
and U1667 (N_1667,In_1866,In_1780);
nand U1668 (N_1668,In_466,In_504);
or U1669 (N_1669,In_1610,In_304);
and U1670 (N_1670,In_902,In_484);
or U1671 (N_1671,In_1443,In_908);
nor U1672 (N_1672,In_1868,In_829);
or U1673 (N_1673,In_1183,In_1938);
and U1674 (N_1674,In_91,In_1057);
and U1675 (N_1675,In_1422,In_474);
and U1676 (N_1676,In_352,In_488);
nand U1677 (N_1677,In_688,In_972);
nor U1678 (N_1678,In_925,In_175);
nor U1679 (N_1679,In_1692,In_676);
or U1680 (N_1680,In_174,In_196);
and U1681 (N_1681,In_173,In_1288);
nor U1682 (N_1682,In_1264,In_1452);
or U1683 (N_1683,In_1570,In_1561);
and U1684 (N_1684,In_235,In_529);
nor U1685 (N_1685,In_979,In_1075);
nand U1686 (N_1686,In_1224,In_434);
nand U1687 (N_1687,In_1297,In_682);
nor U1688 (N_1688,In_199,In_1131);
nor U1689 (N_1689,In_1011,In_615);
nand U1690 (N_1690,In_1966,In_812);
nor U1691 (N_1691,In_337,In_1317);
or U1692 (N_1692,In_1964,In_549);
or U1693 (N_1693,In_1209,In_376);
and U1694 (N_1694,In_525,In_1930);
nor U1695 (N_1695,In_1044,In_586);
or U1696 (N_1696,In_255,In_1666);
or U1697 (N_1697,In_247,In_990);
and U1698 (N_1698,In_1553,In_428);
or U1699 (N_1699,In_758,In_200);
nand U1700 (N_1700,In_1505,In_716);
and U1701 (N_1701,In_190,In_988);
nor U1702 (N_1702,In_761,In_1051);
nor U1703 (N_1703,In_565,In_1229);
nor U1704 (N_1704,In_1476,In_1858);
or U1705 (N_1705,In_74,In_257);
nor U1706 (N_1706,In_1393,In_434);
nand U1707 (N_1707,In_335,In_735);
and U1708 (N_1708,In_1928,In_528);
and U1709 (N_1709,In_1485,In_296);
nand U1710 (N_1710,In_1825,In_1082);
nor U1711 (N_1711,In_69,In_407);
nand U1712 (N_1712,In_1117,In_170);
nand U1713 (N_1713,In_641,In_1624);
nor U1714 (N_1714,In_8,In_352);
nand U1715 (N_1715,In_589,In_849);
xnor U1716 (N_1716,In_1762,In_586);
nand U1717 (N_1717,In_473,In_790);
nand U1718 (N_1718,In_964,In_1571);
and U1719 (N_1719,In_232,In_1294);
nand U1720 (N_1720,In_764,In_1550);
nand U1721 (N_1721,In_1855,In_257);
nor U1722 (N_1722,In_1871,In_1041);
nand U1723 (N_1723,In_1157,In_998);
and U1724 (N_1724,In_1564,In_1471);
or U1725 (N_1725,In_1244,In_7);
or U1726 (N_1726,In_668,In_114);
nand U1727 (N_1727,In_777,In_411);
or U1728 (N_1728,In_393,In_157);
or U1729 (N_1729,In_1160,In_1579);
nand U1730 (N_1730,In_1977,In_530);
nand U1731 (N_1731,In_1812,In_556);
nor U1732 (N_1732,In_221,In_775);
nand U1733 (N_1733,In_1071,In_562);
nand U1734 (N_1734,In_856,In_331);
and U1735 (N_1735,In_1771,In_408);
and U1736 (N_1736,In_1682,In_1489);
nand U1737 (N_1737,In_1308,In_168);
nor U1738 (N_1738,In_1167,In_1225);
nand U1739 (N_1739,In_1325,In_24);
and U1740 (N_1740,In_1980,In_1732);
and U1741 (N_1741,In_1103,In_1824);
nand U1742 (N_1742,In_1782,In_793);
nor U1743 (N_1743,In_381,In_470);
nor U1744 (N_1744,In_721,In_1230);
or U1745 (N_1745,In_415,In_531);
and U1746 (N_1746,In_1772,In_1608);
nand U1747 (N_1747,In_528,In_322);
or U1748 (N_1748,In_829,In_741);
nor U1749 (N_1749,In_1538,In_179);
or U1750 (N_1750,In_459,In_1787);
nor U1751 (N_1751,In_379,In_392);
nor U1752 (N_1752,In_289,In_581);
nor U1753 (N_1753,In_122,In_1890);
or U1754 (N_1754,In_1771,In_256);
nor U1755 (N_1755,In_1968,In_1100);
nor U1756 (N_1756,In_534,In_396);
or U1757 (N_1757,In_84,In_120);
and U1758 (N_1758,In_1704,In_1962);
or U1759 (N_1759,In_556,In_728);
or U1760 (N_1760,In_57,In_577);
nand U1761 (N_1761,In_1080,In_1690);
nor U1762 (N_1762,In_184,In_775);
nor U1763 (N_1763,In_262,In_1467);
and U1764 (N_1764,In_189,In_1154);
nand U1765 (N_1765,In_688,In_1616);
or U1766 (N_1766,In_808,In_1425);
nand U1767 (N_1767,In_1650,In_200);
and U1768 (N_1768,In_552,In_732);
nand U1769 (N_1769,In_886,In_1985);
or U1770 (N_1770,In_1456,In_1721);
and U1771 (N_1771,In_903,In_1000);
or U1772 (N_1772,In_725,In_313);
or U1773 (N_1773,In_1853,In_98);
nand U1774 (N_1774,In_811,In_80);
nand U1775 (N_1775,In_613,In_348);
xor U1776 (N_1776,In_671,In_959);
or U1777 (N_1777,In_1668,In_734);
or U1778 (N_1778,In_155,In_1884);
nor U1779 (N_1779,In_1345,In_989);
and U1780 (N_1780,In_777,In_1866);
nand U1781 (N_1781,In_1898,In_1059);
xor U1782 (N_1782,In_1367,In_787);
nand U1783 (N_1783,In_433,In_1908);
nand U1784 (N_1784,In_336,In_480);
nor U1785 (N_1785,In_1315,In_1972);
nand U1786 (N_1786,In_207,In_140);
nor U1787 (N_1787,In_965,In_1988);
or U1788 (N_1788,In_823,In_1009);
nand U1789 (N_1789,In_287,In_1950);
and U1790 (N_1790,In_78,In_1177);
nand U1791 (N_1791,In_606,In_1909);
or U1792 (N_1792,In_1843,In_278);
nor U1793 (N_1793,In_807,In_1625);
and U1794 (N_1794,In_1703,In_1670);
or U1795 (N_1795,In_264,In_105);
nor U1796 (N_1796,In_166,In_252);
nand U1797 (N_1797,In_574,In_1172);
or U1798 (N_1798,In_755,In_16);
nand U1799 (N_1799,In_1844,In_1106);
nor U1800 (N_1800,In_1304,In_834);
or U1801 (N_1801,In_1582,In_83);
or U1802 (N_1802,In_921,In_1368);
or U1803 (N_1803,In_770,In_646);
or U1804 (N_1804,In_1137,In_878);
nor U1805 (N_1805,In_1558,In_782);
nor U1806 (N_1806,In_1859,In_1798);
nor U1807 (N_1807,In_1353,In_182);
nand U1808 (N_1808,In_1440,In_465);
or U1809 (N_1809,In_63,In_298);
xnor U1810 (N_1810,In_1130,In_1841);
xor U1811 (N_1811,In_789,In_205);
nor U1812 (N_1812,In_1820,In_1019);
nand U1813 (N_1813,In_1643,In_1238);
nor U1814 (N_1814,In_1700,In_1617);
or U1815 (N_1815,In_1064,In_1362);
and U1816 (N_1816,In_1865,In_579);
nand U1817 (N_1817,In_906,In_1234);
and U1818 (N_1818,In_669,In_999);
nor U1819 (N_1819,In_664,In_1193);
nand U1820 (N_1820,In_322,In_429);
nor U1821 (N_1821,In_1929,In_1749);
and U1822 (N_1822,In_1043,In_1939);
and U1823 (N_1823,In_1213,In_510);
or U1824 (N_1824,In_559,In_1839);
nor U1825 (N_1825,In_325,In_1822);
nand U1826 (N_1826,In_1210,In_282);
or U1827 (N_1827,In_869,In_1673);
or U1828 (N_1828,In_1265,In_484);
or U1829 (N_1829,In_1032,In_864);
nand U1830 (N_1830,In_802,In_78);
and U1831 (N_1831,In_1843,In_1252);
nand U1832 (N_1832,In_778,In_762);
or U1833 (N_1833,In_509,In_900);
or U1834 (N_1834,In_821,In_1756);
nand U1835 (N_1835,In_1682,In_65);
and U1836 (N_1836,In_673,In_1903);
or U1837 (N_1837,In_1603,In_610);
or U1838 (N_1838,In_1436,In_1082);
nand U1839 (N_1839,In_1991,In_1223);
nor U1840 (N_1840,In_308,In_1446);
nand U1841 (N_1841,In_1620,In_1128);
nand U1842 (N_1842,In_917,In_88);
nand U1843 (N_1843,In_562,In_560);
and U1844 (N_1844,In_1281,In_34);
or U1845 (N_1845,In_545,In_1804);
nor U1846 (N_1846,In_1151,In_1213);
nand U1847 (N_1847,In_1152,In_685);
nor U1848 (N_1848,In_1294,In_733);
nor U1849 (N_1849,In_143,In_609);
or U1850 (N_1850,In_204,In_579);
or U1851 (N_1851,In_499,In_616);
or U1852 (N_1852,In_1604,In_417);
nand U1853 (N_1853,In_456,In_1335);
nand U1854 (N_1854,In_512,In_1499);
and U1855 (N_1855,In_669,In_1272);
or U1856 (N_1856,In_793,In_303);
nand U1857 (N_1857,In_143,In_289);
or U1858 (N_1858,In_1485,In_1710);
and U1859 (N_1859,In_1309,In_1050);
or U1860 (N_1860,In_7,In_1812);
nand U1861 (N_1861,In_452,In_852);
and U1862 (N_1862,In_669,In_1706);
and U1863 (N_1863,In_201,In_99);
or U1864 (N_1864,In_1673,In_594);
nand U1865 (N_1865,In_1528,In_1190);
or U1866 (N_1866,In_1805,In_74);
nand U1867 (N_1867,In_294,In_1084);
and U1868 (N_1868,In_864,In_821);
nor U1869 (N_1869,In_753,In_1607);
and U1870 (N_1870,In_214,In_1743);
nor U1871 (N_1871,In_1999,In_140);
and U1872 (N_1872,In_550,In_1914);
and U1873 (N_1873,In_1617,In_1223);
nand U1874 (N_1874,In_930,In_1921);
nor U1875 (N_1875,In_459,In_946);
and U1876 (N_1876,In_357,In_1006);
nand U1877 (N_1877,In_409,In_320);
nor U1878 (N_1878,In_635,In_257);
and U1879 (N_1879,In_13,In_1487);
and U1880 (N_1880,In_149,In_92);
and U1881 (N_1881,In_240,In_1205);
nor U1882 (N_1882,In_694,In_719);
nor U1883 (N_1883,In_1310,In_1447);
nand U1884 (N_1884,In_1766,In_1555);
xor U1885 (N_1885,In_1495,In_1346);
and U1886 (N_1886,In_875,In_1749);
nand U1887 (N_1887,In_712,In_72);
or U1888 (N_1888,In_1036,In_397);
nor U1889 (N_1889,In_1285,In_389);
and U1890 (N_1890,In_238,In_1430);
or U1891 (N_1891,In_1496,In_693);
nand U1892 (N_1892,In_895,In_107);
and U1893 (N_1893,In_1134,In_344);
or U1894 (N_1894,In_1939,In_1194);
and U1895 (N_1895,In_1119,In_717);
and U1896 (N_1896,In_342,In_1835);
nor U1897 (N_1897,In_1454,In_1556);
and U1898 (N_1898,In_3,In_1046);
nor U1899 (N_1899,In_1591,In_621);
or U1900 (N_1900,In_1414,In_503);
or U1901 (N_1901,In_1086,In_1404);
or U1902 (N_1902,In_930,In_931);
nand U1903 (N_1903,In_742,In_471);
or U1904 (N_1904,In_933,In_162);
nand U1905 (N_1905,In_1156,In_1975);
or U1906 (N_1906,In_606,In_266);
xnor U1907 (N_1907,In_1332,In_467);
nor U1908 (N_1908,In_849,In_1059);
and U1909 (N_1909,In_1485,In_341);
or U1910 (N_1910,In_1571,In_1014);
nor U1911 (N_1911,In_1000,In_1884);
nand U1912 (N_1912,In_338,In_509);
nand U1913 (N_1913,In_1357,In_1573);
and U1914 (N_1914,In_1407,In_238);
or U1915 (N_1915,In_620,In_1372);
and U1916 (N_1916,In_1759,In_350);
nand U1917 (N_1917,In_1796,In_1045);
or U1918 (N_1918,In_1909,In_1210);
xnor U1919 (N_1919,In_1489,In_1016);
or U1920 (N_1920,In_797,In_1689);
nor U1921 (N_1921,In_255,In_1610);
nor U1922 (N_1922,In_310,In_393);
or U1923 (N_1923,In_1966,In_883);
nor U1924 (N_1924,In_569,In_1128);
and U1925 (N_1925,In_1781,In_1829);
nand U1926 (N_1926,In_947,In_1247);
nor U1927 (N_1927,In_1820,In_1422);
and U1928 (N_1928,In_1776,In_363);
nand U1929 (N_1929,In_896,In_1878);
and U1930 (N_1930,In_926,In_184);
or U1931 (N_1931,In_150,In_1352);
and U1932 (N_1932,In_1223,In_1640);
nor U1933 (N_1933,In_760,In_21);
nand U1934 (N_1934,In_15,In_480);
nand U1935 (N_1935,In_1058,In_851);
nor U1936 (N_1936,In_767,In_390);
and U1937 (N_1937,In_942,In_1637);
and U1938 (N_1938,In_1402,In_549);
nand U1939 (N_1939,In_579,In_1398);
and U1940 (N_1940,In_268,In_1220);
nor U1941 (N_1941,In_1241,In_29);
and U1942 (N_1942,In_1827,In_332);
nand U1943 (N_1943,In_844,In_638);
or U1944 (N_1944,In_1799,In_75);
nand U1945 (N_1945,In_1865,In_272);
and U1946 (N_1946,In_401,In_1599);
or U1947 (N_1947,In_1182,In_832);
nand U1948 (N_1948,In_1064,In_105);
nand U1949 (N_1949,In_884,In_1999);
nand U1950 (N_1950,In_68,In_800);
nand U1951 (N_1951,In_151,In_719);
nor U1952 (N_1952,In_1445,In_1053);
nor U1953 (N_1953,In_966,In_1402);
or U1954 (N_1954,In_719,In_1639);
nand U1955 (N_1955,In_1469,In_613);
nand U1956 (N_1956,In_675,In_1751);
nand U1957 (N_1957,In_466,In_986);
nand U1958 (N_1958,In_1898,In_1250);
nor U1959 (N_1959,In_844,In_999);
nand U1960 (N_1960,In_204,In_1798);
or U1961 (N_1961,In_85,In_1680);
xnor U1962 (N_1962,In_1516,In_146);
nor U1963 (N_1963,In_106,In_335);
nor U1964 (N_1964,In_1390,In_464);
and U1965 (N_1965,In_1384,In_688);
nand U1966 (N_1966,In_826,In_805);
nor U1967 (N_1967,In_1123,In_1992);
or U1968 (N_1968,In_940,In_938);
or U1969 (N_1969,In_1932,In_1370);
or U1970 (N_1970,In_1440,In_200);
and U1971 (N_1971,In_1965,In_1960);
or U1972 (N_1972,In_1805,In_1164);
nor U1973 (N_1973,In_947,In_168);
and U1974 (N_1974,In_385,In_49);
and U1975 (N_1975,In_1229,In_375);
nor U1976 (N_1976,In_1776,In_1380);
nand U1977 (N_1977,In_595,In_749);
nor U1978 (N_1978,In_1399,In_236);
and U1979 (N_1979,In_606,In_892);
nand U1980 (N_1980,In_1724,In_1423);
nand U1981 (N_1981,In_889,In_1256);
nand U1982 (N_1982,In_229,In_1176);
and U1983 (N_1983,In_1338,In_174);
or U1984 (N_1984,In_340,In_69);
and U1985 (N_1985,In_852,In_1366);
nor U1986 (N_1986,In_1192,In_681);
and U1987 (N_1987,In_59,In_1850);
and U1988 (N_1988,In_882,In_662);
and U1989 (N_1989,In_1674,In_75);
nand U1990 (N_1990,In_1284,In_1460);
or U1991 (N_1991,In_806,In_230);
nand U1992 (N_1992,In_590,In_1408);
or U1993 (N_1993,In_577,In_1123);
and U1994 (N_1994,In_151,In_338);
and U1995 (N_1995,In_118,In_378);
or U1996 (N_1996,In_1571,In_396);
nand U1997 (N_1997,In_345,In_1332);
nor U1998 (N_1998,In_743,In_589);
nor U1999 (N_1999,In_468,In_1319);
or U2000 (N_2000,In_1436,In_332);
nand U2001 (N_2001,In_1417,In_1507);
and U2002 (N_2002,In_309,In_1418);
nand U2003 (N_2003,In_1182,In_1063);
or U2004 (N_2004,In_1114,In_1970);
and U2005 (N_2005,In_1524,In_1326);
nor U2006 (N_2006,In_1913,In_843);
nand U2007 (N_2007,In_1188,In_546);
nor U2008 (N_2008,In_121,In_1579);
and U2009 (N_2009,In_450,In_1755);
and U2010 (N_2010,In_1110,In_709);
or U2011 (N_2011,In_1454,In_472);
nand U2012 (N_2012,In_1022,In_1040);
or U2013 (N_2013,In_1899,In_1924);
or U2014 (N_2014,In_1929,In_383);
nand U2015 (N_2015,In_939,In_1127);
nand U2016 (N_2016,In_225,In_919);
or U2017 (N_2017,In_1575,In_1258);
nand U2018 (N_2018,In_1128,In_1788);
and U2019 (N_2019,In_594,In_981);
and U2020 (N_2020,In_506,In_1755);
or U2021 (N_2021,In_1710,In_888);
and U2022 (N_2022,In_576,In_1806);
nand U2023 (N_2023,In_155,In_212);
and U2024 (N_2024,In_606,In_563);
nor U2025 (N_2025,In_517,In_1840);
and U2026 (N_2026,In_1650,In_1557);
and U2027 (N_2027,In_910,In_1337);
nand U2028 (N_2028,In_1786,In_686);
nand U2029 (N_2029,In_627,In_1578);
or U2030 (N_2030,In_1470,In_1510);
nor U2031 (N_2031,In_440,In_99);
nand U2032 (N_2032,In_1882,In_1778);
and U2033 (N_2033,In_474,In_54);
or U2034 (N_2034,In_968,In_1326);
and U2035 (N_2035,In_829,In_1228);
nand U2036 (N_2036,In_1336,In_627);
nor U2037 (N_2037,In_790,In_137);
or U2038 (N_2038,In_427,In_1792);
or U2039 (N_2039,In_1075,In_1325);
and U2040 (N_2040,In_1852,In_832);
and U2041 (N_2041,In_1600,In_636);
nor U2042 (N_2042,In_451,In_585);
and U2043 (N_2043,In_621,In_326);
or U2044 (N_2044,In_984,In_485);
and U2045 (N_2045,In_1194,In_1474);
or U2046 (N_2046,In_484,In_752);
and U2047 (N_2047,In_1241,In_850);
nor U2048 (N_2048,In_732,In_564);
nor U2049 (N_2049,In_1468,In_1855);
nor U2050 (N_2050,In_1641,In_1866);
nor U2051 (N_2051,In_1019,In_1983);
nor U2052 (N_2052,In_533,In_607);
and U2053 (N_2053,In_1392,In_1535);
nand U2054 (N_2054,In_163,In_1028);
nor U2055 (N_2055,In_150,In_1907);
or U2056 (N_2056,In_1317,In_1962);
and U2057 (N_2057,In_356,In_1133);
or U2058 (N_2058,In_411,In_426);
nand U2059 (N_2059,In_379,In_1511);
and U2060 (N_2060,In_1216,In_356);
or U2061 (N_2061,In_445,In_1603);
nand U2062 (N_2062,In_1197,In_358);
or U2063 (N_2063,In_82,In_1159);
nor U2064 (N_2064,In_1762,In_1743);
or U2065 (N_2065,In_424,In_415);
nor U2066 (N_2066,In_762,In_291);
and U2067 (N_2067,In_1443,In_168);
and U2068 (N_2068,In_502,In_1233);
nor U2069 (N_2069,In_1695,In_324);
or U2070 (N_2070,In_936,In_537);
and U2071 (N_2071,In_319,In_371);
and U2072 (N_2072,In_1456,In_68);
and U2073 (N_2073,In_283,In_1871);
or U2074 (N_2074,In_1972,In_246);
and U2075 (N_2075,In_1496,In_272);
nor U2076 (N_2076,In_593,In_904);
nor U2077 (N_2077,In_1224,In_716);
nand U2078 (N_2078,In_555,In_1964);
and U2079 (N_2079,In_160,In_366);
or U2080 (N_2080,In_1452,In_1128);
or U2081 (N_2081,In_1434,In_462);
nor U2082 (N_2082,In_1564,In_248);
and U2083 (N_2083,In_1016,In_1410);
nand U2084 (N_2084,In_1620,In_647);
xnor U2085 (N_2085,In_1537,In_1040);
nand U2086 (N_2086,In_73,In_841);
or U2087 (N_2087,In_581,In_1113);
nor U2088 (N_2088,In_53,In_301);
nand U2089 (N_2089,In_534,In_114);
nand U2090 (N_2090,In_1576,In_698);
nor U2091 (N_2091,In_612,In_1837);
or U2092 (N_2092,In_1525,In_1219);
nand U2093 (N_2093,In_52,In_1281);
or U2094 (N_2094,In_576,In_1836);
or U2095 (N_2095,In_885,In_19);
and U2096 (N_2096,In_1167,In_1886);
or U2097 (N_2097,In_562,In_183);
nand U2098 (N_2098,In_1204,In_573);
nor U2099 (N_2099,In_1081,In_1431);
nand U2100 (N_2100,In_57,In_1429);
or U2101 (N_2101,In_1774,In_1279);
or U2102 (N_2102,In_1443,In_818);
and U2103 (N_2103,In_1894,In_1231);
nand U2104 (N_2104,In_1417,In_1278);
nand U2105 (N_2105,In_519,In_578);
and U2106 (N_2106,In_1968,In_896);
nand U2107 (N_2107,In_56,In_885);
or U2108 (N_2108,In_573,In_485);
and U2109 (N_2109,In_260,In_1379);
and U2110 (N_2110,In_224,In_1392);
nand U2111 (N_2111,In_1907,In_1797);
or U2112 (N_2112,In_1336,In_1207);
nor U2113 (N_2113,In_1642,In_94);
or U2114 (N_2114,In_916,In_1987);
nand U2115 (N_2115,In_1843,In_1127);
and U2116 (N_2116,In_542,In_886);
nor U2117 (N_2117,In_1969,In_279);
and U2118 (N_2118,In_1518,In_926);
and U2119 (N_2119,In_395,In_1529);
nand U2120 (N_2120,In_1027,In_921);
or U2121 (N_2121,In_115,In_1231);
or U2122 (N_2122,In_1404,In_1464);
nand U2123 (N_2123,In_238,In_94);
nand U2124 (N_2124,In_1925,In_116);
and U2125 (N_2125,In_785,In_697);
nand U2126 (N_2126,In_128,In_230);
and U2127 (N_2127,In_727,In_499);
nor U2128 (N_2128,In_1294,In_175);
and U2129 (N_2129,In_1414,In_1386);
nand U2130 (N_2130,In_269,In_754);
nand U2131 (N_2131,In_8,In_729);
and U2132 (N_2132,In_876,In_888);
and U2133 (N_2133,In_181,In_1098);
and U2134 (N_2134,In_245,In_1158);
and U2135 (N_2135,In_1401,In_1762);
and U2136 (N_2136,In_1710,In_710);
and U2137 (N_2137,In_1297,In_1523);
xor U2138 (N_2138,In_1317,In_1873);
nand U2139 (N_2139,In_712,In_1515);
or U2140 (N_2140,In_22,In_884);
nor U2141 (N_2141,In_1112,In_1757);
and U2142 (N_2142,In_1669,In_1809);
nand U2143 (N_2143,In_1273,In_246);
or U2144 (N_2144,In_1084,In_1559);
nor U2145 (N_2145,In_649,In_1098);
nand U2146 (N_2146,In_1082,In_1360);
or U2147 (N_2147,In_1872,In_869);
and U2148 (N_2148,In_879,In_1849);
or U2149 (N_2149,In_375,In_1962);
nand U2150 (N_2150,In_1150,In_87);
and U2151 (N_2151,In_1471,In_408);
or U2152 (N_2152,In_752,In_1661);
nand U2153 (N_2153,In_1055,In_664);
nor U2154 (N_2154,In_1494,In_248);
and U2155 (N_2155,In_1746,In_371);
or U2156 (N_2156,In_1781,In_1992);
nor U2157 (N_2157,In_1481,In_1518);
nor U2158 (N_2158,In_850,In_1930);
xnor U2159 (N_2159,In_1775,In_629);
and U2160 (N_2160,In_108,In_239);
or U2161 (N_2161,In_777,In_1834);
or U2162 (N_2162,In_885,In_934);
nor U2163 (N_2163,In_892,In_1359);
nor U2164 (N_2164,In_887,In_19);
and U2165 (N_2165,In_343,In_1018);
and U2166 (N_2166,In_1149,In_1588);
and U2167 (N_2167,In_1842,In_439);
xnor U2168 (N_2168,In_1786,In_1109);
or U2169 (N_2169,In_1146,In_879);
nor U2170 (N_2170,In_1966,In_1060);
nor U2171 (N_2171,In_1946,In_845);
and U2172 (N_2172,In_1606,In_1761);
and U2173 (N_2173,In_1956,In_1844);
nor U2174 (N_2174,In_175,In_977);
nor U2175 (N_2175,In_1135,In_1440);
nor U2176 (N_2176,In_1532,In_1283);
and U2177 (N_2177,In_1112,In_885);
or U2178 (N_2178,In_937,In_1405);
nor U2179 (N_2179,In_491,In_1585);
xnor U2180 (N_2180,In_970,In_1718);
nand U2181 (N_2181,In_1369,In_380);
or U2182 (N_2182,In_891,In_1077);
nand U2183 (N_2183,In_1584,In_1408);
or U2184 (N_2184,In_1775,In_1999);
nor U2185 (N_2185,In_791,In_198);
and U2186 (N_2186,In_1112,In_270);
xor U2187 (N_2187,In_925,In_1858);
or U2188 (N_2188,In_1165,In_1422);
nand U2189 (N_2189,In_1142,In_1867);
nor U2190 (N_2190,In_514,In_1003);
and U2191 (N_2191,In_1850,In_1737);
nand U2192 (N_2192,In_43,In_430);
and U2193 (N_2193,In_1225,In_650);
nor U2194 (N_2194,In_1721,In_424);
and U2195 (N_2195,In_930,In_1341);
nor U2196 (N_2196,In_1547,In_622);
nor U2197 (N_2197,In_267,In_389);
and U2198 (N_2198,In_1035,In_392);
nand U2199 (N_2199,In_600,In_37);
or U2200 (N_2200,In_1464,In_1356);
or U2201 (N_2201,In_1746,In_36);
or U2202 (N_2202,In_352,In_369);
xor U2203 (N_2203,In_1131,In_1442);
nor U2204 (N_2204,In_926,In_1012);
or U2205 (N_2205,In_485,In_702);
or U2206 (N_2206,In_1527,In_1707);
and U2207 (N_2207,In_738,In_328);
or U2208 (N_2208,In_27,In_278);
and U2209 (N_2209,In_644,In_1241);
or U2210 (N_2210,In_1115,In_1931);
nor U2211 (N_2211,In_452,In_996);
and U2212 (N_2212,In_1095,In_1513);
or U2213 (N_2213,In_1389,In_1585);
and U2214 (N_2214,In_1227,In_110);
and U2215 (N_2215,In_709,In_1157);
nand U2216 (N_2216,In_988,In_968);
or U2217 (N_2217,In_1808,In_958);
nand U2218 (N_2218,In_1181,In_1126);
nand U2219 (N_2219,In_1990,In_1377);
and U2220 (N_2220,In_1221,In_1684);
or U2221 (N_2221,In_992,In_283);
nor U2222 (N_2222,In_1965,In_784);
nor U2223 (N_2223,In_1056,In_950);
and U2224 (N_2224,In_487,In_1281);
nor U2225 (N_2225,In_1521,In_104);
nor U2226 (N_2226,In_241,In_1329);
or U2227 (N_2227,In_272,In_1702);
nor U2228 (N_2228,In_1743,In_976);
nand U2229 (N_2229,In_40,In_110);
or U2230 (N_2230,In_1937,In_863);
nor U2231 (N_2231,In_1077,In_255);
and U2232 (N_2232,In_1134,In_1949);
or U2233 (N_2233,In_1048,In_1649);
and U2234 (N_2234,In_1888,In_1792);
or U2235 (N_2235,In_610,In_911);
nor U2236 (N_2236,In_1573,In_707);
and U2237 (N_2237,In_1116,In_1782);
nand U2238 (N_2238,In_777,In_1683);
nand U2239 (N_2239,In_630,In_1531);
and U2240 (N_2240,In_1158,In_1865);
xor U2241 (N_2241,In_836,In_817);
nand U2242 (N_2242,In_271,In_1821);
or U2243 (N_2243,In_600,In_833);
nand U2244 (N_2244,In_1766,In_1040);
or U2245 (N_2245,In_12,In_1363);
or U2246 (N_2246,In_1685,In_1162);
or U2247 (N_2247,In_1678,In_362);
or U2248 (N_2248,In_1582,In_1371);
nand U2249 (N_2249,In_924,In_388);
nand U2250 (N_2250,In_276,In_1789);
nor U2251 (N_2251,In_535,In_750);
and U2252 (N_2252,In_850,In_890);
and U2253 (N_2253,In_1408,In_39);
or U2254 (N_2254,In_14,In_923);
nor U2255 (N_2255,In_1948,In_16);
and U2256 (N_2256,In_783,In_1042);
nand U2257 (N_2257,In_1370,In_1484);
nor U2258 (N_2258,In_71,In_1385);
or U2259 (N_2259,In_1166,In_1460);
and U2260 (N_2260,In_892,In_1760);
nor U2261 (N_2261,In_1727,In_1307);
nand U2262 (N_2262,In_755,In_116);
nor U2263 (N_2263,In_491,In_348);
nand U2264 (N_2264,In_1968,In_496);
nand U2265 (N_2265,In_561,In_318);
nor U2266 (N_2266,In_615,In_1022);
or U2267 (N_2267,In_1474,In_575);
nand U2268 (N_2268,In_970,In_1280);
and U2269 (N_2269,In_354,In_1208);
or U2270 (N_2270,In_166,In_460);
nand U2271 (N_2271,In_466,In_967);
nor U2272 (N_2272,In_393,In_275);
or U2273 (N_2273,In_1437,In_780);
nor U2274 (N_2274,In_452,In_300);
nand U2275 (N_2275,In_851,In_1311);
xnor U2276 (N_2276,In_1504,In_1774);
and U2277 (N_2277,In_667,In_1908);
or U2278 (N_2278,In_994,In_302);
nor U2279 (N_2279,In_1703,In_956);
or U2280 (N_2280,In_1256,In_1694);
nor U2281 (N_2281,In_1200,In_177);
or U2282 (N_2282,In_1954,In_16);
and U2283 (N_2283,In_994,In_1237);
or U2284 (N_2284,In_184,In_435);
or U2285 (N_2285,In_727,In_1315);
and U2286 (N_2286,In_1424,In_174);
nor U2287 (N_2287,In_409,In_1698);
nor U2288 (N_2288,In_327,In_479);
nand U2289 (N_2289,In_623,In_748);
or U2290 (N_2290,In_1128,In_1333);
nor U2291 (N_2291,In_846,In_1666);
nor U2292 (N_2292,In_184,In_345);
and U2293 (N_2293,In_358,In_1395);
and U2294 (N_2294,In_1669,In_64);
nor U2295 (N_2295,In_8,In_480);
or U2296 (N_2296,In_1144,In_725);
nand U2297 (N_2297,In_1715,In_473);
nor U2298 (N_2298,In_138,In_657);
nor U2299 (N_2299,In_131,In_1852);
and U2300 (N_2300,In_1581,In_1795);
and U2301 (N_2301,In_1514,In_385);
nor U2302 (N_2302,In_880,In_1527);
nor U2303 (N_2303,In_1059,In_1336);
nor U2304 (N_2304,In_1605,In_1177);
xor U2305 (N_2305,In_1794,In_229);
and U2306 (N_2306,In_301,In_1411);
nor U2307 (N_2307,In_522,In_1074);
or U2308 (N_2308,In_1373,In_1287);
or U2309 (N_2309,In_101,In_383);
or U2310 (N_2310,In_500,In_1868);
and U2311 (N_2311,In_554,In_1370);
nand U2312 (N_2312,In_1745,In_869);
and U2313 (N_2313,In_731,In_1299);
nor U2314 (N_2314,In_1067,In_624);
nor U2315 (N_2315,In_6,In_106);
and U2316 (N_2316,In_415,In_1925);
or U2317 (N_2317,In_186,In_538);
and U2318 (N_2318,In_888,In_1452);
nand U2319 (N_2319,In_573,In_102);
nor U2320 (N_2320,In_1802,In_525);
nand U2321 (N_2321,In_1473,In_1587);
or U2322 (N_2322,In_1874,In_1305);
and U2323 (N_2323,In_196,In_762);
nand U2324 (N_2324,In_201,In_1161);
nand U2325 (N_2325,In_530,In_1066);
nand U2326 (N_2326,In_778,In_237);
nand U2327 (N_2327,In_714,In_584);
and U2328 (N_2328,In_1219,In_620);
nand U2329 (N_2329,In_958,In_571);
nand U2330 (N_2330,In_1777,In_836);
nor U2331 (N_2331,In_1222,In_335);
or U2332 (N_2332,In_1787,In_613);
and U2333 (N_2333,In_739,In_1012);
nor U2334 (N_2334,In_977,In_1363);
nand U2335 (N_2335,In_513,In_1045);
nor U2336 (N_2336,In_1361,In_1994);
nand U2337 (N_2337,In_1672,In_853);
or U2338 (N_2338,In_784,In_360);
and U2339 (N_2339,In_1269,In_1999);
xor U2340 (N_2340,In_927,In_1697);
nor U2341 (N_2341,In_1561,In_96);
and U2342 (N_2342,In_1079,In_105);
or U2343 (N_2343,In_1335,In_655);
xor U2344 (N_2344,In_1127,In_230);
nor U2345 (N_2345,In_1021,In_1105);
xnor U2346 (N_2346,In_531,In_1189);
or U2347 (N_2347,In_54,In_1698);
nand U2348 (N_2348,In_1098,In_997);
and U2349 (N_2349,In_1009,In_1875);
and U2350 (N_2350,In_257,In_1922);
nand U2351 (N_2351,In_1585,In_1751);
and U2352 (N_2352,In_1894,In_1124);
nand U2353 (N_2353,In_1924,In_1828);
nand U2354 (N_2354,In_1708,In_427);
or U2355 (N_2355,In_878,In_1864);
or U2356 (N_2356,In_218,In_1455);
or U2357 (N_2357,In_1638,In_1835);
nor U2358 (N_2358,In_150,In_1399);
and U2359 (N_2359,In_848,In_1683);
nor U2360 (N_2360,In_1924,In_630);
xor U2361 (N_2361,In_1673,In_395);
nand U2362 (N_2362,In_1921,In_1867);
xnor U2363 (N_2363,In_301,In_970);
and U2364 (N_2364,In_1353,In_220);
nand U2365 (N_2365,In_1544,In_1193);
nand U2366 (N_2366,In_33,In_588);
nand U2367 (N_2367,In_1794,In_716);
nand U2368 (N_2368,In_14,In_428);
nand U2369 (N_2369,In_143,In_44);
nand U2370 (N_2370,In_986,In_151);
and U2371 (N_2371,In_622,In_282);
nor U2372 (N_2372,In_1946,In_85);
and U2373 (N_2373,In_1774,In_1489);
or U2374 (N_2374,In_1413,In_1700);
and U2375 (N_2375,In_132,In_1778);
and U2376 (N_2376,In_1781,In_195);
xnor U2377 (N_2377,In_1451,In_1697);
or U2378 (N_2378,In_1938,In_1775);
nand U2379 (N_2379,In_1069,In_65);
xor U2380 (N_2380,In_17,In_1792);
or U2381 (N_2381,In_852,In_778);
nor U2382 (N_2382,In_311,In_1698);
nand U2383 (N_2383,In_1721,In_187);
or U2384 (N_2384,In_1364,In_1185);
and U2385 (N_2385,In_1675,In_650);
or U2386 (N_2386,In_834,In_1207);
nor U2387 (N_2387,In_645,In_119);
and U2388 (N_2388,In_1607,In_91);
nand U2389 (N_2389,In_1275,In_903);
and U2390 (N_2390,In_918,In_937);
nand U2391 (N_2391,In_437,In_344);
nand U2392 (N_2392,In_1070,In_941);
and U2393 (N_2393,In_515,In_1799);
nand U2394 (N_2394,In_1166,In_253);
nor U2395 (N_2395,In_255,In_776);
and U2396 (N_2396,In_888,In_424);
and U2397 (N_2397,In_1138,In_1668);
or U2398 (N_2398,In_774,In_1207);
nor U2399 (N_2399,In_1688,In_864);
and U2400 (N_2400,In_1925,In_21);
nand U2401 (N_2401,In_1703,In_1655);
and U2402 (N_2402,In_1995,In_143);
nor U2403 (N_2403,In_1211,In_787);
nor U2404 (N_2404,In_323,In_967);
nand U2405 (N_2405,In_1549,In_1460);
nand U2406 (N_2406,In_816,In_1473);
nor U2407 (N_2407,In_884,In_876);
nor U2408 (N_2408,In_1581,In_629);
nand U2409 (N_2409,In_115,In_1167);
nand U2410 (N_2410,In_70,In_1391);
or U2411 (N_2411,In_1649,In_1640);
nor U2412 (N_2412,In_1248,In_942);
nor U2413 (N_2413,In_1868,In_1704);
and U2414 (N_2414,In_298,In_1686);
or U2415 (N_2415,In_1796,In_1849);
nor U2416 (N_2416,In_544,In_1166);
nand U2417 (N_2417,In_1490,In_814);
nand U2418 (N_2418,In_351,In_1664);
nand U2419 (N_2419,In_676,In_1687);
or U2420 (N_2420,In_790,In_913);
nor U2421 (N_2421,In_73,In_416);
nand U2422 (N_2422,In_1276,In_1737);
or U2423 (N_2423,In_1634,In_943);
nand U2424 (N_2424,In_1446,In_1532);
nor U2425 (N_2425,In_1465,In_104);
or U2426 (N_2426,In_11,In_1398);
or U2427 (N_2427,In_1114,In_1403);
nand U2428 (N_2428,In_148,In_19);
nor U2429 (N_2429,In_1892,In_226);
or U2430 (N_2430,In_1267,In_73);
nand U2431 (N_2431,In_1761,In_1446);
or U2432 (N_2432,In_938,In_1839);
and U2433 (N_2433,In_1529,In_1013);
or U2434 (N_2434,In_953,In_1918);
or U2435 (N_2435,In_1210,In_1234);
or U2436 (N_2436,In_30,In_742);
or U2437 (N_2437,In_93,In_546);
and U2438 (N_2438,In_1046,In_914);
and U2439 (N_2439,In_1445,In_220);
nand U2440 (N_2440,In_583,In_901);
nand U2441 (N_2441,In_1805,In_279);
and U2442 (N_2442,In_653,In_428);
nor U2443 (N_2443,In_1824,In_590);
or U2444 (N_2444,In_205,In_1779);
and U2445 (N_2445,In_1898,In_565);
or U2446 (N_2446,In_191,In_1246);
nor U2447 (N_2447,In_895,In_70);
and U2448 (N_2448,In_1467,In_317);
or U2449 (N_2449,In_1984,In_1143);
nand U2450 (N_2450,In_1858,In_230);
nand U2451 (N_2451,In_1846,In_66);
or U2452 (N_2452,In_1627,In_1084);
nor U2453 (N_2453,In_1728,In_495);
and U2454 (N_2454,In_1295,In_976);
or U2455 (N_2455,In_641,In_451);
nor U2456 (N_2456,In_579,In_468);
and U2457 (N_2457,In_1779,In_544);
nand U2458 (N_2458,In_951,In_476);
nand U2459 (N_2459,In_1312,In_1692);
nor U2460 (N_2460,In_959,In_1006);
nand U2461 (N_2461,In_1532,In_468);
and U2462 (N_2462,In_1924,In_370);
or U2463 (N_2463,In_1439,In_1237);
nor U2464 (N_2464,In_1544,In_5);
nand U2465 (N_2465,In_294,In_1449);
xor U2466 (N_2466,In_618,In_127);
nor U2467 (N_2467,In_1132,In_497);
and U2468 (N_2468,In_1442,In_655);
or U2469 (N_2469,In_434,In_120);
or U2470 (N_2470,In_165,In_340);
nor U2471 (N_2471,In_1623,In_1522);
and U2472 (N_2472,In_320,In_541);
nor U2473 (N_2473,In_754,In_270);
and U2474 (N_2474,In_1245,In_959);
and U2475 (N_2475,In_1743,In_274);
xor U2476 (N_2476,In_686,In_1898);
nand U2477 (N_2477,In_749,In_1487);
nand U2478 (N_2478,In_1608,In_488);
nor U2479 (N_2479,In_1927,In_1892);
nand U2480 (N_2480,In_793,In_230);
nor U2481 (N_2481,In_1896,In_1470);
nor U2482 (N_2482,In_657,In_1876);
and U2483 (N_2483,In_1219,In_1227);
nand U2484 (N_2484,In_1208,In_1356);
and U2485 (N_2485,In_190,In_321);
and U2486 (N_2486,In_635,In_401);
nand U2487 (N_2487,In_649,In_1468);
nand U2488 (N_2488,In_1746,In_874);
nor U2489 (N_2489,In_724,In_953);
or U2490 (N_2490,In_1217,In_1411);
xnor U2491 (N_2491,In_1599,In_709);
and U2492 (N_2492,In_42,In_871);
and U2493 (N_2493,In_1343,In_1202);
and U2494 (N_2494,In_1571,In_736);
nand U2495 (N_2495,In_968,In_1496);
and U2496 (N_2496,In_1655,In_1474);
and U2497 (N_2497,In_1429,In_319);
nand U2498 (N_2498,In_633,In_1173);
nor U2499 (N_2499,In_768,In_652);
and U2500 (N_2500,In_1795,In_367);
or U2501 (N_2501,In_1594,In_1718);
nor U2502 (N_2502,In_1454,In_1677);
nand U2503 (N_2503,In_1707,In_124);
and U2504 (N_2504,In_1901,In_1451);
xor U2505 (N_2505,In_1931,In_127);
nor U2506 (N_2506,In_760,In_297);
or U2507 (N_2507,In_1868,In_605);
or U2508 (N_2508,In_1292,In_484);
or U2509 (N_2509,In_1951,In_429);
or U2510 (N_2510,In_1589,In_640);
or U2511 (N_2511,In_1296,In_1570);
and U2512 (N_2512,In_360,In_1825);
or U2513 (N_2513,In_1040,In_285);
and U2514 (N_2514,In_1297,In_416);
and U2515 (N_2515,In_114,In_560);
nor U2516 (N_2516,In_1859,In_1125);
and U2517 (N_2517,In_1036,In_46);
and U2518 (N_2518,In_815,In_128);
nor U2519 (N_2519,In_1408,In_250);
nand U2520 (N_2520,In_53,In_146);
or U2521 (N_2521,In_1096,In_1708);
nand U2522 (N_2522,In_764,In_1447);
and U2523 (N_2523,In_170,In_1453);
and U2524 (N_2524,In_1484,In_40);
nand U2525 (N_2525,In_1573,In_1871);
nand U2526 (N_2526,In_383,In_1999);
nor U2527 (N_2527,In_1833,In_794);
nor U2528 (N_2528,In_780,In_1029);
xor U2529 (N_2529,In_718,In_1800);
nor U2530 (N_2530,In_879,In_1624);
or U2531 (N_2531,In_1044,In_726);
and U2532 (N_2532,In_116,In_1647);
nor U2533 (N_2533,In_1756,In_1845);
or U2534 (N_2534,In_388,In_986);
nor U2535 (N_2535,In_1196,In_1711);
nor U2536 (N_2536,In_79,In_1236);
nand U2537 (N_2537,In_1315,In_963);
or U2538 (N_2538,In_322,In_146);
nor U2539 (N_2539,In_1199,In_1765);
and U2540 (N_2540,In_1832,In_457);
nor U2541 (N_2541,In_87,In_1371);
xor U2542 (N_2542,In_1341,In_699);
and U2543 (N_2543,In_602,In_776);
nor U2544 (N_2544,In_1406,In_204);
nor U2545 (N_2545,In_988,In_406);
nand U2546 (N_2546,In_1095,In_1129);
nand U2547 (N_2547,In_98,In_124);
or U2548 (N_2548,In_1633,In_411);
and U2549 (N_2549,In_254,In_1162);
and U2550 (N_2550,In_819,In_151);
and U2551 (N_2551,In_622,In_1108);
nand U2552 (N_2552,In_1924,In_1637);
nand U2553 (N_2553,In_21,In_450);
and U2554 (N_2554,In_1144,In_1281);
or U2555 (N_2555,In_1504,In_666);
nor U2556 (N_2556,In_1663,In_679);
or U2557 (N_2557,In_884,In_466);
nor U2558 (N_2558,In_1126,In_1577);
and U2559 (N_2559,In_1251,In_1383);
nor U2560 (N_2560,In_577,In_1591);
nand U2561 (N_2561,In_1389,In_1797);
and U2562 (N_2562,In_1076,In_148);
and U2563 (N_2563,In_65,In_445);
nand U2564 (N_2564,In_720,In_1460);
nand U2565 (N_2565,In_303,In_1916);
nand U2566 (N_2566,In_1398,In_1586);
or U2567 (N_2567,In_183,In_237);
nand U2568 (N_2568,In_1969,In_1496);
and U2569 (N_2569,In_1754,In_837);
nor U2570 (N_2570,In_225,In_1270);
nor U2571 (N_2571,In_1643,In_1826);
nor U2572 (N_2572,In_1240,In_1731);
nand U2573 (N_2573,In_1563,In_1170);
nand U2574 (N_2574,In_1985,In_439);
and U2575 (N_2575,In_438,In_1878);
nor U2576 (N_2576,In_906,In_643);
and U2577 (N_2577,In_1746,In_167);
or U2578 (N_2578,In_1914,In_53);
or U2579 (N_2579,In_945,In_384);
and U2580 (N_2580,In_330,In_713);
or U2581 (N_2581,In_1605,In_76);
xnor U2582 (N_2582,In_1379,In_782);
nand U2583 (N_2583,In_1777,In_1007);
nand U2584 (N_2584,In_1520,In_263);
nand U2585 (N_2585,In_1409,In_988);
or U2586 (N_2586,In_226,In_1463);
nand U2587 (N_2587,In_1266,In_156);
nor U2588 (N_2588,In_680,In_795);
nor U2589 (N_2589,In_1168,In_1472);
nor U2590 (N_2590,In_24,In_1650);
nand U2591 (N_2591,In_956,In_86);
nor U2592 (N_2592,In_959,In_13);
or U2593 (N_2593,In_1323,In_446);
nand U2594 (N_2594,In_708,In_403);
and U2595 (N_2595,In_285,In_1726);
and U2596 (N_2596,In_775,In_784);
nor U2597 (N_2597,In_415,In_1444);
and U2598 (N_2598,In_1908,In_1206);
nor U2599 (N_2599,In_33,In_751);
nor U2600 (N_2600,In_413,In_1677);
or U2601 (N_2601,In_348,In_818);
nor U2602 (N_2602,In_1307,In_40);
and U2603 (N_2603,In_481,In_1720);
or U2604 (N_2604,In_1381,In_1411);
or U2605 (N_2605,In_1317,In_1094);
and U2606 (N_2606,In_1238,In_949);
nor U2607 (N_2607,In_127,In_1689);
or U2608 (N_2608,In_1912,In_1819);
nor U2609 (N_2609,In_309,In_1515);
and U2610 (N_2610,In_1917,In_1484);
and U2611 (N_2611,In_1511,In_1953);
nor U2612 (N_2612,In_215,In_270);
or U2613 (N_2613,In_1438,In_751);
nand U2614 (N_2614,In_1628,In_692);
and U2615 (N_2615,In_668,In_130);
nand U2616 (N_2616,In_1742,In_1761);
or U2617 (N_2617,In_1050,In_1483);
nor U2618 (N_2618,In_1095,In_1952);
nor U2619 (N_2619,In_1685,In_820);
or U2620 (N_2620,In_1609,In_1032);
and U2621 (N_2621,In_293,In_1380);
nand U2622 (N_2622,In_1537,In_398);
nor U2623 (N_2623,In_629,In_1397);
or U2624 (N_2624,In_1980,In_1599);
and U2625 (N_2625,In_1091,In_1065);
and U2626 (N_2626,In_1156,In_1293);
or U2627 (N_2627,In_673,In_478);
nor U2628 (N_2628,In_328,In_369);
and U2629 (N_2629,In_1955,In_595);
or U2630 (N_2630,In_662,In_1755);
or U2631 (N_2631,In_1079,In_123);
nor U2632 (N_2632,In_1992,In_723);
or U2633 (N_2633,In_1655,In_1478);
and U2634 (N_2634,In_812,In_317);
nand U2635 (N_2635,In_1051,In_857);
nand U2636 (N_2636,In_562,In_1432);
nand U2637 (N_2637,In_1159,In_155);
and U2638 (N_2638,In_760,In_1926);
nand U2639 (N_2639,In_791,In_1934);
and U2640 (N_2640,In_759,In_870);
nor U2641 (N_2641,In_117,In_1062);
nand U2642 (N_2642,In_291,In_1180);
nand U2643 (N_2643,In_1846,In_1874);
and U2644 (N_2644,In_1635,In_393);
nor U2645 (N_2645,In_1102,In_50);
or U2646 (N_2646,In_1557,In_1068);
nand U2647 (N_2647,In_408,In_624);
nor U2648 (N_2648,In_33,In_573);
nor U2649 (N_2649,In_1778,In_1903);
or U2650 (N_2650,In_1573,In_1308);
or U2651 (N_2651,In_1734,In_1964);
and U2652 (N_2652,In_116,In_548);
and U2653 (N_2653,In_815,In_1765);
nand U2654 (N_2654,In_176,In_45);
and U2655 (N_2655,In_1953,In_55);
and U2656 (N_2656,In_928,In_595);
nand U2657 (N_2657,In_1413,In_1232);
nor U2658 (N_2658,In_1409,In_1743);
and U2659 (N_2659,In_1001,In_113);
and U2660 (N_2660,In_1261,In_1270);
nor U2661 (N_2661,In_1840,In_1875);
and U2662 (N_2662,In_588,In_613);
nor U2663 (N_2663,In_1224,In_227);
nand U2664 (N_2664,In_715,In_1139);
and U2665 (N_2665,In_1189,In_1811);
and U2666 (N_2666,In_1315,In_918);
and U2667 (N_2667,In_1181,In_1644);
nand U2668 (N_2668,In_1602,In_1686);
nand U2669 (N_2669,In_1099,In_835);
and U2670 (N_2670,In_305,In_1655);
nand U2671 (N_2671,In_712,In_1215);
or U2672 (N_2672,In_928,In_183);
nand U2673 (N_2673,In_1589,In_937);
and U2674 (N_2674,In_196,In_1857);
nor U2675 (N_2675,In_274,In_272);
nor U2676 (N_2676,In_1870,In_1865);
nand U2677 (N_2677,In_833,In_1646);
and U2678 (N_2678,In_1139,In_727);
or U2679 (N_2679,In_105,In_1082);
nor U2680 (N_2680,In_1630,In_688);
and U2681 (N_2681,In_1030,In_1966);
nor U2682 (N_2682,In_768,In_1159);
or U2683 (N_2683,In_1631,In_1970);
and U2684 (N_2684,In_548,In_1910);
xor U2685 (N_2685,In_537,In_294);
or U2686 (N_2686,In_1172,In_126);
nor U2687 (N_2687,In_1206,In_1134);
nor U2688 (N_2688,In_511,In_408);
and U2689 (N_2689,In_1343,In_117);
and U2690 (N_2690,In_894,In_1752);
and U2691 (N_2691,In_1398,In_1566);
xor U2692 (N_2692,In_1461,In_1342);
nand U2693 (N_2693,In_128,In_927);
or U2694 (N_2694,In_392,In_1913);
xnor U2695 (N_2695,In_1058,In_493);
nand U2696 (N_2696,In_748,In_947);
nand U2697 (N_2697,In_1924,In_1809);
nand U2698 (N_2698,In_1787,In_1203);
or U2699 (N_2699,In_1645,In_615);
nor U2700 (N_2700,In_836,In_519);
nor U2701 (N_2701,In_1941,In_1186);
and U2702 (N_2702,In_882,In_1549);
nor U2703 (N_2703,In_1979,In_1009);
nor U2704 (N_2704,In_786,In_518);
or U2705 (N_2705,In_839,In_1153);
nand U2706 (N_2706,In_370,In_1599);
nor U2707 (N_2707,In_470,In_1470);
or U2708 (N_2708,In_1273,In_1203);
nor U2709 (N_2709,In_150,In_1850);
and U2710 (N_2710,In_11,In_1976);
and U2711 (N_2711,In_1598,In_1846);
nand U2712 (N_2712,In_1196,In_1511);
or U2713 (N_2713,In_894,In_1337);
or U2714 (N_2714,In_790,In_1247);
and U2715 (N_2715,In_634,In_1136);
or U2716 (N_2716,In_96,In_760);
or U2717 (N_2717,In_315,In_1641);
or U2718 (N_2718,In_299,In_1186);
nor U2719 (N_2719,In_1695,In_1493);
or U2720 (N_2720,In_1650,In_1239);
nor U2721 (N_2721,In_1036,In_149);
xor U2722 (N_2722,In_1821,In_1908);
nor U2723 (N_2723,In_1988,In_450);
and U2724 (N_2724,In_1867,In_1914);
and U2725 (N_2725,In_615,In_229);
nand U2726 (N_2726,In_1492,In_1792);
or U2727 (N_2727,In_1923,In_1332);
or U2728 (N_2728,In_1595,In_1896);
nand U2729 (N_2729,In_610,In_73);
and U2730 (N_2730,In_1946,In_1486);
nand U2731 (N_2731,In_483,In_256);
or U2732 (N_2732,In_1390,In_1598);
nand U2733 (N_2733,In_423,In_1465);
and U2734 (N_2734,In_1106,In_1796);
or U2735 (N_2735,In_704,In_1113);
nand U2736 (N_2736,In_694,In_970);
or U2737 (N_2737,In_1151,In_419);
nand U2738 (N_2738,In_1517,In_300);
nor U2739 (N_2739,In_586,In_230);
nor U2740 (N_2740,In_622,In_1058);
nand U2741 (N_2741,In_892,In_1699);
and U2742 (N_2742,In_1858,In_200);
nand U2743 (N_2743,In_1415,In_878);
and U2744 (N_2744,In_518,In_1991);
or U2745 (N_2745,In_1266,In_859);
nand U2746 (N_2746,In_1900,In_1722);
or U2747 (N_2747,In_639,In_59);
xor U2748 (N_2748,In_1281,In_226);
nand U2749 (N_2749,In_1926,In_15);
and U2750 (N_2750,In_1623,In_128);
and U2751 (N_2751,In_1959,In_585);
and U2752 (N_2752,In_1573,In_1361);
or U2753 (N_2753,In_695,In_34);
and U2754 (N_2754,In_729,In_1784);
nor U2755 (N_2755,In_1261,In_1853);
and U2756 (N_2756,In_65,In_792);
xor U2757 (N_2757,In_1483,In_835);
nor U2758 (N_2758,In_756,In_1135);
nand U2759 (N_2759,In_1344,In_1007);
or U2760 (N_2760,In_358,In_470);
or U2761 (N_2761,In_1185,In_416);
nor U2762 (N_2762,In_396,In_975);
and U2763 (N_2763,In_893,In_1636);
or U2764 (N_2764,In_664,In_19);
nor U2765 (N_2765,In_1436,In_1136);
nor U2766 (N_2766,In_923,In_1140);
or U2767 (N_2767,In_764,In_1718);
nor U2768 (N_2768,In_1203,In_1471);
and U2769 (N_2769,In_853,In_323);
or U2770 (N_2770,In_1062,In_865);
nor U2771 (N_2771,In_747,In_280);
nor U2772 (N_2772,In_870,In_513);
xor U2773 (N_2773,In_1128,In_808);
nor U2774 (N_2774,In_1151,In_65);
or U2775 (N_2775,In_953,In_195);
nand U2776 (N_2776,In_537,In_1700);
nand U2777 (N_2777,In_1384,In_790);
and U2778 (N_2778,In_241,In_889);
or U2779 (N_2779,In_846,In_1392);
nand U2780 (N_2780,In_1316,In_1248);
nand U2781 (N_2781,In_296,In_1827);
nor U2782 (N_2782,In_1780,In_1879);
nor U2783 (N_2783,In_893,In_2);
nand U2784 (N_2784,In_1782,In_1139);
nor U2785 (N_2785,In_1226,In_1340);
nor U2786 (N_2786,In_1950,In_409);
and U2787 (N_2787,In_272,In_221);
nand U2788 (N_2788,In_781,In_34);
nand U2789 (N_2789,In_375,In_1119);
or U2790 (N_2790,In_1111,In_1115);
nand U2791 (N_2791,In_725,In_1064);
nor U2792 (N_2792,In_1651,In_1163);
nor U2793 (N_2793,In_892,In_690);
nand U2794 (N_2794,In_1842,In_823);
nor U2795 (N_2795,In_1486,In_1634);
and U2796 (N_2796,In_399,In_1792);
nor U2797 (N_2797,In_323,In_719);
and U2798 (N_2798,In_1464,In_1780);
nor U2799 (N_2799,In_366,In_1118);
nand U2800 (N_2800,In_131,In_1701);
nor U2801 (N_2801,In_1231,In_832);
or U2802 (N_2802,In_1973,In_1581);
and U2803 (N_2803,In_1102,In_198);
nand U2804 (N_2804,In_272,In_639);
and U2805 (N_2805,In_1787,In_952);
nor U2806 (N_2806,In_1166,In_1834);
or U2807 (N_2807,In_395,In_364);
nor U2808 (N_2808,In_760,In_1681);
nor U2809 (N_2809,In_972,In_410);
nand U2810 (N_2810,In_87,In_1992);
nor U2811 (N_2811,In_196,In_1816);
and U2812 (N_2812,In_1764,In_5);
and U2813 (N_2813,In_1456,In_191);
nand U2814 (N_2814,In_1629,In_739);
or U2815 (N_2815,In_997,In_1902);
nor U2816 (N_2816,In_1700,In_967);
and U2817 (N_2817,In_1662,In_1494);
or U2818 (N_2818,In_1844,In_1791);
nand U2819 (N_2819,In_1379,In_1455);
or U2820 (N_2820,In_1978,In_806);
nand U2821 (N_2821,In_954,In_925);
or U2822 (N_2822,In_185,In_1476);
nor U2823 (N_2823,In_595,In_1569);
nor U2824 (N_2824,In_1653,In_384);
and U2825 (N_2825,In_1299,In_656);
nor U2826 (N_2826,In_1137,In_1084);
or U2827 (N_2827,In_629,In_628);
or U2828 (N_2828,In_775,In_738);
and U2829 (N_2829,In_517,In_24);
and U2830 (N_2830,In_981,In_1474);
nand U2831 (N_2831,In_1189,In_1066);
and U2832 (N_2832,In_197,In_1252);
and U2833 (N_2833,In_1688,In_1906);
or U2834 (N_2834,In_339,In_163);
and U2835 (N_2835,In_135,In_1549);
nor U2836 (N_2836,In_221,In_95);
nor U2837 (N_2837,In_1482,In_1803);
nand U2838 (N_2838,In_1479,In_1754);
nand U2839 (N_2839,In_1720,In_1904);
nand U2840 (N_2840,In_1474,In_701);
nand U2841 (N_2841,In_654,In_1586);
or U2842 (N_2842,In_798,In_1070);
nor U2843 (N_2843,In_186,In_1409);
nand U2844 (N_2844,In_658,In_1952);
nor U2845 (N_2845,In_1641,In_480);
or U2846 (N_2846,In_1063,In_735);
nor U2847 (N_2847,In_885,In_1101);
nor U2848 (N_2848,In_1332,In_476);
nor U2849 (N_2849,In_1367,In_960);
nand U2850 (N_2850,In_698,In_234);
nand U2851 (N_2851,In_1823,In_1170);
xnor U2852 (N_2852,In_94,In_1654);
nand U2853 (N_2853,In_1588,In_250);
nand U2854 (N_2854,In_935,In_1732);
nor U2855 (N_2855,In_259,In_575);
or U2856 (N_2856,In_969,In_1762);
and U2857 (N_2857,In_1062,In_1856);
nand U2858 (N_2858,In_1567,In_1096);
and U2859 (N_2859,In_996,In_1891);
and U2860 (N_2860,In_79,In_1371);
nor U2861 (N_2861,In_1713,In_1493);
and U2862 (N_2862,In_1255,In_1432);
or U2863 (N_2863,In_760,In_632);
and U2864 (N_2864,In_552,In_439);
and U2865 (N_2865,In_1368,In_1282);
nand U2866 (N_2866,In_1128,In_20);
or U2867 (N_2867,In_354,In_532);
or U2868 (N_2868,In_1376,In_621);
nor U2869 (N_2869,In_1593,In_251);
nand U2870 (N_2870,In_1487,In_1072);
and U2871 (N_2871,In_1871,In_1872);
or U2872 (N_2872,In_377,In_350);
nand U2873 (N_2873,In_435,In_1311);
nor U2874 (N_2874,In_915,In_322);
nand U2875 (N_2875,In_1154,In_1883);
nand U2876 (N_2876,In_1493,In_144);
nor U2877 (N_2877,In_1056,In_770);
nor U2878 (N_2878,In_1074,In_1669);
nor U2879 (N_2879,In_188,In_856);
nand U2880 (N_2880,In_1096,In_22);
and U2881 (N_2881,In_934,In_1580);
and U2882 (N_2882,In_1964,In_522);
nand U2883 (N_2883,In_1789,In_873);
nor U2884 (N_2884,In_712,In_327);
and U2885 (N_2885,In_1176,In_766);
nand U2886 (N_2886,In_1615,In_849);
and U2887 (N_2887,In_695,In_1604);
or U2888 (N_2888,In_805,In_857);
nand U2889 (N_2889,In_1978,In_31);
and U2890 (N_2890,In_1777,In_368);
nand U2891 (N_2891,In_1570,In_1090);
or U2892 (N_2892,In_1360,In_681);
or U2893 (N_2893,In_724,In_1241);
nor U2894 (N_2894,In_1021,In_1578);
nand U2895 (N_2895,In_1710,In_1140);
or U2896 (N_2896,In_1242,In_811);
xor U2897 (N_2897,In_395,In_1024);
nor U2898 (N_2898,In_408,In_997);
nand U2899 (N_2899,In_29,In_1496);
or U2900 (N_2900,In_19,In_1990);
nand U2901 (N_2901,In_847,In_673);
or U2902 (N_2902,In_264,In_612);
or U2903 (N_2903,In_1659,In_933);
and U2904 (N_2904,In_1896,In_1916);
and U2905 (N_2905,In_1911,In_55);
or U2906 (N_2906,In_1166,In_1667);
or U2907 (N_2907,In_1406,In_437);
or U2908 (N_2908,In_786,In_172);
or U2909 (N_2909,In_1075,In_611);
or U2910 (N_2910,In_434,In_1985);
nor U2911 (N_2911,In_604,In_744);
nand U2912 (N_2912,In_1711,In_1107);
nor U2913 (N_2913,In_1865,In_167);
nand U2914 (N_2914,In_881,In_149);
xor U2915 (N_2915,In_518,In_1671);
or U2916 (N_2916,In_1261,In_154);
nand U2917 (N_2917,In_1986,In_56);
nand U2918 (N_2918,In_610,In_715);
or U2919 (N_2919,In_1097,In_1756);
or U2920 (N_2920,In_1293,In_645);
nand U2921 (N_2921,In_889,In_1627);
and U2922 (N_2922,In_1077,In_1487);
nor U2923 (N_2923,In_1008,In_1320);
nor U2924 (N_2924,In_398,In_1025);
or U2925 (N_2925,In_188,In_1937);
nand U2926 (N_2926,In_913,In_1907);
and U2927 (N_2927,In_1180,In_475);
and U2928 (N_2928,In_1493,In_145);
or U2929 (N_2929,In_430,In_1126);
and U2930 (N_2930,In_1743,In_378);
nor U2931 (N_2931,In_571,In_936);
or U2932 (N_2932,In_61,In_85);
nor U2933 (N_2933,In_1192,In_1495);
or U2934 (N_2934,In_1716,In_1536);
nor U2935 (N_2935,In_1557,In_1372);
nand U2936 (N_2936,In_1435,In_925);
nand U2937 (N_2937,In_133,In_1169);
nor U2938 (N_2938,In_744,In_764);
nand U2939 (N_2939,In_756,In_146);
nor U2940 (N_2940,In_1637,In_1662);
and U2941 (N_2941,In_1334,In_939);
xor U2942 (N_2942,In_1904,In_1009);
or U2943 (N_2943,In_367,In_728);
nand U2944 (N_2944,In_763,In_437);
nor U2945 (N_2945,In_1778,In_765);
nor U2946 (N_2946,In_1085,In_701);
and U2947 (N_2947,In_1143,In_1767);
or U2948 (N_2948,In_885,In_703);
nor U2949 (N_2949,In_825,In_886);
nand U2950 (N_2950,In_1586,In_491);
and U2951 (N_2951,In_1105,In_207);
or U2952 (N_2952,In_1307,In_1270);
and U2953 (N_2953,In_1201,In_287);
and U2954 (N_2954,In_24,In_946);
or U2955 (N_2955,In_1005,In_690);
or U2956 (N_2956,In_1189,In_258);
nand U2957 (N_2957,In_1977,In_79);
nand U2958 (N_2958,In_1272,In_725);
or U2959 (N_2959,In_380,In_251);
or U2960 (N_2960,In_439,In_1511);
nand U2961 (N_2961,In_837,In_615);
nor U2962 (N_2962,In_1799,In_608);
nand U2963 (N_2963,In_437,In_961);
nand U2964 (N_2964,In_1012,In_1427);
and U2965 (N_2965,In_1862,In_1970);
xnor U2966 (N_2966,In_643,In_1676);
or U2967 (N_2967,In_480,In_1785);
nor U2968 (N_2968,In_1262,In_1626);
nor U2969 (N_2969,In_662,In_26);
or U2970 (N_2970,In_1411,In_1283);
or U2971 (N_2971,In_1821,In_596);
nor U2972 (N_2972,In_787,In_934);
and U2973 (N_2973,In_1893,In_730);
or U2974 (N_2974,In_946,In_877);
or U2975 (N_2975,In_1241,In_1202);
nor U2976 (N_2976,In_69,In_1594);
or U2977 (N_2977,In_1591,In_1779);
or U2978 (N_2978,In_565,In_440);
or U2979 (N_2979,In_199,In_87);
nor U2980 (N_2980,In_844,In_596);
and U2981 (N_2981,In_1208,In_1095);
nor U2982 (N_2982,In_1338,In_146);
nor U2983 (N_2983,In_144,In_916);
nor U2984 (N_2984,In_1926,In_1044);
nor U2985 (N_2985,In_1217,In_1331);
nand U2986 (N_2986,In_1131,In_1878);
nor U2987 (N_2987,In_547,In_1717);
nand U2988 (N_2988,In_1694,In_979);
nand U2989 (N_2989,In_1345,In_1920);
xor U2990 (N_2990,In_223,In_1884);
nand U2991 (N_2991,In_622,In_115);
nand U2992 (N_2992,In_522,In_1113);
nor U2993 (N_2993,In_1399,In_1032);
nand U2994 (N_2994,In_1682,In_1614);
and U2995 (N_2995,In_371,In_803);
nand U2996 (N_2996,In_810,In_975);
or U2997 (N_2997,In_1269,In_111);
nor U2998 (N_2998,In_967,In_1567);
or U2999 (N_2999,In_1692,In_727);
and U3000 (N_3000,In_703,In_1473);
nor U3001 (N_3001,In_552,In_1520);
nand U3002 (N_3002,In_488,In_1800);
nor U3003 (N_3003,In_977,In_813);
or U3004 (N_3004,In_1359,In_1117);
nor U3005 (N_3005,In_1365,In_336);
and U3006 (N_3006,In_619,In_905);
or U3007 (N_3007,In_285,In_1026);
and U3008 (N_3008,In_1458,In_279);
and U3009 (N_3009,In_257,In_1539);
and U3010 (N_3010,In_1477,In_782);
or U3011 (N_3011,In_782,In_1937);
and U3012 (N_3012,In_1670,In_1142);
and U3013 (N_3013,In_885,In_1606);
or U3014 (N_3014,In_1395,In_1908);
or U3015 (N_3015,In_246,In_1247);
and U3016 (N_3016,In_45,In_1724);
or U3017 (N_3017,In_1006,In_498);
nor U3018 (N_3018,In_1732,In_745);
nand U3019 (N_3019,In_953,In_1815);
or U3020 (N_3020,In_1996,In_1803);
nand U3021 (N_3021,In_886,In_1571);
and U3022 (N_3022,In_1852,In_1615);
nand U3023 (N_3023,In_958,In_1421);
and U3024 (N_3024,In_380,In_242);
and U3025 (N_3025,In_913,In_1422);
nand U3026 (N_3026,In_683,In_1096);
and U3027 (N_3027,In_620,In_1954);
nand U3028 (N_3028,In_1586,In_1290);
xor U3029 (N_3029,In_774,In_1291);
nor U3030 (N_3030,In_595,In_1863);
and U3031 (N_3031,In_314,In_1490);
nand U3032 (N_3032,In_1569,In_805);
or U3033 (N_3033,In_1809,In_1931);
or U3034 (N_3034,In_1628,In_1880);
nand U3035 (N_3035,In_806,In_389);
or U3036 (N_3036,In_1519,In_1197);
or U3037 (N_3037,In_477,In_746);
or U3038 (N_3038,In_1252,In_455);
and U3039 (N_3039,In_1067,In_1590);
or U3040 (N_3040,In_238,In_1729);
nand U3041 (N_3041,In_1540,In_529);
nor U3042 (N_3042,In_1058,In_1709);
nor U3043 (N_3043,In_450,In_940);
and U3044 (N_3044,In_1820,In_1575);
nor U3045 (N_3045,In_980,In_0);
nand U3046 (N_3046,In_1931,In_693);
nand U3047 (N_3047,In_1583,In_590);
or U3048 (N_3048,In_1428,In_607);
nand U3049 (N_3049,In_398,In_665);
or U3050 (N_3050,In_1687,In_1997);
nand U3051 (N_3051,In_662,In_269);
or U3052 (N_3052,In_574,In_1276);
and U3053 (N_3053,In_1328,In_129);
nand U3054 (N_3054,In_1158,In_1367);
nand U3055 (N_3055,In_639,In_737);
and U3056 (N_3056,In_766,In_1296);
nor U3057 (N_3057,In_840,In_478);
or U3058 (N_3058,In_1610,In_81);
or U3059 (N_3059,In_782,In_1973);
and U3060 (N_3060,In_48,In_622);
nand U3061 (N_3061,In_772,In_112);
and U3062 (N_3062,In_938,In_876);
or U3063 (N_3063,In_749,In_1616);
or U3064 (N_3064,In_1406,In_1651);
and U3065 (N_3065,In_710,In_809);
and U3066 (N_3066,In_1064,In_1583);
nand U3067 (N_3067,In_594,In_275);
nand U3068 (N_3068,In_1072,In_92);
nand U3069 (N_3069,In_159,In_1028);
and U3070 (N_3070,In_1893,In_1111);
nor U3071 (N_3071,In_803,In_791);
nor U3072 (N_3072,In_619,In_1676);
nor U3073 (N_3073,In_1212,In_682);
or U3074 (N_3074,In_538,In_866);
nor U3075 (N_3075,In_486,In_433);
nand U3076 (N_3076,In_1855,In_1278);
or U3077 (N_3077,In_1267,In_1179);
or U3078 (N_3078,In_445,In_1876);
and U3079 (N_3079,In_502,In_1570);
nand U3080 (N_3080,In_1270,In_1454);
or U3081 (N_3081,In_622,In_1695);
nand U3082 (N_3082,In_630,In_860);
nand U3083 (N_3083,In_1834,In_1474);
or U3084 (N_3084,In_145,In_857);
or U3085 (N_3085,In_453,In_1176);
or U3086 (N_3086,In_1444,In_1487);
nor U3087 (N_3087,In_380,In_1933);
nand U3088 (N_3088,In_1289,In_1713);
nor U3089 (N_3089,In_610,In_3);
nor U3090 (N_3090,In_1409,In_1574);
or U3091 (N_3091,In_1416,In_880);
nand U3092 (N_3092,In_1496,In_1827);
nor U3093 (N_3093,In_1345,In_1437);
nor U3094 (N_3094,In_887,In_1108);
nand U3095 (N_3095,In_217,In_1208);
and U3096 (N_3096,In_1101,In_931);
or U3097 (N_3097,In_1680,In_1295);
nor U3098 (N_3098,In_582,In_1766);
or U3099 (N_3099,In_651,In_1543);
and U3100 (N_3100,In_994,In_217);
nor U3101 (N_3101,In_216,In_348);
or U3102 (N_3102,In_1536,In_1968);
nand U3103 (N_3103,In_291,In_1313);
nor U3104 (N_3104,In_573,In_1128);
or U3105 (N_3105,In_131,In_1140);
nor U3106 (N_3106,In_786,In_1393);
and U3107 (N_3107,In_219,In_220);
nor U3108 (N_3108,In_935,In_1228);
or U3109 (N_3109,In_943,In_1215);
and U3110 (N_3110,In_1191,In_1702);
or U3111 (N_3111,In_275,In_759);
nand U3112 (N_3112,In_247,In_1422);
or U3113 (N_3113,In_1354,In_589);
and U3114 (N_3114,In_1647,In_308);
nand U3115 (N_3115,In_758,In_728);
nor U3116 (N_3116,In_201,In_770);
nor U3117 (N_3117,In_132,In_1243);
and U3118 (N_3118,In_1030,In_1723);
nor U3119 (N_3119,In_964,In_942);
nor U3120 (N_3120,In_1031,In_1230);
and U3121 (N_3121,In_754,In_648);
nand U3122 (N_3122,In_689,In_1391);
nand U3123 (N_3123,In_139,In_484);
or U3124 (N_3124,In_422,In_603);
and U3125 (N_3125,In_634,In_1331);
nor U3126 (N_3126,In_1239,In_132);
nor U3127 (N_3127,In_37,In_1969);
nor U3128 (N_3128,In_408,In_731);
nor U3129 (N_3129,In_801,In_963);
nor U3130 (N_3130,In_1479,In_583);
nor U3131 (N_3131,In_231,In_491);
and U3132 (N_3132,In_953,In_1901);
xor U3133 (N_3133,In_433,In_328);
and U3134 (N_3134,In_185,In_641);
and U3135 (N_3135,In_966,In_1493);
nor U3136 (N_3136,In_1553,In_892);
xor U3137 (N_3137,In_1102,In_1584);
nor U3138 (N_3138,In_18,In_1893);
or U3139 (N_3139,In_1938,In_1289);
or U3140 (N_3140,In_321,In_888);
or U3141 (N_3141,In_1970,In_1398);
and U3142 (N_3142,In_1504,In_1428);
nor U3143 (N_3143,In_1293,In_122);
nor U3144 (N_3144,In_506,In_1017);
nand U3145 (N_3145,In_1509,In_1455);
nand U3146 (N_3146,In_570,In_183);
and U3147 (N_3147,In_529,In_48);
xnor U3148 (N_3148,In_1690,In_921);
nand U3149 (N_3149,In_1726,In_565);
nand U3150 (N_3150,In_819,In_1948);
nand U3151 (N_3151,In_749,In_1058);
or U3152 (N_3152,In_1465,In_979);
nand U3153 (N_3153,In_34,In_230);
nor U3154 (N_3154,In_583,In_1287);
nor U3155 (N_3155,In_982,In_1875);
or U3156 (N_3156,In_1260,In_790);
nor U3157 (N_3157,In_1016,In_559);
nand U3158 (N_3158,In_403,In_1343);
nand U3159 (N_3159,In_1881,In_1520);
and U3160 (N_3160,In_1296,In_1314);
or U3161 (N_3161,In_1718,In_1522);
nand U3162 (N_3162,In_1651,In_1112);
and U3163 (N_3163,In_445,In_1790);
and U3164 (N_3164,In_309,In_432);
or U3165 (N_3165,In_935,In_1128);
and U3166 (N_3166,In_1042,In_1141);
nand U3167 (N_3167,In_1602,In_352);
and U3168 (N_3168,In_1751,In_1358);
or U3169 (N_3169,In_1483,In_1482);
nor U3170 (N_3170,In_754,In_120);
and U3171 (N_3171,In_516,In_1955);
xor U3172 (N_3172,In_392,In_1523);
nand U3173 (N_3173,In_1498,In_1552);
and U3174 (N_3174,In_314,In_1344);
nor U3175 (N_3175,In_216,In_1513);
nor U3176 (N_3176,In_689,In_1519);
or U3177 (N_3177,In_1499,In_1784);
or U3178 (N_3178,In_872,In_1784);
or U3179 (N_3179,In_351,In_1877);
or U3180 (N_3180,In_1506,In_920);
and U3181 (N_3181,In_1789,In_126);
and U3182 (N_3182,In_1470,In_927);
nand U3183 (N_3183,In_1542,In_571);
nand U3184 (N_3184,In_1847,In_107);
and U3185 (N_3185,In_1185,In_692);
or U3186 (N_3186,In_24,In_977);
nand U3187 (N_3187,In_1122,In_1730);
nand U3188 (N_3188,In_405,In_350);
or U3189 (N_3189,In_506,In_1534);
nor U3190 (N_3190,In_847,In_740);
and U3191 (N_3191,In_448,In_1659);
nand U3192 (N_3192,In_767,In_774);
and U3193 (N_3193,In_827,In_817);
and U3194 (N_3194,In_313,In_293);
nor U3195 (N_3195,In_621,In_1671);
and U3196 (N_3196,In_303,In_382);
nor U3197 (N_3197,In_209,In_883);
nand U3198 (N_3198,In_923,In_1730);
nand U3199 (N_3199,In_470,In_1627);
nand U3200 (N_3200,In_1006,In_226);
nor U3201 (N_3201,In_526,In_713);
nand U3202 (N_3202,In_1431,In_1406);
and U3203 (N_3203,In_297,In_493);
and U3204 (N_3204,In_1394,In_702);
nor U3205 (N_3205,In_1402,In_1240);
and U3206 (N_3206,In_571,In_1761);
nor U3207 (N_3207,In_1120,In_1591);
nand U3208 (N_3208,In_1764,In_1685);
or U3209 (N_3209,In_1433,In_1114);
and U3210 (N_3210,In_989,In_1325);
nor U3211 (N_3211,In_1430,In_1221);
or U3212 (N_3212,In_413,In_1777);
nand U3213 (N_3213,In_621,In_492);
nand U3214 (N_3214,In_1395,In_1085);
and U3215 (N_3215,In_927,In_1801);
or U3216 (N_3216,In_1060,In_1352);
nor U3217 (N_3217,In_1461,In_397);
or U3218 (N_3218,In_1416,In_1111);
or U3219 (N_3219,In_1057,In_1909);
and U3220 (N_3220,In_1809,In_1190);
and U3221 (N_3221,In_1768,In_1108);
or U3222 (N_3222,In_639,In_1677);
nand U3223 (N_3223,In_1107,In_1282);
nand U3224 (N_3224,In_1796,In_619);
nand U3225 (N_3225,In_50,In_141);
and U3226 (N_3226,In_1625,In_605);
nor U3227 (N_3227,In_1874,In_317);
and U3228 (N_3228,In_803,In_1116);
and U3229 (N_3229,In_419,In_716);
and U3230 (N_3230,In_801,In_513);
or U3231 (N_3231,In_1454,In_1831);
nor U3232 (N_3232,In_1243,In_186);
nor U3233 (N_3233,In_1922,In_1866);
or U3234 (N_3234,In_1026,In_496);
nor U3235 (N_3235,In_650,In_189);
and U3236 (N_3236,In_1593,In_362);
nor U3237 (N_3237,In_1038,In_1099);
nand U3238 (N_3238,In_1963,In_137);
nand U3239 (N_3239,In_1269,In_899);
nand U3240 (N_3240,In_34,In_1464);
nand U3241 (N_3241,In_913,In_1473);
and U3242 (N_3242,In_395,In_1192);
or U3243 (N_3243,In_1597,In_867);
nand U3244 (N_3244,In_474,In_522);
nand U3245 (N_3245,In_1152,In_779);
nor U3246 (N_3246,In_681,In_580);
nor U3247 (N_3247,In_491,In_431);
nand U3248 (N_3248,In_1747,In_1849);
nor U3249 (N_3249,In_1355,In_1081);
nor U3250 (N_3250,In_792,In_1877);
or U3251 (N_3251,In_1358,In_1210);
xor U3252 (N_3252,In_1705,In_916);
nor U3253 (N_3253,In_1472,In_451);
nand U3254 (N_3254,In_516,In_1374);
or U3255 (N_3255,In_1923,In_1625);
or U3256 (N_3256,In_1965,In_1590);
or U3257 (N_3257,In_162,In_1718);
and U3258 (N_3258,In_1572,In_125);
nor U3259 (N_3259,In_367,In_842);
or U3260 (N_3260,In_129,In_695);
nand U3261 (N_3261,In_1799,In_1416);
nand U3262 (N_3262,In_848,In_1579);
nor U3263 (N_3263,In_1286,In_1263);
and U3264 (N_3264,In_1789,In_1197);
or U3265 (N_3265,In_1952,In_1586);
xor U3266 (N_3266,In_832,In_983);
nand U3267 (N_3267,In_826,In_1935);
nand U3268 (N_3268,In_603,In_292);
nor U3269 (N_3269,In_262,In_1079);
nand U3270 (N_3270,In_664,In_652);
or U3271 (N_3271,In_67,In_366);
nand U3272 (N_3272,In_1237,In_1677);
and U3273 (N_3273,In_814,In_1594);
nand U3274 (N_3274,In_1326,In_1620);
or U3275 (N_3275,In_1523,In_1517);
nand U3276 (N_3276,In_984,In_1228);
nor U3277 (N_3277,In_1305,In_1293);
nor U3278 (N_3278,In_36,In_400);
xor U3279 (N_3279,In_1575,In_1063);
and U3280 (N_3280,In_733,In_1005);
and U3281 (N_3281,In_244,In_250);
and U3282 (N_3282,In_1028,In_883);
nor U3283 (N_3283,In_1181,In_1945);
or U3284 (N_3284,In_1111,In_338);
nor U3285 (N_3285,In_1852,In_961);
xor U3286 (N_3286,In_15,In_351);
nand U3287 (N_3287,In_1299,In_1297);
or U3288 (N_3288,In_1790,In_1599);
or U3289 (N_3289,In_1100,In_1934);
xor U3290 (N_3290,In_891,In_992);
and U3291 (N_3291,In_799,In_1565);
nand U3292 (N_3292,In_1127,In_1105);
and U3293 (N_3293,In_857,In_662);
nor U3294 (N_3294,In_496,In_359);
and U3295 (N_3295,In_324,In_50);
and U3296 (N_3296,In_627,In_1362);
nand U3297 (N_3297,In_1035,In_410);
nor U3298 (N_3298,In_694,In_841);
nand U3299 (N_3299,In_1059,In_1271);
or U3300 (N_3300,In_65,In_595);
or U3301 (N_3301,In_795,In_1698);
nor U3302 (N_3302,In_1707,In_518);
or U3303 (N_3303,In_775,In_1580);
or U3304 (N_3304,In_488,In_922);
nand U3305 (N_3305,In_397,In_1747);
nor U3306 (N_3306,In_1989,In_1616);
nor U3307 (N_3307,In_27,In_1653);
and U3308 (N_3308,In_1465,In_1437);
nand U3309 (N_3309,In_1196,In_954);
nand U3310 (N_3310,In_1152,In_1663);
and U3311 (N_3311,In_297,In_665);
and U3312 (N_3312,In_1339,In_929);
nor U3313 (N_3313,In_936,In_1216);
and U3314 (N_3314,In_744,In_225);
and U3315 (N_3315,In_1625,In_397);
nor U3316 (N_3316,In_813,In_891);
nand U3317 (N_3317,In_1176,In_1333);
and U3318 (N_3318,In_135,In_934);
and U3319 (N_3319,In_1259,In_500);
nor U3320 (N_3320,In_1296,In_1276);
and U3321 (N_3321,In_863,In_1206);
nand U3322 (N_3322,In_663,In_811);
and U3323 (N_3323,In_311,In_75);
or U3324 (N_3324,In_1444,In_668);
and U3325 (N_3325,In_422,In_667);
nor U3326 (N_3326,In_1900,In_1036);
nand U3327 (N_3327,In_1944,In_283);
nand U3328 (N_3328,In_1825,In_1068);
and U3329 (N_3329,In_531,In_1999);
nor U3330 (N_3330,In_1686,In_769);
and U3331 (N_3331,In_625,In_169);
and U3332 (N_3332,In_436,In_843);
xor U3333 (N_3333,In_819,In_263);
nand U3334 (N_3334,In_1276,In_1203);
and U3335 (N_3335,In_717,In_591);
and U3336 (N_3336,In_924,In_1472);
and U3337 (N_3337,In_1535,In_1601);
nand U3338 (N_3338,In_693,In_230);
and U3339 (N_3339,In_635,In_1171);
and U3340 (N_3340,In_212,In_1547);
or U3341 (N_3341,In_896,In_809);
nand U3342 (N_3342,In_1049,In_1014);
and U3343 (N_3343,In_1648,In_976);
or U3344 (N_3344,In_1059,In_1565);
nand U3345 (N_3345,In_611,In_1218);
nand U3346 (N_3346,In_1812,In_1827);
or U3347 (N_3347,In_774,In_1603);
and U3348 (N_3348,In_328,In_20);
or U3349 (N_3349,In_1853,In_1784);
or U3350 (N_3350,In_902,In_1545);
nand U3351 (N_3351,In_1570,In_210);
nand U3352 (N_3352,In_1028,In_1482);
nand U3353 (N_3353,In_61,In_908);
or U3354 (N_3354,In_1965,In_1451);
nor U3355 (N_3355,In_1124,In_506);
or U3356 (N_3356,In_1835,In_895);
or U3357 (N_3357,In_554,In_1261);
nand U3358 (N_3358,In_896,In_651);
and U3359 (N_3359,In_1992,In_832);
and U3360 (N_3360,In_201,In_1992);
and U3361 (N_3361,In_1197,In_1403);
nand U3362 (N_3362,In_1531,In_1888);
or U3363 (N_3363,In_897,In_1178);
nand U3364 (N_3364,In_712,In_1699);
and U3365 (N_3365,In_1623,In_1529);
nand U3366 (N_3366,In_834,In_1938);
nand U3367 (N_3367,In_1967,In_334);
and U3368 (N_3368,In_802,In_1911);
or U3369 (N_3369,In_650,In_1447);
or U3370 (N_3370,In_364,In_1317);
or U3371 (N_3371,In_1293,In_1256);
nand U3372 (N_3372,In_1060,In_799);
nor U3373 (N_3373,In_99,In_1525);
or U3374 (N_3374,In_911,In_1947);
and U3375 (N_3375,In_1450,In_1625);
or U3376 (N_3376,In_1892,In_1006);
or U3377 (N_3377,In_1306,In_259);
and U3378 (N_3378,In_928,In_832);
nand U3379 (N_3379,In_489,In_102);
or U3380 (N_3380,In_1328,In_939);
nand U3381 (N_3381,In_228,In_1338);
nand U3382 (N_3382,In_866,In_1125);
and U3383 (N_3383,In_361,In_45);
nor U3384 (N_3384,In_750,In_1832);
or U3385 (N_3385,In_937,In_268);
nand U3386 (N_3386,In_240,In_1174);
nor U3387 (N_3387,In_350,In_1563);
nand U3388 (N_3388,In_849,In_1727);
or U3389 (N_3389,In_347,In_1286);
or U3390 (N_3390,In_1361,In_1922);
nand U3391 (N_3391,In_860,In_1321);
nor U3392 (N_3392,In_972,In_879);
or U3393 (N_3393,In_1392,In_1442);
nand U3394 (N_3394,In_171,In_519);
nor U3395 (N_3395,In_259,In_504);
nor U3396 (N_3396,In_369,In_991);
nor U3397 (N_3397,In_206,In_1959);
nand U3398 (N_3398,In_1933,In_1015);
and U3399 (N_3399,In_1497,In_1058);
nand U3400 (N_3400,In_392,In_159);
or U3401 (N_3401,In_486,In_800);
nor U3402 (N_3402,In_1025,In_1885);
and U3403 (N_3403,In_1374,In_105);
or U3404 (N_3404,In_1614,In_1510);
and U3405 (N_3405,In_706,In_1231);
or U3406 (N_3406,In_64,In_1520);
nor U3407 (N_3407,In_183,In_1549);
and U3408 (N_3408,In_1965,In_1037);
xnor U3409 (N_3409,In_1013,In_1544);
or U3410 (N_3410,In_1839,In_1420);
or U3411 (N_3411,In_867,In_1021);
nand U3412 (N_3412,In_1975,In_217);
nor U3413 (N_3413,In_864,In_64);
nor U3414 (N_3414,In_1639,In_908);
nor U3415 (N_3415,In_270,In_1870);
and U3416 (N_3416,In_872,In_514);
or U3417 (N_3417,In_568,In_716);
or U3418 (N_3418,In_125,In_279);
nand U3419 (N_3419,In_1889,In_58);
and U3420 (N_3420,In_124,In_794);
and U3421 (N_3421,In_1368,In_1734);
nand U3422 (N_3422,In_1405,In_607);
nor U3423 (N_3423,In_1832,In_133);
or U3424 (N_3424,In_1752,In_1224);
nand U3425 (N_3425,In_217,In_865);
nand U3426 (N_3426,In_1097,In_163);
or U3427 (N_3427,In_1404,In_836);
nor U3428 (N_3428,In_508,In_1405);
or U3429 (N_3429,In_281,In_1480);
nor U3430 (N_3430,In_281,In_1629);
nor U3431 (N_3431,In_1962,In_495);
and U3432 (N_3432,In_464,In_58);
or U3433 (N_3433,In_1567,In_1073);
nor U3434 (N_3434,In_1957,In_639);
nand U3435 (N_3435,In_1974,In_824);
or U3436 (N_3436,In_747,In_372);
nor U3437 (N_3437,In_1711,In_219);
and U3438 (N_3438,In_1212,In_890);
and U3439 (N_3439,In_1795,In_141);
or U3440 (N_3440,In_215,In_1103);
or U3441 (N_3441,In_268,In_676);
nor U3442 (N_3442,In_1242,In_674);
xnor U3443 (N_3443,In_1366,In_328);
nand U3444 (N_3444,In_781,In_1161);
nor U3445 (N_3445,In_1265,In_1094);
nand U3446 (N_3446,In_1645,In_1858);
nor U3447 (N_3447,In_88,In_1068);
nor U3448 (N_3448,In_880,In_1666);
or U3449 (N_3449,In_652,In_359);
nand U3450 (N_3450,In_0,In_1174);
and U3451 (N_3451,In_1462,In_481);
nand U3452 (N_3452,In_1538,In_1340);
and U3453 (N_3453,In_378,In_1985);
or U3454 (N_3454,In_1963,In_539);
and U3455 (N_3455,In_1726,In_1032);
nor U3456 (N_3456,In_1855,In_1254);
nor U3457 (N_3457,In_243,In_1564);
nor U3458 (N_3458,In_1089,In_454);
nand U3459 (N_3459,In_342,In_790);
nor U3460 (N_3460,In_1070,In_1837);
nor U3461 (N_3461,In_752,In_1562);
or U3462 (N_3462,In_468,In_1886);
or U3463 (N_3463,In_1105,In_1238);
and U3464 (N_3464,In_691,In_68);
nor U3465 (N_3465,In_603,In_1430);
nand U3466 (N_3466,In_1071,In_1872);
and U3467 (N_3467,In_210,In_1486);
nor U3468 (N_3468,In_854,In_1198);
nor U3469 (N_3469,In_96,In_1505);
and U3470 (N_3470,In_986,In_570);
nand U3471 (N_3471,In_444,In_1969);
and U3472 (N_3472,In_988,In_1321);
nand U3473 (N_3473,In_1350,In_935);
nand U3474 (N_3474,In_730,In_1305);
nand U3475 (N_3475,In_805,In_91);
and U3476 (N_3476,In_295,In_366);
nor U3477 (N_3477,In_1266,In_201);
or U3478 (N_3478,In_1976,In_431);
nand U3479 (N_3479,In_1773,In_1799);
or U3480 (N_3480,In_793,In_1289);
and U3481 (N_3481,In_941,In_944);
nor U3482 (N_3482,In_569,In_773);
nand U3483 (N_3483,In_444,In_1394);
or U3484 (N_3484,In_473,In_1696);
or U3485 (N_3485,In_1334,In_479);
or U3486 (N_3486,In_1616,In_625);
nor U3487 (N_3487,In_1028,In_1861);
nand U3488 (N_3488,In_1868,In_1525);
or U3489 (N_3489,In_1223,In_220);
nor U3490 (N_3490,In_1575,In_694);
nor U3491 (N_3491,In_321,In_706);
and U3492 (N_3492,In_739,In_548);
nand U3493 (N_3493,In_1768,In_454);
nand U3494 (N_3494,In_165,In_1849);
nor U3495 (N_3495,In_419,In_1888);
nor U3496 (N_3496,In_1281,In_365);
nor U3497 (N_3497,In_1652,In_1802);
nand U3498 (N_3498,In_1855,In_597);
and U3499 (N_3499,In_1486,In_1753);
nand U3500 (N_3500,In_1521,In_794);
and U3501 (N_3501,In_115,In_679);
or U3502 (N_3502,In_667,In_1850);
or U3503 (N_3503,In_948,In_606);
or U3504 (N_3504,In_140,In_1042);
or U3505 (N_3505,In_31,In_1227);
nand U3506 (N_3506,In_1075,In_215);
and U3507 (N_3507,In_1133,In_1001);
and U3508 (N_3508,In_1646,In_1089);
nand U3509 (N_3509,In_315,In_1080);
nor U3510 (N_3510,In_1357,In_1748);
or U3511 (N_3511,In_1667,In_308);
or U3512 (N_3512,In_733,In_1822);
and U3513 (N_3513,In_180,In_1842);
nand U3514 (N_3514,In_619,In_1014);
or U3515 (N_3515,In_1866,In_1513);
and U3516 (N_3516,In_1599,In_1827);
and U3517 (N_3517,In_802,In_1200);
and U3518 (N_3518,In_846,In_1964);
nand U3519 (N_3519,In_172,In_1168);
or U3520 (N_3520,In_997,In_1996);
or U3521 (N_3521,In_373,In_965);
nor U3522 (N_3522,In_1262,In_40);
and U3523 (N_3523,In_1784,In_862);
nor U3524 (N_3524,In_866,In_1810);
nor U3525 (N_3525,In_1349,In_442);
or U3526 (N_3526,In_982,In_673);
nor U3527 (N_3527,In_991,In_754);
nor U3528 (N_3528,In_216,In_1074);
or U3529 (N_3529,In_792,In_804);
nand U3530 (N_3530,In_672,In_1645);
and U3531 (N_3531,In_987,In_1384);
nand U3532 (N_3532,In_962,In_937);
nor U3533 (N_3533,In_752,In_1917);
and U3534 (N_3534,In_1559,In_972);
nand U3535 (N_3535,In_614,In_817);
and U3536 (N_3536,In_1935,In_1378);
or U3537 (N_3537,In_801,In_362);
and U3538 (N_3538,In_525,In_748);
or U3539 (N_3539,In_326,In_891);
nand U3540 (N_3540,In_1806,In_792);
and U3541 (N_3541,In_1123,In_1881);
nor U3542 (N_3542,In_1021,In_982);
or U3543 (N_3543,In_359,In_1414);
nand U3544 (N_3544,In_227,In_527);
and U3545 (N_3545,In_905,In_412);
or U3546 (N_3546,In_404,In_445);
nor U3547 (N_3547,In_1868,In_494);
and U3548 (N_3548,In_243,In_12);
nor U3549 (N_3549,In_1900,In_874);
and U3550 (N_3550,In_252,In_177);
and U3551 (N_3551,In_1069,In_1117);
xor U3552 (N_3552,In_947,In_884);
nor U3553 (N_3553,In_1069,In_566);
nor U3554 (N_3554,In_1521,In_407);
nand U3555 (N_3555,In_972,In_942);
and U3556 (N_3556,In_1028,In_193);
nand U3557 (N_3557,In_270,In_168);
nand U3558 (N_3558,In_1331,In_1361);
and U3559 (N_3559,In_1901,In_1133);
nor U3560 (N_3560,In_716,In_764);
or U3561 (N_3561,In_503,In_842);
and U3562 (N_3562,In_1302,In_1399);
nand U3563 (N_3563,In_207,In_753);
and U3564 (N_3564,In_795,In_1673);
and U3565 (N_3565,In_1687,In_704);
nor U3566 (N_3566,In_1522,In_1686);
or U3567 (N_3567,In_387,In_627);
or U3568 (N_3568,In_337,In_1968);
nand U3569 (N_3569,In_130,In_1741);
nor U3570 (N_3570,In_165,In_1783);
and U3571 (N_3571,In_767,In_799);
nand U3572 (N_3572,In_749,In_983);
and U3573 (N_3573,In_633,In_925);
nor U3574 (N_3574,In_1412,In_1143);
or U3575 (N_3575,In_1212,In_580);
xor U3576 (N_3576,In_613,In_128);
and U3577 (N_3577,In_1984,In_1464);
and U3578 (N_3578,In_291,In_955);
and U3579 (N_3579,In_278,In_224);
nor U3580 (N_3580,In_521,In_150);
nor U3581 (N_3581,In_1292,In_1274);
nor U3582 (N_3582,In_81,In_1818);
nor U3583 (N_3583,In_1317,In_660);
nand U3584 (N_3584,In_745,In_595);
and U3585 (N_3585,In_58,In_1303);
and U3586 (N_3586,In_307,In_1802);
nor U3587 (N_3587,In_1462,In_1576);
nand U3588 (N_3588,In_144,In_607);
or U3589 (N_3589,In_267,In_1783);
nor U3590 (N_3590,In_1491,In_1024);
nor U3591 (N_3591,In_251,In_1841);
or U3592 (N_3592,In_1638,In_447);
and U3593 (N_3593,In_1214,In_1679);
nor U3594 (N_3594,In_1298,In_411);
nand U3595 (N_3595,In_169,In_250);
nor U3596 (N_3596,In_359,In_1392);
and U3597 (N_3597,In_1048,In_1762);
and U3598 (N_3598,In_1750,In_1768);
nor U3599 (N_3599,In_1353,In_1875);
nand U3600 (N_3600,In_73,In_405);
nand U3601 (N_3601,In_1579,In_1831);
nand U3602 (N_3602,In_570,In_492);
nor U3603 (N_3603,In_1983,In_1935);
nor U3604 (N_3604,In_1529,In_953);
or U3605 (N_3605,In_1188,In_580);
nand U3606 (N_3606,In_636,In_1786);
nor U3607 (N_3607,In_168,In_1995);
xnor U3608 (N_3608,In_500,In_1467);
nand U3609 (N_3609,In_1836,In_366);
nor U3610 (N_3610,In_1912,In_1964);
and U3611 (N_3611,In_827,In_1704);
nand U3612 (N_3612,In_1136,In_1630);
or U3613 (N_3613,In_358,In_192);
and U3614 (N_3614,In_910,In_289);
nor U3615 (N_3615,In_1296,In_1165);
nor U3616 (N_3616,In_276,In_873);
nor U3617 (N_3617,In_827,In_856);
nor U3618 (N_3618,In_1316,In_1802);
or U3619 (N_3619,In_398,In_1160);
or U3620 (N_3620,In_1581,In_1230);
or U3621 (N_3621,In_1741,In_1546);
nor U3622 (N_3622,In_1018,In_1733);
xnor U3623 (N_3623,In_1802,In_1012);
nand U3624 (N_3624,In_1,In_965);
or U3625 (N_3625,In_530,In_1166);
xor U3626 (N_3626,In_1285,In_999);
or U3627 (N_3627,In_1554,In_1221);
nor U3628 (N_3628,In_1843,In_1110);
or U3629 (N_3629,In_818,In_1775);
nand U3630 (N_3630,In_1985,In_1342);
nand U3631 (N_3631,In_315,In_1757);
nor U3632 (N_3632,In_283,In_802);
and U3633 (N_3633,In_417,In_601);
nor U3634 (N_3634,In_494,In_1680);
or U3635 (N_3635,In_654,In_1023);
or U3636 (N_3636,In_1852,In_1935);
nor U3637 (N_3637,In_1983,In_293);
or U3638 (N_3638,In_1623,In_1954);
or U3639 (N_3639,In_856,In_260);
nand U3640 (N_3640,In_944,In_1227);
nor U3641 (N_3641,In_1931,In_1894);
nor U3642 (N_3642,In_383,In_1126);
nand U3643 (N_3643,In_594,In_1419);
and U3644 (N_3644,In_970,In_664);
or U3645 (N_3645,In_1090,In_1266);
nand U3646 (N_3646,In_180,In_1345);
and U3647 (N_3647,In_1278,In_390);
nand U3648 (N_3648,In_1603,In_899);
xnor U3649 (N_3649,In_112,In_358);
nand U3650 (N_3650,In_3,In_54);
nor U3651 (N_3651,In_461,In_1652);
nor U3652 (N_3652,In_1159,In_1994);
nor U3653 (N_3653,In_1891,In_1183);
and U3654 (N_3654,In_357,In_907);
nand U3655 (N_3655,In_1513,In_1862);
or U3656 (N_3656,In_827,In_511);
or U3657 (N_3657,In_1214,In_40);
and U3658 (N_3658,In_1473,In_1943);
and U3659 (N_3659,In_447,In_384);
nor U3660 (N_3660,In_859,In_1308);
nor U3661 (N_3661,In_1102,In_1754);
nand U3662 (N_3662,In_1261,In_865);
or U3663 (N_3663,In_1857,In_1216);
nand U3664 (N_3664,In_253,In_1835);
and U3665 (N_3665,In_845,In_1750);
or U3666 (N_3666,In_789,In_1051);
nand U3667 (N_3667,In_287,In_1580);
nand U3668 (N_3668,In_1093,In_293);
nor U3669 (N_3669,In_1864,In_1463);
and U3670 (N_3670,In_1345,In_240);
nor U3671 (N_3671,In_1382,In_362);
nor U3672 (N_3672,In_1693,In_1143);
nand U3673 (N_3673,In_1987,In_815);
nand U3674 (N_3674,In_337,In_1591);
and U3675 (N_3675,In_1099,In_539);
and U3676 (N_3676,In_236,In_627);
or U3677 (N_3677,In_692,In_1086);
nor U3678 (N_3678,In_1175,In_1598);
nand U3679 (N_3679,In_1375,In_1350);
nand U3680 (N_3680,In_1622,In_1191);
nor U3681 (N_3681,In_803,In_1299);
nor U3682 (N_3682,In_1193,In_946);
nand U3683 (N_3683,In_143,In_841);
nor U3684 (N_3684,In_1074,In_1787);
or U3685 (N_3685,In_1029,In_620);
or U3686 (N_3686,In_554,In_1193);
and U3687 (N_3687,In_1887,In_73);
nand U3688 (N_3688,In_1652,In_1675);
or U3689 (N_3689,In_386,In_1583);
or U3690 (N_3690,In_4,In_1509);
nand U3691 (N_3691,In_629,In_1147);
nor U3692 (N_3692,In_1793,In_1775);
and U3693 (N_3693,In_755,In_1171);
or U3694 (N_3694,In_836,In_910);
and U3695 (N_3695,In_52,In_393);
or U3696 (N_3696,In_1543,In_404);
or U3697 (N_3697,In_1265,In_607);
or U3698 (N_3698,In_1002,In_879);
nand U3699 (N_3699,In_1799,In_1889);
nand U3700 (N_3700,In_1319,In_817);
and U3701 (N_3701,In_1117,In_771);
and U3702 (N_3702,In_238,In_1665);
xnor U3703 (N_3703,In_895,In_688);
and U3704 (N_3704,In_1788,In_55);
and U3705 (N_3705,In_1915,In_1365);
and U3706 (N_3706,In_523,In_1528);
xor U3707 (N_3707,In_123,In_907);
nor U3708 (N_3708,In_1338,In_1748);
nor U3709 (N_3709,In_1715,In_551);
and U3710 (N_3710,In_1748,In_432);
nand U3711 (N_3711,In_86,In_522);
or U3712 (N_3712,In_64,In_355);
or U3713 (N_3713,In_996,In_1625);
nor U3714 (N_3714,In_625,In_1230);
nand U3715 (N_3715,In_536,In_335);
or U3716 (N_3716,In_1234,In_1562);
nand U3717 (N_3717,In_579,In_1295);
and U3718 (N_3718,In_238,In_825);
and U3719 (N_3719,In_428,In_1369);
nand U3720 (N_3720,In_232,In_1086);
nor U3721 (N_3721,In_1498,In_499);
nand U3722 (N_3722,In_446,In_69);
or U3723 (N_3723,In_827,In_1629);
and U3724 (N_3724,In_1604,In_701);
nand U3725 (N_3725,In_1665,In_610);
nand U3726 (N_3726,In_79,In_418);
xor U3727 (N_3727,In_222,In_691);
or U3728 (N_3728,In_689,In_1205);
nor U3729 (N_3729,In_804,In_908);
nand U3730 (N_3730,In_1537,In_794);
nand U3731 (N_3731,In_615,In_444);
or U3732 (N_3732,In_35,In_1774);
nand U3733 (N_3733,In_17,In_1085);
nor U3734 (N_3734,In_46,In_888);
nor U3735 (N_3735,In_856,In_34);
nor U3736 (N_3736,In_1796,In_1100);
nand U3737 (N_3737,In_965,In_951);
and U3738 (N_3738,In_677,In_1889);
nand U3739 (N_3739,In_966,In_523);
nand U3740 (N_3740,In_531,In_630);
nor U3741 (N_3741,In_1714,In_979);
and U3742 (N_3742,In_129,In_932);
or U3743 (N_3743,In_67,In_1436);
nand U3744 (N_3744,In_683,In_1637);
nor U3745 (N_3745,In_783,In_255);
and U3746 (N_3746,In_860,In_1183);
nor U3747 (N_3747,In_760,In_1989);
and U3748 (N_3748,In_212,In_377);
nand U3749 (N_3749,In_1046,In_1391);
nor U3750 (N_3750,In_1542,In_1230);
and U3751 (N_3751,In_697,In_1503);
nor U3752 (N_3752,In_1081,In_1912);
nand U3753 (N_3753,In_1379,In_1155);
nor U3754 (N_3754,In_394,In_475);
nor U3755 (N_3755,In_1287,In_1292);
and U3756 (N_3756,In_201,In_1926);
nor U3757 (N_3757,In_1360,In_1804);
or U3758 (N_3758,In_1935,In_1785);
or U3759 (N_3759,In_1569,In_1006);
nor U3760 (N_3760,In_604,In_1430);
or U3761 (N_3761,In_1483,In_1027);
nor U3762 (N_3762,In_943,In_873);
nor U3763 (N_3763,In_1670,In_1000);
nand U3764 (N_3764,In_153,In_1423);
nand U3765 (N_3765,In_960,In_1996);
or U3766 (N_3766,In_1077,In_1060);
nand U3767 (N_3767,In_1046,In_107);
nand U3768 (N_3768,In_462,In_1773);
nand U3769 (N_3769,In_970,In_1840);
nand U3770 (N_3770,In_1496,In_581);
nor U3771 (N_3771,In_1234,In_1283);
or U3772 (N_3772,In_1826,In_1001);
or U3773 (N_3773,In_1399,In_1273);
nor U3774 (N_3774,In_904,In_1233);
nand U3775 (N_3775,In_1548,In_1556);
or U3776 (N_3776,In_1402,In_591);
xor U3777 (N_3777,In_946,In_1319);
nand U3778 (N_3778,In_679,In_183);
and U3779 (N_3779,In_107,In_861);
nor U3780 (N_3780,In_669,In_522);
and U3781 (N_3781,In_489,In_1492);
or U3782 (N_3782,In_534,In_1905);
and U3783 (N_3783,In_1581,In_361);
and U3784 (N_3784,In_831,In_1200);
and U3785 (N_3785,In_1904,In_88);
or U3786 (N_3786,In_1334,In_1300);
nand U3787 (N_3787,In_1098,In_1891);
nand U3788 (N_3788,In_1781,In_141);
nor U3789 (N_3789,In_1319,In_1815);
nand U3790 (N_3790,In_880,In_87);
and U3791 (N_3791,In_59,In_452);
nor U3792 (N_3792,In_1256,In_1263);
and U3793 (N_3793,In_1869,In_403);
nand U3794 (N_3794,In_159,In_1503);
nand U3795 (N_3795,In_479,In_33);
or U3796 (N_3796,In_500,In_1189);
or U3797 (N_3797,In_116,In_1287);
and U3798 (N_3798,In_1142,In_726);
or U3799 (N_3799,In_1019,In_1449);
nor U3800 (N_3800,In_781,In_65);
or U3801 (N_3801,In_263,In_1364);
nor U3802 (N_3802,In_697,In_1325);
and U3803 (N_3803,In_65,In_1755);
nand U3804 (N_3804,In_1104,In_1398);
or U3805 (N_3805,In_1606,In_1925);
or U3806 (N_3806,In_1999,In_1063);
nor U3807 (N_3807,In_1575,In_271);
nand U3808 (N_3808,In_575,In_377);
nand U3809 (N_3809,In_240,In_1126);
nor U3810 (N_3810,In_1813,In_1654);
or U3811 (N_3811,In_1734,In_979);
nand U3812 (N_3812,In_405,In_772);
or U3813 (N_3813,In_1612,In_440);
and U3814 (N_3814,In_104,In_1437);
or U3815 (N_3815,In_335,In_1648);
or U3816 (N_3816,In_419,In_1668);
nor U3817 (N_3817,In_435,In_1661);
or U3818 (N_3818,In_1535,In_920);
or U3819 (N_3819,In_1412,In_1063);
nor U3820 (N_3820,In_756,In_244);
xnor U3821 (N_3821,In_1966,In_870);
or U3822 (N_3822,In_1385,In_154);
xnor U3823 (N_3823,In_1193,In_700);
nor U3824 (N_3824,In_491,In_1026);
nand U3825 (N_3825,In_1860,In_295);
or U3826 (N_3826,In_1769,In_1053);
or U3827 (N_3827,In_502,In_549);
and U3828 (N_3828,In_341,In_1619);
or U3829 (N_3829,In_825,In_20);
and U3830 (N_3830,In_1119,In_119);
nor U3831 (N_3831,In_1712,In_878);
and U3832 (N_3832,In_720,In_1501);
or U3833 (N_3833,In_1932,In_1803);
nor U3834 (N_3834,In_1538,In_1727);
nor U3835 (N_3835,In_594,In_1444);
nand U3836 (N_3836,In_617,In_1120);
or U3837 (N_3837,In_753,In_184);
xnor U3838 (N_3838,In_962,In_812);
nor U3839 (N_3839,In_1149,In_984);
nand U3840 (N_3840,In_1757,In_1555);
nand U3841 (N_3841,In_1145,In_968);
and U3842 (N_3842,In_801,In_326);
and U3843 (N_3843,In_1960,In_1187);
nand U3844 (N_3844,In_1389,In_235);
nand U3845 (N_3845,In_532,In_1721);
or U3846 (N_3846,In_327,In_1864);
or U3847 (N_3847,In_1296,In_503);
and U3848 (N_3848,In_541,In_260);
or U3849 (N_3849,In_843,In_1526);
or U3850 (N_3850,In_1058,In_912);
and U3851 (N_3851,In_1572,In_1447);
nand U3852 (N_3852,In_1539,In_1787);
or U3853 (N_3853,In_179,In_505);
and U3854 (N_3854,In_1932,In_310);
nand U3855 (N_3855,In_1426,In_640);
or U3856 (N_3856,In_740,In_137);
and U3857 (N_3857,In_345,In_1330);
and U3858 (N_3858,In_1071,In_522);
nand U3859 (N_3859,In_1424,In_1038);
and U3860 (N_3860,In_1727,In_1079);
and U3861 (N_3861,In_65,In_1267);
or U3862 (N_3862,In_19,In_1394);
or U3863 (N_3863,In_108,In_1543);
and U3864 (N_3864,In_1597,In_863);
and U3865 (N_3865,In_1246,In_312);
and U3866 (N_3866,In_693,In_1246);
or U3867 (N_3867,In_1478,In_870);
nand U3868 (N_3868,In_486,In_1864);
or U3869 (N_3869,In_1629,In_1259);
xor U3870 (N_3870,In_747,In_1307);
nor U3871 (N_3871,In_266,In_1824);
or U3872 (N_3872,In_191,In_1080);
nand U3873 (N_3873,In_91,In_453);
or U3874 (N_3874,In_300,In_963);
and U3875 (N_3875,In_1904,In_300);
nand U3876 (N_3876,In_280,In_1505);
nor U3877 (N_3877,In_12,In_1633);
nand U3878 (N_3878,In_1154,In_156);
nand U3879 (N_3879,In_38,In_700);
nand U3880 (N_3880,In_903,In_1148);
and U3881 (N_3881,In_1355,In_1176);
xor U3882 (N_3882,In_337,In_62);
or U3883 (N_3883,In_970,In_1451);
or U3884 (N_3884,In_1140,In_1337);
nand U3885 (N_3885,In_963,In_1462);
nand U3886 (N_3886,In_280,In_1824);
and U3887 (N_3887,In_1419,In_1479);
or U3888 (N_3888,In_1900,In_1065);
and U3889 (N_3889,In_1786,In_1591);
or U3890 (N_3890,In_1633,In_418);
xnor U3891 (N_3891,In_290,In_1962);
and U3892 (N_3892,In_1735,In_615);
and U3893 (N_3893,In_1086,In_1667);
nand U3894 (N_3894,In_902,In_1532);
xnor U3895 (N_3895,In_1715,In_122);
nand U3896 (N_3896,In_536,In_1035);
nor U3897 (N_3897,In_468,In_135);
or U3898 (N_3898,In_1132,In_682);
or U3899 (N_3899,In_157,In_485);
or U3900 (N_3900,In_1383,In_1601);
or U3901 (N_3901,In_1,In_1341);
nor U3902 (N_3902,In_1770,In_35);
and U3903 (N_3903,In_1726,In_363);
nor U3904 (N_3904,In_1908,In_772);
nand U3905 (N_3905,In_1192,In_1291);
nand U3906 (N_3906,In_522,In_557);
nor U3907 (N_3907,In_146,In_575);
nand U3908 (N_3908,In_1926,In_792);
nand U3909 (N_3909,In_694,In_1053);
and U3910 (N_3910,In_981,In_170);
nor U3911 (N_3911,In_133,In_1195);
and U3912 (N_3912,In_1692,In_1373);
and U3913 (N_3913,In_1071,In_80);
or U3914 (N_3914,In_279,In_323);
or U3915 (N_3915,In_360,In_1021);
and U3916 (N_3916,In_1950,In_1519);
nor U3917 (N_3917,In_1850,In_780);
nand U3918 (N_3918,In_1468,In_1446);
or U3919 (N_3919,In_455,In_1576);
nor U3920 (N_3920,In_149,In_1274);
and U3921 (N_3921,In_501,In_1145);
or U3922 (N_3922,In_1555,In_937);
nand U3923 (N_3923,In_891,In_1558);
nor U3924 (N_3924,In_718,In_942);
nand U3925 (N_3925,In_1273,In_1724);
and U3926 (N_3926,In_1426,In_202);
or U3927 (N_3927,In_1460,In_58);
nor U3928 (N_3928,In_795,In_553);
or U3929 (N_3929,In_1784,In_1210);
or U3930 (N_3930,In_1997,In_514);
or U3931 (N_3931,In_437,In_1519);
and U3932 (N_3932,In_295,In_679);
nor U3933 (N_3933,In_468,In_1138);
nor U3934 (N_3934,In_755,In_1849);
or U3935 (N_3935,In_115,In_118);
nor U3936 (N_3936,In_1224,In_1240);
nand U3937 (N_3937,In_1217,In_1141);
or U3938 (N_3938,In_853,In_195);
nand U3939 (N_3939,In_1129,In_1592);
nand U3940 (N_3940,In_1178,In_1199);
nand U3941 (N_3941,In_784,In_128);
and U3942 (N_3942,In_954,In_1654);
and U3943 (N_3943,In_943,In_1080);
and U3944 (N_3944,In_22,In_817);
nor U3945 (N_3945,In_982,In_1027);
and U3946 (N_3946,In_184,In_1745);
nand U3947 (N_3947,In_1172,In_1404);
and U3948 (N_3948,In_1875,In_1804);
nor U3949 (N_3949,In_1253,In_51);
and U3950 (N_3950,In_1148,In_1287);
and U3951 (N_3951,In_385,In_112);
or U3952 (N_3952,In_1133,In_1733);
and U3953 (N_3953,In_1100,In_1313);
nand U3954 (N_3954,In_522,In_1283);
nand U3955 (N_3955,In_836,In_224);
nand U3956 (N_3956,In_1916,In_836);
or U3957 (N_3957,In_661,In_33);
xnor U3958 (N_3958,In_1338,In_175);
nand U3959 (N_3959,In_53,In_224);
nor U3960 (N_3960,In_1009,In_993);
nand U3961 (N_3961,In_1629,In_186);
or U3962 (N_3962,In_1990,In_1613);
and U3963 (N_3963,In_637,In_127);
or U3964 (N_3964,In_1073,In_1718);
and U3965 (N_3965,In_1709,In_1366);
nand U3966 (N_3966,In_275,In_1906);
and U3967 (N_3967,In_184,In_1517);
nor U3968 (N_3968,In_1254,In_1108);
and U3969 (N_3969,In_1655,In_816);
or U3970 (N_3970,In_1155,In_1780);
nor U3971 (N_3971,In_341,In_165);
nand U3972 (N_3972,In_1532,In_691);
nor U3973 (N_3973,In_989,In_674);
or U3974 (N_3974,In_1089,In_807);
nor U3975 (N_3975,In_665,In_875);
nand U3976 (N_3976,In_1686,In_1085);
nand U3977 (N_3977,In_1525,In_653);
nor U3978 (N_3978,In_1817,In_1574);
and U3979 (N_3979,In_100,In_1180);
nand U3980 (N_3980,In_231,In_430);
or U3981 (N_3981,In_290,In_1423);
nand U3982 (N_3982,In_1653,In_1579);
nor U3983 (N_3983,In_1745,In_499);
xnor U3984 (N_3984,In_744,In_420);
or U3985 (N_3985,In_881,In_1654);
and U3986 (N_3986,In_1161,In_439);
or U3987 (N_3987,In_628,In_443);
and U3988 (N_3988,In_921,In_136);
and U3989 (N_3989,In_1374,In_119);
nor U3990 (N_3990,In_542,In_1740);
and U3991 (N_3991,In_1571,In_1227);
nor U3992 (N_3992,In_149,In_257);
or U3993 (N_3993,In_1416,In_1084);
or U3994 (N_3994,In_406,In_1547);
or U3995 (N_3995,In_657,In_279);
or U3996 (N_3996,In_1238,In_1990);
or U3997 (N_3997,In_528,In_1123);
or U3998 (N_3998,In_1602,In_1579);
and U3999 (N_3999,In_1593,In_530);
nand U4000 (N_4000,N_2023,N_2054);
or U4001 (N_4001,N_1132,N_199);
and U4002 (N_4002,N_2289,N_2490);
and U4003 (N_4003,N_1272,N_3046);
and U4004 (N_4004,N_2193,N_1677);
nand U4005 (N_4005,N_3317,N_384);
nor U4006 (N_4006,N_3224,N_3088);
nor U4007 (N_4007,N_389,N_1489);
or U4008 (N_4008,N_3754,N_1765);
or U4009 (N_4009,N_1046,N_1153);
or U4010 (N_4010,N_1012,N_2301);
nor U4011 (N_4011,N_3261,N_382);
or U4012 (N_4012,N_2581,N_824);
nand U4013 (N_4013,N_2218,N_2880);
or U4014 (N_4014,N_1081,N_1374);
nor U4015 (N_4015,N_3844,N_147);
and U4016 (N_4016,N_3057,N_2883);
or U4017 (N_4017,N_2322,N_235);
nor U4018 (N_4018,N_1303,N_2374);
and U4019 (N_4019,N_2814,N_2402);
and U4020 (N_4020,N_2905,N_247);
or U4021 (N_4021,N_28,N_785);
and U4022 (N_4022,N_3839,N_2793);
or U4023 (N_4023,N_3586,N_372);
or U4024 (N_4024,N_530,N_1842);
or U4025 (N_4025,N_3535,N_2435);
xnor U4026 (N_4026,N_313,N_1898);
nor U4027 (N_4027,N_2889,N_821);
nand U4028 (N_4028,N_3903,N_2148);
or U4029 (N_4029,N_712,N_3333);
and U4030 (N_4030,N_933,N_221);
or U4031 (N_4031,N_3705,N_2760);
nor U4032 (N_4032,N_2418,N_3939);
or U4033 (N_4033,N_3611,N_604);
or U4034 (N_4034,N_2354,N_1942);
nor U4035 (N_4035,N_1028,N_1950);
xnor U4036 (N_4036,N_2529,N_85);
nand U4037 (N_4037,N_1503,N_2671);
or U4038 (N_4038,N_3455,N_1360);
xor U4039 (N_4039,N_248,N_3554);
and U4040 (N_4040,N_1876,N_2875);
nor U4041 (N_4041,N_1596,N_1837);
nand U4042 (N_4042,N_1983,N_1205);
or U4043 (N_4043,N_153,N_829);
or U4044 (N_4044,N_2752,N_1108);
and U4045 (N_4045,N_2300,N_2429);
nor U4046 (N_4046,N_1770,N_2086);
or U4047 (N_4047,N_383,N_1748);
nand U4048 (N_4048,N_1970,N_3485);
or U4049 (N_4049,N_3559,N_2226);
or U4050 (N_4050,N_3159,N_1252);
nor U4051 (N_4051,N_2488,N_84);
nor U4052 (N_4052,N_490,N_1952);
or U4053 (N_4053,N_168,N_718);
or U4054 (N_4054,N_511,N_1811);
or U4055 (N_4055,N_3603,N_112);
nor U4056 (N_4056,N_2820,N_913);
nand U4057 (N_4057,N_207,N_2634);
and U4058 (N_4058,N_2512,N_1756);
and U4059 (N_4059,N_3030,N_356);
and U4060 (N_4060,N_537,N_3096);
nand U4061 (N_4061,N_1921,N_569);
nor U4062 (N_4062,N_3583,N_2776);
nor U4063 (N_4063,N_3541,N_2768);
or U4064 (N_4064,N_2405,N_100);
nand U4065 (N_4065,N_1783,N_1328);
or U4066 (N_4066,N_3923,N_1008);
nor U4067 (N_4067,N_2244,N_2932);
and U4068 (N_4068,N_2697,N_2773);
nor U4069 (N_4069,N_3153,N_752);
nand U4070 (N_4070,N_1137,N_1248);
or U4071 (N_4071,N_3548,N_981);
nand U4072 (N_4072,N_231,N_1389);
nor U4073 (N_4073,N_3335,N_3824);
nor U4074 (N_4074,N_332,N_2891);
or U4075 (N_4075,N_425,N_872);
and U4076 (N_4076,N_1135,N_1126);
and U4077 (N_4077,N_2770,N_1804);
and U4078 (N_4078,N_3790,N_1053);
and U4079 (N_4079,N_2794,N_1242);
nor U4080 (N_4080,N_1738,N_3181);
nor U4081 (N_4081,N_1468,N_1515);
nand U4082 (N_4082,N_3276,N_1334);
and U4083 (N_4083,N_1199,N_2598);
and U4084 (N_4084,N_1647,N_150);
or U4085 (N_4085,N_1999,N_2310);
or U4086 (N_4086,N_1814,N_721);
or U4087 (N_4087,N_3066,N_155);
nor U4088 (N_4088,N_2135,N_2816);
or U4089 (N_4089,N_395,N_438);
nand U4090 (N_4090,N_246,N_2040);
and U4091 (N_4091,N_2616,N_2569);
nand U4092 (N_4092,N_454,N_2319);
nor U4093 (N_4093,N_3841,N_3697);
nand U4094 (N_4094,N_1116,N_539);
and U4095 (N_4095,N_2214,N_3174);
or U4096 (N_4096,N_1339,N_3718);
and U4097 (N_4097,N_3119,N_141);
and U4098 (N_4098,N_1160,N_698);
xnor U4099 (N_4099,N_1522,N_3629);
and U4100 (N_4100,N_1196,N_1279);
and U4101 (N_4101,N_2041,N_573);
nor U4102 (N_4102,N_720,N_3749);
nor U4103 (N_4103,N_2727,N_949);
or U4104 (N_4104,N_3454,N_2309);
and U4105 (N_4105,N_1225,N_892);
nor U4106 (N_4106,N_1107,N_781);
nor U4107 (N_4107,N_3378,N_368);
or U4108 (N_4108,N_3807,N_2571);
nor U4109 (N_4109,N_1971,N_1332);
nand U4110 (N_4110,N_1250,N_2828);
nand U4111 (N_4111,N_1633,N_2717);
and U4112 (N_4112,N_729,N_3550);
nand U4113 (N_4113,N_1749,N_503);
nor U4114 (N_4114,N_3873,N_2120);
or U4115 (N_4115,N_1384,N_607);
nand U4116 (N_4116,N_1678,N_411);
nand U4117 (N_4117,N_3228,N_1056);
nand U4118 (N_4118,N_2747,N_3917);
nand U4119 (N_4119,N_423,N_982);
nor U4120 (N_4120,N_1266,N_955);
nor U4121 (N_4121,N_2343,N_2272);
nand U4122 (N_4122,N_2293,N_2826);
or U4123 (N_4123,N_1015,N_2583);
nor U4124 (N_4124,N_2792,N_268);
nor U4125 (N_4125,N_629,N_3644);
nor U4126 (N_4126,N_2029,N_1085);
and U4127 (N_4127,N_188,N_518);
and U4128 (N_4128,N_2779,N_189);
or U4129 (N_4129,N_2712,N_3270);
xor U4130 (N_4130,N_1230,N_1855);
xor U4131 (N_4131,N_1551,N_3205);
and U4132 (N_4132,N_916,N_1792);
nand U4133 (N_4133,N_678,N_253);
and U4134 (N_4134,N_1895,N_2213);
nor U4135 (N_4135,N_2075,N_2073);
and U4136 (N_4136,N_3955,N_2657);
and U4137 (N_4137,N_804,N_3471);
or U4138 (N_4138,N_2335,N_1307);
and U4139 (N_4139,N_1350,N_462);
nor U4140 (N_4140,N_703,N_828);
nor U4141 (N_4141,N_2686,N_2927);
and U4142 (N_4142,N_2548,N_622);
nand U4143 (N_4143,N_2359,N_2922);
xor U4144 (N_4144,N_1233,N_3125);
and U4145 (N_4145,N_324,N_3290);
and U4146 (N_4146,N_2401,N_2476);
nand U4147 (N_4147,N_3770,N_1101);
nor U4148 (N_4148,N_2325,N_2945);
and U4149 (N_4149,N_1484,N_3621);
or U4150 (N_4150,N_1818,N_2497);
and U4151 (N_4151,N_1431,N_3695);
nand U4152 (N_4152,N_1645,N_637);
nand U4153 (N_4153,N_1306,N_1905);
and U4154 (N_4154,N_3899,N_2524);
and U4155 (N_4155,N_840,N_2454);
nor U4156 (N_4156,N_544,N_1962);
nor U4157 (N_4157,N_1165,N_1981);
and U4158 (N_4158,N_3085,N_1669);
or U4159 (N_4159,N_2140,N_2898);
nor U4160 (N_4160,N_1093,N_2234);
nor U4161 (N_4161,N_1612,N_2582);
nor U4162 (N_4162,N_364,N_3528);
and U4163 (N_4163,N_3787,N_2836);
nand U4164 (N_4164,N_1414,N_405);
and U4165 (N_4165,N_1260,N_2229);
and U4166 (N_4166,N_3287,N_1540);
nor U4167 (N_4167,N_1002,N_1603);
nand U4168 (N_4168,N_512,N_780);
nand U4169 (N_4169,N_2378,N_2566);
nor U4170 (N_4170,N_1967,N_1773);
nor U4171 (N_4171,N_1437,N_2132);
nand U4172 (N_4172,N_1371,N_2740);
and U4173 (N_4173,N_3590,N_1941);
or U4174 (N_4174,N_1675,N_2703);
and U4175 (N_4175,N_1278,N_289);
nor U4176 (N_4176,N_3039,N_3896);
nor U4177 (N_4177,N_1890,N_1760);
nor U4178 (N_4178,N_521,N_2643);
and U4179 (N_4179,N_360,N_2459);
or U4180 (N_4180,N_3238,N_1398);
nor U4181 (N_4181,N_2406,N_1104);
and U4182 (N_4182,N_3376,N_1471);
nor U4183 (N_4183,N_3431,N_853);
and U4184 (N_4184,N_3552,N_1672);
or U4185 (N_4185,N_1822,N_789);
nand U4186 (N_4186,N_3874,N_1395);
nand U4187 (N_4187,N_889,N_186);
or U4188 (N_4188,N_2388,N_16);
xor U4189 (N_4189,N_3828,N_3625);
and U4190 (N_4190,N_2978,N_2101);
nor U4191 (N_4191,N_448,N_2914);
and U4192 (N_4192,N_1416,N_3043);
nand U4193 (N_4193,N_2166,N_3194);
or U4194 (N_4194,N_2312,N_3734);
nand U4195 (N_4195,N_3010,N_1387);
xor U4196 (N_4196,N_434,N_3231);
and U4197 (N_4197,N_3155,N_200);
xor U4198 (N_4198,N_3446,N_2267);
or U4199 (N_4199,N_3257,N_398);
or U4200 (N_4200,N_3493,N_2552);
nand U4201 (N_4201,N_3916,N_2735);
nor U4202 (N_4202,N_1314,N_922);
and U4203 (N_4203,N_798,N_394);
or U4204 (N_4204,N_3669,N_1772);
or U4205 (N_4205,N_3936,N_414);
nand U4206 (N_4206,N_1826,N_2726);
nand U4207 (N_4207,N_103,N_2540);
or U4208 (N_4208,N_3819,N_2573);
and U4209 (N_4209,N_2645,N_3064);
and U4210 (N_4210,N_2460,N_1894);
nor U4211 (N_4211,N_1936,N_1537);
nor U4212 (N_4212,N_3112,N_2580);
xor U4213 (N_4213,N_225,N_652);
nor U4214 (N_4214,N_82,N_764);
or U4215 (N_4215,N_2420,N_3750);
or U4216 (N_4216,N_1037,N_3310);
nand U4217 (N_4217,N_3211,N_3392);
nand U4218 (N_4218,N_3811,N_3608);
and U4219 (N_4219,N_1327,N_165);
and U4220 (N_4220,N_2980,N_1400);
or U4221 (N_4221,N_2757,N_1906);
nand U4222 (N_4222,N_3143,N_1102);
nor U4223 (N_4223,N_2655,N_2968);
nand U4224 (N_4224,N_2926,N_1901);
or U4225 (N_4225,N_3018,N_309);
nor U4226 (N_4226,N_3078,N_1179);
nor U4227 (N_4227,N_3626,N_3662);
nand U4228 (N_4228,N_192,N_2186);
nand U4229 (N_4229,N_292,N_3624);
nor U4230 (N_4230,N_2182,N_1685);
nand U4231 (N_4231,N_3262,N_2038);
nand U4232 (N_4232,N_3729,N_2147);
and U4233 (N_4233,N_1791,N_3022);
and U4234 (N_4234,N_3459,N_3145);
and U4235 (N_4235,N_3236,N_3822);
and U4236 (N_4236,N_19,N_2844);
nand U4237 (N_4237,N_353,N_3977);
nor U4238 (N_4238,N_1009,N_592);
or U4239 (N_4239,N_571,N_3014);
and U4240 (N_4240,N_3,N_1361);
nor U4241 (N_4241,N_3052,N_2434);
or U4242 (N_4242,N_3881,N_3645);
or U4243 (N_4243,N_1476,N_2651);
or U4244 (N_4244,N_1530,N_33);
xnor U4245 (N_4245,N_457,N_1638);
nor U4246 (N_4246,N_610,N_1907);
and U4247 (N_4247,N_3732,N_3233);
or U4248 (N_4248,N_3715,N_583);
and U4249 (N_4249,N_2323,N_1594);
nor U4250 (N_4250,N_2718,N_1899);
or U4251 (N_4251,N_3038,N_208);
xor U4252 (N_4252,N_567,N_2840);
nor U4253 (N_4253,N_2257,N_1316);
nor U4254 (N_4254,N_868,N_2425);
nand U4255 (N_4255,N_2610,N_1459);
xnor U4256 (N_4256,N_1203,N_1856);
nor U4257 (N_4257,N_2494,N_2924);
or U4258 (N_4258,N_3445,N_2282);
nand U4259 (N_4259,N_3515,N_2992);
nor U4260 (N_4260,N_838,N_1340);
and U4261 (N_4261,N_2242,N_3756);
or U4262 (N_4262,N_426,N_174);
and U4263 (N_4263,N_2827,N_1946);
nor U4264 (N_4264,N_31,N_2716);
and U4265 (N_4265,N_3938,N_3968);
nor U4266 (N_4266,N_3309,N_3922);
or U4267 (N_4267,N_790,N_2129);
or U4268 (N_4268,N_2500,N_2138);
and U4269 (N_4269,N_3539,N_627);
nand U4270 (N_4270,N_3544,N_391);
and U4271 (N_4271,N_3855,N_1172);
xor U4272 (N_4272,N_3967,N_1824);
or U4273 (N_4273,N_3373,N_588);
nor U4274 (N_4274,N_3131,N_3067);
or U4275 (N_4275,N_1070,N_1428);
nor U4276 (N_4276,N_3104,N_1424);
xor U4277 (N_4277,N_3651,N_224);
and U4278 (N_4278,N_2404,N_3845);
and U4279 (N_4279,N_527,N_1246);
and U4280 (N_4280,N_990,N_3792);
or U4281 (N_4281,N_119,N_1615);
or U4282 (N_4282,N_418,N_3053);
nor U4283 (N_4283,N_1680,N_2611);
or U4284 (N_4284,N_2764,N_707);
and U4285 (N_4285,N_3793,N_3639);
and U4286 (N_4286,N_3566,N_1308);
or U4287 (N_4287,N_1485,N_1665);
and U4288 (N_4288,N_3154,N_3298);
or U4289 (N_4289,N_582,N_2155);
nand U4290 (N_4290,N_1805,N_2094);
nand U4291 (N_4291,N_2277,N_3109);
and U4292 (N_4292,N_3138,N_2532);
and U4293 (N_4293,N_687,N_1376);
nand U4294 (N_4294,N_2266,N_3612);
and U4295 (N_4295,N_2884,N_494);
nand U4296 (N_4296,N_1174,N_996);
or U4297 (N_4297,N_1052,N_3398);
or U4298 (N_4298,N_2991,N_2984);
nor U4299 (N_4299,N_1573,N_1456);
nor U4300 (N_4300,N_1682,N_603);
or U4301 (N_4301,N_506,N_3008);
nand U4302 (N_4302,N_879,N_2360);
and U4303 (N_4303,N_867,N_3274);
or U4304 (N_4304,N_1202,N_965);
nor U4305 (N_4305,N_1336,N_3685);
nor U4306 (N_4306,N_3055,N_624);
nor U4307 (N_4307,N_1114,N_270);
and U4308 (N_4308,N_1741,N_3217);
or U4309 (N_4309,N_1227,N_3707);
or U4310 (N_4310,N_3998,N_668);
and U4311 (N_4311,N_311,N_3420);
nor U4312 (N_4312,N_338,N_3883);
nand U4313 (N_4313,N_815,N_2625);
nor U4314 (N_4314,N_3489,N_3306);
nand U4315 (N_4315,N_3688,N_412);
nand U4316 (N_4316,N_3061,N_1852);
nor U4317 (N_4317,N_3383,N_3268);
and U4318 (N_4318,N_1061,N_377);
nand U4319 (N_4319,N_3313,N_2595);
or U4320 (N_4320,N_677,N_1069);
nand U4321 (N_4321,N_2578,N_3964);
nor U4322 (N_4322,N_1452,N_615);
xnor U4323 (N_4323,N_1018,N_3056);
nor U4324 (N_4324,N_86,N_3779);
nor U4325 (N_4325,N_1536,N_3269);
xnor U4326 (N_4326,N_859,N_644);
nor U4327 (N_4327,N_3457,N_3180);
nand U4328 (N_4328,N_670,N_1978);
nor U4329 (N_4329,N_2422,N_1211);
nor U4330 (N_4330,N_2302,N_1917);
nor U4331 (N_4331,N_2077,N_279);
or U4332 (N_4332,N_3585,N_3843);
nand U4333 (N_4333,N_3385,N_1925);
and U4334 (N_4334,N_1241,N_2877);
or U4335 (N_4335,N_3912,N_3854);
or U4336 (N_4336,N_2846,N_198);
nand U4337 (N_4337,N_3555,N_3797);
nand U4338 (N_4338,N_3579,N_685);
or U4339 (N_4339,N_1695,N_1825);
or U4340 (N_4340,N_69,N_2367);
and U4341 (N_4341,N_848,N_3692);
nand U4342 (N_4342,N_2079,N_3432);
and U4343 (N_4343,N_1446,N_495);
and U4344 (N_4344,N_1236,N_38);
nand U4345 (N_4345,N_710,N_525);
or U4346 (N_4346,N_3108,N_2538);
or U4347 (N_4347,N_3725,N_3635);
or U4348 (N_4348,N_3777,N_1684);
and U4349 (N_4349,N_380,N_3696);
nand U4350 (N_4350,N_1284,N_1560);
xnor U4351 (N_4351,N_1257,N_1930);
or U4352 (N_4352,N_29,N_736);
and U4353 (N_4353,N_1388,N_2894);
nand U4354 (N_4354,N_2585,N_3142);
nand U4355 (N_4355,N_3470,N_726);
nor U4356 (N_4356,N_2004,N_57);
or U4357 (N_4357,N_745,N_2890);
nand U4358 (N_4358,N_3524,N_3375);
nand U4359 (N_4359,N_1105,N_3760);
nor U4360 (N_4360,N_971,N_1091);
or U4361 (N_4361,N_1819,N_3202);
xor U4362 (N_4362,N_167,N_580);
or U4363 (N_4363,N_2925,N_941);
nor U4364 (N_4364,N_3122,N_3694);
xor U4365 (N_4365,N_2204,N_3935);
nor U4366 (N_4366,N_267,N_1466);
and U4367 (N_4367,N_271,N_541);
or U4368 (N_4368,N_2111,N_1863);
and U4369 (N_4369,N_1687,N_2142);
and U4370 (N_4370,N_2803,N_1705);
nand U4371 (N_4371,N_3124,N_2505);
and U4372 (N_4372,N_754,N_3486);
and U4373 (N_4373,N_2192,N_3927);
nor U4374 (N_4374,N_2996,N_1535);
nand U4375 (N_4375,N_915,N_20);
nand U4376 (N_4376,N_2995,N_1832);
and U4377 (N_4377,N_3263,N_2307);
nand U4378 (N_4378,N_3965,N_1088);
nand U4379 (N_4379,N_406,N_1106);
and U4380 (N_4380,N_963,N_3011);
or U4381 (N_4381,N_44,N_3895);
xnor U4382 (N_4382,N_2919,N_3944);
and U4383 (N_4383,N_1673,N_3774);
or U4384 (N_4384,N_466,N_1419);
or U4385 (N_4385,N_929,N_1382);
nand U4386 (N_4386,N_3160,N_1843);
and U4387 (N_4387,N_2543,N_3784);
xor U4388 (N_4388,N_3752,N_694);
nand U4389 (N_4389,N_1933,N_2334);
nor U4390 (N_4390,N_3768,N_3834);
or U4391 (N_4391,N_2839,N_1963);
nand U4392 (N_4392,N_645,N_2818);
and U4393 (N_4393,N_433,N_113);
or U4394 (N_4394,N_1555,N_58);
nand U4395 (N_4395,N_706,N_2994);
nand U4396 (N_4396,N_2184,N_2949);
or U4397 (N_4397,N_2713,N_1755);
and U4398 (N_4398,N_2921,N_2346);
and U4399 (N_4399,N_612,N_3092);
or U4400 (N_4400,N_3337,N_2613);
and U4401 (N_4401,N_3002,N_866);
or U4402 (N_4402,N_2461,N_304);
or U4403 (N_4403,N_3817,N_1816);
or U4404 (N_4404,N_2896,N_2276);
or U4405 (N_4405,N_301,N_171);
nand U4406 (N_4406,N_522,N_2862);
nor U4407 (N_4407,N_327,N_683);
nand U4408 (N_4408,N_3571,N_3703);
xor U4409 (N_4409,N_621,N_2108);
and U4410 (N_4410,N_3213,N_1637);
nor U4411 (N_4411,N_430,N_3886);
and U4412 (N_4412,N_458,N_1984);
nor U4413 (N_4413,N_2572,N_449);
or U4414 (N_4414,N_1130,N_2666);
nor U4415 (N_4415,N_2369,N_3389);
and U4416 (N_4416,N_1482,N_2899);
nor U4417 (N_4417,N_2467,N_3832);
or U4418 (N_4418,N_2270,N_1838);
nor U4419 (N_4419,N_1142,N_792);
nor U4420 (N_4420,N_1289,N_3381);
and U4421 (N_4421,N_954,N_2593);
nand U4422 (N_4422,N_1062,N_2551);
or U4423 (N_4423,N_3478,N_2834);
nor U4424 (N_4424,N_1644,N_375);
nand U4425 (N_4425,N_648,N_777);
nand U4426 (N_4426,N_126,N_134);
nor U4427 (N_4427,N_3821,N_3163);
nand U4428 (N_4428,N_146,N_1293);
nor U4429 (N_4429,N_1888,N_1910);
nand U4430 (N_4430,N_2442,N_379);
and U4431 (N_4431,N_3435,N_1977);
nor U4432 (N_4432,N_1063,N_1193);
and U4433 (N_4433,N_3168,N_3032);
and U4434 (N_4434,N_2897,N_3012);
and U4435 (N_4435,N_1457,N_3034);
nor U4436 (N_4436,N_2384,N_3058);
and U4437 (N_4437,N_993,N_1486);
and U4438 (N_4438,N_96,N_2305);
nor U4439 (N_4439,N_1239,N_1996);
and U4440 (N_4440,N_3556,N_1604);
nand U4441 (N_4441,N_318,N_222);
or U4442 (N_4442,N_3812,N_118);
nand U4443 (N_4443,N_1924,N_1606);
nand U4444 (N_4444,N_299,N_1393);
nor U4445 (N_4445,N_2102,N_984);
nand U4446 (N_4446,N_3746,N_1874);
and U4447 (N_4447,N_1681,N_1976);
nor U4448 (N_4448,N_464,N_3201);
nand U4449 (N_4449,N_3506,N_2414);
and U4450 (N_4450,N_3818,N_106);
and U4451 (N_4451,N_601,N_839);
nand U4452 (N_4452,N_809,N_2046);
or U4453 (N_4453,N_133,N_3670);
nand U4454 (N_4454,N_2971,N_3364);
nand U4455 (N_4455,N_1251,N_3837);
or U4456 (N_4456,N_2190,N_3733);
nor U4457 (N_4457,N_3962,N_937);
nand U4458 (N_4458,N_811,N_1432);
or U4459 (N_4459,N_3350,N_316);
or U4460 (N_4460,N_3204,N_87);
or U4461 (N_4461,N_2621,N_442);
nand U4462 (N_4462,N_1571,N_1462);
nor U4463 (N_4463,N_3177,N_953);
and U4464 (N_4464,N_1379,N_1143);
nand U4465 (N_4465,N_2531,N_3116);
nand U4466 (N_4466,N_3076,N_3570);
xnor U4467 (N_4467,N_2523,N_3026);
nor U4468 (N_4468,N_2791,N_3315);
nor U4469 (N_4469,N_2262,N_3588);
or U4470 (N_4470,N_1528,N_3241);
nor U4471 (N_4471,N_1483,N_2471);
nor U4472 (N_4472,N_2953,N_3465);
xor U4473 (N_4473,N_856,N_2944);
and U4474 (N_4474,N_1733,N_2099);
nand U4475 (N_4475,N_2084,N_2853);
and U4476 (N_4476,N_326,N_1525);
nor U4477 (N_4477,N_3135,N_2855);
nor U4478 (N_4478,N_1312,N_3141);
or U4479 (N_4479,N_1879,N_2409);
and U4480 (N_4480,N_2096,N_3864);
and U4481 (N_4481,N_3618,N_1017);
nand U4482 (N_4482,N_3123,N_2246);
or U4483 (N_4483,N_3007,N_223);
or U4484 (N_4484,N_2854,N_203);
and U4485 (N_4485,N_3607,N_759);
and U4486 (N_4486,N_911,N_966);
and U4487 (N_4487,N_3074,N_3456);
nor U4488 (N_4488,N_3722,N_672);
nor U4489 (N_4489,N_553,N_2134);
nand U4490 (N_4490,N_1583,N_1858);
or U4491 (N_4491,N_3945,N_3304);
nor U4492 (N_4492,N_3103,N_197);
nor U4493 (N_4493,N_1399,N_4);
nand U4494 (N_4494,N_2823,N_2954);
nand U4495 (N_4495,N_2380,N_2179);
and U4496 (N_4496,N_2368,N_1508);
nand U4497 (N_4497,N_597,N_3995);
nand U4498 (N_4498,N_300,N_566);
nor U4499 (N_4499,N_381,N_2649);
nand U4500 (N_4500,N_3134,N_2599);
nor U4501 (N_4501,N_2131,N_3331);
nand U4502 (N_4502,N_2231,N_2462);
nor U4503 (N_4503,N_2588,N_1469);
nor U4504 (N_4504,N_2145,N_2088);
nand U4505 (N_4505,N_1763,N_3082);
nor U4506 (N_4506,N_3743,N_3069);
or U4507 (N_4507,N_517,N_1348);
and U4508 (N_4508,N_1690,N_3341);
nor U4509 (N_4509,N_3656,N_337);
nand U4510 (N_4510,N_2070,N_1718);
nor U4511 (N_4511,N_594,N_3152);
nor U4512 (N_4512,N_1566,N_3617);
xor U4513 (N_4513,N_3164,N_137);
nand U4514 (N_4514,N_2688,N_773);
or U4515 (N_4515,N_979,N_1402);
nor U4516 (N_4516,N_1329,N_2376);
nor U4517 (N_4517,N_1585,N_2714);
nor U4518 (N_4518,N_2181,N_3149);
nor U4519 (N_4519,N_2357,N_2452);
and U4520 (N_4520,N_2158,N_1993);
nor U4521 (N_4521,N_3305,N_887);
nor U4522 (N_4522,N_1192,N_2876);
nor U4523 (N_4523,N_2473,N_2603);
nor U4524 (N_4524,N_1627,N_705);
nor U4525 (N_4525,N_920,N_1703);
or U4526 (N_4526,N_3243,N_42);
nand U4527 (N_4527,N_3426,N_3804);
nand U4528 (N_4528,N_2985,N_3156);
or U4529 (N_4529,N_1164,N_3396);
nor U4530 (N_4530,N_1785,N_2344);
and U4531 (N_4531,N_501,N_1722);
nand U4532 (N_4532,N_74,N_3963);
nand U4533 (N_4533,N_1848,N_2423);
and U4534 (N_4534,N_2617,N_3953);
nor U4535 (N_4535,N_234,N_574);
or U4536 (N_4536,N_404,N_1287);
and U4537 (N_4537,N_2444,N_2050);
or U4538 (N_4538,N_1207,N_2910);
nor U4539 (N_4539,N_1719,N_56);
or U4540 (N_4540,N_1159,N_376);
nand U4541 (N_4541,N_2164,N_3724);
and U4542 (N_4542,N_385,N_1403);
and U4543 (N_4543,N_800,N_378);
and U4544 (N_4544,N_882,N_1441);
or U4545 (N_4545,N_2465,N_613);
nor U4546 (N_4546,N_3023,N_1189);
and U4547 (N_4547,N_3993,N_1417);
and U4548 (N_4548,N_1781,N_2769);
and U4549 (N_4549,N_7,N_2661);
nor U4550 (N_4550,N_156,N_1478);
or U4551 (N_4551,N_3551,N_2230);
nor U4552 (N_4552,N_2455,N_663);
nand U4553 (N_4553,N_2482,N_1198);
or U4554 (N_4554,N_1707,N_2126);
nand U4555 (N_4555,N_1157,N_3488);
or U4556 (N_4556,N_1529,N_148);
xnor U4557 (N_4557,N_3372,N_3356);
nand U4558 (N_4558,N_1454,N_1578);
nand U4559 (N_4559,N_2183,N_702);
nor U4560 (N_4560,N_3748,N_697);
nor U4561 (N_4561,N_2872,N_2081);
nand U4562 (N_4562,N_144,N_505);
nand U4563 (N_4563,N_325,N_631);
nand U4564 (N_4564,N_1200,N_2295);
nand U4565 (N_4565,N_3147,N_1881);
or U4566 (N_4566,N_2245,N_1181);
nand U4567 (N_4567,N_456,N_2200);
nor U4568 (N_4568,N_2169,N_761);
or U4569 (N_4569,N_802,N_3848);
or U4570 (N_4570,N_1026,N_1505);
xor U4571 (N_4571,N_986,N_2513);
nand U4572 (N_4572,N_2391,N_1068);
nor U4573 (N_4573,N_1351,N_1);
and U4574 (N_4574,N_3250,N_3979);
and U4575 (N_4575,N_3460,N_504);
nor U4576 (N_4576,N_2232,N_2669);
and U4577 (N_4577,N_806,N_1768);
nand U4578 (N_4578,N_2195,N_283);
and U4579 (N_4579,N_734,N_1857);
nand U4580 (N_4580,N_3780,N_181);
or U4581 (N_4581,N_1514,N_229);
or U4582 (N_4582,N_2412,N_3781);
and U4583 (N_4583,N_3636,N_1247);
or U4584 (N_4584,N_1405,N_2489);
nor U4585 (N_4585,N_3773,N_1591);
nor U4586 (N_4586,N_3437,N_1039);
or U4587 (N_4587,N_3782,N_657);
or U4588 (N_4588,N_794,N_121);
and U4589 (N_4589,N_640,N_487);
and U4590 (N_4590,N_2177,N_3235);
nand U4591 (N_4591,N_3678,N_408);
nor U4592 (N_4592,N_641,N_2563);
or U4593 (N_4593,N_1488,N_3740);
and U4594 (N_4594,N_54,N_543);
nand U4595 (N_4595,N_3706,N_2918);
or U4596 (N_4596,N_3862,N_475);
or U4597 (N_4597,N_2408,N_2100);
or U4598 (N_4598,N_2016,N_1273);
nand U4599 (N_4599,N_578,N_2981);
and U4600 (N_4600,N_1958,N_688);
nor U4601 (N_4601,N_2579,N_2674);
or U4602 (N_4602,N_595,N_485);
nor U4603 (N_4603,N_3424,N_3390);
and U4604 (N_4604,N_1470,N_3464);
and U4605 (N_4605,N_73,N_1296);
or U4606 (N_4606,N_2256,N_3139);
nor U4607 (N_4607,N_2052,N_2542);
nor U4608 (N_4608,N_814,N_139);
or U4609 (N_4609,N_2911,N_3189);
or U4610 (N_4610,N_1162,N_2732);
nor U4611 (N_4611,N_808,N_3190);
or U4612 (N_4612,N_2342,N_951);
or U4613 (N_4613,N_1083,N_1543);
or U4614 (N_4614,N_1372,N_2199);
and U4615 (N_4615,N_3942,N_3683);
and U4616 (N_4616,N_214,N_50);
and U4617 (N_4617,N_827,N_3910);
nor U4618 (N_4618,N_3300,N_575);
or U4619 (N_4619,N_1980,N_3004);
and U4620 (N_4620,N_348,N_782);
and U4621 (N_4621,N_3137,N_3671);
and U4622 (N_4622,N_2762,N_1709);
nor U4623 (N_4623,N_542,N_2701);
nor U4624 (N_4624,N_3025,N_861);
and U4625 (N_4625,N_2670,N_1493);
nor U4626 (N_4626,N_642,N_2665);
or U4627 (N_4627,N_770,N_1865);
nand U4628 (N_4628,N_3887,N_2537);
nor U4629 (N_4629,N_771,N_1846);
and U4630 (N_4630,N_2520,N_297);
nor U4631 (N_4631,N_1620,N_3596);
nor U4632 (N_4632,N_696,N_2515);
and U4633 (N_4633,N_3713,N_2832);
nor U4634 (N_4634,N_3869,N_170);
xor U4635 (N_4635,N_1623,N_1290);
or U4636 (N_4636,N_2336,N_959);
nor U4637 (N_4637,N_1343,N_3642);
nor U4638 (N_4638,N_2239,N_2110);
and U4639 (N_4639,N_534,N_3207);
and U4640 (N_4640,N_1531,N_3643);
or U4641 (N_4641,N_2136,N_3690);
and U4642 (N_4642,N_2594,N_273);
nand U4643 (N_4643,N_1067,N_3393);
nor U4644 (N_4644,N_2264,N_440);
nand U4645 (N_4645,N_646,N_1533);
nor U4646 (N_4646,N_2410,N_2392);
nand U4647 (N_4647,N_321,N_2011);
nand U4648 (N_4648,N_2445,N_1170);
and U4649 (N_4649,N_614,N_2092);
nor U4650 (N_4650,N_2511,N_158);
xor U4651 (N_4651,N_3831,N_769);
nand U4652 (N_4652,N_2206,N_3495);
or U4653 (N_4653,N_870,N_2091);
or U4654 (N_4654,N_2672,N_184);
or U4655 (N_4655,N_926,N_1830);
nand U4656 (N_4656,N_2268,N_12);
and U4657 (N_4657,N_826,N_1442);
or U4658 (N_4658,N_739,N_3438);
and U4659 (N_4659,N_1286,N_3829);
nor U4660 (N_4660,N_250,N_1982);
and U4661 (N_4661,N_3609,N_2753);
and U4662 (N_4662,N_2692,N_2729);
nor U4663 (N_4663,N_2350,N_2351);
nor U4664 (N_4664,N_2930,N_1504);
and U4665 (N_4665,N_2385,N_3271);
nand U4666 (N_4666,N_3117,N_676);
nand U4667 (N_4667,N_3753,N_2804);
nand U4668 (N_4668,N_2976,N_2225);
or U4669 (N_4669,N_1667,N_1556);
nor U4670 (N_4670,N_3195,N_3536);
and U4671 (N_4671,N_417,N_2887);
nand U4672 (N_4672,N_498,N_1264);
nor U4673 (N_4673,N_2650,N_2711);
and U4674 (N_4674,N_1282,N_3657);
nor U4675 (N_4675,N_2660,N_2125);
and U4676 (N_4676,N_122,N_958);
or U4677 (N_4677,N_2759,N_863);
nand U4678 (N_4678,N_742,N_1120);
or U4679 (N_4679,N_3425,N_943);
or U4680 (N_4680,N_1860,N_3266);
nand U4681 (N_4681,N_1447,N_1224);
or U4682 (N_4682,N_1323,N_1953);
and U4683 (N_4683,N_1268,N_3518);
nor U4684 (N_4684,N_3237,N_1346);
or U4685 (N_4685,N_2493,N_3599);
and U4686 (N_4686,N_1119,N_2825);
nor U4687 (N_4687,N_2358,N_3332);
or U4688 (N_4688,N_2781,N_1883);
nor U4689 (N_4689,N_927,N_909);
or U4690 (N_4690,N_3736,N_2294);
and U4691 (N_4691,N_473,N_989);
or U4692 (N_4692,N_1746,N_1050);
nor U4693 (N_4693,N_1201,N_3301);
nor U4694 (N_4694,N_2684,N_2039);
nor U4695 (N_4695,N_453,N_3291);
and U4696 (N_4696,N_2950,N_733);
nor U4697 (N_4697,N_2287,N_3846);
nor U4698 (N_4698,N_2977,N_2030);
and U4699 (N_4699,N_779,N_3986);
nand U4700 (N_4700,N_1909,N_635);
or U4701 (N_4701,N_2062,N_2530);
nor U4702 (N_4702,N_1373,N_3254);
and U4703 (N_4703,N_1380,N_2989);
nand U4704 (N_4704,N_446,N_3712);
nand U4705 (N_4705,N_2058,N_3484);
or U4706 (N_4706,N_2936,N_1550);
and U4707 (N_4707,N_3741,N_142);
nor U4708 (N_4708,N_2281,N_1902);
or U4709 (N_4709,N_3308,N_1025);
and U4710 (N_4710,N_1803,N_328);
xnor U4711 (N_4711,N_3654,N_623);
and U4712 (N_4712,N_3288,N_731);
and U4713 (N_4713,N_3162,N_2215);
nor U4714 (N_4714,N_923,N_2253);
and U4715 (N_4715,N_719,N_3472);
and U4716 (N_4716,N_114,N_3884);
nor U4717 (N_4717,N_1990,N_2208);
nand U4718 (N_4718,N_2328,N_3127);
or U4719 (N_4719,N_3297,N_3036);
nand U4720 (N_4720,N_903,N_709);
or U4721 (N_4721,N_2685,N_1743);
or U4722 (N_4722,N_1850,N_459);
or U4723 (N_4723,N_1775,N_1711);
or U4724 (N_4724,N_1960,N_3809);
nand U4725 (N_4725,N_1761,N_3188);
nor U4726 (N_4726,N_3118,N_2326);
and U4727 (N_4727,N_1599,N_2061);
nand U4728 (N_4728,N_1213,N_2372);
and U4729 (N_4729,N_2786,N_625);
or U4730 (N_4730,N_2998,N_547);
nor U4731 (N_4731,N_3397,N_2366);
or U4732 (N_4732,N_2049,N_3689);
or U4733 (N_4733,N_2498,N_3897);
and U4734 (N_4734,N_3028,N_3946);
or U4735 (N_4735,N_568,N_159);
and U4736 (N_4736,N_2441,N_1628);
nand U4737 (N_4737,N_820,N_227);
nand U4738 (N_4738,N_3042,N_1989);
and U4739 (N_4739,N_3623,N_886);
nor U4740 (N_4740,N_935,N_2106);
and U4741 (N_4741,N_210,N_2963);
nand U4742 (N_4742,N_1926,N_3033);
and U4743 (N_4743,N_3680,N_2093);
nor U4744 (N_4744,N_3380,N_2576);
nor U4745 (N_4745,N_1568,N_1509);
xor U4746 (N_4746,N_3496,N_2741);
and U4747 (N_4747,N_1121,N_2260);
or U4748 (N_4748,N_1048,N_2112);
nor U4749 (N_4749,N_2708,N_3653);
nor U4750 (N_4750,N_1892,N_682);
nand U4751 (N_4751,N_532,N_1590);
nand U4752 (N_4752,N_2830,N_3830);
or U4753 (N_4753,N_1517,N_3661);
and U4754 (N_4754,N_421,N_3747);
or U4755 (N_4755,N_900,N_917);
or U4756 (N_4756,N_2123,N_3704);
nand U4757 (N_4757,N_2533,N_2042);
nor U4758 (N_4758,N_3606,N_1139);
or U4759 (N_4759,N_1654,N_1129);
or U4760 (N_4760,N_3399,N_2623);
nor U4761 (N_4761,N_1782,N_1891);
nand U4762 (N_4762,N_1363,N_1877);
nand U4763 (N_4763,N_3200,N_2211);
or U4764 (N_4764,N_1968,N_2948);
or U4765 (N_4765,N_711,N_564);
nor U4766 (N_4766,N_1465,N_2715);
nand U4767 (N_4767,N_536,N_3448);
nor U4768 (N_4768,N_90,N_2178);
and U4769 (N_4769,N_2223,N_3299);
and U4770 (N_4770,N_2487,N_1735);
and U4771 (N_4771,N_738,N_1125);
and U4772 (N_4772,N_3835,N_2063);
nand U4773 (N_4773,N_2608,N_2197);
nand U4774 (N_4774,N_1261,N_1443);
and U4775 (N_4775,N_3650,N_2838);
nor U4776 (N_4776,N_2440,N_883);
nand U4777 (N_4777,N_437,N_3186);
nand U4778 (N_4778,N_2060,N_2541);
xor U4779 (N_4779,N_254,N_2025);
or U4780 (N_4780,N_2694,N_3958);
and U4781 (N_4781,N_823,N_2265);
nand U4782 (N_4782,N_2861,N_232);
or U4783 (N_4783,N_3111,N_2427);
nor U4784 (N_4784,N_1754,N_484);
and U4785 (N_4785,N_2349,N_3369);
or U4786 (N_4786,N_211,N_3226);
nand U4787 (N_4787,N_3320,N_1047);
and U4788 (N_4788,N_2782,N_950);
nand U4789 (N_4789,N_3987,N_3314);
nand U4790 (N_4790,N_228,N_2124);
xor U4791 (N_4791,N_143,N_13);
nand U4792 (N_4792,N_3087,N_3312);
or U4793 (N_4793,N_509,N_1277);
nand U4794 (N_4794,N_2469,N_3871);
or U4795 (N_4795,N_1689,N_2048);
or U4796 (N_4796,N_2730,N_486);
nand U4797 (N_4797,N_713,N_3853);
nand U4798 (N_4798,N_3719,N_2127);
xnor U4799 (N_4799,N_1911,N_1758);
nor U4800 (N_4800,N_2553,N_419);
or U4801 (N_4801,N_3950,N_2561);
or U4802 (N_4802,N_699,N_1629);
nand U4803 (N_4803,N_3569,N_1720);
nand U4804 (N_4804,N_1014,N_3342);
nand U4805 (N_4805,N_1322,N_215);
nor U4806 (N_4806,N_3996,N_2055);
and U4807 (N_4807,N_1030,N_2503);
nor U4808 (N_4808,N_3462,N_362);
and U4809 (N_4809,N_51,N_704);
and U4810 (N_4810,N_2290,N_1985);
and U4811 (N_4811,N_2939,N_1255);
and U4812 (N_4812,N_3441,N_3622);
and U4813 (N_4813,N_99,N_3591);
nand U4814 (N_4814,N_1561,N_3762);
and U4815 (N_4815,N_2419,N_2114);
nand U4816 (N_4816,N_1275,N_2986);
nor U4817 (N_4817,N_3500,N_1800);
and U4818 (N_4818,N_1650,N_343);
and U4819 (N_4819,N_3547,N_3847);
nor U4820 (N_4820,N_2878,N_2640);
nor U4821 (N_4821,N_1495,N_1082);
or U4822 (N_4822,N_3319,N_1292);
or U4823 (N_4823,N_845,N_765);
and U4824 (N_4824,N_3295,N_968);
nand U4825 (N_4825,N_2766,N_1000);
and U4826 (N_4826,N_132,N_1954);
nor U4827 (N_4827,N_2915,N_957);
nand U4828 (N_4828,N_1161,N_3562);
nor U4829 (N_4829,N_1074,N_1152);
and U4830 (N_4830,N_659,N_303);
and U4831 (N_4831,N_3481,N_2470);
nand U4832 (N_4832,N_1702,N_3717);
and U4833 (N_4833,N_3796,N_1674);
nand U4834 (N_4834,N_2118,N_1592);
and U4835 (N_4835,N_2577,N_2033);
or U4836 (N_4836,N_1096,N_2798);
nor U4837 (N_4837,N_3789,N_2612);
and U4838 (N_4838,N_1580,N_750);
and U4839 (N_4839,N_2706,N_3940);
nand U4840 (N_4840,N_3311,N_3165);
and U4841 (N_4841,N_3574,N_3763);
and U4842 (N_4842,N_3490,N_1058);
nand U4843 (N_4843,N_3336,N_2241);
nand U4844 (N_4844,N_2291,N_336);
nand U4845 (N_4845,N_674,N_1799);
nand U4846 (N_4846,N_409,N_3795);
and U4847 (N_4847,N_1586,N_2090);
and U4848 (N_4848,N_2528,N_312);
nand U4849 (N_4849,N_3400,N_3592);
nor U4850 (N_4850,N_550,N_3003);
or U4851 (N_4851,N_795,N_502);
and U4852 (N_4852,N_1226,N_1362);
or U4853 (N_4853,N_2034,N_1778);
nor U4854 (N_4854,N_2501,N_755);
and U4855 (N_4855,N_2031,N_556);
and U4856 (N_4856,N_2397,N_2678);
xor U4857 (N_4857,N_163,N_962);
or U4858 (N_4858,N_2037,N_3277);
nand U4859 (N_4859,N_2066,N_3983);
or U4860 (N_4860,N_2499,N_2690);
or U4861 (N_4861,N_40,N_1972);
and U4862 (N_4862,N_851,N_3294);
or U4863 (N_4863,N_3672,N_1657);
or U4864 (N_4864,N_2122,N_102);
or U4865 (N_4865,N_1966,N_744);
and U4866 (N_4866,N_91,N_3388);
or U4867 (N_4867,N_416,N_157);
or U4868 (N_4868,N_3070,N_3648);
nand U4869 (N_4869,N_1011,N_1280);
or U4870 (N_4870,N_88,N_2421);
xor U4871 (N_4871,N_1127,N_2345);
or U4872 (N_4872,N_2386,N_1234);
and U4873 (N_4873,N_1214,N_1502);
nor U4874 (N_4874,N_76,N_1238);
and U4875 (N_4875,N_1944,N_3913);
and U4876 (N_4876,N_700,N_298);
nand U4877 (N_4877,N_239,N_2733);
and U4878 (N_4878,N_901,N_918);
and U4879 (N_4879,N_62,N_125);
or U4880 (N_4880,N_489,N_1786);
and U4881 (N_4881,N_496,N_53);
nor U4882 (N_4882,N_3323,N_3932);
nand U4883 (N_4883,N_1408,N_784);
and U4884 (N_4884,N_1676,N_2098);
or U4885 (N_4885,N_2504,N_3737);
nand U4886 (N_4886,N_3889,N_884);
nor U4887 (N_4887,N_2203,N_1169);
and U4888 (N_4888,N_3852,N_175);
and U4889 (N_4889,N_1455,N_274);
and U4890 (N_4890,N_1923,N_1496);
nor U4891 (N_4891,N_519,N_1195);
nor U4892 (N_4892,N_632,N_1079);
nand U4893 (N_4893,N_2904,N_1145);
nor U4894 (N_4894,N_2702,N_1430);
nor U4895 (N_4895,N_1777,N_2704);
or U4896 (N_4896,N_1518,N_3560);
nand U4897 (N_4897,N_3197,N_1059);
or U4898 (N_4898,N_71,N_124);
nand U4899 (N_4899,N_1784,N_3387);
or U4900 (N_4900,N_2316,N_2162);
nor U4901 (N_4901,N_314,N_1163);
nand U4902 (N_4902,N_1410,N_1715);
and U4903 (N_4903,N_1448,N_3206);
and U4904 (N_4904,N_1131,N_2849);
or U4905 (N_4905,N_2361,N_3751);
nor U4906 (N_4906,N_3172,N_138);
or U4907 (N_4907,N_3814,N_1166);
or U4908 (N_4908,N_3503,N_3422);
nand U4909 (N_4909,N_1084,N_1563);
nand U4910 (N_4910,N_528,N_2920);
and U4911 (N_4911,N_2738,N_1191);
nand U4912 (N_4912,N_3150,N_275);
nand U4913 (N_4913,N_3015,N_1964);
or U4914 (N_4914,N_3423,N_584);
or U4915 (N_4915,N_747,N_3242);
and U4916 (N_4916,N_361,N_1487);
and U4917 (N_4917,N_346,N_2352);
nor U4918 (N_4918,N_2510,N_2586);
nand U4919 (N_4919,N_2982,N_2956);
nand U4920 (N_4920,N_701,N_2387);
nand U4921 (N_4921,N_2247,N_891);
or U4922 (N_4922,N_3498,N_2767);
or U4923 (N_4923,N_786,N_2749);
or U4924 (N_4924,N_3791,N_1961);
and U4925 (N_4925,N_1723,N_3245);
nand U4926 (N_4926,N_634,N_1222);
nor U4927 (N_4927,N_1574,N_1572);
or U4928 (N_4928,N_3876,N_3584);
and U4929 (N_4929,N_647,N_972);
or U4930 (N_4930,N_1378,N_18);
or U4931 (N_4931,N_857,N_1815);
nor U4932 (N_4932,N_1031,N_1249);
nor U4933 (N_4933,N_2619,N_3613);
nand U4934 (N_4934,N_3051,N_1270);
nand U4935 (N_4935,N_94,N_3384);
xnor U4936 (N_4936,N_2001,N_3664);
or U4937 (N_4937,N_2007,N_3416);
or U4938 (N_4938,N_1262,N_914);
xnor U4939 (N_4939,N_3575,N_3068);
xnor U4940 (N_4940,N_63,N_2065);
or U4941 (N_4941,N_1413,N_2235);
nand U4942 (N_4942,N_529,N_1019);
nor U4943 (N_4943,N_3355,N_2297);
nand U4944 (N_4944,N_78,N_1429);
nand U4945 (N_4945,N_3930,N_1662);
or U4946 (N_4946,N_2941,N_2189);
or U4947 (N_4947,N_1994,N_1696);
or U4948 (N_4948,N_470,N_2801);
or U4949 (N_4949,N_3915,N_3615);
nand U4950 (N_4950,N_1291,N_2026);
nand U4951 (N_4951,N_24,N_3788);
nand U4952 (N_4952,N_2687,N_2559);
or U4953 (N_4953,N_2519,N_2456);
or U4954 (N_4954,N_2864,N_491);
nand U4955 (N_4955,N_630,N_351);
xnor U4956 (N_4956,N_2448,N_1183);
nand U4957 (N_4957,N_1995,N_2654);
nor U4958 (N_4958,N_1742,N_236);
or U4959 (N_4959,N_3283,N_2144);
nor U4960 (N_4960,N_492,N_77);
and U4961 (N_4961,N_1802,N_2509);
nor U4962 (N_4962,N_2415,N_816);
nand U4963 (N_4963,N_1652,N_242);
xor U4964 (N_4964,N_1390,N_1115);
nand U4965 (N_4965,N_2705,N_835);
and U4966 (N_4966,N_152,N_3193);
nor U4967 (N_4967,N_2168,N_1510);
xnor U4968 (N_4968,N_2858,N_760);
nor U4969 (N_4969,N_2314,N_0);
and U4970 (N_4970,N_2338,N_269);
and U4971 (N_4971,N_1661,N_1171);
nor U4972 (N_4972,N_469,N_2154);
nor U4973 (N_4973,N_533,N_2159);
and U4974 (N_4974,N_3130,N_3196);
nand U4975 (N_4975,N_3009,N_1820);
or U4976 (N_4976,N_1136,N_1004);
and U4977 (N_4977,N_2139,N_2095);
xnor U4978 (N_4978,N_2824,N_3840);
or U4979 (N_4979,N_3395,N_3419);
and U4980 (N_4980,N_46,N_1956);
nand U4981 (N_4981,N_1147,N_2153);
nor U4982 (N_4982,N_3581,N_881);
and U4983 (N_4983,N_2085,N_3778);
nand U4984 (N_4984,N_3386,N_2584);
nor U4985 (N_4985,N_3783,N_3577);
and U4986 (N_4986,N_3045,N_1896);
nand U4987 (N_4987,N_193,N_2641);
or U4988 (N_4988,N_3906,N_259);
nand U4989 (N_4989,N_1117,N_1423);
and U4990 (N_4990,N_305,N_2765);
nand U4991 (N_4991,N_493,N_1729);
nor U4992 (N_4992,N_1807,N_2907);
or U4993 (N_4993,N_3285,N_2721);
nor U4994 (N_4994,N_1317,N_3776);
nand U4995 (N_4995,N_3595,N_3169);
nand U4996 (N_4996,N_633,N_743);
nor U4997 (N_4997,N_1281,N_2999);
nor U4998 (N_4998,N_2074,N_1732);
or U4999 (N_4999,N_910,N_2522);
nor U5000 (N_5000,N_128,N_2043);
nand U5001 (N_5001,N_2810,N_1112);
and U5002 (N_5002,N_2843,N_3861);
nand U5003 (N_5003,N_552,N_2217);
nand U5004 (N_5004,N_1893,N_3702);
nand U5005 (N_5005,N_2008,N_1725);
nand U5006 (N_5006,N_1407,N_1182);
nor U5007 (N_5007,N_2464,N_3699);
nand U5008 (N_5008,N_3474,N_3533);
and U5009 (N_5009,N_1751,N_2479);
nor U5010 (N_5010,N_2389,N_401);
or U5011 (N_5011,N_1365,N_287);
and U5012 (N_5012,N_2258,N_3512);
nand U5013 (N_5013,N_2851,N_1150);
nor U5014 (N_5014,N_2755,N_2795);
and U5015 (N_5015,N_2167,N_579);
nor U5016 (N_5016,N_3820,N_413);
nor U5017 (N_5017,N_393,N_3540);
nand U5018 (N_5018,N_366,N_3101);
or U5019 (N_5019,N_600,N_2318);
nand U5020 (N_5020,N_177,N_3062);
or U5021 (N_5021,N_3658,N_497);
or U5022 (N_5022,N_1216,N_3379);
nand U5023 (N_5023,N_1320,N_3933);
nand U5024 (N_5024,N_1655,N_2592);
nand U5025 (N_5025,N_2627,N_1658);
nand U5026 (N_5026,N_3409,N_1766);
and U5027 (N_5027,N_2847,N_1366);
and U5028 (N_5028,N_3507,N_2116);
or U5029 (N_5029,N_400,N_1045);
or U5030 (N_5030,N_1474,N_3701);
and U5031 (N_5031,N_2128,N_164);
or U5032 (N_5032,N_2356,N_2156);
nor U5033 (N_5033,N_3628,N_2652);
nor U5034 (N_5034,N_3674,N_1639);
nand U5035 (N_5035,N_1197,N_3976);
or U5036 (N_5036,N_2064,N_1175);
nand U5037 (N_5037,N_2935,N_1411);
nand U5038 (N_5038,N_2973,N_3765);
nor U5039 (N_5039,N_3382,N_520);
or U5040 (N_5040,N_757,N_3047);
nand U5041 (N_5041,N_3904,N_468);
and U5042 (N_5042,N_3203,N_1319);
nand U5043 (N_5043,N_3097,N_2675);
or U5044 (N_5044,N_3081,N_17);
xnor U5045 (N_5045,N_3289,N_1020);
and U5046 (N_5046,N_2010,N_3934);
xor U5047 (N_5047,N_1959,N_3075);
nand U5048 (N_5048,N_2045,N_1258);
or U5049 (N_5049,N_3275,N_3710);
or U5050 (N_5050,N_2152,N_1664);
and U5051 (N_5051,N_285,N_2564);
nor U5052 (N_5052,N_323,N_1769);
and U5053 (N_5053,N_1237,N_3248);
nor U5054 (N_5054,N_3349,N_1716);
xnor U5055 (N_5055,N_1259,N_649);
nor U5056 (N_5056,N_3610,N_319);
nand U5057 (N_5057,N_1027,N_315);
and U5058 (N_5058,N_1796,N_1098);
or U5059 (N_5059,N_1712,N_1094);
and U5060 (N_5060,N_3280,N_3060);
or U5061 (N_5061,N_1636,N_2719);
nor U5062 (N_5062,N_897,N_865);
and U5063 (N_5063,N_961,N_3745);
or U5064 (N_5064,N_774,N_3394);
or U5065 (N_5065,N_1232,N_3173);
or U5066 (N_5066,N_1269,N_427);
or U5067 (N_5067,N_1285,N_70);
nor U5068 (N_5068,N_1040,N_768);
nand U5069 (N_5069,N_1567,N_1245);
or U5070 (N_5070,N_2724,N_1158);
nand U5071 (N_5071,N_675,N_2353);
and U5072 (N_5072,N_875,N_3667);
nor U5073 (N_5073,N_1344,N_238);
nor U5074 (N_5074,N_1683,N_945);
nor U5075 (N_5075,N_2436,N_15);
nor U5076 (N_5076,N_1436,N_3024);
nor U5077 (N_5077,N_776,N_1375);
and U5078 (N_5078,N_2433,N_893);
nand U5079 (N_5079,N_2296,N_2778);
or U5080 (N_5080,N_1304,N_3604);
or U5081 (N_5081,N_403,N_791);
nand U5082 (N_5082,N_1798,N_952);
or U5083 (N_5083,N_1184,N_2815);
nor U5084 (N_5084,N_2416,N_390);
or U5085 (N_5085,N_708,N_3286);
nand U5086 (N_5086,N_357,N_3764);
nor U5087 (N_5087,N_551,N_737);
and U5088 (N_5088,N_2746,N_345);
nor U5089 (N_5089,N_2539,N_3041);
or U5090 (N_5090,N_3857,N_3215);
nand U5091 (N_5091,N_3999,N_450);
or U5092 (N_5092,N_465,N_2014);
and U5093 (N_5093,N_2381,N_1180);
nor U5094 (N_5094,N_1177,N_1790);
and U5095 (N_5095,N_1310,N_3370);
nor U5096 (N_5096,N_3411,N_638);
nand U5097 (N_5097,N_2394,N_805);
nand U5098 (N_5098,N_431,N_507);
or U5099 (N_5099,N_105,N_692);
nor U5100 (N_5100,N_2723,N_3757);
or U5101 (N_5101,N_3063,N_833);
and U5102 (N_5102,N_1065,N_1554);
or U5103 (N_5103,N_1829,N_2362);
or U5104 (N_5104,N_1609,N_2842);
nand U5105 (N_5105,N_3029,N_3144);
or U5106 (N_5106,N_331,N_3602);
and U5107 (N_5107,N_3902,N_2928);
or U5108 (N_5108,N_878,N_2848);
and U5109 (N_5109,N_173,N_3686);
and U5110 (N_5110,N_651,N_3739);
nand U5111 (N_5111,N_3402,N_3909);
nor U5112 (N_5112,N_3079,N_2805);
and U5113 (N_5113,N_2624,N_204);
nand U5114 (N_5114,N_2044,N_3114);
nor U5115 (N_5115,N_2974,N_3514);
or U5116 (N_5116,N_1801,N_1975);
or U5117 (N_5117,N_444,N_2748);
nor U5118 (N_5118,N_284,N_2535);
nor U5119 (N_5119,N_2632,N_3327);
xor U5120 (N_5120,N_2496,N_2547);
nor U5121 (N_5121,N_728,N_399);
or U5122 (N_5122,N_2635,N_2331);
nand U5123 (N_5123,N_2317,N_2789);
nand U5124 (N_5124,N_508,N_75);
or U5125 (N_5125,N_2868,N_1325);
nand U5126 (N_5126,N_265,N_1113);
or U5127 (N_5127,N_3048,N_2480);
nor U5128 (N_5128,N_1401,N_1271);
or U5129 (N_5129,N_628,N_1463);
and U5130 (N_5130,N_2710,N_3265);
and U5131 (N_5131,N_3878,N_176);
nand U5132 (N_5132,N_2438,N_3802);
xnor U5133 (N_5133,N_1753,N_2173);
or U5134 (N_5134,N_2591,N_3214);
and U5135 (N_5135,N_810,N_2115);
xnor U5136 (N_5136,N_930,N_3321);
and U5137 (N_5137,N_2602,N_3482);
or U5138 (N_5138,N_1836,N_3742);
and U5139 (N_5139,N_1708,N_898);
and U5140 (N_5140,N_2492,N_1793);
nor U5141 (N_5141,N_3919,N_2653);
and U5142 (N_5142,N_1267,N_2067);
nand U5143 (N_5143,N_3709,N_2895);
or U5144 (N_5144,N_1532,N_2163);
nand U5145 (N_5145,N_201,N_104);
or U5146 (N_5146,N_8,N_2032);
and U5147 (N_5147,N_3875,N_499);
or U5148 (N_5148,N_2857,N_1095);
or U5149 (N_5149,N_127,N_3593);
nand U5150 (N_5150,N_3230,N_1653);
or U5151 (N_5151,N_1427,N_3758);
nor U5152 (N_5152,N_263,N_2036);
or U5153 (N_5153,N_855,N_767);
nor U5154 (N_5154,N_1007,N_3619);
nor U5155 (N_5155,N_3361,N_2105);
nand U5156 (N_5156,N_2709,N_340);
nor U5157 (N_5157,N_183,N_2775);
nand U5158 (N_5158,N_3966,N_108);
or U5159 (N_5159,N_3850,N_2327);
or U5160 (N_5160,N_2119,N_1490);
nor U5161 (N_5161,N_2486,N_1997);
nand U5162 (N_5162,N_606,N_531);
or U5163 (N_5163,N_3412,N_2829);
or U5164 (N_5164,N_2562,N_2076);
nor U5165 (N_5165,N_2558,N_306);
and U5166 (N_5166,N_3000,N_3805);
xnor U5167 (N_5167,N_3044,N_367);
nor U5168 (N_5168,N_3620,N_1859);
nand U5169 (N_5169,N_1077,N_717);
or U5170 (N_5170,N_2606,N_3178);
nor U5171 (N_5171,N_3508,N_3351);
nand U5172 (N_5172,N_995,N_169);
nand U5173 (N_5173,N_1581,N_1607);
or U5174 (N_5174,N_1370,N_83);
nand U5175 (N_5175,N_3247,N_3665);
and U5176 (N_5176,N_662,N_3973);
or U5177 (N_5177,N_2628,N_1527);
nand U5178 (N_5178,N_693,N_975);
nand U5179 (N_5179,N_1345,N_2274);
and U5180 (N_5180,N_3362,N_874);
nand U5181 (N_5181,N_877,N_1033);
and U5182 (N_5182,N_1935,N_2534);
nand U5183 (N_5183,N_1438,N_2589);
and U5184 (N_5184,N_3347,N_907);
nor U5185 (N_5185,N_1577,N_2549);
nor U5186 (N_5186,N_1412,N_3918);
nor U5187 (N_5187,N_680,N_3405);
or U5188 (N_5188,N_350,N_3589);
and U5189 (N_5189,N_3343,N_445);
and U5190 (N_5190,N_3561,N_286);
or U5191 (N_5191,N_3867,N_3049);
and U5192 (N_5192,N_724,N_1885);
or U5193 (N_5193,N_439,N_64);
or U5194 (N_5194,N_2975,N_3511);
or U5195 (N_5195,N_2216,N_756);
and U5196 (N_5196,N_1521,N_2901);
nor U5197 (N_5197,N_476,N_2151);
or U5198 (N_5198,N_2615,N_1461);
nand U5199 (N_5199,N_344,N_3907);
or U5200 (N_5200,N_2736,N_333);
and U5201 (N_5201,N_940,N_420);
nor U5202 (N_5202,N_1433,N_2969);
nand U5203 (N_5203,N_3466,N_1840);
or U5204 (N_5204,N_513,N_1545);
nor U5205 (N_5205,N_1833,N_277);
and U5206 (N_5206,N_3256,N_1986);
and U5207 (N_5207,N_1562,N_2874);
or U5208 (N_5208,N_3505,N_2248);
nor U5209 (N_5209,N_1737,N_2888);
or U5210 (N_5210,N_977,N_1186);
nor U5211 (N_5211,N_3893,N_2417);
nor U5212 (N_5212,N_980,N_25);
or U5213 (N_5213,N_3318,N_2507);
nor U5214 (N_5214,N_3253,N_3652);
nor U5215 (N_5215,N_2850,N_1821);
and U5216 (N_5216,N_3251,N_3937);
or U5217 (N_5217,N_3497,N_2209);
nand U5218 (N_5218,N_2841,N_2700);
nor U5219 (N_5219,N_1221,N_1445);
nand U5220 (N_5220,N_161,N_447);
or U5221 (N_5221,N_2900,N_258);
nand U5222 (N_5222,N_560,N_3941);
and U5223 (N_5223,N_185,N_179);
nor U5224 (N_5224,N_716,N_667);
or U5225 (N_5225,N_1055,N_1043);
or U5226 (N_5226,N_2263,N_2970);
and U5227 (N_5227,N_974,N_463);
or U5228 (N_5228,N_1844,N_3557);
or U5229 (N_5229,N_2280,N_3527);
nand U5230 (N_5230,N_1918,N_2567);
nand U5231 (N_5231,N_3359,N_1100);
or U5232 (N_5232,N_2068,N_3278);
and U5233 (N_5233,N_3240,N_2453);
xnor U5234 (N_5234,N_2174,N_218);
nor U5235 (N_5235,N_3345,N_1900);
or U5236 (N_5236,N_1358,N_3414);
nor U5237 (N_5237,N_1872,N_3943);
nand U5238 (N_5238,N_3365,N_2620);
nor U5239 (N_5239,N_1878,N_2955);
nand U5240 (N_5240,N_415,N_1640);
nand U5241 (N_5241,N_1324,N_1908);
and U5242 (N_5242,N_1134,N_3990);
or U5243 (N_5243,N_2626,N_89);
nor U5244 (N_5244,N_1693,N_2141);
nor U5245 (N_5245,N_1651,N_2751);
nor U5246 (N_5246,N_1524,N_1032);
nand U5247 (N_5247,N_3537,N_3813);
nor U5248 (N_5248,N_2078,N_558);
nand U5249 (N_5249,N_2550,N_946);
or U5250 (N_5250,N_2695,N_2002);
or U5251 (N_5251,N_2220,N_1276);
nor U5252 (N_5252,N_2320,N_2979);
and U5253 (N_5253,N_276,N_2691);
nor U5254 (N_5254,N_3105,N_1913);
nand U5255 (N_5255,N_2398,N_3084);
and U5256 (N_5256,N_249,N_1632);
or U5257 (N_5257,N_1133,N_3017);
nor U5258 (N_5258,N_658,N_1066);
nand U5259 (N_5259,N_2527,N_2279);
nand U5260 (N_5260,N_2859,N_136);
nor U5261 (N_5261,N_3072,N_295);
nor U5262 (N_5262,N_2083,N_2972);
and U5263 (N_5263,N_664,N_2987);
or U5264 (N_5264,N_1739,N_3259);
and U5265 (N_5265,N_3218,N_1789);
and U5266 (N_5266,N_3293,N_1464);
or U5267 (N_5267,N_942,N_2614);
and U5268 (N_5268,N_831,N_2771);
and U5269 (N_5269,N_1616,N_3815);
nand U5270 (N_5270,N_1506,N_643);
nand U5271 (N_5271,N_2259,N_2662);
xnor U5272 (N_5272,N_1223,N_746);
and U5273 (N_5273,N_1920,N_2906);
or U5274 (N_5274,N_1565,N_2348);
nand U5275 (N_5275,N_282,N_619);
nor U5276 (N_5276,N_2750,N_3597);
or U5277 (N_5277,N_1700,N_2780);
and U5278 (N_5278,N_47,N_3823);
nor U5279 (N_5279,N_3255,N_1513);
nand U5280 (N_5280,N_609,N_472);
nor U5281 (N_5281,N_1762,N_1072);
and U5282 (N_5282,N_3679,N_402);
nand U5283 (N_5283,N_374,N_455);
nand U5284 (N_5284,N_49,N_451);
nand U5285 (N_5285,N_3614,N_1010);
and U5286 (N_5286,N_1064,N_817);
nor U5287 (N_5287,N_3985,N_3452);
and U5288 (N_5288,N_1726,N_1847);
or U5289 (N_5289,N_3948,N_2390);
and U5290 (N_5290,N_1110,N_145);
or U5291 (N_5291,N_206,N_2450);
nor U5292 (N_5292,N_2271,N_2682);
nor U5293 (N_5293,N_3981,N_1880);
nand U5294 (N_5294,N_1167,N_190);
nand U5295 (N_5295,N_2379,N_3898);
or U5296 (N_5296,N_3429,N_3148);
or U5297 (N_5297,N_1302,N_515);
xor U5298 (N_5298,N_1003,N_1450);
nor U5299 (N_5299,N_3494,N_3363);
and U5300 (N_5300,N_1229,N_825);
xor U5301 (N_5301,N_3404,N_3549);
and U5302 (N_5302,N_2908,N_1071);
and U5303 (N_5303,N_3526,N_317);
and U5304 (N_5304,N_3929,N_1614);
nor U5305 (N_5305,N_129,N_1188);
nor U5306 (N_5306,N_2508,N_130);
nand U5307 (N_5307,N_1794,N_2570);
or U5308 (N_5308,N_1500,N_2745);
nand U5309 (N_5309,N_347,N_2056);
and U5310 (N_5310,N_1299,N_618);
nand U5311 (N_5311,N_3001,N_591);
and U5312 (N_5312,N_1060,N_2656);
nor U5313 (N_5313,N_1512,N_2254);
or U5314 (N_5314,N_2224,N_1934);
nand U5315 (N_5315,N_3928,N_3877);
or U5316 (N_5316,N_352,N_1882);
or U5317 (N_5317,N_1731,N_2893);
nor U5318 (N_5318,N_3868,N_1948);
nand U5319 (N_5319,N_2250,N_3655);
and U5320 (N_5320,N_2495,N_2431);
or U5321 (N_5321,N_2261,N_2283);
or U5322 (N_5322,N_3851,N_3467);
and U5323 (N_5323,N_2865,N_3960);
or U5324 (N_5324,N_1927,N_938);
nor U5325 (N_5325,N_2993,N_960);
and U5326 (N_5326,N_1204,N_1355);
xor U5327 (N_5327,N_151,N_3175);
and U5328 (N_5328,N_876,N_2311);
and U5329 (N_5329,N_3860,N_1209);
and U5330 (N_5330,N_187,N_2809);
and U5331 (N_5331,N_554,N_549);
and U5332 (N_5332,N_1943,N_3677);
nand U5333 (N_5333,N_479,N_665);
nor U5334 (N_5334,N_3982,N_535);
xnor U5335 (N_5335,N_107,N_1947);
or U5336 (N_5336,N_1118,N_1156);
or U5337 (N_5337,N_967,N_3340);
or U5338 (N_5338,N_1587,N_1449);
and U5339 (N_5339,N_2646,N_2699);
nor U5340 (N_5340,N_3638,N_1481);
and U5341 (N_5341,N_2557,N_1619);
and U5342 (N_5342,N_585,N_3284);
and U5343 (N_5343,N_2638,N_1305);
nand U5344 (N_5344,N_3543,N_1035);
and U5345 (N_5345,N_2633,N_280);
or U5346 (N_5346,N_3358,N_1823);
and U5347 (N_5347,N_605,N_807);
nand U5348 (N_5348,N_661,N_3330);
nand U5349 (N_5349,N_1386,N_2047);
nor U5350 (N_5350,N_3468,N_3905);
xor U5351 (N_5351,N_2150,N_1354);
nand U5352 (N_5352,N_2546,N_3951);
nor U5353 (N_5353,N_1713,N_2080);
and U5354 (N_5354,N_813,N_2961);
nor U5355 (N_5355,N_3632,N_3640);
nor U5356 (N_5356,N_365,N_1185);
nand U5357 (N_5357,N_3249,N_559);
nor U5358 (N_5358,N_3799,N_1618);
or U5359 (N_5359,N_885,N_3182);
and U5360 (N_5360,N_1331,N_939);
or U5361 (N_5361,N_135,N_34);
nand U5362 (N_5362,N_1300,N_1759);
nor U5363 (N_5363,N_1023,N_2017);
or U5364 (N_5364,N_3483,N_2035);
or U5365 (N_5365,N_3693,N_3675);
nor U5366 (N_5366,N_191,N_3542);
nand U5367 (N_5367,N_101,N_2837);
and U5368 (N_5368,N_1075,N_3427);
and U5369 (N_5369,N_1670,N_818);
nand U5370 (N_5370,N_2113,N_2806);
nor U5371 (N_5371,N_3587,N_545);
nand U5372 (N_5372,N_3324,N_1582);
or U5373 (N_5373,N_3433,N_2902);
nor U5374 (N_5374,N_2886,N_131);
and U5375 (N_5375,N_1744,N_1479);
and U5376 (N_5376,N_1534,N_991);
and U5377 (N_5377,N_894,N_1569);
or U5378 (N_5378,N_1955,N_3073);
or U5379 (N_5379,N_2720,N_3099);
nor U5380 (N_5380,N_1146,N_2053);
nor U5381 (N_5381,N_3921,N_3339);
nand U5382 (N_5382,N_2188,N_1710);
or U5383 (N_5383,N_2693,N_2545);
nor U5384 (N_5384,N_730,N_1914);
nor U5385 (N_5385,N_1078,N_3232);
nor U5386 (N_5386,N_2333,N_3568);
nor U5387 (N_5387,N_3436,N_55);
and U5388 (N_5388,N_586,N_3357);
nand U5389 (N_5389,N_1548,N_1057);
and U5390 (N_5390,N_1557,N_3100);
or U5391 (N_5391,N_1721,N_1103);
nor U5392 (N_5392,N_3377,N_371);
nor U5393 (N_5393,N_363,N_1764);
or U5394 (N_5394,N_1477,N_3094);
or U5395 (N_5395,N_2149,N_1492);
and U5396 (N_5396,N_1928,N_572);
nand U5397 (N_5397,N_3176,N_3209);
and U5398 (N_5398,N_3663,N_81);
nor U5399 (N_5399,N_3098,N_723);
or U5400 (N_5400,N_1049,N_1625);
or U5401 (N_5401,N_3723,N_43);
nand U5402 (N_5402,N_3292,N_1624);
nand U5403 (N_5403,N_233,N_2642);
and U5404 (N_5404,N_79,N_3273);
and U5405 (N_5405,N_349,N_748);
and U5406 (N_5406,N_3997,N_2443);
or U5407 (N_5407,N_3735,N_1549);
or U5408 (N_5408,N_2821,N_1643);
nor U5409 (N_5409,N_1038,N_1646);
and U5410 (N_5410,N_488,N_3971);
nor U5411 (N_5411,N_1155,N_3220);
nor U5412 (N_5412,N_1215,N_1538);
nor U5413 (N_5413,N_1086,N_1558);
nand U5414 (N_5414,N_3229,N_2399);
nand U5415 (N_5415,N_596,N_1610);
nor U5416 (N_5416,N_896,N_3727);
and U5417 (N_5417,N_3975,N_998);
nor U5418 (N_5418,N_11,N_2233);
or U5419 (N_5419,N_2219,N_117);
nand U5420 (N_5420,N_854,N_3475);
nand U5421 (N_5421,N_1051,N_2172);
nor U5422 (N_5422,N_2286,N_1774);
xor U5423 (N_5423,N_2536,N_732);
or U5424 (N_5424,N_1666,N_1364);
and U5425 (N_5425,N_1073,N_2796);
nor U5426 (N_5426,N_3020,N_452);
xnor U5427 (N_5427,N_443,N_341);
or U5428 (N_5428,N_976,N_1367);
nor U5429 (N_5429,N_2019,N_461);
nand U5430 (N_5430,N_1584,N_2866);
and U5431 (N_5431,N_3091,N_1021);
or U5432 (N_5432,N_3473,N_1692);
nand U5433 (N_5433,N_2252,N_3684);
and U5434 (N_5434,N_290,N_3885);
and U5435 (N_5435,N_195,N_310);
or U5436 (N_5436,N_1922,N_1635);
or U5437 (N_5437,N_2502,N_2658);
nand U5438 (N_5438,N_2957,N_557);
nor U5439 (N_5439,N_2097,N_1520);
and U5440 (N_5440,N_3759,N_3731);
nand U5441 (N_5441,N_2236,N_3430);
nand U5442 (N_5442,N_1274,N_2396);
or U5443 (N_5443,N_904,N_2375);
nor U5444 (N_5444,N_660,N_3279);
or U5445 (N_5445,N_308,N_2284);
nand U5446 (N_5446,N_3682,N_695);
nand U5447 (N_5447,N_3576,N_1294);
or U5448 (N_5448,N_2555,N_2802);
or U5449 (N_5449,N_3171,N_1458);
nor U5450 (N_5450,N_2298,N_655);
xnor U5451 (N_5451,N_3192,N_1318);
nand U5452 (N_5452,N_2171,N_3221);
or U5453 (N_5453,N_3947,N_252);
or U5454 (N_5454,N_3179,N_355);
and U5455 (N_5455,N_1979,N_1369);
or U5456 (N_5456,N_2228,N_1099);
nor U5457 (N_5457,N_2130,N_1089);
and U5458 (N_5458,N_1868,N_2722);
nand U5459 (N_5459,N_3184,N_1575);
and U5460 (N_5460,N_1231,N_3988);
and U5461 (N_5461,N_1656,N_1776);
or U5462 (N_5462,N_3077,N_1253);
nand U5463 (N_5463,N_1834,N_1602);
nand U5464 (N_5464,N_3726,N_3633);
or U5465 (N_5465,N_59,N_3827);
or U5466 (N_5466,N_2916,N_3328);
nor U5467 (N_5467,N_2647,N_546);
or U5468 (N_5468,N_864,N_788);
nand U5469 (N_5469,N_1808,N_2249);
nor U5470 (N_5470,N_3730,N_1854);
and U5471 (N_5471,N_66,N_1243);
nand U5472 (N_5472,N_2997,N_474);
nand U5473 (N_5473,N_3509,N_3970);
or U5474 (N_5474,N_1915,N_2629);
or U5475 (N_5475,N_251,N_160);
xnor U5476 (N_5476,N_908,N_1254);
nor U5477 (N_5477,N_590,N_1016);
nor U5478 (N_5478,N_934,N_172);
or U5479 (N_5479,N_2870,N_1123);
nand U5480 (N_5480,N_2133,N_1757);
nand U5481 (N_5481,N_3371,N_237);
nor U5482 (N_5482,N_1397,N_1668);
nor U5483 (N_5483,N_1404,N_2491);
nor U5484 (N_5484,N_2931,N_2483);
nor U5485 (N_5485,N_1542,N_2146);
nor U5486 (N_5486,N_243,N_1547);
nor U5487 (N_5487,N_3888,N_3565);
and U5488 (N_5488,N_1988,N_2554);
nand U5489 (N_5489,N_514,N_3325);
nor U5490 (N_5490,N_477,N_1553);
and U5491 (N_5491,N_656,N_2315);
nand U5492 (N_5492,N_1780,N_1870);
and U5493 (N_5493,N_3491,N_3071);
and U5494 (N_5494,N_471,N_2292);
and U5495 (N_5495,N_3668,N_354);
nor U5496 (N_5496,N_262,N_3234);
nor U5497 (N_5497,N_906,N_994);
or U5498 (N_5498,N_2737,N_1042);
and U5499 (N_5499,N_3140,N_2946);
and U5500 (N_5500,N_3458,N_460);
or U5501 (N_5501,N_3901,N_1422);
and U5502 (N_5502,N_2707,N_1864);
and U5503 (N_5503,N_1795,N_481);
nor U5504 (N_5504,N_3421,N_1111);
nand U5505 (N_5505,N_2107,N_2196);
or U5506 (N_5506,N_3065,N_3744);
nand U5507 (N_5507,N_3086,N_1597);
nand U5508 (N_5508,N_3027,N_2437);
nand U5509 (N_5509,N_194,N_3798);
and U5510 (N_5510,N_2951,N_2340);
or U5511 (N_5511,N_2201,N_1173);
nand U5512 (N_5512,N_2006,N_1686);
nand U5513 (N_5513,N_1333,N_3598);
or U5514 (N_5514,N_387,N_2089);
or U5515 (N_5515,N_1698,N_2728);
nor U5516 (N_5516,N_1579,N_369);
nand U5517 (N_5517,N_3476,N_1141);
or U5518 (N_5518,N_3037,N_636);
or U5519 (N_5519,N_1138,N_1740);
or U5520 (N_5520,N_862,N_1570);
or U5521 (N_5521,N_1688,N_110);
or U5522 (N_5522,N_617,N_1889);
or U5523 (N_5523,N_2237,N_2556);
nor U5524 (N_5524,N_3516,N_3637);
nor U5525 (N_5525,N_3630,N_2506);
and U5526 (N_5526,N_3720,N_3956);
and U5527 (N_5527,N_3949,N_1178);
or U5528 (N_5528,N_2069,N_2964);
nand U5529 (N_5529,N_111,N_1600);
nor U5530 (N_5530,N_288,N_2959);
and U5531 (N_5531,N_3634,N_895);
or U5532 (N_5532,N_2673,N_654);
nor U5533 (N_5533,N_1973,N_1097);
xor U5534 (N_5534,N_1663,N_2299);
or U5535 (N_5535,N_3870,N_1552);
nand U5536 (N_5536,N_2689,N_3856);
nor U5537 (N_5537,N_1866,N_1140);
nand U5538 (N_5538,N_783,N_3649);
nor U5539 (N_5539,N_599,N_626);
and U5540 (N_5540,N_3089,N_565);
nand U5541 (N_5541,N_2015,N_373);
and U5542 (N_5542,N_2330,N_435);
nor U5543 (N_5543,N_1435,N_1631);
nor U5544 (N_5544,N_2667,N_2306);
nor U5545 (N_5545,N_230,N_2400);
and U5546 (N_5546,N_1391,N_2407);
and U5547 (N_5547,N_3920,N_2609);
and U5548 (N_5548,N_1377,N_3627);
nand U5549 (N_5549,N_763,N_2087);
or U5550 (N_5550,N_2251,N_3563);
nor U5551 (N_5551,N_3187,N_841);
and U5552 (N_5552,N_1342,N_2761);
or U5553 (N_5553,N_1076,N_2355);
nand U5554 (N_5554,N_3767,N_1949);
nor U5555 (N_5555,N_2269,N_3185);
nor U5556 (N_5556,N_1206,N_2867);
or U5557 (N_5557,N_2605,N_1991);
and U5558 (N_5558,N_852,N_2021);
nor U5559 (N_5559,N_562,N_1475);
and U5560 (N_5560,N_255,N_3785);
or U5561 (N_5561,N_3338,N_3031);
and U5562 (N_5562,N_1491,N_3183);
and U5563 (N_5563,N_2424,N_1897);
nor U5564 (N_5564,N_120,N_2377);
and U5565 (N_5565,N_2157,N_1335);
and U5566 (N_5566,N_1473,N_735);
or U5567 (N_5567,N_2845,N_1426);
nand U5568 (N_5568,N_751,N_2285);
and U5569 (N_5569,N_1244,N_3641);
or U5570 (N_5570,N_2909,N_931);
and U5571 (N_5571,N_3892,N_3129);
and U5572 (N_5572,N_2180,N_3418);
and U5573 (N_5573,N_162,N_1969);
nor U5574 (N_5574,N_581,N_3891);
nand U5575 (N_5575,N_1187,N_2);
or U5576 (N_5576,N_928,N_608);
or U5577 (N_5577,N_832,N_293);
or U5578 (N_5578,N_2879,N_241);
and U5579 (N_5579,N_2176,N_2525);
xnor U5580 (N_5580,N_3170,N_2772);
and U5581 (N_5581,N_3132,N_1109);
nor U5582 (N_5582,N_3959,N_2811);
nand U5583 (N_5583,N_1828,N_548);
nor U5584 (N_5584,N_2784,N_27);
nand U5585 (N_5585,N_2965,N_3836);
nor U5586 (N_5586,N_1867,N_3772);
and U5587 (N_5587,N_3128,N_3151);
nor U5588 (N_5588,N_2059,N_149);
and U5589 (N_5589,N_2005,N_182);
and U5590 (N_5590,N_244,N_2137);
nand U5591 (N_5591,N_2966,N_2403);
and U5592 (N_5592,N_576,N_37);
or U5593 (N_5593,N_178,N_2303);
nand U5594 (N_5594,N_261,N_2382);
nand U5595 (N_5595,N_2618,N_988);
or U5596 (N_5596,N_690,N_3761);
nor U5597 (N_5597,N_3711,N_2637);
or U5598 (N_5598,N_2365,N_3329);
and U5599 (N_5599,N_969,N_1544);
nor U5600 (N_5600,N_749,N_1168);
and U5601 (N_5601,N_3126,N_1511);
nand U5602 (N_5602,N_899,N_1916);
or U5603 (N_5603,N_905,N_3716);
nand U5604 (N_5604,N_2071,N_2278);
nor U5605 (N_5605,N_524,N_482);
nor U5606 (N_5606,N_587,N_890);
or U5607 (N_5607,N_2194,N_3914);
nor U5608 (N_5608,N_3978,N_1845);
xor U5609 (N_5609,N_593,N_320);
nand U5610 (N_5610,N_1451,N_3673);
and U5611 (N_5611,N_1903,N_985);
nand U5612 (N_5612,N_3444,N_3992);
and U5613 (N_5613,N_1288,N_3417);
and U5614 (N_5614,N_1611,N_2273);
or U5615 (N_5615,N_3401,N_1210);
and U5616 (N_5616,N_92,N_478);
nor U5617 (N_5617,N_2432,N_2601);
and U5618 (N_5618,N_1806,N_2446);
and U5619 (N_5619,N_48,N_98);
and U5620 (N_5620,N_1453,N_2648);
and U5621 (N_5621,N_335,N_3353);
nor U5622 (N_5622,N_68,N_240);
nor U5623 (N_5623,N_846,N_2788);
xor U5624 (N_5624,N_2308,N_3005);
nand U5625 (N_5625,N_93,N_3825);
xor U5626 (N_5626,N_3775,N_216);
nand U5627 (N_5627,N_1736,N_3307);
nor U5628 (N_5628,N_109,N_2983);
or U5629 (N_5629,N_3415,N_2205);
nor U5630 (N_5630,N_2952,N_3502);
and U5631 (N_5631,N_2938,N_3477);
or U5632 (N_5632,N_2960,N_919);
nor U5633 (N_5633,N_3520,N_1220);
and U5634 (N_5634,N_2739,N_3954);
nand U5635 (N_5635,N_3925,N_3517);
nand U5636 (N_5636,N_997,N_1494);
nor U5637 (N_5637,N_715,N_3407);
or U5638 (N_5638,N_3219,N_1240);
nand U5639 (N_5639,N_1945,N_52);
or U5640 (N_5640,N_2923,N_441);
nor U5641 (N_5641,N_2313,N_3013);
nor U5642 (N_5642,N_3403,N_342);
or U5643 (N_5643,N_3354,N_801);
nand U5644 (N_5644,N_843,N_2227);
and U5645 (N_5645,N_3721,N_1394);
nand U5646 (N_5646,N_1605,N_2833);
or U5647 (N_5647,N_1480,N_3882);
nand U5648 (N_5648,N_2639,N_1219);
nand U5649 (N_5649,N_2852,N_2822);
and U5650 (N_5650,N_3521,N_26);
or U5651 (N_5651,N_2631,N_196);
and U5652 (N_5652,N_1660,N_1588);
nand U5653 (N_5653,N_3572,N_2860);
nand U5654 (N_5654,N_2943,N_2790);
nand U5655 (N_5655,N_3391,N_1717);
and U5656 (N_5656,N_844,N_1595);
and U5657 (N_5657,N_2873,N_1704);
or U5658 (N_5658,N_3080,N_1396);
and U5659 (N_5659,N_1747,N_1937);
nor U5660 (N_5660,N_35,N_3258);
nor U5661 (N_5661,N_921,N_1385);
and U5662 (N_5662,N_3059,N_669);
or U5663 (N_5663,N_987,N_3216);
nand U5664 (N_5664,N_3198,N_1853);
and U5665 (N_5665,N_3158,N_2807);
nand U5666 (N_5666,N_396,N_2426);
and U5667 (N_5667,N_3974,N_762);
and U5668 (N_5668,N_2413,N_1875);
nor U5669 (N_5669,N_1940,N_202);
nor U5670 (N_5670,N_339,N_2468);
or U5671 (N_5671,N_2744,N_2072);
or U5672 (N_5672,N_1931,N_1176);
nand U5673 (N_5673,N_3016,N_1965);
and U5674 (N_5674,N_2222,N_2800);
nand U5675 (N_5675,N_602,N_2947);
nor U5676 (N_5676,N_2371,N_2869);
xor U5677 (N_5677,N_3513,N_2912);
nand U5678 (N_5678,N_598,N_932);
or U5679 (N_5679,N_2942,N_1649);
and U5680 (N_5680,N_725,N_1392);
or U5681 (N_5681,N_1642,N_589);
xnor U5682 (N_5682,N_2329,N_1315);
or U5683 (N_5683,N_1831,N_639);
and U5684 (N_5684,N_3833,N_3442);
and U5685 (N_5685,N_2170,N_3808);
nor U5686 (N_5686,N_3800,N_797);
nor U5687 (N_5687,N_2607,N_2457);
nand U5688 (N_5688,N_3838,N_3083);
nand U5689 (N_5689,N_2221,N_999);
nor U5690 (N_5690,N_2514,N_3522);
or U5691 (N_5691,N_1434,N_2447);
and U5692 (N_5692,N_1779,N_1813);
nor U5693 (N_5693,N_2012,N_1034);
nor U5694 (N_5694,N_2185,N_3146);
and U5695 (N_5695,N_2103,N_1005);
nor U5696 (N_5696,N_2799,N_888);
and U5697 (N_5697,N_3631,N_3866);
or U5698 (N_5698,N_1256,N_2680);
or U5699 (N_5699,N_483,N_3157);
and U5700 (N_5700,N_2937,N_3054);
nand U5701 (N_5701,N_3698,N_1724);
or U5702 (N_5702,N_577,N_944);
nor U5703 (N_5703,N_2337,N_3647);
or U5704 (N_5704,N_753,N_3133);
or U5705 (N_5705,N_3504,N_766);
nand U5706 (N_5706,N_256,N_2109);
nor U5707 (N_5707,N_3687,N_3546);
nand U5708 (N_5708,N_2198,N_2393);
and U5709 (N_5709,N_1295,N_1576);
and U5710 (N_5710,N_2484,N_1887);
nor U5711 (N_5711,N_2363,N_1861);
nor U5712 (N_5712,N_1812,N_3252);
and U5713 (N_5713,N_14,N_2207);
nand U5714 (N_5714,N_2819,N_2364);
or U5715 (N_5715,N_21,N_3880);
or U5716 (N_5716,N_2777,N_3120);
and U5717 (N_5717,N_219,N_41);
and U5718 (N_5718,N_1036,N_924);
and U5719 (N_5719,N_480,N_758);
or U5720 (N_5720,N_1418,N_2057);
nor U5721 (N_5721,N_620,N_2475);
nand U5722 (N_5722,N_2742,N_3366);
or U5723 (N_5723,N_3244,N_1974);
or U5724 (N_5724,N_2255,N_2596);
nand U5725 (N_5725,N_3322,N_1745);
or U5726 (N_5726,N_3858,N_686);
and U5727 (N_5727,N_803,N_869);
nor U5728 (N_5728,N_2472,N_3538);
nor U5729 (N_5729,N_1497,N_2481);
nand U5730 (N_5730,N_2477,N_3567);
or U5731 (N_5731,N_213,N_2238);
and U5732 (N_5732,N_2774,N_209);
nor U5733 (N_5733,N_2808,N_3534);
nand U5734 (N_5734,N_2885,N_2395);
or U5735 (N_5735,N_1714,N_1767);
nor U5736 (N_5736,N_1228,N_3826);
nand U5737 (N_5737,N_2518,N_1987);
xor U5738 (N_5738,N_1626,N_2304);
and U5739 (N_5739,N_2587,N_334);
and U5740 (N_5740,N_2160,N_2967);
nor U5741 (N_5741,N_1912,N_740);
and U5742 (N_5742,N_1608,N_836);
and U5743 (N_5743,N_1406,N_3223);
or U5744 (N_5744,N_1871,N_3816);
and U5745 (N_5745,N_2758,N_812);
and U5746 (N_5746,N_2892,N_436);
and U5747 (N_5747,N_1788,N_2187);
nand U5748 (N_5748,N_1190,N_912);
nor U5749 (N_5749,N_2449,N_2929);
and U5750 (N_5750,N_370,N_1444);
or U5751 (N_5751,N_1041,N_3890);
nand U5752 (N_5752,N_1381,N_3106);
nor U5753 (N_5753,N_2463,N_1301);
nand U5754 (N_5754,N_1154,N_3849);
nor U5755 (N_5755,N_2797,N_1341);
and U5756 (N_5756,N_180,N_2787);
nand U5757 (N_5757,N_3019,N_956);
and U5758 (N_5758,N_1727,N_3766);
and U5759 (N_5759,N_3810,N_2009);
or U5760 (N_5760,N_2439,N_1622);
or U5761 (N_5761,N_722,N_3451);
nor U5762 (N_5762,N_1752,N_2370);
nand U5763 (N_5763,N_3529,N_294);
nand U5764 (N_5764,N_3728,N_2659);
or U5765 (N_5765,N_1613,N_837);
or U5766 (N_5766,N_1092,N_3660);
and U5767 (N_5767,N_850,N_3302);
or U5768 (N_5768,N_3786,N_2590);
or U5769 (N_5769,N_936,N_2517);
xnor U5770 (N_5770,N_1439,N_2988);
or U5771 (N_5771,N_3994,N_3040);
nor U5772 (N_5772,N_3594,N_2962);
nand U5773 (N_5773,N_39,N_1054);
and U5774 (N_5774,N_1359,N_3246);
and U5775 (N_5775,N_281,N_1235);
nor U5776 (N_5776,N_3900,N_500);
and U5777 (N_5777,N_3646,N_3530);
nor U5778 (N_5778,N_1265,N_1541);
nor U5779 (N_5779,N_3161,N_3136);
nor U5780 (N_5780,N_2783,N_2466);
xnor U5781 (N_5781,N_2024,N_2597);
or U5782 (N_5782,N_23,N_2575);
nand U5783 (N_5783,N_671,N_2763);
nor U5784 (N_5784,N_1080,N_1516);
or U5785 (N_5785,N_3926,N_540);
nand U5786 (N_5786,N_2000,N_1519);
or U5787 (N_5787,N_2668,N_3107);
or U5788 (N_5788,N_2240,N_428);
or U5789 (N_5789,N_2663,N_2696);
nand U5790 (N_5790,N_3115,N_2743);
nand U5791 (N_5791,N_3210,N_2835);
and U5792 (N_5792,N_1810,N_2022);
or U5793 (N_5793,N_278,N_2676);
or U5794 (N_5794,N_3344,N_1499);
xor U5795 (N_5795,N_2636,N_2347);
or U5796 (N_5796,N_60,N_3110);
or U5797 (N_5797,N_3191,N_2028);
or U5798 (N_5798,N_3691,N_3499);
nand U5799 (N_5799,N_410,N_2288);
or U5800 (N_5800,N_1827,N_3553);
nor U5801 (N_5801,N_67,N_2831);
and U5802 (N_5802,N_1044,N_611);
nand U5803 (N_5803,N_2664,N_429);
or U5804 (N_5804,N_2785,N_1297);
or U5805 (N_5805,N_3428,N_2544);
nand U5806 (N_5806,N_964,N_1787);
or U5807 (N_5807,N_3806,N_1353);
or U5808 (N_5808,N_10,N_397);
or U5809 (N_5809,N_3360,N_3510);
nor U5810 (N_5810,N_1617,N_154);
nand U5811 (N_5811,N_2734,N_681);
or U5812 (N_5812,N_1326,N_1298);
nor U5813 (N_5813,N_2903,N_1124);
or U5814 (N_5814,N_260,N_30);
nor U5815 (N_5815,N_72,N_1932);
and U5816 (N_5816,N_1090,N_1352);
nor U5817 (N_5817,N_3801,N_2917);
nor U5818 (N_5818,N_1420,N_329);
nand U5819 (N_5819,N_1919,N_653);
nor U5820 (N_5820,N_2430,N_3406);
nand U5821 (N_5821,N_1998,N_830);
nor U5822 (N_5822,N_1467,N_1564);
and U5823 (N_5823,N_3879,N_3199);
nand U5824 (N_5824,N_3859,N_947);
nor U5825 (N_5825,N_3267,N_3957);
nor U5826 (N_5826,N_1347,N_140);
or U5827 (N_5827,N_3281,N_3479);
nand U5828 (N_5828,N_847,N_1884);
and U5829 (N_5829,N_1771,N_1006);
and U5830 (N_5830,N_1208,N_3439);
nand U5831 (N_5831,N_1357,N_2630);
nor U5832 (N_5832,N_3769,N_1349);
nor U5833 (N_5833,N_2191,N_873);
and U5834 (N_5834,N_80,N_3006);
nor U5835 (N_5835,N_3666,N_3519);
or U5836 (N_5836,N_1992,N_272);
nand U5837 (N_5837,N_2574,N_3264);
and U5838 (N_5838,N_1862,N_2003);
nand U5839 (N_5839,N_1440,N_2516);
nor U5840 (N_5840,N_3050,N_422);
nand U5841 (N_5841,N_2013,N_61);
or U5842 (N_5842,N_3469,N_2600);
nor U5843 (N_5843,N_842,N_3755);
nor U5844 (N_5844,N_1425,N_3872);
nor U5845 (N_5845,N_424,N_570);
or U5846 (N_5846,N_2560,N_2451);
nand U5847 (N_5847,N_2754,N_302);
and U5848 (N_5848,N_386,N_2243);
nand U5849 (N_5849,N_2104,N_3374);
nand U5850 (N_5850,N_1029,N_330);
or U5851 (N_5851,N_2683,N_3434);
and U5852 (N_5852,N_3212,N_3443);
nand U5853 (N_5853,N_3303,N_2604);
nor U5854 (N_5854,N_1598,N_3969);
or U5855 (N_5855,N_3531,N_3558);
or U5856 (N_5856,N_3095,N_2990);
nand U5857 (N_5857,N_3348,N_2324);
and U5858 (N_5858,N_2474,N_2568);
and U5859 (N_5859,N_3659,N_3564);
nor U5860 (N_5860,N_902,N_3492);
or U5861 (N_5861,N_1873,N_1194);
nor U5862 (N_5862,N_691,N_392);
nand U5863 (N_5863,N_3605,N_1809);
nand U5864 (N_5864,N_3239,N_2933);
nand U5865 (N_5865,N_6,N_3794);
and U5866 (N_5866,N_1218,N_796);
and U5867 (N_5867,N_3501,N_2681);
xor U5868 (N_5868,N_97,N_1929);
nor U5869 (N_5869,N_563,N_2813);
or U5870 (N_5870,N_1368,N_3090);
or U5871 (N_5871,N_3167,N_3865);
nand U5872 (N_5872,N_2411,N_2677);
nand U5873 (N_5873,N_1144,N_2121);
nor U5874 (N_5874,N_291,N_2321);
or U5875 (N_5875,N_1122,N_432);
nand U5876 (N_5876,N_1526,N_36);
or U5877 (N_5877,N_616,N_1694);
nor U5878 (N_5878,N_2521,N_2175);
nor U5879 (N_5879,N_2027,N_3616);
nand U5880 (N_5880,N_2856,N_2082);
nand U5881 (N_5881,N_3545,N_822);
or U5882 (N_5882,N_1311,N_2428);
or U5883 (N_5883,N_3166,N_3803);
nand U5884 (N_5884,N_205,N_1851);
and U5885 (N_5885,N_3450,N_3681);
nand U5886 (N_5886,N_727,N_1730);
and U5887 (N_5887,N_1212,N_2913);
nor U5888 (N_5888,N_3121,N_296);
xor U5889 (N_5889,N_1938,N_2478);
nor U5890 (N_5890,N_65,N_1546);
nor U5891 (N_5891,N_3582,N_3863);
nor U5892 (N_5892,N_1001,N_3771);
xnor U5893 (N_5893,N_3113,N_2332);
nor U5894 (N_5894,N_3894,N_1951);
or U5895 (N_5895,N_1839,N_1659);
and U5896 (N_5896,N_3035,N_264);
and U5897 (N_5897,N_799,N_1309);
and U5898 (N_5898,N_3924,N_1539);
nor U5899 (N_5899,N_22,N_1957);
or U5900 (N_5900,N_2863,N_2756);
nor U5901 (N_5901,N_358,N_992);
nor U5902 (N_5902,N_1621,N_2812);
nand U5903 (N_5903,N_3601,N_1421);
or U5904 (N_5904,N_2565,N_2117);
nor U5905 (N_5905,N_1356,N_1337);
or U5906 (N_5906,N_3316,N_388);
nand U5907 (N_5907,N_3208,N_2051);
or U5908 (N_5908,N_1507,N_3440);
and U5909 (N_5909,N_3368,N_3272);
or U5910 (N_5910,N_1589,N_2143);
and U5911 (N_5911,N_3972,N_3480);
nor U5912 (N_5912,N_1148,N_3578);
and U5913 (N_5913,N_970,N_561);
or U5914 (N_5914,N_925,N_787);
or U5915 (N_5915,N_3227,N_3676);
and U5916 (N_5916,N_1383,N_115);
nor U5917 (N_5917,N_3991,N_1691);
nor U5918 (N_5918,N_1648,N_3447);
nor U5919 (N_5919,N_679,N_1024);
nor U5920 (N_5920,N_1321,N_2275);
and U5921 (N_5921,N_226,N_3714);
xnor U5922 (N_5922,N_858,N_2958);
nand U5923 (N_5923,N_793,N_1559);
and U5924 (N_5924,N_555,N_1797);
nand U5925 (N_5925,N_1699,N_1313);
and U5926 (N_5926,N_217,N_772);
nor U5927 (N_5927,N_1013,N_467);
and U5928 (N_5928,N_1817,N_1330);
and U5929 (N_5929,N_322,N_2018);
nor U5930 (N_5930,N_1263,N_45);
and U5931 (N_5931,N_1706,N_516);
nor U5932 (N_5932,N_3842,N_2698);
nand U5933 (N_5933,N_307,N_1498);
nor U5934 (N_5934,N_2679,N_983);
and U5935 (N_5935,N_123,N_819);
nor U5936 (N_5936,N_3346,N_2458);
and U5937 (N_5937,N_973,N_1728);
and U5938 (N_5938,N_2202,N_257);
and U5939 (N_5939,N_1750,N_3600);
or U5940 (N_5940,N_1601,N_359);
xor U5941 (N_5941,N_871,N_538);
nand U5942 (N_5942,N_1472,N_3260);
and U5943 (N_5943,N_741,N_1338);
nand U5944 (N_5944,N_650,N_1128);
or U5945 (N_5945,N_166,N_2622);
nor U5946 (N_5946,N_2020,N_3367);
and U5947 (N_5947,N_2341,N_3326);
nand U5948 (N_5948,N_1217,N_3700);
and U5949 (N_5949,N_2644,N_1501);
and U5950 (N_5950,N_2339,N_3984);
nor U5951 (N_5951,N_860,N_978);
nor U5952 (N_5952,N_1634,N_3102);
nand U5953 (N_5953,N_3580,N_2934);
nand U5954 (N_5954,N_220,N_1523);
nor U5955 (N_5955,N_3908,N_3021);
xor U5956 (N_5956,N_2881,N_3410);
nand U5957 (N_5957,N_1283,N_3487);
nor U5958 (N_5958,N_1415,N_3408);
and U5959 (N_5959,N_1022,N_407);
or U5960 (N_5960,N_3980,N_849);
nand U5961 (N_5961,N_3296,N_1630);
nor U5962 (N_5962,N_2485,N_2882);
nor U5963 (N_5963,N_3952,N_1939);
nand U5964 (N_5964,N_714,N_510);
nor U5965 (N_5965,N_948,N_1087);
nor U5966 (N_5966,N_3449,N_2210);
nor U5967 (N_5967,N_1869,N_3225);
nor U5968 (N_5968,N_1841,N_3093);
nor U5969 (N_5969,N_1151,N_3413);
nor U5970 (N_5970,N_2871,N_3525);
nor U5971 (N_5971,N_1734,N_1701);
nor U5972 (N_5972,N_1697,N_3708);
nand U5973 (N_5973,N_523,N_3573);
nor U5974 (N_5974,N_778,N_116);
and U5975 (N_5975,N_3931,N_3352);
and U5976 (N_5976,N_1679,N_1849);
or U5977 (N_5977,N_3911,N_666);
nand U5978 (N_5978,N_3738,N_2725);
and U5979 (N_5979,N_1460,N_3282);
and U5980 (N_5980,N_3989,N_1641);
or U5981 (N_5981,N_32,N_1904);
and U5982 (N_5982,N_2817,N_2526);
nand U5983 (N_5983,N_3463,N_212);
nand U5984 (N_5984,N_775,N_2940);
and U5985 (N_5985,N_1409,N_266);
or U5986 (N_5986,N_3453,N_2383);
nor U5987 (N_5987,N_526,N_3961);
nor U5988 (N_5988,N_689,N_3532);
or U5989 (N_5989,N_2161,N_1671);
or U5990 (N_5990,N_1886,N_2165);
nor U5991 (N_5991,N_3222,N_880);
xnor U5992 (N_5992,N_3334,N_1593);
nor U5993 (N_5993,N_9,N_2731);
or U5994 (N_5994,N_5,N_673);
nor U5995 (N_5995,N_2373,N_3461);
and U5996 (N_5996,N_245,N_684);
or U5997 (N_5997,N_1149,N_2212);
xor U5998 (N_5998,N_1835,N_3523);
nand U5999 (N_5999,N_834,N_95);
nand U6000 (N_6000,N_2757,N_1137);
nor U6001 (N_6001,N_2969,N_3430);
nand U6002 (N_6002,N_1060,N_3065);
nand U6003 (N_6003,N_3629,N_2480);
or U6004 (N_6004,N_3967,N_2364);
or U6005 (N_6005,N_3099,N_3353);
nor U6006 (N_6006,N_3482,N_390);
or U6007 (N_6007,N_31,N_3455);
and U6008 (N_6008,N_3698,N_2266);
nor U6009 (N_6009,N_832,N_251);
or U6010 (N_6010,N_1360,N_1097);
and U6011 (N_6011,N_447,N_200);
or U6012 (N_6012,N_709,N_560);
nand U6013 (N_6013,N_1737,N_1653);
nor U6014 (N_6014,N_3888,N_3279);
nor U6015 (N_6015,N_3759,N_3281);
nand U6016 (N_6016,N_2503,N_2008);
or U6017 (N_6017,N_3021,N_3111);
nand U6018 (N_6018,N_3838,N_2532);
and U6019 (N_6019,N_3106,N_352);
or U6020 (N_6020,N_207,N_1938);
and U6021 (N_6021,N_3869,N_436);
nand U6022 (N_6022,N_2647,N_194);
and U6023 (N_6023,N_2280,N_697);
nand U6024 (N_6024,N_1602,N_1657);
nand U6025 (N_6025,N_2856,N_203);
or U6026 (N_6026,N_1712,N_3240);
or U6027 (N_6027,N_1809,N_2420);
and U6028 (N_6028,N_2739,N_189);
and U6029 (N_6029,N_383,N_2677);
and U6030 (N_6030,N_638,N_3913);
or U6031 (N_6031,N_2698,N_3157);
nand U6032 (N_6032,N_1355,N_8);
nand U6033 (N_6033,N_2239,N_1563);
nor U6034 (N_6034,N_1772,N_3886);
nand U6035 (N_6035,N_3029,N_3431);
nand U6036 (N_6036,N_2712,N_1558);
nor U6037 (N_6037,N_1386,N_276);
or U6038 (N_6038,N_524,N_3702);
nand U6039 (N_6039,N_1170,N_2262);
nand U6040 (N_6040,N_2722,N_3452);
or U6041 (N_6041,N_2014,N_3425);
nor U6042 (N_6042,N_2920,N_3352);
nand U6043 (N_6043,N_1070,N_1816);
nor U6044 (N_6044,N_2466,N_1253);
nor U6045 (N_6045,N_1170,N_1242);
and U6046 (N_6046,N_144,N_2159);
and U6047 (N_6047,N_1749,N_1264);
xor U6048 (N_6048,N_56,N_3754);
nand U6049 (N_6049,N_289,N_1396);
nand U6050 (N_6050,N_19,N_24);
and U6051 (N_6051,N_474,N_3818);
and U6052 (N_6052,N_763,N_354);
nor U6053 (N_6053,N_3671,N_640);
and U6054 (N_6054,N_2250,N_2959);
or U6055 (N_6055,N_3179,N_1887);
nor U6056 (N_6056,N_2157,N_2547);
or U6057 (N_6057,N_2646,N_3692);
nor U6058 (N_6058,N_2552,N_2640);
xnor U6059 (N_6059,N_2119,N_812);
or U6060 (N_6060,N_3356,N_820);
or U6061 (N_6061,N_907,N_2277);
or U6062 (N_6062,N_820,N_2223);
xnor U6063 (N_6063,N_874,N_1927);
nor U6064 (N_6064,N_686,N_3613);
nor U6065 (N_6065,N_3914,N_2475);
and U6066 (N_6066,N_3144,N_3065);
nand U6067 (N_6067,N_2470,N_3747);
and U6068 (N_6068,N_3197,N_1775);
nand U6069 (N_6069,N_1161,N_126);
or U6070 (N_6070,N_3613,N_1107);
and U6071 (N_6071,N_2388,N_692);
and U6072 (N_6072,N_2262,N_2177);
or U6073 (N_6073,N_3117,N_1755);
nand U6074 (N_6074,N_2774,N_591);
and U6075 (N_6075,N_1219,N_2479);
nand U6076 (N_6076,N_3016,N_1229);
nor U6077 (N_6077,N_685,N_2525);
nand U6078 (N_6078,N_2515,N_461);
nor U6079 (N_6079,N_510,N_753);
and U6080 (N_6080,N_3950,N_661);
or U6081 (N_6081,N_479,N_528);
and U6082 (N_6082,N_1488,N_3716);
or U6083 (N_6083,N_36,N_1946);
and U6084 (N_6084,N_2450,N_3658);
and U6085 (N_6085,N_2282,N_3681);
and U6086 (N_6086,N_1630,N_3624);
nor U6087 (N_6087,N_2837,N_1927);
and U6088 (N_6088,N_3139,N_3874);
or U6089 (N_6089,N_2812,N_2061);
nand U6090 (N_6090,N_1829,N_3054);
and U6091 (N_6091,N_368,N_1569);
or U6092 (N_6092,N_1588,N_1838);
and U6093 (N_6093,N_1372,N_3680);
xor U6094 (N_6094,N_2293,N_3200);
and U6095 (N_6095,N_1794,N_730);
and U6096 (N_6096,N_113,N_3760);
or U6097 (N_6097,N_2296,N_598);
nand U6098 (N_6098,N_1275,N_2171);
or U6099 (N_6099,N_1974,N_839);
or U6100 (N_6100,N_819,N_2424);
nor U6101 (N_6101,N_184,N_3907);
nor U6102 (N_6102,N_3332,N_3762);
xnor U6103 (N_6103,N_650,N_1323);
or U6104 (N_6104,N_18,N_3683);
xor U6105 (N_6105,N_2294,N_3998);
nor U6106 (N_6106,N_350,N_2718);
nor U6107 (N_6107,N_908,N_185);
or U6108 (N_6108,N_2713,N_2599);
nor U6109 (N_6109,N_1321,N_3717);
and U6110 (N_6110,N_3400,N_2445);
nor U6111 (N_6111,N_310,N_3299);
nor U6112 (N_6112,N_1821,N_1458);
or U6113 (N_6113,N_1545,N_1775);
nor U6114 (N_6114,N_3714,N_1958);
nor U6115 (N_6115,N_2672,N_2277);
and U6116 (N_6116,N_2376,N_3195);
nand U6117 (N_6117,N_185,N_213);
and U6118 (N_6118,N_1056,N_1536);
nand U6119 (N_6119,N_2421,N_1505);
and U6120 (N_6120,N_1038,N_3477);
nand U6121 (N_6121,N_2040,N_1570);
or U6122 (N_6122,N_3723,N_3404);
and U6123 (N_6123,N_449,N_1743);
nor U6124 (N_6124,N_3747,N_3425);
nand U6125 (N_6125,N_1455,N_1478);
nand U6126 (N_6126,N_3810,N_794);
nor U6127 (N_6127,N_2663,N_450);
and U6128 (N_6128,N_638,N_3227);
nor U6129 (N_6129,N_3153,N_1584);
nand U6130 (N_6130,N_1637,N_3113);
or U6131 (N_6131,N_1232,N_1879);
or U6132 (N_6132,N_1010,N_1865);
nand U6133 (N_6133,N_575,N_1340);
and U6134 (N_6134,N_367,N_3570);
and U6135 (N_6135,N_3789,N_2828);
nor U6136 (N_6136,N_3757,N_2126);
or U6137 (N_6137,N_1357,N_2445);
and U6138 (N_6138,N_1220,N_353);
or U6139 (N_6139,N_1315,N_248);
or U6140 (N_6140,N_3014,N_3882);
nor U6141 (N_6141,N_486,N_39);
nand U6142 (N_6142,N_729,N_484);
xor U6143 (N_6143,N_2842,N_1384);
or U6144 (N_6144,N_1557,N_2454);
nor U6145 (N_6145,N_251,N_1728);
and U6146 (N_6146,N_3401,N_97);
and U6147 (N_6147,N_1577,N_1441);
nor U6148 (N_6148,N_2752,N_1261);
and U6149 (N_6149,N_220,N_615);
nand U6150 (N_6150,N_588,N_1900);
nor U6151 (N_6151,N_2857,N_1787);
nand U6152 (N_6152,N_855,N_1384);
and U6153 (N_6153,N_1701,N_250);
or U6154 (N_6154,N_1798,N_3532);
nand U6155 (N_6155,N_1529,N_2718);
and U6156 (N_6156,N_827,N_3570);
nand U6157 (N_6157,N_3749,N_2454);
or U6158 (N_6158,N_1637,N_1015);
or U6159 (N_6159,N_1293,N_2043);
or U6160 (N_6160,N_2369,N_1675);
or U6161 (N_6161,N_1948,N_2970);
nand U6162 (N_6162,N_93,N_2146);
or U6163 (N_6163,N_2253,N_2287);
and U6164 (N_6164,N_2809,N_3272);
or U6165 (N_6165,N_3756,N_3522);
nand U6166 (N_6166,N_3429,N_1384);
nand U6167 (N_6167,N_241,N_979);
or U6168 (N_6168,N_2347,N_3219);
and U6169 (N_6169,N_2352,N_2692);
or U6170 (N_6170,N_1897,N_2065);
or U6171 (N_6171,N_1366,N_3585);
nand U6172 (N_6172,N_2555,N_1627);
and U6173 (N_6173,N_1554,N_85);
nand U6174 (N_6174,N_1701,N_1272);
and U6175 (N_6175,N_458,N_1981);
and U6176 (N_6176,N_2006,N_3513);
nor U6177 (N_6177,N_974,N_1838);
nor U6178 (N_6178,N_847,N_2114);
or U6179 (N_6179,N_1713,N_1306);
and U6180 (N_6180,N_1236,N_2169);
or U6181 (N_6181,N_594,N_1825);
nor U6182 (N_6182,N_937,N_803);
and U6183 (N_6183,N_2338,N_783);
and U6184 (N_6184,N_2463,N_1844);
and U6185 (N_6185,N_1268,N_3207);
nor U6186 (N_6186,N_427,N_3426);
and U6187 (N_6187,N_1857,N_2474);
nand U6188 (N_6188,N_3305,N_235);
nor U6189 (N_6189,N_710,N_3875);
nand U6190 (N_6190,N_1007,N_3303);
xnor U6191 (N_6191,N_3622,N_3826);
nor U6192 (N_6192,N_3987,N_1983);
and U6193 (N_6193,N_3779,N_1602);
nor U6194 (N_6194,N_3988,N_1157);
nand U6195 (N_6195,N_3690,N_1886);
or U6196 (N_6196,N_2665,N_2617);
or U6197 (N_6197,N_1081,N_2861);
nor U6198 (N_6198,N_2304,N_603);
nor U6199 (N_6199,N_186,N_2972);
nand U6200 (N_6200,N_153,N_2593);
nand U6201 (N_6201,N_190,N_3836);
and U6202 (N_6202,N_3882,N_1987);
and U6203 (N_6203,N_1166,N_88);
nor U6204 (N_6204,N_1047,N_1441);
nor U6205 (N_6205,N_1683,N_2364);
or U6206 (N_6206,N_766,N_392);
nand U6207 (N_6207,N_1767,N_3667);
nor U6208 (N_6208,N_509,N_3124);
and U6209 (N_6209,N_3948,N_549);
and U6210 (N_6210,N_452,N_474);
xnor U6211 (N_6211,N_1007,N_2973);
or U6212 (N_6212,N_1358,N_267);
and U6213 (N_6213,N_3019,N_3462);
xnor U6214 (N_6214,N_2119,N_3528);
or U6215 (N_6215,N_499,N_90);
nand U6216 (N_6216,N_1635,N_1685);
and U6217 (N_6217,N_1906,N_1487);
and U6218 (N_6218,N_232,N_1261);
nor U6219 (N_6219,N_2423,N_1608);
nand U6220 (N_6220,N_397,N_760);
xor U6221 (N_6221,N_1765,N_465);
and U6222 (N_6222,N_1892,N_2913);
and U6223 (N_6223,N_55,N_48);
nand U6224 (N_6224,N_469,N_2686);
nand U6225 (N_6225,N_3025,N_1060);
nor U6226 (N_6226,N_1536,N_3930);
nand U6227 (N_6227,N_57,N_3071);
or U6228 (N_6228,N_277,N_1298);
or U6229 (N_6229,N_2758,N_2599);
or U6230 (N_6230,N_378,N_2772);
or U6231 (N_6231,N_3922,N_2683);
nand U6232 (N_6232,N_1217,N_1602);
or U6233 (N_6233,N_3094,N_258);
nor U6234 (N_6234,N_2809,N_3056);
nor U6235 (N_6235,N_726,N_1013);
nand U6236 (N_6236,N_1760,N_1180);
and U6237 (N_6237,N_1783,N_1603);
nand U6238 (N_6238,N_3724,N_2468);
nand U6239 (N_6239,N_2130,N_2881);
nand U6240 (N_6240,N_1947,N_3187);
nor U6241 (N_6241,N_3388,N_3269);
and U6242 (N_6242,N_1024,N_1759);
and U6243 (N_6243,N_3421,N_2068);
and U6244 (N_6244,N_2334,N_1621);
and U6245 (N_6245,N_3281,N_1389);
nand U6246 (N_6246,N_3426,N_526);
nor U6247 (N_6247,N_1434,N_932);
nor U6248 (N_6248,N_3960,N_3291);
nor U6249 (N_6249,N_809,N_2977);
or U6250 (N_6250,N_2805,N_1162);
nor U6251 (N_6251,N_3870,N_204);
or U6252 (N_6252,N_1273,N_2336);
nor U6253 (N_6253,N_2513,N_2499);
or U6254 (N_6254,N_1631,N_3499);
and U6255 (N_6255,N_3081,N_888);
nand U6256 (N_6256,N_2181,N_3077);
or U6257 (N_6257,N_1910,N_2613);
and U6258 (N_6258,N_1915,N_2094);
nor U6259 (N_6259,N_1177,N_793);
and U6260 (N_6260,N_14,N_2911);
nand U6261 (N_6261,N_3802,N_3925);
and U6262 (N_6262,N_707,N_2831);
nand U6263 (N_6263,N_3721,N_1369);
or U6264 (N_6264,N_3204,N_2938);
or U6265 (N_6265,N_526,N_3199);
nand U6266 (N_6266,N_1750,N_3004);
nand U6267 (N_6267,N_1125,N_1105);
nand U6268 (N_6268,N_3674,N_1776);
nand U6269 (N_6269,N_3128,N_3618);
and U6270 (N_6270,N_2463,N_2582);
and U6271 (N_6271,N_288,N_3626);
and U6272 (N_6272,N_3990,N_1642);
or U6273 (N_6273,N_229,N_524);
or U6274 (N_6274,N_3672,N_2776);
and U6275 (N_6275,N_592,N_1565);
nand U6276 (N_6276,N_1695,N_971);
or U6277 (N_6277,N_1404,N_1707);
or U6278 (N_6278,N_2987,N_3080);
or U6279 (N_6279,N_3578,N_2290);
nand U6280 (N_6280,N_348,N_243);
nor U6281 (N_6281,N_2200,N_1636);
nand U6282 (N_6282,N_3968,N_364);
nor U6283 (N_6283,N_1237,N_1616);
and U6284 (N_6284,N_995,N_3984);
nand U6285 (N_6285,N_3768,N_3800);
and U6286 (N_6286,N_1128,N_3982);
xnor U6287 (N_6287,N_2203,N_2623);
and U6288 (N_6288,N_619,N_3524);
or U6289 (N_6289,N_239,N_3307);
nand U6290 (N_6290,N_402,N_1236);
nand U6291 (N_6291,N_1776,N_3493);
and U6292 (N_6292,N_2422,N_1417);
and U6293 (N_6293,N_1725,N_3130);
nand U6294 (N_6294,N_1017,N_1193);
or U6295 (N_6295,N_2362,N_1837);
nand U6296 (N_6296,N_3675,N_1218);
or U6297 (N_6297,N_2076,N_3473);
or U6298 (N_6298,N_2578,N_1524);
nor U6299 (N_6299,N_1815,N_2053);
and U6300 (N_6300,N_2841,N_851);
nor U6301 (N_6301,N_2895,N_1898);
or U6302 (N_6302,N_311,N_3207);
nor U6303 (N_6303,N_3995,N_1100);
nor U6304 (N_6304,N_148,N_1996);
nand U6305 (N_6305,N_3935,N_1725);
nor U6306 (N_6306,N_2415,N_1784);
nand U6307 (N_6307,N_92,N_2726);
and U6308 (N_6308,N_3289,N_2311);
nand U6309 (N_6309,N_2454,N_1073);
nand U6310 (N_6310,N_2805,N_3254);
nor U6311 (N_6311,N_3902,N_3838);
or U6312 (N_6312,N_2566,N_1508);
nor U6313 (N_6313,N_1449,N_389);
nand U6314 (N_6314,N_1387,N_2269);
nor U6315 (N_6315,N_309,N_1602);
nor U6316 (N_6316,N_277,N_699);
or U6317 (N_6317,N_3092,N_60);
and U6318 (N_6318,N_1346,N_1360);
and U6319 (N_6319,N_106,N_3514);
nor U6320 (N_6320,N_1641,N_3723);
and U6321 (N_6321,N_508,N_3566);
or U6322 (N_6322,N_2847,N_675);
or U6323 (N_6323,N_2065,N_1613);
and U6324 (N_6324,N_1724,N_1151);
and U6325 (N_6325,N_2967,N_3135);
nor U6326 (N_6326,N_3245,N_626);
and U6327 (N_6327,N_2708,N_126);
nor U6328 (N_6328,N_3319,N_3720);
and U6329 (N_6329,N_933,N_2240);
or U6330 (N_6330,N_1792,N_2132);
nand U6331 (N_6331,N_1851,N_129);
and U6332 (N_6332,N_3902,N_1843);
nor U6333 (N_6333,N_2727,N_1647);
or U6334 (N_6334,N_860,N_1198);
and U6335 (N_6335,N_146,N_610);
nor U6336 (N_6336,N_3867,N_1553);
nand U6337 (N_6337,N_2007,N_523);
and U6338 (N_6338,N_1047,N_1992);
or U6339 (N_6339,N_1050,N_3219);
nand U6340 (N_6340,N_1087,N_252);
or U6341 (N_6341,N_135,N_3257);
or U6342 (N_6342,N_2300,N_309);
or U6343 (N_6343,N_2262,N_3545);
xnor U6344 (N_6344,N_2746,N_2714);
nand U6345 (N_6345,N_2088,N_298);
nand U6346 (N_6346,N_2168,N_653);
nor U6347 (N_6347,N_1771,N_1309);
nand U6348 (N_6348,N_3936,N_3770);
nand U6349 (N_6349,N_247,N_848);
or U6350 (N_6350,N_319,N_2464);
nand U6351 (N_6351,N_2999,N_3871);
and U6352 (N_6352,N_3301,N_1266);
or U6353 (N_6353,N_350,N_2445);
nand U6354 (N_6354,N_1091,N_3604);
and U6355 (N_6355,N_2017,N_1808);
nand U6356 (N_6356,N_858,N_1002);
nor U6357 (N_6357,N_3034,N_1705);
and U6358 (N_6358,N_1550,N_1597);
nor U6359 (N_6359,N_99,N_1584);
nor U6360 (N_6360,N_401,N_1283);
and U6361 (N_6361,N_969,N_787);
or U6362 (N_6362,N_2800,N_508);
and U6363 (N_6363,N_1737,N_290);
nor U6364 (N_6364,N_2500,N_1015);
or U6365 (N_6365,N_2940,N_779);
and U6366 (N_6366,N_73,N_2760);
nand U6367 (N_6367,N_2569,N_3712);
nor U6368 (N_6368,N_675,N_792);
nor U6369 (N_6369,N_1439,N_1705);
or U6370 (N_6370,N_1000,N_667);
and U6371 (N_6371,N_881,N_1569);
nor U6372 (N_6372,N_930,N_2072);
or U6373 (N_6373,N_3169,N_3932);
nand U6374 (N_6374,N_3662,N_1970);
and U6375 (N_6375,N_2881,N_1216);
or U6376 (N_6376,N_1875,N_1765);
xnor U6377 (N_6377,N_3431,N_2995);
nand U6378 (N_6378,N_3205,N_848);
and U6379 (N_6379,N_564,N_1983);
nor U6380 (N_6380,N_3867,N_1169);
xnor U6381 (N_6381,N_1540,N_3242);
nor U6382 (N_6382,N_1533,N_2586);
or U6383 (N_6383,N_3551,N_2926);
and U6384 (N_6384,N_3652,N_1909);
and U6385 (N_6385,N_3445,N_760);
nand U6386 (N_6386,N_3870,N_3370);
nand U6387 (N_6387,N_2900,N_1031);
or U6388 (N_6388,N_1705,N_2335);
nand U6389 (N_6389,N_814,N_3345);
or U6390 (N_6390,N_2260,N_1532);
or U6391 (N_6391,N_2499,N_696);
nor U6392 (N_6392,N_790,N_1227);
nand U6393 (N_6393,N_3732,N_3340);
and U6394 (N_6394,N_3734,N_456);
nand U6395 (N_6395,N_3896,N_3235);
nor U6396 (N_6396,N_216,N_884);
nand U6397 (N_6397,N_3994,N_3606);
nor U6398 (N_6398,N_3151,N_3929);
nor U6399 (N_6399,N_829,N_1458);
nor U6400 (N_6400,N_27,N_739);
and U6401 (N_6401,N_3224,N_1903);
and U6402 (N_6402,N_3699,N_2739);
and U6403 (N_6403,N_1799,N_2976);
nand U6404 (N_6404,N_3857,N_1153);
and U6405 (N_6405,N_3368,N_3101);
nand U6406 (N_6406,N_2652,N_2463);
xor U6407 (N_6407,N_2478,N_967);
or U6408 (N_6408,N_363,N_2509);
nor U6409 (N_6409,N_1637,N_2518);
nor U6410 (N_6410,N_1246,N_2284);
or U6411 (N_6411,N_2276,N_3487);
and U6412 (N_6412,N_783,N_2717);
xor U6413 (N_6413,N_1339,N_53);
nor U6414 (N_6414,N_2723,N_253);
nand U6415 (N_6415,N_3570,N_431);
nor U6416 (N_6416,N_1740,N_2530);
nor U6417 (N_6417,N_3215,N_1717);
and U6418 (N_6418,N_3379,N_1770);
nor U6419 (N_6419,N_2692,N_1500);
or U6420 (N_6420,N_2348,N_884);
nand U6421 (N_6421,N_23,N_2727);
nor U6422 (N_6422,N_1853,N_2089);
nor U6423 (N_6423,N_2892,N_2695);
nor U6424 (N_6424,N_3389,N_1135);
nand U6425 (N_6425,N_2898,N_746);
nor U6426 (N_6426,N_1223,N_13);
or U6427 (N_6427,N_1302,N_280);
or U6428 (N_6428,N_1739,N_479);
and U6429 (N_6429,N_742,N_1617);
and U6430 (N_6430,N_1731,N_524);
nand U6431 (N_6431,N_3779,N_3660);
nor U6432 (N_6432,N_1274,N_3860);
and U6433 (N_6433,N_335,N_2556);
nand U6434 (N_6434,N_1543,N_2201);
and U6435 (N_6435,N_2124,N_2014);
and U6436 (N_6436,N_160,N_555);
or U6437 (N_6437,N_2051,N_2950);
or U6438 (N_6438,N_3922,N_2756);
xor U6439 (N_6439,N_3574,N_2523);
nor U6440 (N_6440,N_1562,N_393);
or U6441 (N_6441,N_2701,N_86);
xnor U6442 (N_6442,N_2370,N_1253);
and U6443 (N_6443,N_3663,N_1915);
or U6444 (N_6444,N_1536,N_2889);
and U6445 (N_6445,N_1458,N_658);
nor U6446 (N_6446,N_1909,N_7);
nor U6447 (N_6447,N_3229,N_3827);
and U6448 (N_6448,N_3456,N_3495);
or U6449 (N_6449,N_91,N_3064);
nand U6450 (N_6450,N_2100,N_481);
or U6451 (N_6451,N_1855,N_369);
nand U6452 (N_6452,N_1060,N_2398);
and U6453 (N_6453,N_2029,N_488);
nor U6454 (N_6454,N_3286,N_3688);
and U6455 (N_6455,N_2176,N_533);
and U6456 (N_6456,N_2168,N_574);
or U6457 (N_6457,N_2555,N_2750);
or U6458 (N_6458,N_2864,N_3272);
nor U6459 (N_6459,N_337,N_2724);
nor U6460 (N_6460,N_828,N_2899);
nor U6461 (N_6461,N_3636,N_3008);
and U6462 (N_6462,N_3412,N_1875);
nand U6463 (N_6463,N_627,N_2502);
and U6464 (N_6464,N_790,N_3242);
nor U6465 (N_6465,N_1671,N_1906);
and U6466 (N_6466,N_283,N_1006);
or U6467 (N_6467,N_2223,N_314);
nand U6468 (N_6468,N_3524,N_3673);
nand U6469 (N_6469,N_197,N_3857);
or U6470 (N_6470,N_18,N_3845);
or U6471 (N_6471,N_2677,N_3103);
or U6472 (N_6472,N_779,N_2900);
nor U6473 (N_6473,N_3455,N_1264);
nand U6474 (N_6474,N_911,N_2776);
or U6475 (N_6475,N_2966,N_3222);
nor U6476 (N_6476,N_936,N_635);
nand U6477 (N_6477,N_3350,N_3141);
or U6478 (N_6478,N_3899,N_2920);
nor U6479 (N_6479,N_977,N_877);
nand U6480 (N_6480,N_2050,N_2710);
nand U6481 (N_6481,N_812,N_988);
nand U6482 (N_6482,N_1143,N_576);
nor U6483 (N_6483,N_2141,N_1831);
and U6484 (N_6484,N_2563,N_3198);
and U6485 (N_6485,N_2992,N_3430);
nor U6486 (N_6486,N_1668,N_2132);
nand U6487 (N_6487,N_1838,N_3284);
nand U6488 (N_6488,N_3514,N_1547);
nand U6489 (N_6489,N_1850,N_855);
and U6490 (N_6490,N_3913,N_3453);
nand U6491 (N_6491,N_1226,N_2298);
and U6492 (N_6492,N_902,N_253);
xnor U6493 (N_6493,N_2374,N_707);
nand U6494 (N_6494,N_2377,N_3301);
nand U6495 (N_6495,N_2380,N_3367);
and U6496 (N_6496,N_3426,N_1491);
nor U6497 (N_6497,N_526,N_3632);
nand U6498 (N_6498,N_2411,N_2605);
or U6499 (N_6499,N_1917,N_1235);
nand U6500 (N_6500,N_1918,N_843);
and U6501 (N_6501,N_3494,N_347);
nor U6502 (N_6502,N_825,N_2149);
or U6503 (N_6503,N_775,N_2271);
or U6504 (N_6504,N_3142,N_3744);
nor U6505 (N_6505,N_361,N_116);
nor U6506 (N_6506,N_3816,N_1114);
nand U6507 (N_6507,N_1020,N_2517);
or U6508 (N_6508,N_3649,N_1603);
nor U6509 (N_6509,N_1163,N_447);
nand U6510 (N_6510,N_76,N_1855);
or U6511 (N_6511,N_828,N_3763);
and U6512 (N_6512,N_3186,N_2856);
and U6513 (N_6513,N_1052,N_1825);
nor U6514 (N_6514,N_2189,N_468);
nand U6515 (N_6515,N_3789,N_3107);
or U6516 (N_6516,N_1531,N_2669);
or U6517 (N_6517,N_2197,N_1972);
nor U6518 (N_6518,N_848,N_35);
and U6519 (N_6519,N_943,N_851);
and U6520 (N_6520,N_643,N_3735);
nand U6521 (N_6521,N_335,N_2106);
and U6522 (N_6522,N_898,N_357);
nand U6523 (N_6523,N_269,N_426);
and U6524 (N_6524,N_2552,N_60);
nand U6525 (N_6525,N_269,N_2512);
nand U6526 (N_6526,N_1226,N_1943);
and U6527 (N_6527,N_3942,N_3448);
and U6528 (N_6528,N_1010,N_2767);
nand U6529 (N_6529,N_938,N_3706);
or U6530 (N_6530,N_1657,N_11);
nor U6531 (N_6531,N_2156,N_3808);
nand U6532 (N_6532,N_3544,N_3509);
and U6533 (N_6533,N_1909,N_1208);
nor U6534 (N_6534,N_3436,N_2976);
or U6535 (N_6535,N_3852,N_2731);
nor U6536 (N_6536,N_2508,N_3845);
nand U6537 (N_6537,N_1216,N_2047);
or U6538 (N_6538,N_3926,N_721);
nand U6539 (N_6539,N_3077,N_3091);
nor U6540 (N_6540,N_2616,N_821);
nand U6541 (N_6541,N_1106,N_3140);
nand U6542 (N_6542,N_1524,N_2470);
and U6543 (N_6543,N_799,N_2630);
nand U6544 (N_6544,N_933,N_2353);
nand U6545 (N_6545,N_1890,N_89);
and U6546 (N_6546,N_2730,N_3737);
nor U6547 (N_6547,N_3526,N_3391);
or U6548 (N_6548,N_2428,N_324);
and U6549 (N_6549,N_3766,N_2053);
and U6550 (N_6550,N_1477,N_1320);
and U6551 (N_6551,N_300,N_998);
and U6552 (N_6552,N_1159,N_803);
nand U6553 (N_6553,N_2826,N_2903);
and U6554 (N_6554,N_2540,N_3577);
and U6555 (N_6555,N_3289,N_2768);
or U6556 (N_6556,N_3799,N_30);
and U6557 (N_6557,N_3681,N_1802);
and U6558 (N_6558,N_3284,N_3268);
nor U6559 (N_6559,N_615,N_872);
nor U6560 (N_6560,N_628,N_435);
nand U6561 (N_6561,N_3741,N_2232);
nand U6562 (N_6562,N_3305,N_317);
nand U6563 (N_6563,N_3995,N_3733);
or U6564 (N_6564,N_2918,N_883);
xor U6565 (N_6565,N_468,N_3504);
and U6566 (N_6566,N_1929,N_3477);
or U6567 (N_6567,N_2524,N_1377);
and U6568 (N_6568,N_1000,N_3529);
nor U6569 (N_6569,N_1316,N_850);
or U6570 (N_6570,N_3345,N_2495);
and U6571 (N_6571,N_1841,N_144);
or U6572 (N_6572,N_3806,N_2342);
or U6573 (N_6573,N_1277,N_2201);
or U6574 (N_6574,N_1421,N_1497);
nand U6575 (N_6575,N_2349,N_428);
or U6576 (N_6576,N_3522,N_3142);
nand U6577 (N_6577,N_224,N_3911);
or U6578 (N_6578,N_2066,N_2777);
or U6579 (N_6579,N_2624,N_3034);
and U6580 (N_6580,N_3715,N_1252);
or U6581 (N_6581,N_3238,N_2647);
or U6582 (N_6582,N_3058,N_1536);
nand U6583 (N_6583,N_1523,N_2362);
or U6584 (N_6584,N_1566,N_779);
or U6585 (N_6585,N_3783,N_2066);
xnor U6586 (N_6586,N_1309,N_3096);
and U6587 (N_6587,N_3967,N_792);
nor U6588 (N_6588,N_3807,N_2165);
nand U6589 (N_6589,N_488,N_616);
nor U6590 (N_6590,N_1856,N_268);
nand U6591 (N_6591,N_2539,N_1624);
and U6592 (N_6592,N_2465,N_1973);
nand U6593 (N_6593,N_2785,N_3826);
or U6594 (N_6594,N_1766,N_3725);
nand U6595 (N_6595,N_1478,N_3157);
xor U6596 (N_6596,N_2724,N_481);
nand U6597 (N_6597,N_215,N_961);
and U6598 (N_6598,N_928,N_284);
and U6599 (N_6599,N_2126,N_1211);
nor U6600 (N_6600,N_697,N_1686);
and U6601 (N_6601,N_508,N_1646);
or U6602 (N_6602,N_3726,N_180);
nand U6603 (N_6603,N_1403,N_1058);
or U6604 (N_6604,N_1333,N_2774);
nor U6605 (N_6605,N_3973,N_3896);
or U6606 (N_6606,N_1624,N_1644);
and U6607 (N_6607,N_283,N_2252);
nor U6608 (N_6608,N_1971,N_1694);
or U6609 (N_6609,N_819,N_3280);
xnor U6610 (N_6610,N_3871,N_1497);
or U6611 (N_6611,N_87,N_186);
nor U6612 (N_6612,N_3827,N_893);
nand U6613 (N_6613,N_119,N_3203);
nor U6614 (N_6614,N_3916,N_2163);
nor U6615 (N_6615,N_2697,N_2819);
nor U6616 (N_6616,N_2505,N_1571);
and U6617 (N_6617,N_2759,N_1183);
nor U6618 (N_6618,N_942,N_174);
nand U6619 (N_6619,N_2977,N_931);
or U6620 (N_6620,N_2317,N_2615);
nand U6621 (N_6621,N_1326,N_1834);
and U6622 (N_6622,N_901,N_1838);
and U6623 (N_6623,N_833,N_2359);
nand U6624 (N_6624,N_3475,N_1119);
nor U6625 (N_6625,N_3848,N_1128);
or U6626 (N_6626,N_1097,N_2992);
nand U6627 (N_6627,N_1997,N_1819);
or U6628 (N_6628,N_3792,N_590);
nand U6629 (N_6629,N_1975,N_3332);
and U6630 (N_6630,N_1482,N_3091);
or U6631 (N_6631,N_2842,N_3898);
nor U6632 (N_6632,N_432,N_3640);
nor U6633 (N_6633,N_2701,N_1663);
nand U6634 (N_6634,N_3091,N_2048);
nand U6635 (N_6635,N_2480,N_63);
and U6636 (N_6636,N_3718,N_2106);
nor U6637 (N_6637,N_1518,N_315);
and U6638 (N_6638,N_1475,N_2061);
nand U6639 (N_6639,N_108,N_705);
and U6640 (N_6640,N_1842,N_3717);
nor U6641 (N_6641,N_2436,N_2898);
nor U6642 (N_6642,N_3191,N_3938);
nor U6643 (N_6643,N_2123,N_2904);
or U6644 (N_6644,N_2987,N_2502);
nand U6645 (N_6645,N_2363,N_3458);
nand U6646 (N_6646,N_738,N_2106);
and U6647 (N_6647,N_874,N_264);
and U6648 (N_6648,N_309,N_2229);
nor U6649 (N_6649,N_1823,N_891);
and U6650 (N_6650,N_2936,N_3609);
and U6651 (N_6651,N_3968,N_2283);
or U6652 (N_6652,N_2213,N_3607);
or U6653 (N_6653,N_3680,N_747);
or U6654 (N_6654,N_92,N_2342);
nor U6655 (N_6655,N_510,N_2342);
and U6656 (N_6656,N_782,N_253);
nor U6657 (N_6657,N_2090,N_3595);
or U6658 (N_6658,N_1081,N_892);
and U6659 (N_6659,N_3843,N_1325);
nand U6660 (N_6660,N_2310,N_903);
and U6661 (N_6661,N_2066,N_225);
nor U6662 (N_6662,N_1945,N_819);
or U6663 (N_6663,N_751,N_3213);
nor U6664 (N_6664,N_3057,N_3385);
nor U6665 (N_6665,N_3682,N_3936);
nand U6666 (N_6666,N_1223,N_1731);
nand U6667 (N_6667,N_1256,N_3784);
nor U6668 (N_6668,N_444,N_289);
nand U6669 (N_6669,N_969,N_1700);
or U6670 (N_6670,N_3784,N_2534);
and U6671 (N_6671,N_154,N_3260);
nor U6672 (N_6672,N_1004,N_3993);
nor U6673 (N_6673,N_3685,N_300);
nor U6674 (N_6674,N_3176,N_1583);
nor U6675 (N_6675,N_3479,N_1321);
nor U6676 (N_6676,N_3410,N_3151);
nand U6677 (N_6677,N_3899,N_2605);
nand U6678 (N_6678,N_3894,N_1113);
and U6679 (N_6679,N_178,N_3906);
nor U6680 (N_6680,N_3963,N_1841);
and U6681 (N_6681,N_3161,N_3297);
nor U6682 (N_6682,N_137,N_3172);
or U6683 (N_6683,N_2879,N_3990);
and U6684 (N_6684,N_1621,N_2984);
or U6685 (N_6685,N_3177,N_2823);
nand U6686 (N_6686,N_2162,N_2518);
nor U6687 (N_6687,N_3631,N_1061);
nor U6688 (N_6688,N_2304,N_1123);
or U6689 (N_6689,N_1406,N_642);
or U6690 (N_6690,N_937,N_2643);
or U6691 (N_6691,N_1349,N_2214);
or U6692 (N_6692,N_628,N_2598);
and U6693 (N_6693,N_2519,N_2741);
and U6694 (N_6694,N_3206,N_2062);
nor U6695 (N_6695,N_1341,N_1164);
or U6696 (N_6696,N_2783,N_3203);
nand U6697 (N_6697,N_1808,N_1910);
or U6698 (N_6698,N_3298,N_3157);
and U6699 (N_6699,N_262,N_3218);
nor U6700 (N_6700,N_1329,N_2772);
nor U6701 (N_6701,N_3992,N_2859);
or U6702 (N_6702,N_1833,N_1965);
nor U6703 (N_6703,N_105,N_2624);
nor U6704 (N_6704,N_1862,N_2266);
nor U6705 (N_6705,N_609,N_3380);
or U6706 (N_6706,N_2715,N_2585);
or U6707 (N_6707,N_2178,N_3764);
or U6708 (N_6708,N_599,N_2691);
and U6709 (N_6709,N_1920,N_509);
nor U6710 (N_6710,N_603,N_3971);
nand U6711 (N_6711,N_1951,N_2589);
and U6712 (N_6712,N_991,N_2206);
or U6713 (N_6713,N_594,N_749);
nand U6714 (N_6714,N_768,N_1946);
and U6715 (N_6715,N_1973,N_358);
nand U6716 (N_6716,N_434,N_3493);
nand U6717 (N_6717,N_3908,N_280);
or U6718 (N_6718,N_3624,N_608);
and U6719 (N_6719,N_1864,N_1898);
nor U6720 (N_6720,N_3954,N_3883);
nand U6721 (N_6721,N_3388,N_734);
and U6722 (N_6722,N_1142,N_3311);
or U6723 (N_6723,N_3184,N_784);
nor U6724 (N_6724,N_1048,N_3699);
nor U6725 (N_6725,N_2951,N_3667);
and U6726 (N_6726,N_880,N_1678);
or U6727 (N_6727,N_3951,N_3161);
or U6728 (N_6728,N_2984,N_175);
nor U6729 (N_6729,N_3969,N_3877);
nand U6730 (N_6730,N_3379,N_3866);
nand U6731 (N_6731,N_849,N_2486);
or U6732 (N_6732,N_2354,N_842);
nor U6733 (N_6733,N_1011,N_1094);
nor U6734 (N_6734,N_2011,N_2162);
nand U6735 (N_6735,N_2449,N_310);
nand U6736 (N_6736,N_2787,N_1869);
or U6737 (N_6737,N_3143,N_157);
nor U6738 (N_6738,N_1109,N_929);
and U6739 (N_6739,N_1842,N_451);
nand U6740 (N_6740,N_3839,N_540);
nor U6741 (N_6741,N_3088,N_2884);
nand U6742 (N_6742,N_2602,N_237);
nor U6743 (N_6743,N_2748,N_1451);
and U6744 (N_6744,N_1687,N_3373);
or U6745 (N_6745,N_3368,N_442);
and U6746 (N_6746,N_944,N_2300);
nor U6747 (N_6747,N_2602,N_3732);
nor U6748 (N_6748,N_1141,N_283);
nand U6749 (N_6749,N_1923,N_414);
nor U6750 (N_6750,N_128,N_533);
nand U6751 (N_6751,N_3238,N_886);
nand U6752 (N_6752,N_3538,N_1333);
or U6753 (N_6753,N_742,N_1013);
nand U6754 (N_6754,N_1160,N_3281);
nor U6755 (N_6755,N_678,N_1608);
or U6756 (N_6756,N_3464,N_2349);
nor U6757 (N_6757,N_2411,N_2008);
nand U6758 (N_6758,N_1661,N_3326);
nor U6759 (N_6759,N_2996,N_1948);
nor U6760 (N_6760,N_993,N_424);
or U6761 (N_6761,N_2303,N_5);
nor U6762 (N_6762,N_1521,N_670);
and U6763 (N_6763,N_3816,N_3949);
or U6764 (N_6764,N_88,N_1308);
and U6765 (N_6765,N_662,N_1447);
nand U6766 (N_6766,N_2506,N_1598);
nand U6767 (N_6767,N_1740,N_3247);
nor U6768 (N_6768,N_2477,N_3338);
or U6769 (N_6769,N_2742,N_493);
or U6770 (N_6770,N_1622,N_2611);
and U6771 (N_6771,N_2853,N_3775);
or U6772 (N_6772,N_646,N_2419);
and U6773 (N_6773,N_2206,N_121);
and U6774 (N_6774,N_1718,N_2418);
and U6775 (N_6775,N_1364,N_643);
nor U6776 (N_6776,N_1652,N_1239);
nand U6777 (N_6777,N_2276,N_1952);
nand U6778 (N_6778,N_3518,N_3281);
nand U6779 (N_6779,N_2058,N_489);
nor U6780 (N_6780,N_2375,N_3273);
and U6781 (N_6781,N_1638,N_750);
nand U6782 (N_6782,N_2494,N_1886);
nor U6783 (N_6783,N_3792,N_3103);
nand U6784 (N_6784,N_2455,N_2593);
xnor U6785 (N_6785,N_2929,N_3509);
or U6786 (N_6786,N_1026,N_2323);
nand U6787 (N_6787,N_3759,N_82);
nor U6788 (N_6788,N_2749,N_2274);
or U6789 (N_6789,N_349,N_1691);
nor U6790 (N_6790,N_1667,N_435);
or U6791 (N_6791,N_1718,N_3891);
or U6792 (N_6792,N_801,N_1336);
or U6793 (N_6793,N_885,N_1205);
or U6794 (N_6794,N_793,N_3243);
nor U6795 (N_6795,N_1156,N_762);
nor U6796 (N_6796,N_3198,N_551);
nor U6797 (N_6797,N_1156,N_727);
and U6798 (N_6798,N_2979,N_1340);
nand U6799 (N_6799,N_2606,N_210);
and U6800 (N_6800,N_1855,N_2321);
or U6801 (N_6801,N_2634,N_1508);
nor U6802 (N_6802,N_2797,N_952);
nor U6803 (N_6803,N_2163,N_3295);
and U6804 (N_6804,N_1073,N_1889);
and U6805 (N_6805,N_558,N_568);
nor U6806 (N_6806,N_2588,N_1680);
nand U6807 (N_6807,N_3651,N_3066);
nand U6808 (N_6808,N_1179,N_1465);
xnor U6809 (N_6809,N_2886,N_43);
or U6810 (N_6810,N_3783,N_1048);
nor U6811 (N_6811,N_3288,N_1402);
nor U6812 (N_6812,N_2332,N_358);
nand U6813 (N_6813,N_2765,N_55);
nor U6814 (N_6814,N_3601,N_1311);
nand U6815 (N_6815,N_361,N_3896);
nor U6816 (N_6816,N_3466,N_3331);
nor U6817 (N_6817,N_3087,N_2878);
nor U6818 (N_6818,N_3870,N_860);
and U6819 (N_6819,N_1635,N_2966);
nor U6820 (N_6820,N_1681,N_466);
and U6821 (N_6821,N_3754,N_2056);
nor U6822 (N_6822,N_412,N_3218);
or U6823 (N_6823,N_1618,N_3386);
and U6824 (N_6824,N_3958,N_806);
nand U6825 (N_6825,N_1293,N_2179);
or U6826 (N_6826,N_200,N_3248);
nand U6827 (N_6827,N_1774,N_3413);
or U6828 (N_6828,N_331,N_3511);
or U6829 (N_6829,N_1096,N_1102);
nand U6830 (N_6830,N_3189,N_2279);
or U6831 (N_6831,N_1044,N_3427);
and U6832 (N_6832,N_2616,N_721);
nand U6833 (N_6833,N_3664,N_2414);
and U6834 (N_6834,N_2778,N_2255);
nor U6835 (N_6835,N_2430,N_2358);
and U6836 (N_6836,N_2743,N_1037);
nand U6837 (N_6837,N_2412,N_1544);
and U6838 (N_6838,N_148,N_3401);
nor U6839 (N_6839,N_3229,N_1);
and U6840 (N_6840,N_632,N_3276);
nor U6841 (N_6841,N_1719,N_2785);
and U6842 (N_6842,N_2510,N_1123);
and U6843 (N_6843,N_165,N_1504);
nand U6844 (N_6844,N_527,N_1754);
or U6845 (N_6845,N_3861,N_2273);
nor U6846 (N_6846,N_2921,N_3966);
or U6847 (N_6847,N_2685,N_2347);
nand U6848 (N_6848,N_230,N_1484);
or U6849 (N_6849,N_1509,N_1322);
or U6850 (N_6850,N_2341,N_1292);
or U6851 (N_6851,N_3698,N_3837);
nor U6852 (N_6852,N_3989,N_1588);
and U6853 (N_6853,N_348,N_2871);
or U6854 (N_6854,N_2972,N_3052);
nor U6855 (N_6855,N_509,N_3410);
and U6856 (N_6856,N_1017,N_2446);
nor U6857 (N_6857,N_2966,N_499);
and U6858 (N_6858,N_939,N_3548);
and U6859 (N_6859,N_2814,N_1809);
nor U6860 (N_6860,N_3707,N_631);
and U6861 (N_6861,N_2290,N_710);
nor U6862 (N_6862,N_3072,N_616);
or U6863 (N_6863,N_398,N_2434);
and U6864 (N_6864,N_1721,N_2120);
or U6865 (N_6865,N_1480,N_1132);
xnor U6866 (N_6866,N_2059,N_1984);
or U6867 (N_6867,N_420,N_450);
nand U6868 (N_6868,N_720,N_3855);
or U6869 (N_6869,N_7,N_3684);
and U6870 (N_6870,N_1301,N_124);
nand U6871 (N_6871,N_1123,N_2202);
nor U6872 (N_6872,N_1773,N_2852);
nor U6873 (N_6873,N_1810,N_946);
nor U6874 (N_6874,N_1640,N_3316);
or U6875 (N_6875,N_1295,N_560);
nor U6876 (N_6876,N_147,N_3518);
and U6877 (N_6877,N_2384,N_2807);
nand U6878 (N_6878,N_1873,N_1912);
or U6879 (N_6879,N_893,N_2349);
or U6880 (N_6880,N_315,N_551);
nor U6881 (N_6881,N_1893,N_1518);
and U6882 (N_6882,N_1723,N_857);
or U6883 (N_6883,N_1826,N_175);
xnor U6884 (N_6884,N_3750,N_1252);
nand U6885 (N_6885,N_330,N_3011);
or U6886 (N_6886,N_3086,N_3665);
and U6887 (N_6887,N_3747,N_924);
nand U6888 (N_6888,N_3597,N_3169);
and U6889 (N_6889,N_1878,N_1542);
nor U6890 (N_6890,N_467,N_3292);
nor U6891 (N_6891,N_3504,N_3357);
nand U6892 (N_6892,N_2505,N_1845);
and U6893 (N_6893,N_1590,N_2599);
or U6894 (N_6894,N_1666,N_957);
or U6895 (N_6895,N_2241,N_1328);
nand U6896 (N_6896,N_896,N_2841);
nand U6897 (N_6897,N_1958,N_2840);
or U6898 (N_6898,N_3612,N_819);
nor U6899 (N_6899,N_768,N_2159);
nor U6900 (N_6900,N_2620,N_3290);
and U6901 (N_6901,N_3780,N_885);
and U6902 (N_6902,N_2428,N_3301);
nor U6903 (N_6903,N_2448,N_2533);
nand U6904 (N_6904,N_2868,N_145);
or U6905 (N_6905,N_2065,N_2994);
and U6906 (N_6906,N_2180,N_2728);
or U6907 (N_6907,N_2765,N_323);
and U6908 (N_6908,N_338,N_3255);
nand U6909 (N_6909,N_870,N_3551);
nand U6910 (N_6910,N_628,N_3658);
or U6911 (N_6911,N_703,N_3689);
and U6912 (N_6912,N_2729,N_3367);
xor U6913 (N_6913,N_890,N_3774);
nand U6914 (N_6914,N_1681,N_3615);
and U6915 (N_6915,N_3714,N_3745);
and U6916 (N_6916,N_3918,N_583);
and U6917 (N_6917,N_690,N_1477);
or U6918 (N_6918,N_3787,N_3433);
xor U6919 (N_6919,N_3882,N_22);
and U6920 (N_6920,N_2646,N_872);
nand U6921 (N_6921,N_3782,N_242);
nor U6922 (N_6922,N_1656,N_3454);
or U6923 (N_6923,N_2520,N_63);
nor U6924 (N_6924,N_1198,N_2951);
or U6925 (N_6925,N_2999,N_2916);
and U6926 (N_6926,N_2275,N_2738);
nand U6927 (N_6927,N_3862,N_2266);
and U6928 (N_6928,N_2660,N_1242);
nor U6929 (N_6929,N_3894,N_1765);
nor U6930 (N_6930,N_3039,N_2143);
nor U6931 (N_6931,N_2761,N_2918);
or U6932 (N_6932,N_708,N_3319);
nor U6933 (N_6933,N_412,N_2689);
and U6934 (N_6934,N_321,N_2916);
nand U6935 (N_6935,N_415,N_1257);
and U6936 (N_6936,N_1089,N_3741);
and U6937 (N_6937,N_1539,N_1967);
or U6938 (N_6938,N_1830,N_2093);
or U6939 (N_6939,N_2744,N_1432);
nor U6940 (N_6940,N_3987,N_416);
and U6941 (N_6941,N_179,N_217);
nor U6942 (N_6942,N_122,N_3928);
or U6943 (N_6943,N_3232,N_1594);
nor U6944 (N_6944,N_2815,N_3454);
nor U6945 (N_6945,N_1887,N_3716);
nand U6946 (N_6946,N_776,N_2368);
or U6947 (N_6947,N_3690,N_3244);
or U6948 (N_6948,N_2599,N_1405);
and U6949 (N_6949,N_463,N_3293);
and U6950 (N_6950,N_3918,N_527);
and U6951 (N_6951,N_3582,N_3549);
nand U6952 (N_6952,N_3574,N_2553);
and U6953 (N_6953,N_3873,N_3761);
nand U6954 (N_6954,N_984,N_587);
nor U6955 (N_6955,N_496,N_1911);
and U6956 (N_6956,N_3377,N_1247);
and U6957 (N_6957,N_2929,N_2124);
and U6958 (N_6958,N_3202,N_2482);
nor U6959 (N_6959,N_92,N_2844);
nand U6960 (N_6960,N_183,N_1745);
or U6961 (N_6961,N_1306,N_232);
and U6962 (N_6962,N_2441,N_1439);
and U6963 (N_6963,N_603,N_2637);
nor U6964 (N_6964,N_2299,N_827);
nor U6965 (N_6965,N_1770,N_650);
and U6966 (N_6966,N_2927,N_1195);
or U6967 (N_6967,N_970,N_3062);
or U6968 (N_6968,N_3265,N_2494);
nand U6969 (N_6969,N_1517,N_677);
and U6970 (N_6970,N_2844,N_1492);
nand U6971 (N_6971,N_2440,N_385);
nor U6972 (N_6972,N_3803,N_3185);
nand U6973 (N_6973,N_3012,N_1458);
nand U6974 (N_6974,N_1537,N_3012);
nand U6975 (N_6975,N_2495,N_2954);
and U6976 (N_6976,N_1092,N_883);
nor U6977 (N_6977,N_333,N_1520);
nand U6978 (N_6978,N_2948,N_558);
or U6979 (N_6979,N_3471,N_26);
and U6980 (N_6980,N_261,N_1401);
or U6981 (N_6981,N_1658,N_2237);
and U6982 (N_6982,N_552,N_3358);
nand U6983 (N_6983,N_3366,N_2148);
and U6984 (N_6984,N_2348,N_2772);
nand U6985 (N_6985,N_3070,N_3033);
and U6986 (N_6986,N_1830,N_3900);
nand U6987 (N_6987,N_1878,N_3741);
nor U6988 (N_6988,N_2013,N_439);
and U6989 (N_6989,N_1198,N_2019);
nand U6990 (N_6990,N_561,N_589);
or U6991 (N_6991,N_3510,N_3589);
and U6992 (N_6992,N_516,N_547);
or U6993 (N_6993,N_2897,N_1608);
and U6994 (N_6994,N_297,N_2598);
or U6995 (N_6995,N_3090,N_243);
nor U6996 (N_6996,N_1953,N_2727);
and U6997 (N_6997,N_2971,N_254);
and U6998 (N_6998,N_2201,N_709);
nand U6999 (N_6999,N_3898,N_2566);
nand U7000 (N_7000,N_2225,N_92);
nor U7001 (N_7001,N_3500,N_1867);
nand U7002 (N_7002,N_1410,N_3952);
or U7003 (N_7003,N_3893,N_3661);
and U7004 (N_7004,N_791,N_1184);
nand U7005 (N_7005,N_3597,N_2992);
or U7006 (N_7006,N_460,N_649);
nand U7007 (N_7007,N_1317,N_958);
nor U7008 (N_7008,N_3375,N_1646);
nor U7009 (N_7009,N_2414,N_1615);
nand U7010 (N_7010,N_3316,N_3630);
nand U7011 (N_7011,N_802,N_659);
or U7012 (N_7012,N_1084,N_2654);
and U7013 (N_7013,N_1967,N_3265);
and U7014 (N_7014,N_1456,N_1802);
nor U7015 (N_7015,N_3202,N_913);
nor U7016 (N_7016,N_3452,N_3236);
nor U7017 (N_7017,N_399,N_2716);
or U7018 (N_7018,N_601,N_1404);
or U7019 (N_7019,N_850,N_364);
nand U7020 (N_7020,N_552,N_2324);
nand U7021 (N_7021,N_3521,N_3614);
and U7022 (N_7022,N_2185,N_3704);
and U7023 (N_7023,N_3335,N_1243);
or U7024 (N_7024,N_274,N_1735);
nor U7025 (N_7025,N_3278,N_3137);
nor U7026 (N_7026,N_879,N_2959);
or U7027 (N_7027,N_744,N_1245);
nand U7028 (N_7028,N_3745,N_562);
nor U7029 (N_7029,N_187,N_1808);
and U7030 (N_7030,N_1702,N_266);
and U7031 (N_7031,N_2598,N_2272);
nor U7032 (N_7032,N_1521,N_3665);
and U7033 (N_7033,N_2128,N_301);
or U7034 (N_7034,N_2042,N_819);
or U7035 (N_7035,N_225,N_2257);
and U7036 (N_7036,N_1185,N_3421);
or U7037 (N_7037,N_3960,N_733);
nand U7038 (N_7038,N_1210,N_2215);
or U7039 (N_7039,N_40,N_212);
nand U7040 (N_7040,N_611,N_17);
nand U7041 (N_7041,N_3097,N_2319);
and U7042 (N_7042,N_1328,N_2212);
or U7043 (N_7043,N_2122,N_3046);
nor U7044 (N_7044,N_2324,N_2585);
or U7045 (N_7045,N_3692,N_3962);
nor U7046 (N_7046,N_359,N_2394);
and U7047 (N_7047,N_2318,N_1336);
and U7048 (N_7048,N_1897,N_1747);
or U7049 (N_7049,N_2050,N_1826);
or U7050 (N_7050,N_3155,N_1552);
nand U7051 (N_7051,N_3363,N_1310);
nand U7052 (N_7052,N_1901,N_2360);
or U7053 (N_7053,N_1974,N_3540);
or U7054 (N_7054,N_546,N_1703);
nand U7055 (N_7055,N_2302,N_2846);
or U7056 (N_7056,N_3748,N_407);
and U7057 (N_7057,N_533,N_3432);
nand U7058 (N_7058,N_1291,N_3810);
or U7059 (N_7059,N_3498,N_1647);
nor U7060 (N_7060,N_1233,N_2729);
nor U7061 (N_7061,N_1205,N_1707);
nand U7062 (N_7062,N_3928,N_3383);
or U7063 (N_7063,N_1155,N_1664);
or U7064 (N_7064,N_1616,N_2575);
nand U7065 (N_7065,N_2463,N_3719);
or U7066 (N_7066,N_1320,N_2422);
nand U7067 (N_7067,N_2428,N_2292);
nand U7068 (N_7068,N_1492,N_2052);
or U7069 (N_7069,N_2234,N_1395);
or U7070 (N_7070,N_2769,N_1472);
and U7071 (N_7071,N_3722,N_2867);
and U7072 (N_7072,N_1205,N_3554);
or U7073 (N_7073,N_1723,N_943);
and U7074 (N_7074,N_1089,N_1451);
nor U7075 (N_7075,N_1708,N_2289);
or U7076 (N_7076,N_2285,N_3258);
or U7077 (N_7077,N_56,N_2129);
or U7078 (N_7078,N_3122,N_2081);
and U7079 (N_7079,N_2402,N_2817);
and U7080 (N_7080,N_2633,N_2103);
or U7081 (N_7081,N_317,N_3720);
and U7082 (N_7082,N_3068,N_2090);
nor U7083 (N_7083,N_3331,N_2201);
or U7084 (N_7084,N_1870,N_3166);
nand U7085 (N_7085,N_3017,N_2912);
or U7086 (N_7086,N_2457,N_2033);
nor U7087 (N_7087,N_1670,N_3309);
and U7088 (N_7088,N_338,N_3337);
nor U7089 (N_7089,N_3199,N_3449);
nor U7090 (N_7090,N_916,N_1523);
and U7091 (N_7091,N_103,N_1838);
nand U7092 (N_7092,N_1740,N_3534);
and U7093 (N_7093,N_1097,N_3553);
nand U7094 (N_7094,N_1891,N_203);
nor U7095 (N_7095,N_3145,N_1943);
nor U7096 (N_7096,N_570,N_2713);
nand U7097 (N_7097,N_232,N_2730);
nor U7098 (N_7098,N_2625,N_3407);
nand U7099 (N_7099,N_2749,N_2635);
and U7100 (N_7100,N_3904,N_2398);
nor U7101 (N_7101,N_2853,N_3876);
nand U7102 (N_7102,N_3961,N_2176);
and U7103 (N_7103,N_3394,N_3259);
nand U7104 (N_7104,N_3494,N_3856);
or U7105 (N_7105,N_3650,N_644);
nand U7106 (N_7106,N_753,N_2239);
nor U7107 (N_7107,N_828,N_2028);
nor U7108 (N_7108,N_2135,N_2958);
nor U7109 (N_7109,N_1499,N_1946);
and U7110 (N_7110,N_565,N_1466);
or U7111 (N_7111,N_2470,N_1755);
nand U7112 (N_7112,N_3372,N_2565);
nand U7113 (N_7113,N_3682,N_2084);
nand U7114 (N_7114,N_1998,N_1970);
or U7115 (N_7115,N_1039,N_3558);
and U7116 (N_7116,N_2013,N_554);
or U7117 (N_7117,N_3046,N_385);
nand U7118 (N_7118,N_3553,N_1966);
nand U7119 (N_7119,N_1790,N_369);
or U7120 (N_7120,N_659,N_2155);
or U7121 (N_7121,N_563,N_177);
nand U7122 (N_7122,N_2856,N_2507);
and U7123 (N_7123,N_2549,N_2336);
and U7124 (N_7124,N_3739,N_1254);
nor U7125 (N_7125,N_1251,N_1395);
or U7126 (N_7126,N_2504,N_230);
and U7127 (N_7127,N_2308,N_256);
nand U7128 (N_7128,N_711,N_3277);
nand U7129 (N_7129,N_3422,N_175);
or U7130 (N_7130,N_1168,N_142);
nand U7131 (N_7131,N_2401,N_2493);
nor U7132 (N_7132,N_3172,N_3889);
and U7133 (N_7133,N_3062,N_2184);
or U7134 (N_7134,N_2403,N_3003);
nor U7135 (N_7135,N_3691,N_1888);
or U7136 (N_7136,N_3190,N_1095);
nor U7137 (N_7137,N_990,N_2414);
and U7138 (N_7138,N_2279,N_78);
and U7139 (N_7139,N_333,N_1174);
or U7140 (N_7140,N_1614,N_2113);
or U7141 (N_7141,N_1117,N_3153);
nor U7142 (N_7142,N_2244,N_1214);
or U7143 (N_7143,N_2307,N_2769);
xor U7144 (N_7144,N_1503,N_1310);
nand U7145 (N_7145,N_2975,N_2523);
xor U7146 (N_7146,N_1847,N_323);
nand U7147 (N_7147,N_3543,N_1098);
and U7148 (N_7148,N_1118,N_612);
or U7149 (N_7149,N_708,N_3199);
and U7150 (N_7150,N_2850,N_2494);
and U7151 (N_7151,N_668,N_1174);
nand U7152 (N_7152,N_3073,N_3017);
nand U7153 (N_7153,N_3075,N_3316);
or U7154 (N_7154,N_2434,N_2314);
and U7155 (N_7155,N_3563,N_2685);
nor U7156 (N_7156,N_1520,N_1123);
and U7157 (N_7157,N_1281,N_1432);
and U7158 (N_7158,N_1196,N_3090);
nor U7159 (N_7159,N_1927,N_2395);
nor U7160 (N_7160,N_1933,N_373);
nand U7161 (N_7161,N_1417,N_3671);
nor U7162 (N_7162,N_3500,N_1537);
nand U7163 (N_7163,N_60,N_3690);
and U7164 (N_7164,N_1815,N_722);
nor U7165 (N_7165,N_2983,N_306);
nor U7166 (N_7166,N_183,N_1695);
nor U7167 (N_7167,N_2844,N_3050);
and U7168 (N_7168,N_1234,N_3563);
or U7169 (N_7169,N_932,N_3648);
nor U7170 (N_7170,N_3447,N_3009);
or U7171 (N_7171,N_3855,N_2178);
nand U7172 (N_7172,N_552,N_284);
nor U7173 (N_7173,N_3690,N_3389);
nand U7174 (N_7174,N_3127,N_3199);
nand U7175 (N_7175,N_3864,N_3175);
nor U7176 (N_7176,N_2083,N_3066);
nand U7177 (N_7177,N_2817,N_2889);
and U7178 (N_7178,N_2750,N_3347);
nand U7179 (N_7179,N_805,N_233);
nor U7180 (N_7180,N_3359,N_196);
and U7181 (N_7181,N_1285,N_3537);
nor U7182 (N_7182,N_2224,N_3159);
nor U7183 (N_7183,N_1330,N_2355);
nand U7184 (N_7184,N_2477,N_1442);
and U7185 (N_7185,N_2045,N_2454);
or U7186 (N_7186,N_179,N_3944);
nand U7187 (N_7187,N_1592,N_540);
nor U7188 (N_7188,N_1437,N_3069);
nor U7189 (N_7189,N_2798,N_1158);
and U7190 (N_7190,N_1621,N_3594);
and U7191 (N_7191,N_2859,N_3543);
or U7192 (N_7192,N_2401,N_572);
nor U7193 (N_7193,N_2393,N_1736);
and U7194 (N_7194,N_3828,N_1909);
nor U7195 (N_7195,N_2192,N_3618);
nor U7196 (N_7196,N_3220,N_2788);
and U7197 (N_7197,N_1745,N_1679);
nor U7198 (N_7198,N_260,N_3506);
xor U7199 (N_7199,N_1819,N_3230);
and U7200 (N_7200,N_1891,N_1135);
nor U7201 (N_7201,N_315,N_575);
nor U7202 (N_7202,N_2722,N_3484);
nand U7203 (N_7203,N_1345,N_2192);
nand U7204 (N_7204,N_2163,N_3002);
and U7205 (N_7205,N_2616,N_568);
nor U7206 (N_7206,N_138,N_3327);
nand U7207 (N_7207,N_903,N_1869);
and U7208 (N_7208,N_1604,N_2399);
or U7209 (N_7209,N_2006,N_236);
and U7210 (N_7210,N_3834,N_3378);
and U7211 (N_7211,N_3399,N_1084);
nor U7212 (N_7212,N_3828,N_1227);
and U7213 (N_7213,N_3755,N_3599);
or U7214 (N_7214,N_863,N_231);
and U7215 (N_7215,N_1972,N_1678);
nor U7216 (N_7216,N_1141,N_2220);
nand U7217 (N_7217,N_1643,N_129);
nor U7218 (N_7218,N_2766,N_137);
xor U7219 (N_7219,N_170,N_3581);
and U7220 (N_7220,N_192,N_900);
or U7221 (N_7221,N_34,N_2430);
nand U7222 (N_7222,N_2406,N_1363);
nand U7223 (N_7223,N_3315,N_2672);
nor U7224 (N_7224,N_2109,N_3319);
nor U7225 (N_7225,N_3217,N_2245);
and U7226 (N_7226,N_1286,N_2429);
and U7227 (N_7227,N_2114,N_1684);
nand U7228 (N_7228,N_3920,N_1677);
nor U7229 (N_7229,N_1266,N_2322);
nor U7230 (N_7230,N_1934,N_3679);
and U7231 (N_7231,N_3813,N_3855);
nand U7232 (N_7232,N_2389,N_810);
or U7233 (N_7233,N_2163,N_3600);
and U7234 (N_7234,N_3840,N_3934);
nand U7235 (N_7235,N_1710,N_344);
or U7236 (N_7236,N_1700,N_1246);
nor U7237 (N_7237,N_3715,N_1258);
nor U7238 (N_7238,N_1926,N_2413);
nand U7239 (N_7239,N_2650,N_2357);
nor U7240 (N_7240,N_1453,N_970);
or U7241 (N_7241,N_1367,N_48);
or U7242 (N_7242,N_2649,N_1906);
or U7243 (N_7243,N_3413,N_3063);
nor U7244 (N_7244,N_106,N_1945);
or U7245 (N_7245,N_2594,N_2036);
nand U7246 (N_7246,N_580,N_429);
and U7247 (N_7247,N_2870,N_3828);
xor U7248 (N_7248,N_1740,N_1454);
and U7249 (N_7249,N_23,N_2283);
nand U7250 (N_7250,N_715,N_2440);
nand U7251 (N_7251,N_3253,N_2938);
or U7252 (N_7252,N_3470,N_412);
or U7253 (N_7253,N_457,N_3729);
or U7254 (N_7254,N_3976,N_1092);
or U7255 (N_7255,N_698,N_1344);
and U7256 (N_7256,N_2106,N_337);
nor U7257 (N_7257,N_33,N_3439);
or U7258 (N_7258,N_3135,N_2727);
nand U7259 (N_7259,N_3774,N_2722);
nor U7260 (N_7260,N_430,N_3977);
and U7261 (N_7261,N_2113,N_1008);
nand U7262 (N_7262,N_3442,N_3457);
and U7263 (N_7263,N_1191,N_1958);
nor U7264 (N_7264,N_2024,N_2679);
and U7265 (N_7265,N_3075,N_2225);
or U7266 (N_7266,N_1898,N_1629);
and U7267 (N_7267,N_1408,N_1442);
nor U7268 (N_7268,N_738,N_605);
nor U7269 (N_7269,N_3081,N_1120);
and U7270 (N_7270,N_1926,N_271);
nand U7271 (N_7271,N_3286,N_1912);
nand U7272 (N_7272,N_34,N_354);
or U7273 (N_7273,N_3019,N_1815);
and U7274 (N_7274,N_172,N_225);
nand U7275 (N_7275,N_1413,N_1200);
or U7276 (N_7276,N_3685,N_2747);
or U7277 (N_7277,N_1152,N_1263);
nor U7278 (N_7278,N_1855,N_906);
nor U7279 (N_7279,N_2766,N_2187);
or U7280 (N_7280,N_1390,N_1681);
or U7281 (N_7281,N_3220,N_1649);
nor U7282 (N_7282,N_2499,N_1735);
nor U7283 (N_7283,N_3711,N_2985);
nor U7284 (N_7284,N_3030,N_865);
nand U7285 (N_7285,N_390,N_3016);
nor U7286 (N_7286,N_2745,N_1077);
or U7287 (N_7287,N_2201,N_2602);
and U7288 (N_7288,N_1676,N_963);
nand U7289 (N_7289,N_2374,N_1199);
or U7290 (N_7290,N_1561,N_675);
nor U7291 (N_7291,N_597,N_2159);
nor U7292 (N_7292,N_3585,N_2181);
nor U7293 (N_7293,N_354,N_2959);
and U7294 (N_7294,N_1356,N_968);
nand U7295 (N_7295,N_1602,N_2203);
and U7296 (N_7296,N_2271,N_202);
nor U7297 (N_7297,N_3963,N_359);
nand U7298 (N_7298,N_633,N_875);
or U7299 (N_7299,N_2535,N_742);
and U7300 (N_7300,N_3606,N_1212);
nor U7301 (N_7301,N_385,N_142);
nand U7302 (N_7302,N_1014,N_661);
or U7303 (N_7303,N_1483,N_657);
nor U7304 (N_7304,N_770,N_715);
or U7305 (N_7305,N_221,N_3502);
nor U7306 (N_7306,N_1964,N_1343);
xnor U7307 (N_7307,N_2717,N_438);
and U7308 (N_7308,N_2598,N_343);
or U7309 (N_7309,N_2680,N_3766);
nor U7310 (N_7310,N_853,N_1406);
and U7311 (N_7311,N_676,N_1895);
and U7312 (N_7312,N_148,N_282);
or U7313 (N_7313,N_454,N_2386);
nand U7314 (N_7314,N_3137,N_2579);
or U7315 (N_7315,N_611,N_1022);
nor U7316 (N_7316,N_1155,N_3287);
and U7317 (N_7317,N_3930,N_2913);
nor U7318 (N_7318,N_3408,N_2800);
or U7319 (N_7319,N_164,N_3767);
and U7320 (N_7320,N_850,N_1883);
and U7321 (N_7321,N_251,N_1244);
or U7322 (N_7322,N_1138,N_960);
nand U7323 (N_7323,N_3966,N_1739);
nor U7324 (N_7324,N_2581,N_823);
or U7325 (N_7325,N_2796,N_169);
nor U7326 (N_7326,N_376,N_2951);
or U7327 (N_7327,N_1594,N_2962);
or U7328 (N_7328,N_1871,N_175);
or U7329 (N_7329,N_1257,N_1448);
nor U7330 (N_7330,N_3733,N_1189);
or U7331 (N_7331,N_2034,N_744);
or U7332 (N_7332,N_1986,N_1334);
nand U7333 (N_7333,N_1799,N_1838);
and U7334 (N_7334,N_884,N_1162);
nor U7335 (N_7335,N_3212,N_3248);
nand U7336 (N_7336,N_550,N_3979);
or U7337 (N_7337,N_2064,N_290);
nor U7338 (N_7338,N_840,N_2745);
nor U7339 (N_7339,N_3369,N_2086);
and U7340 (N_7340,N_2257,N_3590);
or U7341 (N_7341,N_2951,N_3322);
and U7342 (N_7342,N_108,N_332);
and U7343 (N_7343,N_279,N_3855);
and U7344 (N_7344,N_2281,N_2905);
and U7345 (N_7345,N_170,N_3950);
xor U7346 (N_7346,N_1852,N_3605);
and U7347 (N_7347,N_3071,N_1867);
or U7348 (N_7348,N_3383,N_2611);
nand U7349 (N_7349,N_2960,N_3608);
or U7350 (N_7350,N_1715,N_2013);
nor U7351 (N_7351,N_1014,N_1470);
xnor U7352 (N_7352,N_2794,N_3774);
and U7353 (N_7353,N_2390,N_2512);
and U7354 (N_7354,N_2372,N_3203);
or U7355 (N_7355,N_2406,N_3987);
nor U7356 (N_7356,N_1614,N_1989);
nor U7357 (N_7357,N_1784,N_2648);
and U7358 (N_7358,N_3734,N_1770);
nand U7359 (N_7359,N_1900,N_1953);
and U7360 (N_7360,N_2292,N_1528);
and U7361 (N_7361,N_490,N_3427);
nor U7362 (N_7362,N_1732,N_1696);
xor U7363 (N_7363,N_1333,N_1365);
and U7364 (N_7364,N_3403,N_936);
or U7365 (N_7365,N_1545,N_3625);
and U7366 (N_7366,N_2072,N_3463);
or U7367 (N_7367,N_2390,N_3478);
nor U7368 (N_7368,N_2312,N_3968);
nor U7369 (N_7369,N_663,N_991);
or U7370 (N_7370,N_101,N_932);
or U7371 (N_7371,N_862,N_1078);
nand U7372 (N_7372,N_2664,N_1688);
nand U7373 (N_7373,N_2923,N_1782);
and U7374 (N_7374,N_2704,N_3326);
nand U7375 (N_7375,N_1533,N_1386);
or U7376 (N_7376,N_3777,N_3446);
or U7377 (N_7377,N_3687,N_1447);
nor U7378 (N_7378,N_757,N_775);
and U7379 (N_7379,N_3769,N_226);
nor U7380 (N_7380,N_205,N_491);
and U7381 (N_7381,N_561,N_3040);
and U7382 (N_7382,N_542,N_28);
and U7383 (N_7383,N_2842,N_181);
nand U7384 (N_7384,N_13,N_590);
nor U7385 (N_7385,N_930,N_1529);
nor U7386 (N_7386,N_553,N_882);
nor U7387 (N_7387,N_890,N_3989);
and U7388 (N_7388,N_1364,N_833);
or U7389 (N_7389,N_2550,N_715);
and U7390 (N_7390,N_2232,N_1440);
or U7391 (N_7391,N_2402,N_3601);
nor U7392 (N_7392,N_3323,N_3342);
nor U7393 (N_7393,N_855,N_3661);
and U7394 (N_7394,N_2812,N_2549);
nor U7395 (N_7395,N_1297,N_3932);
and U7396 (N_7396,N_876,N_2589);
nor U7397 (N_7397,N_2525,N_17);
nand U7398 (N_7398,N_2419,N_1216);
and U7399 (N_7399,N_1653,N_3225);
xnor U7400 (N_7400,N_3700,N_2285);
nand U7401 (N_7401,N_1877,N_1891);
nor U7402 (N_7402,N_3184,N_2912);
and U7403 (N_7403,N_430,N_606);
nor U7404 (N_7404,N_208,N_1118);
nand U7405 (N_7405,N_1023,N_3991);
or U7406 (N_7406,N_2539,N_3798);
nor U7407 (N_7407,N_3601,N_3415);
or U7408 (N_7408,N_1207,N_2461);
nor U7409 (N_7409,N_2584,N_1190);
nor U7410 (N_7410,N_3630,N_653);
and U7411 (N_7411,N_989,N_3531);
and U7412 (N_7412,N_1109,N_1143);
and U7413 (N_7413,N_2307,N_1681);
nand U7414 (N_7414,N_2350,N_410);
and U7415 (N_7415,N_20,N_1606);
and U7416 (N_7416,N_1744,N_1895);
nand U7417 (N_7417,N_1647,N_3770);
nor U7418 (N_7418,N_3574,N_2202);
or U7419 (N_7419,N_1547,N_2666);
or U7420 (N_7420,N_493,N_3489);
nand U7421 (N_7421,N_1058,N_1544);
nor U7422 (N_7422,N_2707,N_2451);
and U7423 (N_7423,N_1930,N_1332);
nand U7424 (N_7424,N_2403,N_1158);
nand U7425 (N_7425,N_435,N_3240);
nand U7426 (N_7426,N_3500,N_3869);
or U7427 (N_7427,N_1766,N_3240);
nand U7428 (N_7428,N_1428,N_3242);
nand U7429 (N_7429,N_2977,N_3228);
or U7430 (N_7430,N_2813,N_2001);
and U7431 (N_7431,N_2202,N_2539);
nor U7432 (N_7432,N_3841,N_3779);
or U7433 (N_7433,N_3248,N_1637);
nor U7434 (N_7434,N_556,N_2128);
nand U7435 (N_7435,N_929,N_2738);
or U7436 (N_7436,N_454,N_3452);
and U7437 (N_7437,N_3059,N_679);
nor U7438 (N_7438,N_963,N_80);
nor U7439 (N_7439,N_1919,N_2440);
nor U7440 (N_7440,N_451,N_1380);
and U7441 (N_7441,N_3801,N_2419);
or U7442 (N_7442,N_1780,N_1337);
nand U7443 (N_7443,N_2041,N_187);
nand U7444 (N_7444,N_3499,N_26);
nand U7445 (N_7445,N_3071,N_1930);
nor U7446 (N_7446,N_169,N_346);
or U7447 (N_7447,N_3483,N_1539);
nor U7448 (N_7448,N_1106,N_2565);
and U7449 (N_7449,N_959,N_2673);
nand U7450 (N_7450,N_3992,N_2540);
and U7451 (N_7451,N_579,N_335);
xor U7452 (N_7452,N_521,N_101);
nand U7453 (N_7453,N_1634,N_2608);
and U7454 (N_7454,N_718,N_3726);
nor U7455 (N_7455,N_2877,N_641);
and U7456 (N_7456,N_2772,N_1016);
nor U7457 (N_7457,N_665,N_1972);
and U7458 (N_7458,N_684,N_3954);
or U7459 (N_7459,N_2234,N_1115);
nand U7460 (N_7460,N_1513,N_1756);
or U7461 (N_7461,N_1031,N_3665);
and U7462 (N_7462,N_3748,N_2430);
or U7463 (N_7463,N_3537,N_1057);
nor U7464 (N_7464,N_3001,N_563);
or U7465 (N_7465,N_2669,N_2562);
nor U7466 (N_7466,N_1648,N_1365);
or U7467 (N_7467,N_2828,N_1509);
nor U7468 (N_7468,N_2711,N_3701);
and U7469 (N_7469,N_3801,N_3604);
and U7470 (N_7470,N_3162,N_325);
and U7471 (N_7471,N_2095,N_1102);
nand U7472 (N_7472,N_3347,N_2996);
and U7473 (N_7473,N_1783,N_2731);
and U7474 (N_7474,N_813,N_42);
nor U7475 (N_7475,N_3527,N_1980);
and U7476 (N_7476,N_2205,N_1029);
or U7477 (N_7477,N_2993,N_2320);
or U7478 (N_7478,N_1935,N_3717);
nor U7479 (N_7479,N_3483,N_1913);
and U7480 (N_7480,N_1488,N_3755);
and U7481 (N_7481,N_3124,N_3818);
and U7482 (N_7482,N_1393,N_1358);
nand U7483 (N_7483,N_119,N_3400);
and U7484 (N_7484,N_8,N_3935);
nor U7485 (N_7485,N_801,N_3928);
and U7486 (N_7486,N_1818,N_2119);
or U7487 (N_7487,N_1691,N_2400);
nand U7488 (N_7488,N_1574,N_1316);
or U7489 (N_7489,N_1544,N_794);
or U7490 (N_7490,N_2266,N_2027);
and U7491 (N_7491,N_1973,N_2876);
nor U7492 (N_7492,N_3739,N_2354);
and U7493 (N_7493,N_537,N_481);
xor U7494 (N_7494,N_507,N_3664);
or U7495 (N_7495,N_3360,N_3036);
and U7496 (N_7496,N_838,N_3844);
nand U7497 (N_7497,N_3594,N_1734);
nand U7498 (N_7498,N_3920,N_445);
or U7499 (N_7499,N_797,N_1027);
xor U7500 (N_7500,N_1306,N_3159);
nand U7501 (N_7501,N_2136,N_1391);
nor U7502 (N_7502,N_1289,N_515);
nand U7503 (N_7503,N_265,N_437);
or U7504 (N_7504,N_3363,N_493);
nor U7505 (N_7505,N_204,N_2758);
and U7506 (N_7506,N_2582,N_362);
and U7507 (N_7507,N_1895,N_3250);
and U7508 (N_7508,N_3984,N_138);
nand U7509 (N_7509,N_1857,N_535);
or U7510 (N_7510,N_1673,N_3135);
or U7511 (N_7511,N_2952,N_1000);
nand U7512 (N_7512,N_144,N_2682);
nand U7513 (N_7513,N_3685,N_1891);
nand U7514 (N_7514,N_2920,N_2265);
or U7515 (N_7515,N_1506,N_1378);
and U7516 (N_7516,N_2449,N_199);
and U7517 (N_7517,N_315,N_2576);
nand U7518 (N_7518,N_3096,N_460);
nor U7519 (N_7519,N_2497,N_1331);
or U7520 (N_7520,N_3940,N_2500);
or U7521 (N_7521,N_828,N_2527);
or U7522 (N_7522,N_2259,N_2600);
and U7523 (N_7523,N_3564,N_73);
nor U7524 (N_7524,N_3756,N_2466);
or U7525 (N_7525,N_3332,N_1667);
and U7526 (N_7526,N_13,N_3632);
nor U7527 (N_7527,N_1526,N_2355);
nand U7528 (N_7528,N_430,N_2329);
nand U7529 (N_7529,N_2668,N_3105);
nand U7530 (N_7530,N_2819,N_2807);
and U7531 (N_7531,N_507,N_849);
nor U7532 (N_7532,N_1817,N_3085);
or U7533 (N_7533,N_1192,N_200);
and U7534 (N_7534,N_3136,N_3279);
nand U7535 (N_7535,N_1659,N_608);
or U7536 (N_7536,N_1742,N_1066);
nand U7537 (N_7537,N_2407,N_525);
nand U7538 (N_7538,N_1950,N_2840);
and U7539 (N_7539,N_558,N_1366);
or U7540 (N_7540,N_40,N_1145);
nand U7541 (N_7541,N_3406,N_2103);
and U7542 (N_7542,N_3235,N_547);
nor U7543 (N_7543,N_88,N_3012);
nor U7544 (N_7544,N_2187,N_2529);
and U7545 (N_7545,N_1435,N_90);
nor U7546 (N_7546,N_1408,N_345);
nor U7547 (N_7547,N_1711,N_670);
or U7548 (N_7548,N_3446,N_1681);
nand U7549 (N_7549,N_3406,N_186);
nand U7550 (N_7550,N_3607,N_461);
or U7551 (N_7551,N_2896,N_81);
nor U7552 (N_7552,N_1006,N_1681);
or U7553 (N_7553,N_1398,N_1060);
nor U7554 (N_7554,N_3375,N_1952);
or U7555 (N_7555,N_3153,N_2935);
nor U7556 (N_7556,N_2183,N_1189);
nor U7557 (N_7557,N_2121,N_930);
nor U7558 (N_7558,N_2216,N_1718);
nor U7559 (N_7559,N_741,N_2658);
nand U7560 (N_7560,N_3447,N_3005);
nor U7561 (N_7561,N_966,N_3558);
or U7562 (N_7562,N_1009,N_1931);
or U7563 (N_7563,N_1126,N_2586);
nand U7564 (N_7564,N_3959,N_3562);
or U7565 (N_7565,N_1832,N_2757);
nor U7566 (N_7566,N_912,N_356);
or U7567 (N_7567,N_144,N_823);
and U7568 (N_7568,N_765,N_1851);
or U7569 (N_7569,N_2049,N_2518);
or U7570 (N_7570,N_3944,N_3410);
nor U7571 (N_7571,N_1432,N_1188);
nor U7572 (N_7572,N_2363,N_1816);
or U7573 (N_7573,N_2992,N_2647);
nor U7574 (N_7574,N_2196,N_1706);
nor U7575 (N_7575,N_3288,N_3435);
and U7576 (N_7576,N_347,N_1995);
nor U7577 (N_7577,N_349,N_2169);
nor U7578 (N_7578,N_2339,N_1338);
and U7579 (N_7579,N_2529,N_3817);
nor U7580 (N_7580,N_602,N_3051);
and U7581 (N_7581,N_91,N_966);
and U7582 (N_7582,N_1776,N_1826);
nand U7583 (N_7583,N_35,N_3046);
nor U7584 (N_7584,N_1473,N_1877);
or U7585 (N_7585,N_3472,N_3634);
nor U7586 (N_7586,N_2689,N_140);
nand U7587 (N_7587,N_2204,N_2490);
nor U7588 (N_7588,N_1248,N_573);
nor U7589 (N_7589,N_3664,N_2846);
and U7590 (N_7590,N_1070,N_2837);
nand U7591 (N_7591,N_2590,N_3266);
nor U7592 (N_7592,N_1582,N_3796);
nor U7593 (N_7593,N_1863,N_3301);
and U7594 (N_7594,N_353,N_827);
nor U7595 (N_7595,N_579,N_1130);
or U7596 (N_7596,N_1169,N_628);
and U7597 (N_7597,N_2268,N_3757);
nand U7598 (N_7598,N_2234,N_286);
or U7599 (N_7599,N_669,N_2411);
xnor U7600 (N_7600,N_1671,N_3802);
or U7601 (N_7601,N_352,N_3916);
nor U7602 (N_7602,N_63,N_3152);
and U7603 (N_7603,N_347,N_485);
and U7604 (N_7604,N_516,N_1968);
xnor U7605 (N_7605,N_3505,N_1551);
nor U7606 (N_7606,N_1426,N_3129);
nand U7607 (N_7607,N_459,N_10);
or U7608 (N_7608,N_1164,N_1831);
nor U7609 (N_7609,N_305,N_3488);
nand U7610 (N_7610,N_625,N_1187);
or U7611 (N_7611,N_1074,N_1354);
nor U7612 (N_7612,N_793,N_1035);
and U7613 (N_7613,N_128,N_473);
nand U7614 (N_7614,N_1824,N_1002);
or U7615 (N_7615,N_2286,N_937);
nand U7616 (N_7616,N_3020,N_525);
xor U7617 (N_7617,N_3107,N_3404);
and U7618 (N_7618,N_3074,N_2511);
xnor U7619 (N_7619,N_2277,N_170);
nand U7620 (N_7620,N_1057,N_1453);
nand U7621 (N_7621,N_3536,N_419);
or U7622 (N_7622,N_1868,N_2133);
and U7623 (N_7623,N_1864,N_727);
and U7624 (N_7624,N_524,N_1003);
xnor U7625 (N_7625,N_2346,N_1281);
and U7626 (N_7626,N_542,N_715);
and U7627 (N_7627,N_2701,N_2673);
nor U7628 (N_7628,N_3746,N_3433);
nand U7629 (N_7629,N_761,N_1925);
or U7630 (N_7630,N_2038,N_2767);
xor U7631 (N_7631,N_1781,N_1587);
nor U7632 (N_7632,N_1522,N_2784);
nand U7633 (N_7633,N_3745,N_1188);
nor U7634 (N_7634,N_229,N_1081);
nor U7635 (N_7635,N_2127,N_2045);
nor U7636 (N_7636,N_695,N_3581);
nor U7637 (N_7637,N_278,N_3763);
and U7638 (N_7638,N_732,N_2881);
nor U7639 (N_7639,N_1790,N_3941);
and U7640 (N_7640,N_2361,N_1993);
or U7641 (N_7641,N_3980,N_3450);
nand U7642 (N_7642,N_3661,N_1716);
nor U7643 (N_7643,N_2804,N_2206);
and U7644 (N_7644,N_695,N_3692);
and U7645 (N_7645,N_3139,N_2362);
or U7646 (N_7646,N_2582,N_2479);
nor U7647 (N_7647,N_677,N_2648);
or U7648 (N_7648,N_754,N_1223);
and U7649 (N_7649,N_1874,N_3908);
nor U7650 (N_7650,N_2797,N_1030);
xnor U7651 (N_7651,N_3326,N_1788);
or U7652 (N_7652,N_2896,N_2952);
or U7653 (N_7653,N_2154,N_977);
nand U7654 (N_7654,N_1941,N_2550);
and U7655 (N_7655,N_452,N_376);
nand U7656 (N_7656,N_3519,N_702);
or U7657 (N_7657,N_1920,N_519);
and U7658 (N_7658,N_948,N_2331);
nand U7659 (N_7659,N_3432,N_2264);
and U7660 (N_7660,N_3155,N_1206);
xor U7661 (N_7661,N_318,N_2825);
or U7662 (N_7662,N_1681,N_1145);
nor U7663 (N_7663,N_3024,N_792);
nand U7664 (N_7664,N_1078,N_3480);
or U7665 (N_7665,N_1078,N_1260);
and U7666 (N_7666,N_549,N_2707);
nor U7667 (N_7667,N_1211,N_373);
nand U7668 (N_7668,N_3129,N_366);
or U7669 (N_7669,N_31,N_3569);
or U7670 (N_7670,N_1848,N_351);
nor U7671 (N_7671,N_2544,N_2864);
nor U7672 (N_7672,N_3296,N_1360);
nand U7673 (N_7673,N_2143,N_1813);
nand U7674 (N_7674,N_3584,N_714);
and U7675 (N_7675,N_179,N_1473);
nand U7676 (N_7676,N_39,N_2938);
and U7677 (N_7677,N_842,N_3203);
nand U7678 (N_7678,N_728,N_3001);
or U7679 (N_7679,N_3096,N_2942);
or U7680 (N_7680,N_1291,N_683);
nand U7681 (N_7681,N_441,N_608);
nor U7682 (N_7682,N_2369,N_2173);
nand U7683 (N_7683,N_243,N_2877);
and U7684 (N_7684,N_3741,N_423);
or U7685 (N_7685,N_2096,N_672);
or U7686 (N_7686,N_3903,N_3128);
nand U7687 (N_7687,N_1573,N_901);
and U7688 (N_7688,N_1231,N_2411);
and U7689 (N_7689,N_236,N_1746);
nor U7690 (N_7690,N_686,N_156);
and U7691 (N_7691,N_1342,N_839);
or U7692 (N_7692,N_1481,N_263);
and U7693 (N_7693,N_2559,N_479);
and U7694 (N_7694,N_1137,N_1261);
and U7695 (N_7695,N_2370,N_2284);
or U7696 (N_7696,N_2818,N_2404);
nand U7697 (N_7697,N_3151,N_1432);
nand U7698 (N_7698,N_1189,N_2771);
or U7699 (N_7699,N_1392,N_1484);
nor U7700 (N_7700,N_2265,N_3837);
nor U7701 (N_7701,N_2929,N_1197);
or U7702 (N_7702,N_647,N_1954);
nand U7703 (N_7703,N_1125,N_1894);
nor U7704 (N_7704,N_3583,N_3800);
nand U7705 (N_7705,N_1142,N_1024);
nor U7706 (N_7706,N_2946,N_1286);
nand U7707 (N_7707,N_3515,N_3672);
nand U7708 (N_7708,N_1168,N_3565);
nor U7709 (N_7709,N_1795,N_1393);
and U7710 (N_7710,N_3820,N_974);
nor U7711 (N_7711,N_2081,N_1990);
or U7712 (N_7712,N_2380,N_1073);
or U7713 (N_7713,N_1011,N_2928);
and U7714 (N_7714,N_3104,N_2445);
nand U7715 (N_7715,N_3695,N_1230);
nor U7716 (N_7716,N_3694,N_164);
nand U7717 (N_7717,N_3878,N_3810);
or U7718 (N_7718,N_3991,N_3702);
nor U7719 (N_7719,N_2241,N_3686);
nor U7720 (N_7720,N_174,N_1507);
and U7721 (N_7721,N_3606,N_3272);
or U7722 (N_7722,N_2727,N_3019);
nor U7723 (N_7723,N_997,N_1719);
and U7724 (N_7724,N_284,N_909);
nor U7725 (N_7725,N_2977,N_2417);
nand U7726 (N_7726,N_872,N_315);
nand U7727 (N_7727,N_3979,N_3322);
nand U7728 (N_7728,N_1762,N_2974);
nor U7729 (N_7729,N_2749,N_918);
nand U7730 (N_7730,N_2858,N_98);
nand U7731 (N_7731,N_3310,N_2504);
or U7732 (N_7732,N_587,N_2382);
nor U7733 (N_7733,N_3770,N_1369);
or U7734 (N_7734,N_563,N_78);
nor U7735 (N_7735,N_1407,N_862);
or U7736 (N_7736,N_3391,N_2579);
nor U7737 (N_7737,N_2901,N_1128);
nor U7738 (N_7738,N_1615,N_3040);
or U7739 (N_7739,N_2758,N_1153);
or U7740 (N_7740,N_317,N_3151);
or U7741 (N_7741,N_3074,N_2076);
and U7742 (N_7742,N_1330,N_1546);
nor U7743 (N_7743,N_3696,N_1252);
and U7744 (N_7744,N_3660,N_2139);
nor U7745 (N_7745,N_2972,N_2458);
nand U7746 (N_7746,N_236,N_2789);
nor U7747 (N_7747,N_3029,N_764);
nor U7748 (N_7748,N_1253,N_3471);
nor U7749 (N_7749,N_3542,N_344);
nand U7750 (N_7750,N_1790,N_2867);
and U7751 (N_7751,N_362,N_2252);
nand U7752 (N_7752,N_1012,N_3646);
nor U7753 (N_7753,N_36,N_742);
or U7754 (N_7754,N_522,N_3882);
nor U7755 (N_7755,N_3096,N_2268);
and U7756 (N_7756,N_322,N_304);
and U7757 (N_7757,N_2269,N_795);
xor U7758 (N_7758,N_2198,N_3074);
nor U7759 (N_7759,N_1184,N_553);
nor U7760 (N_7760,N_907,N_1646);
or U7761 (N_7761,N_204,N_3927);
or U7762 (N_7762,N_2587,N_1016);
xnor U7763 (N_7763,N_3563,N_3816);
nand U7764 (N_7764,N_1754,N_1024);
nor U7765 (N_7765,N_3204,N_2572);
or U7766 (N_7766,N_3047,N_3848);
nor U7767 (N_7767,N_2549,N_2354);
nor U7768 (N_7768,N_2222,N_3267);
nand U7769 (N_7769,N_2540,N_702);
or U7770 (N_7770,N_3091,N_861);
nor U7771 (N_7771,N_3069,N_2391);
and U7772 (N_7772,N_1015,N_3744);
and U7773 (N_7773,N_1094,N_15);
or U7774 (N_7774,N_347,N_3048);
nand U7775 (N_7775,N_3705,N_3305);
and U7776 (N_7776,N_3997,N_3537);
or U7777 (N_7777,N_2173,N_3031);
and U7778 (N_7778,N_3777,N_426);
or U7779 (N_7779,N_2628,N_112);
nor U7780 (N_7780,N_3309,N_195);
nand U7781 (N_7781,N_3421,N_2615);
or U7782 (N_7782,N_2211,N_2136);
nand U7783 (N_7783,N_1883,N_90);
and U7784 (N_7784,N_2350,N_2272);
or U7785 (N_7785,N_2969,N_2198);
nand U7786 (N_7786,N_2680,N_2765);
and U7787 (N_7787,N_1906,N_14);
or U7788 (N_7788,N_2904,N_3819);
and U7789 (N_7789,N_624,N_3482);
nand U7790 (N_7790,N_1460,N_3683);
or U7791 (N_7791,N_1504,N_2022);
or U7792 (N_7792,N_1391,N_2158);
nor U7793 (N_7793,N_3156,N_828);
and U7794 (N_7794,N_3787,N_1841);
or U7795 (N_7795,N_3031,N_299);
and U7796 (N_7796,N_3018,N_1400);
and U7797 (N_7797,N_2766,N_1949);
nor U7798 (N_7798,N_3814,N_2556);
or U7799 (N_7799,N_2913,N_2128);
xnor U7800 (N_7800,N_982,N_3303);
and U7801 (N_7801,N_104,N_1163);
xor U7802 (N_7802,N_1952,N_3424);
nor U7803 (N_7803,N_832,N_2640);
nand U7804 (N_7804,N_1741,N_1714);
or U7805 (N_7805,N_156,N_2044);
and U7806 (N_7806,N_1486,N_2328);
nor U7807 (N_7807,N_2491,N_3190);
or U7808 (N_7808,N_1443,N_3064);
or U7809 (N_7809,N_2179,N_2819);
nor U7810 (N_7810,N_2246,N_2425);
and U7811 (N_7811,N_358,N_1004);
or U7812 (N_7812,N_3863,N_2965);
and U7813 (N_7813,N_3603,N_1298);
and U7814 (N_7814,N_749,N_3456);
or U7815 (N_7815,N_3732,N_426);
nand U7816 (N_7816,N_2816,N_2527);
nand U7817 (N_7817,N_3073,N_1480);
and U7818 (N_7818,N_2448,N_1242);
nor U7819 (N_7819,N_1181,N_2447);
and U7820 (N_7820,N_1368,N_3264);
or U7821 (N_7821,N_3119,N_3433);
nor U7822 (N_7822,N_696,N_856);
nand U7823 (N_7823,N_2051,N_433);
nand U7824 (N_7824,N_899,N_508);
nand U7825 (N_7825,N_1615,N_1180);
or U7826 (N_7826,N_2908,N_3165);
nor U7827 (N_7827,N_1888,N_2775);
or U7828 (N_7828,N_3171,N_3384);
or U7829 (N_7829,N_1271,N_1768);
and U7830 (N_7830,N_269,N_3873);
or U7831 (N_7831,N_2852,N_48);
nor U7832 (N_7832,N_551,N_362);
nand U7833 (N_7833,N_3852,N_2131);
and U7834 (N_7834,N_1800,N_3902);
or U7835 (N_7835,N_1980,N_2984);
and U7836 (N_7836,N_1223,N_1739);
nor U7837 (N_7837,N_1167,N_364);
or U7838 (N_7838,N_3080,N_2613);
or U7839 (N_7839,N_3283,N_3700);
nand U7840 (N_7840,N_635,N_2470);
nand U7841 (N_7841,N_3791,N_1659);
nand U7842 (N_7842,N_3686,N_868);
or U7843 (N_7843,N_2958,N_2821);
nor U7844 (N_7844,N_2433,N_3954);
or U7845 (N_7845,N_2057,N_1809);
nor U7846 (N_7846,N_1409,N_1037);
and U7847 (N_7847,N_3716,N_2147);
and U7848 (N_7848,N_586,N_3563);
or U7849 (N_7849,N_3615,N_621);
or U7850 (N_7850,N_3233,N_3864);
nand U7851 (N_7851,N_702,N_747);
nand U7852 (N_7852,N_2127,N_2035);
and U7853 (N_7853,N_2694,N_3904);
and U7854 (N_7854,N_375,N_384);
and U7855 (N_7855,N_1734,N_959);
xnor U7856 (N_7856,N_502,N_163);
nand U7857 (N_7857,N_1415,N_1475);
nand U7858 (N_7858,N_2867,N_1355);
or U7859 (N_7859,N_2924,N_2296);
nor U7860 (N_7860,N_3468,N_3092);
or U7861 (N_7861,N_3956,N_3099);
nand U7862 (N_7862,N_2251,N_3799);
nor U7863 (N_7863,N_3529,N_613);
and U7864 (N_7864,N_2382,N_2367);
and U7865 (N_7865,N_2250,N_3618);
or U7866 (N_7866,N_444,N_3634);
nor U7867 (N_7867,N_3714,N_3194);
and U7868 (N_7868,N_865,N_1078);
and U7869 (N_7869,N_2934,N_3579);
nand U7870 (N_7870,N_3468,N_241);
nand U7871 (N_7871,N_3396,N_2604);
or U7872 (N_7872,N_2557,N_3097);
nor U7873 (N_7873,N_1162,N_78);
nor U7874 (N_7874,N_1097,N_2867);
nor U7875 (N_7875,N_1666,N_1307);
nor U7876 (N_7876,N_949,N_2858);
nand U7877 (N_7877,N_1489,N_577);
nor U7878 (N_7878,N_2021,N_1204);
or U7879 (N_7879,N_953,N_3205);
nand U7880 (N_7880,N_2170,N_3830);
and U7881 (N_7881,N_3965,N_3440);
nand U7882 (N_7882,N_990,N_734);
nor U7883 (N_7883,N_19,N_3511);
nand U7884 (N_7884,N_3083,N_1034);
xnor U7885 (N_7885,N_880,N_2619);
and U7886 (N_7886,N_102,N_3537);
nor U7887 (N_7887,N_2876,N_468);
or U7888 (N_7888,N_324,N_2253);
nor U7889 (N_7889,N_469,N_3845);
nand U7890 (N_7890,N_2227,N_197);
and U7891 (N_7891,N_3592,N_3255);
nand U7892 (N_7892,N_1534,N_515);
xor U7893 (N_7893,N_2417,N_1467);
and U7894 (N_7894,N_3427,N_1970);
nand U7895 (N_7895,N_542,N_1480);
nand U7896 (N_7896,N_552,N_2517);
nand U7897 (N_7897,N_1537,N_1972);
xnor U7898 (N_7898,N_947,N_3289);
nor U7899 (N_7899,N_1264,N_2782);
nand U7900 (N_7900,N_920,N_3491);
and U7901 (N_7901,N_2118,N_411);
and U7902 (N_7902,N_3316,N_3080);
nand U7903 (N_7903,N_1987,N_413);
nand U7904 (N_7904,N_2883,N_3759);
nand U7905 (N_7905,N_2988,N_1302);
nor U7906 (N_7906,N_1039,N_3387);
nor U7907 (N_7907,N_473,N_443);
or U7908 (N_7908,N_1126,N_3540);
nand U7909 (N_7909,N_3374,N_3783);
and U7910 (N_7910,N_3033,N_2812);
nand U7911 (N_7911,N_2642,N_54);
and U7912 (N_7912,N_2928,N_485);
nand U7913 (N_7913,N_1737,N_1535);
and U7914 (N_7914,N_3889,N_890);
or U7915 (N_7915,N_1247,N_2364);
nor U7916 (N_7916,N_2164,N_1680);
and U7917 (N_7917,N_649,N_3303);
nor U7918 (N_7918,N_3622,N_1776);
nand U7919 (N_7919,N_1939,N_2972);
nor U7920 (N_7920,N_2431,N_2661);
or U7921 (N_7921,N_406,N_487);
and U7922 (N_7922,N_2168,N_2722);
nor U7923 (N_7923,N_3443,N_3072);
nand U7924 (N_7924,N_2424,N_3331);
nor U7925 (N_7925,N_1180,N_855);
or U7926 (N_7926,N_3035,N_2164);
nor U7927 (N_7927,N_3596,N_1084);
nand U7928 (N_7928,N_3900,N_663);
nand U7929 (N_7929,N_420,N_2710);
or U7930 (N_7930,N_3111,N_790);
or U7931 (N_7931,N_2962,N_713);
nor U7932 (N_7932,N_401,N_1730);
nor U7933 (N_7933,N_1906,N_997);
nand U7934 (N_7934,N_2954,N_3571);
nand U7935 (N_7935,N_3488,N_3370);
nand U7936 (N_7936,N_2276,N_3324);
or U7937 (N_7937,N_3373,N_838);
or U7938 (N_7938,N_489,N_2364);
nor U7939 (N_7939,N_252,N_2479);
and U7940 (N_7940,N_3460,N_3053);
nor U7941 (N_7941,N_2669,N_2367);
and U7942 (N_7942,N_3154,N_1990);
and U7943 (N_7943,N_2608,N_2493);
nand U7944 (N_7944,N_1756,N_2384);
nor U7945 (N_7945,N_2959,N_1154);
nand U7946 (N_7946,N_3176,N_2109);
nor U7947 (N_7947,N_2014,N_1925);
and U7948 (N_7948,N_1079,N_2816);
or U7949 (N_7949,N_3665,N_3230);
or U7950 (N_7950,N_3166,N_3987);
nor U7951 (N_7951,N_1819,N_3668);
nand U7952 (N_7952,N_751,N_391);
nor U7953 (N_7953,N_864,N_2042);
nor U7954 (N_7954,N_314,N_3877);
nor U7955 (N_7955,N_206,N_2297);
or U7956 (N_7956,N_529,N_2037);
nor U7957 (N_7957,N_1879,N_383);
nor U7958 (N_7958,N_2991,N_1493);
nor U7959 (N_7959,N_116,N_2248);
nor U7960 (N_7960,N_2639,N_3005);
or U7961 (N_7961,N_3943,N_935);
or U7962 (N_7962,N_1387,N_1145);
nor U7963 (N_7963,N_1474,N_1042);
and U7964 (N_7964,N_2949,N_1487);
nand U7965 (N_7965,N_542,N_2093);
and U7966 (N_7966,N_721,N_3251);
or U7967 (N_7967,N_3759,N_2433);
nor U7968 (N_7968,N_2814,N_3174);
and U7969 (N_7969,N_754,N_1032);
and U7970 (N_7970,N_3656,N_1142);
nor U7971 (N_7971,N_1968,N_2642);
or U7972 (N_7972,N_6,N_3771);
or U7973 (N_7973,N_1285,N_1670);
nor U7974 (N_7974,N_2869,N_3028);
or U7975 (N_7975,N_2201,N_3874);
nand U7976 (N_7976,N_882,N_1723);
nor U7977 (N_7977,N_1910,N_90);
or U7978 (N_7978,N_46,N_2378);
and U7979 (N_7979,N_1482,N_3757);
nor U7980 (N_7980,N_3904,N_1886);
or U7981 (N_7981,N_2763,N_1005);
nor U7982 (N_7982,N_1690,N_3697);
xnor U7983 (N_7983,N_3766,N_2068);
nand U7984 (N_7984,N_3358,N_3257);
nor U7985 (N_7985,N_1400,N_117);
or U7986 (N_7986,N_1224,N_2483);
nand U7987 (N_7987,N_445,N_2950);
nand U7988 (N_7988,N_2186,N_3119);
nand U7989 (N_7989,N_2644,N_976);
nor U7990 (N_7990,N_2515,N_475);
nor U7991 (N_7991,N_3113,N_823);
or U7992 (N_7992,N_2478,N_3501);
and U7993 (N_7993,N_456,N_3894);
nor U7994 (N_7994,N_739,N_3276);
nor U7995 (N_7995,N_3947,N_729);
nor U7996 (N_7996,N_271,N_3546);
nor U7997 (N_7997,N_1557,N_1838);
nand U7998 (N_7998,N_2914,N_1423);
nand U7999 (N_7999,N_3965,N_394);
nand U8000 (N_8000,N_5823,N_7461);
nand U8001 (N_8001,N_4942,N_6968);
and U8002 (N_8002,N_4006,N_7989);
nand U8003 (N_8003,N_4127,N_7698);
nor U8004 (N_8004,N_5977,N_4517);
nor U8005 (N_8005,N_5042,N_4966);
nand U8006 (N_8006,N_4888,N_6250);
nand U8007 (N_8007,N_4373,N_5473);
and U8008 (N_8008,N_6994,N_7939);
nand U8009 (N_8009,N_5663,N_7747);
nand U8010 (N_8010,N_5273,N_6533);
nand U8011 (N_8011,N_4069,N_6448);
nor U8012 (N_8012,N_5645,N_4163);
nor U8013 (N_8013,N_5896,N_4145);
nand U8014 (N_8014,N_7202,N_4179);
nor U8015 (N_8015,N_4495,N_7595);
nor U8016 (N_8016,N_6975,N_5798);
and U8017 (N_8017,N_7699,N_4435);
or U8018 (N_8018,N_4235,N_4247);
nor U8019 (N_8019,N_5999,N_7280);
nand U8020 (N_8020,N_5375,N_4051);
or U8021 (N_8021,N_4479,N_5703);
nor U8022 (N_8022,N_4246,N_6151);
or U8023 (N_8023,N_7804,N_5722);
nor U8024 (N_8024,N_7648,N_6142);
and U8025 (N_8025,N_6768,N_4868);
nor U8026 (N_8026,N_6038,N_4560);
nor U8027 (N_8027,N_6338,N_5480);
nor U8028 (N_8028,N_4340,N_6271);
and U8029 (N_8029,N_5598,N_7117);
and U8030 (N_8030,N_5537,N_7673);
nand U8031 (N_8031,N_6444,N_6590);
nor U8032 (N_8032,N_7677,N_7009);
and U8033 (N_8033,N_6293,N_7971);
nor U8034 (N_8034,N_5214,N_7608);
and U8035 (N_8035,N_7314,N_5884);
nand U8036 (N_8036,N_4183,N_5370);
nor U8037 (N_8037,N_4763,N_6595);
nand U8038 (N_8038,N_4583,N_7669);
or U8039 (N_8039,N_4896,N_4335);
nand U8040 (N_8040,N_4515,N_6729);
or U8041 (N_8041,N_4122,N_7169);
nand U8042 (N_8042,N_4672,N_4241);
nor U8043 (N_8043,N_5837,N_4605);
or U8044 (N_8044,N_4107,N_6294);
nor U8045 (N_8045,N_4253,N_7089);
nor U8046 (N_8046,N_4550,N_7775);
nor U8047 (N_8047,N_7359,N_5257);
or U8048 (N_8048,N_5254,N_4131);
and U8049 (N_8049,N_7509,N_6800);
or U8050 (N_8050,N_5964,N_4167);
or U8051 (N_8051,N_7080,N_7030);
and U8052 (N_8052,N_5326,N_5835);
nor U8053 (N_8053,N_7703,N_6769);
or U8054 (N_8054,N_4879,N_7491);
nand U8055 (N_8055,N_6535,N_5074);
nand U8056 (N_8056,N_7445,N_5384);
or U8057 (N_8057,N_4432,N_6086);
nor U8058 (N_8058,N_5763,N_4033);
nand U8059 (N_8059,N_4255,N_6613);
and U8060 (N_8060,N_7610,N_5959);
and U8061 (N_8061,N_5578,N_4574);
nor U8062 (N_8062,N_6346,N_7094);
nor U8063 (N_8063,N_5551,N_4626);
nor U8064 (N_8064,N_4083,N_5543);
and U8065 (N_8065,N_6229,N_4624);
or U8066 (N_8066,N_6721,N_6664);
or U8067 (N_8067,N_7439,N_5724);
nor U8068 (N_8068,N_5617,N_4451);
xor U8069 (N_8069,N_6561,N_5653);
nor U8070 (N_8070,N_7734,N_4618);
or U8071 (N_8071,N_5250,N_7731);
nand U8072 (N_8072,N_6388,N_5531);
or U8073 (N_8073,N_6368,N_4393);
or U8074 (N_8074,N_5713,N_4042);
or U8075 (N_8075,N_7936,N_5987);
and U8076 (N_8076,N_5846,N_6493);
and U8077 (N_8077,N_6688,N_7497);
and U8078 (N_8078,N_5595,N_4477);
or U8079 (N_8079,N_7163,N_4237);
nand U8080 (N_8080,N_5008,N_6034);
or U8081 (N_8081,N_5600,N_4439);
or U8082 (N_8082,N_5237,N_4073);
or U8083 (N_8083,N_4749,N_4882);
nand U8084 (N_8084,N_5574,N_4846);
nor U8085 (N_8085,N_7861,N_5817);
nor U8086 (N_8086,N_4342,N_4512);
or U8087 (N_8087,N_5201,N_6818);
and U8088 (N_8088,N_7296,N_7988);
nand U8089 (N_8089,N_5101,N_4249);
or U8090 (N_8090,N_4712,N_5196);
and U8091 (N_8091,N_6801,N_5850);
and U8092 (N_8092,N_5168,N_7575);
nor U8093 (N_8093,N_6504,N_5686);
nor U8094 (N_8094,N_6720,N_4487);
and U8095 (N_8095,N_6371,N_7000);
or U8096 (N_8096,N_7612,N_4684);
and U8097 (N_8097,N_5677,N_4797);
and U8098 (N_8098,N_5532,N_4429);
or U8099 (N_8099,N_6989,N_6006);
nor U8100 (N_8100,N_6694,N_4243);
or U8101 (N_8101,N_4032,N_7859);
and U8102 (N_8102,N_7954,N_5943);
nand U8103 (N_8103,N_6364,N_4236);
nor U8104 (N_8104,N_4196,N_7417);
xor U8105 (N_8105,N_4481,N_4284);
nand U8106 (N_8106,N_7842,N_5380);
nand U8107 (N_8107,N_6681,N_5744);
nand U8108 (N_8108,N_5833,N_4799);
and U8109 (N_8109,N_7847,N_6358);
and U8110 (N_8110,N_7700,N_6269);
or U8111 (N_8111,N_5156,N_6712);
or U8112 (N_8112,N_7985,N_7334);
nand U8113 (N_8113,N_4115,N_4076);
and U8114 (N_8114,N_4627,N_5090);
nand U8115 (N_8115,N_6016,N_7161);
nor U8116 (N_8116,N_5826,N_4368);
nand U8117 (N_8117,N_7603,N_5199);
nor U8118 (N_8118,N_6013,N_7875);
and U8119 (N_8119,N_4058,N_6360);
and U8120 (N_8120,N_6410,N_7548);
or U8121 (N_8121,N_7654,N_6242);
nand U8122 (N_8122,N_4741,N_4589);
nand U8123 (N_8123,N_7421,N_4724);
or U8124 (N_8124,N_5770,N_4467);
or U8125 (N_8125,N_6702,N_4141);
and U8126 (N_8126,N_4314,N_5918);
or U8127 (N_8127,N_5401,N_7145);
or U8128 (N_8128,N_5174,N_4556);
and U8129 (N_8129,N_6866,N_4385);
or U8130 (N_8130,N_6017,N_4162);
or U8131 (N_8131,N_6891,N_6121);
nor U8132 (N_8132,N_5939,N_4187);
nand U8133 (N_8133,N_5172,N_6486);
or U8134 (N_8134,N_6884,N_4168);
nor U8135 (N_8135,N_6566,N_6012);
or U8136 (N_8136,N_5501,N_6734);
nand U8137 (N_8137,N_7887,N_4952);
nor U8138 (N_8138,N_5003,N_7776);
nand U8139 (N_8139,N_6287,N_7283);
nor U8140 (N_8140,N_7868,N_7542);
and U8141 (N_8141,N_5312,N_7362);
or U8142 (N_8142,N_6123,N_4416);
or U8143 (N_8143,N_4600,N_5961);
nor U8144 (N_8144,N_6265,N_4878);
and U8145 (N_8145,N_7377,N_5382);
or U8146 (N_8146,N_6683,N_6191);
or U8147 (N_8147,N_6862,N_7075);
and U8148 (N_8148,N_7708,N_5980);
nor U8149 (N_8149,N_6437,N_6926);
or U8150 (N_8150,N_4981,N_7401);
and U8151 (N_8151,N_7801,N_5671);
nor U8152 (N_8152,N_5970,N_4016);
nor U8153 (N_8153,N_4005,N_5742);
and U8154 (N_8154,N_6606,N_5762);
nand U8155 (N_8155,N_6028,N_5468);
or U8156 (N_8156,N_4388,N_7239);
nor U8157 (N_8157,N_4003,N_7164);
or U8158 (N_8158,N_5284,N_5586);
or U8159 (N_8159,N_7824,N_5181);
nand U8160 (N_8160,N_4395,N_5444);
and U8161 (N_8161,N_4787,N_5700);
and U8162 (N_8162,N_6266,N_6159);
nand U8163 (N_8163,N_6495,N_4527);
and U8164 (N_8164,N_7690,N_6983);
and U8165 (N_8165,N_7081,N_4662);
or U8166 (N_8166,N_4655,N_7771);
nand U8167 (N_8167,N_7388,N_5754);
and U8168 (N_8168,N_6666,N_4984);
and U8169 (N_8169,N_6218,N_6379);
nor U8170 (N_8170,N_7504,N_7532);
nor U8171 (N_8171,N_7286,N_7781);
nor U8172 (N_8172,N_5769,N_5550);
nor U8173 (N_8173,N_6095,N_7343);
or U8174 (N_8174,N_6275,N_7273);
and U8175 (N_8175,N_7136,N_4200);
and U8176 (N_8176,N_7079,N_5136);
or U8177 (N_8177,N_6436,N_5979);
nor U8178 (N_8178,N_5327,N_5052);
nand U8179 (N_8179,N_4802,N_4631);
or U8180 (N_8180,N_7885,N_7526);
nor U8181 (N_8181,N_4054,N_7645);
nand U8182 (N_8182,N_7931,N_4833);
nand U8183 (N_8183,N_5056,N_4424);
or U8184 (N_8184,N_6193,N_7162);
nor U8185 (N_8185,N_7990,N_5809);
nand U8186 (N_8186,N_5441,N_6829);
or U8187 (N_8187,N_6982,N_7996);
and U8188 (N_8188,N_7746,N_5832);
or U8189 (N_8189,N_4976,N_7973);
or U8190 (N_8190,N_5981,N_5492);
nor U8191 (N_8191,N_6319,N_7611);
or U8192 (N_8192,N_6995,N_6903);
nand U8193 (N_8193,N_4795,N_6053);
or U8194 (N_8194,N_5357,N_4931);
or U8195 (N_8195,N_7250,N_7469);
nor U8196 (N_8196,N_6967,N_7835);
nand U8197 (N_8197,N_6745,N_5889);
nor U8198 (N_8198,N_4172,N_5830);
nand U8199 (N_8199,N_5587,N_6794);
and U8200 (N_8200,N_5291,N_6585);
or U8201 (N_8201,N_7253,N_4336);
nor U8202 (N_8202,N_4806,N_4800);
nand U8203 (N_8203,N_5973,N_6166);
and U8204 (N_8204,N_7065,N_6161);
nor U8205 (N_8205,N_5041,N_5572);
nand U8206 (N_8206,N_6676,N_5938);
or U8207 (N_8207,N_7390,N_4372);
nand U8208 (N_8208,N_6747,N_6043);
or U8209 (N_8209,N_6211,N_4281);
nor U8210 (N_8210,N_7123,N_5394);
xor U8211 (N_8211,N_5496,N_5554);
nor U8212 (N_8212,N_5530,N_5180);
nand U8213 (N_8213,N_6010,N_4520);
and U8214 (N_8214,N_6460,N_5126);
or U8215 (N_8215,N_7862,N_7529);
or U8216 (N_8216,N_6552,N_5089);
nor U8217 (N_8217,N_7800,N_6812);
and U8218 (N_8218,N_7033,N_7400);
nor U8219 (N_8219,N_7368,N_6213);
or U8220 (N_8220,N_4238,N_7977);
or U8221 (N_8221,N_7440,N_6108);
and U8222 (N_8222,N_4607,N_6179);
nand U8223 (N_8223,N_7705,N_6523);
and U8224 (N_8224,N_4320,N_6872);
or U8225 (N_8225,N_5517,N_5355);
nand U8226 (N_8226,N_5428,N_4557);
nor U8227 (N_8227,N_7932,N_4581);
nor U8228 (N_8228,N_7658,N_4842);
and U8229 (N_8229,N_6517,N_4497);
nor U8230 (N_8230,N_6935,N_6393);
or U8231 (N_8231,N_4616,N_6612);
or U8232 (N_8232,N_5526,N_4921);
or U8233 (N_8233,N_6913,N_7053);
and U8234 (N_8234,N_7642,N_5911);
nor U8235 (N_8235,N_7451,N_6065);
nor U8236 (N_8236,N_4291,N_6069);
nor U8237 (N_8237,N_4022,N_7938);
nand U8238 (N_8238,N_6785,N_7070);
nand U8239 (N_8239,N_4035,N_5780);
and U8240 (N_8240,N_4551,N_4650);
and U8241 (N_8241,N_4519,N_4217);
nand U8242 (N_8242,N_7363,N_7992);
and U8243 (N_8243,N_6224,N_6744);
nor U8244 (N_8244,N_4608,N_5723);
nand U8245 (N_8245,N_6573,N_6646);
and U8246 (N_8246,N_6588,N_4754);
or U8247 (N_8247,N_5400,N_7981);
or U8248 (N_8248,N_5975,N_7599);
or U8249 (N_8249,N_4577,N_7688);
or U8250 (N_8250,N_4328,N_5229);
nand U8251 (N_8251,N_4904,N_7028);
or U8252 (N_8252,N_7966,N_7342);
or U8253 (N_8253,N_7178,N_4468);
or U8254 (N_8254,N_5462,N_5466);
nor U8255 (N_8255,N_7718,N_4779);
nor U8256 (N_8256,N_6449,N_4635);
nor U8257 (N_8257,N_6751,N_5616);
nor U8258 (N_8258,N_7662,N_5505);
nand U8259 (N_8259,N_7633,N_7455);
nor U8260 (N_8260,N_7546,N_4177);
nand U8261 (N_8261,N_7737,N_4188);
nand U8262 (N_8262,N_7810,N_6007);
or U8263 (N_8263,N_4370,N_7017);
nand U8264 (N_8264,N_5442,N_6934);
nor U8265 (N_8265,N_6656,N_4184);
nor U8266 (N_8266,N_7722,N_6753);
xnor U8267 (N_8267,N_4760,N_5681);
nor U8268 (N_8268,N_7750,N_7796);
nand U8269 (N_8269,N_6519,N_4986);
or U8270 (N_8270,N_5608,N_5418);
or U8271 (N_8271,N_5408,N_6336);
nand U8272 (N_8272,N_4294,N_4817);
or U8273 (N_8273,N_4908,N_7027);
nand U8274 (N_8274,N_4598,N_7551);
and U8275 (N_8275,N_5046,N_4965);
and U8276 (N_8276,N_7606,N_5398);
nand U8277 (N_8277,N_5210,N_5870);
and U8278 (N_8278,N_4860,N_5377);
nand U8279 (N_8279,N_6231,N_6788);
nand U8280 (N_8280,N_4265,N_5140);
or U8281 (N_8281,N_7849,N_5290);
and U8282 (N_8282,N_6759,N_4152);
or U8283 (N_8283,N_4398,N_7066);
nand U8284 (N_8284,N_7381,N_5272);
nor U8285 (N_8285,N_7130,N_6897);
xnor U8286 (N_8286,N_4832,N_5746);
and U8287 (N_8287,N_4024,N_5697);
or U8288 (N_8288,N_7900,N_4933);
and U8289 (N_8289,N_4160,N_6133);
and U8290 (N_8290,N_6855,N_5880);
nand U8291 (N_8291,N_7371,N_4982);
nand U8292 (N_8292,N_6987,N_6570);
and U8293 (N_8293,N_7126,N_7841);
or U8294 (N_8294,N_7727,N_4660);
and U8295 (N_8295,N_4937,N_7046);
nor U8296 (N_8296,N_7099,N_4776);
or U8297 (N_8297,N_6302,N_6578);
and U8298 (N_8298,N_7918,N_4677);
nand U8299 (N_8299,N_6171,N_5103);
and U8300 (N_8300,N_7090,N_4820);
nor U8301 (N_8301,N_6576,N_5672);
or U8302 (N_8302,N_6550,N_5864);
nand U8303 (N_8303,N_6555,N_5555);
nor U8304 (N_8304,N_7873,N_7236);
nand U8305 (N_8305,N_6654,N_5361);
and U8306 (N_8306,N_7528,N_6509);
nor U8307 (N_8307,N_7815,N_5463);
nor U8308 (N_8308,N_7015,N_7715);
or U8309 (N_8309,N_6472,N_5552);
or U8310 (N_8310,N_5100,N_5396);
nand U8311 (N_8311,N_6649,N_5892);
nand U8312 (N_8312,N_5072,N_5208);
nand U8313 (N_8313,N_4278,N_4590);
nand U8314 (N_8314,N_6343,N_5869);
or U8315 (N_8315,N_7225,N_4214);
or U8316 (N_8316,N_7949,N_7284);
or U8317 (N_8317,N_5483,N_6684);
or U8318 (N_8318,N_6541,N_4601);
nor U8319 (N_8319,N_6950,N_4475);
or U8320 (N_8320,N_5399,N_4504);
nand U8321 (N_8321,N_5528,N_5323);
and U8322 (N_8322,N_6580,N_7092);
or U8323 (N_8323,N_7624,N_5612);
nor U8324 (N_8324,N_6630,N_7503);
nand U8325 (N_8325,N_6109,N_4951);
or U8326 (N_8326,N_6369,N_6426);
or U8327 (N_8327,N_5359,N_5651);
xnor U8328 (N_8328,N_6423,N_7720);
nand U8329 (N_8329,N_7723,N_4268);
or U8330 (N_8330,N_5271,N_4926);
nand U8331 (N_8331,N_4205,N_4169);
and U8332 (N_8332,N_5756,N_6079);
and U8333 (N_8333,N_6977,N_6244);
or U8334 (N_8334,N_5731,N_4652);
or U8335 (N_8335,N_4793,N_6249);
nor U8336 (N_8336,N_7186,N_6096);
or U8337 (N_8337,N_4159,N_7508);
nor U8338 (N_8338,N_7257,N_5030);
nor U8339 (N_8339,N_7054,N_7158);
or U8340 (N_8340,N_5840,N_4227);
and U8341 (N_8341,N_6365,N_4838);
and U8342 (N_8342,N_7454,N_4383);
nor U8343 (N_8343,N_4544,N_7809);
and U8344 (N_8344,N_5856,N_4474);
or U8345 (N_8345,N_6257,N_6045);
or U8346 (N_8346,N_5784,N_7958);
xor U8347 (N_8347,N_7402,N_4004);
nand U8348 (N_8348,N_7278,N_6996);
nand U8349 (N_8349,N_6300,N_5258);
nand U8350 (N_8350,N_4105,N_6616);
nand U8351 (N_8351,N_6584,N_7067);
nand U8352 (N_8352,N_4441,N_4286);
nor U8353 (N_8353,N_6766,N_6883);
nor U8354 (N_8354,N_4453,N_7322);
or U8355 (N_8355,N_7170,N_6985);
and U8356 (N_8356,N_4546,N_7347);
nor U8357 (N_8357,N_6317,N_7056);
nand U8358 (N_8358,N_4647,N_5706);
and U8359 (N_8359,N_7372,N_5010);
or U8360 (N_8360,N_5356,N_5637);
and U8361 (N_8361,N_6383,N_4566);
nor U8362 (N_8362,N_5236,N_5913);
nand U8363 (N_8363,N_4613,N_6039);
or U8364 (N_8364,N_5488,N_7518);
and U8365 (N_8365,N_7083,N_7318);
nand U8366 (N_8366,N_6280,N_5871);
and U8367 (N_8367,N_7730,N_5144);
or U8368 (N_8368,N_5684,N_5139);
nand U8369 (N_8369,N_6959,N_4442);
or U8370 (N_8370,N_4514,N_5047);
nand U8371 (N_8371,N_5500,N_6691);
or U8372 (N_8372,N_6088,N_5482);
xor U8373 (N_8373,N_7562,N_5591);
nand U8374 (N_8374,N_4394,N_4056);
and U8375 (N_8375,N_5226,N_6810);
and U8376 (N_8376,N_4444,N_4762);
and U8377 (N_8377,N_5265,N_5534);
nand U8378 (N_8378,N_4427,N_6430);
and U8379 (N_8379,N_5286,N_4358);
nand U8380 (N_8380,N_4097,N_6483);
nor U8381 (N_8381,N_6152,N_4591);
nor U8382 (N_8382,N_4554,N_6839);
nor U8383 (N_8383,N_7558,N_4509);
nand U8384 (N_8384,N_7206,N_5866);
nand U8385 (N_8385,N_5387,N_4198);
nand U8386 (N_8386,N_7657,N_5661);
or U8387 (N_8387,N_7324,N_5508);
nand U8388 (N_8388,N_6310,N_6868);
nand U8389 (N_8389,N_4967,N_7210);
or U8390 (N_8390,N_4106,N_5969);
nand U8391 (N_8391,N_7860,N_6377);
nor U8392 (N_8392,N_7147,N_6169);
nor U8393 (N_8393,N_4599,N_5506);
nor U8394 (N_8394,N_4496,N_7184);
and U8395 (N_8395,N_4109,N_5717);
or U8396 (N_8396,N_5390,N_4176);
nor U8397 (N_8397,N_6886,N_5538);
and U8398 (N_8398,N_5879,N_4958);
nor U8399 (N_8399,N_6237,N_4446);
or U8400 (N_8400,N_4050,N_6814);
and U8401 (N_8401,N_6411,N_7391);
and U8402 (N_8402,N_5082,N_4791);
or U8403 (N_8403,N_4941,N_6227);
nand U8404 (N_8404,N_5544,N_5097);
nand U8405 (N_8405,N_5433,N_5926);
xor U8406 (N_8406,N_5908,N_4212);
and U8407 (N_8407,N_6037,N_5794);
or U8408 (N_8408,N_5026,N_6617);
and U8409 (N_8409,N_7930,N_6757);
nor U8410 (N_8410,N_6046,N_6626);
xnor U8411 (N_8411,N_7179,N_6796);
and U8412 (N_8412,N_6635,N_4082);
nor U8413 (N_8413,N_6873,N_7758);
or U8414 (N_8414,N_5450,N_4737);
and U8415 (N_8415,N_4440,N_4459);
nand U8416 (N_8416,N_4257,N_7753);
nor U8417 (N_8417,N_4490,N_4856);
and U8418 (N_8418,N_4100,N_4869);
nand U8419 (N_8419,N_6998,N_4824);
nand U8420 (N_8420,N_4017,N_4074);
and U8421 (N_8421,N_5549,N_7837);
nor U8422 (N_8422,N_7668,N_7002);
and U8423 (N_8423,N_5388,N_7133);
or U8424 (N_8424,N_7907,N_5863);
or U8425 (N_8425,N_6727,N_4654);
and U8426 (N_8426,N_5623,N_6515);
nor U8427 (N_8427,N_5475,N_4139);
nor U8428 (N_8428,N_7261,N_6148);
and U8429 (N_8429,N_7615,N_5602);
nor U8430 (N_8430,N_7336,N_4841);
nand U8431 (N_8431,N_5922,N_5788);
and U8432 (N_8432,N_4645,N_4571);
nor U8433 (N_8433,N_4743,N_6205);
nand U8434 (N_8434,N_4234,N_6156);
nand U8435 (N_8435,N_5927,N_5247);
nor U8436 (N_8436,N_6333,N_6979);
nand U8437 (N_8437,N_7640,N_4002);
nor U8438 (N_8438,N_4748,N_6147);
nor U8439 (N_8439,N_6204,N_7834);
nand U8440 (N_8440,N_7375,N_7913);
or U8441 (N_8441,N_4630,N_7507);
nand U8442 (N_8442,N_7116,N_5293);
nand U8443 (N_8443,N_6480,N_5197);
nand U8444 (N_8444,N_5639,N_6802);
or U8445 (N_8445,N_5547,N_6971);
nor U8446 (N_8446,N_5243,N_5426);
and U8447 (N_8447,N_4270,N_5031);
nor U8448 (N_8448,N_4646,N_4818);
nand U8449 (N_8449,N_7772,N_5749);
nor U8450 (N_8450,N_4364,N_4189);
or U8451 (N_8451,N_4576,N_5662);
nand U8452 (N_8452,N_7195,N_5045);
and U8453 (N_8453,N_7408,N_5460);
nor U8454 (N_8454,N_6922,N_7622);
nor U8455 (N_8455,N_4804,N_5157);
and U8456 (N_8456,N_4957,N_4085);
and U8457 (N_8457,N_7916,N_5594);
nand U8458 (N_8458,N_6706,N_4485);
and U8459 (N_8459,N_6619,N_6236);
or U8460 (N_8460,N_6723,N_7577);
or U8461 (N_8461,N_4470,N_4615);
and U8462 (N_8462,N_6748,N_7379);
and U8463 (N_8463,N_7742,N_6755);
nor U8464 (N_8464,N_7495,N_6197);
or U8465 (N_8465,N_5069,N_5890);
nor U8466 (N_8466,N_6381,N_5940);
nor U8467 (N_8467,N_5317,N_5274);
and U8468 (N_8468,N_7923,N_5750);
or U8469 (N_8469,N_6041,N_7249);
and U8470 (N_8470,N_7159,N_6542);
or U8471 (N_8471,N_4404,N_7071);
nor U8472 (N_8472,N_6022,N_4088);
nor U8473 (N_8473,N_7951,N_7706);
or U8474 (N_8474,N_7952,N_6914);
nand U8475 (N_8475,N_5123,N_6513);
and U8476 (N_8476,N_7755,N_6190);
and U8477 (N_8477,N_5134,N_5704);
nand U8478 (N_8478,N_7018,N_4801);
nor U8479 (N_8479,N_5527,N_7049);
nor U8480 (N_8480,N_4990,N_6604);
nand U8481 (N_8481,N_7434,N_5955);
nor U8482 (N_8482,N_4678,N_5105);
nor U8483 (N_8483,N_5563,N_7997);
nor U8484 (N_8484,N_5667,N_6173);
nor U8485 (N_8485,N_7986,N_5086);
and U8486 (N_8486,N_5194,N_7807);
nor U8487 (N_8487,N_4889,N_5231);
and U8488 (N_8488,N_5409,N_4772);
nand U8489 (N_8489,N_4559,N_6507);
or U8490 (N_8490,N_6895,N_4430);
or U8491 (N_8491,N_4309,N_7741);
nor U8492 (N_8492,N_7486,N_7693);
xnor U8493 (N_8493,N_5934,N_7139);
nor U8494 (N_8494,N_4536,N_4478);
and U8495 (N_8495,N_5655,N_4319);
nand U8496 (N_8496,N_4771,N_5303);
nor U8497 (N_8497,N_5122,N_7514);
nor U8498 (N_8498,N_6732,N_7665);
or U8499 (N_8499,N_5013,N_5486);
and U8500 (N_8500,N_4526,N_4421);
nand U8501 (N_8501,N_4825,N_4715);
or U8502 (N_8502,N_6246,N_7506);
nand U8503 (N_8503,N_5137,N_4185);
or U8504 (N_8504,N_6438,N_6132);
nor U8505 (N_8505,N_6948,N_5410);
or U8506 (N_8506,N_5102,N_5504);
nor U8507 (N_8507,N_4498,N_4053);
or U8508 (N_8508,N_7448,N_4756);
or U8509 (N_8509,N_6024,N_7927);
nand U8510 (N_8510,N_5485,N_5687);
nor U8511 (N_8511,N_7275,N_5446);
or U8512 (N_8512,N_5541,N_5949);
or U8513 (N_8513,N_5991,N_6367);
and U8514 (N_8514,N_7452,N_4850);
or U8515 (N_8515,N_7216,N_6482);
nand U8516 (N_8516,N_4166,N_7237);
nor U8517 (N_8517,N_6400,N_5730);
nand U8518 (N_8518,N_4277,N_6463);
or U8519 (N_8519,N_6716,N_7101);
or U8520 (N_8520,N_7512,N_5903);
nor U8521 (N_8521,N_6587,N_5718);
or U8522 (N_8522,N_7374,N_7413);
and U8523 (N_8523,N_7244,N_4697);
nor U8524 (N_8524,N_6072,N_5330);
or U8525 (N_8525,N_4323,N_6880);
nor U8526 (N_8526,N_6005,N_6413);
or U8527 (N_8527,N_7821,N_7243);
nor U8528 (N_8528,N_4578,N_5834);
and U8529 (N_8529,N_5381,N_7903);
nand U8530 (N_8530,N_4326,N_4351);
nand U8531 (N_8531,N_4714,N_7369);
nand U8532 (N_8532,N_7479,N_4325);
and U8533 (N_8533,N_4147,N_4930);
and U8534 (N_8534,N_4473,N_7387);
xor U8535 (N_8535,N_6230,N_6731);
or U8536 (N_8536,N_5842,N_5715);
xor U8537 (N_8537,N_5130,N_6481);
or U8538 (N_8538,N_7467,N_7108);
and U8539 (N_8539,N_4669,N_4521);
nand U8540 (N_8540,N_5148,N_7203);
and U8541 (N_8541,N_5407,N_5000);
nor U8542 (N_8542,N_7441,N_6908);
and U8543 (N_8543,N_7282,N_5191);
and U8544 (N_8544,N_6864,N_6910);
and U8545 (N_8545,N_5575,N_6990);
and U8546 (N_8546,N_4740,N_5028);
nand U8547 (N_8547,N_6629,N_4668);
nand U8548 (N_8548,N_4734,N_6544);
or U8549 (N_8549,N_6842,N_4095);
nand U8550 (N_8550,N_6678,N_4847);
nand U8551 (N_8551,N_5511,N_5822);
xor U8552 (N_8552,N_4923,N_6981);
and U8553 (N_8553,N_5115,N_5057);
or U8554 (N_8554,N_5688,N_5386);
or U8555 (N_8555,N_6451,N_6239);
or U8556 (N_8556,N_7626,N_7880);
or U8557 (N_8557,N_7306,N_7928);
or U8558 (N_8558,N_7129,N_4254);
nor U8559 (N_8559,N_6409,N_4584);
or U8560 (N_8560,N_6308,N_7259);
or U8561 (N_8561,N_6391,N_6915);
nor U8562 (N_8562,N_7045,N_4494);
nor U8563 (N_8563,N_7544,N_7326);
nand U8564 (N_8564,N_4118,N_7780);
and U8565 (N_8565,N_7650,N_7319);
nor U8566 (N_8566,N_5368,N_4903);
nand U8567 (N_8567,N_4658,N_4907);
nand U8568 (N_8568,N_5024,N_5339);
nor U8569 (N_8569,N_7462,N_4400);
or U8570 (N_8570,N_7480,N_6980);
or U8571 (N_8571,N_4233,N_6077);
nand U8572 (N_8572,N_4343,N_7235);
xnor U8573 (N_8573,N_4489,N_7102);
nand U8574 (N_8574,N_7478,N_7666);
nor U8575 (N_8575,N_7517,N_7743);
and U8576 (N_8576,N_5402,N_6663);
and U8577 (N_8577,N_7305,N_7211);
nand U8578 (N_8578,N_7255,N_5867);
nor U8579 (N_8579,N_4471,N_6264);
xor U8580 (N_8580,N_4653,N_4642);
and U8581 (N_8581,N_6878,N_5557);
or U8582 (N_8582,N_7857,N_7078);
nand U8583 (N_8583,N_5984,N_5957);
nor U8584 (N_8584,N_5347,N_4300);
or U8585 (N_8585,N_6650,N_5478);
and U8586 (N_8586,N_7414,N_6083);
nor U8587 (N_8587,N_4777,N_7404);
nor U8588 (N_8588,N_6911,N_4745);
and U8589 (N_8589,N_6454,N_5307);
and U8590 (N_8590,N_7224,N_5771);
or U8591 (N_8591,N_7521,N_7912);
nor U8592 (N_8592,N_7614,N_5657);
or U8593 (N_8593,N_5675,N_5065);
and U8594 (N_8594,N_4260,N_6125);
nand U8595 (N_8595,N_4572,N_5607);
nand U8596 (N_8596,N_6898,N_5354);
nand U8597 (N_8597,N_7010,N_4307);
and U8598 (N_8598,N_6315,N_4983);
nor U8599 (N_8599,N_5423,N_7198);
or U8600 (N_8600,N_5811,N_5752);
and U8601 (N_8601,N_4575,N_7199);
xnor U8602 (N_8602,N_7604,N_7122);
or U8603 (N_8603,N_7185,N_5033);
xor U8604 (N_8604,N_6540,N_7153);
nand U8605 (N_8605,N_5479,N_6462);
nor U8606 (N_8606,N_5519,N_5588);
nor U8607 (N_8607,N_7713,N_4788);
nor U8608 (N_8608,N_4414,N_4086);
and U8609 (N_8609,N_4000,N_6004);
nand U8610 (N_8610,N_6141,N_4969);
nand U8611 (N_8611,N_4659,N_7309);
or U8612 (N_8612,N_7453,N_7762);
and U8613 (N_8613,N_6809,N_5152);
nor U8614 (N_8614,N_4037,N_6025);
or U8615 (N_8615,N_7157,N_7327);
nand U8616 (N_8616,N_7909,N_5133);
nor U8617 (N_8617,N_5945,N_4092);
and U8618 (N_8618,N_5994,N_6060);
or U8619 (N_8619,N_7373,N_6565);
or U8620 (N_8620,N_5251,N_6091);
or U8621 (N_8621,N_7915,N_5084);
nand U8622 (N_8622,N_7472,N_7424);
nand U8623 (N_8623,N_4464,N_4014);
nand U8624 (N_8624,N_5343,N_4707);
and U8625 (N_8625,N_4055,N_6305);
and U8626 (N_8626,N_4289,N_6347);
nand U8627 (N_8627,N_6567,N_7717);
xnor U8628 (N_8628,N_7035,N_4640);
nand U8629 (N_8629,N_7616,N_4425);
or U8630 (N_8630,N_7189,N_5195);
nor U8631 (N_8631,N_6687,N_4588);
and U8632 (N_8632,N_5099,N_4894);
nor U8633 (N_8633,N_6306,N_7968);
nor U8634 (N_8634,N_5472,N_5783);
nand U8635 (N_8635,N_6421,N_6714);
or U8636 (N_8636,N_6180,N_5393);
or U8637 (N_8637,N_7201,N_4158);
nor U8638 (N_8638,N_7596,N_5114);
nor U8639 (N_8639,N_5539,N_6099);
nand U8640 (N_8640,N_4486,N_4331);
nand U8641 (N_8641,N_4493,N_7048);
or U8642 (N_8642,N_4413,N_7822);
and U8643 (N_8643,N_7525,N_7355);
nor U8644 (N_8644,N_6089,N_6348);
nor U8645 (N_8645,N_5650,N_7197);
or U8646 (N_8646,N_6964,N_4711);
and U8647 (N_8647,N_6813,N_7566);
nor U8648 (N_8648,N_7987,N_6304);
xor U8649 (N_8649,N_4831,N_7338);
and U8650 (N_8650,N_4597,N_5736);
or U8651 (N_8651,N_4633,N_6527);
nor U8652 (N_8652,N_6583,N_5848);
and U8653 (N_8653,N_7778,N_4780);
nand U8654 (N_8654,N_6798,N_6207);
and U8655 (N_8655,N_4732,N_7765);
or U8656 (N_8656,N_4622,N_4700);
and U8657 (N_8657,N_4950,N_5853);
nor U8658 (N_8658,N_5668,N_4324);
nand U8659 (N_8659,N_5235,N_4310);
xnor U8660 (N_8660,N_5219,N_7358);
or U8661 (N_8661,N_6960,N_6906);
nand U8662 (N_8662,N_5825,N_6644);
or U8663 (N_8663,N_5696,N_6076);
nor U8664 (N_8664,N_5135,N_4318);
or U8665 (N_8665,N_7538,N_6081);
and U8666 (N_8666,N_6313,N_6636);
or U8667 (N_8667,N_4040,N_6708);
or U8668 (N_8668,N_4094,N_7132);
and U8669 (N_8669,N_7697,N_7095);
and U8670 (N_8670,N_4103,N_4871);
or U8671 (N_8671,N_5253,N_6894);
or U8672 (N_8672,N_7466,N_4542);
and U8673 (N_8673,N_7999,N_6176);
nand U8674 (N_8674,N_4381,N_4462);
and U8675 (N_8675,N_6496,N_4993);
nand U8676 (N_8676,N_4944,N_7220);
nor U8677 (N_8677,N_5440,N_6784);
nand U8678 (N_8678,N_5664,N_5413);
and U8679 (N_8679,N_4482,N_6742);
or U8680 (N_8680,N_5342,N_5790);
or U8681 (N_8681,N_5039,N_7625);
nor U8682 (N_8682,N_6201,N_7475);
or U8683 (N_8683,N_4798,N_4781);
nand U8684 (N_8684,N_4228,N_5520);
nand U8685 (N_8685,N_7838,N_7811);
xor U8686 (N_8686,N_4349,N_6647);
nor U8687 (N_8687,N_5606,N_6641);
and U8688 (N_8688,N_4506,N_4736);
nand U8689 (N_8689,N_4267,N_6155);
and U8690 (N_8690,N_6274,N_4239);
xor U8691 (N_8691,N_4330,N_4365);
nor U8692 (N_8692,N_4125,N_6247);
and U8693 (N_8693,N_7232,N_5565);
or U8694 (N_8694,N_5020,N_5392);
nor U8695 (N_8695,N_4312,N_4202);
nand U8696 (N_8696,N_5094,N_6445);
nand U8697 (N_8697,N_4354,N_6172);
or U8698 (N_8698,N_4116,N_6696);
nand U8699 (N_8699,N_7797,N_7473);
or U8700 (N_8700,N_5857,N_6547);
nand U8701 (N_8701,N_7144,N_5659);
and U8702 (N_8702,N_5509,N_6820);
and U8703 (N_8703,N_5819,N_6221);
nor U8704 (N_8704,N_5230,N_6611);
nand U8705 (N_8705,N_6049,N_5620);
nand U8706 (N_8706,N_7395,N_5562);
xnor U8707 (N_8707,N_7794,N_7269);
and U8708 (N_8708,N_7960,N_6733);
and U8709 (N_8709,N_5222,N_4380);
nand U8710 (N_8710,N_7899,N_6568);
nand U8711 (N_8711,N_4311,N_7003);
and U8712 (N_8712,N_4962,N_6847);
nor U8713 (N_8713,N_6932,N_5111);
or U8714 (N_8714,N_4592,N_6021);
nor U8715 (N_8715,N_7292,N_6488);
nor U8716 (N_8716,N_4858,N_6399);
and U8717 (N_8717,N_7569,N_6586);
nor U8718 (N_8718,N_6354,N_6564);
and U8719 (N_8719,N_7866,N_5974);
and U8720 (N_8720,N_5032,N_7840);
and U8721 (N_8721,N_5535,N_6440);
nand U8722 (N_8722,N_4783,N_7264);
xnor U8723 (N_8723,N_7166,N_6780);
nand U8724 (N_8724,N_5928,N_6033);
or U8725 (N_8725,N_7635,N_6828);
and U8726 (N_8726,N_7587,N_4988);
or U8727 (N_8727,N_5944,N_7376);
and U8728 (N_8728,N_5907,N_5119);
nor U8729 (N_8729,N_4656,N_6129);
nor U8730 (N_8730,N_4706,N_6836);
nand U8731 (N_8731,N_5861,N_5277);
and U8732 (N_8732,N_5690,N_4367);
or U8733 (N_8733,N_5893,N_5149);
and U8734 (N_8734,N_5206,N_7594);
or U8735 (N_8735,N_6285,N_4350);
nor U8736 (N_8736,N_5986,N_5431);
nand U8737 (N_8737,N_6879,N_4436);
or U8738 (N_8738,N_6321,N_5034);
nand U8739 (N_8739,N_6832,N_4855);
nor U8740 (N_8740,N_6210,N_7105);
nand U8741 (N_8741,N_7738,N_7001);
nor U8742 (N_8742,N_6791,N_7082);
and U8743 (N_8743,N_6750,N_7077);
or U8744 (N_8744,N_4195,N_7819);
and U8745 (N_8745,N_4693,N_6182);
nor U8746 (N_8746,N_6177,N_7876);
nor U8747 (N_8747,N_4376,N_4244);
nor U8748 (N_8748,N_4805,N_5281);
and U8749 (N_8749,N_4028,N_6402);
and U8750 (N_8750,N_7394,N_6673);
nor U8751 (N_8751,N_7729,N_4870);
or U8752 (N_8752,N_4199,N_7831);
and U8753 (N_8753,N_4066,N_6162);
or U8754 (N_8754,N_4469,N_5685);
or U8755 (N_8755,N_5753,N_4126);
or U8756 (N_8756,N_6642,N_4523);
nor U8757 (N_8757,N_6638,N_5495);
and U8758 (N_8758,N_4991,N_4359);
nor U8759 (N_8759,N_5417,N_6887);
and U8760 (N_8760,N_5378,N_5533);
nand U8761 (N_8761,N_6503,N_7393);
nor U8762 (N_8762,N_5897,N_7739);
or U8763 (N_8763,N_6846,N_7352);
nor U8764 (N_8764,N_5510,N_4333);
and U8765 (N_8765,N_7933,N_5054);
and U8766 (N_8766,N_4596,N_7590);
nand U8767 (N_8767,N_6120,N_7591);
nand U8768 (N_8768,N_7629,N_6329);
xor U8769 (N_8769,N_5349,N_6145);
and U8770 (N_8770,N_4104,N_6395);
or U8771 (N_8771,N_6050,N_6394);
nand U8772 (N_8772,N_6634,N_6150);
nor U8773 (N_8773,N_6209,N_6817);
nor U8774 (N_8774,N_4569,N_7982);
nand U8775 (N_8775,N_4690,N_7247);
nor U8776 (N_8776,N_6455,N_6026);
and U8777 (N_8777,N_7403,N_5778);
nor U8778 (N_8778,N_5451,N_4973);
and U8779 (N_8779,N_4587,N_4296);
and U8780 (N_8780,N_4463,N_6139);
or U8781 (N_8781,N_7516,N_4075);
nand U8782 (N_8782,N_5420,N_5767);
nor U8783 (N_8783,N_5239,N_7683);
or U8784 (N_8784,N_6861,N_5193);
nor U8785 (N_8785,N_5077,N_7712);
and U8786 (N_8786,N_5985,N_4488);
nor U8787 (N_8787,N_7134,N_7142);
or U8788 (N_8788,N_5002,N_5909);
and U8789 (N_8789,N_7721,N_5331);
and U8790 (N_8790,N_4492,N_4619);
or U8791 (N_8791,N_5404,N_5300);
and U8792 (N_8792,N_5751,N_5693);
nand U8793 (N_8793,N_6396,N_4522);
nand U8794 (N_8794,N_5593,N_6937);
nor U8795 (N_8795,N_6728,N_6116);
nand U8796 (N_8796,N_4043,N_6537);
nor U8797 (N_8797,N_4012,N_6514);
and U8798 (N_8798,N_6961,N_6157);
and U8799 (N_8799,N_7911,N_4874);
and U8800 (N_8800,N_4443,N_6558);
nand U8801 (N_8801,N_4945,N_7346);
nand U8802 (N_8802,N_7681,N_7953);
or U8803 (N_8803,N_6484,N_4676);
nor U8804 (N_8804,N_6299,N_6052);
or U8805 (N_8805,N_4720,N_4410);
or U8806 (N_8806,N_5683,N_4124);
and U8807 (N_8807,N_6774,N_6610);
nor U8808 (N_8808,N_4687,N_4995);
nor U8809 (N_8809,N_5872,N_6467);
nand U8810 (N_8810,N_6592,N_4164);
nor U8811 (N_8811,N_7212,N_6625);
or U8812 (N_8812,N_5951,N_7962);
or U8813 (N_8813,N_6743,N_7846);
nand U8814 (N_8814,N_6951,N_6243);
or U8815 (N_8815,N_4899,N_6082);
or U8816 (N_8816,N_7023,N_6185);
nand U8817 (N_8817,N_5815,N_5891);
nor U8818 (N_8818,N_4823,N_7444);
and U8819 (N_8819,N_4977,N_6003);
nand U8820 (N_8820,N_7586,N_5828);
and U8821 (N_8821,N_7006,N_7274);
nor U8822 (N_8822,N_6375,N_5705);
nor U8823 (N_8823,N_5424,N_6530);
nand U8824 (N_8824,N_5873,N_4866);
nor U8825 (N_8825,N_5865,N_7143);
nand U8826 (N_8826,N_4251,N_5553);
nand U8827 (N_8827,N_4839,N_7628);
nor U8828 (N_8828,N_4213,N_5721);
or U8829 (N_8829,N_4857,N_7442);
and U8830 (N_8830,N_5843,N_5336);
and U8831 (N_8831,N_5048,N_6372);
and U8832 (N_8832,N_7709,N_5329);
nor U8833 (N_8833,N_7748,N_6871);
nor U8834 (N_8834,N_7680,N_6607);
nor U8835 (N_8835,N_6704,N_4843);
nand U8836 (N_8836,N_7692,N_5728);
and U8837 (N_8837,N_7151,N_5429);
nor U8838 (N_8838,N_6860,N_6353);
or U8839 (N_8839,N_5829,N_7788);
and U8840 (N_8840,N_6303,N_6078);
or U8841 (N_8841,N_5876,N_5712);
and U8842 (N_8842,N_5477,N_7345);
or U8843 (N_8843,N_6772,N_4063);
or U8844 (N_8844,N_4609,N_4438);
nor U8845 (N_8845,N_7180,N_4961);
nand U8846 (N_8846,N_7839,N_7993);
nor U8847 (N_8847,N_5108,N_6856);
and U8848 (N_8848,N_6675,N_5207);
or U8849 (N_8849,N_5205,N_6464);
nand U8850 (N_8850,N_5470,N_4090);
nand U8851 (N_8851,N_4081,N_5905);
and U8852 (N_8852,N_6941,N_4279);
nor U8853 (N_8853,N_4390,N_7019);
nor U8854 (N_8854,N_7025,N_7728);
nand U8855 (N_8855,N_5040,N_7285);
nor U8856 (N_8856,N_5773,N_5345);
nand U8857 (N_8857,N_7805,N_4864);
or U8858 (N_8858,N_5252,N_7574);
nand U8859 (N_8859,N_6797,N_4834);
and U8860 (N_8860,N_4698,N_5276);
nor U8861 (N_8861,N_5249,N_6330);
nand U8862 (N_8862,N_7174,N_5147);
or U8863 (N_8863,N_7488,N_4786);
nand U8864 (N_8864,N_4796,N_7656);
nor U8865 (N_8865,N_6397,N_4694);
nor U8866 (N_8866,N_6923,N_5716);
and U8867 (N_8867,N_5295,N_4457);
and U8868 (N_8868,N_4769,N_6422);
and U8869 (N_8869,N_5405,N_5670);
nor U8870 (N_8870,N_6268,N_5383);
nor U8871 (N_8871,N_6840,N_4766);
and U8872 (N_8872,N_5406,N_6874);
nand U8873 (N_8873,N_7103,N_5464);
nand U8874 (N_8874,N_5582,N_4203);
or U8875 (N_8875,N_5452,N_7564);
and U8876 (N_8876,N_6787,N_4298);
or U8877 (N_8877,N_4355,N_4761);
nor U8878 (N_8878,N_7213,N_7074);
nand U8879 (N_8879,N_7125,N_7233);
nand U8880 (N_8880,N_5646,N_5200);
or U8881 (N_8881,N_7917,N_4230);
nor U8882 (N_8882,N_6008,N_7493);
nor U8883 (N_8883,N_5209,N_6548);
nand U8884 (N_8884,N_6479,N_7024);
or U8885 (N_8885,N_6900,N_7008);
nor U8886 (N_8886,N_7904,N_5443);
nand U8887 (N_8887,N_6615,N_7886);
and U8888 (N_8888,N_7217,N_6485);
nor U8889 (N_8889,N_7530,N_4946);
nor U8890 (N_8890,N_7791,N_6863);
or U8891 (N_8891,N_6128,N_4890);
nand U8892 (N_8892,N_4271,N_6323);
nand U8893 (N_8893,N_4407,N_6944);
or U8894 (N_8894,N_6909,N_6165);
and U8895 (N_8895,N_6853,N_7965);
and U8896 (N_8896,N_4563,N_6251);
and U8897 (N_8897,N_4010,N_6848);
nor U8898 (N_8898,N_6457,N_6603);
or U8899 (N_8899,N_4285,N_5894);
and U8900 (N_8900,N_5958,N_6453);
nand U8901 (N_8901,N_7638,N_6633);
nor U8902 (N_8902,N_5225,N_7471);
nor U8903 (N_8903,N_7152,N_5344);
and U8904 (N_8904,N_4637,N_4175);
xnor U8905 (N_8905,N_6127,N_7191);
nand U8906 (N_8906,N_6707,N_4530);
and U8907 (N_8907,N_4980,N_4625);
and U8908 (N_8908,N_4001,N_5614);
nand U8909 (N_8909,N_5184,N_6953);
nor U8910 (N_8910,N_6976,N_7412);
nor U8911 (N_8911,N_7685,N_6328);
or U8912 (N_8912,N_7934,N_4258);
nor U8913 (N_8913,N_7975,N_4114);
or U8914 (N_8914,N_6135,N_5457);
and U8915 (N_8915,N_6854,N_5131);
and U8916 (N_8916,N_7851,N_5567);
and U8917 (N_8917,N_7332,N_4437);
nor U8918 (N_8918,N_6594,N_5297);
or U8919 (N_8919,N_7043,N_4369);
nand U8920 (N_8920,N_7937,N_6212);
nand U8921 (N_8921,N_5971,N_4332);
nand U8922 (N_8922,N_7784,N_7736);
nand U8923 (N_8923,N_6048,N_7925);
nor U8924 (N_8924,N_4282,N_6805);
nor U8925 (N_8925,N_6949,N_7883);
nand U8926 (N_8926,N_6334,N_5238);
nor U8927 (N_8927,N_7307,N_5881);
and U8928 (N_8928,N_5737,N_6441);
and U8929 (N_8929,N_7578,N_4674);
nor U8930 (N_8930,N_4211,N_5925);
and U8931 (N_8931,N_4555,N_4194);
or U8932 (N_8932,N_4445,N_5051);
nand U8933 (N_8933,N_7617,N_5921);
or U8934 (N_8934,N_7613,N_4272);
and U8935 (N_8935,N_5818,N_5839);
and U8936 (N_8936,N_5571,N_6528);
and U8937 (N_8937,N_6107,N_6739);
xnor U8938 (N_8938,N_5795,N_5542);
nor U8939 (N_8939,N_5525,N_7802);
or U8940 (N_8940,N_6031,N_5592);
nor U8941 (N_8941,N_6973,N_4744);
and U8942 (N_8942,N_6557,N_6764);
and U8943 (N_8943,N_4361,N_4840);
or U8944 (N_8944,N_5445,N_5076);
or U8945 (N_8945,N_5827,N_5515);
nand U8946 (N_8946,N_6137,N_7969);
nand U8947 (N_8947,N_5335,N_4371);
nand U8948 (N_8948,N_4940,N_7223);
and U8949 (N_8949,N_4755,N_5178);
and U8950 (N_8950,N_5658,N_6877);
nand U8951 (N_8951,N_7443,N_4865);
or U8952 (N_8952,N_6289,N_4960);
nand U8953 (N_8953,N_5568,N_4192);
nor U8954 (N_8954,N_7260,N_6153);
and U8955 (N_8955,N_5502,N_7344);
nand U8956 (N_8956,N_6414,N_5093);
and U8957 (N_8957,N_6042,N_6331);
or U8958 (N_8958,N_4998,N_4927);
or U8959 (N_8959,N_7808,N_7012);
nor U8960 (N_8960,N_5484,N_6420);
or U8961 (N_8961,N_4299,N_5022);
or U8962 (N_8962,N_4916,N_6401);
nor U8963 (N_8963,N_7176,N_7156);
or U8964 (N_8964,N_6154,N_6756);
nor U8965 (N_8965,N_5379,N_4460);
and U8966 (N_8966,N_6408,N_5145);
nand U8967 (N_8967,N_7052,N_6831);
nand U8968 (N_8968,N_4529,N_4648);
nand U8969 (N_8969,N_6931,N_4339);
and U8970 (N_8970,N_7754,N_5786);
or U8971 (N_8971,N_4295,N_5768);
and U8972 (N_8972,N_6560,N_4675);
nor U8973 (N_8973,N_6332,N_7337);
and U8974 (N_8974,N_7298,N_6602);
nand U8975 (N_8975,N_7539,N_5302);
or U8976 (N_8976,N_6815,N_5217);
and U8977 (N_8977,N_4867,N_5601);
or U8978 (N_8978,N_5216,N_7527);
nor U8979 (N_8979,N_5636,N_6778);
or U8980 (N_8980,N_5888,N_7330);
nand U8981 (N_8981,N_4898,N_6418);
or U8982 (N_8982,N_7816,N_4503);
and U8983 (N_8983,N_6341,N_7420);
or U8984 (N_8984,N_5234,N_4182);
and U8985 (N_8985,N_6254,N_5814);
nor U8986 (N_8986,N_4346,N_6986);
or U8987 (N_8987,N_5314,N_5761);
nand U8988 (N_8988,N_7795,N_7118);
nor U8989 (N_8989,N_4153,N_7970);
nor U8990 (N_8990,N_5953,N_6763);
or U8991 (N_8991,N_6677,N_7609);
nor U8992 (N_8992,N_7812,N_5680);
nand U8993 (N_8993,N_6581,N_7291);
or U8994 (N_8994,N_6556,N_4181);
and U8995 (N_8995,N_5649,N_4276);
and U8996 (N_8996,N_4641,N_4705);
nor U8997 (N_8997,N_5454,N_4938);
and U8998 (N_8998,N_5597,N_5758);
nor U8999 (N_8999,N_6845,N_4422);
and U9000 (N_9000,N_7310,N_6235);
and U9001 (N_9001,N_5996,N_4634);
nand U9002 (N_9002,N_5647,N_6378);
nor U9003 (N_9003,N_7759,N_6019);
and U9004 (N_9004,N_6066,N_5512);
nand U9005 (N_9005,N_7924,N_5240);
nor U9006 (N_9006,N_6387,N_6808);
or U9007 (N_9007,N_5807,N_7589);
or U9008 (N_9008,N_5177,N_5183);
xnor U9009 (N_9009,N_5067,N_5989);
nor U9010 (N_9010,N_6094,N_5228);
nand U9011 (N_9011,N_4638,N_6433);
and U9012 (N_9012,N_4815,N_5315);
nor U9013 (N_9013,N_7789,N_6522);
or U9014 (N_9014,N_6940,N_5150);
nand U9015 (N_9015,N_6737,N_7661);
nand U9016 (N_9016,N_5071,N_7265);
and U9017 (N_9017,N_4876,N_7906);
nor U9018 (N_9018,N_7155,N_4686);
xor U9019 (N_9019,N_4845,N_5306);
nand U9020 (N_9020,N_7221,N_5064);
or U9021 (N_9021,N_7929,N_6893);
nand U9022 (N_9022,N_5367,N_5029);
nor U9023 (N_9023,N_7272,N_4093);
nor U9024 (N_9024,N_7450,N_5995);
nor U9025 (N_9025,N_7349,N_5710);
nor U9026 (N_9026,N_7537,N_6623);
and U9027 (N_9027,N_6357,N_4165);
xnor U9028 (N_9028,N_6248,N_4250);
and U9029 (N_9029,N_6298,N_5261);
or U9030 (N_9030,N_6439,N_7914);
or U9031 (N_9031,N_4925,N_5632);
or U9032 (N_9032,N_5860,N_7483);
or U9033 (N_9033,N_7761,N_5066);
and U9034 (N_9034,N_6256,N_5411);
and U9035 (N_9035,N_5507,N_5800);
nand U9036 (N_9036,N_7552,N_7559);
and U9037 (N_9037,N_6632,N_7489);
and U9038 (N_9038,N_5545,N_7321);
nand U9039 (N_9039,N_7109,N_6474);
nor U9040 (N_9040,N_4280,N_5628);
nand U9041 (N_9041,N_7663,N_4747);
and U9042 (N_9042,N_6111,N_6261);
nand U9043 (N_9043,N_6888,N_7058);
and U9044 (N_9044,N_4363,N_6773);
and U9045 (N_9045,N_4764,N_4345);
xor U9046 (N_9046,N_7263,N_4606);
or U9047 (N_9047,N_5609,N_5993);
nor U9048 (N_9048,N_5781,N_5494);
or U9049 (N_9049,N_7980,N_7465);
nand U9050 (N_9050,N_4297,N_4757);
nand U9051 (N_9051,N_5966,N_7817);
or U9052 (N_9052,N_7733,N_6374);
and U9053 (N_9053,N_5109,N_6508);
nand U9054 (N_9054,N_7686,N_4378);
nor U9055 (N_9055,N_6339,N_7051);
nand U9056 (N_9056,N_4955,N_6966);
and U9057 (N_9057,N_4552,N_6628);
nor U9058 (N_9058,N_6754,N_5098);
nand U9059 (N_9059,N_6380,N_6722);
and U9060 (N_9060,N_4322,N_6090);
and U9061 (N_9061,N_6282,N_6792);
xor U9062 (N_9062,N_4084,N_6984);
nand U9063 (N_9063,N_7317,N_6667);
nor U9064 (N_9064,N_5287,N_7406);
nor U9065 (N_9065,N_7647,N_5107);
nor U9066 (N_9066,N_6875,N_7695);
nor U9067 (N_9067,N_7303,N_4208);
and U9068 (N_9068,N_5080,N_4020);
and U9069 (N_9069,N_7430,N_7477);
and U9070 (N_9070,N_7293,N_6777);
nor U9071 (N_9071,N_7026,N_7131);
nand U9072 (N_9072,N_4502,N_6803);
and U9073 (N_9073,N_4067,N_4665);
and U9074 (N_9074,N_5719,N_4848);
nor U9075 (N_9075,N_5011,N_4775);
nor U9076 (N_9076,N_6760,N_7121);
nor U9077 (N_9077,N_6067,N_7005);
or U9078 (N_9078,N_4275,N_6491);
and U9079 (N_9079,N_5845,N_6215);
and U9080 (N_9080,N_7832,N_4099);
nor U9081 (N_9081,N_5173,N_7435);
nor U9082 (N_9082,N_6849,N_6102);
nand U9083 (N_9083,N_5633,N_7234);
nand U9084 (N_9084,N_5155,N_6838);
nand U9085 (N_9085,N_4362,N_6672);
nor U9086 (N_9086,N_6071,N_6896);
nor U9087 (N_9087,N_6164,N_6912);
or U9088 (N_9088,N_7463,N_6730);
or U9089 (N_9089,N_4893,N_6882);
or U9090 (N_9090,N_4651,N_6539);
nor U9091 (N_9091,N_7716,N_6119);
nand U9092 (N_9092,N_7331,N_4417);
and U9093 (N_9093,N_6653,N_4009);
nand U9094 (N_9094,N_4352,N_5371);
nand U9095 (N_9095,N_4007,N_7304);
or U9096 (N_9096,N_4561,N_5255);
nand U9097 (N_9097,N_5775,N_5038);
or U9098 (N_9098,N_5596,N_7830);
nand U9099 (N_9099,N_4533,N_5682);
nor U9100 (N_9100,N_5319,N_7146);
xnor U9101 (N_9101,N_6040,N_5430);
or U9102 (N_9102,N_5316,N_5091);
nor U9103 (N_9103,N_6869,N_5006);
and U9104 (N_9104,N_6532,N_5419);
nand U9105 (N_9105,N_6114,N_4098);
and U9106 (N_9106,N_7557,N_7877);
and U9107 (N_9107,N_5403,N_7767);
nor U9108 (N_9108,N_7882,N_4681);
nand U9109 (N_9109,N_5179,N_4735);
or U9110 (N_9110,N_6233,N_6459);
or U9111 (N_9111,N_6097,N_4742);
nand U9112 (N_9112,N_4287,N_6149);
or U9113 (N_9113,N_5223,N_6032);
or U9114 (N_9114,N_6363,N_6804);
or U9115 (N_9115,N_5296,N_7300);
nor U9116 (N_9116,N_6920,N_4327);
and U9117 (N_9117,N_7165,N_5333);
nor U9118 (N_9118,N_7511,N_7963);
or U9119 (N_9119,N_6988,N_7173);
and U9120 (N_9120,N_6925,N_7214);
nand U9121 (N_9121,N_6789,N_7149);
and U9122 (N_9122,N_4547,N_4447);
or U9123 (N_9123,N_5902,N_5882);
and U9124 (N_9124,N_4305,N_7431);
or U9125 (N_9125,N_4829,N_4614);
nor U9126 (N_9126,N_7055,N_6370);
nand U9127 (N_9127,N_5652,N_4891);
nand U9128 (N_9128,N_4682,N_7764);
or U9129 (N_9129,N_7059,N_5036);
nor U9130 (N_9130,N_6705,N_7634);
nor U9131 (N_9131,N_4288,N_6865);
nor U9132 (N_9132,N_4595,N_5282);
nand U9133 (N_9133,N_5269,N_5898);
nor U9134 (N_9134,N_5923,N_4702);
nand U9135 (N_9135,N_5416,N_7704);
nand U9136 (N_9136,N_4612,N_4396);
and U9137 (N_9137,N_6417,N_6458);
or U9138 (N_9138,N_4389,N_5522);
nand U9139 (N_9139,N_7476,N_4347);
or U9140 (N_9140,N_4015,N_5062);
nand U9141 (N_9141,N_4044,N_4767);
nand U9142 (N_9142,N_7902,N_6811);
nor U9143 (N_9143,N_6267,N_5916);
and U9144 (N_9144,N_6559,N_4018);
nor U9145 (N_9145,N_7267,N_7995);
and U9146 (N_9146,N_5497,N_5625);
and U9147 (N_9147,N_7515,N_4065);
xor U9148 (N_9148,N_5885,N_6892);
or U9149 (N_9149,N_5666,N_6452);
and U9150 (N_9150,N_7757,N_6200);
nand U9151 (N_9151,N_7620,N_4814);
or U9152 (N_9152,N_6703,N_5154);
xor U9153 (N_9153,N_5166,N_6605);
nor U9154 (N_9154,N_5435,N_7627);
nor U9155 (N_9155,N_6446,N_6531);
nor U9156 (N_9156,N_6325,N_4204);
and U9157 (N_9157,N_7944,N_7534);
nand U9158 (N_9158,N_4628,N_6962);
or U9159 (N_9159,N_6525,N_4695);
or U9160 (N_9160,N_5931,N_6824);
or U9161 (N_9161,N_6228,N_4580);
or U9162 (N_9162,N_6058,N_6724);
and U9163 (N_9163,N_4191,N_5895);
and U9164 (N_9164,N_7744,N_4201);
or U9165 (N_9165,N_4906,N_5299);
and U9166 (N_9166,N_6245,N_7585);
nor U9167 (N_9167,N_7865,N_6098);
or U9168 (N_9168,N_4450,N_4629);
nor U9169 (N_9169,N_7825,N_5621);
and U9170 (N_9170,N_6859,N_6957);
nor U9171 (N_9171,N_6056,N_5997);
or U9172 (N_9172,N_7941,N_4031);
nor U9173 (N_9173,N_5900,N_7088);
or U9174 (N_9174,N_5001,N_5340);
nor U9175 (N_9175,N_6429,N_6279);
or U9176 (N_9176,N_4215,N_4835);
and U9177 (N_9177,N_6698,N_4120);
nand U9178 (N_9178,N_4411,N_5727);
nor U9179 (N_9179,N_4218,N_4956);
or U9180 (N_9180,N_7607,N_7711);
and U9181 (N_9181,N_4047,N_7565);
or U9182 (N_9182,N_7513,N_4431);
nand U9183 (N_9183,N_4564,N_4223);
and U9184 (N_9184,N_6188,N_4397);
or U9185 (N_9185,N_6389,N_7852);
and U9186 (N_9186,N_4900,N_6765);
nor U9187 (N_9187,N_5432,N_4434);
nor U9188 (N_9188,N_5707,N_5270);
and U9189 (N_9189,N_5806,N_7432);
or U9190 (N_9190,N_7792,N_7409);
nor U9191 (N_9191,N_5747,N_5564);
and U9192 (N_9192,N_5151,N_5310);
and U9193 (N_9193,N_7014,N_6187);
nor U9194 (N_9194,N_5708,N_6679);
or U9195 (N_9195,N_4068,N_6278);
nand U9196 (N_9196,N_6238,N_6907);
or U9197 (N_9197,N_5453,N_7751);
nand U9198 (N_9198,N_4108,N_5521);
xor U9199 (N_9199,N_7582,N_5427);
nand U9200 (N_9200,N_6686,N_7288);
or U9201 (N_9201,N_7120,N_4510);
nand U9202 (N_9202,N_5142,N_6419);
or U9203 (N_9203,N_7571,N_7245);
or U9204 (N_9204,N_6183,N_4729);
nand U9205 (N_9205,N_5855,N_7763);
nand U9206 (N_9206,N_6385,N_7871);
and U9207 (N_9207,N_6589,N_4836);
nand U9208 (N_9208,N_7464,N_6551);
and U9209 (N_9209,N_7725,N_4038);
nor U9210 (N_9210,N_6992,N_5391);
nor U9211 (N_9211,N_7676,N_5412);
nand U9212 (N_9212,N_5007,N_4997);
nor U9213 (N_9213,N_4884,N_7207);
or U9214 (N_9214,N_4041,N_7060);
or U9215 (N_9215,N_5182,N_4357);
and U9216 (N_9216,N_6921,N_4412);
or U9217 (N_9217,N_4785,N_4154);
and U9218 (N_9218,N_6105,N_7869);
nand U9219 (N_9219,N_6170,N_5218);
nand U9220 (N_9220,N_4087,N_6011);
nand U9221 (N_9221,N_7299,N_4423);
nor U9222 (N_9222,N_6240,N_5611);
nor U9223 (N_9223,N_7942,N_7097);
nand U9224 (N_9224,N_4150,N_6510);
and U9225 (N_9225,N_6697,N_6643);
or U9226 (N_9226,N_4077,N_6047);
or U9227 (N_9227,N_5104,N_6362);
nor U9228 (N_9228,N_4768,N_7651);
nor U9229 (N_9229,N_6501,N_7266);
or U9230 (N_9230,N_6036,N_5070);
and U9231 (N_9231,N_7770,N_6946);
or U9232 (N_9232,N_5362,N_5789);
and U9233 (N_9233,N_4290,N_6113);
nand U9234 (N_9234,N_5456,N_4499);
nand U9235 (N_9235,N_7085,N_5622);
or U9236 (N_9236,N_6577,N_7320);
and U9237 (N_9237,N_7702,N_4516);
nand U9238 (N_9238,N_4225,N_5695);
nand U9239 (N_9239,N_6631,N_4353);
or U9240 (N_9240,N_5005,N_6270);
and U9241 (N_9241,N_6122,N_5275);
or U9242 (N_9242,N_6138,N_4994);
and U9243 (N_9243,N_6928,N_6062);
and U9244 (N_9244,N_4263,N_6516);
or U9245 (N_9245,N_4545,N_7459);
and U9246 (N_9246,N_6255,N_4685);
and U9247 (N_9247,N_6100,N_7935);
nor U9248 (N_9248,N_6092,N_7160);
and U9249 (N_9249,N_7492,N_5518);
or U9250 (N_9250,N_7897,N_4880);
and U9251 (N_9251,N_7485,N_5169);
or U9252 (N_9252,N_4491,N_7482);
nor U9253 (N_9253,N_7360,N_5524);
nor U9254 (N_9254,N_7664,N_6620);
nand U9255 (N_9255,N_7790,N_4418);
nor U9256 (N_9256,N_7039,N_7460);
or U9257 (N_9257,N_5397,N_5060);
or U9258 (N_9258,N_5810,N_5467);
or U9259 (N_9259,N_4713,N_6506);
and U9260 (N_9260,N_6061,N_6852);
nor U9261 (N_9261,N_5802,N_7799);
and U9262 (N_9262,N_6112,N_6652);
or U9263 (N_9263,N_6489,N_6349);
nand U9264 (N_9264,N_4091,N_7222);
nand U9265 (N_9265,N_7367,N_7779);
nor U9266 (N_9266,N_6974,N_7945);
nor U9267 (N_9267,N_4644,N_6993);
nor U9268 (N_9268,N_6554,N_5937);
and U9269 (N_9269,N_7639,N_4827);
and U9270 (N_9270,N_6301,N_5755);
or U9271 (N_9271,N_4852,N_4209);
and U9272 (N_9272,N_6466,N_5764);
nand U9273 (N_9273,N_5702,N_6899);
or U9274 (N_9274,N_6307,N_6283);
and U9275 (N_9275,N_6146,N_4079);
nand U9276 (N_9276,N_5304,N_6103);
or U9277 (N_9277,N_6057,N_6761);
nor U9278 (N_9278,N_4979,N_5603);
and U9279 (N_9279,N_5556,N_7896);
and U9280 (N_9280,N_4924,N_4059);
and U9281 (N_9281,N_7905,N_4029);
nor U9282 (N_9282,N_5904,N_6741);
or U9283 (N_9283,N_7955,N_6087);
nor U9284 (N_9284,N_4360,N_6009);
nor U9285 (N_9285,N_5037,N_6598);
or U9286 (N_9286,N_4579,N_4726);
or U9287 (N_9287,N_7505,N_6281);
or U9288 (N_9288,N_4025,N_6521);
nand U9289 (N_9289,N_4770,N_7560);
nor U9290 (N_9290,N_6035,N_4315);
or U9291 (N_9291,N_5159,N_6232);
nor U9292 (N_9292,N_4119,N_4752);
xor U9293 (N_9293,N_6158,N_6746);
nor U9294 (N_9294,N_5932,N_5190);
nor U9295 (N_9295,N_7976,N_5021);
or U9296 (N_9296,N_6916,N_7536);
nor U9297 (N_9297,N_4978,N_4822);
nor U9298 (N_9298,N_6478,N_6292);
and U9299 (N_9299,N_7959,N_7351);
and U9300 (N_9300,N_4570,N_4210);
and U9301 (N_9301,N_5583,N_4525);
nand U9302 (N_9302,N_6740,N_6569);
or U9303 (N_9303,N_4419,N_4692);
nor U9304 (N_9304,N_5787,N_4190);
xnor U9305 (N_9305,N_6826,N_4338);
or U9306 (N_9306,N_7140,N_4959);
and U9307 (N_9307,N_6295,N_4549);
or U9308 (N_9308,N_6355,N_4543);
and U9309 (N_9309,N_5776,N_7848);
or U9310 (N_9310,N_7111,N_7684);
nand U9311 (N_9311,N_4914,N_4456);
nand U9312 (N_9312,N_4632,N_5590);
nor U9313 (N_9313,N_5163,N_5558);
nand U9314 (N_9314,N_4792,N_4913);
or U9315 (N_9315,N_4963,N_4180);
nor U9316 (N_9316,N_6168,N_4810);
nor U9317 (N_9317,N_7418,N_5779);
and U9318 (N_9318,N_5395,N_7556);
nand U9319 (N_9319,N_6575,N_6203);
and U9320 (N_9320,N_6219,N_7392);
or U9321 (N_9321,N_7087,N_7823);
nor U9322 (N_9322,N_7457,N_7192);
nand U9323 (N_9323,N_5352,N_6690);
and U9324 (N_9324,N_6020,N_7294);
nor U9325 (N_9325,N_6351,N_5004);
nand U9326 (N_9326,N_6876,N_7652);
nand U9327 (N_9327,N_5735,N_5619);
or U9328 (N_9328,N_5782,N_5118);
nand U9329 (N_9329,N_6101,N_4863);
nand U9330 (N_9330,N_6384,N_5305);
or U9331 (N_9331,N_5774,N_7325);
nor U9332 (N_9332,N_7908,N_7678);
and U9333 (N_9333,N_6465,N_6214);
and U9334 (N_9334,N_5332,N_6536);
nor U9335 (N_9335,N_5972,N_7093);
nor U9336 (N_9336,N_7572,N_5610);
nor U9337 (N_9337,N_7276,N_5095);
or U9338 (N_9338,N_4718,N_7204);
nand U9339 (N_9339,N_4593,N_6526);
nor U9340 (N_9340,N_5063,N_5068);
or U9341 (N_9341,N_7870,N_4535);
or U9342 (N_9342,N_6701,N_4224);
or U9343 (N_9343,N_6392,N_5268);
nand U9344 (N_9344,N_6015,N_7036);
or U9345 (N_9345,N_4883,N_5844);
nor U9346 (N_9346,N_5604,N_4480);
and U9347 (N_9347,N_4129,N_7593);
nor U9348 (N_9348,N_7740,N_5701);
nand U9349 (N_9349,N_7228,N_4928);
nor U9350 (N_9350,N_5836,N_7581);
or U9351 (N_9351,N_4303,N_4731);
nand U9352 (N_9352,N_4089,N_7084);
or U9353 (N_9353,N_4193,N_5025);
or U9354 (N_9354,N_4853,N_4008);
or U9355 (N_9355,N_4366,N_6044);
nor U9356 (N_9356,N_7076,N_7490);
and U9357 (N_9357,N_6502,N_4138);
and U9358 (N_9358,N_7845,N_4301);
nand U9359 (N_9359,N_5474,N_4341);
nand U9360 (N_9360,N_5914,N_4408);
nand U9361 (N_9361,N_6695,N_6857);
and U9362 (N_9362,N_6178,N_7670);
nor U9363 (N_9363,N_5246,N_6494);
nand U9364 (N_9364,N_5198,N_5950);
xnor U9365 (N_9365,N_6284,N_7752);
nor U9366 (N_9366,N_7630,N_4242);
or U9367 (N_9367,N_7290,N_4121);
nor U9368 (N_9368,N_4386,N_6889);
and U9369 (N_9369,N_5085,N_6668);
or U9370 (N_9370,N_6059,N_7946);
nand U9371 (N_9371,N_7308,N_4382);
nor U9372 (N_9372,N_5414,N_6080);
nand U9373 (N_9373,N_7853,N_7749);
xor U9374 (N_9374,N_6263,N_6671);
nand U9375 (N_9375,N_5679,N_6442);
or U9376 (N_9376,N_6241,N_5852);
xor U9377 (N_9377,N_7854,N_5709);
and U9378 (N_9378,N_6795,N_5260);
nand U9379 (N_9379,N_4897,N_4261);
or U9380 (N_9380,N_7921,N_4222);
nor U9381 (N_9381,N_6762,N_5748);
nand U9382 (N_9382,N_5232,N_7498);
nor U9383 (N_9383,N_5164,N_6661);
or U9384 (N_9384,N_5353,N_7407);
xnor U9385 (N_9385,N_7827,N_6427);
nand U9386 (N_9386,N_6956,N_4013);
nor U9387 (N_9387,N_7175,N_6276);
xnor U9388 (N_9388,N_7605,N_6834);
or U9389 (N_9389,N_7710,N_7230);
and U9390 (N_9390,N_6312,N_7069);
nor U9391 (N_9391,N_5162,N_6659);
or U9392 (N_9392,N_4123,N_7215);
or U9393 (N_9393,N_4920,N_5624);
or U9394 (N_9394,N_6520,N_5854);
nor U9395 (N_9395,N_5503,N_4657);
nor U9396 (N_9396,N_6160,N_7277);
nand U9397 (N_9397,N_6562,N_5962);
nor U9398 (N_9398,N_4391,N_7196);
or U9399 (N_9399,N_4140,N_5757);
or U9400 (N_9400,N_6779,N_7844);
nand U9401 (N_9401,N_7311,N_7438);
and U9402 (N_9402,N_7535,N_6640);
or U9403 (N_9403,N_5627,N_6924);
nor U9404 (N_9404,N_5859,N_4379);
nand U9405 (N_9405,N_7115,N_4999);
or U9406 (N_9406,N_6715,N_5185);
nand U9407 (N_9407,N_4221,N_6657);
and U9408 (N_9408,N_4895,N_7894);
nor U9409 (N_9409,N_6790,N_4293);
nand U9410 (N_9410,N_6597,N_6991);
nor U9411 (N_9411,N_7545,N_6682);
and U9412 (N_9412,N_6749,N_5437);
and U9413 (N_9413,N_6674,N_7774);
or U9414 (N_9414,N_4026,N_6143);
or U9415 (N_9415,N_6549,N_5447);
or U9416 (N_9416,N_7701,N_7231);
nor U9417 (N_9417,N_5267,N_7631);
and U9418 (N_9418,N_4538,N_7783);
or U9419 (N_9419,N_7798,N_5263);
nor U9420 (N_9420,N_4679,N_7295);
nor U9421 (N_9421,N_7707,N_7328);
or U9422 (N_9422,N_5324,N_5915);
nand U9423 (N_9423,N_6662,N_5469);
or U9424 (N_9424,N_6837,N_4971);
nand U9425 (N_9425,N_4670,N_4582);
and U9426 (N_9426,N_6669,N_7050);
or U9427 (N_9427,N_5053,N_4774);
and U9428 (N_9428,N_7150,N_4750);
and U9429 (N_9429,N_6366,N_6645);
or U9430 (N_9430,N_6851,N_6054);
and U9431 (N_9431,N_7580,N_6767);
nand U9432 (N_9432,N_6027,N_7972);
nand U9433 (N_9433,N_4262,N_7519);
nor U9434 (N_9434,N_7874,N_6001);
xnor U9435 (N_9435,N_5009,N_4811);
nor U9436 (N_9436,N_5711,N_7021);
and U9437 (N_9437,N_7732,N_4723);
and U9438 (N_9438,N_5487,N_7124);
and U9439 (N_9439,N_6919,N_6002);
and U9440 (N_9440,N_4216,N_4992);
nor U9441 (N_9441,N_7168,N_6206);
or U9442 (N_9442,N_7553,N_4274);
nand U9443 (N_9443,N_6063,N_5739);
and U9444 (N_9444,N_4062,N_6450);
and U9445 (N_9445,N_4245,N_7687);
nand U9446 (N_9446,N_5689,N_6352);
and U9447 (N_9447,N_5801,N_6106);
nor U9448 (N_9448,N_6958,N_7137);
or U9449 (N_9449,N_4465,N_5073);
or U9450 (N_9450,N_7531,N_6621);
or U9451 (N_9451,N_4602,N_7380);
and U9452 (N_9452,N_5952,N_7389);
nand U9453 (N_9453,N_6905,N_7855);
and U9454 (N_9454,N_4534,N_4133);
nand U9455 (N_9455,N_4308,N_7766);
or U9456 (N_9456,N_4905,N_4691);
nand U9457 (N_9457,N_6827,N_4039);
and U9458 (N_9458,N_6608,N_7073);
nor U9459 (N_9459,N_5158,N_7672);
nor U9460 (N_9460,N_6954,N_5570);
nor U9461 (N_9461,N_7653,N_7570);
and U9462 (N_9462,N_4455,N_5560);
and U9463 (N_9463,N_5729,N_7127);
and U9464 (N_9464,N_6648,N_7086);
nor U9465 (N_9465,N_6927,N_6512);
nor U9466 (N_9466,N_5288,N_6885);
nand U9467 (N_9467,N_4518,N_6134);
xor U9468 (N_9468,N_5043,N_6997);
or U9469 (N_9469,N_4375,N_6074);
and U9470 (N_9470,N_4273,N_5878);
and U9471 (N_9471,N_4134,N_4252);
and U9472 (N_9472,N_7714,N_7062);
or U9473 (N_9473,N_4812,N_4399);
nor U9474 (N_9474,N_7694,N_6252);
xnor U9475 (N_9475,N_5654,N_6783);
or U9476 (N_9476,N_5851,N_6073);
nand U9477 (N_9477,N_6775,N_4875);
nor U9478 (N_9478,N_7964,N_4710);
or U9479 (N_9479,N_4329,N_5278);
nand U9480 (N_9480,N_4021,N_4128);
nor U9481 (N_9481,N_5581,N_5325);
nand U9482 (N_9482,N_6424,N_7719);
and U9483 (N_9483,N_4765,N_5791);
nor U9484 (N_9484,N_5186,N_7967);
or U9485 (N_9485,N_6192,N_6689);
and U9486 (N_9486,N_6018,N_5350);
nor U9487 (N_9487,N_7785,N_6658);
or U9488 (N_9488,N_6175,N_5203);
or U9489 (N_9489,N_6867,N_6340);
nand U9490 (N_9490,N_4500,N_7229);
nand U9491 (N_9491,N_5824,N_4704);
and U9492 (N_9492,N_6226,N_5847);
nand U9493 (N_9493,N_6163,N_6601);
nand U9494 (N_9494,N_5309,N_6945);
nand U9495 (N_9495,N_7978,N_7579);
or U9496 (N_9496,N_4048,N_4663);
nand U9497 (N_9497,N_4113,N_5132);
or U9498 (N_9498,N_4699,N_4813);
nor U9499 (N_9499,N_4603,N_7181);
nor U9500 (N_9500,N_4426,N_5490);
nor U9501 (N_9501,N_7068,N_4171);
or U9502 (N_9502,N_5294,N_5421);
and U9503 (N_9503,N_4207,N_6194);
nor U9504 (N_9504,N_7415,N_6806);
or U9505 (N_9505,N_6534,N_6816);
nand U9506 (N_9506,N_4558,N_5256);
and U9507 (N_9507,N_7433,N_7385);
nor U9508 (N_9508,N_5211,N_5772);
xor U9509 (N_9509,N_4060,N_7867);
and U9510 (N_9510,N_5153,N_7353);
or U9511 (N_9511,N_7251,N_4929);
or U9512 (N_9512,N_6415,N_7113);
nand U9513 (N_9513,N_6553,N_7782);
or U9514 (N_9514,N_5561,N_4513);
or U9515 (N_9515,N_4507,N_7550);
and U9516 (N_9516,N_6447,N_5983);
or U9517 (N_9517,N_4226,N_5188);
nor U9518 (N_9518,N_7428,N_7919);
or U9519 (N_9519,N_7501,N_4142);
or U9520 (N_9520,N_7037,N_4671);
nand U9521 (N_9521,N_5493,N_6326);
and U9522 (N_9522,N_7554,N_7348);
or U9523 (N_9523,N_7646,N_7279);
or U9524 (N_9524,N_4406,N_6793);
nor U9525 (N_9525,N_6947,N_4932);
xnor U9526 (N_9526,N_5422,N_5813);
and U9527 (N_9527,N_6579,N_6500);
nand U9528 (N_9528,N_6140,N_5796);
nor U9529 (N_9529,N_6234,N_4594);
nand U9530 (N_9530,N_4717,N_6425);
or U9531 (N_9531,N_7281,N_5516);
nor U9532 (N_9532,N_4972,N_5935);
nand U9533 (N_9533,N_6345,N_4392);
and U9534 (N_9534,N_6952,N_7895);
and U9535 (N_9535,N_6290,N_7597);
and U9536 (N_9536,N_5127,N_4117);
or U9537 (N_9537,N_7474,N_4078);
nor U9538 (N_9538,N_5699,N_4701);
and U9539 (N_9539,N_5113,N_5138);
and U9540 (N_9540,N_4036,N_5212);
nor U9541 (N_9541,N_7399,N_6131);
nor U9542 (N_9542,N_6000,N_6939);
nand U9543 (N_9543,N_7659,N_6870);
nor U9544 (N_9544,N_4302,N_4348);
and U9545 (N_9545,N_4321,N_5259);
and U9546 (N_9546,N_4531,N_7598);
nand U9547 (N_9547,N_6821,N_7119);
nand U9548 (N_9548,N_4649,N_7619);
nor U9549 (N_9549,N_6639,N_7044);
nand U9550 (N_9550,N_5948,N_4939);
nor U9551 (N_9551,N_7041,N_5803);
and U9552 (N_9552,N_6524,N_4821);
nand U9553 (N_9553,N_7366,N_6819);
or U9554 (N_9554,N_6468,N_6609);
xor U9555 (N_9555,N_4374,N_6272);
and U9556 (N_9556,N_7063,N_5714);
nor U9557 (N_9557,N_6030,N_5580);
or U9558 (N_9558,N_5471,N_5589);
or U9559 (N_9559,N_7806,N_5055);
or U9560 (N_9560,N_5990,N_5376);
nor U9561 (N_9561,N_5476,N_6843);
nand U9562 (N_9562,N_7901,N_7370);
nor U9563 (N_9563,N_5369,N_4220);
or U9564 (N_9564,N_4725,N_4730);
nand U9565 (N_9565,N_6627,N_4409);
or U9566 (N_9566,N_4156,N_4344);
nor U9567 (N_9567,N_4045,N_7756);
and U9568 (N_9568,N_4789,N_6297);
or U9569 (N_9569,N_5615,N_4433);
xor U9570 (N_9570,N_6670,N_6511);
or U9571 (N_9571,N_6431,N_7940);
xnor U9572 (N_9572,N_7383,N_6700);
nor U9573 (N_9573,N_4356,N_7148);
and U9574 (N_9574,N_4808,N_5202);
or U9575 (N_9575,N_7208,N_5548);
nand U9576 (N_9576,N_4666,N_7983);
or U9577 (N_9577,N_7636,N_6490);
xnor U9578 (N_9578,N_6546,N_7411);
or U9579 (N_9579,N_5875,N_6719);
nand U9580 (N_9580,N_7878,N_6359);
or U9581 (N_9581,N_4562,N_4861);
nor U9582 (N_9582,N_4405,N_6752);
nand U9583 (N_9583,N_7190,N_7910);
nor U9584 (N_9584,N_5027,N_5365);
nor U9585 (N_9585,N_5698,N_5777);
nor U9586 (N_9586,N_7356,N_4256);
and U9587 (N_9587,N_4161,N_5116);
nand U9588 (N_9588,N_5322,N_7602);
and U9589 (N_9589,N_5338,N_7850);
nor U9590 (N_9590,N_7829,N_7499);
nand U9591 (N_9591,N_4816,N_7098);
and U9592 (N_9592,N_7038,N_4466);
nand U9593 (N_9593,N_5341,N_4454);
nand U9594 (N_9594,N_5014,N_6291);
xor U9595 (N_9595,N_7004,N_6356);
and U9596 (N_9596,N_7240,N_7427);
and U9597 (N_9597,N_4954,N_7858);
nand U9598 (N_9598,N_4508,N_5569);
nand U9599 (N_9599,N_6699,N_5917);
nand U9600 (N_9600,N_4809,N_4449);
and U9601 (N_9601,N_6253,N_5289);
or U9602 (N_9602,N_5760,N_4996);
nor U9603 (N_9603,N_5691,N_4420);
nor U9604 (N_9604,N_7892,N_7029);
nor U9605 (N_9605,N_5301,N_6469);
or U9606 (N_9606,N_5947,N_4739);
and U9607 (N_9607,N_5481,N_5613);
nand U9608 (N_9608,N_6167,N_6104);
or U9609 (N_9609,N_4830,N_5204);
nor U9610 (N_9610,N_5279,N_6195);
nand U9611 (N_9611,N_7618,N_6386);
and U9612 (N_9612,N_4264,N_4072);
and U9613 (N_9613,N_5083,N_7200);
nor U9614 (N_9614,N_4877,N_5176);
nand U9615 (N_9615,N_7114,N_4585);
or U9616 (N_9616,N_6978,N_7760);
nand U9617 (N_9617,N_4623,N_4643);
nand U9618 (N_9618,N_7446,N_6199);
nor U9619 (N_9619,N_4887,N_5514);
nand U9620 (N_9620,N_4071,N_6563);
nor U9621 (N_9621,N_5187,N_7323);
nand U9622 (N_9622,N_5901,N_4758);
nand U9623 (N_9623,N_7643,N_6262);
nor U9624 (N_9624,N_4415,N_5887);
xor U9625 (N_9625,N_5665,N_7333);
or U9626 (N_9626,N_4872,N_6093);
and U9627 (N_9627,N_4248,N_4266);
nand U9628 (N_9628,N_6807,N_5334);
nand U9629 (N_9629,N_5954,N_4553);
or U9630 (N_9630,N_7891,N_5455);
nor U9631 (N_9631,N_4915,N_6680);
nor U9632 (N_9632,N_7268,N_5812);
and U9633 (N_9633,N_6473,N_6342);
and U9634 (N_9634,N_5141,N_5635);
nor U9635 (N_9635,N_7194,N_6970);
nor U9636 (N_9636,N_5629,N_7623);
or U9637 (N_9637,N_4716,N_5992);
nor U9638 (N_9638,N_5266,N_7110);
nand U9639 (N_9639,N_7382,N_6434);
nor U9640 (N_9640,N_7872,N_6318);
or U9641 (N_9641,N_5221,N_6023);
or U9642 (N_9642,N_6637,N_7948);
nor U9643 (N_9643,N_6117,N_5019);
or U9644 (N_9644,N_5919,N_5643);
nor U9645 (N_9645,N_4901,N_4541);
nor U9646 (N_9646,N_4773,N_4987);
and U9647 (N_9647,N_6543,N_7032);
nand U9648 (N_9648,N_6963,N_5641);
nor U9649 (N_9649,N_4046,N_6692);
nor U9650 (N_9650,N_5498,N_4173);
nor U9651 (N_9651,N_6309,N_5936);
and U9652 (N_9652,N_5321,N_4586);
or U9653 (N_9653,N_4873,N_6382);
nor U9654 (N_9654,N_5192,N_7984);
or U9655 (N_9655,N_4784,N_5831);
and U9656 (N_9656,N_7813,N_6918);
nand U9657 (N_9657,N_5110,N_6498);
and U9658 (N_9658,N_5328,N_5968);
nor U9659 (N_9659,N_5167,N_5743);
nand U9660 (N_9660,N_7350,N_5804);
or U9661 (N_9661,N_5808,N_6314);
nor U9662 (N_9662,N_4149,N_4170);
or U9663 (N_9663,N_7956,N_7943);
and U9664 (N_9664,N_6126,N_7361);
nand U9665 (N_9665,N_7691,N_4719);
or U9666 (N_9666,N_7386,N_5092);
nor U9667 (N_9667,N_7419,N_5120);
nand U9668 (N_9668,N_6618,N_5924);
and U9669 (N_9669,N_7584,N_4746);
or U9670 (N_9670,N_6936,N_7814);
nor U9671 (N_9671,N_4528,N_5360);
or U9672 (N_9672,N_5523,N_4483);
and U9673 (N_9673,N_7957,N_6600);
and U9674 (N_9674,N_7258,N_4862);
or U9675 (N_9675,N_4231,N_7449);
nor U9676 (N_9676,N_6844,N_7547);
nor U9677 (N_9677,N_7922,N_5337);
or U9678 (N_9678,N_6476,N_6665);
nor U9679 (N_9679,N_5899,N_7637);
and U9680 (N_9680,N_5642,N_7540);
nor U9681 (N_9681,N_7573,N_7470);
and U9682 (N_9682,N_7011,N_6124);
or U9683 (N_9683,N_5930,N_7600);
nand U9684 (N_9684,N_4636,N_4403);
or U9685 (N_9685,N_7154,N_4144);
nand U9686 (N_9686,N_4721,N_7820);
or U9687 (N_9687,N_7660,N_6260);
and U9688 (N_9688,N_4753,N_6850);
nor U9689 (N_9689,N_4844,N_4269);
nand U9690 (N_9690,N_4146,N_5956);
nand U9691 (N_9691,N_4794,N_4837);
nand U9692 (N_9692,N_7458,N_4854);
and U9693 (N_9693,N_5529,N_5449);
or U9694 (N_9694,N_5023,N_4034);
nor U9695 (N_9695,N_5946,N_6969);
and U9696 (N_9696,N_4722,N_5425);
nor U9697 (N_9697,N_5838,N_5694);
or U9698 (N_9698,N_7138,N_6735);
xor U9699 (N_9699,N_5805,N_5960);
nor U9700 (N_9700,N_7696,N_4807);
and U9701 (N_9701,N_7141,N_7312);
and U9702 (N_9702,N_7456,N_6833);
nand U9703 (N_9703,N_5128,N_7679);
nor U9704 (N_9704,N_7246,N_4778);
nor U9705 (N_9705,N_6208,N_6085);
or U9706 (N_9706,N_7384,N_7104);
or U9707 (N_9707,N_4886,N_6904);
and U9708 (N_9708,N_4027,N_4540);
nand U9709 (N_9709,N_4667,N_7675);
or U9710 (N_9710,N_6110,N_7998);
or U9711 (N_9711,N_5465,N_5017);
nor U9712 (N_9712,N_7644,N_4019);
or U9713 (N_9713,N_5244,N_6202);
nor U9714 (N_9714,N_4934,N_5978);
nor U9715 (N_9715,N_5489,N_7378);
and U9716 (N_9716,N_5233,N_5920);
and U9717 (N_9717,N_4912,N_6198);
nand U9718 (N_9718,N_5821,N_5669);
nand U9719 (N_9719,N_4174,N_5765);
or U9720 (N_9720,N_6320,N_5745);
nor U9721 (N_9721,N_7583,N_6572);
nor U9722 (N_9722,N_5241,N_4782);
or U9723 (N_9723,N_6064,N_4402);
or U9724 (N_9724,N_7339,N_7803);
nand U9725 (N_9725,N_4970,N_5434);
nand U9726 (N_9726,N_6492,N_6538);
and U9727 (N_9727,N_7884,N_6858);
or U9728 (N_9728,N_7107,N_4985);
nand U9729 (N_9729,N_5820,N_7863);
nand U9730 (N_9730,N_4102,N_7889);
xor U9731 (N_9731,N_7020,N_4110);
xor U9732 (N_9732,N_5436,N_4548);
or U9733 (N_9733,N_7826,N_5599);
or U9734 (N_9734,N_7447,N_4968);
nor U9735 (N_9735,N_6186,N_7879);
or U9736 (N_9736,N_5348,N_4680);
xnor U9737 (N_9737,N_7248,N_5797);
nand U9738 (N_9738,N_4859,N_6406);
and U9739 (N_9739,N_4057,N_5546);
nor U9740 (N_9740,N_5841,N_7436);
or U9741 (N_9741,N_5726,N_6324);
and U9742 (N_9742,N_6403,N_6296);
nand U9743 (N_9743,N_4476,N_5605);
and U9744 (N_9744,N_5227,N_4727);
nand U9745 (N_9745,N_5673,N_7042);
and U9746 (N_9746,N_5792,N_5559);
nand U9747 (N_9747,N_4111,N_5373);
or U9748 (N_9748,N_5015,N_5886);
or U9749 (N_9749,N_7991,N_6327);
xor U9750 (N_9750,N_4524,N_5579);
or U9751 (N_9751,N_4974,N_6344);
nand U9752 (N_9752,N_7769,N_5982);
nand U9753 (N_9753,N_4849,N_7568);
or U9754 (N_9754,N_7031,N_5766);
and U9755 (N_9755,N_7950,N_5078);
and U9756 (N_9756,N_7543,N_4448);
and U9757 (N_9757,N_4696,N_6782);
and U9758 (N_9758,N_7423,N_5143);
nor U9759 (N_9759,N_7316,N_6174);
and U9760 (N_9760,N_7241,N_7818);
or U9761 (N_9761,N_4567,N_4283);
and U9762 (N_9762,N_5121,N_6416);
and U9763 (N_9763,N_6770,N_4936);
or U9764 (N_9764,N_6881,N_4953);
or U9765 (N_9765,N_7974,N_4240);
or U9766 (N_9766,N_6709,N_4568);
nor U9767 (N_9767,N_7422,N_7187);
nor U9768 (N_9768,N_6404,N_7329);
nand U9769 (N_9769,N_6443,N_5988);
nor U9770 (N_9770,N_6184,N_6614);
nand U9771 (N_9771,N_5318,N_5170);
and U9772 (N_9772,N_7238,N_5906);
nand U9773 (N_9773,N_5075,N_7533);
and U9774 (N_9774,N_4885,N_4219);
and U9775 (N_9775,N_4061,N_4337);
nor U9776 (N_9776,N_7061,N_6136);
nand U9777 (N_9777,N_6286,N_7522);
or U9778 (N_9778,N_4304,N_4664);
and U9779 (N_9779,N_5877,N_4229);
and U9780 (N_9780,N_6505,N_6217);
nand U9781 (N_9781,N_7632,N_7262);
nand U9782 (N_9782,N_7227,N_5618);
nand U9783 (N_9783,N_7726,N_4259);
nand U9784 (N_9784,N_6487,N_6622);
or U9785 (N_9785,N_6776,N_4137);
or U9786 (N_9786,N_5759,N_6222);
and U9787 (N_9787,N_4030,N_7667);
nand U9788 (N_9788,N_7218,N_4317);
or U9789 (N_9789,N_4689,N_5634);
nor U9790 (N_9790,N_4975,N_7773);
nand U9791 (N_9791,N_5883,N_5280);
nand U9792 (N_9792,N_4206,N_5942);
and U9793 (N_9793,N_4892,N_6786);
or U9794 (N_9794,N_7410,N_4461);
or U9795 (N_9795,N_7689,N_6475);
and U9796 (N_9796,N_7398,N_5308);
or U9797 (N_9797,N_5358,N_7649);
or U9798 (N_9798,N_6771,N_4639);
and U9799 (N_9799,N_4728,N_5248);
nand U9800 (N_9800,N_4023,N_7188);
xor U9801 (N_9801,N_6582,N_7106);
and U9802 (N_9802,N_4112,N_5058);
or U9803 (N_9803,N_4621,N_7100);
or U9804 (N_9804,N_5385,N_7979);
nand U9805 (N_9805,N_4733,N_4387);
nor U9806 (N_9806,N_5674,N_5720);
nand U9807 (N_9807,N_5448,N_5311);
and U9808 (N_9808,N_5573,N_5584);
nand U9809 (N_9809,N_5816,N_4132);
nand U9810 (N_9810,N_7242,N_6841);
xnor U9811 (N_9811,N_6407,N_7437);
nor U9812 (N_9812,N_6651,N_4306);
nand U9813 (N_9813,N_7655,N_5929);
nor U9814 (N_9814,N_4157,N_5313);
and U9815 (N_9815,N_7405,N_4909);
or U9816 (N_9816,N_7777,N_5081);
or U9817 (N_9817,N_6435,N_5785);
nand U9818 (N_9818,N_7893,N_5631);
nor U9819 (N_9819,N_4703,N_6736);
nand U9820 (N_9820,N_7172,N_6725);
nand U9821 (N_9821,N_6830,N_4948);
or U9822 (N_9822,N_5125,N_6361);
and U9823 (N_9823,N_7252,N_7397);
or U9824 (N_9824,N_4511,N_7182);
and U9825 (N_9825,N_7890,N_7484);
nor U9826 (N_9826,N_5499,N_6196);
nor U9827 (N_9827,N_5540,N_7520);
nor U9828 (N_9828,N_4484,N_7429);
and U9829 (N_9829,N_7576,N_7682);
and U9830 (N_9830,N_7341,N_5458);
nor U9831 (N_9831,N_6412,N_4064);
and U9832 (N_9832,N_4917,N_4101);
or U9833 (N_9833,N_6972,N_5912);
or U9834 (N_9834,N_6901,N_4738);
or U9835 (N_9835,N_6055,N_6029);
and U9836 (N_9836,N_5438,N_4505);
nand U9837 (N_9837,N_5160,N_5461);
or U9838 (N_9838,N_7287,N_7091);
xor U9839 (N_9839,N_6593,N_5292);
nor U9840 (N_9840,N_7072,N_6258);
nor U9841 (N_9841,N_7787,N_4919);
nand U9842 (N_9842,N_6350,N_4316);
or U9843 (N_9843,N_6497,N_7396);
nand U9844 (N_9844,N_6376,N_6316);
and U9845 (N_9845,N_7007,N_6471);
and U9846 (N_9846,N_4537,N_7013);
and U9847 (N_9847,N_5124,N_5215);
nor U9848 (N_9848,N_7786,N_5049);
and U9849 (N_9849,N_7205,N_6335);
or U9850 (N_9850,N_6225,N_5364);
and U9851 (N_9851,N_7034,N_7219);
nand U9852 (N_9852,N_7926,N_6189);
and U9853 (N_9853,N_6823,N_5459);
nor U9854 (N_9854,N_7487,N_6398);
xor U9855 (N_9855,N_7601,N_7022);
nand U9856 (N_9856,N_4011,N_7256);
xor U9857 (N_9857,N_4826,N_6288);
or U9858 (N_9858,N_7226,N_4532);
nand U9859 (N_9859,N_4709,N_7563);
and U9860 (N_9860,N_4143,N_5346);
nand U9861 (N_9861,N_4539,N_7271);
nor U9862 (N_9862,N_7340,N_5638);
or U9863 (N_9863,N_7641,N_6799);
nor U9864 (N_9864,N_5129,N_7745);
or U9865 (N_9865,N_7315,N_6390);
xor U9866 (N_9866,N_4313,N_4130);
nand U9867 (N_9867,N_7047,N_6216);
or U9868 (N_9868,N_6718,N_4151);
and U9869 (N_9869,N_7833,N_5264);
nand U9870 (N_9870,N_5374,N_5165);
or U9871 (N_9871,N_7289,N_5112);
and U9872 (N_9872,N_5088,N_5640);
and U9873 (N_9873,N_5439,N_5050);
nor U9874 (N_9874,N_5146,N_5320);
and U9875 (N_9875,N_5220,N_7524);
or U9876 (N_9876,N_5298,N_6726);
nand U9877 (N_9877,N_7836,N_4935);
or U9878 (N_9878,N_4197,N_7354);
nor U9879 (N_9879,N_6529,N_6599);
or U9880 (N_9880,N_7843,N_4178);
or U9881 (N_9881,N_5366,N_7416);
or U9882 (N_9882,N_7209,N_7096);
or U9883 (N_9883,N_5171,N_7496);
nand U9884 (N_9884,N_7297,N_7177);
or U9885 (N_9885,N_5175,N_4661);
nor U9886 (N_9886,N_7549,N_6273);
nand U9887 (N_9887,N_4501,N_4851);
nand U9888 (N_9888,N_4918,N_6835);
xor U9889 (N_9889,N_5262,N_5965);
nand U9890 (N_9890,N_6277,N_5285);
or U9891 (N_9891,N_5941,N_5858);
nor U9892 (N_9892,N_6259,N_5245);
and U9893 (N_9893,N_7567,N_7856);
or U9894 (N_9894,N_6545,N_5656);
nor U9895 (N_9895,N_7920,N_5079);
nor U9896 (N_9896,N_7057,N_5849);
and U9897 (N_9897,N_7426,N_6070);
nand U9898 (N_9898,N_6322,N_4708);
or U9899 (N_9899,N_6571,N_4617);
nor U9900 (N_9900,N_4688,N_6938);
or U9901 (N_9901,N_7016,N_5351);
nand U9902 (N_9902,N_4604,N_6075);
nand U9903 (N_9903,N_7541,N_6929);
or U9904 (N_9904,N_4881,N_4673);
nand U9905 (N_9905,N_5630,N_7335);
nand U9906 (N_9906,N_5242,N_5660);
nor U9907 (N_9907,N_6574,N_6405);
nand U9908 (N_9908,N_5967,N_4070);
and U9909 (N_9909,N_7674,N_6499);
nor U9910 (N_9910,N_5566,N_7621);
nand U9911 (N_9911,N_6223,N_6014);
or U9912 (N_9912,N_6220,N_7994);
xor U9913 (N_9913,N_5096,N_4803);
xor U9914 (N_9914,N_6181,N_7270);
nor U9915 (N_9915,N_4910,N_5868);
and U9916 (N_9916,N_7183,N_5732);
nand U9917 (N_9917,N_6373,N_7040);
nand U9918 (N_9918,N_7888,N_4334);
or U9919 (N_9919,N_5963,N_6084);
and U9920 (N_9920,N_4819,N_6917);
nor U9921 (N_9921,N_7502,N_7357);
nand U9922 (N_9922,N_5513,N_7193);
nor U9923 (N_9923,N_4947,N_4135);
nor U9924 (N_9924,N_6115,N_4401);
and U9925 (N_9925,N_6965,N_7724);
and U9926 (N_9926,N_4611,N_5910);
nor U9927 (N_9927,N_4052,N_6051);
and U9928 (N_9928,N_6955,N_5734);
and U9929 (N_9929,N_6930,N_4683);
or U9930 (N_9930,N_5799,N_6470);
nor U9931 (N_9931,N_4080,N_7135);
nand U9932 (N_9932,N_5741,N_6660);
or U9933 (N_9933,N_6738,N_6337);
and U9934 (N_9934,N_5224,N_5061);
and U9935 (N_9935,N_6461,N_5576);
nand U9936 (N_9936,N_7500,N_4922);
xnor U9937 (N_9937,N_4828,N_6118);
or U9938 (N_9938,N_5644,N_7171);
or U9939 (N_9939,N_7167,N_5585);
or U9940 (N_9940,N_5161,N_6596);
and U9941 (N_9941,N_6624,N_7302);
nor U9942 (N_9942,N_7735,N_6890);
nand U9943 (N_9943,N_4186,N_5738);
nand U9944 (N_9944,N_5692,N_4148);
and U9945 (N_9945,N_6711,N_7947);
nor U9946 (N_9946,N_6144,N_7561);
nor U9947 (N_9947,N_5626,N_6311);
or U9948 (N_9948,N_6518,N_5577);
and U9949 (N_9949,N_7128,N_6825);
and U9950 (N_9950,N_5363,N_6942);
and U9951 (N_9951,N_5389,N_5793);
nor U9952 (N_9952,N_5874,N_7112);
and U9953 (N_9953,N_5035,N_5059);
nor U9954 (N_9954,N_6713,N_6943);
nand U9955 (N_9955,N_5372,N_6591);
and U9956 (N_9956,N_7510,N_7592);
and U9957 (N_9957,N_4136,N_4610);
or U9958 (N_9958,N_6068,N_7364);
nor U9959 (N_9959,N_7898,N_5016);
or U9960 (N_9960,N_6685,N_4949);
nor U9961 (N_9961,N_5491,N_6710);
and U9962 (N_9962,N_5415,N_5106);
nor U9963 (N_9963,N_7555,N_4751);
nand U9964 (N_9964,N_4620,N_5536);
and U9965 (N_9965,N_7313,N_6933);
nand U9966 (N_9966,N_4472,N_4049);
and U9967 (N_9967,N_4790,N_5676);
nand U9968 (N_9968,N_5976,N_7828);
nand U9969 (N_9969,N_5213,N_7793);
or U9970 (N_9970,N_5012,N_7365);
nand U9971 (N_9971,N_4573,N_5087);
nor U9972 (N_9972,N_4096,N_5998);
or U9973 (N_9973,N_7425,N_5678);
nand U9974 (N_9974,N_4384,N_6456);
nor U9975 (N_9975,N_7864,N_6717);
nor U9976 (N_9976,N_4377,N_5740);
or U9977 (N_9977,N_4943,N_6428);
or U9978 (N_9978,N_7671,N_6999);
nor U9979 (N_9979,N_4452,N_4565);
nand U9980 (N_9980,N_4292,N_7961);
nand U9981 (N_9981,N_5044,N_6432);
nand U9982 (N_9982,N_6130,N_6822);
nand U9983 (N_9983,N_4989,N_6902);
or U9984 (N_9984,N_5283,N_6781);
nand U9985 (N_9985,N_4902,N_7481);
and U9986 (N_9986,N_4428,N_7468);
nand U9987 (N_9987,N_4759,N_6477);
and U9988 (N_9988,N_7523,N_5018);
and U9989 (N_9989,N_6693,N_7301);
nand U9990 (N_9990,N_7588,N_5117);
nand U9991 (N_9991,N_4458,N_7494);
nor U9992 (N_9992,N_5725,N_7254);
nor U9993 (N_9993,N_6655,N_5189);
or U9994 (N_9994,N_7768,N_6758);
nor U9995 (N_9995,N_4232,N_7064);
nand U9996 (N_9996,N_5862,N_4911);
and U9997 (N_9997,N_5933,N_4155);
nand U9998 (N_9998,N_5733,N_4964);
nor U9999 (N_9999,N_7881,N_5648);
or U10000 (N_10000,N_6217,N_7750);
nor U10001 (N_10001,N_7239,N_6438);
or U10002 (N_10002,N_6106,N_7779);
or U10003 (N_10003,N_5708,N_5691);
nor U10004 (N_10004,N_7287,N_7092);
nand U10005 (N_10005,N_6639,N_4604);
or U10006 (N_10006,N_5960,N_6794);
nand U10007 (N_10007,N_4892,N_5440);
nor U10008 (N_10008,N_7205,N_7526);
or U10009 (N_10009,N_7573,N_4762);
or U10010 (N_10010,N_6126,N_7117);
nor U10011 (N_10011,N_5177,N_4767);
and U10012 (N_10012,N_5738,N_4416);
and U10013 (N_10013,N_7984,N_5631);
nor U10014 (N_10014,N_7303,N_4679);
nand U10015 (N_10015,N_6587,N_7830);
nand U10016 (N_10016,N_6192,N_6852);
xnor U10017 (N_10017,N_6851,N_6799);
xnor U10018 (N_10018,N_6840,N_7489);
nor U10019 (N_10019,N_6558,N_4518);
or U10020 (N_10020,N_4923,N_7018);
and U10021 (N_10021,N_7348,N_6744);
nand U10022 (N_10022,N_7302,N_6931);
nor U10023 (N_10023,N_4321,N_6504);
or U10024 (N_10024,N_7217,N_7567);
and U10025 (N_10025,N_4284,N_5828);
and U10026 (N_10026,N_6976,N_5457);
nand U10027 (N_10027,N_7540,N_6011);
or U10028 (N_10028,N_7604,N_5743);
nor U10029 (N_10029,N_6926,N_6694);
or U10030 (N_10030,N_7784,N_7922);
nand U10031 (N_10031,N_5030,N_5137);
nand U10032 (N_10032,N_4802,N_6787);
or U10033 (N_10033,N_7937,N_5650);
nand U10034 (N_10034,N_5436,N_7373);
and U10035 (N_10035,N_4909,N_7865);
nand U10036 (N_10036,N_6684,N_4516);
nor U10037 (N_10037,N_4034,N_4823);
or U10038 (N_10038,N_4472,N_7519);
nand U10039 (N_10039,N_6407,N_6760);
nor U10040 (N_10040,N_5241,N_7496);
nor U10041 (N_10041,N_7912,N_6872);
nand U10042 (N_10042,N_4398,N_7092);
or U10043 (N_10043,N_4125,N_7675);
nand U10044 (N_10044,N_5596,N_7817);
nor U10045 (N_10045,N_4413,N_4760);
nand U10046 (N_10046,N_7342,N_7493);
nor U10047 (N_10047,N_5130,N_6750);
nand U10048 (N_10048,N_6519,N_4261);
nand U10049 (N_10049,N_6593,N_5906);
nor U10050 (N_10050,N_7704,N_7997);
and U10051 (N_10051,N_4401,N_6076);
or U10052 (N_10052,N_7985,N_7587);
nor U10053 (N_10053,N_5227,N_4823);
or U10054 (N_10054,N_6947,N_5786);
or U10055 (N_10055,N_7112,N_7229);
and U10056 (N_10056,N_6876,N_5477);
nand U10057 (N_10057,N_6492,N_7851);
and U10058 (N_10058,N_7647,N_6198);
and U10059 (N_10059,N_6561,N_4335);
and U10060 (N_10060,N_4170,N_7871);
and U10061 (N_10061,N_4990,N_6599);
or U10062 (N_10062,N_5505,N_7091);
nand U10063 (N_10063,N_6673,N_5894);
and U10064 (N_10064,N_7072,N_4935);
nor U10065 (N_10065,N_4254,N_7116);
nand U10066 (N_10066,N_4921,N_7419);
or U10067 (N_10067,N_4337,N_4300);
or U10068 (N_10068,N_7861,N_5094);
nor U10069 (N_10069,N_6016,N_6561);
nor U10070 (N_10070,N_5012,N_5967);
and U10071 (N_10071,N_7268,N_4633);
nand U10072 (N_10072,N_6946,N_6485);
and U10073 (N_10073,N_7253,N_6333);
and U10074 (N_10074,N_6567,N_7820);
nor U10075 (N_10075,N_5558,N_6845);
and U10076 (N_10076,N_6999,N_5602);
or U10077 (N_10077,N_4980,N_5834);
nor U10078 (N_10078,N_7777,N_6701);
and U10079 (N_10079,N_5397,N_6433);
and U10080 (N_10080,N_6755,N_4011);
nor U10081 (N_10081,N_4662,N_5715);
or U10082 (N_10082,N_5163,N_4712);
and U10083 (N_10083,N_4955,N_4414);
nand U10084 (N_10084,N_4526,N_6332);
nor U10085 (N_10085,N_6643,N_5658);
nor U10086 (N_10086,N_4584,N_7082);
nor U10087 (N_10087,N_5844,N_6472);
nor U10088 (N_10088,N_6654,N_7131);
nor U10089 (N_10089,N_6127,N_7054);
or U10090 (N_10090,N_5830,N_4319);
nor U10091 (N_10091,N_5808,N_6928);
nor U10092 (N_10092,N_5759,N_4306);
and U10093 (N_10093,N_5458,N_5343);
nand U10094 (N_10094,N_5746,N_6051);
nor U10095 (N_10095,N_7579,N_7550);
nand U10096 (N_10096,N_7107,N_4885);
nor U10097 (N_10097,N_4874,N_6661);
nand U10098 (N_10098,N_5805,N_7359);
and U10099 (N_10099,N_7433,N_6258);
or U10100 (N_10100,N_7915,N_6310);
xor U10101 (N_10101,N_7150,N_4288);
nand U10102 (N_10102,N_4560,N_4976);
and U10103 (N_10103,N_7740,N_5150);
nand U10104 (N_10104,N_7755,N_6778);
or U10105 (N_10105,N_6844,N_6685);
nor U10106 (N_10106,N_5316,N_5516);
nor U10107 (N_10107,N_4972,N_7603);
or U10108 (N_10108,N_4170,N_6848);
and U10109 (N_10109,N_6970,N_4595);
or U10110 (N_10110,N_7410,N_4801);
nor U10111 (N_10111,N_6892,N_6833);
nor U10112 (N_10112,N_7871,N_5045);
nor U10113 (N_10113,N_4212,N_7957);
nand U10114 (N_10114,N_6569,N_5173);
nand U10115 (N_10115,N_5037,N_5312);
or U10116 (N_10116,N_6170,N_6102);
and U10117 (N_10117,N_6412,N_7841);
or U10118 (N_10118,N_6911,N_6235);
nand U10119 (N_10119,N_6835,N_5098);
nand U10120 (N_10120,N_6300,N_7461);
or U10121 (N_10121,N_5459,N_4589);
and U10122 (N_10122,N_7700,N_6800);
and U10123 (N_10123,N_7981,N_4935);
or U10124 (N_10124,N_6485,N_7478);
nand U10125 (N_10125,N_4436,N_4747);
or U10126 (N_10126,N_5613,N_6528);
or U10127 (N_10127,N_4071,N_5762);
or U10128 (N_10128,N_5432,N_4946);
and U10129 (N_10129,N_7042,N_4781);
and U10130 (N_10130,N_5618,N_6560);
and U10131 (N_10131,N_6193,N_7845);
or U10132 (N_10132,N_6452,N_5974);
nand U10133 (N_10133,N_7587,N_4617);
and U10134 (N_10134,N_5350,N_4397);
and U10135 (N_10135,N_6717,N_7004);
nor U10136 (N_10136,N_4099,N_4594);
and U10137 (N_10137,N_5488,N_7302);
nand U10138 (N_10138,N_4217,N_5401);
or U10139 (N_10139,N_7221,N_6291);
nand U10140 (N_10140,N_7686,N_4898);
xnor U10141 (N_10141,N_6346,N_4960);
nand U10142 (N_10142,N_6574,N_4587);
nor U10143 (N_10143,N_5476,N_4794);
or U10144 (N_10144,N_4949,N_5271);
nand U10145 (N_10145,N_7432,N_5654);
xor U10146 (N_10146,N_6074,N_7393);
nand U10147 (N_10147,N_5646,N_7533);
and U10148 (N_10148,N_6125,N_4062);
or U10149 (N_10149,N_6972,N_6903);
nand U10150 (N_10150,N_6221,N_7045);
and U10151 (N_10151,N_5788,N_4825);
nand U10152 (N_10152,N_5668,N_7587);
nand U10153 (N_10153,N_4324,N_4375);
nor U10154 (N_10154,N_4360,N_4837);
and U10155 (N_10155,N_4688,N_4183);
and U10156 (N_10156,N_7774,N_4704);
or U10157 (N_10157,N_5625,N_7592);
or U10158 (N_10158,N_4392,N_5602);
and U10159 (N_10159,N_7996,N_4064);
nand U10160 (N_10160,N_6331,N_6584);
or U10161 (N_10161,N_5422,N_7153);
and U10162 (N_10162,N_4437,N_4899);
and U10163 (N_10163,N_4673,N_6467);
and U10164 (N_10164,N_6247,N_6729);
or U10165 (N_10165,N_5890,N_4852);
and U10166 (N_10166,N_5523,N_5241);
nand U10167 (N_10167,N_5225,N_6604);
or U10168 (N_10168,N_5389,N_5100);
and U10169 (N_10169,N_5128,N_6937);
and U10170 (N_10170,N_4481,N_5334);
and U10171 (N_10171,N_4929,N_4221);
and U10172 (N_10172,N_6461,N_6540);
nand U10173 (N_10173,N_6325,N_5812);
or U10174 (N_10174,N_5436,N_7464);
or U10175 (N_10175,N_5739,N_5688);
nand U10176 (N_10176,N_5120,N_7724);
nor U10177 (N_10177,N_6085,N_4959);
or U10178 (N_10178,N_6729,N_5060);
nor U10179 (N_10179,N_4523,N_5176);
and U10180 (N_10180,N_7576,N_6935);
or U10181 (N_10181,N_7468,N_4159);
and U10182 (N_10182,N_7269,N_4927);
nand U10183 (N_10183,N_6651,N_4751);
nand U10184 (N_10184,N_4294,N_6119);
or U10185 (N_10185,N_4007,N_4098);
and U10186 (N_10186,N_7052,N_5244);
xor U10187 (N_10187,N_4241,N_7639);
or U10188 (N_10188,N_7151,N_6941);
nand U10189 (N_10189,N_7156,N_7534);
or U10190 (N_10190,N_4362,N_5337);
or U10191 (N_10191,N_4575,N_7130);
or U10192 (N_10192,N_5325,N_4187);
nand U10193 (N_10193,N_5205,N_5524);
or U10194 (N_10194,N_4336,N_6981);
and U10195 (N_10195,N_7253,N_7545);
and U10196 (N_10196,N_4823,N_6789);
nand U10197 (N_10197,N_4725,N_7098);
nor U10198 (N_10198,N_4933,N_7353);
or U10199 (N_10199,N_7714,N_4589);
nor U10200 (N_10200,N_7762,N_5235);
or U10201 (N_10201,N_6509,N_4354);
or U10202 (N_10202,N_4716,N_6668);
nor U10203 (N_10203,N_7334,N_7942);
nor U10204 (N_10204,N_6364,N_7849);
or U10205 (N_10205,N_6915,N_6464);
or U10206 (N_10206,N_6626,N_4811);
nor U10207 (N_10207,N_7953,N_7992);
nor U10208 (N_10208,N_5841,N_4065);
or U10209 (N_10209,N_5629,N_4909);
and U10210 (N_10210,N_7779,N_6959);
nand U10211 (N_10211,N_4584,N_7853);
and U10212 (N_10212,N_6699,N_7025);
nor U10213 (N_10213,N_7311,N_4783);
and U10214 (N_10214,N_7835,N_5926);
nor U10215 (N_10215,N_5355,N_6450);
nand U10216 (N_10216,N_4061,N_5940);
nor U10217 (N_10217,N_5488,N_6959);
nor U10218 (N_10218,N_4865,N_5639);
or U10219 (N_10219,N_4575,N_6121);
or U10220 (N_10220,N_4432,N_7646);
and U10221 (N_10221,N_7003,N_7311);
nand U10222 (N_10222,N_6243,N_6599);
nor U10223 (N_10223,N_6747,N_6814);
nor U10224 (N_10224,N_4085,N_7364);
nand U10225 (N_10225,N_5729,N_5478);
xnor U10226 (N_10226,N_4176,N_7752);
or U10227 (N_10227,N_5144,N_5240);
nand U10228 (N_10228,N_4957,N_4706);
or U10229 (N_10229,N_5173,N_4344);
nor U10230 (N_10230,N_4760,N_5447);
nor U10231 (N_10231,N_7096,N_4684);
and U10232 (N_10232,N_4645,N_6125);
nand U10233 (N_10233,N_7396,N_6498);
and U10234 (N_10234,N_5612,N_5592);
nand U10235 (N_10235,N_6834,N_7302);
or U10236 (N_10236,N_6396,N_4931);
nor U10237 (N_10237,N_4537,N_6266);
or U10238 (N_10238,N_6617,N_7077);
and U10239 (N_10239,N_7147,N_6100);
nor U10240 (N_10240,N_5091,N_5559);
nand U10241 (N_10241,N_5880,N_5819);
and U10242 (N_10242,N_5888,N_4744);
nand U10243 (N_10243,N_7499,N_7341);
and U10244 (N_10244,N_4115,N_5310);
or U10245 (N_10245,N_7127,N_5799);
nor U10246 (N_10246,N_4869,N_7377);
nand U10247 (N_10247,N_6036,N_5624);
or U10248 (N_10248,N_5542,N_4888);
nor U10249 (N_10249,N_6776,N_4376);
nand U10250 (N_10250,N_7936,N_4203);
nand U10251 (N_10251,N_7058,N_6430);
or U10252 (N_10252,N_4154,N_5185);
nor U10253 (N_10253,N_7769,N_4144);
nand U10254 (N_10254,N_6187,N_5751);
or U10255 (N_10255,N_4197,N_4479);
and U10256 (N_10256,N_7392,N_4109);
and U10257 (N_10257,N_7813,N_5413);
or U10258 (N_10258,N_4295,N_7229);
nor U10259 (N_10259,N_6719,N_7703);
and U10260 (N_10260,N_6425,N_6305);
nand U10261 (N_10261,N_6738,N_6393);
or U10262 (N_10262,N_6721,N_5925);
nand U10263 (N_10263,N_4867,N_7481);
or U10264 (N_10264,N_6782,N_5522);
and U10265 (N_10265,N_4328,N_6264);
nor U10266 (N_10266,N_7141,N_7406);
nand U10267 (N_10267,N_4498,N_7652);
and U10268 (N_10268,N_6212,N_4338);
nand U10269 (N_10269,N_7028,N_4798);
nor U10270 (N_10270,N_5569,N_6475);
and U10271 (N_10271,N_6953,N_7697);
and U10272 (N_10272,N_7681,N_4589);
and U10273 (N_10273,N_7077,N_6464);
nor U10274 (N_10274,N_7877,N_5727);
and U10275 (N_10275,N_6621,N_6240);
nor U10276 (N_10276,N_6437,N_6172);
nand U10277 (N_10277,N_5664,N_5779);
or U10278 (N_10278,N_5799,N_7364);
nand U10279 (N_10279,N_5909,N_4892);
and U10280 (N_10280,N_4419,N_6925);
nand U10281 (N_10281,N_4349,N_7152);
and U10282 (N_10282,N_4230,N_4198);
or U10283 (N_10283,N_5437,N_4394);
nand U10284 (N_10284,N_7260,N_7833);
and U10285 (N_10285,N_7046,N_4413);
nand U10286 (N_10286,N_6897,N_7778);
nand U10287 (N_10287,N_4313,N_5966);
nor U10288 (N_10288,N_7211,N_7725);
or U10289 (N_10289,N_5805,N_5034);
nor U10290 (N_10290,N_7668,N_7829);
or U10291 (N_10291,N_5269,N_6408);
or U10292 (N_10292,N_4490,N_4634);
nor U10293 (N_10293,N_6035,N_5514);
nor U10294 (N_10294,N_5949,N_7150);
nor U10295 (N_10295,N_7545,N_7177);
nor U10296 (N_10296,N_7640,N_7006);
nor U10297 (N_10297,N_4245,N_6297);
xnor U10298 (N_10298,N_4130,N_7697);
nand U10299 (N_10299,N_7001,N_5925);
nand U10300 (N_10300,N_5653,N_7444);
nand U10301 (N_10301,N_4147,N_5939);
nand U10302 (N_10302,N_6421,N_5139);
and U10303 (N_10303,N_4736,N_5591);
or U10304 (N_10304,N_5040,N_6153);
and U10305 (N_10305,N_4604,N_5800);
nor U10306 (N_10306,N_7893,N_4958);
nor U10307 (N_10307,N_5526,N_4273);
and U10308 (N_10308,N_6870,N_5537);
nor U10309 (N_10309,N_7736,N_5792);
nand U10310 (N_10310,N_4989,N_5780);
nand U10311 (N_10311,N_5298,N_4488);
nor U10312 (N_10312,N_6362,N_4094);
nand U10313 (N_10313,N_5001,N_4926);
nand U10314 (N_10314,N_4769,N_7220);
or U10315 (N_10315,N_7258,N_6226);
and U10316 (N_10316,N_7449,N_4278);
nor U10317 (N_10317,N_4400,N_6963);
and U10318 (N_10318,N_4341,N_7641);
or U10319 (N_10319,N_5514,N_6854);
nand U10320 (N_10320,N_4556,N_5683);
and U10321 (N_10321,N_5497,N_5290);
and U10322 (N_10322,N_4143,N_7172);
nand U10323 (N_10323,N_5239,N_5363);
nor U10324 (N_10324,N_6598,N_7034);
nand U10325 (N_10325,N_6879,N_4579);
nand U10326 (N_10326,N_7634,N_5635);
nand U10327 (N_10327,N_6439,N_5143);
nor U10328 (N_10328,N_5779,N_4305);
nand U10329 (N_10329,N_5269,N_6755);
or U10330 (N_10330,N_4307,N_7965);
nand U10331 (N_10331,N_6008,N_7848);
or U10332 (N_10332,N_7200,N_6459);
nand U10333 (N_10333,N_4174,N_4642);
or U10334 (N_10334,N_7659,N_4158);
nand U10335 (N_10335,N_4487,N_5049);
and U10336 (N_10336,N_6144,N_6012);
or U10337 (N_10337,N_5260,N_7407);
nand U10338 (N_10338,N_6767,N_6321);
and U10339 (N_10339,N_4133,N_7171);
nand U10340 (N_10340,N_5896,N_4150);
and U10341 (N_10341,N_6740,N_6532);
nor U10342 (N_10342,N_5458,N_4415);
and U10343 (N_10343,N_4265,N_5662);
and U10344 (N_10344,N_7211,N_4062);
nand U10345 (N_10345,N_7527,N_7114);
and U10346 (N_10346,N_6776,N_7292);
or U10347 (N_10347,N_5708,N_6762);
and U10348 (N_10348,N_5850,N_5537);
nor U10349 (N_10349,N_4456,N_6811);
xor U10350 (N_10350,N_6978,N_6084);
nor U10351 (N_10351,N_6418,N_7866);
nor U10352 (N_10352,N_5699,N_4176);
and U10353 (N_10353,N_4211,N_5036);
nor U10354 (N_10354,N_6756,N_5378);
nor U10355 (N_10355,N_4173,N_7408);
or U10356 (N_10356,N_5306,N_6970);
nand U10357 (N_10357,N_6669,N_4287);
nand U10358 (N_10358,N_5074,N_6213);
or U10359 (N_10359,N_5238,N_6691);
or U10360 (N_10360,N_5794,N_4594);
nand U10361 (N_10361,N_5993,N_4031);
and U10362 (N_10362,N_5943,N_4457);
or U10363 (N_10363,N_5301,N_4869);
and U10364 (N_10364,N_4386,N_4260);
and U10365 (N_10365,N_7790,N_7261);
or U10366 (N_10366,N_6364,N_6530);
nand U10367 (N_10367,N_7105,N_6470);
and U10368 (N_10368,N_5965,N_5508);
and U10369 (N_10369,N_6523,N_6985);
nand U10370 (N_10370,N_7820,N_5450);
nand U10371 (N_10371,N_4295,N_5299);
or U10372 (N_10372,N_4801,N_7961);
or U10373 (N_10373,N_4249,N_4482);
nor U10374 (N_10374,N_4411,N_4245);
or U10375 (N_10375,N_7527,N_5950);
nand U10376 (N_10376,N_6565,N_7490);
nand U10377 (N_10377,N_7413,N_7002);
and U10378 (N_10378,N_5597,N_5371);
nand U10379 (N_10379,N_6112,N_7750);
nand U10380 (N_10380,N_7812,N_4348);
and U10381 (N_10381,N_7907,N_7222);
or U10382 (N_10382,N_6272,N_5816);
nand U10383 (N_10383,N_7425,N_4784);
nor U10384 (N_10384,N_7864,N_7488);
and U10385 (N_10385,N_6037,N_7094);
nor U10386 (N_10386,N_7853,N_4866);
nand U10387 (N_10387,N_4215,N_5324);
or U10388 (N_10388,N_4406,N_7550);
or U10389 (N_10389,N_5427,N_5408);
xor U10390 (N_10390,N_7902,N_6320);
and U10391 (N_10391,N_6604,N_6199);
or U10392 (N_10392,N_6946,N_4282);
nand U10393 (N_10393,N_6187,N_7864);
or U10394 (N_10394,N_7852,N_6016);
nor U10395 (N_10395,N_6967,N_5507);
and U10396 (N_10396,N_4611,N_5791);
and U10397 (N_10397,N_7789,N_7916);
and U10398 (N_10398,N_5804,N_6378);
nand U10399 (N_10399,N_7464,N_6745);
and U10400 (N_10400,N_7531,N_7883);
nor U10401 (N_10401,N_6783,N_4958);
or U10402 (N_10402,N_7769,N_7675);
nor U10403 (N_10403,N_4243,N_5217);
nor U10404 (N_10404,N_5579,N_5539);
or U10405 (N_10405,N_7924,N_7860);
and U10406 (N_10406,N_5543,N_4569);
nor U10407 (N_10407,N_5426,N_4115);
and U10408 (N_10408,N_5393,N_4820);
and U10409 (N_10409,N_5993,N_7675);
nand U10410 (N_10410,N_5558,N_7803);
nor U10411 (N_10411,N_6588,N_4368);
nor U10412 (N_10412,N_7486,N_7697);
nor U10413 (N_10413,N_6846,N_7409);
and U10414 (N_10414,N_7451,N_5510);
or U10415 (N_10415,N_6061,N_6748);
nand U10416 (N_10416,N_4810,N_6724);
nand U10417 (N_10417,N_6592,N_4465);
nand U10418 (N_10418,N_4785,N_7771);
or U10419 (N_10419,N_5503,N_7299);
and U10420 (N_10420,N_5168,N_4463);
or U10421 (N_10421,N_4414,N_6367);
nand U10422 (N_10422,N_4675,N_7120);
and U10423 (N_10423,N_7041,N_6906);
nor U10424 (N_10424,N_5864,N_4760);
and U10425 (N_10425,N_4105,N_5619);
nand U10426 (N_10426,N_5626,N_5746);
and U10427 (N_10427,N_6398,N_5053);
nand U10428 (N_10428,N_7640,N_4256);
and U10429 (N_10429,N_4796,N_4340);
or U10430 (N_10430,N_7449,N_4695);
nor U10431 (N_10431,N_5884,N_7768);
or U10432 (N_10432,N_7585,N_4741);
nor U10433 (N_10433,N_5255,N_4262);
nand U10434 (N_10434,N_6971,N_7940);
nand U10435 (N_10435,N_7828,N_6507);
or U10436 (N_10436,N_4615,N_5470);
nand U10437 (N_10437,N_6412,N_6185);
nand U10438 (N_10438,N_7989,N_7174);
or U10439 (N_10439,N_5131,N_6518);
nor U10440 (N_10440,N_4856,N_5157);
nand U10441 (N_10441,N_7350,N_7569);
and U10442 (N_10442,N_4382,N_6511);
nand U10443 (N_10443,N_4103,N_6758);
nand U10444 (N_10444,N_6559,N_6943);
nor U10445 (N_10445,N_4371,N_5610);
nor U10446 (N_10446,N_5910,N_5497);
or U10447 (N_10447,N_7902,N_5766);
nand U10448 (N_10448,N_5781,N_7169);
nor U10449 (N_10449,N_7997,N_5016);
or U10450 (N_10450,N_6765,N_7824);
nand U10451 (N_10451,N_5704,N_6132);
or U10452 (N_10452,N_6795,N_7984);
or U10453 (N_10453,N_4841,N_5589);
nor U10454 (N_10454,N_7573,N_7544);
nand U10455 (N_10455,N_4007,N_6377);
nand U10456 (N_10456,N_7926,N_6046);
nand U10457 (N_10457,N_5281,N_4005);
and U10458 (N_10458,N_4218,N_5129);
and U10459 (N_10459,N_6338,N_7271);
and U10460 (N_10460,N_4099,N_4509);
nand U10461 (N_10461,N_7170,N_6046);
and U10462 (N_10462,N_6649,N_7009);
or U10463 (N_10463,N_6802,N_6761);
xnor U10464 (N_10464,N_5217,N_4174);
and U10465 (N_10465,N_6220,N_5906);
nor U10466 (N_10466,N_5169,N_4262);
nor U10467 (N_10467,N_7127,N_7609);
nor U10468 (N_10468,N_4557,N_4656);
nor U10469 (N_10469,N_4240,N_4209);
and U10470 (N_10470,N_6519,N_7883);
nor U10471 (N_10471,N_7084,N_5852);
or U10472 (N_10472,N_4030,N_7264);
nand U10473 (N_10473,N_5546,N_7234);
xnor U10474 (N_10474,N_6644,N_7486);
nor U10475 (N_10475,N_6068,N_5484);
nand U10476 (N_10476,N_7057,N_4029);
or U10477 (N_10477,N_4929,N_6085);
and U10478 (N_10478,N_5657,N_5866);
nand U10479 (N_10479,N_5440,N_5845);
or U10480 (N_10480,N_5662,N_7414);
nand U10481 (N_10481,N_5931,N_6261);
nor U10482 (N_10482,N_4413,N_5860);
nor U10483 (N_10483,N_4506,N_5104);
or U10484 (N_10484,N_6879,N_7999);
and U10485 (N_10485,N_5277,N_6067);
xor U10486 (N_10486,N_7213,N_4736);
nor U10487 (N_10487,N_5636,N_4843);
nor U10488 (N_10488,N_5618,N_7927);
and U10489 (N_10489,N_4226,N_4049);
or U10490 (N_10490,N_4920,N_6294);
nand U10491 (N_10491,N_6714,N_4957);
nor U10492 (N_10492,N_5696,N_4715);
or U10493 (N_10493,N_5028,N_4382);
nand U10494 (N_10494,N_5793,N_7270);
or U10495 (N_10495,N_5579,N_7091);
nand U10496 (N_10496,N_4585,N_7448);
and U10497 (N_10497,N_5124,N_5264);
nand U10498 (N_10498,N_6600,N_4594);
or U10499 (N_10499,N_4242,N_7016);
and U10500 (N_10500,N_6377,N_5554);
or U10501 (N_10501,N_6605,N_6429);
and U10502 (N_10502,N_4375,N_5494);
and U10503 (N_10503,N_4773,N_6219);
or U10504 (N_10504,N_5478,N_4174);
or U10505 (N_10505,N_6605,N_4289);
and U10506 (N_10506,N_5594,N_6378);
or U10507 (N_10507,N_4110,N_6749);
nor U10508 (N_10508,N_6453,N_6855);
or U10509 (N_10509,N_6333,N_4069);
and U10510 (N_10510,N_7212,N_7219);
nor U10511 (N_10511,N_7861,N_5396);
nor U10512 (N_10512,N_6041,N_4904);
or U10513 (N_10513,N_6617,N_7164);
nor U10514 (N_10514,N_6402,N_6332);
and U10515 (N_10515,N_6338,N_5689);
and U10516 (N_10516,N_6381,N_7424);
and U10517 (N_10517,N_7903,N_6568);
and U10518 (N_10518,N_4751,N_4101);
and U10519 (N_10519,N_7453,N_4183);
and U10520 (N_10520,N_5932,N_6969);
or U10521 (N_10521,N_5826,N_6179);
nor U10522 (N_10522,N_5401,N_4259);
and U10523 (N_10523,N_5486,N_5782);
and U10524 (N_10524,N_4685,N_6139);
nor U10525 (N_10525,N_6254,N_5002);
and U10526 (N_10526,N_4737,N_4376);
nor U10527 (N_10527,N_4350,N_7355);
nor U10528 (N_10528,N_6833,N_4209);
nand U10529 (N_10529,N_6948,N_6559);
or U10530 (N_10530,N_5852,N_7952);
nand U10531 (N_10531,N_6428,N_7344);
xor U10532 (N_10532,N_4930,N_5846);
nand U10533 (N_10533,N_6418,N_4178);
nor U10534 (N_10534,N_7933,N_6366);
and U10535 (N_10535,N_7862,N_5855);
nand U10536 (N_10536,N_4999,N_6353);
nor U10537 (N_10537,N_6356,N_7144);
nor U10538 (N_10538,N_4441,N_7520);
nand U10539 (N_10539,N_7014,N_6387);
nor U10540 (N_10540,N_7873,N_5672);
and U10541 (N_10541,N_6231,N_5883);
and U10542 (N_10542,N_6684,N_6825);
nand U10543 (N_10543,N_7261,N_4557);
nor U10544 (N_10544,N_6011,N_4214);
nand U10545 (N_10545,N_7707,N_4569);
nand U10546 (N_10546,N_6855,N_6260);
or U10547 (N_10547,N_4686,N_4184);
xnor U10548 (N_10548,N_7409,N_6955);
and U10549 (N_10549,N_6288,N_7369);
nor U10550 (N_10550,N_6050,N_4187);
and U10551 (N_10551,N_7911,N_4861);
nand U10552 (N_10552,N_6919,N_4245);
nor U10553 (N_10553,N_4914,N_7231);
and U10554 (N_10554,N_5321,N_6154);
nand U10555 (N_10555,N_6947,N_5679);
nand U10556 (N_10556,N_4740,N_7808);
or U10557 (N_10557,N_7890,N_5201);
nor U10558 (N_10558,N_7229,N_5497);
and U10559 (N_10559,N_6733,N_5344);
or U10560 (N_10560,N_7309,N_4336);
nor U10561 (N_10561,N_4222,N_5001);
nor U10562 (N_10562,N_4198,N_4489);
nor U10563 (N_10563,N_5602,N_5208);
or U10564 (N_10564,N_4084,N_4757);
nor U10565 (N_10565,N_6539,N_6472);
nand U10566 (N_10566,N_4433,N_5790);
nand U10567 (N_10567,N_4301,N_6571);
or U10568 (N_10568,N_6267,N_6460);
nand U10569 (N_10569,N_6542,N_4597);
nand U10570 (N_10570,N_6622,N_7501);
or U10571 (N_10571,N_7129,N_6301);
nor U10572 (N_10572,N_7543,N_4479);
nand U10573 (N_10573,N_7664,N_4689);
or U10574 (N_10574,N_4776,N_6978);
nor U10575 (N_10575,N_6265,N_4904);
nand U10576 (N_10576,N_5212,N_5965);
or U10577 (N_10577,N_5288,N_5467);
nand U10578 (N_10578,N_5351,N_7687);
or U10579 (N_10579,N_5241,N_7688);
and U10580 (N_10580,N_5361,N_5017);
or U10581 (N_10581,N_5337,N_4173);
nor U10582 (N_10582,N_5890,N_7638);
nand U10583 (N_10583,N_7795,N_4264);
nor U10584 (N_10584,N_4277,N_4040);
and U10585 (N_10585,N_4275,N_5381);
xor U10586 (N_10586,N_4676,N_4966);
or U10587 (N_10587,N_5222,N_5172);
nor U10588 (N_10588,N_4796,N_5296);
and U10589 (N_10589,N_4315,N_6723);
nand U10590 (N_10590,N_7219,N_7974);
nand U10591 (N_10591,N_6902,N_7832);
or U10592 (N_10592,N_6692,N_4739);
and U10593 (N_10593,N_5980,N_4038);
nor U10594 (N_10594,N_6917,N_6591);
nor U10595 (N_10595,N_4657,N_4347);
or U10596 (N_10596,N_5915,N_4855);
xnor U10597 (N_10597,N_5574,N_4053);
or U10598 (N_10598,N_7441,N_5124);
and U10599 (N_10599,N_6829,N_5388);
or U10600 (N_10600,N_5924,N_6796);
or U10601 (N_10601,N_5641,N_4757);
and U10602 (N_10602,N_7719,N_6792);
or U10603 (N_10603,N_6537,N_7195);
nor U10604 (N_10604,N_7547,N_5270);
and U10605 (N_10605,N_5318,N_7685);
nand U10606 (N_10606,N_7148,N_5969);
or U10607 (N_10607,N_5708,N_5391);
nor U10608 (N_10608,N_6528,N_6284);
and U10609 (N_10609,N_4877,N_5446);
or U10610 (N_10610,N_4885,N_4431);
and U10611 (N_10611,N_4297,N_5715);
xnor U10612 (N_10612,N_6741,N_4397);
nand U10613 (N_10613,N_5334,N_4574);
nor U10614 (N_10614,N_5486,N_5862);
nor U10615 (N_10615,N_5683,N_5953);
nor U10616 (N_10616,N_6511,N_6076);
nor U10617 (N_10617,N_4703,N_7878);
nand U10618 (N_10618,N_6192,N_7325);
nor U10619 (N_10619,N_4031,N_5637);
nor U10620 (N_10620,N_4792,N_7582);
nor U10621 (N_10621,N_7509,N_4033);
or U10622 (N_10622,N_5606,N_5447);
nand U10623 (N_10623,N_6485,N_5902);
nand U10624 (N_10624,N_5036,N_6842);
nor U10625 (N_10625,N_7296,N_7312);
nand U10626 (N_10626,N_5034,N_6098);
and U10627 (N_10627,N_5855,N_4399);
and U10628 (N_10628,N_7072,N_6688);
and U10629 (N_10629,N_7137,N_5644);
and U10630 (N_10630,N_6663,N_4748);
and U10631 (N_10631,N_5323,N_4484);
nor U10632 (N_10632,N_5387,N_5767);
nor U10633 (N_10633,N_6717,N_4263);
nor U10634 (N_10634,N_6374,N_5861);
and U10635 (N_10635,N_7560,N_4306);
nand U10636 (N_10636,N_7568,N_6747);
nor U10637 (N_10637,N_5712,N_6322);
and U10638 (N_10638,N_6108,N_7409);
nand U10639 (N_10639,N_7768,N_5038);
nand U10640 (N_10640,N_6135,N_4070);
and U10641 (N_10641,N_6751,N_7497);
and U10642 (N_10642,N_6032,N_6527);
nor U10643 (N_10643,N_7751,N_5315);
and U10644 (N_10644,N_7648,N_7424);
or U10645 (N_10645,N_5571,N_4956);
nor U10646 (N_10646,N_7323,N_6978);
nand U10647 (N_10647,N_5853,N_7406);
or U10648 (N_10648,N_6445,N_5622);
and U10649 (N_10649,N_5605,N_6014);
and U10650 (N_10650,N_4503,N_5996);
nor U10651 (N_10651,N_7146,N_7170);
nor U10652 (N_10652,N_4211,N_5228);
and U10653 (N_10653,N_6795,N_4002);
nand U10654 (N_10654,N_5405,N_5187);
or U10655 (N_10655,N_6014,N_4665);
or U10656 (N_10656,N_6697,N_6623);
nor U10657 (N_10657,N_5499,N_4265);
and U10658 (N_10658,N_7859,N_6565);
nor U10659 (N_10659,N_5082,N_5547);
nand U10660 (N_10660,N_6974,N_7809);
or U10661 (N_10661,N_4142,N_4020);
nor U10662 (N_10662,N_4246,N_6720);
and U10663 (N_10663,N_4258,N_5537);
or U10664 (N_10664,N_7800,N_5053);
nor U10665 (N_10665,N_6322,N_5593);
nor U10666 (N_10666,N_7795,N_6963);
nand U10667 (N_10667,N_6111,N_6408);
and U10668 (N_10668,N_6877,N_6517);
or U10669 (N_10669,N_4648,N_7540);
and U10670 (N_10670,N_5761,N_6849);
nor U10671 (N_10671,N_5443,N_4789);
and U10672 (N_10672,N_7139,N_7233);
and U10673 (N_10673,N_7117,N_5123);
nor U10674 (N_10674,N_4516,N_6886);
nor U10675 (N_10675,N_5978,N_7036);
nand U10676 (N_10676,N_5641,N_4603);
nand U10677 (N_10677,N_7344,N_4103);
nand U10678 (N_10678,N_4965,N_6287);
and U10679 (N_10679,N_5456,N_4125);
and U10680 (N_10680,N_6555,N_5944);
or U10681 (N_10681,N_7594,N_6051);
or U10682 (N_10682,N_5974,N_4579);
or U10683 (N_10683,N_5706,N_7072);
or U10684 (N_10684,N_4989,N_4094);
nor U10685 (N_10685,N_4865,N_4160);
nor U10686 (N_10686,N_5351,N_5525);
or U10687 (N_10687,N_5828,N_4627);
nand U10688 (N_10688,N_7481,N_6788);
and U10689 (N_10689,N_4033,N_4889);
nor U10690 (N_10690,N_7381,N_7916);
or U10691 (N_10691,N_6852,N_4551);
nand U10692 (N_10692,N_5200,N_5719);
and U10693 (N_10693,N_7519,N_4938);
nand U10694 (N_10694,N_5204,N_4479);
or U10695 (N_10695,N_4396,N_4442);
nor U10696 (N_10696,N_5582,N_7169);
nor U10697 (N_10697,N_4506,N_7038);
and U10698 (N_10698,N_5780,N_7720);
nor U10699 (N_10699,N_4142,N_6791);
nor U10700 (N_10700,N_7259,N_6295);
and U10701 (N_10701,N_7097,N_7078);
nor U10702 (N_10702,N_5901,N_7486);
and U10703 (N_10703,N_6597,N_5266);
and U10704 (N_10704,N_6232,N_5857);
nand U10705 (N_10705,N_6444,N_4916);
nand U10706 (N_10706,N_4699,N_6522);
or U10707 (N_10707,N_5184,N_4587);
nor U10708 (N_10708,N_4049,N_6530);
and U10709 (N_10709,N_7346,N_6788);
nand U10710 (N_10710,N_6062,N_7878);
or U10711 (N_10711,N_6261,N_7200);
or U10712 (N_10712,N_6580,N_4923);
or U10713 (N_10713,N_7718,N_6131);
nor U10714 (N_10714,N_7545,N_5284);
nor U10715 (N_10715,N_5958,N_4163);
and U10716 (N_10716,N_7995,N_5725);
or U10717 (N_10717,N_7490,N_5988);
or U10718 (N_10718,N_4098,N_4803);
and U10719 (N_10719,N_7617,N_4827);
nor U10720 (N_10720,N_6388,N_6114);
and U10721 (N_10721,N_6309,N_5527);
or U10722 (N_10722,N_6249,N_6565);
and U10723 (N_10723,N_5469,N_7994);
nor U10724 (N_10724,N_4574,N_4955);
and U10725 (N_10725,N_7626,N_6235);
and U10726 (N_10726,N_5163,N_5878);
and U10727 (N_10727,N_4057,N_7727);
nor U10728 (N_10728,N_7608,N_5479);
and U10729 (N_10729,N_4257,N_5617);
nand U10730 (N_10730,N_6898,N_5400);
or U10731 (N_10731,N_6446,N_5883);
nand U10732 (N_10732,N_4542,N_7090);
and U10733 (N_10733,N_5020,N_6671);
and U10734 (N_10734,N_6045,N_4355);
nor U10735 (N_10735,N_5321,N_4247);
and U10736 (N_10736,N_4436,N_6008);
nor U10737 (N_10737,N_7731,N_7696);
nor U10738 (N_10738,N_6260,N_4120);
nor U10739 (N_10739,N_6746,N_4550);
and U10740 (N_10740,N_5448,N_5787);
xnor U10741 (N_10741,N_4894,N_7995);
or U10742 (N_10742,N_7824,N_7673);
and U10743 (N_10743,N_4429,N_6561);
or U10744 (N_10744,N_5736,N_5519);
nor U10745 (N_10745,N_5281,N_6464);
and U10746 (N_10746,N_4643,N_6580);
and U10747 (N_10747,N_7419,N_7051);
or U10748 (N_10748,N_6770,N_7316);
nand U10749 (N_10749,N_7992,N_5018);
xor U10750 (N_10750,N_4062,N_7764);
and U10751 (N_10751,N_4645,N_6741);
or U10752 (N_10752,N_6268,N_5421);
or U10753 (N_10753,N_7352,N_7516);
nor U10754 (N_10754,N_7865,N_7012);
and U10755 (N_10755,N_7939,N_5011);
and U10756 (N_10756,N_4492,N_4543);
and U10757 (N_10757,N_6944,N_5408);
or U10758 (N_10758,N_7503,N_5962);
nand U10759 (N_10759,N_5898,N_7098);
or U10760 (N_10760,N_4354,N_7997);
nor U10761 (N_10761,N_7518,N_7654);
and U10762 (N_10762,N_4371,N_5771);
and U10763 (N_10763,N_7973,N_4928);
nor U10764 (N_10764,N_4886,N_5491);
nor U10765 (N_10765,N_4526,N_7029);
nor U10766 (N_10766,N_5308,N_6182);
or U10767 (N_10767,N_5801,N_5845);
nor U10768 (N_10768,N_5293,N_6355);
nand U10769 (N_10769,N_4520,N_6416);
or U10770 (N_10770,N_6630,N_5380);
and U10771 (N_10771,N_4311,N_7569);
and U10772 (N_10772,N_6105,N_6889);
or U10773 (N_10773,N_5806,N_4386);
xor U10774 (N_10774,N_6508,N_5018);
or U10775 (N_10775,N_5898,N_6912);
nor U10776 (N_10776,N_6070,N_6452);
nor U10777 (N_10777,N_7321,N_7556);
or U10778 (N_10778,N_7880,N_6775);
or U10779 (N_10779,N_4107,N_4703);
xnor U10780 (N_10780,N_6820,N_4836);
xor U10781 (N_10781,N_7963,N_7980);
nor U10782 (N_10782,N_6833,N_7944);
nor U10783 (N_10783,N_4770,N_6092);
and U10784 (N_10784,N_5472,N_6973);
nor U10785 (N_10785,N_7756,N_7138);
nand U10786 (N_10786,N_7858,N_7574);
and U10787 (N_10787,N_4876,N_7404);
nand U10788 (N_10788,N_4593,N_4259);
or U10789 (N_10789,N_7330,N_4446);
or U10790 (N_10790,N_6108,N_7557);
and U10791 (N_10791,N_7542,N_7374);
and U10792 (N_10792,N_4464,N_7771);
and U10793 (N_10793,N_5512,N_4644);
or U10794 (N_10794,N_6834,N_4878);
or U10795 (N_10795,N_7476,N_5283);
and U10796 (N_10796,N_4741,N_6356);
nand U10797 (N_10797,N_4246,N_5906);
nand U10798 (N_10798,N_7971,N_5166);
nand U10799 (N_10799,N_7663,N_4980);
nor U10800 (N_10800,N_7020,N_6585);
nand U10801 (N_10801,N_4663,N_6094);
nor U10802 (N_10802,N_7241,N_7836);
nand U10803 (N_10803,N_4009,N_6140);
and U10804 (N_10804,N_4008,N_5995);
nor U10805 (N_10805,N_4367,N_6408);
and U10806 (N_10806,N_6198,N_6361);
nand U10807 (N_10807,N_7826,N_6926);
nand U10808 (N_10808,N_5776,N_6656);
and U10809 (N_10809,N_4130,N_4393);
and U10810 (N_10810,N_4426,N_5851);
nor U10811 (N_10811,N_4641,N_5920);
nor U10812 (N_10812,N_6743,N_4558);
nand U10813 (N_10813,N_7084,N_4478);
nand U10814 (N_10814,N_6656,N_7962);
and U10815 (N_10815,N_4909,N_7188);
or U10816 (N_10816,N_5852,N_6730);
nand U10817 (N_10817,N_6435,N_5813);
nand U10818 (N_10818,N_5091,N_6622);
xnor U10819 (N_10819,N_4630,N_6743);
nor U10820 (N_10820,N_5854,N_5485);
nor U10821 (N_10821,N_6439,N_4638);
nor U10822 (N_10822,N_7880,N_5241);
and U10823 (N_10823,N_7601,N_6297);
xnor U10824 (N_10824,N_6034,N_5787);
and U10825 (N_10825,N_6671,N_5167);
and U10826 (N_10826,N_5731,N_5529);
nand U10827 (N_10827,N_4016,N_7634);
nand U10828 (N_10828,N_6248,N_6408);
and U10829 (N_10829,N_5977,N_4411);
nor U10830 (N_10830,N_4964,N_6725);
nor U10831 (N_10831,N_4741,N_4598);
nand U10832 (N_10832,N_5602,N_4323);
and U10833 (N_10833,N_7175,N_6099);
nor U10834 (N_10834,N_6236,N_7279);
and U10835 (N_10835,N_4372,N_4962);
and U10836 (N_10836,N_4966,N_7017);
or U10837 (N_10837,N_7294,N_6411);
xor U10838 (N_10838,N_5624,N_4181);
nor U10839 (N_10839,N_7025,N_6963);
and U10840 (N_10840,N_6417,N_6402);
nor U10841 (N_10841,N_5302,N_7742);
nand U10842 (N_10842,N_5539,N_4862);
and U10843 (N_10843,N_6573,N_7258);
nor U10844 (N_10844,N_7610,N_5787);
and U10845 (N_10845,N_5151,N_5944);
xnor U10846 (N_10846,N_6307,N_6761);
and U10847 (N_10847,N_5863,N_7622);
nand U10848 (N_10848,N_7887,N_6705);
nand U10849 (N_10849,N_7138,N_4977);
nand U10850 (N_10850,N_6718,N_4654);
or U10851 (N_10851,N_7023,N_5631);
nor U10852 (N_10852,N_5830,N_6103);
and U10853 (N_10853,N_5024,N_6354);
or U10854 (N_10854,N_7968,N_6863);
and U10855 (N_10855,N_6125,N_4280);
nor U10856 (N_10856,N_6468,N_4902);
or U10857 (N_10857,N_7452,N_4412);
or U10858 (N_10858,N_7513,N_5361);
nor U10859 (N_10859,N_5651,N_7695);
nand U10860 (N_10860,N_4057,N_6976);
or U10861 (N_10861,N_7221,N_6721);
nand U10862 (N_10862,N_7192,N_7865);
nor U10863 (N_10863,N_4889,N_4765);
xnor U10864 (N_10864,N_6539,N_6177);
or U10865 (N_10865,N_6903,N_7223);
or U10866 (N_10866,N_7100,N_7933);
nor U10867 (N_10867,N_6643,N_7053);
nor U10868 (N_10868,N_6244,N_5453);
nand U10869 (N_10869,N_7281,N_5523);
nand U10870 (N_10870,N_4645,N_4341);
or U10871 (N_10871,N_5154,N_4414);
and U10872 (N_10872,N_7849,N_7857);
and U10873 (N_10873,N_6687,N_6106);
nand U10874 (N_10874,N_5820,N_7672);
nand U10875 (N_10875,N_4654,N_6504);
nand U10876 (N_10876,N_7908,N_4128);
or U10877 (N_10877,N_4161,N_7308);
nor U10878 (N_10878,N_7186,N_6007);
or U10879 (N_10879,N_6158,N_5196);
or U10880 (N_10880,N_5640,N_6845);
nand U10881 (N_10881,N_6847,N_7566);
or U10882 (N_10882,N_5903,N_6758);
nor U10883 (N_10883,N_6118,N_5175);
nand U10884 (N_10884,N_6928,N_7419);
xor U10885 (N_10885,N_5930,N_4768);
and U10886 (N_10886,N_6031,N_5689);
and U10887 (N_10887,N_4707,N_4987);
nor U10888 (N_10888,N_6766,N_6944);
or U10889 (N_10889,N_4176,N_6870);
and U10890 (N_10890,N_4749,N_7633);
and U10891 (N_10891,N_7359,N_7150);
nor U10892 (N_10892,N_5056,N_5175);
nand U10893 (N_10893,N_4183,N_5831);
and U10894 (N_10894,N_7827,N_6550);
nand U10895 (N_10895,N_5766,N_5228);
and U10896 (N_10896,N_4925,N_4257);
nand U10897 (N_10897,N_6445,N_7394);
nand U10898 (N_10898,N_4008,N_6336);
nor U10899 (N_10899,N_7349,N_5373);
nand U10900 (N_10900,N_6328,N_4115);
nand U10901 (N_10901,N_6008,N_4956);
nand U10902 (N_10902,N_7754,N_7370);
and U10903 (N_10903,N_4547,N_5786);
or U10904 (N_10904,N_5898,N_4889);
nor U10905 (N_10905,N_6277,N_7639);
nor U10906 (N_10906,N_6197,N_4861);
nand U10907 (N_10907,N_4063,N_4470);
and U10908 (N_10908,N_5591,N_6116);
nand U10909 (N_10909,N_7260,N_4541);
and U10910 (N_10910,N_5677,N_7847);
and U10911 (N_10911,N_4456,N_4284);
nand U10912 (N_10912,N_4983,N_5774);
and U10913 (N_10913,N_7270,N_4859);
nand U10914 (N_10914,N_7958,N_6247);
nand U10915 (N_10915,N_4534,N_4851);
and U10916 (N_10916,N_5473,N_6704);
and U10917 (N_10917,N_4306,N_5570);
nand U10918 (N_10918,N_6518,N_5729);
nor U10919 (N_10919,N_6852,N_4031);
and U10920 (N_10920,N_5852,N_4130);
and U10921 (N_10921,N_4195,N_7999);
nand U10922 (N_10922,N_6079,N_6646);
and U10923 (N_10923,N_4921,N_6775);
nand U10924 (N_10924,N_4123,N_7311);
nand U10925 (N_10925,N_6363,N_5083);
nand U10926 (N_10926,N_5162,N_7884);
nor U10927 (N_10927,N_5308,N_6714);
or U10928 (N_10928,N_6715,N_5056);
nor U10929 (N_10929,N_5679,N_7926);
nand U10930 (N_10930,N_4611,N_6809);
nor U10931 (N_10931,N_5749,N_7684);
nand U10932 (N_10932,N_6853,N_7509);
and U10933 (N_10933,N_4349,N_4675);
or U10934 (N_10934,N_5421,N_5015);
and U10935 (N_10935,N_4532,N_6113);
and U10936 (N_10936,N_7875,N_7296);
nor U10937 (N_10937,N_5681,N_7273);
and U10938 (N_10938,N_6462,N_4639);
xor U10939 (N_10939,N_6915,N_5336);
or U10940 (N_10940,N_4759,N_4946);
nand U10941 (N_10941,N_7788,N_7868);
or U10942 (N_10942,N_6336,N_5288);
nor U10943 (N_10943,N_6687,N_5975);
and U10944 (N_10944,N_5278,N_5789);
nand U10945 (N_10945,N_4888,N_6982);
nor U10946 (N_10946,N_6008,N_6629);
nand U10947 (N_10947,N_6659,N_5803);
or U10948 (N_10948,N_5209,N_7830);
and U10949 (N_10949,N_6829,N_4725);
nor U10950 (N_10950,N_5845,N_4815);
or U10951 (N_10951,N_4431,N_6375);
nor U10952 (N_10952,N_5923,N_7422);
and U10953 (N_10953,N_5111,N_5839);
nor U10954 (N_10954,N_4592,N_4964);
and U10955 (N_10955,N_5051,N_5059);
nand U10956 (N_10956,N_6435,N_4809);
nand U10957 (N_10957,N_7602,N_5596);
nand U10958 (N_10958,N_7595,N_6004);
nand U10959 (N_10959,N_4043,N_7628);
nand U10960 (N_10960,N_4772,N_4958);
nor U10961 (N_10961,N_7844,N_5940);
xnor U10962 (N_10962,N_4634,N_4000);
nor U10963 (N_10963,N_7431,N_7763);
nand U10964 (N_10964,N_6643,N_6948);
or U10965 (N_10965,N_6797,N_4545);
or U10966 (N_10966,N_7822,N_6227);
and U10967 (N_10967,N_6559,N_4890);
and U10968 (N_10968,N_5410,N_6640);
nand U10969 (N_10969,N_6301,N_4868);
nand U10970 (N_10970,N_5449,N_4072);
nand U10971 (N_10971,N_7045,N_4821);
and U10972 (N_10972,N_5858,N_5608);
nand U10973 (N_10973,N_7502,N_4038);
or U10974 (N_10974,N_7238,N_5367);
nand U10975 (N_10975,N_4015,N_5314);
nor U10976 (N_10976,N_7460,N_4093);
and U10977 (N_10977,N_6942,N_5583);
and U10978 (N_10978,N_7143,N_7966);
nand U10979 (N_10979,N_5169,N_7451);
or U10980 (N_10980,N_4394,N_5004);
nand U10981 (N_10981,N_5030,N_5117);
or U10982 (N_10982,N_5369,N_5142);
and U10983 (N_10983,N_6976,N_7552);
and U10984 (N_10984,N_7223,N_4663);
nor U10985 (N_10985,N_7704,N_6178);
or U10986 (N_10986,N_6816,N_5112);
nand U10987 (N_10987,N_6105,N_6740);
nor U10988 (N_10988,N_4591,N_4621);
nor U10989 (N_10989,N_6121,N_4600);
or U10990 (N_10990,N_4665,N_7293);
nor U10991 (N_10991,N_7402,N_4082);
nand U10992 (N_10992,N_4642,N_4147);
or U10993 (N_10993,N_7297,N_6144);
and U10994 (N_10994,N_4132,N_5088);
or U10995 (N_10995,N_5213,N_6785);
xnor U10996 (N_10996,N_5179,N_6045);
and U10997 (N_10997,N_7719,N_4646);
xor U10998 (N_10998,N_5170,N_6816);
nor U10999 (N_10999,N_4348,N_6154);
and U11000 (N_11000,N_6065,N_5605);
nor U11001 (N_11001,N_6235,N_6234);
nor U11002 (N_11002,N_7556,N_5638);
or U11003 (N_11003,N_7797,N_7775);
nor U11004 (N_11004,N_6514,N_4990);
or U11005 (N_11005,N_7581,N_4165);
or U11006 (N_11006,N_4630,N_5187);
nand U11007 (N_11007,N_4691,N_6304);
and U11008 (N_11008,N_4563,N_6865);
and U11009 (N_11009,N_7022,N_7302);
nor U11010 (N_11010,N_6245,N_7562);
and U11011 (N_11011,N_7707,N_7047);
nand U11012 (N_11012,N_4842,N_7506);
or U11013 (N_11013,N_5117,N_4081);
or U11014 (N_11014,N_5155,N_5559);
or U11015 (N_11015,N_4101,N_6745);
nor U11016 (N_11016,N_4567,N_7982);
nor U11017 (N_11017,N_7481,N_7048);
xnor U11018 (N_11018,N_5853,N_5154);
nor U11019 (N_11019,N_4649,N_4845);
nand U11020 (N_11020,N_7381,N_7667);
xor U11021 (N_11021,N_4437,N_6641);
nand U11022 (N_11022,N_5305,N_5100);
and U11023 (N_11023,N_6489,N_5563);
nand U11024 (N_11024,N_5586,N_6754);
nand U11025 (N_11025,N_4705,N_7967);
or U11026 (N_11026,N_4976,N_5002);
or U11027 (N_11027,N_6132,N_7540);
or U11028 (N_11028,N_7796,N_7508);
and U11029 (N_11029,N_5632,N_4596);
nand U11030 (N_11030,N_6607,N_4205);
or U11031 (N_11031,N_4474,N_6341);
nand U11032 (N_11032,N_7501,N_4599);
nor U11033 (N_11033,N_4127,N_7505);
nand U11034 (N_11034,N_6254,N_6372);
or U11035 (N_11035,N_5483,N_6580);
or U11036 (N_11036,N_4540,N_4073);
and U11037 (N_11037,N_7846,N_7781);
nor U11038 (N_11038,N_7334,N_4411);
nand U11039 (N_11039,N_6729,N_6156);
nor U11040 (N_11040,N_5498,N_7454);
nand U11041 (N_11041,N_4738,N_4156);
or U11042 (N_11042,N_6192,N_6506);
and U11043 (N_11043,N_4562,N_4530);
nand U11044 (N_11044,N_6745,N_6936);
nor U11045 (N_11045,N_5382,N_5117);
or U11046 (N_11046,N_6874,N_6155);
nor U11047 (N_11047,N_5617,N_5028);
nand U11048 (N_11048,N_7065,N_5700);
nand U11049 (N_11049,N_4705,N_4068);
nor U11050 (N_11050,N_5841,N_7399);
or U11051 (N_11051,N_6428,N_6756);
and U11052 (N_11052,N_5946,N_5979);
and U11053 (N_11053,N_7037,N_4919);
and U11054 (N_11054,N_7195,N_7207);
nor U11055 (N_11055,N_4170,N_5993);
nand U11056 (N_11056,N_5714,N_5094);
and U11057 (N_11057,N_7025,N_4980);
or U11058 (N_11058,N_4343,N_4154);
and U11059 (N_11059,N_4503,N_7447);
xnor U11060 (N_11060,N_6091,N_5120);
nor U11061 (N_11061,N_4752,N_6022);
nor U11062 (N_11062,N_6788,N_7109);
or U11063 (N_11063,N_7428,N_6865);
or U11064 (N_11064,N_4615,N_5215);
and U11065 (N_11065,N_5198,N_4856);
and U11066 (N_11066,N_6847,N_6387);
xnor U11067 (N_11067,N_6047,N_5366);
nor U11068 (N_11068,N_6064,N_7662);
nand U11069 (N_11069,N_4528,N_6446);
and U11070 (N_11070,N_5186,N_5773);
nand U11071 (N_11071,N_4383,N_4812);
nand U11072 (N_11072,N_5133,N_4005);
nor U11073 (N_11073,N_4469,N_4488);
or U11074 (N_11074,N_5790,N_5478);
or U11075 (N_11075,N_7361,N_7221);
or U11076 (N_11076,N_4638,N_7172);
nor U11077 (N_11077,N_4775,N_7383);
nor U11078 (N_11078,N_4102,N_4078);
and U11079 (N_11079,N_7806,N_5807);
nand U11080 (N_11080,N_4141,N_7069);
and U11081 (N_11081,N_5187,N_7436);
xor U11082 (N_11082,N_6449,N_4198);
nor U11083 (N_11083,N_4134,N_5715);
or U11084 (N_11084,N_7978,N_7380);
nand U11085 (N_11085,N_7617,N_7129);
or U11086 (N_11086,N_7178,N_6934);
or U11087 (N_11087,N_4219,N_5717);
and U11088 (N_11088,N_5273,N_7085);
and U11089 (N_11089,N_7352,N_5021);
nor U11090 (N_11090,N_5307,N_6607);
nand U11091 (N_11091,N_7047,N_5263);
xor U11092 (N_11092,N_5118,N_7605);
nand U11093 (N_11093,N_5527,N_6046);
nor U11094 (N_11094,N_5936,N_7413);
or U11095 (N_11095,N_7235,N_7293);
nand U11096 (N_11096,N_7656,N_4034);
nand U11097 (N_11097,N_7564,N_7878);
or U11098 (N_11098,N_7865,N_7923);
or U11099 (N_11099,N_7544,N_6831);
nor U11100 (N_11100,N_5967,N_4866);
or U11101 (N_11101,N_7203,N_5970);
or U11102 (N_11102,N_4187,N_6442);
nor U11103 (N_11103,N_5783,N_4652);
and U11104 (N_11104,N_5811,N_4239);
nor U11105 (N_11105,N_7897,N_4694);
nand U11106 (N_11106,N_4013,N_4288);
nand U11107 (N_11107,N_7027,N_7881);
and U11108 (N_11108,N_5283,N_7219);
xor U11109 (N_11109,N_6266,N_5668);
xnor U11110 (N_11110,N_7598,N_4432);
or U11111 (N_11111,N_7823,N_6339);
nor U11112 (N_11112,N_4485,N_4045);
nor U11113 (N_11113,N_4756,N_6161);
and U11114 (N_11114,N_6142,N_5605);
nand U11115 (N_11115,N_5813,N_7516);
nand U11116 (N_11116,N_6461,N_4745);
nand U11117 (N_11117,N_7046,N_6657);
or U11118 (N_11118,N_4272,N_7319);
or U11119 (N_11119,N_7763,N_6393);
nand U11120 (N_11120,N_4233,N_5343);
xor U11121 (N_11121,N_6812,N_4759);
nor U11122 (N_11122,N_6169,N_5760);
and U11123 (N_11123,N_7030,N_7417);
nand U11124 (N_11124,N_7026,N_5051);
nand U11125 (N_11125,N_7592,N_5635);
or U11126 (N_11126,N_5469,N_5433);
or U11127 (N_11127,N_6705,N_7934);
nor U11128 (N_11128,N_5451,N_5499);
and U11129 (N_11129,N_4445,N_4752);
and U11130 (N_11130,N_6717,N_7771);
nand U11131 (N_11131,N_5532,N_4425);
or U11132 (N_11132,N_4666,N_7987);
nor U11133 (N_11133,N_4625,N_4578);
or U11134 (N_11134,N_4018,N_5209);
and U11135 (N_11135,N_5800,N_7564);
or U11136 (N_11136,N_5979,N_6100);
or U11137 (N_11137,N_4739,N_6117);
or U11138 (N_11138,N_7025,N_7148);
xnor U11139 (N_11139,N_4763,N_5852);
nor U11140 (N_11140,N_5883,N_4693);
nand U11141 (N_11141,N_5479,N_5930);
nor U11142 (N_11142,N_4578,N_7407);
or U11143 (N_11143,N_4170,N_7179);
or U11144 (N_11144,N_6462,N_4205);
nor U11145 (N_11145,N_6349,N_5612);
and U11146 (N_11146,N_6311,N_4005);
nand U11147 (N_11147,N_6876,N_5451);
nand U11148 (N_11148,N_7619,N_4017);
nand U11149 (N_11149,N_5072,N_6641);
nand U11150 (N_11150,N_4637,N_5301);
and U11151 (N_11151,N_6583,N_4531);
nor U11152 (N_11152,N_4146,N_4884);
or U11153 (N_11153,N_5249,N_7016);
and U11154 (N_11154,N_7282,N_6275);
and U11155 (N_11155,N_6896,N_5623);
and U11156 (N_11156,N_5831,N_6852);
nand U11157 (N_11157,N_4793,N_5561);
or U11158 (N_11158,N_5920,N_5179);
and U11159 (N_11159,N_6941,N_7732);
nor U11160 (N_11160,N_6786,N_4190);
nor U11161 (N_11161,N_5735,N_4745);
nand U11162 (N_11162,N_5345,N_4573);
and U11163 (N_11163,N_6357,N_5371);
nor U11164 (N_11164,N_6412,N_4578);
nand U11165 (N_11165,N_4712,N_5355);
and U11166 (N_11166,N_7206,N_7308);
nand U11167 (N_11167,N_6291,N_4874);
nor U11168 (N_11168,N_7801,N_6680);
nand U11169 (N_11169,N_7666,N_4940);
and U11170 (N_11170,N_5110,N_5235);
and U11171 (N_11171,N_5494,N_4786);
or U11172 (N_11172,N_5678,N_4716);
nor U11173 (N_11173,N_5720,N_6186);
nand U11174 (N_11174,N_5315,N_5032);
and U11175 (N_11175,N_4051,N_6057);
xor U11176 (N_11176,N_7698,N_7355);
nor U11177 (N_11177,N_7933,N_6580);
nand U11178 (N_11178,N_5208,N_5324);
and U11179 (N_11179,N_7607,N_5375);
and U11180 (N_11180,N_6677,N_4201);
xnor U11181 (N_11181,N_6296,N_7607);
and U11182 (N_11182,N_5569,N_4709);
nor U11183 (N_11183,N_7045,N_7346);
and U11184 (N_11184,N_7780,N_6277);
nand U11185 (N_11185,N_4457,N_5964);
and U11186 (N_11186,N_5654,N_7287);
or U11187 (N_11187,N_5777,N_4691);
nand U11188 (N_11188,N_4017,N_7620);
xnor U11189 (N_11189,N_6056,N_4506);
nor U11190 (N_11190,N_6402,N_6320);
nor U11191 (N_11191,N_6420,N_4562);
nor U11192 (N_11192,N_4218,N_6995);
and U11193 (N_11193,N_6863,N_5289);
and U11194 (N_11194,N_4049,N_7080);
or U11195 (N_11195,N_7634,N_7615);
nor U11196 (N_11196,N_7305,N_4579);
nor U11197 (N_11197,N_7290,N_4753);
or U11198 (N_11198,N_5600,N_7122);
nand U11199 (N_11199,N_7611,N_7666);
nand U11200 (N_11200,N_5823,N_4732);
xor U11201 (N_11201,N_6555,N_4116);
and U11202 (N_11202,N_5469,N_7271);
and U11203 (N_11203,N_7011,N_4900);
nor U11204 (N_11204,N_4008,N_4958);
nor U11205 (N_11205,N_6193,N_4978);
or U11206 (N_11206,N_7565,N_7287);
nand U11207 (N_11207,N_4693,N_5036);
nand U11208 (N_11208,N_5824,N_6976);
and U11209 (N_11209,N_7954,N_7485);
and U11210 (N_11210,N_5105,N_4404);
and U11211 (N_11211,N_5694,N_5085);
nor U11212 (N_11212,N_5626,N_4670);
or U11213 (N_11213,N_5429,N_5402);
nand U11214 (N_11214,N_7918,N_5237);
and U11215 (N_11215,N_4799,N_7179);
nand U11216 (N_11216,N_5258,N_6724);
and U11217 (N_11217,N_6319,N_7054);
and U11218 (N_11218,N_7926,N_4796);
nor U11219 (N_11219,N_7219,N_6336);
or U11220 (N_11220,N_4628,N_5607);
nor U11221 (N_11221,N_6771,N_5308);
nor U11222 (N_11222,N_6655,N_4490);
nand U11223 (N_11223,N_5657,N_5479);
and U11224 (N_11224,N_5036,N_7898);
nor U11225 (N_11225,N_4956,N_5808);
or U11226 (N_11226,N_7111,N_7093);
and U11227 (N_11227,N_4035,N_4849);
or U11228 (N_11228,N_6671,N_5441);
and U11229 (N_11229,N_4386,N_6216);
or U11230 (N_11230,N_6223,N_5664);
and U11231 (N_11231,N_7398,N_4661);
nand U11232 (N_11232,N_4913,N_6619);
or U11233 (N_11233,N_7287,N_5129);
or U11234 (N_11234,N_4008,N_6831);
nor U11235 (N_11235,N_6584,N_6346);
nor U11236 (N_11236,N_7520,N_5948);
or U11237 (N_11237,N_5850,N_7137);
nor U11238 (N_11238,N_5312,N_6539);
nor U11239 (N_11239,N_7574,N_4712);
nand U11240 (N_11240,N_5148,N_4688);
and U11241 (N_11241,N_7758,N_7852);
nor U11242 (N_11242,N_5808,N_4893);
and U11243 (N_11243,N_7199,N_5355);
nor U11244 (N_11244,N_5582,N_6351);
nor U11245 (N_11245,N_4426,N_6337);
or U11246 (N_11246,N_5413,N_5749);
or U11247 (N_11247,N_6926,N_7040);
nor U11248 (N_11248,N_7453,N_7121);
nand U11249 (N_11249,N_6195,N_6049);
or U11250 (N_11250,N_4149,N_7099);
and U11251 (N_11251,N_4637,N_7707);
nor U11252 (N_11252,N_6189,N_7001);
and U11253 (N_11253,N_6452,N_4230);
nor U11254 (N_11254,N_6067,N_5338);
and U11255 (N_11255,N_4263,N_7499);
nand U11256 (N_11256,N_5310,N_4641);
and U11257 (N_11257,N_4829,N_5015);
and U11258 (N_11258,N_4849,N_5834);
and U11259 (N_11259,N_4989,N_6823);
nand U11260 (N_11260,N_6569,N_6852);
and U11261 (N_11261,N_7727,N_7887);
and U11262 (N_11262,N_4846,N_7382);
and U11263 (N_11263,N_6208,N_6506);
nand U11264 (N_11264,N_5966,N_6615);
and U11265 (N_11265,N_6567,N_6023);
and U11266 (N_11266,N_4379,N_7864);
nand U11267 (N_11267,N_6659,N_5569);
nand U11268 (N_11268,N_5490,N_5088);
and U11269 (N_11269,N_5910,N_5328);
and U11270 (N_11270,N_7136,N_7179);
and U11271 (N_11271,N_5048,N_7980);
xnor U11272 (N_11272,N_7615,N_5968);
xnor U11273 (N_11273,N_6591,N_4825);
xor U11274 (N_11274,N_5293,N_5572);
nor U11275 (N_11275,N_5114,N_4718);
nor U11276 (N_11276,N_4644,N_6221);
nor U11277 (N_11277,N_7001,N_6481);
or U11278 (N_11278,N_5950,N_6046);
nand U11279 (N_11279,N_6009,N_4982);
nor U11280 (N_11280,N_7334,N_4950);
or U11281 (N_11281,N_6942,N_5035);
nor U11282 (N_11282,N_7199,N_6848);
or U11283 (N_11283,N_7128,N_5646);
nor U11284 (N_11284,N_4020,N_7977);
nor U11285 (N_11285,N_5984,N_7265);
and U11286 (N_11286,N_6145,N_4307);
nor U11287 (N_11287,N_4639,N_6968);
and U11288 (N_11288,N_7509,N_6916);
nand U11289 (N_11289,N_5288,N_7265);
and U11290 (N_11290,N_7424,N_6810);
nand U11291 (N_11291,N_5871,N_7509);
or U11292 (N_11292,N_5447,N_5139);
and U11293 (N_11293,N_5091,N_5871);
and U11294 (N_11294,N_6779,N_6590);
nand U11295 (N_11295,N_7875,N_5800);
nor U11296 (N_11296,N_6358,N_5418);
and U11297 (N_11297,N_6451,N_6991);
nor U11298 (N_11298,N_4297,N_7862);
xor U11299 (N_11299,N_6637,N_4652);
nand U11300 (N_11300,N_4219,N_6121);
or U11301 (N_11301,N_7013,N_5316);
or U11302 (N_11302,N_6259,N_7920);
or U11303 (N_11303,N_4028,N_5460);
nor U11304 (N_11304,N_5805,N_4317);
nor U11305 (N_11305,N_6474,N_5783);
or U11306 (N_11306,N_7743,N_7301);
nor U11307 (N_11307,N_5654,N_4690);
and U11308 (N_11308,N_7651,N_5713);
xor U11309 (N_11309,N_7215,N_5090);
nor U11310 (N_11310,N_6878,N_4679);
nand U11311 (N_11311,N_5265,N_7256);
or U11312 (N_11312,N_7047,N_6035);
nor U11313 (N_11313,N_5160,N_7110);
or U11314 (N_11314,N_7358,N_7794);
and U11315 (N_11315,N_4758,N_6557);
nor U11316 (N_11316,N_6532,N_5386);
nand U11317 (N_11317,N_6590,N_6430);
nand U11318 (N_11318,N_6866,N_7194);
xor U11319 (N_11319,N_7302,N_5295);
xnor U11320 (N_11320,N_7043,N_4835);
nand U11321 (N_11321,N_7777,N_4220);
nor U11322 (N_11322,N_7203,N_4593);
nand U11323 (N_11323,N_4895,N_6068);
or U11324 (N_11324,N_6799,N_7419);
nor U11325 (N_11325,N_5624,N_6462);
nand U11326 (N_11326,N_5613,N_5656);
nand U11327 (N_11327,N_6554,N_7104);
nand U11328 (N_11328,N_7511,N_5323);
nand U11329 (N_11329,N_7979,N_4087);
and U11330 (N_11330,N_4070,N_5680);
xnor U11331 (N_11331,N_5726,N_5045);
nand U11332 (N_11332,N_4318,N_7252);
and U11333 (N_11333,N_6439,N_4831);
and U11334 (N_11334,N_7624,N_4262);
nor U11335 (N_11335,N_4098,N_5886);
nand U11336 (N_11336,N_4212,N_7006);
or U11337 (N_11337,N_4312,N_5840);
and U11338 (N_11338,N_4553,N_5214);
nor U11339 (N_11339,N_5288,N_7963);
or U11340 (N_11340,N_7161,N_5307);
and U11341 (N_11341,N_5420,N_6042);
or U11342 (N_11342,N_5104,N_7055);
or U11343 (N_11343,N_4783,N_4458);
nor U11344 (N_11344,N_6094,N_7454);
nand U11345 (N_11345,N_7703,N_7915);
nor U11346 (N_11346,N_4665,N_4685);
nand U11347 (N_11347,N_7721,N_5381);
nand U11348 (N_11348,N_6579,N_4777);
xor U11349 (N_11349,N_6762,N_5102);
and U11350 (N_11350,N_7724,N_6402);
or U11351 (N_11351,N_5296,N_4496);
nor U11352 (N_11352,N_5448,N_7440);
and U11353 (N_11353,N_7152,N_6697);
nor U11354 (N_11354,N_5550,N_4217);
or U11355 (N_11355,N_6924,N_5287);
nor U11356 (N_11356,N_5546,N_6127);
nand U11357 (N_11357,N_6623,N_6144);
and U11358 (N_11358,N_7190,N_7466);
xor U11359 (N_11359,N_7760,N_7554);
or U11360 (N_11360,N_4288,N_4817);
xnor U11361 (N_11361,N_7160,N_5097);
nor U11362 (N_11362,N_6369,N_4324);
or U11363 (N_11363,N_7372,N_6845);
or U11364 (N_11364,N_5774,N_6188);
nor U11365 (N_11365,N_6489,N_7929);
and U11366 (N_11366,N_7988,N_7295);
and U11367 (N_11367,N_7330,N_5361);
or U11368 (N_11368,N_6382,N_5305);
and U11369 (N_11369,N_6881,N_5526);
nor U11370 (N_11370,N_4493,N_6793);
or U11371 (N_11371,N_4749,N_7735);
nand U11372 (N_11372,N_5725,N_4196);
or U11373 (N_11373,N_5215,N_5546);
and U11374 (N_11374,N_5911,N_7547);
or U11375 (N_11375,N_7298,N_6058);
and U11376 (N_11376,N_6602,N_7194);
and U11377 (N_11377,N_7796,N_4766);
nor U11378 (N_11378,N_7221,N_6608);
nand U11379 (N_11379,N_6951,N_6273);
nor U11380 (N_11380,N_4647,N_6213);
or U11381 (N_11381,N_6227,N_5028);
nor U11382 (N_11382,N_5498,N_5260);
or U11383 (N_11383,N_4798,N_5696);
nor U11384 (N_11384,N_7641,N_5633);
xor U11385 (N_11385,N_6276,N_6692);
or U11386 (N_11386,N_5852,N_5811);
xnor U11387 (N_11387,N_7291,N_7112);
or U11388 (N_11388,N_7731,N_7830);
nand U11389 (N_11389,N_6763,N_6896);
or U11390 (N_11390,N_4642,N_6355);
or U11391 (N_11391,N_4552,N_5244);
nor U11392 (N_11392,N_6899,N_5311);
nor U11393 (N_11393,N_6432,N_7076);
nand U11394 (N_11394,N_5940,N_6285);
nand U11395 (N_11395,N_4050,N_5754);
nand U11396 (N_11396,N_6825,N_6875);
and U11397 (N_11397,N_6602,N_5544);
and U11398 (N_11398,N_5152,N_6191);
nor U11399 (N_11399,N_4808,N_7095);
nand U11400 (N_11400,N_5171,N_5076);
and U11401 (N_11401,N_4899,N_5521);
nand U11402 (N_11402,N_4537,N_7536);
and U11403 (N_11403,N_4151,N_6085);
nor U11404 (N_11404,N_5940,N_4350);
nor U11405 (N_11405,N_5355,N_4665);
nand U11406 (N_11406,N_6637,N_4923);
nor U11407 (N_11407,N_7834,N_4048);
and U11408 (N_11408,N_4704,N_6824);
or U11409 (N_11409,N_7708,N_5494);
xor U11410 (N_11410,N_6635,N_6070);
nand U11411 (N_11411,N_5275,N_4589);
and U11412 (N_11412,N_7181,N_5605);
and U11413 (N_11413,N_4109,N_7050);
nand U11414 (N_11414,N_7956,N_7488);
xor U11415 (N_11415,N_4146,N_7484);
or U11416 (N_11416,N_5733,N_5570);
or U11417 (N_11417,N_5232,N_7386);
or U11418 (N_11418,N_7606,N_5510);
and U11419 (N_11419,N_7660,N_4799);
and U11420 (N_11420,N_6092,N_5352);
nor U11421 (N_11421,N_7825,N_4304);
nand U11422 (N_11422,N_7014,N_6907);
or U11423 (N_11423,N_4592,N_7321);
or U11424 (N_11424,N_7292,N_6919);
or U11425 (N_11425,N_6247,N_5890);
nand U11426 (N_11426,N_6251,N_6970);
or U11427 (N_11427,N_5737,N_7071);
nand U11428 (N_11428,N_6353,N_6360);
nor U11429 (N_11429,N_4384,N_7704);
or U11430 (N_11430,N_4380,N_6794);
nand U11431 (N_11431,N_7734,N_4423);
nor U11432 (N_11432,N_6116,N_4530);
or U11433 (N_11433,N_5787,N_5638);
or U11434 (N_11434,N_7369,N_4086);
and U11435 (N_11435,N_5537,N_5973);
nand U11436 (N_11436,N_4788,N_7682);
nand U11437 (N_11437,N_5091,N_4835);
nand U11438 (N_11438,N_4853,N_7878);
nand U11439 (N_11439,N_4933,N_6271);
xor U11440 (N_11440,N_7105,N_4695);
and U11441 (N_11441,N_5112,N_5070);
or U11442 (N_11442,N_4999,N_4077);
nor U11443 (N_11443,N_7746,N_7806);
nand U11444 (N_11444,N_5711,N_4701);
and U11445 (N_11445,N_6635,N_6884);
nand U11446 (N_11446,N_7179,N_6521);
nand U11447 (N_11447,N_6732,N_4915);
and U11448 (N_11448,N_7277,N_6122);
nor U11449 (N_11449,N_6963,N_5104);
and U11450 (N_11450,N_7256,N_7106);
nor U11451 (N_11451,N_7085,N_4289);
nor U11452 (N_11452,N_6331,N_6035);
nand U11453 (N_11453,N_7873,N_6323);
nor U11454 (N_11454,N_5998,N_4314);
and U11455 (N_11455,N_7424,N_6543);
or U11456 (N_11456,N_5222,N_4019);
nor U11457 (N_11457,N_7910,N_6785);
nor U11458 (N_11458,N_7617,N_6449);
nand U11459 (N_11459,N_5121,N_5539);
and U11460 (N_11460,N_5208,N_4007);
nor U11461 (N_11461,N_7425,N_6854);
nor U11462 (N_11462,N_4874,N_7651);
nand U11463 (N_11463,N_7877,N_4621);
or U11464 (N_11464,N_5882,N_4129);
and U11465 (N_11465,N_6556,N_6700);
or U11466 (N_11466,N_6752,N_5164);
nand U11467 (N_11467,N_5464,N_4053);
nor U11468 (N_11468,N_7187,N_7543);
or U11469 (N_11469,N_4896,N_5008);
nand U11470 (N_11470,N_4597,N_6825);
nor U11471 (N_11471,N_5842,N_6157);
and U11472 (N_11472,N_4276,N_4343);
nor U11473 (N_11473,N_6370,N_5925);
and U11474 (N_11474,N_4989,N_4337);
nand U11475 (N_11475,N_7581,N_7488);
nand U11476 (N_11476,N_6375,N_6606);
nand U11477 (N_11477,N_5528,N_4726);
nand U11478 (N_11478,N_7676,N_5058);
and U11479 (N_11479,N_7963,N_4495);
and U11480 (N_11480,N_7903,N_4901);
and U11481 (N_11481,N_6428,N_6446);
nor U11482 (N_11482,N_5542,N_7112);
nor U11483 (N_11483,N_7816,N_6689);
nor U11484 (N_11484,N_6782,N_4085);
nand U11485 (N_11485,N_5706,N_5495);
and U11486 (N_11486,N_5375,N_7742);
nand U11487 (N_11487,N_7625,N_5299);
xor U11488 (N_11488,N_7678,N_6407);
nand U11489 (N_11489,N_4725,N_4997);
or U11490 (N_11490,N_4202,N_6658);
nand U11491 (N_11491,N_5906,N_7769);
nand U11492 (N_11492,N_4312,N_5866);
nor U11493 (N_11493,N_4925,N_7705);
nor U11494 (N_11494,N_5427,N_7178);
or U11495 (N_11495,N_4507,N_6765);
nand U11496 (N_11496,N_7325,N_6881);
or U11497 (N_11497,N_7416,N_5347);
xor U11498 (N_11498,N_6416,N_4290);
nor U11499 (N_11499,N_4512,N_5123);
nor U11500 (N_11500,N_5425,N_6299);
or U11501 (N_11501,N_7814,N_7587);
nor U11502 (N_11502,N_4066,N_4059);
nand U11503 (N_11503,N_6085,N_5331);
and U11504 (N_11504,N_7564,N_7615);
nor U11505 (N_11505,N_4861,N_4077);
or U11506 (N_11506,N_5376,N_4994);
nand U11507 (N_11507,N_6559,N_4161);
nand U11508 (N_11508,N_7521,N_5565);
and U11509 (N_11509,N_4959,N_5891);
nand U11510 (N_11510,N_5792,N_7325);
and U11511 (N_11511,N_5282,N_5440);
nor U11512 (N_11512,N_4013,N_6664);
nand U11513 (N_11513,N_5198,N_4218);
nor U11514 (N_11514,N_7447,N_5147);
and U11515 (N_11515,N_7655,N_7993);
or U11516 (N_11516,N_6289,N_7511);
or U11517 (N_11517,N_6409,N_6358);
nor U11518 (N_11518,N_5524,N_5579);
or U11519 (N_11519,N_7480,N_5109);
and U11520 (N_11520,N_5582,N_5581);
or U11521 (N_11521,N_7231,N_5781);
and U11522 (N_11522,N_4817,N_6282);
or U11523 (N_11523,N_6847,N_4110);
and U11524 (N_11524,N_5976,N_6806);
and U11525 (N_11525,N_5538,N_5412);
xor U11526 (N_11526,N_4824,N_4992);
and U11527 (N_11527,N_4422,N_7894);
nor U11528 (N_11528,N_6701,N_7716);
nand U11529 (N_11529,N_5238,N_6242);
or U11530 (N_11530,N_4204,N_7853);
or U11531 (N_11531,N_6671,N_5572);
nor U11532 (N_11532,N_7191,N_6640);
nor U11533 (N_11533,N_6386,N_4606);
and U11534 (N_11534,N_4916,N_4923);
nand U11535 (N_11535,N_7467,N_7583);
nand U11536 (N_11536,N_4370,N_5988);
and U11537 (N_11537,N_7882,N_5579);
or U11538 (N_11538,N_7104,N_5057);
nand U11539 (N_11539,N_4820,N_6804);
and U11540 (N_11540,N_6273,N_5558);
or U11541 (N_11541,N_4682,N_5629);
xnor U11542 (N_11542,N_6676,N_5250);
nor U11543 (N_11543,N_7207,N_4049);
nor U11544 (N_11544,N_7791,N_4959);
nand U11545 (N_11545,N_5900,N_7816);
and U11546 (N_11546,N_5724,N_6672);
or U11547 (N_11547,N_4232,N_4847);
nand U11548 (N_11548,N_5114,N_4898);
or U11549 (N_11549,N_4240,N_4321);
or U11550 (N_11550,N_5461,N_4801);
nor U11551 (N_11551,N_5460,N_6652);
or U11552 (N_11552,N_6916,N_5091);
nand U11553 (N_11553,N_7370,N_7385);
or U11554 (N_11554,N_5319,N_5836);
nor U11555 (N_11555,N_6131,N_6725);
nor U11556 (N_11556,N_4902,N_7050);
and U11557 (N_11557,N_7383,N_7313);
nor U11558 (N_11558,N_5520,N_7415);
nor U11559 (N_11559,N_5890,N_7382);
nand U11560 (N_11560,N_6596,N_7301);
or U11561 (N_11561,N_6962,N_7681);
nand U11562 (N_11562,N_5147,N_6102);
and U11563 (N_11563,N_5570,N_4346);
or U11564 (N_11564,N_7463,N_6979);
or U11565 (N_11565,N_4801,N_6635);
nor U11566 (N_11566,N_5928,N_6853);
or U11567 (N_11567,N_5664,N_7847);
nor U11568 (N_11568,N_6384,N_4669);
nor U11569 (N_11569,N_6549,N_5984);
nor U11570 (N_11570,N_4517,N_6584);
and U11571 (N_11571,N_6612,N_4272);
nor U11572 (N_11572,N_4148,N_6151);
and U11573 (N_11573,N_5494,N_7174);
nor U11574 (N_11574,N_4486,N_5156);
and U11575 (N_11575,N_7633,N_4700);
nand U11576 (N_11576,N_4792,N_7859);
nor U11577 (N_11577,N_6683,N_5576);
nand U11578 (N_11578,N_4677,N_5522);
or U11579 (N_11579,N_5717,N_4726);
and U11580 (N_11580,N_6924,N_6365);
nand U11581 (N_11581,N_5675,N_4698);
and U11582 (N_11582,N_7269,N_6709);
and U11583 (N_11583,N_4775,N_6293);
or U11584 (N_11584,N_4076,N_4375);
nor U11585 (N_11585,N_5961,N_5782);
nor U11586 (N_11586,N_5601,N_7233);
nor U11587 (N_11587,N_7775,N_6012);
and U11588 (N_11588,N_6116,N_4212);
nand U11589 (N_11589,N_5136,N_6752);
or U11590 (N_11590,N_7136,N_7738);
nand U11591 (N_11591,N_5793,N_4613);
or U11592 (N_11592,N_7608,N_5569);
nor U11593 (N_11593,N_7326,N_6618);
and U11594 (N_11594,N_4572,N_6382);
or U11595 (N_11595,N_4660,N_4489);
nor U11596 (N_11596,N_5673,N_6779);
nor U11597 (N_11597,N_7481,N_7662);
xor U11598 (N_11598,N_4327,N_6746);
and U11599 (N_11599,N_7717,N_4271);
nand U11600 (N_11600,N_5119,N_7340);
or U11601 (N_11601,N_6560,N_5559);
nand U11602 (N_11602,N_6939,N_5773);
and U11603 (N_11603,N_4505,N_7937);
and U11604 (N_11604,N_5243,N_6575);
or U11605 (N_11605,N_6705,N_4647);
nor U11606 (N_11606,N_5382,N_6631);
nand U11607 (N_11607,N_7706,N_6037);
xnor U11608 (N_11608,N_5523,N_7790);
xor U11609 (N_11609,N_6753,N_5263);
and U11610 (N_11610,N_4002,N_7115);
nor U11611 (N_11611,N_4397,N_4558);
or U11612 (N_11612,N_4327,N_6800);
and U11613 (N_11613,N_7683,N_7002);
nor U11614 (N_11614,N_5282,N_7726);
nor U11615 (N_11615,N_6087,N_7228);
nor U11616 (N_11616,N_7911,N_6215);
or U11617 (N_11617,N_6557,N_4960);
or U11618 (N_11618,N_5146,N_7323);
or U11619 (N_11619,N_7645,N_5792);
or U11620 (N_11620,N_6531,N_5164);
nand U11621 (N_11621,N_4421,N_7909);
and U11622 (N_11622,N_5342,N_7577);
nor U11623 (N_11623,N_5243,N_6254);
or U11624 (N_11624,N_7375,N_7737);
and U11625 (N_11625,N_6468,N_7649);
nand U11626 (N_11626,N_6445,N_6239);
or U11627 (N_11627,N_4498,N_5908);
nor U11628 (N_11628,N_7514,N_6646);
nand U11629 (N_11629,N_4497,N_5432);
or U11630 (N_11630,N_7167,N_6294);
nand U11631 (N_11631,N_7511,N_4920);
nor U11632 (N_11632,N_5297,N_5709);
and U11633 (N_11633,N_7839,N_7774);
and U11634 (N_11634,N_6661,N_5073);
nor U11635 (N_11635,N_5995,N_6438);
nand U11636 (N_11636,N_7868,N_6516);
and U11637 (N_11637,N_7779,N_4111);
and U11638 (N_11638,N_5155,N_7163);
nand U11639 (N_11639,N_6802,N_4897);
and U11640 (N_11640,N_4817,N_5214);
nor U11641 (N_11641,N_5889,N_6203);
and U11642 (N_11642,N_6146,N_7509);
and U11643 (N_11643,N_7500,N_5809);
xor U11644 (N_11644,N_4869,N_6619);
nor U11645 (N_11645,N_5496,N_4859);
or U11646 (N_11646,N_7252,N_7714);
nand U11647 (N_11647,N_4506,N_5761);
nor U11648 (N_11648,N_6399,N_5215);
nand U11649 (N_11649,N_6686,N_6931);
or U11650 (N_11650,N_4771,N_6168);
or U11651 (N_11651,N_4702,N_6681);
and U11652 (N_11652,N_7763,N_4176);
nand U11653 (N_11653,N_6172,N_5822);
or U11654 (N_11654,N_4756,N_5999);
or U11655 (N_11655,N_7415,N_5048);
or U11656 (N_11656,N_4029,N_7241);
and U11657 (N_11657,N_5777,N_4738);
xnor U11658 (N_11658,N_6895,N_6853);
nand U11659 (N_11659,N_4951,N_4532);
or U11660 (N_11660,N_5135,N_6124);
nand U11661 (N_11661,N_4337,N_5440);
nand U11662 (N_11662,N_5321,N_5864);
nand U11663 (N_11663,N_5162,N_6562);
nand U11664 (N_11664,N_4923,N_5092);
nor U11665 (N_11665,N_4656,N_7858);
nor U11666 (N_11666,N_5225,N_7437);
nor U11667 (N_11667,N_7135,N_4341);
and U11668 (N_11668,N_7189,N_7403);
or U11669 (N_11669,N_7089,N_6938);
nand U11670 (N_11670,N_6019,N_6547);
nand U11671 (N_11671,N_5245,N_6881);
xor U11672 (N_11672,N_7959,N_5458);
or U11673 (N_11673,N_5121,N_7938);
or U11674 (N_11674,N_5484,N_6091);
nand U11675 (N_11675,N_4333,N_4997);
nor U11676 (N_11676,N_6258,N_5825);
or U11677 (N_11677,N_7191,N_7541);
or U11678 (N_11678,N_4292,N_4956);
nor U11679 (N_11679,N_7725,N_4910);
nor U11680 (N_11680,N_4437,N_7468);
or U11681 (N_11681,N_6897,N_7857);
or U11682 (N_11682,N_6629,N_5916);
and U11683 (N_11683,N_6143,N_6371);
nor U11684 (N_11684,N_4539,N_5243);
nand U11685 (N_11685,N_5805,N_7966);
nor U11686 (N_11686,N_7758,N_5742);
or U11687 (N_11687,N_4528,N_4134);
nand U11688 (N_11688,N_4070,N_5113);
nand U11689 (N_11689,N_4009,N_7858);
nand U11690 (N_11690,N_5156,N_5044);
nor U11691 (N_11691,N_5249,N_7781);
and U11692 (N_11692,N_6449,N_5542);
nor U11693 (N_11693,N_5864,N_5349);
or U11694 (N_11694,N_6459,N_5982);
nor U11695 (N_11695,N_6923,N_6135);
nand U11696 (N_11696,N_4509,N_4664);
or U11697 (N_11697,N_6192,N_6994);
xnor U11698 (N_11698,N_6023,N_7751);
nor U11699 (N_11699,N_5100,N_5483);
nand U11700 (N_11700,N_6893,N_4811);
nor U11701 (N_11701,N_5839,N_4033);
and U11702 (N_11702,N_5928,N_4918);
or U11703 (N_11703,N_5900,N_5093);
and U11704 (N_11704,N_4344,N_7068);
nand U11705 (N_11705,N_4296,N_6264);
xor U11706 (N_11706,N_5615,N_4623);
nor U11707 (N_11707,N_4830,N_7103);
and U11708 (N_11708,N_6394,N_7510);
nand U11709 (N_11709,N_6882,N_4473);
nor U11710 (N_11710,N_6032,N_5764);
and U11711 (N_11711,N_5734,N_7775);
and U11712 (N_11712,N_4542,N_5568);
and U11713 (N_11713,N_5633,N_6288);
nand U11714 (N_11714,N_6677,N_6334);
or U11715 (N_11715,N_6250,N_7475);
and U11716 (N_11716,N_5484,N_4748);
xor U11717 (N_11717,N_4242,N_5015);
and U11718 (N_11718,N_5114,N_5619);
or U11719 (N_11719,N_6323,N_7220);
nand U11720 (N_11720,N_4777,N_6054);
nor U11721 (N_11721,N_5192,N_7563);
nand U11722 (N_11722,N_6269,N_4922);
or U11723 (N_11723,N_6567,N_6047);
xnor U11724 (N_11724,N_5122,N_7448);
and U11725 (N_11725,N_7447,N_6031);
or U11726 (N_11726,N_7121,N_4590);
nor U11727 (N_11727,N_4431,N_6981);
or U11728 (N_11728,N_5438,N_5887);
nand U11729 (N_11729,N_6116,N_7311);
nor U11730 (N_11730,N_7401,N_7146);
or U11731 (N_11731,N_4046,N_7933);
and U11732 (N_11732,N_5993,N_4422);
and U11733 (N_11733,N_6233,N_5758);
nor U11734 (N_11734,N_6797,N_4484);
nand U11735 (N_11735,N_7101,N_7146);
nor U11736 (N_11736,N_4575,N_4673);
and U11737 (N_11737,N_4566,N_5583);
nor U11738 (N_11738,N_6510,N_6346);
or U11739 (N_11739,N_7639,N_4305);
nor U11740 (N_11740,N_5989,N_5769);
nand U11741 (N_11741,N_7587,N_6386);
nand U11742 (N_11742,N_7219,N_4652);
nor U11743 (N_11743,N_5886,N_4674);
or U11744 (N_11744,N_5889,N_7037);
and U11745 (N_11745,N_7431,N_7642);
nand U11746 (N_11746,N_7338,N_4152);
nor U11747 (N_11747,N_5192,N_7748);
nand U11748 (N_11748,N_4105,N_5607);
nor U11749 (N_11749,N_7631,N_7766);
nand U11750 (N_11750,N_4600,N_5966);
xnor U11751 (N_11751,N_7857,N_7055);
or U11752 (N_11752,N_4203,N_4091);
and U11753 (N_11753,N_7698,N_7864);
nand U11754 (N_11754,N_5680,N_7428);
nand U11755 (N_11755,N_5434,N_6820);
nor U11756 (N_11756,N_7303,N_4410);
nand U11757 (N_11757,N_6642,N_6321);
or U11758 (N_11758,N_6298,N_6234);
or U11759 (N_11759,N_4074,N_6252);
nor U11760 (N_11760,N_4563,N_7894);
or U11761 (N_11761,N_7209,N_4285);
nand U11762 (N_11762,N_7476,N_6441);
or U11763 (N_11763,N_4302,N_7614);
nand U11764 (N_11764,N_6104,N_6536);
or U11765 (N_11765,N_5549,N_4207);
and U11766 (N_11766,N_5427,N_7068);
or U11767 (N_11767,N_5510,N_4115);
nand U11768 (N_11768,N_4750,N_6341);
or U11769 (N_11769,N_4795,N_4034);
nor U11770 (N_11770,N_4357,N_6718);
or U11771 (N_11771,N_4716,N_5454);
nand U11772 (N_11772,N_5179,N_5143);
and U11773 (N_11773,N_4529,N_4140);
or U11774 (N_11774,N_5079,N_7640);
or U11775 (N_11775,N_7701,N_5739);
nor U11776 (N_11776,N_7926,N_7427);
and U11777 (N_11777,N_5876,N_7451);
nand U11778 (N_11778,N_4596,N_7798);
nand U11779 (N_11779,N_7611,N_7080);
nand U11780 (N_11780,N_4561,N_4328);
nor U11781 (N_11781,N_7286,N_5669);
and U11782 (N_11782,N_6396,N_5071);
and U11783 (N_11783,N_7455,N_7656);
or U11784 (N_11784,N_4380,N_5817);
nor U11785 (N_11785,N_7765,N_6155);
or U11786 (N_11786,N_5586,N_6335);
nor U11787 (N_11787,N_7021,N_6155);
and U11788 (N_11788,N_7387,N_6588);
and U11789 (N_11789,N_5945,N_5930);
nand U11790 (N_11790,N_7961,N_6419);
and U11791 (N_11791,N_6155,N_4700);
or U11792 (N_11792,N_5875,N_6986);
nor U11793 (N_11793,N_4649,N_6767);
nand U11794 (N_11794,N_7801,N_5303);
and U11795 (N_11795,N_7355,N_4940);
nor U11796 (N_11796,N_4653,N_7052);
and U11797 (N_11797,N_7289,N_5910);
and U11798 (N_11798,N_4674,N_5466);
nor U11799 (N_11799,N_7978,N_7961);
nor U11800 (N_11800,N_5401,N_4673);
nor U11801 (N_11801,N_4687,N_6191);
or U11802 (N_11802,N_5339,N_7472);
nand U11803 (N_11803,N_7985,N_6975);
or U11804 (N_11804,N_5349,N_7811);
or U11805 (N_11805,N_6210,N_6904);
nor U11806 (N_11806,N_5323,N_6405);
nor U11807 (N_11807,N_5451,N_5684);
nand U11808 (N_11808,N_6498,N_4693);
nand U11809 (N_11809,N_5189,N_4359);
nor U11810 (N_11810,N_5020,N_4514);
xor U11811 (N_11811,N_7116,N_4460);
and U11812 (N_11812,N_7019,N_4807);
or U11813 (N_11813,N_6990,N_7809);
xor U11814 (N_11814,N_6957,N_4809);
nor U11815 (N_11815,N_7687,N_4511);
and U11816 (N_11816,N_6452,N_7627);
and U11817 (N_11817,N_4525,N_5569);
nand U11818 (N_11818,N_6685,N_4911);
nor U11819 (N_11819,N_5063,N_4057);
or U11820 (N_11820,N_7317,N_5542);
nand U11821 (N_11821,N_5100,N_5798);
and U11822 (N_11822,N_4210,N_6275);
or U11823 (N_11823,N_4382,N_4910);
or U11824 (N_11824,N_6710,N_5734);
or U11825 (N_11825,N_5608,N_4343);
nand U11826 (N_11826,N_6815,N_7396);
or U11827 (N_11827,N_5605,N_4006);
nor U11828 (N_11828,N_5062,N_5954);
or U11829 (N_11829,N_7346,N_4222);
nand U11830 (N_11830,N_6500,N_6922);
nor U11831 (N_11831,N_4238,N_7240);
nand U11832 (N_11832,N_6536,N_7467);
or U11833 (N_11833,N_4797,N_5943);
nand U11834 (N_11834,N_6001,N_4083);
or U11835 (N_11835,N_4767,N_4354);
or U11836 (N_11836,N_7476,N_5154);
nor U11837 (N_11837,N_4613,N_6334);
nor U11838 (N_11838,N_5070,N_6532);
or U11839 (N_11839,N_5397,N_7087);
or U11840 (N_11840,N_7662,N_6210);
or U11841 (N_11841,N_6041,N_7677);
nor U11842 (N_11842,N_6823,N_7425);
nor U11843 (N_11843,N_6508,N_5958);
nand U11844 (N_11844,N_4513,N_4593);
or U11845 (N_11845,N_4038,N_6878);
nor U11846 (N_11846,N_4252,N_4748);
and U11847 (N_11847,N_7109,N_7008);
or U11848 (N_11848,N_6897,N_6330);
xnor U11849 (N_11849,N_5194,N_4861);
and U11850 (N_11850,N_7265,N_4614);
and U11851 (N_11851,N_4913,N_6686);
nand U11852 (N_11852,N_6295,N_7766);
or U11853 (N_11853,N_7898,N_5935);
or U11854 (N_11854,N_5643,N_7948);
and U11855 (N_11855,N_5828,N_4201);
nand U11856 (N_11856,N_7530,N_7206);
or U11857 (N_11857,N_5786,N_7275);
nor U11858 (N_11858,N_6139,N_4027);
or U11859 (N_11859,N_6672,N_5803);
nand U11860 (N_11860,N_4279,N_6926);
xnor U11861 (N_11861,N_5133,N_7115);
nor U11862 (N_11862,N_4550,N_7348);
nor U11863 (N_11863,N_7833,N_5602);
nor U11864 (N_11864,N_4811,N_6082);
nand U11865 (N_11865,N_4550,N_4248);
nand U11866 (N_11866,N_6613,N_4854);
nand U11867 (N_11867,N_4416,N_4953);
nor U11868 (N_11868,N_7657,N_4904);
xnor U11869 (N_11869,N_6679,N_5792);
nor U11870 (N_11870,N_5296,N_4071);
and U11871 (N_11871,N_7234,N_4227);
and U11872 (N_11872,N_7618,N_7591);
nor U11873 (N_11873,N_4031,N_6349);
and U11874 (N_11874,N_6526,N_4403);
and U11875 (N_11875,N_7088,N_6046);
nor U11876 (N_11876,N_6786,N_6778);
nor U11877 (N_11877,N_7195,N_5727);
and U11878 (N_11878,N_5200,N_4683);
nand U11879 (N_11879,N_6663,N_6362);
nand U11880 (N_11880,N_4753,N_5186);
or U11881 (N_11881,N_4691,N_5961);
or U11882 (N_11882,N_6047,N_7302);
and U11883 (N_11883,N_4802,N_6737);
nor U11884 (N_11884,N_7330,N_6917);
or U11885 (N_11885,N_6305,N_5845);
nand U11886 (N_11886,N_6435,N_5486);
and U11887 (N_11887,N_7019,N_5343);
or U11888 (N_11888,N_4794,N_7537);
and U11889 (N_11889,N_6118,N_4576);
nor U11890 (N_11890,N_7725,N_4192);
and U11891 (N_11891,N_6936,N_4622);
and U11892 (N_11892,N_5935,N_7620);
or U11893 (N_11893,N_5469,N_5500);
nor U11894 (N_11894,N_7494,N_5470);
or U11895 (N_11895,N_7752,N_7236);
nor U11896 (N_11896,N_6645,N_7225);
nand U11897 (N_11897,N_7348,N_4015);
and U11898 (N_11898,N_7475,N_4606);
or U11899 (N_11899,N_4676,N_4365);
nand U11900 (N_11900,N_4398,N_4444);
nor U11901 (N_11901,N_7291,N_7190);
nand U11902 (N_11902,N_7805,N_4305);
nand U11903 (N_11903,N_5334,N_6529);
and U11904 (N_11904,N_7257,N_4171);
nand U11905 (N_11905,N_6837,N_7382);
nand U11906 (N_11906,N_4121,N_7769);
and U11907 (N_11907,N_6715,N_7994);
nor U11908 (N_11908,N_4258,N_6203);
nand U11909 (N_11909,N_7125,N_5238);
nand U11910 (N_11910,N_4037,N_5742);
and U11911 (N_11911,N_6694,N_7846);
nand U11912 (N_11912,N_6083,N_5453);
nand U11913 (N_11913,N_5636,N_6010);
and U11914 (N_11914,N_7427,N_4541);
nand U11915 (N_11915,N_4714,N_6187);
nor U11916 (N_11916,N_6627,N_5790);
nand U11917 (N_11917,N_7873,N_6450);
or U11918 (N_11918,N_7966,N_7402);
and U11919 (N_11919,N_7306,N_5958);
and U11920 (N_11920,N_5429,N_5461);
nand U11921 (N_11921,N_6864,N_4280);
and U11922 (N_11922,N_7442,N_6406);
nor U11923 (N_11923,N_7044,N_5548);
nand U11924 (N_11924,N_7222,N_5551);
nand U11925 (N_11925,N_4601,N_4248);
nor U11926 (N_11926,N_6509,N_5459);
nor U11927 (N_11927,N_4421,N_5696);
or U11928 (N_11928,N_7004,N_6327);
or U11929 (N_11929,N_4962,N_7161);
nand U11930 (N_11930,N_7044,N_6661);
nand U11931 (N_11931,N_6642,N_5174);
nand U11932 (N_11932,N_7818,N_7832);
and U11933 (N_11933,N_5861,N_4372);
and U11934 (N_11934,N_4923,N_6753);
or U11935 (N_11935,N_4620,N_7947);
nand U11936 (N_11936,N_6485,N_5535);
nor U11937 (N_11937,N_6921,N_4755);
nand U11938 (N_11938,N_7736,N_5829);
and U11939 (N_11939,N_6714,N_7525);
nor U11940 (N_11940,N_6573,N_5200);
nor U11941 (N_11941,N_6308,N_4610);
nand U11942 (N_11942,N_6930,N_4966);
nand U11943 (N_11943,N_6928,N_6497);
and U11944 (N_11944,N_7626,N_7619);
nor U11945 (N_11945,N_6247,N_6934);
or U11946 (N_11946,N_6580,N_6648);
and U11947 (N_11947,N_5672,N_7206);
and U11948 (N_11948,N_5803,N_5590);
nand U11949 (N_11949,N_4901,N_7484);
or U11950 (N_11950,N_6534,N_6248);
or U11951 (N_11951,N_6196,N_4279);
nor U11952 (N_11952,N_5573,N_5086);
nor U11953 (N_11953,N_6993,N_5280);
or U11954 (N_11954,N_5794,N_7213);
and U11955 (N_11955,N_5263,N_5005);
nor U11956 (N_11956,N_4853,N_7233);
and U11957 (N_11957,N_7974,N_7531);
and U11958 (N_11958,N_5793,N_4832);
nand U11959 (N_11959,N_4888,N_7517);
nand U11960 (N_11960,N_4521,N_7824);
nor U11961 (N_11961,N_6862,N_5281);
or U11962 (N_11962,N_6480,N_7298);
or U11963 (N_11963,N_5186,N_6477);
or U11964 (N_11964,N_6618,N_5500);
or U11965 (N_11965,N_7797,N_4748);
nor U11966 (N_11966,N_4850,N_7283);
nand U11967 (N_11967,N_5874,N_6459);
and U11968 (N_11968,N_5270,N_7433);
xnor U11969 (N_11969,N_5342,N_5027);
nor U11970 (N_11970,N_5975,N_6691);
or U11971 (N_11971,N_7062,N_5573);
nor U11972 (N_11972,N_7712,N_7099);
nor U11973 (N_11973,N_7385,N_7613);
nor U11974 (N_11974,N_4981,N_6111);
nor U11975 (N_11975,N_4260,N_4177);
nand U11976 (N_11976,N_4203,N_7603);
nor U11977 (N_11977,N_5217,N_5673);
nand U11978 (N_11978,N_4909,N_7729);
and U11979 (N_11979,N_5581,N_6820);
and U11980 (N_11980,N_5031,N_5947);
or U11981 (N_11981,N_5110,N_4313);
nor U11982 (N_11982,N_7279,N_4421);
or U11983 (N_11983,N_6610,N_7167);
or U11984 (N_11984,N_4415,N_6502);
nand U11985 (N_11985,N_5608,N_6576);
or U11986 (N_11986,N_7359,N_7503);
and U11987 (N_11987,N_5093,N_7438);
or U11988 (N_11988,N_7393,N_7157);
nor U11989 (N_11989,N_7851,N_7350);
nand U11990 (N_11990,N_7754,N_5861);
nand U11991 (N_11991,N_4161,N_7435);
nor U11992 (N_11992,N_7203,N_7207);
nand U11993 (N_11993,N_7059,N_6498);
nor U11994 (N_11994,N_7746,N_5487);
and U11995 (N_11995,N_6136,N_6808);
nand U11996 (N_11996,N_4647,N_6905);
nor U11997 (N_11997,N_4597,N_7773);
and U11998 (N_11998,N_7916,N_5370);
or U11999 (N_11999,N_7368,N_5637);
and U12000 (N_12000,N_10385,N_8093);
or U12001 (N_12001,N_10567,N_10862);
nor U12002 (N_12002,N_11570,N_9177);
and U12003 (N_12003,N_9751,N_9091);
or U12004 (N_12004,N_10530,N_8373);
nor U12005 (N_12005,N_8656,N_11348);
nand U12006 (N_12006,N_10750,N_8718);
nor U12007 (N_12007,N_11700,N_10569);
nor U12008 (N_12008,N_10179,N_10905);
and U12009 (N_12009,N_9489,N_9030);
or U12010 (N_12010,N_8307,N_10037);
nor U12011 (N_12011,N_8902,N_9031);
or U12012 (N_12012,N_10985,N_11222);
or U12013 (N_12013,N_8658,N_9998);
and U12014 (N_12014,N_10816,N_10394);
or U12015 (N_12015,N_8281,N_11175);
nor U12016 (N_12016,N_11772,N_9036);
nand U12017 (N_12017,N_10747,N_9678);
nor U12018 (N_12018,N_8524,N_10998);
or U12019 (N_12019,N_9529,N_11828);
or U12020 (N_12020,N_11007,N_11301);
or U12021 (N_12021,N_8827,N_11477);
and U12022 (N_12022,N_8435,N_11227);
and U12023 (N_12023,N_8572,N_11894);
nand U12024 (N_12024,N_8810,N_9522);
nand U12025 (N_12025,N_9835,N_10267);
and U12026 (N_12026,N_11687,N_11487);
and U12027 (N_12027,N_10430,N_11034);
nand U12028 (N_12028,N_9558,N_8650);
nand U12029 (N_12029,N_11978,N_10201);
or U12030 (N_12030,N_8198,N_10587);
nor U12031 (N_12031,N_11986,N_10525);
nand U12032 (N_12032,N_10200,N_11784);
or U12033 (N_12033,N_8331,N_11145);
nor U12034 (N_12034,N_8360,N_10344);
nor U12035 (N_12035,N_8151,N_9782);
nand U12036 (N_12036,N_11091,N_10528);
nand U12037 (N_12037,N_11383,N_10938);
or U12038 (N_12038,N_9092,N_8762);
nand U12039 (N_12039,N_9926,N_11401);
or U12040 (N_12040,N_8688,N_8088);
nand U12041 (N_12041,N_8239,N_11272);
and U12042 (N_12042,N_11172,N_8903);
nor U12043 (N_12043,N_8941,N_11470);
nor U12044 (N_12044,N_11742,N_9222);
xnor U12045 (N_12045,N_8595,N_10029);
nor U12046 (N_12046,N_11992,N_8452);
and U12047 (N_12047,N_11727,N_11333);
nand U12048 (N_12048,N_10011,N_8060);
and U12049 (N_12049,N_9130,N_11887);
and U12050 (N_12050,N_11170,N_10239);
or U12051 (N_12051,N_8104,N_10506);
nor U12052 (N_12052,N_9714,N_10081);
nor U12053 (N_12053,N_10433,N_10763);
and U12054 (N_12054,N_10994,N_8953);
and U12055 (N_12055,N_11443,N_11220);
nor U12056 (N_12056,N_10323,N_8070);
or U12057 (N_12057,N_10142,N_10890);
or U12058 (N_12058,N_11631,N_9661);
nand U12059 (N_12059,N_10184,N_8448);
and U12060 (N_12060,N_10228,N_10602);
or U12061 (N_12061,N_8900,N_8698);
nand U12062 (N_12062,N_8474,N_9243);
and U12063 (N_12063,N_9015,N_10275);
nor U12064 (N_12064,N_11239,N_11540);
nor U12065 (N_12065,N_9963,N_10290);
nor U12066 (N_12066,N_10926,N_11962);
or U12067 (N_12067,N_11778,N_10366);
or U12068 (N_12068,N_8608,N_8115);
nor U12069 (N_12069,N_8712,N_9220);
nand U12070 (N_12070,N_10893,N_11505);
and U12071 (N_12071,N_10552,N_10393);
or U12072 (N_12072,N_8132,N_9893);
and U12073 (N_12073,N_8199,N_11511);
nor U12074 (N_12074,N_9607,N_10683);
xnor U12075 (N_12075,N_11711,N_10751);
or U12076 (N_12076,N_10818,N_8032);
nand U12077 (N_12077,N_8432,N_11226);
or U12078 (N_12078,N_8125,N_9350);
and U12079 (N_12079,N_11783,N_9076);
or U12080 (N_12080,N_8250,N_11524);
nand U12081 (N_12081,N_10513,N_10606);
nand U12082 (N_12082,N_8910,N_8426);
nor U12083 (N_12083,N_11902,N_8407);
or U12084 (N_12084,N_9160,N_11840);
nor U12085 (N_12085,N_11782,N_10349);
nand U12086 (N_12086,N_9448,N_9388);
or U12087 (N_12087,N_11110,N_8570);
xor U12088 (N_12088,N_9333,N_8927);
or U12089 (N_12089,N_9827,N_10934);
nand U12090 (N_12090,N_10671,N_8583);
and U12091 (N_12091,N_11102,N_8803);
nand U12092 (N_12092,N_9563,N_11770);
nor U12093 (N_12093,N_9271,N_11943);
xnor U12094 (N_12094,N_9635,N_8057);
nand U12095 (N_12095,N_9737,N_8215);
nand U12096 (N_12096,N_8922,N_9949);
nand U12097 (N_12097,N_8556,N_11389);
nor U12098 (N_12098,N_9007,N_9857);
and U12099 (N_12099,N_8613,N_11789);
nand U12100 (N_12100,N_11623,N_10988);
and U12101 (N_12101,N_9624,N_9037);
nand U12102 (N_12102,N_9372,N_10016);
nand U12103 (N_12103,N_8555,N_8732);
nand U12104 (N_12104,N_8495,N_10266);
nand U12105 (N_12105,N_8787,N_8591);
or U12106 (N_12106,N_9469,N_8358);
and U12107 (N_12107,N_11530,N_11653);
nor U12108 (N_12108,N_8429,N_9139);
or U12109 (N_12109,N_8870,N_10071);
and U12110 (N_12110,N_8867,N_10279);
nand U12111 (N_12111,N_10743,N_11276);
xnor U12112 (N_12112,N_11686,N_11982);
nand U12113 (N_12113,N_8794,N_11247);
nor U12114 (N_12114,N_8574,N_9593);
nor U12115 (N_12115,N_8559,N_9476);
and U12116 (N_12116,N_11406,N_9959);
nor U12117 (N_12117,N_9877,N_11039);
and U12118 (N_12118,N_11868,N_9648);
nor U12119 (N_12119,N_8341,N_8837);
nor U12120 (N_12120,N_11205,N_8222);
nand U12121 (N_12121,N_8348,N_10832);
nor U12122 (N_12122,N_9933,N_10064);
and U12123 (N_12123,N_9394,N_10965);
and U12124 (N_12124,N_9109,N_10821);
or U12125 (N_12125,N_10702,N_8587);
and U12126 (N_12126,N_9509,N_10805);
nand U12127 (N_12127,N_9019,N_11682);
nor U12128 (N_12128,N_9767,N_11891);
nand U12129 (N_12129,N_11599,N_8871);
or U12130 (N_12130,N_8036,N_9807);
nor U12131 (N_12131,N_8451,N_9916);
nor U12132 (N_12132,N_11837,N_8736);
nor U12133 (N_12133,N_11269,N_8883);
and U12134 (N_12134,N_10610,N_11280);
and U12135 (N_12135,N_11850,N_11201);
nor U12136 (N_12136,N_9851,N_9823);
and U12137 (N_12137,N_8631,N_10539);
or U12138 (N_12138,N_10744,N_9490);
or U12139 (N_12139,N_9174,N_8702);
nor U12140 (N_12140,N_8445,N_10262);
nor U12141 (N_12141,N_8720,N_8911);
nand U12142 (N_12142,N_8383,N_9942);
nor U12143 (N_12143,N_8691,N_8487);
or U12144 (N_12144,N_11278,N_11958);
or U12145 (N_12145,N_11225,N_9517);
nor U12146 (N_12146,N_9217,N_9708);
or U12147 (N_12147,N_9687,N_10629);
and U12148 (N_12148,N_11701,N_11000);
nor U12149 (N_12149,N_10535,N_9176);
nand U12150 (N_12150,N_10878,N_8097);
or U12151 (N_12151,N_11413,N_9148);
and U12152 (N_12152,N_11564,N_11569);
nand U12153 (N_12153,N_9623,N_10450);
or U12154 (N_12154,N_10304,N_9586);
and U12155 (N_12155,N_10109,N_10792);
nor U12156 (N_12156,N_8368,N_8007);
or U12157 (N_12157,N_8447,N_11402);
nor U12158 (N_12158,N_11922,N_11409);
and U12159 (N_12159,N_10462,N_10054);
or U12160 (N_12160,N_8805,N_8386);
and U12161 (N_12161,N_8991,N_11529);
nor U12162 (N_12162,N_9214,N_10800);
nand U12163 (N_12163,N_9016,N_11664);
and U12164 (N_12164,N_8783,N_10216);
nor U12165 (N_12165,N_8512,N_8262);
or U12166 (N_12166,N_10557,N_10864);
nor U12167 (N_12167,N_8039,N_11849);
and U12168 (N_12168,N_8716,N_8066);
nand U12169 (N_12169,N_9918,N_11604);
and U12170 (N_12170,N_10674,N_11748);
nand U12171 (N_12171,N_9254,N_11805);
and U12172 (N_12172,N_9227,N_10360);
nor U12173 (N_12173,N_8010,N_9716);
nand U12174 (N_12174,N_11353,N_8844);
and U12175 (N_12175,N_10568,N_10426);
or U12176 (N_12176,N_8601,N_9669);
or U12177 (N_12177,N_10693,N_11467);
nor U12178 (N_12178,N_8935,N_9314);
nor U12179 (N_12179,N_11160,N_11014);
or U12180 (N_12180,N_8567,N_10100);
nand U12181 (N_12181,N_11036,N_9673);
nor U12182 (N_12182,N_11498,N_9233);
or U12183 (N_12183,N_8117,N_9183);
and U12184 (N_12184,N_10570,N_10692);
or U12185 (N_12185,N_9798,N_10456);
nor U12186 (N_12186,N_8390,N_8237);
nand U12187 (N_12187,N_10155,N_9609);
xnor U12188 (N_12188,N_9154,N_8232);
and U12189 (N_12189,N_10466,N_9017);
and U12190 (N_12190,N_10065,N_8836);
nand U12191 (N_12191,N_8674,N_9001);
and U12192 (N_12192,N_10645,N_9791);
or U12193 (N_12193,N_10622,N_8054);
xnor U12194 (N_12194,N_8897,N_11606);
nand U12195 (N_12195,N_9184,N_10617);
or U12196 (N_12196,N_8596,N_11520);
nor U12197 (N_12197,N_8138,N_10901);
nand U12198 (N_12198,N_8327,N_8534);
and U12199 (N_12199,N_10654,N_8682);
nor U12200 (N_12200,N_8073,N_8764);
xor U12201 (N_12201,N_10390,N_9417);
or U12202 (N_12202,N_11066,N_9523);
nor U12203 (N_12203,N_8485,N_8486);
or U12204 (N_12204,N_8318,N_9844);
nor U12205 (N_12205,N_9068,N_10869);
nor U12206 (N_12206,N_10440,N_10149);
or U12207 (N_12207,N_9799,N_10108);
and U12208 (N_12208,N_8284,N_9083);
nor U12209 (N_12209,N_8645,N_11508);
and U12210 (N_12210,N_10399,N_10590);
nand U12211 (N_12211,N_11720,N_8663);
nand U12212 (N_12212,N_10746,N_11869);
and U12213 (N_12213,N_8380,N_10565);
nor U12214 (N_12214,N_9119,N_11185);
and U12215 (N_12215,N_9287,N_11150);
and U12216 (N_12216,N_8995,N_11703);
and U12217 (N_12217,N_9003,N_10580);
or U12218 (N_12218,N_9599,N_9867);
and U12219 (N_12219,N_9058,N_8742);
nand U12220 (N_12220,N_10190,N_11440);
and U12221 (N_12221,N_8760,N_8547);
and U12222 (N_12222,N_10953,N_10555);
or U12223 (N_12223,N_10949,N_11515);
nand U12224 (N_12224,N_9571,N_9142);
nand U12225 (N_12225,N_11399,N_8956);
nor U12226 (N_12226,N_9014,N_10457);
nor U12227 (N_12227,N_10300,N_9616);
nand U12228 (N_12228,N_10742,N_11715);
or U12229 (N_12229,N_10461,N_9568);
and U12230 (N_12230,N_10055,N_11182);
or U12231 (N_12231,N_11268,N_9895);
nor U12232 (N_12232,N_10043,N_11643);
nand U12233 (N_12233,N_11331,N_10002);
nand U12234 (N_12234,N_8826,N_11549);
nand U12235 (N_12235,N_8108,N_9230);
and U12236 (N_12236,N_10915,N_11108);
or U12237 (N_12237,N_11147,N_11735);
nor U12238 (N_12238,N_8116,N_9114);
nor U12239 (N_12239,N_8276,N_11547);
and U12240 (N_12240,N_9574,N_11306);
nor U12241 (N_12241,N_11527,N_10761);
and U12242 (N_12242,N_9501,N_11836);
or U12243 (N_12243,N_8785,N_11075);
or U12244 (N_12244,N_8179,N_9371);
or U12245 (N_12245,N_10181,N_11574);
nand U12246 (N_12246,N_8012,N_11058);
nor U12247 (N_12247,N_8210,N_10336);
or U12248 (N_12248,N_11873,N_9817);
or U12249 (N_12249,N_10755,N_8471);
and U12250 (N_12250,N_9284,N_11284);
nor U12251 (N_12251,N_10607,N_10357);
or U12252 (N_12252,N_11590,N_10971);
nor U12253 (N_12253,N_11372,N_10014);
nand U12254 (N_12254,N_10130,N_8385);
and U12255 (N_12255,N_10589,N_9738);
or U12256 (N_12256,N_8816,N_9059);
nand U12257 (N_12257,N_11612,N_9659);
nor U12258 (N_12258,N_10233,N_9706);
and U12259 (N_12259,N_9885,N_8080);
nand U12260 (N_12260,N_11636,N_8023);
or U12261 (N_12261,N_11461,N_10022);
nand U12262 (N_12262,N_10386,N_9210);
nand U12263 (N_12263,N_8016,N_9644);
nor U12264 (N_12264,N_8183,N_9471);
and U12265 (N_12265,N_8172,N_10854);
and U12266 (N_12266,N_8299,N_10019);
nand U12267 (N_12267,N_10479,N_10989);
and U12268 (N_12268,N_8295,N_10235);
nand U12269 (N_12269,N_11924,N_8413);
and U12270 (N_12270,N_10137,N_9821);
and U12271 (N_12271,N_8599,N_9125);
nor U12272 (N_12272,N_9202,N_11038);
nand U12273 (N_12273,N_8424,N_11342);
nand U12274 (N_12274,N_9793,N_9968);
and U12275 (N_12275,N_8632,N_8503);
or U12276 (N_12276,N_9620,N_9355);
nand U12277 (N_12277,N_8800,N_10085);
nand U12278 (N_12278,N_11688,N_10937);
and U12279 (N_12279,N_9131,N_8157);
xor U12280 (N_12280,N_8293,N_10904);
or U12281 (N_12281,N_8192,N_11138);
xor U12282 (N_12282,N_9377,N_9225);
xor U12283 (N_12283,N_10132,N_8978);
nand U12284 (N_12284,N_9118,N_9790);
and U12285 (N_12285,N_10895,N_9294);
and U12286 (N_12286,N_11362,N_10280);
and U12287 (N_12287,N_9047,N_9600);
nor U12288 (N_12288,N_9163,N_11886);
or U12289 (N_12289,N_11369,N_11394);
nor U12290 (N_12290,N_10882,N_9773);
and U12291 (N_12291,N_10863,N_9424);
nand U12292 (N_12292,N_9858,N_11290);
and U12293 (N_12293,N_9820,N_10253);
nor U12294 (N_12294,N_11806,N_8392);
nand U12295 (N_12295,N_8517,N_11626);
nand U12296 (N_12296,N_10401,N_11573);
nor U12297 (N_12297,N_10355,N_9997);
or U12298 (N_12298,N_11340,N_9402);
or U12299 (N_12299,N_11258,N_11006);
or U12300 (N_12300,N_11499,N_10082);
and U12301 (N_12301,N_10489,N_8319);
nor U12302 (N_12302,N_10773,N_11457);
or U12303 (N_12303,N_10665,N_11318);
nor U12304 (N_12304,N_11001,N_11624);
nor U12305 (N_12305,N_11017,N_8029);
nand U12306 (N_12306,N_10306,N_11486);
or U12307 (N_12307,N_8045,N_10911);
nand U12308 (N_12308,N_10198,N_8796);
or U12309 (N_12309,N_10448,N_9438);
or U12310 (N_12310,N_10775,N_11531);
or U12311 (N_12311,N_8003,N_9265);
or U12312 (N_12312,N_8363,N_11536);
or U12313 (N_12313,N_10490,N_11684);
or U12314 (N_12314,N_11602,N_8751);
and U12315 (N_12315,N_10368,N_10110);
and U12316 (N_12316,N_9179,N_9164);
or U12317 (N_12317,N_8706,N_9038);
and U12318 (N_12318,N_11708,N_10260);
nor U12319 (N_12319,N_10000,N_9513);
nand U12320 (N_12320,N_9994,N_11293);
nor U12321 (N_12321,N_10648,N_11810);
or U12322 (N_12322,N_10739,N_9248);
or U12323 (N_12323,N_11853,N_11552);
or U12324 (N_12324,N_10546,N_10397);
and U12325 (N_12325,N_8538,N_9946);
and U12326 (N_12326,N_8858,N_9507);
and U12327 (N_12327,N_8161,N_8456);
nor U12328 (N_12328,N_8376,N_10205);
and U12329 (N_12329,N_9508,N_10678);
or U12330 (N_12330,N_10951,N_9537);
or U12331 (N_12331,N_9457,N_8843);
nand U12332 (N_12332,N_10619,N_10125);
and U12333 (N_12333,N_11725,N_11244);
or U12334 (N_12334,N_9805,N_8711);
nor U12335 (N_12335,N_11618,N_9084);
nor U12336 (N_12336,N_9715,N_11099);
nand U12337 (N_12337,N_8223,N_10302);
nor U12338 (N_12338,N_11469,N_11378);
nand U12339 (N_12339,N_9707,N_9080);
or U12340 (N_12340,N_11667,N_9010);
and U12341 (N_12341,N_11941,N_11193);
nand U12342 (N_12342,N_9944,N_8668);
nand U12343 (N_12343,N_10710,N_8067);
nand U12344 (N_12344,N_9645,N_8387);
and U12345 (N_12345,N_8347,N_9069);
or U12346 (N_12346,N_11442,N_9231);
and U12347 (N_12347,N_11171,N_9679);
or U12348 (N_12348,N_11230,N_11827);
nand U12349 (N_12349,N_10049,N_10340);
and U12350 (N_12350,N_9432,N_11198);
nand U12351 (N_12351,N_10767,N_8278);
nor U12352 (N_12352,N_10494,N_11031);
xor U12353 (N_12353,N_8554,N_11944);
and U12354 (N_12354,N_9911,N_10026);
and U12355 (N_12355,N_8196,N_8100);
or U12356 (N_12356,N_8047,N_11365);
nand U12357 (N_12357,N_10406,N_9257);
nor U12358 (N_12358,N_9194,N_10036);
nand U12359 (N_12359,N_10066,N_11003);
nand U12360 (N_12360,N_11468,N_10636);
nand U12361 (N_12361,N_8197,N_11330);
and U12362 (N_12362,N_8932,N_8735);
and U12363 (N_12363,N_10059,N_8779);
nor U12364 (N_12364,N_9397,N_9411);
or U12365 (N_12365,N_11656,N_9928);
nor U12366 (N_12366,N_11263,N_10993);
and U12367 (N_12367,N_8807,N_11070);
nor U12368 (N_12368,N_10122,N_11156);
or U12369 (N_12369,N_11181,N_10416);
and U12370 (N_12370,N_10141,N_10412);
nor U12371 (N_12371,N_9796,N_10229);
nand U12372 (N_12372,N_11803,N_8838);
or U12373 (N_12373,N_10786,N_11747);
or U12374 (N_12374,N_10135,N_11859);
or U12375 (N_12375,N_11396,N_11051);
or U12376 (N_12376,N_8131,N_8946);
or U12377 (N_12377,N_9369,N_11423);
or U12378 (N_12378,N_8315,N_11454);
and U12379 (N_12379,N_9259,N_9903);
and U12380 (N_12380,N_9153,N_10270);
or U12381 (N_12381,N_9956,N_8337);
nor U12382 (N_12382,N_10512,N_8549);
or U12383 (N_12383,N_11358,N_8257);
nor U12384 (N_12384,N_10236,N_10756);
nor U12385 (N_12385,N_11266,N_8737);
nand U12386 (N_12386,N_10738,N_8825);
and U12387 (N_12387,N_10644,N_10417);
and U12388 (N_12388,N_10312,N_9633);
and U12389 (N_12389,N_10987,N_11609);
and U12390 (N_12390,N_9876,N_10460);
nand U12391 (N_12391,N_9358,N_8063);
nand U12392 (N_12392,N_9731,N_11286);
and U12393 (N_12393,N_11165,N_8026);
and U12394 (N_12394,N_11525,N_9362);
xor U12395 (N_12395,N_10234,N_8030);
or U12396 (N_12396,N_11951,N_11503);
nor U12397 (N_12397,N_9423,N_10363);
and U12398 (N_12398,N_11839,N_9165);
and U12399 (N_12399,N_11802,N_9374);
or U12400 (N_12400,N_8884,N_9026);
or U12401 (N_12401,N_8312,N_8440);
and U12402 (N_12402,N_10757,N_11645);
nor U12403 (N_12403,N_9258,N_8968);
or U12404 (N_12404,N_10396,N_8344);
and U12405 (N_12405,N_10913,N_9831);
nand U12406 (N_12406,N_11509,N_8297);
nand U12407 (N_12407,N_10405,N_10701);
nor U12408 (N_12408,N_8111,N_10923);
nand U12409 (N_12409,N_8494,N_11862);
nor U12410 (N_12410,N_8561,N_11680);
or U12411 (N_12411,N_9481,N_10389);
nor U12412 (N_12412,N_9988,N_11831);
and U12413 (N_12413,N_8925,N_8694);
or U12414 (N_12414,N_9376,N_8072);
nand U12415 (N_12415,N_9102,N_10928);
nand U12416 (N_12416,N_9575,N_10099);
nand U12417 (N_12417,N_11973,N_8689);
nand U12418 (N_12418,N_10810,N_11288);
and U12419 (N_12419,N_10851,N_10917);
and U12420 (N_12420,N_10483,N_8042);
nand U12421 (N_12421,N_11398,N_10296);
or U12422 (N_12422,N_10735,N_10966);
or U12423 (N_12423,N_11062,N_8869);
nor U12424 (N_12424,N_11814,N_10365);
nor U12425 (N_12425,N_11760,N_8382);
nor U12426 (N_12426,N_10331,N_11240);
nor U12427 (N_12427,N_9193,N_10127);
or U12428 (N_12428,N_9646,N_11421);
or U12429 (N_12429,N_10929,N_8573);
nand U12430 (N_12430,N_10319,N_10486);
nand U12431 (N_12431,N_9234,N_10660);
nand U12432 (N_12432,N_10898,N_11065);
or U12433 (N_12433,N_10025,N_11692);
and U12434 (N_12434,N_11625,N_10620);
or U12435 (N_12435,N_9240,N_8264);
and U12436 (N_12436,N_9764,N_9781);
nor U12437 (N_12437,N_9601,N_11542);
and U12438 (N_12438,N_8401,N_9078);
or U12439 (N_12439,N_9541,N_8926);
or U12440 (N_12440,N_8562,N_9875);
or U12441 (N_12441,N_9450,N_10615);
nor U12442 (N_12442,N_10721,N_10910);
or U12443 (N_12443,N_9710,N_10837);
nand U12444 (N_12444,N_9533,N_11950);
or U12445 (N_12445,N_8168,N_10601);
and U12446 (N_12446,N_10498,N_10139);
or U12447 (N_12447,N_11094,N_8819);
nor U12448 (N_12448,N_11723,N_8181);
nor U12449 (N_12449,N_11119,N_10400);
or U12450 (N_12450,N_11431,N_11676);
xnor U12451 (N_12451,N_8552,N_11654);
xnor U12452 (N_12452,N_10885,N_9011);
and U12453 (N_12453,N_11011,N_11513);
xor U12454 (N_12454,N_11610,N_9236);
or U12455 (N_12455,N_8644,N_10307);
or U12456 (N_12456,N_9880,N_8078);
nand U12457 (N_12457,N_9307,N_10154);
or U12458 (N_12458,N_11100,N_9639);
nor U12459 (N_12459,N_8541,N_10045);
and U12460 (N_12460,N_8896,N_9052);
and U12461 (N_12461,N_10481,N_10611);
nand U12462 (N_12462,N_8763,N_9954);
and U12463 (N_12463,N_10586,N_10733);
or U12464 (N_12464,N_9467,N_11722);
nand U12465 (N_12465,N_10484,N_10421);
nand U12466 (N_12466,N_10255,N_8335);
and U12467 (N_12467,N_9292,N_8890);
and U12468 (N_12468,N_10825,N_8614);
nand U12469 (N_12469,N_10585,N_9381);
nand U12470 (N_12470,N_9288,N_11086);
nor U12471 (N_12471,N_8498,N_11303);
nand U12472 (N_12472,N_11002,N_8277);
nor U12473 (N_12473,N_9213,N_8643);
nand U12474 (N_12474,N_9426,N_9811);
nand U12475 (N_12475,N_11166,N_8155);
and U12476 (N_12476,N_8346,N_9693);
or U12477 (N_12477,N_8921,N_11641);
or U12478 (N_12478,N_11644,N_8960);
nor U12479 (N_12479,N_8038,N_11865);
and U12480 (N_12480,N_9856,N_8345);
nor U12481 (N_12481,N_11129,N_10380);
nor U12482 (N_12482,N_9524,N_9306);
or U12483 (N_12483,N_10437,N_8412);
nor U12484 (N_12484,N_8544,N_9634);
or U12485 (N_12485,N_8449,N_9800);
or U12486 (N_12486,N_10439,N_9311);
or U12487 (N_12487,N_11219,N_9697);
and U12488 (N_12488,N_8727,N_9349);
or U12489 (N_12489,N_10553,N_9705);
or U12490 (N_12490,N_10291,N_10298);
nor U12491 (N_12491,N_9181,N_8714);
and U12492 (N_12492,N_8962,N_9526);
and U12493 (N_12493,N_8798,N_11285);
nand U12494 (N_12494,N_11673,N_11140);
and U12495 (N_12495,N_10826,N_9939);
or U12496 (N_12496,N_11955,N_9486);
or U12497 (N_12497,N_10058,N_11134);
nor U12498 (N_12498,N_9770,N_11658);
nor U12499 (N_12499,N_9447,N_8062);
nor U12500 (N_12500,N_11382,N_9115);
and U12501 (N_12501,N_8976,N_11364);
nor U12502 (N_12502,N_11890,N_9106);
or U12503 (N_12503,N_8229,N_8831);
nor U12504 (N_12504,N_11047,N_8349);
or U12505 (N_12505,N_11972,N_9352);
or U12506 (N_12506,N_11112,N_8142);
or U12507 (N_12507,N_11638,N_10752);
nand U12508 (N_12508,N_11907,N_9548);
or U12509 (N_12509,N_8961,N_9694);
or U12510 (N_12510,N_8004,N_8667);
or U12511 (N_12511,N_10372,N_9463);
and U12512 (N_12512,N_9188,N_11718);
and U12513 (N_12513,N_9290,N_9162);
nor U12514 (N_12514,N_11123,N_11153);
nand U12515 (N_12515,N_10517,N_8126);
or U12516 (N_12516,N_9690,N_10543);
or U12517 (N_12517,N_10537,N_10423);
and U12518 (N_12518,N_11111,N_8227);
nor U12519 (N_12519,N_10131,N_9000);
and U12520 (N_12520,N_8865,N_9096);
and U12521 (N_12521,N_9536,N_11337);
and U12522 (N_12522,N_10801,N_9110);
or U12523 (N_12523,N_8610,N_10865);
and U12524 (N_12524,N_8411,N_8289);
or U12525 (N_12525,N_11127,N_11143);
nor U12526 (N_12526,N_8765,N_9925);
and U12527 (N_12527,N_10695,N_9497);
and U12528 (N_12528,N_10112,N_8450);
and U12529 (N_12529,N_8988,N_11852);
nor U12530 (N_12530,N_9120,N_8367);
or U12531 (N_12531,N_9229,N_9562);
xor U12532 (N_12532,N_10215,N_10010);
and U12533 (N_12533,N_10754,N_11072);
and U12534 (N_12534,N_8272,N_9395);
nand U12535 (N_12535,N_10070,N_8464);
nor U12536 (N_12536,N_8258,N_11203);
and U12537 (N_12537,N_11872,N_9878);
nor U12538 (N_12538,N_11121,N_11825);
or U12539 (N_12539,N_9121,N_9027);
xor U12540 (N_12540,N_9853,N_10133);
nor U12541 (N_12541,N_10244,N_11555);
xnor U12542 (N_12542,N_8928,N_10724);
nand U12543 (N_12543,N_10327,N_10653);
nor U12544 (N_12544,N_9849,N_9180);
or U12545 (N_12545,N_10097,N_8120);
nor U12546 (N_12546,N_9342,N_8421);
or U12547 (N_12547,N_10514,N_8577);
and U12548 (N_12548,N_9219,N_10325);
or U12549 (N_12549,N_10158,N_11546);
nand U12550 (N_12550,N_9466,N_8539);
nor U12551 (N_12551,N_10700,N_10548);
and U12552 (N_12552,N_10123,N_10712);
nor U12553 (N_12553,N_11940,N_11412);
nand U12554 (N_12554,N_9122,N_10519);
and U12555 (N_12555,N_8937,N_9825);
nand U12556 (N_12556,N_11375,N_10762);
or U12557 (N_12557,N_11107,N_11287);
nor U12558 (N_12558,N_9309,N_11238);
nand U12559 (N_12559,N_11035,N_9657);
nand U12560 (N_12560,N_8766,N_9757);
nor U12561 (N_12561,N_10633,N_9367);
nor U12562 (N_12562,N_11595,N_10624);
or U12563 (N_12563,N_11518,N_9830);
or U12564 (N_12564,N_8158,N_8954);
or U12565 (N_12565,N_9896,N_9062);
nor U12566 (N_12566,N_11124,N_9488);
and U12567 (N_12567,N_10688,N_8334);
nand U12568 (N_12568,N_9129,N_9128);
or U12569 (N_12569,N_9921,N_9649);
nand U12570 (N_12570,N_10402,N_8499);
nand U12571 (N_12571,N_9753,N_10523);
nand U12572 (N_12572,N_8887,N_10277);
or U12573 (N_12573,N_10899,N_11428);
and U12574 (N_12574,N_8781,N_8374);
and U12575 (N_12575,N_9865,N_11122);
or U12576 (N_12576,N_9503,N_8009);
or U12577 (N_12577,N_11550,N_9505);
and U12578 (N_12578,N_10497,N_11324);
or U12579 (N_12579,N_9116,N_10441);
or U12580 (N_12580,N_10652,N_11261);
nor U12581 (N_12581,N_10425,N_9774);
nand U12582 (N_12582,N_11101,N_8880);
or U12583 (N_12583,N_9277,N_10278);
and U12584 (N_12584,N_11693,N_11496);
xnor U12585 (N_12585,N_9957,N_11282);
nand U12586 (N_12586,N_8860,N_8321);
nand U12587 (N_12587,N_9146,N_8994);
nor U12588 (N_12588,N_8273,N_9126);
nand U12589 (N_12589,N_11300,N_9766);
or U12590 (N_12590,N_8502,N_8841);
nand U12591 (N_12591,N_11728,N_9018);
and U12592 (N_12592,N_8015,N_10467);
nand U12593 (N_12593,N_8579,N_10959);
nand U12594 (N_12594,N_9462,N_8920);
or U12595 (N_12595,N_10667,N_10948);
xor U12596 (N_12596,N_11584,N_8989);
nand U12597 (N_12597,N_9917,N_10942);
nor U12598 (N_12598,N_10670,N_11652);
nor U12599 (N_12599,N_10076,N_10114);
or U12600 (N_12600,N_10732,N_11874);
nor U12601 (N_12601,N_8877,N_11816);
nor U12602 (N_12602,N_11927,N_9855);
and U12603 (N_12603,N_11298,N_11560);
nand U12604 (N_12604,N_8221,N_9384);
nor U12605 (N_12605,N_9683,N_11947);
or U12606 (N_12606,N_9260,N_10173);
and U12607 (N_12607,N_9555,N_9067);
or U12608 (N_12608,N_9682,N_11329);
nor U12609 (N_12609,N_9317,N_10876);
nor U12610 (N_12610,N_9984,N_8384);
or U12611 (N_12611,N_9403,N_9869);
or U12612 (N_12612,N_11196,N_11906);
nor U12613 (N_12613,N_9598,N_11705);
xor U12614 (N_12614,N_9012,N_9323);
and U12615 (N_12615,N_10939,N_8513);
or U12616 (N_12616,N_8279,N_8467);
and U12617 (N_12617,N_10242,N_11593);
nor U12618 (N_12618,N_10473,N_11968);
nor U12619 (N_12619,N_8906,N_10007);
nand U12620 (N_12620,N_9709,N_9747);
nand U12621 (N_12621,N_10374,N_10772);
or U12622 (N_12622,N_10258,N_8990);
nand U12623 (N_12623,N_11154,N_9502);
nand U12624 (N_12624,N_10807,N_9285);
nor U12625 (N_12625,N_10074,N_10935);
and U12626 (N_12626,N_11420,N_9797);
or U12627 (N_12627,N_11339,N_8930);
nand U12628 (N_12628,N_8664,N_11452);
nand U12629 (N_12629,N_8235,N_10219);
and U12630 (N_12630,N_11714,N_9546);
or U12631 (N_12631,N_8965,N_11126);
or U12632 (N_12632,N_10838,N_11146);
or U12633 (N_12633,N_8854,N_10995);
or U12634 (N_12634,N_8848,N_9980);
nor U12635 (N_12635,N_10315,N_9777);
nand U12636 (N_12636,N_8832,N_11297);
nor U12637 (N_12637,N_10614,N_10824);
nor U12638 (N_12638,N_9135,N_8634);
nor U12639 (N_12639,N_8697,N_11834);
and U12640 (N_12640,N_8641,N_9638);
nand U12641 (N_12641,N_11743,N_11233);
nor U12642 (N_12642,N_9578,N_11472);
nand U12643 (N_12643,N_11884,N_9653);
nand U12644 (N_12644,N_8690,N_10111);
nor U12645 (N_12645,N_9676,N_11662);
nand U12646 (N_12646,N_10193,N_8955);
and U12647 (N_12647,N_10286,N_10276);
and U12648 (N_12648,N_10272,N_8923);
or U12649 (N_12649,N_8035,N_9573);
and U12650 (N_12650,N_11242,N_11309);
or U12651 (N_12651,N_11013,N_9866);
nand U12652 (N_12652,N_10886,N_10984);
nand U12653 (N_12653,N_10577,N_8455);
or U12654 (N_12654,N_9385,N_10954);
nor U12655 (N_12655,N_10811,N_9688);
nor U12656 (N_12656,N_9979,N_9618);
nor U12657 (N_12657,N_11691,N_9982);
nand U12658 (N_12658,N_8233,N_8895);
and U12659 (N_12659,N_9204,N_10453);
and U12660 (N_12660,N_9868,N_11404);
nand U12661 (N_12661,N_8489,N_9413);
or U12662 (N_12662,N_11104,N_9216);
or U12663 (N_12663,N_9945,N_10978);
or U12664 (N_12664,N_10347,N_8777);
and U12665 (N_12665,N_10495,N_11841);
nand U12666 (N_12666,N_11679,N_10875);
nand U12667 (N_12667,N_10737,N_11585);
nand U12668 (N_12668,N_10465,N_9544);
nor U12669 (N_12669,N_11912,N_10769);
and U12670 (N_12670,N_10310,N_11575);
nor U12671 (N_12671,N_9742,N_11535);
xor U12672 (N_12672,N_10573,N_11554);
nand U12673 (N_12673,N_9098,N_9404);
xor U12674 (N_12674,N_10608,N_9822);
nor U12675 (N_12675,N_11795,N_11114);
and U12676 (N_12676,N_8379,N_8758);
or U12677 (N_12677,N_9654,N_8338);
nand U12678 (N_12678,N_8528,N_11501);
or U12679 (N_12679,N_8693,N_8913);
nand U12680 (N_12680,N_11311,N_10314);
or U12681 (N_12681,N_8420,N_9594);
nor U12682 (N_12682,N_9398,N_11236);
or U12683 (N_12683,N_10716,N_9379);
nand U12684 (N_12684,N_11050,N_8022);
nand U12685 (N_12685,N_10521,N_9723);
or U12686 (N_12686,N_11338,N_8463);
or U12687 (N_12687,N_8749,N_9932);
nor U12688 (N_12688,N_11844,N_8862);
nand U12689 (N_12689,N_9244,N_10933);
nand U12690 (N_12690,N_10030,N_9434);
and U12691 (N_12691,N_8571,N_11731);
and U12692 (N_12692,N_8231,N_9802);
or U12693 (N_12693,N_8745,N_10658);
nand U12694 (N_12694,N_10880,N_8280);
and U12695 (N_12695,N_11494,N_9433);
nand U12696 (N_12696,N_9409,N_8027);
or U12697 (N_12697,N_9675,N_10650);
nand U12698 (N_12698,N_10153,N_9953);
nand U12699 (N_12699,N_9343,N_11589);
nor U12700 (N_12700,N_8908,N_11040);
and U12701 (N_12701,N_8952,N_9086);
or U12702 (N_12702,N_10474,N_9322);
and U12703 (N_12703,N_9066,N_9378);
nor U12704 (N_12704,N_8761,N_11565);
nor U12705 (N_12705,N_9630,N_8692);
nor U12706 (N_12706,N_8446,N_9029);
and U12707 (N_12707,N_9478,N_11786);
or U12708 (N_12708,N_8557,N_9771);
and U12709 (N_12709,N_9701,N_8680);
nand U12710 (N_12710,N_8861,N_8167);
nand U12711 (N_12711,N_9293,N_10999);
nand U12712 (N_12712,N_8529,N_9167);
and U12713 (N_12713,N_9406,N_9725);
nor U12714 (N_12714,N_8687,N_9389);
or U12715 (N_12715,N_10501,N_10717);
nor U12716 (N_12716,N_11489,N_11934);
or U12717 (N_12717,N_9960,N_11074);
and U12718 (N_12718,N_9241,N_10859);
nor U12719 (N_12719,N_9787,N_11553);
nand U12720 (N_12720,N_11732,N_11824);
or U12721 (N_12721,N_8416,N_11241);
and U12722 (N_12722,N_10874,N_10974);
or U12723 (N_12723,N_10765,N_11041);
or U12724 (N_12724,N_8532,N_10210);
or U12725 (N_12725,N_11079,N_10496);
nand U12726 (N_12726,N_9819,N_10245);
and U12727 (N_12727,N_11870,N_10264);
or U12728 (N_12728,N_11754,N_10211);
and U12729 (N_12729,N_11188,N_11519);
nor U12730 (N_12730,N_10057,N_10593);
nand U12731 (N_12731,N_11334,N_9662);
and U12732 (N_12732,N_10361,N_8788);
nand U12733 (N_12733,N_11885,N_9941);
nor U12734 (N_12734,N_9872,N_10072);
and U12735 (N_12735,N_11777,N_8717);
nand U12736 (N_12736,N_10618,N_11510);
nor U12737 (N_12737,N_8943,N_10844);
and U12738 (N_12738,N_10980,N_9514);
xor U12739 (N_12739,N_10338,N_11347);
nor U12740 (N_12740,N_9940,N_11082);
or U12741 (N_12741,N_11925,N_11370);
and U12742 (N_12742,N_10680,N_9581);
or U12743 (N_12743,N_9606,N_10088);
nand U12744 (N_12744,N_11228,N_10388);
nor U12745 (N_12745,N_9310,N_11999);
nand U12746 (N_12746,N_11580,N_11097);
or U12747 (N_12747,N_11639,N_11085);
or U12748 (N_12748,N_9993,N_9304);
nor U12749 (N_12749,N_8958,N_8713);
nor U12750 (N_12750,N_8069,N_8313);
nor U12751 (N_12751,N_10558,N_9582);
or U12752 (N_12752,N_8907,N_11733);
or U12753 (N_12753,N_10579,N_10828);
or U12754 (N_12754,N_8225,N_10656);
xor U12755 (N_12755,N_11876,N_10785);
nand U12756 (N_12756,N_9484,N_9923);
and U12757 (N_12757,N_10729,N_8362);
or U12758 (N_12758,N_10500,N_10809);
nand U12759 (N_12759,N_9414,N_8568);
nand U12760 (N_12760,N_9642,N_10220);
nand U12761 (N_12761,N_10842,N_8018);
or U12762 (N_12762,N_10759,N_9622);
nor U12763 (N_12763,N_10776,N_11466);
nor U12764 (N_12764,N_11744,N_11586);
or U12765 (N_12765,N_8951,N_10098);
nand U12766 (N_12766,N_11043,N_8287);
nor U12767 (N_12767,N_11771,N_9881);
nor U12768 (N_12768,N_8008,N_11908);
or U12769 (N_12769,N_9585,N_10176);
nand U12770 (N_12770,N_10551,N_9667);
nand U12771 (N_12771,N_9415,N_11577);
xnor U12772 (N_12772,N_11952,N_8784);
nand U12773 (N_12773,N_10962,N_10664);
nor U12774 (N_12774,N_8970,N_9760);
nand U12775 (N_12775,N_8443,N_8590);
nand U12776 (N_12776,N_11168,N_9351);
and U12777 (N_12777,N_10326,N_9572);
nor U12778 (N_12778,N_10884,N_11155);
and U12779 (N_12779,N_9494,N_8616);
nand U12780 (N_12780,N_8772,N_8578);
nand U12781 (N_12781,N_9272,N_11710);
nand U12782 (N_12782,N_10163,N_9421);
and U12783 (N_12783,N_9208,N_11817);
nand U12784 (N_12784,N_8705,N_9981);
nor U12785 (N_12785,N_10877,N_11507);
nand U12786 (N_12786,N_9221,N_10078);
and U12787 (N_12787,N_11133,N_8089);
and U12788 (N_12788,N_9340,N_9143);
and U12789 (N_12789,N_11901,N_10147);
xnor U12790 (N_12790,N_9383,N_8771);
nand U12791 (N_12791,N_10909,N_8516);
nand U12792 (N_12792,N_9740,N_8031);
nor U12793 (N_12793,N_10562,N_10313);
nor U12794 (N_12794,N_8226,N_10860);
and U12795 (N_12795,N_11766,N_10963);
or U12796 (N_12796,N_11120,N_8056);
or U12797 (N_12797,N_11210,N_10080);
xor U12798 (N_12798,N_11914,N_8423);
and U12799 (N_12799,N_11379,N_8260);
xor U12800 (N_12800,N_8249,N_11152);
xor U12801 (N_12801,N_10912,N_8101);
or U12802 (N_12802,N_9113,N_8569);
nand U12803 (N_12803,N_8789,N_8092);
and U12804 (N_12804,N_11456,N_9475);
xor U12805 (N_12805,N_11713,N_10061);
or U12806 (N_12806,N_8845,N_9854);
nor U12807 (N_12807,N_10592,N_11438);
or U12808 (N_12808,N_11229,N_11308);
nor U12809 (N_12809,N_11916,N_10480);
or U12810 (N_12810,N_8355,N_11186);
nor U12811 (N_12811,N_9952,N_11532);
and U12812 (N_12812,N_9053,N_10572);
and U12813 (N_12813,N_9717,N_11073);
or U12814 (N_12814,N_9977,N_8410);
nand U12815 (N_12815,N_10445,N_11796);
and U12816 (N_12816,N_11232,N_11250);
nand U12817 (N_12817,N_9882,N_9792);
or U12818 (N_12818,N_11502,N_10311);
or U12819 (N_12819,N_10134,N_11480);
and U12820 (N_12820,N_11991,N_9632);
nand U12821 (N_12821,N_9028,N_8786);
or U12822 (N_12822,N_11668,N_10715);
nor U12823 (N_12823,N_10187,N_8185);
nand U12824 (N_12824,N_11963,N_8719);
and U12825 (N_12825,N_10841,N_10943);
nand U12826 (N_12826,N_8320,N_11455);
and U12827 (N_12827,N_11202,N_9579);
nand U12828 (N_12828,N_9611,N_11367);
nand U12829 (N_12829,N_9992,N_9660);
nor U12830 (N_12830,N_8780,N_8381);
and U12831 (N_12831,N_9628,N_9138);
and U12832 (N_12832,N_10042,N_8164);
nand U12833 (N_12833,N_8208,N_8102);
and U12834 (N_12834,N_8488,N_8465);
and U12835 (N_12835,N_11895,N_11611);
xnor U12836 (N_12836,N_11335,N_11323);
nor U12837 (N_12837,N_9775,N_11709);
nor U12838 (N_12838,N_10335,N_10672);
xor U12839 (N_12839,N_8851,N_10766);
or U12840 (N_12840,N_11648,N_8241);
and U12841 (N_12841,N_11197,N_11964);
xnor U12842 (N_12842,N_8715,N_11304);
nand U12843 (N_12843,N_9564,N_8734);
or U12844 (N_12844,N_10282,N_11909);
and U12845 (N_12845,N_11649,N_10538);
and U12846 (N_12846,N_8404,N_9024);
or U12847 (N_12847,N_8635,N_9927);
or U12848 (N_12848,N_10293,N_8201);
nand U12849 (N_12849,N_8149,N_9108);
xor U12850 (N_12850,N_9089,N_9665);
or U12851 (N_12851,N_8773,N_11260);
xnor U12852 (N_12852,N_9891,N_11561);
or U12853 (N_12853,N_9399,N_9088);
or U12854 (N_12854,N_10796,N_9810);
and U12855 (N_12855,N_8997,N_10846);
nand U12856 (N_12856,N_11523,N_8814);
and U12857 (N_12857,N_8177,N_11939);
or U12858 (N_12858,N_11790,N_10378);
or U12859 (N_12859,N_8852,N_9542);
or U12860 (N_12860,N_8625,N_11932);
or U12861 (N_12861,N_8077,N_9899);
and U12862 (N_12862,N_9527,N_8002);
nor U12863 (N_12863,N_11619,N_10161);
nor U12864 (N_12864,N_9094,N_8987);
or U12865 (N_12865,N_8815,N_9761);
and U12866 (N_12866,N_11354,N_11368);
or U12867 (N_12867,N_8143,N_10803);
nand U12868 (N_12868,N_8135,N_9223);
xnor U12869 (N_12869,N_10728,N_11436);
or U12870 (N_12870,N_11016,N_9677);
or U12871 (N_12871,N_10578,N_11215);
and U12872 (N_12872,N_10748,N_8846);
nor U12873 (N_12873,N_8043,N_10164);
nand U12874 (N_12874,N_10346,N_10468);
xor U12875 (N_12875,N_9591,N_11449);
nand U12876 (N_12876,N_8626,N_9336);
nor U12877 (N_12877,N_10391,N_11843);
or U12878 (N_12878,N_8095,N_8051);
nor U12879 (N_12879,N_8442,N_9299);
nor U12880 (N_12880,N_8220,N_8300);
nor U12881 (N_12881,N_10947,N_9270);
nand U12882 (N_12882,N_10192,N_9420);
and U12883 (N_12883,N_8723,N_10850);
nor U12884 (N_12884,N_10060,N_10067);
nor U12885 (N_12885,N_10156,N_8756);
and U12886 (N_12886,N_9689,N_11264);
or U12887 (N_12887,N_8809,N_8079);
or U12888 (N_12888,N_8673,N_10249);
and U12889 (N_12889,N_8129,N_8640);
nor U12890 (N_12890,N_10294,N_8329);
and U12891 (N_12891,N_8017,N_11366);
nor U12892 (N_12892,N_8099,N_10655);
or U12893 (N_12893,N_11292,N_9074);
nand U12894 (N_12894,N_9612,N_9251);
and U12895 (N_12895,N_11384,N_9297);
and U12896 (N_12896,N_8898,N_8082);
nor U12897 (N_12897,N_8879,N_8377);
and U12898 (N_12898,N_8847,N_8041);
nor U12899 (N_12899,N_10852,N_11183);
nor U12900 (N_12900,N_11637,N_11028);
nand U12901 (N_12901,N_9674,N_8460);
nand U12902 (N_12902,N_9008,N_10458);
and U12903 (N_12903,N_9550,N_10777);
nor U12904 (N_12904,N_9739,N_8136);
nor U12905 (N_12905,N_8457,N_10118);
and U12906 (N_12906,N_11551,N_8408);
or U12907 (N_12907,N_11221,N_10364);
nor U12908 (N_12908,N_10529,N_10464);
nand U12909 (N_12909,N_9212,N_11899);
nand U12910 (N_12910,N_8828,N_8085);
and U12911 (N_12911,N_11726,N_11279);
nand U12912 (N_12912,N_11326,N_8255);
or U12913 (N_12913,N_11768,N_9206);
nor U12914 (N_12914,N_11993,N_9641);
nand U12915 (N_12915,N_8985,N_11756);
or U12916 (N_12916,N_9703,N_9283);
nor U12917 (N_12917,N_8655,N_11429);
nand U12918 (N_12918,N_8940,N_10316);
nand U12919 (N_12919,N_11716,N_10318);
and U12920 (N_12920,N_10195,N_10681);
or U12921 (N_12921,N_8236,N_8931);
or U12922 (N_12922,N_11979,N_8919);
and U12923 (N_12923,N_9039,N_8400);
and U12924 (N_12924,N_9499,N_10392);
nand U12925 (N_12925,N_9719,N_11162);
and U12926 (N_12926,N_8491,N_8011);
nand U12927 (N_12927,N_10784,N_9991);
xnor U12928 (N_12928,N_8909,N_8332);
nor U12929 (N_12929,N_9779,N_8388);
nor U12930 (N_12930,N_9736,N_10144);
and U12931 (N_12931,N_10903,N_11488);
nand U12932 (N_12932,N_10119,N_11981);
and U12933 (N_12933,N_9528,N_8589);
or U12934 (N_12934,N_9495,N_11218);
xor U12935 (N_12935,N_11033,N_8314);
and U12936 (N_12936,N_8563,N_11416);
or U12937 (N_12937,N_8156,N_11819);
and U12938 (N_12938,N_9535,N_8253);
xor U12939 (N_12939,N_9493,N_9565);
or U12940 (N_12940,N_9602,N_8793);
and U12941 (N_12941,N_10749,N_10705);
and U12942 (N_12942,N_9430,N_11302);
nor U12943 (N_12943,N_8548,N_9477);
and U12944 (N_12944,N_10940,N_10265);
and U12945 (N_12945,N_11794,N_10647);
or U12946 (N_12946,N_10381,N_11336);
or U12947 (N_12947,N_11976,N_10791);
and U12948 (N_12948,N_11888,N_9104);
or U12949 (N_12949,N_11672,N_9211);
and U12950 (N_12950,N_10612,N_10268);
or U12951 (N_12951,N_11179,N_9894);
nand U12952 (N_12952,N_9357,N_8818);
nor U12953 (N_12953,N_10986,N_8657);
nand U12954 (N_12954,N_10896,N_10689);
and U12955 (N_12955,N_9525,N_11694);
nand U12956 (N_12956,N_8207,N_11414);
nand U12957 (N_12957,N_11441,N_9390);
or U12958 (N_12958,N_10600,N_11475);
and U12959 (N_12959,N_10871,N_8438);
nor U12960 (N_12960,N_11478,N_9734);
and U12961 (N_12961,N_11281,N_11320);
nand U12962 (N_12962,N_8333,N_11897);
nand U12963 (N_12963,N_9730,N_10541);
nor U12964 (N_12964,N_10398,N_10952);
and U12965 (N_12965,N_10833,N_10789);
nor U12966 (N_12966,N_9137,N_10718);
nand U12967 (N_12967,N_9879,N_11217);
and U12968 (N_12968,N_11130,N_11444);
or U12969 (N_12969,N_10536,N_9990);
nand U12970 (N_12970,N_10269,N_8829);
or U12971 (N_12971,N_8915,N_9566);
xnor U12972 (N_12972,N_9989,N_9626);
nand U12973 (N_12973,N_11675,N_8623);
nor U12974 (N_12974,N_10727,N_11424);
nor U12975 (N_12975,N_9983,N_9804);
and U12976 (N_12976,N_11214,N_10379);
nand U12977 (N_12977,N_10855,N_11135);
and U12978 (N_12978,N_10493,N_10827);
nor U12979 (N_12979,N_8904,N_8098);
or U12980 (N_12980,N_8998,N_9040);
and U12981 (N_12981,N_10183,N_8274);
and U12982 (N_12982,N_11283,N_10428);
nor U12983 (N_12983,N_8992,N_11793);
and U12984 (N_12984,N_8811,N_11204);
nor U12985 (N_12985,N_9735,N_11719);
nor U12986 (N_12986,N_8593,N_10964);
or U12987 (N_12987,N_9075,N_9839);
or U12988 (N_12988,N_11918,N_11889);
xnor U12989 (N_12989,N_9836,N_11346);
nor U12990 (N_12990,N_8558,N_8252);
or U12991 (N_12991,N_8243,N_9022);
and U12992 (N_12992,N_8091,N_10646);
xnor U12993 (N_12993,N_9816,N_10505);
and U12994 (N_12994,N_8103,N_11548);
xor U12995 (N_12995,N_10867,N_10476);
or U12996 (N_12996,N_11608,N_11804);
nand U12997 (N_12997,N_8743,N_9658);
or U12998 (N_12998,N_9107,N_11349);
nand U12999 (N_12999,N_11763,N_10544);
or U13000 (N_13000,N_8523,N_11759);
nand U13001 (N_13001,N_8310,N_11008);
nor U13002 (N_13002,N_9032,N_11434);
or U13003 (N_13003,N_11180,N_9393);
or U13004 (N_13004,N_9042,N_11484);
and U13005 (N_13005,N_10442,N_8055);
and U13006 (N_13006,N_11665,N_9595);
and U13007 (N_13007,N_9848,N_11741);
nand U13008 (N_13008,N_8600,N_11647);
nand U13009 (N_13009,N_11098,N_8482);
or U13010 (N_13010,N_9534,N_11009);
nor U13011 (N_13011,N_8654,N_10410);
or U13012 (N_13012,N_8148,N_8206);
nor U13013 (N_13013,N_10591,N_11848);
or U13014 (N_13014,N_9065,N_11601);
and U13015 (N_13015,N_9887,N_11481);
and U13016 (N_13016,N_8704,N_10955);
nand U13017 (N_13017,N_11157,N_11212);
nand U13018 (N_13018,N_11929,N_11640);
and U13019 (N_13019,N_10730,N_9077);
nor U13020 (N_13020,N_8822,N_10031);
nand U13021 (N_13021,N_10289,N_10849);
nor U13022 (N_13022,N_9081,N_8892);
nor U13023 (N_13023,N_8597,N_10804);
or U13024 (N_13024,N_9320,N_11752);
nand U13025 (N_13025,N_11923,N_11967);
nand U13026 (N_13026,N_8891,N_9095);
or U13027 (N_13027,N_9276,N_9584);
xnor U13028 (N_13028,N_8021,N_9082);
or U13029 (N_13029,N_9935,N_8481);
or U13030 (N_13030,N_9803,N_11578);
and U13031 (N_13031,N_10820,N_9691);
nand U13032 (N_13032,N_9833,N_11257);
nor U13033 (N_13033,N_9419,N_11985);
nand U13034 (N_13034,N_9947,N_9686);
or U13035 (N_13035,N_11811,N_8675);
or U13036 (N_13036,N_8959,N_9439);
or U13037 (N_13037,N_8323,N_11842);
or U13038 (N_13038,N_10509,N_8969);
nand U13039 (N_13039,N_10780,N_11893);
nor U13040 (N_13040,N_9530,N_11764);
nand U13041 (N_13041,N_11562,N_9843);
or U13042 (N_13042,N_10367,N_11933);
or U13043 (N_13043,N_9387,N_11903);
and U13044 (N_13044,N_10919,N_9905);
or U13045 (N_13045,N_9604,N_10982);
and U13046 (N_13046,N_8518,N_9915);
or U13047 (N_13047,N_10086,N_8418);
nand U13048 (N_13048,N_11917,N_11433);
nand U13049 (N_13049,N_10107,N_10214);
nor U13050 (N_13050,N_8728,N_8187);
nor U13051 (N_13051,N_9291,N_8275);
nor U13052 (N_13052,N_10455,N_9449);
nor U13053 (N_13053,N_9301,N_8434);
nor U13054 (N_13054,N_9748,N_11628);
or U13055 (N_13055,N_9556,N_9133);
or U13056 (N_13056,N_9950,N_8121);
and U13057 (N_13057,N_10413,N_9354);
and U13058 (N_13058,N_10001,N_11954);
and U13059 (N_13059,N_11371,N_11274);
nand U13060 (N_13060,N_9576,N_10373);
nor U13061 (N_13061,N_8947,N_11256);
nand U13062 (N_13062,N_11262,N_11137);
and U13063 (N_13063,N_11990,N_10559);
or U13064 (N_13064,N_9465,N_11237);
nand U13065 (N_13065,N_8899,N_10936);
nand U13066 (N_13066,N_10764,N_11696);
nor U13067 (N_13067,N_9720,N_9702);
and U13068 (N_13068,N_8195,N_10287);
nand U13069 (N_13069,N_10221,N_8096);
nand U13070 (N_13070,N_11583,N_9117);
and U13071 (N_13071,N_8086,N_11148);
nand U13072 (N_13072,N_10883,N_9073);
or U13073 (N_13073,N_10643,N_11387);
nand U13074 (N_13074,N_10527,N_9883);
nor U13075 (N_13075,N_8545,N_8917);
and U13076 (N_13076,N_9934,N_11448);
nand U13077 (N_13077,N_9834,N_11249);
nor U13078 (N_13078,N_9712,N_8286);
nand U13079 (N_13079,N_9144,N_11975);
nand U13080 (N_13080,N_10709,N_10554);
nand U13081 (N_13081,N_10736,N_10160);
or U13082 (N_13082,N_11400,N_10434);
nor U13083 (N_13083,N_9446,N_8924);
nor U13084 (N_13084,N_10595,N_10446);
and U13085 (N_13085,N_9621,N_10549);
nand U13086 (N_13086,N_9904,N_9280);
nand U13087 (N_13087,N_10051,N_11164);
or U13088 (N_13088,N_9443,N_10408);
or U13089 (N_13089,N_8707,N_10424);
or U13090 (N_13090,N_9132,N_10252);
and U13091 (N_13091,N_11750,N_11020);
nor U13092 (N_13092,N_9431,N_8857);
xnor U13093 (N_13093,N_11858,N_9268);
or U13094 (N_13094,N_11190,N_9762);
and U13095 (N_13095,N_9920,N_9266);
and U13096 (N_13096,N_11712,N_9302);
xnor U13097 (N_13097,N_11131,N_10925);
and U13098 (N_13098,N_10024,N_10642);
or U13099 (N_13099,N_10069,N_8084);
or U13100 (N_13100,N_9056,N_9597);
nand U13101 (N_13101,N_8324,N_9515);
and U13102 (N_13102,N_9239,N_10227);
nor U13103 (N_13103,N_11089,N_11621);
nand U13104 (N_13104,N_8754,N_8216);
nor U13105 (N_13105,N_8160,N_9422);
nor U13106 (N_13106,N_10907,N_10676);
and U13107 (N_13107,N_8399,N_10817);
nor U13108 (N_13108,N_9048,N_11801);
or U13109 (N_13109,N_11957,N_8175);
xor U13110 (N_13110,N_8006,N_8980);
nand U13111 (N_13111,N_10096,N_11178);
or U13112 (N_13112,N_8982,N_8375);
and U13113 (N_13113,N_9961,N_11603);
nand U13114 (N_13114,N_9021,N_9111);
nand U13115 (N_13115,N_9064,N_11787);
nor U13116 (N_13116,N_8808,N_9824);
and U13117 (N_13117,N_8350,N_9801);
and U13118 (N_13118,N_11391,N_10677);
and U13119 (N_13119,N_8974,N_8731);
and U13120 (N_13120,N_11355,N_9704);
nand U13121 (N_13121,N_9370,N_8914);
xnor U13122 (N_13122,N_11004,N_9668);
and U13123 (N_13123,N_8087,N_8514);
and U13124 (N_13124,N_9874,N_10257);
nor U13125 (N_13125,N_10436,N_9161);
nor U13126 (N_13126,N_8228,N_10812);
and U13127 (N_13127,N_11635,N_8725);
nor U13128 (N_13128,N_9964,N_9699);
nand U13129 (N_13129,N_11386,N_9274);
or U13130 (N_13130,N_8005,N_8283);
and U13131 (N_13131,N_8436,N_11689);
nor U13132 (N_13132,N_8637,N_10834);
nand U13133 (N_13133,N_8592,N_10308);
nand U13134 (N_13134,N_11905,N_10299);
nand U13135 (N_13135,N_10916,N_10930);
and U13136 (N_13136,N_11019,N_8259);
and U13137 (N_13137,N_9785,N_9672);
nand U13138 (N_13138,N_11027,N_8166);
or U13139 (N_13139,N_9051,N_9455);
nor U13140 (N_13140,N_11328,N_9670);
and U13141 (N_13141,N_9436,N_8444);
xor U13142 (N_13142,N_11464,N_8081);
nand U13143 (N_13143,N_9973,N_11627);
or U13144 (N_13144,N_9105,N_8648);
nand U13145 (N_13145,N_8202,N_11871);
nor U13146 (N_13146,N_8458,N_10631);
or U13147 (N_13147,N_8322,N_8317);
xor U13148 (N_13148,N_11930,N_8395);
nand U13149 (N_13149,N_11650,N_10077);
nand U13150 (N_13150,N_9860,N_8521);
or U13151 (N_13151,N_9603,N_11417);
and U13152 (N_13152,N_11024,N_10918);
nor U13153 (N_13153,N_11655,N_10725);
and U13154 (N_13154,N_9464,N_10194);
or U13155 (N_13155,N_11312,N_9197);
or U13156 (N_13156,N_10970,N_8311);
or U13157 (N_13157,N_9327,N_11299);
or U13158 (N_13158,N_9589,N_9328);
nand U13159 (N_13159,N_8963,N_9784);
nor U13160 (N_13160,N_9366,N_10143);
or U13161 (N_13161,N_8537,N_8365);
nor U13162 (N_13162,N_8669,N_10320);
or U13163 (N_13163,N_10018,N_9965);
nand U13164 (N_13164,N_9729,N_10597);
nor U13165 (N_13165,N_9886,N_10698);
nand U13166 (N_13166,N_9359,N_11393);
nor U13167 (N_13167,N_11497,N_10522);
nor U13168 (N_13168,N_11392,N_8685);
or U13169 (N_13169,N_9680,N_10781);
nor U13170 (N_13170,N_9832,N_11755);
or U13171 (N_13171,N_8812,N_11076);
nor U13172 (N_13172,N_10516,N_10956);
nor U13173 (N_13173,N_11419,N_9910);
or U13174 (N_13174,N_10469,N_8061);
and U13175 (N_13175,N_10224,N_10487);
nor U13176 (N_13176,N_10177,N_8894);
and U13177 (N_13177,N_11690,N_9655);
or U13178 (N_13178,N_10787,N_9617);
nand U13179 (N_13179,N_9382,N_8094);
and U13180 (N_13180,N_11579,N_8553);
and U13181 (N_13181,N_10040,N_11208);
nor U13182 (N_13182,N_8480,N_11022);
and U13183 (N_13183,N_11115,N_11835);
or U13184 (N_13184,N_10802,N_10206);
and U13185 (N_13185,N_9846,N_11698);
and U13186 (N_13186,N_9267,N_10124);
nor U13187 (N_13187,N_8171,N_11847);
nor U13188 (N_13188,N_10330,N_9684);
or U13189 (N_13189,N_11418,N_11898);
or U13190 (N_13190,N_11830,N_11928);
and U13191 (N_13191,N_10686,N_10719);
nand U13192 (N_13192,N_8752,N_11191);
nor U13193 (N_13193,N_11113,N_9168);
and U13194 (N_13194,N_11558,N_9545);
or U13195 (N_13195,N_10699,N_8560);
nand U13196 (N_13196,N_11106,N_10382);
and U13197 (N_13197,N_8638,N_8064);
xnor U13198 (N_13198,N_10741,N_10204);
nor U13199 (N_13199,N_8214,N_9914);
or U13200 (N_13200,N_9986,N_8708);
and U13201 (N_13201,N_8144,N_8188);
or U13202 (N_13202,N_9441,N_8767);
or U13203 (N_13203,N_8878,N_11799);
xor U13204 (N_13204,N_8501,N_11243);
nor U13205 (N_13205,N_10758,N_11289);
nand U13206 (N_13206,N_8152,N_10407);
and U13207 (N_13207,N_11251,N_10897);
nand U13208 (N_13208,N_10768,N_11857);
and U13209 (N_13209,N_10032,N_10197);
nand U13210 (N_13210,N_8013,N_9900);
or U13211 (N_13211,N_11435,N_8357);
nor U13212 (N_13212,N_10351,N_11971);
and U13213 (N_13213,N_10116,N_8306);
and U13214 (N_13214,N_8224,N_9861);
nor U13215 (N_13215,N_9278,N_10831);
and U13216 (N_13216,N_9605,N_8609);
and U13217 (N_13217,N_11078,N_8676);
nor U13218 (N_13218,N_10668,N_11116);
nor U13219 (N_13219,N_11966,N_8403);
nand U13220 (N_13220,N_8409,N_9580);
nor U13221 (N_13221,N_10616,N_11305);
and U13222 (N_13222,N_8948,N_8999);
nor U13223 (N_13223,N_10605,N_11465);
nor U13224 (N_13224,N_11534,N_11500);
and U13225 (N_13225,N_8839,N_8840);
and U13226 (N_13226,N_9640,N_8551);
or U13227 (N_13227,N_9237,N_8912);
or U13228 (N_13228,N_8130,N_8550);
or U13229 (N_13229,N_11861,N_11674);
nand U13230 (N_13230,N_8340,N_11490);
and U13231 (N_13231,N_10333,N_11385);
and U13232 (N_13232,N_11037,N_9789);
nand U13233 (N_13233,N_8881,N_8633);
and U13234 (N_13234,N_9127,N_10178);
and U13235 (N_13235,N_8738,N_8046);
nor U13236 (N_13236,N_11587,N_10171);
and U13237 (N_13237,N_10324,N_10120);
or U13238 (N_13238,N_10021,N_10477);
and U13239 (N_13239,N_10533,N_10226);
nor U13240 (N_13240,N_11377,N_11945);
and U13241 (N_13241,N_11451,N_11463);
nand U13242 (N_13242,N_8977,N_10419);
or U13243 (N_13243,N_10203,N_9743);
and U13244 (N_13244,N_8427,N_8459);
nor U13245 (N_13245,N_8740,N_9746);
nand U13246 (N_13246,N_9054,N_9185);
or U13247 (N_13247,N_9498,N_11541);
or U13248 (N_13248,N_11314,N_9261);
nor U13249 (N_13249,N_11717,N_10162);
or U13250 (N_13250,N_11666,N_8217);
or U13251 (N_13251,N_8603,N_11271);
or U13252 (N_13252,N_10159,N_8050);
and U13253 (N_13253,N_10050,N_11659);
xnor U13254 (N_13254,N_10793,N_11521);
nor U13255 (N_13255,N_9975,N_8533);
and U13256 (N_13256,N_8627,N_10443);
or U13257 (N_13257,N_11596,N_9346);
nand U13258 (N_13258,N_9901,N_9060);
nand U13259 (N_13259,N_11563,N_11556);
nor U13260 (N_13260,N_8000,N_10121);
nand U13261 (N_13261,N_11151,N_8918);
or U13262 (N_13262,N_10708,N_11661);
or U13263 (N_13263,N_10020,N_8052);
nand U13264 (N_13264,N_9337,N_11295);
nor U13265 (N_13265,N_8876,N_8270);
and U13266 (N_13266,N_10661,N_10250);
and U13267 (N_13267,N_11582,N_9847);
and U13268 (N_13268,N_11125,N_11522);
or U13269 (N_13269,N_11512,N_9396);
nor U13270 (N_13270,N_10013,N_8984);
and U13271 (N_13271,N_10662,N_10369);
nor U13272 (N_13272,N_8150,N_9055);
nor U13273 (N_13273,N_9013,N_8476);
nand U13274 (N_13274,N_9487,N_10813);
nand U13275 (N_13275,N_9930,N_9561);
nor U13276 (N_13276,N_10997,N_9962);
nor U13277 (N_13277,N_8775,N_8025);
nand U13278 (N_13278,N_11460,N_9482);
and U13279 (N_13279,N_8721,N_8744);
and U13280 (N_13280,N_8802,N_9685);
or U13281 (N_13281,N_11798,N_11495);
or U13282 (N_13282,N_11322,N_10696);
nand U13283 (N_13283,N_9698,N_8271);
or U13284 (N_13284,N_10508,N_10212);
and U13285 (N_13285,N_8620,N_10770);
and U13286 (N_13286,N_9156,N_11813);
nor U13287 (N_13287,N_8372,N_10113);
or U13288 (N_13288,N_8361,N_10172);
nor U13289 (N_13289,N_10492,N_10459);
nor U13290 (N_13290,N_8326,N_11427);
or U13291 (N_13291,N_10691,N_8659);
or U13292 (N_13292,N_11984,N_9189);
or U13293 (N_13293,N_11067,N_10707);
or U13294 (N_13294,N_11699,N_11921);
or U13295 (N_13295,N_10990,N_8525);
nand U13296 (N_13296,N_10068,N_11740);
and U13297 (N_13297,N_9711,N_11252);
or U13298 (N_13298,N_10659,N_8371);
nand U13299 (N_13299,N_9491,N_8981);
or U13300 (N_13300,N_8254,N_9929);
or U13301 (N_13301,N_10540,N_10180);
or U13302 (N_13302,N_11882,N_8298);
and U13303 (N_13303,N_11176,N_10628);
nand U13304 (N_13304,N_8034,N_9873);
or U13305 (N_13305,N_10475,N_9338);
or U13306 (N_13306,N_8733,N_10868);
nand U13307 (N_13307,N_9006,N_10887);
nand U13308 (N_13308,N_9331,N_10105);
or U13309 (N_13309,N_8256,N_10377);
and U13310 (N_13310,N_9035,N_11739);
and U13311 (N_13311,N_10182,N_11184);
nand U13312 (N_13312,N_9496,N_8269);
nor U13313 (N_13313,N_11267,N_10950);
nand U13314 (N_13314,N_11970,N_8246);
nor U13315 (N_13315,N_11594,N_10783);
or U13316 (N_13316,N_9199,N_11926);
or U13317 (N_13317,N_8431,N_9141);
xor U13318 (N_13318,N_8646,N_8505);
and U13319 (N_13319,N_10545,N_8535);
xnor U13320 (N_13320,N_11052,N_10207);
and U13321 (N_13321,N_9692,N_10471);
and U13322 (N_13322,N_8791,N_8389);
nand U13323 (N_13323,N_9305,N_8686);
nor U13324 (N_13324,N_11994,N_8200);
nor U13325 (N_13325,N_9281,N_10515);
nand U13326 (N_13326,N_11996,N_10403);
nor U13327 (N_13327,N_10092,N_9741);
nor U13328 (N_13328,N_9025,N_11864);
nor U13329 (N_13329,N_8366,N_8137);
and U13330 (N_13330,N_10231,N_8302);
nand U13331 (N_13331,N_11453,N_10321);
and U13332 (N_13332,N_10713,N_10774);
and U13333 (N_13333,N_8303,N_11253);
nand U13334 (N_13334,N_10117,N_9772);
nand U13335 (N_13335,N_11432,N_8629);
and U13336 (N_13336,N_9425,N_11234);
nor U13337 (N_13337,N_10927,N_10411);
nor U13338 (N_13338,N_8343,N_9169);
or U13339 (N_13339,N_8393,N_11053);
or U13340 (N_13340,N_9429,N_8415);
nand U13341 (N_13341,N_8124,N_10856);
nand U13342 (N_13342,N_10779,N_11757);
and U13343 (N_13343,N_10003,N_9518);
and U13344 (N_13344,N_10621,N_9269);
or U13345 (N_13345,N_11132,N_10463);
or U13346 (N_13346,N_8425,N_9226);
nor U13347 (N_13347,N_8147,N_11677);
and U13348 (N_13348,N_11910,N_11707);
or U13349 (N_13349,N_11380,N_10148);
nand U13350 (N_13350,N_10798,N_9958);
nand U13351 (N_13351,N_8824,N_9613);
and U13352 (N_13352,N_8391,N_9631);
and U13353 (N_13353,N_10507,N_11012);
nor U13354 (N_13354,N_10975,N_8462);
and U13355 (N_13355,N_9512,N_8753);
or U13356 (N_13356,N_11838,N_8757);
nor U13357 (N_13357,N_11753,N_11815);
xor U13358 (N_13358,N_8170,N_9353);
nor U13359 (N_13359,N_11158,N_8248);
nand U13360 (N_13360,N_10673,N_9516);
and U13361 (N_13361,N_10230,N_10682);
nor U13362 (N_13362,N_8219,N_11974);
and U13363 (N_13363,N_11544,N_10922);
nand U13364 (N_13364,N_9776,N_8024);
nor U13365 (N_13365,N_10062,N_11960);
nand U13366 (N_13366,N_11259,N_9134);
nand U13367 (N_13367,N_8267,N_8510);
and U13368 (N_13368,N_9412,N_11068);
and U13369 (N_13369,N_9198,N_11405);
and U13370 (N_13370,N_8174,N_10603);
nand U13371 (N_13371,N_10259,N_9852);
and U13372 (N_13372,N_11528,N_10843);
and U13373 (N_13373,N_8059,N_9209);
and U13374 (N_13374,N_8979,N_8875);
nor U13375 (N_13375,N_11077,N_8872);
nor U13376 (N_13376,N_9046,N_8291);
or U13377 (N_13377,N_8509,N_11774);
nand U13378 (N_13378,N_11821,N_11174);
nand U13379 (N_13379,N_9643,N_9970);
and U13380 (N_13380,N_8169,N_8417);
and U13381 (N_13381,N_11734,N_11491);
or U13382 (N_13382,N_10630,N_9543);
or U13383 (N_13383,N_11826,N_8584);
and U13384 (N_13384,N_10640,N_9778);
or U13385 (N_13385,N_10967,N_8759);
and U13386 (N_13386,N_9837,N_11937);
nand U13387 (N_13387,N_10574,N_8044);
and U13388 (N_13388,N_8996,N_8885);
nor U13389 (N_13389,N_10703,N_9224);
nor U13390 (N_13390,N_9324,N_8068);
or U13391 (N_13391,N_11316,N_9726);
and U13392 (N_13392,N_11408,N_10023);
nor U13393 (N_13393,N_9427,N_10808);
and U13394 (N_13394,N_11395,N_9532);
and U13395 (N_13395,N_11878,N_8123);
and U13396 (N_13396,N_11877,N_9479);
nand U13397 (N_13397,N_10305,N_11516);
and U13398 (N_13398,N_10246,N_8782);
and U13399 (N_13399,N_11833,N_11474);
nand U13400 (N_13400,N_8193,N_9005);
or U13401 (N_13401,N_8821,N_11136);
nand U13402 (N_13402,N_8422,N_8823);
or U13403 (N_13403,N_11961,N_9303);
or U13404 (N_13404,N_11613,N_9695);
or U13405 (N_13405,N_8886,N_8354);
and U13406 (N_13406,N_9452,N_9045);
and U13407 (N_13407,N_10186,N_11779);
or U13408 (N_13408,N_10914,N_9884);
nor U13409 (N_13409,N_8119,N_10657);
nor U13410 (N_13410,N_10679,N_9560);
and U13411 (N_13411,N_11651,N_9201);
nand U13412 (N_13412,N_10063,N_9150);
or U13413 (N_13413,N_8483,N_10575);
nor U13414 (N_13414,N_10271,N_11109);
or U13415 (N_13415,N_11245,N_10745);
or U13416 (N_13416,N_10981,N_8076);
nand U13417 (N_13417,N_9713,N_11633);
xnor U13418 (N_13418,N_10247,N_9610);
nand U13419 (N_13419,N_11706,N_9145);
or U13420 (N_13420,N_10152,N_11080);
or U13421 (N_13421,N_9325,N_8178);
and U13422 (N_13422,N_11046,N_10427);
nor U13423 (N_13423,N_11142,N_9908);
xnor U13424 (N_13424,N_8090,N_8466);
and U13425 (N_13425,N_11149,N_9892);
and U13426 (N_13426,N_9500,N_9044);
or U13427 (N_13427,N_8114,N_10217);
or U13428 (N_13428,N_9400,N_11892);
or U13429 (N_13429,N_9898,N_10889);
or U13430 (N_13430,N_8670,N_8497);
and U13431 (N_13431,N_9531,N_11025);
nand U13432 (N_13432,N_10920,N_8679);
nor U13433 (N_13433,N_8405,N_10778);
nand U13434 (N_13434,N_11646,N_8461);
nand U13435 (N_13435,N_9410,N_9401);
nor U13436 (N_13436,N_8106,N_9814);
nor U13437 (N_13437,N_10526,N_11977);
nand U13438 (N_13438,N_11061,N_9348);
nand U13439 (N_13439,N_11758,N_10309);
and U13440 (N_13440,N_11721,N_11657);
nand U13441 (N_13441,N_9173,N_11622);
and U13442 (N_13442,N_9862,N_10872);
or U13443 (N_13443,N_10478,N_8594);
and U13444 (N_13444,N_9583,N_10992);
nand U13445 (N_13445,N_11998,N_9435);
or U13446 (N_13446,N_10248,N_8769);
or U13447 (N_13447,N_11270,N_8624);
nand U13448 (N_13448,N_11483,N_9727);
or U13449 (N_13449,N_9826,N_11141);
nand U13450 (N_13450,N_10996,N_11422);
or U13451 (N_13451,N_8661,N_8353);
nor U13452 (N_13452,N_10771,N_10641);
or U13453 (N_13453,N_11900,N_9235);
nor U13454 (N_13454,N_9590,N_11965);
nor U13455 (N_13455,N_8028,N_9754);
or U13456 (N_13456,N_9752,N_10006);
or U13457 (N_13457,N_8630,N_10944);
nand U13458 (N_13458,N_9097,N_11471);
or U13459 (N_13459,N_10788,N_9061);
nor U13460 (N_13460,N_10251,N_11729);
and U13461 (N_13461,N_11081,N_9275);
or U13462 (N_13462,N_11315,N_11187);
or U13463 (N_13463,N_8699,N_10632);
nor U13464 (N_13464,N_9485,N_9242);
and U13465 (N_13465,N_11683,N_11069);
nand U13466 (N_13466,N_10582,N_10196);
nand U13467 (N_13467,N_9744,N_10337);
xor U13468 (N_13468,N_9971,N_8842);
nand U13469 (N_13469,N_9136,N_8636);
and U13470 (N_13470,N_11617,N_8905);
or U13471 (N_13471,N_8543,N_10303);
nand U13472 (N_13472,N_8020,N_8508);
nand U13473 (N_13473,N_11189,N_9728);
nor U13474 (N_13474,N_10694,N_11207);
nand U13475 (N_13475,N_11588,N_8033);
nor U13476 (N_13476,N_8866,N_9361);
and U13477 (N_13477,N_8662,N_9912);
and U13478 (N_13478,N_10858,N_9087);
nor U13479 (N_13479,N_9093,N_9319);
or U13480 (N_13480,N_11543,N_9755);
and U13481 (N_13481,N_11357,N_9339);
nor U13482 (N_13482,N_8889,N_10819);
nor U13483 (N_13483,N_9256,N_10946);
or U13484 (N_13484,N_10488,N_10438);
and U13485 (N_13485,N_10285,N_10115);
nor U13486 (N_13486,N_8750,N_10556);
and U13487 (N_13487,N_9551,N_9341);
nand U13488 (N_13488,N_11105,N_10814);
or U13489 (N_13489,N_9763,N_9344);
nor U13490 (N_13490,N_8203,N_10084);
and U13491 (N_13491,N_9637,N_9838);
or U13492 (N_13492,N_11936,N_9870);
or U13493 (N_13493,N_9101,N_8833);
or U13494 (N_13494,N_11571,N_8153);
nor U13495 (N_13495,N_10873,N_9808);
nand U13496 (N_13496,N_8801,N_11983);
nor U13497 (N_13497,N_8565,N_10760);
nor U13498 (N_13498,N_9995,N_9321);
or U13499 (N_13499,N_8053,N_9330);
nand U13500 (N_13500,N_9252,N_11390);
or U13501 (N_13501,N_9567,N_11745);
nand U13502 (N_13502,N_10891,N_9316);
nor U13503 (N_13503,N_9090,N_11341);
and U13504 (N_13504,N_11042,N_10830);
or U13505 (N_13505,N_8540,N_9405);
or U13506 (N_13506,N_8180,N_11195);
nand U13507 (N_13507,N_10627,N_8154);
and U13508 (N_13508,N_11863,N_8105);
nand U13509 (N_13509,N_10932,N_8364);
nand U13510 (N_13510,N_11948,N_8901);
or U13511 (N_13511,N_10623,N_8242);
and U13512 (N_13512,N_9085,N_9549);
nand U13513 (N_13513,N_11064,N_10969);
or U13514 (N_13514,N_11671,N_8209);
and U13515 (N_13515,N_11397,N_10531);
xnor U13516 (N_13516,N_10240,N_10371);
nand U13517 (N_13517,N_10991,N_8134);
and U13518 (N_13518,N_11325,N_11920);
nand U13519 (N_13519,N_11822,N_10829);
and U13520 (N_13520,N_8176,N_8339);
xnor U13521 (N_13521,N_10596,N_10352);
and U13522 (N_13522,N_10317,N_10104);
nor U13523 (N_13523,N_10087,N_11856);
nand U13524 (N_13524,N_11054,N_9943);
and U13525 (N_13525,N_9099,N_10697);
or U13526 (N_13526,N_8722,N_11751);
or U13527 (N_13527,N_8581,N_9615);
nor U13528 (N_13528,N_8710,N_9937);
and U13529 (N_13529,N_10894,N_9408);
and U13530 (N_13530,N_10027,N_11056);
or U13531 (N_13531,N_11566,N_11049);
nor U13532 (N_13532,N_9966,N_9041);
nand U13533 (N_13533,N_10638,N_9629);
nor U13534 (N_13534,N_8768,N_11265);
or U13535 (N_13535,N_10342,N_11090);
nand U13536 (N_13536,N_10447,N_10332);
nor U13537 (N_13537,N_8606,N_10520);
nor U13538 (N_13538,N_11829,N_11913);
nand U13539 (N_13539,N_11533,N_9453);
nand U13540 (N_13540,N_8582,N_8936);
nor U13541 (N_13541,N_9759,N_9460);
nor U13542 (N_13542,N_9972,N_10823);
nor U13543 (N_13543,N_10649,N_10472);
or U13544 (N_13544,N_10669,N_10594);
nor U13545 (N_13545,N_9286,N_9519);
nand U13546 (N_13546,N_8864,N_9890);
and U13547 (N_13547,N_10384,N_11439);
nand U13548 (N_13548,N_9407,N_8402);
and U13549 (N_13549,N_10415,N_9238);
or U13550 (N_13550,N_10870,N_11345);
and U13551 (N_13551,N_9931,N_8945);
nand U13552 (N_13552,N_10128,N_10409);
and U13553 (N_13553,N_8048,N_11780);
nand U13554 (N_13554,N_10906,N_11071);
nor U13555 (N_13555,N_9345,N_10274);
or U13556 (N_13556,N_11867,N_9985);
xor U13557 (N_13557,N_11356,N_11381);
nand U13558 (N_13558,N_9070,N_8678);
and U13559 (N_13559,N_11597,N_11695);
nor U13560 (N_13560,N_10208,N_9897);
nor U13561 (N_13561,N_10564,N_9978);
nor U13562 (N_13562,N_9009,N_10979);
nor U13563 (N_13563,N_11045,N_9356);
nor U13564 (N_13564,N_10039,N_11632);
and U13565 (N_13565,N_10511,N_8700);
nor U13566 (N_13566,N_9625,N_11095);
and U13567 (N_13567,N_11854,N_9806);
nand U13568 (N_13568,N_11255,N_10209);
or U13569 (N_13569,N_8617,N_8263);
nand U13570 (N_13570,N_8194,N_9553);
nand U13571 (N_13571,N_8776,N_8159);
nor U13572 (N_13572,N_10151,N_8647);
nor U13573 (N_13573,N_11450,N_11026);
or U13574 (N_13574,N_9300,N_8957);
or U13575 (N_13575,N_11360,N_8019);
or U13576 (N_13576,N_10362,N_10651);
nor U13577 (N_13577,N_8500,N_10288);
nor U13578 (N_13578,N_8308,N_11118);
nand U13579 (N_13579,N_11462,N_11946);
nand U13580 (N_13580,N_10165,N_11730);
nand U13581 (N_13581,N_9318,N_8703);
or U13582 (N_13582,N_9123,N_8484);
nand U13583 (N_13583,N_8709,N_11023);
or U13584 (N_13584,N_11144,N_10711);
nor U13585 (N_13585,N_11846,N_10383);
nand U13586 (N_13586,N_11769,N_11773);
and U13587 (N_13587,N_10598,N_8542);
nor U13588 (N_13588,N_9033,N_8856);
and U13589 (N_13589,N_11997,N_11620);
and U13590 (N_13590,N_9373,N_8139);
and U13591 (N_13591,N_9418,N_8778);
and U13592 (N_13592,N_8014,N_10157);
or U13593 (N_13593,N_8470,N_9812);
nand U13594 (N_13594,N_8304,N_9733);
nor U13595 (N_13595,N_9034,N_8428);
and U13596 (N_13596,N_11598,N_9049);
nand U13597 (N_13597,N_8893,N_8615);
nand U13598 (N_13598,N_8522,N_10017);
or U13599 (N_13599,N_9470,N_11159);
nand U13600 (N_13600,N_10706,N_11736);
nor U13601 (N_13601,N_9652,N_10012);
and U13602 (N_13602,N_10532,N_8619);
nor U13603 (N_13603,N_10284,N_8515);
nand U13604 (N_13604,N_8397,N_8075);
nand U13605 (N_13605,N_9976,N_11818);
nor U13606 (N_13606,N_10482,N_11581);
nor U13607 (N_13607,N_11296,N_10731);
and U13608 (N_13608,N_9152,N_8746);
and U13609 (N_13609,N_9329,N_10075);
nor U13610 (N_13610,N_11224,N_9888);
nor U13611 (N_13611,N_11223,N_11388);
or U13612 (N_13612,N_10790,N_10375);
nand U13613 (N_13613,N_11139,N_11319);
nand U13614 (N_13614,N_10583,N_9364);
or U13615 (N_13615,N_9335,N_11592);
nand U13616 (N_13616,N_9375,N_11059);
nand U13617 (N_13617,N_10840,N_8971);
and U13618 (N_13618,N_11504,N_10957);
xnor U13619 (N_13619,N_8261,N_9577);
nand U13620 (N_13620,N_8336,N_8370);
and U13621 (N_13621,N_10723,N_10273);
nor U13622 (N_13622,N_11277,N_8526);
or U13623 (N_13623,N_10720,N_9818);
nand U13624 (N_13624,N_8813,N_11911);
nor U13625 (N_13625,N_9079,N_10879);
or U13626 (N_13626,N_8001,N_11018);
nor U13627 (N_13627,N_11211,N_10753);
or U13628 (N_13628,N_8868,N_10888);
or U13629 (N_13629,N_8184,N_8290);
or U13630 (N_13630,N_11614,N_10101);
nand U13631 (N_13631,N_9721,N_11363);
nor U13632 (N_13632,N_10090,N_8301);
nor U13633 (N_13633,N_8580,N_8265);
nor U13634 (N_13634,N_9200,N_10238);
nand U13635 (N_13635,N_9758,N_10902);
nand U13636 (N_13636,N_11167,N_9996);
or U13637 (N_13637,N_8724,N_11200);
and U13638 (N_13638,N_8213,N_10857);
and U13639 (N_13639,N_10322,N_9289);
nor U13640 (N_13640,N_9468,N_9850);
or U13641 (N_13641,N_8398,N_8730);
nand U13642 (N_13642,N_8453,N_8939);
nand U13643 (N_13643,N_9828,N_9228);
or U13644 (N_13644,N_9671,N_10599);
nand U13645 (N_13645,N_10218,N_8666);
nor U13646 (N_13646,N_11938,N_8433);
or U13647 (N_13647,N_8681,N_9786);
nand U13648 (N_13648,N_10799,N_11493);
nor U13649 (N_13649,N_10740,N_9380);
nand U13650 (N_13650,N_10053,N_11327);
nand U13651 (N_13651,N_8642,N_11881);
and U13652 (N_13652,N_10435,N_11572);
and U13653 (N_13653,N_11761,N_11048);
and U13654 (N_13654,N_11447,N_8546);
nor U13655 (N_13655,N_9841,N_8855);
and U13656 (N_13656,N_11860,N_9170);
nor U13657 (N_13657,N_9416,N_10542);
nor U13658 (N_13658,N_10138,N_11959);
and U13659 (N_13659,N_9724,N_11093);
nor U13660 (N_13660,N_9864,N_10861);
nand U13661 (N_13661,N_11746,N_8475);
nor U13662 (N_13662,N_8378,N_11630);
or U13663 (N_13663,N_10281,N_11812);
or U13664 (N_13664,N_11615,N_9588);
and U13665 (N_13665,N_8266,N_10684);
or U13666 (N_13666,N_11087,N_8282);
nor U13667 (N_13667,N_11737,N_10345);
nor U13668 (N_13668,N_9480,N_8605);
nor U13669 (N_13669,N_11403,N_8477);
or U13670 (N_13670,N_11231,N_8944);
or U13671 (N_13671,N_10136,N_8190);
or U13672 (N_13672,N_9794,N_9769);
or U13673 (N_13673,N_8439,N_10454);
nor U13674 (N_13674,N_11005,N_9203);
nand U13675 (N_13675,N_10908,N_11931);
or U13676 (N_13676,N_9539,N_11883);
and U13677 (N_13677,N_9859,N_10550);
nand U13678 (N_13678,N_11591,N_8330);
nand U13679 (N_13679,N_10983,N_8527);
nor U13680 (N_13680,N_9218,N_8109);
xnor U13681 (N_13681,N_8651,N_11060);
nor U13682 (N_13682,N_8588,N_10370);
or U13683 (N_13683,N_10283,N_9205);
nand U13684 (N_13684,N_9938,N_8729);
or U13685 (N_13685,N_8621,N_10126);
nor U13686 (N_13686,N_9765,N_9157);
and U13687 (N_13687,N_9570,N_9750);
or U13688 (N_13688,N_8665,N_8112);
nand U13689 (N_13689,N_9195,N_8649);
or U13690 (N_13690,N_11161,N_8205);
and U13691 (N_13691,N_8530,N_10350);
nor U13692 (N_13692,N_10243,N_8083);
nand U13693 (N_13693,N_10254,N_8173);
nand U13694 (N_13694,N_10604,N_10395);
and U13695 (N_13695,N_9295,N_10223);
or U13696 (N_13696,N_11539,N_11537);
nor U13697 (N_13697,N_10613,N_9298);
nor U13698 (N_13698,N_9020,N_9186);
nand U13699 (N_13699,N_8652,N_8128);
or U13700 (N_13700,N_10376,N_8140);
or U13701 (N_13701,N_10334,N_11988);
or U13702 (N_13702,N_8964,N_10047);
xor U13703 (N_13703,N_8695,N_11785);
nor U13704 (N_13704,N_9511,N_8247);
nor U13705 (N_13705,N_9050,N_11275);
and U13706 (N_13706,N_9510,N_9246);
or U13707 (N_13707,N_11194,N_11254);
nand U13708 (N_13708,N_10976,N_10005);
nand U13709 (N_13709,N_10960,N_11704);
nand U13710 (N_13710,N_11321,N_10170);
or U13711 (N_13711,N_11411,N_10663);
nand U13712 (N_13712,N_10726,N_9308);
nand U13713 (N_13713,N_9732,N_11492);
nand U13714 (N_13714,N_9951,N_8726);
nand U13715 (N_13715,N_11969,N_9559);
and U13716 (N_13716,N_10145,N_11738);
nand U13717 (N_13717,N_10292,N_11808);
and U13718 (N_13718,N_8468,N_9569);
and U13719 (N_13719,N_11344,N_9650);
nor U13720 (N_13720,N_10359,N_8162);
nor U13721 (N_13721,N_8942,N_8141);
nor U13722 (N_13722,N_8916,N_10089);
nor U13723 (N_13723,N_9063,N_10449);
nand U13724 (N_13724,N_10524,N_10836);
nand U13725 (N_13725,N_8853,N_10106);
or U13726 (N_13726,N_9540,N_8850);
nor U13727 (N_13727,N_8218,N_10977);
nand U13728 (N_13728,N_10566,N_10637);
nor U13729 (N_13729,N_11246,N_9587);
and U13730 (N_13730,N_8519,N_10687);
and U13731 (N_13731,N_8949,N_9663);
or U13732 (N_13732,N_10199,N_8430);
nand U13733 (N_13733,N_8873,N_10348);
nand U13734 (N_13734,N_10222,N_10191);
nor U13735 (N_13735,N_11485,N_8107);
nand U13736 (N_13736,N_9255,N_10560);
nand U13737 (N_13737,N_8607,N_11749);
xnor U13738 (N_13738,N_9368,N_10073);
or U13739 (N_13739,N_9263,N_10034);
and U13740 (N_13740,N_9445,N_8437);
and U13741 (N_13741,N_8817,N_9647);
nor U13742 (N_13742,N_10576,N_11866);
and U13743 (N_13743,N_10188,N_10213);
or U13744 (N_13744,N_9829,N_11987);
nor U13745 (N_13745,N_9296,N_10202);
or U13746 (N_13746,N_11044,N_10420);
nand U13747 (N_13747,N_8294,N_10626);
nor U13748 (N_13748,N_8414,N_10033);
nor U13749 (N_13749,N_11352,N_11021);
and U13750 (N_13750,N_10129,N_9863);
or U13751 (N_13751,N_10797,N_11374);
nand U13752 (N_13752,N_10503,N_10429);
or U13753 (N_13753,N_9215,N_9681);
nor U13754 (N_13754,N_10431,N_11600);
or U13755 (N_13755,N_9247,N_9392);
or U13756 (N_13756,N_11425,N_11559);
nor U13757 (N_13757,N_9557,N_9159);
nand U13758 (N_13758,N_10563,N_8628);
and U13759 (N_13759,N_10675,N_8268);
nor U13760 (N_13760,N_9043,N_8874);
nor U13761 (N_13761,N_10847,N_10329);
or U13762 (N_13762,N_8118,N_8441);
or U13763 (N_13763,N_9071,N_10690);
nor U13764 (N_13764,N_11273,N_11820);
or U13765 (N_13765,N_10588,N_9813);
nand U13766 (N_13766,N_11765,N_8189);
nor U13767 (N_13767,N_9902,N_8238);
nand U13768 (N_13768,N_8182,N_11206);
nor U13769 (N_13769,N_9249,N_9437);
nor U13770 (N_13770,N_8585,N_8639);
and U13771 (N_13771,N_8325,N_9140);
xnor U13772 (N_13772,N_11373,N_9171);
nor U13773 (N_13773,N_11030,N_10358);
and U13774 (N_13774,N_10485,N_11781);
nand U13775 (N_13775,N_10052,N_8406);
nand U13776 (N_13776,N_8244,N_8882);
nand U13777 (N_13777,N_10056,N_11351);
nand U13778 (N_13778,N_8531,N_11642);
nor U13779 (N_13779,N_9175,N_11209);
nor U13780 (N_13780,N_8394,N_10609);
and U13781 (N_13781,N_10048,N_11332);
or U13782 (N_13782,N_10103,N_9458);
and U13783 (N_13783,N_8211,N_11517);
and U13784 (N_13784,N_10008,N_9809);
nand U13785 (N_13785,N_8797,N_11317);
or U13786 (N_13786,N_11702,N_9907);
or U13787 (N_13787,N_9279,N_11989);
nor U13788 (N_13788,N_11845,N_10432);
nand U13789 (N_13789,N_10041,N_10625);
or U13790 (N_13790,N_11415,N_8186);
or U13791 (N_13791,N_9768,N_11407);
or U13792 (N_13792,N_11875,N_8973);
nand U13793 (N_13793,N_11634,N_11376);
nor U13794 (N_13794,N_11029,N_8672);
nand U13795 (N_13795,N_8683,N_11935);
and U13796 (N_13796,N_11291,N_8342);
nor U13797 (N_13797,N_11169,N_9456);
nand U13798 (N_13798,N_9919,N_8163);
nor U13799 (N_13799,N_9428,N_8454);
nand U13800 (N_13800,N_9313,N_9780);
nor U13801 (N_13801,N_9889,N_11807);
nor U13802 (N_13802,N_8755,N_11896);
and U13803 (N_13803,N_11163,N_10634);
nor U13804 (N_13804,N_10452,N_9520);
and U13805 (N_13805,N_8506,N_9232);
nand U13806 (N_13806,N_10339,N_11915);
and U13807 (N_13807,N_8975,N_11343);
nor U13808 (N_13808,N_9504,N_11294);
nor U13809 (N_13809,N_8972,N_10968);
nand U13810 (N_13810,N_8058,N_11545);
nor U13811 (N_13811,N_11088,N_8504);
nor U13812 (N_13812,N_8507,N_9347);
and U13813 (N_13813,N_11538,N_10356);
nand U13814 (N_13814,N_9636,N_9253);
xnor U13815 (N_13815,N_8352,N_10853);
nand U13816 (N_13816,N_9312,N_11980);
and U13817 (N_13817,N_9614,N_9155);
nor U13818 (N_13818,N_11567,N_11445);
nor U13819 (N_13819,N_11473,N_8602);
nor U13820 (N_13820,N_8967,N_11177);
or U13821 (N_13821,N_8305,N_8230);
nand U13822 (N_13822,N_9365,N_8888);
xnor U13823 (N_13823,N_8671,N_8511);
or U13824 (N_13824,N_8653,N_9282);
and U13825 (N_13825,N_8113,N_8660);
and U13826 (N_13826,N_11792,N_10945);
and U13827 (N_13827,N_8165,N_8747);
or U13828 (N_13828,N_10168,N_10491);
nor U13829 (N_13829,N_8586,N_9521);
nor U13830 (N_13830,N_8611,N_11313);
and U13831 (N_13831,N_11446,N_10504);
or U13832 (N_13832,N_10038,N_10225);
and U13833 (N_13833,N_10639,N_9913);
and U13834 (N_13834,N_9158,N_10900);
nor U13835 (N_13835,N_9187,N_10973);
or U13836 (N_13836,N_11919,N_8490);
and U13837 (N_13837,N_9472,N_8806);
nand U13838 (N_13838,N_10387,N_8285);
nor U13839 (N_13839,N_9151,N_9072);
nand U13840 (N_13840,N_8677,N_10093);
or U13841 (N_13841,N_9948,N_10263);
or U13842 (N_13842,N_8292,N_10822);
nand U13843 (N_13843,N_10035,N_10261);
and U13844 (N_13844,N_8133,N_8834);
nand U13845 (N_13845,N_10561,N_8934);
nor U13846 (N_13846,N_8983,N_11904);
nor U13847 (N_13847,N_10470,N_11942);
nand U13848 (N_13848,N_11084,N_9444);
and U13849 (N_13849,N_9608,N_8849);
and U13850 (N_13850,N_9987,N_10166);
or U13851 (N_13851,N_11482,N_9245);
nand U13852 (N_13852,N_9057,N_10734);
or U13853 (N_13853,N_8040,N_11526);
nor U13854 (N_13854,N_8830,N_8037);
nor U13855 (N_13855,N_11083,N_8316);
nand U13856 (N_13856,N_8251,N_9955);
nor U13857 (N_13857,N_10722,N_8598);
and U13858 (N_13858,N_10418,N_8795);
nor U13859 (N_13859,N_9103,N_11506);
or U13860 (N_13860,N_9845,N_8622);
nor U13861 (N_13861,N_9483,N_8296);
and U13862 (N_13862,N_10961,N_11055);
and U13863 (N_13863,N_8478,N_9492);
or U13864 (N_13864,N_11092,N_9264);
and U13865 (N_13865,N_11605,N_11762);
nand U13866 (N_13866,N_9936,N_11678);
and U13867 (N_13867,N_10422,N_8799);
xor U13868 (N_13868,N_9332,N_11800);
xnor U13869 (N_13869,N_8204,N_9967);
and U13870 (N_13870,N_8127,N_8245);
nand U13871 (N_13871,N_11426,N_11117);
nand U13872 (N_13872,N_11216,N_9459);
nor U13873 (N_13873,N_9112,N_8473);
or U13874 (N_13874,N_10175,N_9718);
and U13875 (N_13875,N_9196,N_11669);
and U13876 (N_13876,N_9178,N_8309);
nor U13877 (N_13877,N_8986,N_9192);
nor U13878 (N_13878,N_9391,N_9922);
nand U13879 (N_13879,N_8520,N_10167);
or U13880 (N_13880,N_10046,N_10815);
or U13881 (N_13881,N_8576,N_8929);
and U13882 (N_13882,N_10241,N_8820);
and U13883 (N_13883,N_9023,N_10015);
xnor U13884 (N_13884,N_9554,N_11809);
nor U13885 (N_13885,N_10044,N_11823);
nor U13886 (N_13886,N_8472,N_8748);
nor U13887 (N_13887,N_8369,N_9262);
and U13888 (N_13888,N_10921,N_11879);
nor U13889 (N_13889,N_9334,N_10444);
nand U13890 (N_13890,N_9124,N_8212);
nor U13891 (N_13891,N_10794,N_9924);
nand U13892 (N_13892,N_10806,N_10028);
or U13893 (N_13893,N_11310,N_11697);
nor U13894 (N_13894,N_10835,N_10414);
and U13895 (N_13895,N_11557,N_11015);
or U13896 (N_13896,N_11953,N_10547);
nor U13897 (N_13897,N_9474,N_9190);
nand U13898 (N_13898,N_8859,N_8419);
nor U13899 (N_13899,N_11660,N_10584);
and U13900 (N_13900,N_8496,N_11576);
nand U13901 (N_13901,N_10353,N_10341);
or U13902 (N_13902,N_10343,N_11956);
or U13903 (N_13903,N_8493,N_9783);
nand U13904 (N_13904,N_9538,N_9906);
or U13905 (N_13905,N_11437,N_8351);
nand U13906 (N_13906,N_8933,N_11458);
nand U13907 (N_13907,N_10502,N_10704);
or U13908 (N_13908,N_9451,N_11032);
and U13909 (N_13909,N_8604,N_9842);
and U13910 (N_13910,N_10354,N_10295);
or U13911 (N_13911,N_9547,N_10941);
nand U13912 (N_13912,N_9002,N_11128);
and U13913 (N_13913,N_9627,N_8950);
and U13914 (N_13914,N_8618,N_9871);
xor U13915 (N_13915,N_8774,N_10094);
and U13916 (N_13916,N_8564,N_9454);
and U13917 (N_13917,N_8966,N_8065);
nand U13918 (N_13918,N_9473,N_11616);
and U13919 (N_13919,N_9182,N_10174);
nor U13920 (N_13920,N_10004,N_10635);
or U13921 (N_13921,N_10328,N_11359);
nor U13922 (N_13922,N_10189,N_8049);
and U13923 (N_13923,N_11514,N_8356);
nor U13924 (N_13924,N_10185,N_8684);
and U13925 (N_13925,N_9700,N_8071);
and U13926 (N_13926,N_11797,N_10079);
nor U13927 (N_13927,N_9651,N_8288);
or U13928 (N_13928,N_11568,N_11173);
and U13929 (N_13929,N_11410,N_9696);
and U13930 (N_13930,N_9969,N_11192);
and U13931 (N_13931,N_8146,N_11459);
nor U13932 (N_13932,N_10256,N_9442);
or U13933 (N_13933,N_8234,N_10451);
nand U13934 (N_13934,N_10924,N_10140);
xnor U13935 (N_13935,N_11851,N_11057);
and U13936 (N_13936,N_11776,N_9592);
nor U13937 (N_13937,N_11607,N_9172);
nor U13938 (N_13938,N_10150,N_9004);
and U13939 (N_13939,N_9749,N_9100);
or U13940 (N_13940,N_10795,N_10571);
nor U13941 (N_13941,N_8469,N_11880);
or U13942 (N_13942,N_9788,N_11670);
nand U13943 (N_13943,N_10404,N_10782);
and U13944 (N_13944,N_9722,N_9974);
or U13945 (N_13945,N_11010,N_8770);
or U13946 (N_13946,N_8701,N_8790);
and U13947 (N_13947,N_9461,N_10499);
and U13948 (N_13948,N_9596,N_10685);
nor U13949 (N_13949,N_9360,N_8191);
nor U13950 (N_13950,N_8359,N_8804);
nand U13951 (N_13951,N_9191,N_11629);
nor U13952 (N_13952,N_9552,N_11479);
nor U13953 (N_13953,N_10169,N_8566);
nor U13954 (N_13954,N_9166,N_11248);
nand U13955 (N_13955,N_11096,N_10931);
and U13956 (N_13956,N_11775,N_8492);
nand U13957 (N_13957,N_10083,N_11213);
nor U13958 (N_13958,N_8110,N_8396);
nor U13959 (N_13959,N_9909,N_8835);
and U13960 (N_13960,N_8122,N_11724);
and U13961 (N_13961,N_11063,N_9315);
or U13962 (N_13962,N_9666,N_9386);
or U13963 (N_13963,N_9795,N_10892);
nand U13964 (N_13964,N_9745,N_11995);
nor U13965 (N_13965,N_10972,N_11361);
nand U13966 (N_13966,N_10301,N_11307);
nand U13967 (N_13967,N_9273,N_10237);
nor U13968 (N_13968,N_11767,N_10881);
nand U13969 (N_13969,N_9149,N_10845);
or U13970 (N_13970,N_10518,N_9664);
or U13971 (N_13971,N_9440,N_9147);
nor U13972 (N_13972,N_9619,N_10102);
and U13973 (N_13973,N_9326,N_10009);
or U13974 (N_13974,N_10146,N_8612);
nor U13975 (N_13975,N_10866,N_8145);
nor U13976 (N_13976,N_9363,N_10839);
nor U13977 (N_13977,N_8696,N_11103);
or U13978 (N_13978,N_11476,N_9756);
or U13979 (N_13979,N_11235,N_10848);
or U13980 (N_13980,N_11681,N_8074);
or U13981 (N_13981,N_11199,N_11791);
nand U13982 (N_13982,N_8536,N_9207);
nand U13983 (N_13983,N_10232,N_8741);
nand U13984 (N_13984,N_9815,N_11832);
nor U13985 (N_13985,N_8792,N_10958);
and U13986 (N_13986,N_9506,N_10666);
xnor U13987 (N_13987,N_11663,N_9840);
nand U13988 (N_13988,N_10091,N_8739);
and U13989 (N_13989,N_11949,N_9999);
nor U13990 (N_13990,N_10297,N_11685);
nand U13991 (N_13991,N_8479,N_10581);
and U13992 (N_13992,N_10510,N_11855);
or U13993 (N_13993,N_8993,N_9250);
nand U13994 (N_13994,N_10714,N_8938);
xnor U13995 (N_13995,N_11430,N_8575);
nor U13996 (N_13996,N_11788,N_10095);
nor U13997 (N_13997,N_8863,N_11350);
nand U13998 (N_13998,N_8240,N_9656);
or U13999 (N_13999,N_10534,N_8328);
or U14000 (N_14000,N_8841,N_11021);
or U14001 (N_14001,N_8222,N_8127);
or U14002 (N_14002,N_9175,N_9379);
nand U14003 (N_14003,N_10537,N_9908);
nor U14004 (N_14004,N_10046,N_10786);
or U14005 (N_14005,N_8637,N_11486);
nor U14006 (N_14006,N_8405,N_8726);
and U14007 (N_14007,N_11020,N_11409);
or U14008 (N_14008,N_9090,N_10673);
and U14009 (N_14009,N_8615,N_11499);
nand U14010 (N_14010,N_10462,N_11801);
nor U14011 (N_14011,N_11572,N_10906);
nor U14012 (N_14012,N_11270,N_8159);
xnor U14013 (N_14013,N_11424,N_10715);
nand U14014 (N_14014,N_9638,N_10148);
nand U14015 (N_14015,N_8505,N_9169);
nand U14016 (N_14016,N_11560,N_11262);
nor U14017 (N_14017,N_9179,N_10328);
and U14018 (N_14018,N_9227,N_10735);
nand U14019 (N_14019,N_9408,N_10222);
and U14020 (N_14020,N_9446,N_11462);
and U14021 (N_14021,N_10013,N_8456);
or U14022 (N_14022,N_11957,N_11068);
and U14023 (N_14023,N_11968,N_10475);
nand U14024 (N_14024,N_11835,N_8823);
and U14025 (N_14025,N_10694,N_11954);
nor U14026 (N_14026,N_10563,N_11844);
nand U14027 (N_14027,N_8622,N_8306);
nor U14028 (N_14028,N_9582,N_8625);
nand U14029 (N_14029,N_10047,N_11306);
nor U14030 (N_14030,N_9389,N_11231);
and U14031 (N_14031,N_10926,N_9074);
and U14032 (N_14032,N_11809,N_10420);
xnor U14033 (N_14033,N_9736,N_11061);
nor U14034 (N_14034,N_10508,N_8909);
nand U14035 (N_14035,N_11568,N_11976);
nor U14036 (N_14036,N_8479,N_8809);
or U14037 (N_14037,N_11063,N_11241);
and U14038 (N_14038,N_11837,N_11177);
xnor U14039 (N_14039,N_10503,N_9554);
and U14040 (N_14040,N_10458,N_9354);
nand U14041 (N_14041,N_10900,N_8209);
nand U14042 (N_14042,N_8755,N_11063);
and U14043 (N_14043,N_8709,N_11069);
nand U14044 (N_14044,N_10246,N_10214);
and U14045 (N_14045,N_9756,N_11690);
and U14046 (N_14046,N_10967,N_11255);
or U14047 (N_14047,N_9597,N_9934);
and U14048 (N_14048,N_9321,N_10183);
and U14049 (N_14049,N_8163,N_9847);
and U14050 (N_14050,N_10859,N_8929);
and U14051 (N_14051,N_8275,N_10024);
or U14052 (N_14052,N_11601,N_11187);
and U14053 (N_14053,N_11448,N_10958);
and U14054 (N_14054,N_8569,N_8035);
xor U14055 (N_14055,N_11612,N_9177);
and U14056 (N_14056,N_10908,N_11793);
nand U14057 (N_14057,N_10461,N_9691);
nand U14058 (N_14058,N_11286,N_8800);
and U14059 (N_14059,N_11698,N_11093);
and U14060 (N_14060,N_9632,N_8618);
nand U14061 (N_14061,N_11556,N_11630);
nand U14062 (N_14062,N_11711,N_9883);
or U14063 (N_14063,N_10841,N_8790);
and U14064 (N_14064,N_8846,N_10161);
nand U14065 (N_14065,N_9517,N_11940);
or U14066 (N_14066,N_8426,N_9269);
and U14067 (N_14067,N_11232,N_8097);
or U14068 (N_14068,N_11990,N_11105);
nor U14069 (N_14069,N_9134,N_11750);
nor U14070 (N_14070,N_9272,N_11522);
and U14071 (N_14071,N_11377,N_10588);
nand U14072 (N_14072,N_10194,N_9070);
nor U14073 (N_14073,N_8795,N_10995);
and U14074 (N_14074,N_11201,N_8784);
or U14075 (N_14075,N_10321,N_11119);
and U14076 (N_14076,N_10771,N_10810);
nand U14077 (N_14077,N_10181,N_10634);
and U14078 (N_14078,N_8717,N_9860);
and U14079 (N_14079,N_9012,N_11067);
nand U14080 (N_14080,N_11579,N_10396);
nor U14081 (N_14081,N_9579,N_10700);
and U14082 (N_14082,N_10435,N_8822);
nor U14083 (N_14083,N_10114,N_8755);
xnor U14084 (N_14084,N_11099,N_11078);
nand U14085 (N_14085,N_9240,N_9081);
nor U14086 (N_14086,N_8888,N_10662);
nand U14087 (N_14087,N_8651,N_11320);
nor U14088 (N_14088,N_9190,N_8223);
nor U14089 (N_14089,N_10406,N_9553);
nand U14090 (N_14090,N_10818,N_9813);
nand U14091 (N_14091,N_9200,N_11483);
nor U14092 (N_14092,N_8767,N_10394);
nand U14093 (N_14093,N_10573,N_8851);
nor U14094 (N_14094,N_11378,N_10539);
nand U14095 (N_14095,N_9167,N_10918);
or U14096 (N_14096,N_9423,N_10511);
nand U14097 (N_14097,N_8806,N_10635);
nand U14098 (N_14098,N_9180,N_10485);
nor U14099 (N_14099,N_9367,N_10890);
nor U14100 (N_14100,N_9121,N_11213);
nor U14101 (N_14101,N_11895,N_11601);
nand U14102 (N_14102,N_8235,N_10421);
and U14103 (N_14103,N_10951,N_8999);
nor U14104 (N_14104,N_10251,N_8326);
and U14105 (N_14105,N_10237,N_8606);
nor U14106 (N_14106,N_8139,N_8214);
and U14107 (N_14107,N_10080,N_8327);
and U14108 (N_14108,N_8060,N_8024);
or U14109 (N_14109,N_11523,N_10472);
and U14110 (N_14110,N_8795,N_9709);
or U14111 (N_14111,N_10653,N_11447);
and U14112 (N_14112,N_8314,N_8093);
nand U14113 (N_14113,N_11056,N_9595);
nand U14114 (N_14114,N_9182,N_10943);
nor U14115 (N_14115,N_8656,N_9483);
nand U14116 (N_14116,N_8033,N_11374);
and U14117 (N_14117,N_11062,N_11204);
and U14118 (N_14118,N_11017,N_8454);
or U14119 (N_14119,N_8585,N_8093);
xor U14120 (N_14120,N_8151,N_8428);
nor U14121 (N_14121,N_8189,N_10685);
nor U14122 (N_14122,N_11510,N_11511);
or U14123 (N_14123,N_8192,N_10371);
or U14124 (N_14124,N_9828,N_9703);
and U14125 (N_14125,N_11602,N_11474);
nor U14126 (N_14126,N_8589,N_8670);
or U14127 (N_14127,N_9174,N_11247);
or U14128 (N_14128,N_9872,N_8340);
nor U14129 (N_14129,N_9985,N_10444);
nor U14130 (N_14130,N_10152,N_10245);
nor U14131 (N_14131,N_10377,N_9086);
or U14132 (N_14132,N_8894,N_10847);
or U14133 (N_14133,N_8547,N_10242);
and U14134 (N_14134,N_8095,N_11116);
nand U14135 (N_14135,N_8207,N_9916);
and U14136 (N_14136,N_11103,N_9741);
or U14137 (N_14137,N_10439,N_10811);
and U14138 (N_14138,N_8003,N_10545);
nand U14139 (N_14139,N_11982,N_8099);
and U14140 (N_14140,N_10636,N_10106);
nand U14141 (N_14141,N_11480,N_9196);
or U14142 (N_14142,N_11422,N_8088);
or U14143 (N_14143,N_9679,N_9289);
nor U14144 (N_14144,N_9624,N_10948);
or U14145 (N_14145,N_11154,N_8741);
nand U14146 (N_14146,N_10246,N_11887);
or U14147 (N_14147,N_10635,N_9492);
or U14148 (N_14148,N_9410,N_9113);
or U14149 (N_14149,N_9699,N_10847);
nor U14150 (N_14150,N_8895,N_10204);
nand U14151 (N_14151,N_10474,N_8559);
or U14152 (N_14152,N_11823,N_8231);
nor U14153 (N_14153,N_10661,N_9266);
or U14154 (N_14154,N_11007,N_11501);
nand U14155 (N_14155,N_10813,N_9881);
nor U14156 (N_14156,N_11262,N_9582);
nor U14157 (N_14157,N_8268,N_8587);
nand U14158 (N_14158,N_8356,N_8992);
and U14159 (N_14159,N_11940,N_8003);
and U14160 (N_14160,N_10912,N_8791);
or U14161 (N_14161,N_10756,N_10393);
or U14162 (N_14162,N_10975,N_10949);
and U14163 (N_14163,N_10088,N_9166);
and U14164 (N_14164,N_9251,N_11851);
nand U14165 (N_14165,N_8605,N_9565);
nand U14166 (N_14166,N_9923,N_8385);
xnor U14167 (N_14167,N_11360,N_10083);
or U14168 (N_14168,N_10917,N_9615);
and U14169 (N_14169,N_9723,N_10002);
or U14170 (N_14170,N_11704,N_8284);
nand U14171 (N_14171,N_9182,N_8601);
nand U14172 (N_14172,N_9708,N_10634);
nand U14173 (N_14173,N_10984,N_8629);
and U14174 (N_14174,N_9466,N_10461);
nor U14175 (N_14175,N_9531,N_8526);
and U14176 (N_14176,N_11085,N_8059);
or U14177 (N_14177,N_9920,N_10366);
nor U14178 (N_14178,N_8697,N_9359);
xnor U14179 (N_14179,N_9929,N_8099);
and U14180 (N_14180,N_10376,N_8849);
and U14181 (N_14181,N_10365,N_10744);
and U14182 (N_14182,N_8440,N_9826);
and U14183 (N_14183,N_11636,N_8327);
or U14184 (N_14184,N_8190,N_10247);
and U14185 (N_14185,N_9105,N_8356);
and U14186 (N_14186,N_10744,N_11141);
nand U14187 (N_14187,N_9080,N_9787);
or U14188 (N_14188,N_10945,N_9007);
and U14189 (N_14189,N_9363,N_10285);
nor U14190 (N_14190,N_9121,N_8943);
nand U14191 (N_14191,N_9897,N_8832);
and U14192 (N_14192,N_10430,N_8198);
nor U14193 (N_14193,N_11480,N_11011);
and U14194 (N_14194,N_9632,N_10897);
and U14195 (N_14195,N_10106,N_11911);
or U14196 (N_14196,N_9137,N_11079);
nand U14197 (N_14197,N_10394,N_10886);
nor U14198 (N_14198,N_8129,N_10650);
nand U14199 (N_14199,N_9890,N_9448);
nand U14200 (N_14200,N_11680,N_9070);
or U14201 (N_14201,N_11875,N_8425);
or U14202 (N_14202,N_8566,N_8419);
nand U14203 (N_14203,N_9030,N_11111);
nand U14204 (N_14204,N_10007,N_8703);
and U14205 (N_14205,N_10330,N_9473);
nor U14206 (N_14206,N_10209,N_9557);
nor U14207 (N_14207,N_11564,N_10441);
nand U14208 (N_14208,N_10775,N_9002);
nor U14209 (N_14209,N_10988,N_10727);
and U14210 (N_14210,N_9233,N_9462);
nand U14211 (N_14211,N_10348,N_11060);
nor U14212 (N_14212,N_8669,N_10157);
or U14213 (N_14213,N_8690,N_9214);
or U14214 (N_14214,N_9976,N_8149);
and U14215 (N_14215,N_9391,N_11866);
nor U14216 (N_14216,N_9454,N_10435);
nor U14217 (N_14217,N_10923,N_10668);
and U14218 (N_14218,N_8712,N_8505);
nor U14219 (N_14219,N_8858,N_8183);
nand U14220 (N_14220,N_10291,N_9212);
or U14221 (N_14221,N_11635,N_11887);
and U14222 (N_14222,N_8012,N_11955);
nor U14223 (N_14223,N_8823,N_11574);
or U14224 (N_14224,N_9085,N_8560);
nand U14225 (N_14225,N_8512,N_9572);
nand U14226 (N_14226,N_8878,N_10506);
and U14227 (N_14227,N_9073,N_8182);
and U14228 (N_14228,N_8966,N_8013);
and U14229 (N_14229,N_11092,N_8743);
and U14230 (N_14230,N_8539,N_10628);
nand U14231 (N_14231,N_11327,N_10895);
and U14232 (N_14232,N_8098,N_10998);
nand U14233 (N_14233,N_9640,N_10447);
or U14234 (N_14234,N_9914,N_9863);
or U14235 (N_14235,N_9639,N_11099);
nor U14236 (N_14236,N_8925,N_8242);
nand U14237 (N_14237,N_9771,N_10944);
or U14238 (N_14238,N_8398,N_8307);
xnor U14239 (N_14239,N_9767,N_10588);
xnor U14240 (N_14240,N_8002,N_9868);
or U14241 (N_14241,N_10134,N_11158);
or U14242 (N_14242,N_9783,N_11850);
nor U14243 (N_14243,N_11219,N_8969);
and U14244 (N_14244,N_10626,N_11706);
nor U14245 (N_14245,N_10687,N_10560);
or U14246 (N_14246,N_8149,N_11222);
nand U14247 (N_14247,N_10090,N_9161);
nor U14248 (N_14248,N_11895,N_11725);
nor U14249 (N_14249,N_9788,N_8284);
or U14250 (N_14250,N_9630,N_10082);
nor U14251 (N_14251,N_11625,N_9946);
nand U14252 (N_14252,N_9771,N_10169);
nand U14253 (N_14253,N_10242,N_11297);
nor U14254 (N_14254,N_8288,N_11201);
nand U14255 (N_14255,N_10440,N_9734);
nor U14256 (N_14256,N_9376,N_11804);
and U14257 (N_14257,N_11204,N_9954);
nor U14258 (N_14258,N_11275,N_9627);
nand U14259 (N_14259,N_11339,N_11413);
or U14260 (N_14260,N_10806,N_9547);
nor U14261 (N_14261,N_11381,N_11312);
nand U14262 (N_14262,N_10569,N_11343);
nor U14263 (N_14263,N_8111,N_11174);
nor U14264 (N_14264,N_10291,N_8477);
and U14265 (N_14265,N_8358,N_10328);
or U14266 (N_14266,N_10687,N_11728);
or U14267 (N_14267,N_11516,N_9735);
nor U14268 (N_14268,N_10707,N_9133);
nor U14269 (N_14269,N_10243,N_9320);
or U14270 (N_14270,N_8948,N_8872);
and U14271 (N_14271,N_8132,N_11534);
or U14272 (N_14272,N_10277,N_8637);
or U14273 (N_14273,N_11113,N_9189);
and U14274 (N_14274,N_9574,N_8912);
nor U14275 (N_14275,N_10689,N_9527);
xnor U14276 (N_14276,N_10154,N_10935);
nand U14277 (N_14277,N_9240,N_8780);
and U14278 (N_14278,N_10664,N_11364);
nand U14279 (N_14279,N_10827,N_10217);
nand U14280 (N_14280,N_9173,N_11602);
or U14281 (N_14281,N_10410,N_11962);
and U14282 (N_14282,N_11160,N_10142);
and U14283 (N_14283,N_8391,N_8947);
and U14284 (N_14284,N_10686,N_8591);
nand U14285 (N_14285,N_8990,N_8431);
and U14286 (N_14286,N_10210,N_9773);
and U14287 (N_14287,N_9110,N_11716);
nand U14288 (N_14288,N_8353,N_8455);
nor U14289 (N_14289,N_10240,N_8695);
or U14290 (N_14290,N_9439,N_11723);
xor U14291 (N_14291,N_11776,N_9522);
and U14292 (N_14292,N_11778,N_9589);
nor U14293 (N_14293,N_8948,N_9828);
nand U14294 (N_14294,N_10821,N_8080);
nor U14295 (N_14295,N_11466,N_9402);
or U14296 (N_14296,N_9187,N_9481);
and U14297 (N_14297,N_9379,N_11598);
or U14298 (N_14298,N_8466,N_9521);
or U14299 (N_14299,N_8323,N_8358);
nor U14300 (N_14300,N_8614,N_8149);
nand U14301 (N_14301,N_10258,N_8290);
nor U14302 (N_14302,N_10875,N_8396);
or U14303 (N_14303,N_11085,N_10895);
nor U14304 (N_14304,N_10364,N_9591);
nor U14305 (N_14305,N_8481,N_9238);
or U14306 (N_14306,N_8881,N_11747);
or U14307 (N_14307,N_8383,N_11158);
nor U14308 (N_14308,N_8066,N_8421);
and U14309 (N_14309,N_8767,N_10784);
and U14310 (N_14310,N_10108,N_11008);
nand U14311 (N_14311,N_8921,N_9016);
and U14312 (N_14312,N_8061,N_10446);
or U14313 (N_14313,N_11613,N_9131);
or U14314 (N_14314,N_8729,N_9116);
nand U14315 (N_14315,N_9847,N_11826);
and U14316 (N_14316,N_11992,N_11396);
nand U14317 (N_14317,N_9934,N_10725);
nand U14318 (N_14318,N_10642,N_10262);
nor U14319 (N_14319,N_10254,N_11778);
and U14320 (N_14320,N_9171,N_10440);
nand U14321 (N_14321,N_8736,N_9277);
nand U14322 (N_14322,N_10768,N_11757);
and U14323 (N_14323,N_8139,N_11986);
and U14324 (N_14324,N_9586,N_10403);
nor U14325 (N_14325,N_8221,N_11162);
nor U14326 (N_14326,N_11062,N_10463);
and U14327 (N_14327,N_11009,N_10623);
nand U14328 (N_14328,N_10291,N_9588);
or U14329 (N_14329,N_9089,N_10745);
nor U14330 (N_14330,N_8105,N_10239);
and U14331 (N_14331,N_8151,N_8450);
and U14332 (N_14332,N_9597,N_10862);
or U14333 (N_14333,N_8352,N_8448);
or U14334 (N_14334,N_8322,N_11570);
and U14335 (N_14335,N_8031,N_11114);
xor U14336 (N_14336,N_11966,N_11991);
xor U14337 (N_14337,N_11919,N_10134);
nand U14338 (N_14338,N_10040,N_9294);
or U14339 (N_14339,N_11538,N_11429);
nand U14340 (N_14340,N_10523,N_8748);
nor U14341 (N_14341,N_8294,N_9958);
or U14342 (N_14342,N_11731,N_8867);
nand U14343 (N_14343,N_10642,N_9211);
and U14344 (N_14344,N_10855,N_10901);
or U14345 (N_14345,N_11549,N_11039);
nand U14346 (N_14346,N_8529,N_9461);
nand U14347 (N_14347,N_9144,N_8587);
or U14348 (N_14348,N_9200,N_9261);
or U14349 (N_14349,N_11917,N_8591);
nor U14350 (N_14350,N_8482,N_8611);
or U14351 (N_14351,N_10504,N_11043);
xor U14352 (N_14352,N_11066,N_9263);
nor U14353 (N_14353,N_11215,N_10988);
nor U14354 (N_14354,N_9994,N_8858);
nand U14355 (N_14355,N_8459,N_10165);
and U14356 (N_14356,N_10844,N_10267);
nand U14357 (N_14357,N_8840,N_8234);
xnor U14358 (N_14358,N_8210,N_8029);
nand U14359 (N_14359,N_11488,N_10197);
nand U14360 (N_14360,N_11057,N_9809);
nand U14361 (N_14361,N_8107,N_9664);
nor U14362 (N_14362,N_11950,N_8432);
xor U14363 (N_14363,N_10836,N_11577);
or U14364 (N_14364,N_11856,N_8936);
and U14365 (N_14365,N_11045,N_9950);
and U14366 (N_14366,N_11144,N_9733);
or U14367 (N_14367,N_8485,N_9437);
nand U14368 (N_14368,N_9777,N_9175);
and U14369 (N_14369,N_8562,N_8863);
nand U14370 (N_14370,N_11220,N_11851);
or U14371 (N_14371,N_10949,N_9772);
nor U14372 (N_14372,N_8557,N_8749);
or U14373 (N_14373,N_9191,N_11819);
and U14374 (N_14374,N_11398,N_9744);
nand U14375 (N_14375,N_9241,N_10839);
nor U14376 (N_14376,N_10883,N_10270);
and U14377 (N_14377,N_9531,N_9572);
xor U14378 (N_14378,N_11137,N_11858);
nand U14379 (N_14379,N_9921,N_10320);
nand U14380 (N_14380,N_11319,N_11820);
and U14381 (N_14381,N_8567,N_8661);
and U14382 (N_14382,N_10867,N_11557);
nand U14383 (N_14383,N_11541,N_9466);
nor U14384 (N_14384,N_10581,N_10794);
nand U14385 (N_14385,N_9030,N_9438);
and U14386 (N_14386,N_8676,N_10648);
nor U14387 (N_14387,N_9629,N_11671);
nor U14388 (N_14388,N_10739,N_11150);
nand U14389 (N_14389,N_10995,N_10717);
nor U14390 (N_14390,N_8434,N_9144);
nor U14391 (N_14391,N_9089,N_9828);
nor U14392 (N_14392,N_10967,N_11825);
and U14393 (N_14393,N_9874,N_9306);
and U14394 (N_14394,N_10657,N_9215);
nand U14395 (N_14395,N_11709,N_9114);
and U14396 (N_14396,N_10943,N_11401);
nand U14397 (N_14397,N_11768,N_11456);
nor U14398 (N_14398,N_11072,N_10421);
xnor U14399 (N_14399,N_10804,N_11878);
nand U14400 (N_14400,N_11275,N_8001);
nand U14401 (N_14401,N_9649,N_8618);
or U14402 (N_14402,N_9474,N_9321);
nor U14403 (N_14403,N_9247,N_11522);
nand U14404 (N_14404,N_9888,N_9898);
and U14405 (N_14405,N_10130,N_9334);
or U14406 (N_14406,N_10722,N_8824);
nor U14407 (N_14407,N_10517,N_8978);
nand U14408 (N_14408,N_9391,N_11138);
and U14409 (N_14409,N_10513,N_10885);
nand U14410 (N_14410,N_9510,N_8931);
or U14411 (N_14411,N_9193,N_11330);
nor U14412 (N_14412,N_10474,N_9134);
or U14413 (N_14413,N_10881,N_10238);
nor U14414 (N_14414,N_10281,N_11682);
and U14415 (N_14415,N_9539,N_10412);
and U14416 (N_14416,N_8338,N_11434);
nand U14417 (N_14417,N_9500,N_8219);
nor U14418 (N_14418,N_8131,N_10967);
nor U14419 (N_14419,N_8097,N_9032);
nor U14420 (N_14420,N_10776,N_8798);
or U14421 (N_14421,N_10916,N_10872);
or U14422 (N_14422,N_11972,N_11389);
or U14423 (N_14423,N_9480,N_8737);
and U14424 (N_14424,N_11000,N_9785);
nand U14425 (N_14425,N_10346,N_9905);
nor U14426 (N_14426,N_11862,N_9627);
and U14427 (N_14427,N_9346,N_11959);
or U14428 (N_14428,N_9488,N_10337);
nand U14429 (N_14429,N_10891,N_9439);
and U14430 (N_14430,N_11586,N_9236);
nand U14431 (N_14431,N_10007,N_10216);
and U14432 (N_14432,N_9411,N_9044);
nor U14433 (N_14433,N_9270,N_8633);
or U14434 (N_14434,N_9012,N_9534);
nand U14435 (N_14435,N_8421,N_8216);
and U14436 (N_14436,N_10953,N_9158);
or U14437 (N_14437,N_9576,N_11585);
or U14438 (N_14438,N_8802,N_9802);
xnor U14439 (N_14439,N_10552,N_8837);
nor U14440 (N_14440,N_10922,N_10124);
and U14441 (N_14441,N_8234,N_8089);
nand U14442 (N_14442,N_11354,N_10948);
and U14443 (N_14443,N_9464,N_10896);
and U14444 (N_14444,N_9511,N_8570);
and U14445 (N_14445,N_9605,N_9077);
and U14446 (N_14446,N_9226,N_11411);
nand U14447 (N_14447,N_11778,N_10962);
xnor U14448 (N_14448,N_11645,N_10322);
nand U14449 (N_14449,N_8597,N_8563);
nor U14450 (N_14450,N_11065,N_9616);
nand U14451 (N_14451,N_8523,N_11385);
or U14452 (N_14452,N_10751,N_11015);
nor U14453 (N_14453,N_8593,N_10432);
or U14454 (N_14454,N_8029,N_11485);
nand U14455 (N_14455,N_11074,N_8337);
nand U14456 (N_14456,N_10835,N_9266);
nor U14457 (N_14457,N_10820,N_10730);
nand U14458 (N_14458,N_9551,N_9351);
nor U14459 (N_14459,N_10499,N_8762);
and U14460 (N_14460,N_10050,N_11520);
or U14461 (N_14461,N_9291,N_11812);
nand U14462 (N_14462,N_9406,N_8770);
nor U14463 (N_14463,N_9142,N_9159);
and U14464 (N_14464,N_9763,N_9559);
nand U14465 (N_14465,N_11533,N_9332);
nand U14466 (N_14466,N_11475,N_11657);
nor U14467 (N_14467,N_8873,N_10553);
nor U14468 (N_14468,N_9609,N_9953);
or U14469 (N_14469,N_11607,N_8512);
and U14470 (N_14470,N_11254,N_9770);
or U14471 (N_14471,N_8225,N_11118);
or U14472 (N_14472,N_9687,N_8326);
and U14473 (N_14473,N_9193,N_10201);
and U14474 (N_14474,N_11662,N_9771);
nand U14475 (N_14475,N_10711,N_9725);
and U14476 (N_14476,N_11816,N_8131);
and U14477 (N_14477,N_8913,N_10017);
nand U14478 (N_14478,N_10302,N_11284);
nand U14479 (N_14479,N_9252,N_11409);
nor U14480 (N_14480,N_9534,N_9860);
or U14481 (N_14481,N_10556,N_8904);
or U14482 (N_14482,N_9035,N_9307);
nor U14483 (N_14483,N_8360,N_11067);
nor U14484 (N_14484,N_10575,N_8076);
nand U14485 (N_14485,N_8027,N_11535);
and U14486 (N_14486,N_9974,N_10383);
and U14487 (N_14487,N_9444,N_10648);
and U14488 (N_14488,N_11141,N_10290);
and U14489 (N_14489,N_9475,N_9221);
nand U14490 (N_14490,N_8998,N_9978);
and U14491 (N_14491,N_10269,N_8440);
or U14492 (N_14492,N_9526,N_11094);
nand U14493 (N_14493,N_8116,N_10450);
nor U14494 (N_14494,N_10998,N_8432);
xor U14495 (N_14495,N_8894,N_10200);
nand U14496 (N_14496,N_8105,N_9953);
or U14497 (N_14497,N_9315,N_10752);
nor U14498 (N_14498,N_10099,N_8024);
and U14499 (N_14499,N_11970,N_9493);
and U14500 (N_14500,N_11518,N_9762);
nand U14501 (N_14501,N_10308,N_9346);
nor U14502 (N_14502,N_11540,N_9370);
nand U14503 (N_14503,N_11464,N_11610);
nand U14504 (N_14504,N_10891,N_8702);
nor U14505 (N_14505,N_9680,N_9899);
nand U14506 (N_14506,N_9084,N_10731);
xor U14507 (N_14507,N_11017,N_8599);
and U14508 (N_14508,N_11656,N_10146);
and U14509 (N_14509,N_11746,N_11041);
nor U14510 (N_14510,N_9891,N_9699);
and U14511 (N_14511,N_9174,N_10337);
and U14512 (N_14512,N_9464,N_8328);
or U14513 (N_14513,N_11623,N_11949);
or U14514 (N_14514,N_10604,N_8609);
or U14515 (N_14515,N_10197,N_8816);
nand U14516 (N_14516,N_9099,N_11299);
and U14517 (N_14517,N_8966,N_9540);
and U14518 (N_14518,N_8455,N_10701);
and U14519 (N_14519,N_10777,N_11558);
nor U14520 (N_14520,N_9006,N_11190);
and U14521 (N_14521,N_10938,N_9794);
and U14522 (N_14522,N_11176,N_11649);
or U14523 (N_14523,N_11692,N_8444);
nor U14524 (N_14524,N_8215,N_8171);
nand U14525 (N_14525,N_11821,N_8187);
and U14526 (N_14526,N_8243,N_11549);
xnor U14527 (N_14527,N_11921,N_8483);
nor U14528 (N_14528,N_9032,N_11733);
and U14529 (N_14529,N_10142,N_10914);
xnor U14530 (N_14530,N_11044,N_9300);
nand U14531 (N_14531,N_8606,N_11862);
and U14532 (N_14532,N_11981,N_10342);
and U14533 (N_14533,N_8435,N_11727);
or U14534 (N_14534,N_10238,N_11305);
and U14535 (N_14535,N_9863,N_8996);
or U14536 (N_14536,N_10606,N_9077);
and U14537 (N_14537,N_10760,N_8380);
or U14538 (N_14538,N_10979,N_9372);
and U14539 (N_14539,N_8873,N_11964);
nand U14540 (N_14540,N_9790,N_11459);
nand U14541 (N_14541,N_8087,N_9541);
nand U14542 (N_14542,N_8171,N_8948);
and U14543 (N_14543,N_9634,N_11137);
nor U14544 (N_14544,N_8965,N_9740);
or U14545 (N_14545,N_8905,N_8795);
or U14546 (N_14546,N_9950,N_10784);
and U14547 (N_14547,N_9444,N_9877);
nor U14548 (N_14548,N_10707,N_8688);
nor U14549 (N_14549,N_11965,N_9389);
and U14550 (N_14550,N_8725,N_9361);
and U14551 (N_14551,N_10700,N_8117);
or U14552 (N_14552,N_10468,N_9936);
nor U14553 (N_14553,N_8046,N_11746);
nor U14554 (N_14554,N_9876,N_9480);
and U14555 (N_14555,N_9150,N_11930);
nand U14556 (N_14556,N_11857,N_9387);
nand U14557 (N_14557,N_8995,N_10738);
and U14558 (N_14558,N_9756,N_10522);
and U14559 (N_14559,N_9567,N_9138);
or U14560 (N_14560,N_9054,N_9377);
and U14561 (N_14561,N_11599,N_11927);
and U14562 (N_14562,N_11462,N_11931);
and U14563 (N_14563,N_11139,N_11196);
nand U14564 (N_14564,N_10726,N_9559);
and U14565 (N_14565,N_8564,N_9643);
or U14566 (N_14566,N_10371,N_11872);
nand U14567 (N_14567,N_9247,N_8965);
and U14568 (N_14568,N_8357,N_11672);
xnor U14569 (N_14569,N_10843,N_9538);
nor U14570 (N_14570,N_10501,N_9880);
nor U14571 (N_14571,N_9921,N_9171);
nand U14572 (N_14572,N_10815,N_10254);
nor U14573 (N_14573,N_10366,N_10491);
or U14574 (N_14574,N_8923,N_8216);
nor U14575 (N_14575,N_10464,N_9125);
nand U14576 (N_14576,N_8964,N_8278);
nand U14577 (N_14577,N_8543,N_9657);
and U14578 (N_14578,N_9281,N_8937);
and U14579 (N_14579,N_9935,N_11831);
and U14580 (N_14580,N_8275,N_9136);
nand U14581 (N_14581,N_9984,N_8866);
nor U14582 (N_14582,N_9021,N_10672);
and U14583 (N_14583,N_9054,N_11576);
and U14584 (N_14584,N_8078,N_11794);
or U14585 (N_14585,N_11827,N_10400);
xnor U14586 (N_14586,N_8957,N_10093);
and U14587 (N_14587,N_11653,N_8124);
nor U14588 (N_14588,N_8613,N_10546);
nor U14589 (N_14589,N_11057,N_8004);
or U14590 (N_14590,N_10197,N_10892);
or U14591 (N_14591,N_8170,N_9331);
nand U14592 (N_14592,N_11851,N_10141);
and U14593 (N_14593,N_10356,N_9406);
nor U14594 (N_14594,N_11255,N_11389);
nor U14595 (N_14595,N_8813,N_11620);
and U14596 (N_14596,N_11997,N_11429);
or U14597 (N_14597,N_11887,N_9218);
nand U14598 (N_14598,N_11717,N_11092);
and U14599 (N_14599,N_10774,N_9975);
nand U14600 (N_14600,N_9162,N_8348);
nor U14601 (N_14601,N_11354,N_10705);
and U14602 (N_14602,N_10015,N_10189);
or U14603 (N_14603,N_9447,N_11602);
or U14604 (N_14604,N_10506,N_9953);
nor U14605 (N_14605,N_8470,N_11910);
nor U14606 (N_14606,N_9580,N_11872);
nand U14607 (N_14607,N_10966,N_11724);
and U14608 (N_14608,N_11901,N_9116);
and U14609 (N_14609,N_10946,N_11722);
and U14610 (N_14610,N_11257,N_11304);
and U14611 (N_14611,N_9018,N_8163);
nor U14612 (N_14612,N_10077,N_8232);
or U14613 (N_14613,N_8424,N_8298);
or U14614 (N_14614,N_11825,N_10879);
and U14615 (N_14615,N_11077,N_11711);
or U14616 (N_14616,N_8882,N_9312);
or U14617 (N_14617,N_9084,N_11113);
and U14618 (N_14618,N_10600,N_8037);
and U14619 (N_14619,N_8727,N_10110);
or U14620 (N_14620,N_11617,N_8263);
nand U14621 (N_14621,N_10007,N_9351);
and U14622 (N_14622,N_11350,N_9274);
or U14623 (N_14623,N_9468,N_8984);
and U14624 (N_14624,N_8202,N_10837);
or U14625 (N_14625,N_8829,N_8782);
xnor U14626 (N_14626,N_11679,N_8292);
or U14627 (N_14627,N_9001,N_9247);
nand U14628 (N_14628,N_10152,N_11580);
xnor U14629 (N_14629,N_10641,N_9402);
nor U14630 (N_14630,N_11707,N_10933);
xor U14631 (N_14631,N_9176,N_11065);
nor U14632 (N_14632,N_8930,N_11893);
or U14633 (N_14633,N_10216,N_11994);
and U14634 (N_14634,N_10308,N_11099);
nand U14635 (N_14635,N_8126,N_10055);
or U14636 (N_14636,N_10917,N_8065);
and U14637 (N_14637,N_10158,N_10732);
nand U14638 (N_14638,N_8720,N_9181);
nand U14639 (N_14639,N_8670,N_11376);
nor U14640 (N_14640,N_10198,N_10911);
nor U14641 (N_14641,N_10629,N_9440);
nor U14642 (N_14642,N_9227,N_9070);
and U14643 (N_14643,N_9651,N_9303);
nor U14644 (N_14644,N_10127,N_9511);
and U14645 (N_14645,N_9197,N_9023);
or U14646 (N_14646,N_10021,N_9954);
nor U14647 (N_14647,N_8289,N_9306);
nand U14648 (N_14648,N_9300,N_10892);
nand U14649 (N_14649,N_10154,N_8090);
nor U14650 (N_14650,N_10399,N_10908);
and U14651 (N_14651,N_11759,N_11550);
nand U14652 (N_14652,N_10549,N_8142);
nand U14653 (N_14653,N_11110,N_10444);
nor U14654 (N_14654,N_11121,N_10509);
nand U14655 (N_14655,N_11050,N_11556);
and U14656 (N_14656,N_8977,N_9496);
nand U14657 (N_14657,N_10028,N_8836);
or U14658 (N_14658,N_8648,N_10371);
nor U14659 (N_14659,N_11519,N_8080);
nor U14660 (N_14660,N_9414,N_10062);
nor U14661 (N_14661,N_11006,N_9433);
nand U14662 (N_14662,N_11994,N_8382);
or U14663 (N_14663,N_11735,N_9155);
and U14664 (N_14664,N_8507,N_9555);
nand U14665 (N_14665,N_8299,N_10739);
nor U14666 (N_14666,N_10867,N_8760);
and U14667 (N_14667,N_11388,N_10457);
or U14668 (N_14668,N_8931,N_10905);
and U14669 (N_14669,N_9383,N_11196);
nand U14670 (N_14670,N_10660,N_10544);
and U14671 (N_14671,N_10091,N_10235);
nor U14672 (N_14672,N_9372,N_9736);
nand U14673 (N_14673,N_11101,N_8736);
and U14674 (N_14674,N_9731,N_10835);
nor U14675 (N_14675,N_9746,N_9695);
and U14676 (N_14676,N_8990,N_10069);
nand U14677 (N_14677,N_11959,N_11786);
nor U14678 (N_14678,N_8643,N_11564);
and U14679 (N_14679,N_10335,N_10003);
nand U14680 (N_14680,N_8888,N_8211);
nand U14681 (N_14681,N_10826,N_8346);
or U14682 (N_14682,N_11672,N_9648);
nor U14683 (N_14683,N_8613,N_8099);
and U14684 (N_14684,N_11374,N_10429);
and U14685 (N_14685,N_11173,N_10413);
and U14686 (N_14686,N_9138,N_11670);
xor U14687 (N_14687,N_9695,N_8953);
and U14688 (N_14688,N_10088,N_9802);
and U14689 (N_14689,N_11565,N_10609);
nand U14690 (N_14690,N_8445,N_11151);
nor U14691 (N_14691,N_11681,N_8820);
and U14692 (N_14692,N_8362,N_8349);
nor U14693 (N_14693,N_11647,N_11654);
nand U14694 (N_14694,N_10697,N_8392);
and U14695 (N_14695,N_11209,N_11808);
or U14696 (N_14696,N_8661,N_9170);
and U14697 (N_14697,N_11954,N_11978);
and U14698 (N_14698,N_10739,N_9583);
and U14699 (N_14699,N_10148,N_8894);
nand U14700 (N_14700,N_11021,N_8215);
or U14701 (N_14701,N_8576,N_8909);
nor U14702 (N_14702,N_9372,N_10945);
or U14703 (N_14703,N_8888,N_8760);
or U14704 (N_14704,N_10150,N_8863);
and U14705 (N_14705,N_11180,N_11142);
and U14706 (N_14706,N_9493,N_9258);
nand U14707 (N_14707,N_9042,N_10322);
nor U14708 (N_14708,N_9639,N_10387);
or U14709 (N_14709,N_10842,N_10027);
and U14710 (N_14710,N_10559,N_9326);
and U14711 (N_14711,N_11412,N_9831);
nor U14712 (N_14712,N_9977,N_10592);
nor U14713 (N_14713,N_10963,N_8112);
nor U14714 (N_14714,N_10387,N_11274);
or U14715 (N_14715,N_10989,N_8631);
or U14716 (N_14716,N_11766,N_10498);
and U14717 (N_14717,N_11728,N_8608);
or U14718 (N_14718,N_10434,N_11575);
nor U14719 (N_14719,N_9535,N_10596);
or U14720 (N_14720,N_11063,N_10526);
or U14721 (N_14721,N_11241,N_10907);
or U14722 (N_14722,N_10477,N_8520);
nor U14723 (N_14723,N_8226,N_11444);
nor U14724 (N_14724,N_8243,N_8622);
nand U14725 (N_14725,N_8148,N_8517);
and U14726 (N_14726,N_8045,N_9774);
nor U14727 (N_14727,N_10596,N_9837);
or U14728 (N_14728,N_11110,N_9724);
nor U14729 (N_14729,N_11403,N_9816);
nand U14730 (N_14730,N_8625,N_11602);
or U14731 (N_14731,N_10047,N_9076);
nand U14732 (N_14732,N_10662,N_11326);
and U14733 (N_14733,N_10967,N_10728);
or U14734 (N_14734,N_9904,N_10107);
or U14735 (N_14735,N_8685,N_11157);
nor U14736 (N_14736,N_9896,N_10102);
nand U14737 (N_14737,N_9076,N_10883);
nor U14738 (N_14738,N_8134,N_10031);
or U14739 (N_14739,N_10320,N_8070);
nor U14740 (N_14740,N_9302,N_11581);
nand U14741 (N_14741,N_10429,N_9928);
nor U14742 (N_14742,N_10508,N_9579);
and U14743 (N_14743,N_9561,N_9889);
or U14744 (N_14744,N_9156,N_10431);
or U14745 (N_14745,N_9907,N_8154);
nand U14746 (N_14746,N_8388,N_8920);
nand U14747 (N_14747,N_10282,N_8623);
or U14748 (N_14748,N_9307,N_11544);
nand U14749 (N_14749,N_8627,N_8905);
nand U14750 (N_14750,N_8144,N_8231);
and U14751 (N_14751,N_8905,N_11511);
nor U14752 (N_14752,N_8917,N_10230);
and U14753 (N_14753,N_10857,N_11057);
and U14754 (N_14754,N_10709,N_8309);
nor U14755 (N_14755,N_11506,N_9830);
nor U14756 (N_14756,N_9747,N_11342);
nor U14757 (N_14757,N_9788,N_8464);
or U14758 (N_14758,N_8194,N_10332);
nand U14759 (N_14759,N_11293,N_11621);
nor U14760 (N_14760,N_11745,N_11773);
and U14761 (N_14761,N_9233,N_11922);
nand U14762 (N_14762,N_11817,N_8987);
nor U14763 (N_14763,N_9829,N_10057);
and U14764 (N_14764,N_10802,N_11365);
or U14765 (N_14765,N_11724,N_9367);
nand U14766 (N_14766,N_9155,N_10083);
nand U14767 (N_14767,N_11300,N_10817);
nand U14768 (N_14768,N_11663,N_9164);
and U14769 (N_14769,N_9322,N_9859);
or U14770 (N_14770,N_11769,N_8636);
nand U14771 (N_14771,N_9624,N_9978);
or U14772 (N_14772,N_10257,N_9628);
nor U14773 (N_14773,N_8823,N_11691);
nand U14774 (N_14774,N_11546,N_11371);
or U14775 (N_14775,N_9996,N_9959);
and U14776 (N_14776,N_11408,N_11933);
nor U14777 (N_14777,N_9664,N_9683);
and U14778 (N_14778,N_9490,N_10569);
and U14779 (N_14779,N_10386,N_10008);
nand U14780 (N_14780,N_8570,N_10757);
or U14781 (N_14781,N_10152,N_10724);
nand U14782 (N_14782,N_8822,N_10812);
and U14783 (N_14783,N_11110,N_9231);
nor U14784 (N_14784,N_8940,N_9896);
and U14785 (N_14785,N_10413,N_8179);
and U14786 (N_14786,N_8621,N_9566);
and U14787 (N_14787,N_10375,N_11561);
and U14788 (N_14788,N_8009,N_9771);
and U14789 (N_14789,N_10339,N_11731);
or U14790 (N_14790,N_9275,N_11393);
and U14791 (N_14791,N_10800,N_8859);
nand U14792 (N_14792,N_9463,N_8810);
nand U14793 (N_14793,N_9147,N_8429);
nand U14794 (N_14794,N_8705,N_10878);
nor U14795 (N_14795,N_10753,N_8062);
nor U14796 (N_14796,N_10666,N_9328);
and U14797 (N_14797,N_10648,N_11621);
nor U14798 (N_14798,N_11573,N_10757);
or U14799 (N_14799,N_9298,N_8492);
and U14800 (N_14800,N_8995,N_9255);
nand U14801 (N_14801,N_11575,N_8507);
or U14802 (N_14802,N_10826,N_11778);
or U14803 (N_14803,N_11027,N_9783);
nand U14804 (N_14804,N_8819,N_10088);
nor U14805 (N_14805,N_10784,N_11965);
nand U14806 (N_14806,N_9884,N_10389);
nand U14807 (N_14807,N_9769,N_10308);
and U14808 (N_14808,N_8127,N_9996);
nor U14809 (N_14809,N_11189,N_11293);
xnor U14810 (N_14810,N_9278,N_8099);
nand U14811 (N_14811,N_9553,N_11044);
nor U14812 (N_14812,N_8336,N_10581);
or U14813 (N_14813,N_8972,N_9717);
nand U14814 (N_14814,N_10490,N_8182);
nand U14815 (N_14815,N_10796,N_10008);
nand U14816 (N_14816,N_11222,N_10693);
and U14817 (N_14817,N_9517,N_8460);
nand U14818 (N_14818,N_9751,N_9007);
nor U14819 (N_14819,N_9300,N_10827);
and U14820 (N_14820,N_11460,N_8485);
xnor U14821 (N_14821,N_8256,N_11506);
nand U14822 (N_14822,N_10829,N_8491);
nand U14823 (N_14823,N_11661,N_11696);
or U14824 (N_14824,N_8226,N_11700);
nand U14825 (N_14825,N_9475,N_11906);
nor U14826 (N_14826,N_9617,N_11071);
and U14827 (N_14827,N_8859,N_8442);
or U14828 (N_14828,N_9884,N_10113);
and U14829 (N_14829,N_11745,N_9253);
and U14830 (N_14830,N_9148,N_9636);
or U14831 (N_14831,N_10092,N_9702);
or U14832 (N_14832,N_9874,N_10067);
or U14833 (N_14833,N_10442,N_9682);
nand U14834 (N_14834,N_10249,N_8451);
nor U14835 (N_14835,N_8985,N_8293);
nand U14836 (N_14836,N_10152,N_11694);
and U14837 (N_14837,N_11630,N_11651);
nand U14838 (N_14838,N_8516,N_11375);
nand U14839 (N_14839,N_8553,N_8569);
and U14840 (N_14840,N_8429,N_8737);
nor U14841 (N_14841,N_9614,N_9145);
nand U14842 (N_14842,N_8702,N_9046);
nand U14843 (N_14843,N_9701,N_10487);
nand U14844 (N_14844,N_11053,N_9586);
and U14845 (N_14845,N_11619,N_8392);
nor U14846 (N_14846,N_11077,N_8041);
nor U14847 (N_14847,N_10152,N_10710);
and U14848 (N_14848,N_8445,N_8808);
nand U14849 (N_14849,N_10668,N_11037);
nand U14850 (N_14850,N_11866,N_8658);
nand U14851 (N_14851,N_11136,N_8926);
nor U14852 (N_14852,N_8465,N_8440);
or U14853 (N_14853,N_8557,N_9904);
and U14854 (N_14854,N_9832,N_10038);
and U14855 (N_14855,N_9376,N_11205);
or U14856 (N_14856,N_9169,N_11092);
nand U14857 (N_14857,N_8459,N_8892);
or U14858 (N_14858,N_9609,N_10506);
nor U14859 (N_14859,N_10971,N_11701);
nand U14860 (N_14860,N_10371,N_11318);
and U14861 (N_14861,N_8523,N_11961);
or U14862 (N_14862,N_9823,N_10423);
nand U14863 (N_14863,N_9773,N_11419);
xnor U14864 (N_14864,N_9668,N_10326);
and U14865 (N_14865,N_8077,N_8375);
xor U14866 (N_14866,N_9924,N_9635);
or U14867 (N_14867,N_9302,N_11842);
nor U14868 (N_14868,N_10168,N_11870);
or U14869 (N_14869,N_10963,N_10937);
and U14870 (N_14870,N_11874,N_8893);
nor U14871 (N_14871,N_9159,N_11971);
or U14872 (N_14872,N_10636,N_9086);
or U14873 (N_14873,N_11290,N_10814);
and U14874 (N_14874,N_8921,N_8027);
or U14875 (N_14875,N_11920,N_8682);
or U14876 (N_14876,N_11676,N_8187);
or U14877 (N_14877,N_10986,N_9129);
nor U14878 (N_14878,N_11122,N_8948);
or U14879 (N_14879,N_11270,N_8013);
nand U14880 (N_14880,N_11165,N_8686);
and U14881 (N_14881,N_9427,N_8930);
xnor U14882 (N_14882,N_9487,N_11930);
or U14883 (N_14883,N_9201,N_8699);
nand U14884 (N_14884,N_9803,N_8335);
or U14885 (N_14885,N_10892,N_11365);
nor U14886 (N_14886,N_11638,N_11124);
or U14887 (N_14887,N_8374,N_8054);
nand U14888 (N_14888,N_8735,N_8723);
nand U14889 (N_14889,N_11551,N_8110);
nand U14890 (N_14890,N_10777,N_10301);
nand U14891 (N_14891,N_9704,N_8290);
nand U14892 (N_14892,N_9467,N_10003);
and U14893 (N_14893,N_9456,N_9831);
or U14894 (N_14894,N_10693,N_10714);
nor U14895 (N_14895,N_11577,N_10232);
nor U14896 (N_14896,N_9332,N_11930);
and U14897 (N_14897,N_8854,N_9515);
nor U14898 (N_14898,N_11829,N_9251);
nor U14899 (N_14899,N_9662,N_8306);
and U14900 (N_14900,N_10457,N_10821);
or U14901 (N_14901,N_9140,N_11081);
or U14902 (N_14902,N_8379,N_11432);
nand U14903 (N_14903,N_10562,N_8756);
nor U14904 (N_14904,N_8629,N_8575);
nand U14905 (N_14905,N_9984,N_9767);
xor U14906 (N_14906,N_10049,N_9166);
or U14907 (N_14907,N_10342,N_11720);
nand U14908 (N_14908,N_11633,N_11074);
and U14909 (N_14909,N_10159,N_10854);
nor U14910 (N_14910,N_8407,N_9554);
and U14911 (N_14911,N_8877,N_11043);
nor U14912 (N_14912,N_10726,N_8265);
or U14913 (N_14913,N_8152,N_8442);
and U14914 (N_14914,N_11984,N_8800);
nand U14915 (N_14915,N_8443,N_8199);
nand U14916 (N_14916,N_9953,N_10621);
nor U14917 (N_14917,N_11823,N_10474);
nor U14918 (N_14918,N_11085,N_10267);
nor U14919 (N_14919,N_11250,N_9815);
nor U14920 (N_14920,N_11258,N_11239);
xor U14921 (N_14921,N_8758,N_11597);
nor U14922 (N_14922,N_9306,N_10302);
nand U14923 (N_14923,N_10720,N_9048);
and U14924 (N_14924,N_8909,N_9689);
nor U14925 (N_14925,N_9959,N_8886);
nor U14926 (N_14926,N_9272,N_9972);
or U14927 (N_14927,N_9252,N_10194);
nand U14928 (N_14928,N_9294,N_11867);
or U14929 (N_14929,N_10728,N_9156);
or U14930 (N_14930,N_8374,N_10287);
nor U14931 (N_14931,N_8945,N_11446);
nor U14932 (N_14932,N_9430,N_11729);
xnor U14933 (N_14933,N_11032,N_11915);
nor U14934 (N_14934,N_11956,N_10358);
xnor U14935 (N_14935,N_8886,N_10817);
and U14936 (N_14936,N_11067,N_8762);
or U14937 (N_14937,N_9359,N_10609);
nor U14938 (N_14938,N_10594,N_8495);
nor U14939 (N_14939,N_11496,N_11354);
or U14940 (N_14940,N_10179,N_9877);
nor U14941 (N_14941,N_10538,N_9161);
and U14942 (N_14942,N_10855,N_10543);
or U14943 (N_14943,N_10460,N_9900);
nor U14944 (N_14944,N_10419,N_10649);
nor U14945 (N_14945,N_9158,N_8058);
or U14946 (N_14946,N_8768,N_10996);
or U14947 (N_14947,N_8251,N_10368);
and U14948 (N_14948,N_11483,N_9089);
xor U14949 (N_14949,N_11381,N_9101);
nand U14950 (N_14950,N_8818,N_9988);
or U14951 (N_14951,N_9940,N_9180);
nand U14952 (N_14952,N_9602,N_11469);
or U14953 (N_14953,N_8854,N_11897);
nor U14954 (N_14954,N_9641,N_9044);
nand U14955 (N_14955,N_11178,N_11078);
nand U14956 (N_14956,N_8237,N_10001);
or U14957 (N_14957,N_11519,N_10609);
or U14958 (N_14958,N_10370,N_9173);
nor U14959 (N_14959,N_10259,N_9469);
nand U14960 (N_14960,N_9786,N_10795);
and U14961 (N_14961,N_8752,N_8406);
nor U14962 (N_14962,N_11495,N_10299);
and U14963 (N_14963,N_10424,N_8150);
or U14964 (N_14964,N_8122,N_9004);
and U14965 (N_14965,N_9474,N_8472);
nand U14966 (N_14966,N_9850,N_8753);
nor U14967 (N_14967,N_11428,N_9742);
nand U14968 (N_14968,N_10154,N_11556);
nand U14969 (N_14969,N_10367,N_10317);
or U14970 (N_14970,N_9667,N_8581);
or U14971 (N_14971,N_11272,N_11746);
or U14972 (N_14972,N_10531,N_9214);
or U14973 (N_14973,N_8910,N_8809);
nand U14974 (N_14974,N_11800,N_9319);
and U14975 (N_14975,N_10883,N_8073);
nor U14976 (N_14976,N_9906,N_11286);
nand U14977 (N_14977,N_9439,N_8530);
or U14978 (N_14978,N_10918,N_9235);
and U14979 (N_14979,N_10205,N_11840);
nand U14980 (N_14980,N_10616,N_10450);
or U14981 (N_14981,N_9784,N_8570);
and U14982 (N_14982,N_9832,N_11790);
and U14983 (N_14983,N_10410,N_11054);
or U14984 (N_14984,N_8703,N_8462);
xnor U14985 (N_14985,N_11984,N_8605);
nor U14986 (N_14986,N_11774,N_10830);
nor U14987 (N_14987,N_11812,N_10357);
nand U14988 (N_14988,N_9006,N_11733);
nand U14989 (N_14989,N_9663,N_8903);
nand U14990 (N_14990,N_11763,N_9710);
nand U14991 (N_14991,N_10648,N_9038);
xnor U14992 (N_14992,N_9529,N_8086);
and U14993 (N_14993,N_9285,N_8498);
nor U14994 (N_14994,N_8153,N_8331);
or U14995 (N_14995,N_10546,N_8819);
nand U14996 (N_14996,N_10272,N_8951);
or U14997 (N_14997,N_8963,N_10938);
or U14998 (N_14998,N_8371,N_9199);
nor U14999 (N_14999,N_10334,N_8576);
nand U15000 (N_15000,N_10073,N_9527);
xor U15001 (N_15001,N_8174,N_11051);
nor U15002 (N_15002,N_8630,N_8676);
and U15003 (N_15003,N_9787,N_11546);
nor U15004 (N_15004,N_11840,N_9207);
nand U15005 (N_15005,N_8569,N_11647);
nor U15006 (N_15006,N_9408,N_10596);
and U15007 (N_15007,N_8971,N_10542);
or U15008 (N_15008,N_8942,N_10987);
nor U15009 (N_15009,N_9076,N_10644);
and U15010 (N_15010,N_9234,N_8791);
and U15011 (N_15011,N_10625,N_11022);
or U15012 (N_15012,N_8538,N_11461);
and U15013 (N_15013,N_8869,N_9566);
or U15014 (N_15014,N_9512,N_9737);
nand U15015 (N_15015,N_8462,N_11721);
nor U15016 (N_15016,N_11570,N_8108);
or U15017 (N_15017,N_9147,N_11862);
and U15018 (N_15018,N_9310,N_8426);
and U15019 (N_15019,N_11871,N_10892);
or U15020 (N_15020,N_9713,N_11542);
or U15021 (N_15021,N_11136,N_8571);
xor U15022 (N_15022,N_10326,N_9018);
and U15023 (N_15023,N_10602,N_8122);
and U15024 (N_15024,N_8877,N_9045);
nand U15025 (N_15025,N_9673,N_10959);
and U15026 (N_15026,N_10759,N_10955);
nor U15027 (N_15027,N_8891,N_11481);
xnor U15028 (N_15028,N_9207,N_8632);
nand U15029 (N_15029,N_8726,N_11519);
and U15030 (N_15030,N_10071,N_10271);
nand U15031 (N_15031,N_10652,N_8422);
and U15032 (N_15032,N_10873,N_10150);
nand U15033 (N_15033,N_8495,N_10414);
nor U15034 (N_15034,N_11103,N_11901);
and U15035 (N_15035,N_9881,N_8617);
and U15036 (N_15036,N_10533,N_8783);
or U15037 (N_15037,N_10200,N_8120);
xnor U15038 (N_15038,N_9541,N_11216);
or U15039 (N_15039,N_9453,N_8084);
nand U15040 (N_15040,N_10406,N_11679);
and U15041 (N_15041,N_10759,N_11862);
nor U15042 (N_15042,N_10460,N_10848);
nor U15043 (N_15043,N_10014,N_10945);
or U15044 (N_15044,N_8303,N_9397);
and U15045 (N_15045,N_11269,N_11074);
or U15046 (N_15046,N_8568,N_9848);
or U15047 (N_15047,N_11052,N_9591);
nor U15048 (N_15048,N_10508,N_11112);
nand U15049 (N_15049,N_11353,N_11399);
or U15050 (N_15050,N_8935,N_11017);
nand U15051 (N_15051,N_11018,N_9640);
or U15052 (N_15052,N_8393,N_10244);
nor U15053 (N_15053,N_11921,N_11548);
and U15054 (N_15054,N_8541,N_8565);
xor U15055 (N_15055,N_8842,N_11854);
or U15056 (N_15056,N_8741,N_11471);
and U15057 (N_15057,N_9986,N_11906);
nor U15058 (N_15058,N_10883,N_9689);
and U15059 (N_15059,N_9856,N_8255);
nand U15060 (N_15060,N_10584,N_10646);
or U15061 (N_15061,N_10558,N_11658);
or U15062 (N_15062,N_9408,N_11651);
and U15063 (N_15063,N_11961,N_8324);
nand U15064 (N_15064,N_11351,N_8487);
nor U15065 (N_15065,N_10530,N_8103);
and U15066 (N_15066,N_9946,N_11910);
nand U15067 (N_15067,N_9238,N_8283);
xnor U15068 (N_15068,N_9300,N_11969);
xnor U15069 (N_15069,N_9975,N_9314);
nand U15070 (N_15070,N_10132,N_11687);
nand U15071 (N_15071,N_9816,N_10111);
or U15072 (N_15072,N_8699,N_8366);
nor U15073 (N_15073,N_8296,N_9171);
and U15074 (N_15074,N_8249,N_11624);
nor U15075 (N_15075,N_10240,N_8550);
nand U15076 (N_15076,N_11848,N_10763);
and U15077 (N_15077,N_9788,N_9160);
nand U15078 (N_15078,N_10894,N_10985);
and U15079 (N_15079,N_10415,N_9977);
xor U15080 (N_15080,N_11015,N_9254);
nand U15081 (N_15081,N_11710,N_9745);
or U15082 (N_15082,N_9180,N_9003);
nor U15083 (N_15083,N_10605,N_9470);
nand U15084 (N_15084,N_11325,N_8577);
nor U15085 (N_15085,N_11365,N_9703);
nor U15086 (N_15086,N_9802,N_11853);
xnor U15087 (N_15087,N_10570,N_8026);
nor U15088 (N_15088,N_8282,N_10334);
nand U15089 (N_15089,N_8977,N_11136);
nor U15090 (N_15090,N_11070,N_9549);
nand U15091 (N_15091,N_11236,N_9461);
or U15092 (N_15092,N_11004,N_8121);
or U15093 (N_15093,N_10043,N_10109);
nor U15094 (N_15094,N_8572,N_10213);
nor U15095 (N_15095,N_11102,N_10909);
nor U15096 (N_15096,N_11333,N_11369);
and U15097 (N_15097,N_11093,N_8269);
or U15098 (N_15098,N_8668,N_9836);
or U15099 (N_15099,N_10352,N_9994);
or U15100 (N_15100,N_10015,N_10689);
and U15101 (N_15101,N_11194,N_11067);
xnor U15102 (N_15102,N_11391,N_9273);
and U15103 (N_15103,N_8383,N_11341);
nand U15104 (N_15104,N_11535,N_11223);
nand U15105 (N_15105,N_9908,N_11439);
nand U15106 (N_15106,N_11982,N_8426);
nor U15107 (N_15107,N_9933,N_8366);
or U15108 (N_15108,N_8195,N_11541);
nand U15109 (N_15109,N_11767,N_8643);
or U15110 (N_15110,N_10006,N_9841);
nor U15111 (N_15111,N_8509,N_9004);
and U15112 (N_15112,N_11064,N_10920);
or U15113 (N_15113,N_8090,N_11493);
nor U15114 (N_15114,N_8349,N_11820);
and U15115 (N_15115,N_8963,N_8942);
nor U15116 (N_15116,N_9478,N_8356);
and U15117 (N_15117,N_11468,N_10095);
nand U15118 (N_15118,N_11039,N_9370);
nor U15119 (N_15119,N_9461,N_11158);
or U15120 (N_15120,N_9216,N_11887);
or U15121 (N_15121,N_8212,N_9042);
and U15122 (N_15122,N_9323,N_10373);
nand U15123 (N_15123,N_10986,N_9476);
nor U15124 (N_15124,N_11700,N_8862);
nor U15125 (N_15125,N_8571,N_8802);
or U15126 (N_15126,N_9449,N_10731);
or U15127 (N_15127,N_11700,N_10538);
nand U15128 (N_15128,N_10444,N_10052);
or U15129 (N_15129,N_9524,N_8586);
nor U15130 (N_15130,N_8733,N_8133);
nand U15131 (N_15131,N_8450,N_11345);
nand U15132 (N_15132,N_9430,N_9954);
nand U15133 (N_15133,N_11849,N_9097);
nand U15134 (N_15134,N_11737,N_11022);
or U15135 (N_15135,N_11902,N_9067);
or U15136 (N_15136,N_10388,N_9310);
nor U15137 (N_15137,N_8014,N_11372);
or U15138 (N_15138,N_11494,N_10000);
and U15139 (N_15139,N_9333,N_9523);
nor U15140 (N_15140,N_9695,N_10753);
or U15141 (N_15141,N_11860,N_10797);
nand U15142 (N_15142,N_8987,N_9934);
or U15143 (N_15143,N_8594,N_10994);
nor U15144 (N_15144,N_11917,N_9006);
or U15145 (N_15145,N_10939,N_9009);
and U15146 (N_15146,N_9831,N_10688);
or U15147 (N_15147,N_10093,N_10216);
nand U15148 (N_15148,N_8620,N_11785);
nor U15149 (N_15149,N_9896,N_10075);
nor U15150 (N_15150,N_10605,N_9407);
and U15151 (N_15151,N_9963,N_9776);
and U15152 (N_15152,N_8358,N_9733);
or U15153 (N_15153,N_10279,N_8323);
nand U15154 (N_15154,N_8021,N_8198);
nor U15155 (N_15155,N_9044,N_8843);
nor U15156 (N_15156,N_11403,N_9478);
and U15157 (N_15157,N_9162,N_9854);
and U15158 (N_15158,N_11014,N_10396);
or U15159 (N_15159,N_11653,N_11492);
and U15160 (N_15160,N_8439,N_9215);
nand U15161 (N_15161,N_11672,N_9973);
or U15162 (N_15162,N_9640,N_9242);
nor U15163 (N_15163,N_11461,N_9779);
or U15164 (N_15164,N_9238,N_11566);
and U15165 (N_15165,N_10060,N_8588);
or U15166 (N_15166,N_10792,N_9956);
nor U15167 (N_15167,N_11605,N_9901);
nor U15168 (N_15168,N_10653,N_11598);
nor U15169 (N_15169,N_10720,N_9676);
or U15170 (N_15170,N_11127,N_11410);
nor U15171 (N_15171,N_9644,N_8670);
or U15172 (N_15172,N_8793,N_8366);
or U15173 (N_15173,N_9865,N_10816);
and U15174 (N_15174,N_10998,N_8321);
nor U15175 (N_15175,N_10273,N_10296);
and U15176 (N_15176,N_11797,N_11181);
or U15177 (N_15177,N_10045,N_9977);
nand U15178 (N_15178,N_9859,N_9406);
nand U15179 (N_15179,N_11864,N_11638);
and U15180 (N_15180,N_8811,N_8688);
nor U15181 (N_15181,N_9686,N_9846);
or U15182 (N_15182,N_8312,N_11847);
nor U15183 (N_15183,N_10130,N_8083);
xor U15184 (N_15184,N_9662,N_11064);
or U15185 (N_15185,N_9282,N_11815);
nand U15186 (N_15186,N_10242,N_9089);
nand U15187 (N_15187,N_10391,N_11793);
or U15188 (N_15188,N_8116,N_9700);
or U15189 (N_15189,N_11742,N_8635);
nor U15190 (N_15190,N_11690,N_10771);
or U15191 (N_15191,N_8490,N_8470);
and U15192 (N_15192,N_8781,N_9868);
nor U15193 (N_15193,N_10687,N_8955);
and U15194 (N_15194,N_9134,N_11391);
nor U15195 (N_15195,N_10389,N_8753);
and U15196 (N_15196,N_11985,N_9051);
or U15197 (N_15197,N_8848,N_11567);
nor U15198 (N_15198,N_10091,N_8070);
or U15199 (N_15199,N_8900,N_9478);
nor U15200 (N_15200,N_11376,N_10744);
and U15201 (N_15201,N_10380,N_10789);
and U15202 (N_15202,N_11567,N_8660);
nor U15203 (N_15203,N_10872,N_10828);
nor U15204 (N_15204,N_8849,N_9036);
or U15205 (N_15205,N_9905,N_8545);
and U15206 (N_15206,N_11301,N_10062);
nand U15207 (N_15207,N_11544,N_8205);
nand U15208 (N_15208,N_10067,N_8792);
xor U15209 (N_15209,N_8890,N_10762);
nor U15210 (N_15210,N_11444,N_11532);
and U15211 (N_15211,N_8347,N_8086);
nor U15212 (N_15212,N_11864,N_11699);
nor U15213 (N_15213,N_8540,N_10276);
nand U15214 (N_15214,N_8945,N_9740);
or U15215 (N_15215,N_10642,N_11926);
xor U15216 (N_15216,N_8622,N_9637);
nor U15217 (N_15217,N_8660,N_10828);
and U15218 (N_15218,N_8134,N_11263);
nand U15219 (N_15219,N_9879,N_8982);
and U15220 (N_15220,N_8474,N_11194);
or U15221 (N_15221,N_11431,N_8492);
or U15222 (N_15222,N_10058,N_10886);
nand U15223 (N_15223,N_8035,N_9466);
nor U15224 (N_15224,N_11137,N_10727);
and U15225 (N_15225,N_8577,N_9587);
nand U15226 (N_15226,N_8337,N_8235);
nor U15227 (N_15227,N_11822,N_8915);
and U15228 (N_15228,N_9294,N_10493);
nand U15229 (N_15229,N_11066,N_10018);
xor U15230 (N_15230,N_11626,N_8629);
nor U15231 (N_15231,N_11102,N_8831);
or U15232 (N_15232,N_11365,N_10524);
nand U15233 (N_15233,N_8424,N_8655);
nand U15234 (N_15234,N_9464,N_9981);
nand U15235 (N_15235,N_9956,N_10219);
nor U15236 (N_15236,N_8804,N_10799);
or U15237 (N_15237,N_8992,N_10489);
and U15238 (N_15238,N_10758,N_9122);
nand U15239 (N_15239,N_10322,N_10385);
nor U15240 (N_15240,N_11898,N_8426);
or U15241 (N_15241,N_11821,N_9340);
or U15242 (N_15242,N_11691,N_8532);
or U15243 (N_15243,N_10523,N_9826);
nand U15244 (N_15244,N_8303,N_8156);
nand U15245 (N_15245,N_10290,N_9087);
nor U15246 (N_15246,N_10532,N_8518);
nand U15247 (N_15247,N_11361,N_10287);
nor U15248 (N_15248,N_8050,N_9735);
or U15249 (N_15249,N_9322,N_11106);
or U15250 (N_15250,N_10637,N_9754);
nor U15251 (N_15251,N_8175,N_9926);
and U15252 (N_15252,N_8167,N_10937);
or U15253 (N_15253,N_8849,N_11397);
nor U15254 (N_15254,N_11132,N_10623);
nand U15255 (N_15255,N_9234,N_9413);
nor U15256 (N_15256,N_8812,N_11847);
and U15257 (N_15257,N_8478,N_9489);
or U15258 (N_15258,N_9240,N_11146);
nor U15259 (N_15259,N_10065,N_11081);
nand U15260 (N_15260,N_11589,N_10262);
nand U15261 (N_15261,N_9492,N_11456);
nor U15262 (N_15262,N_10927,N_8511);
nand U15263 (N_15263,N_9292,N_11695);
and U15264 (N_15264,N_10465,N_9208);
nand U15265 (N_15265,N_10299,N_10343);
or U15266 (N_15266,N_10212,N_9909);
and U15267 (N_15267,N_10968,N_11090);
and U15268 (N_15268,N_9335,N_8616);
or U15269 (N_15269,N_10882,N_10317);
or U15270 (N_15270,N_11394,N_8072);
nor U15271 (N_15271,N_9768,N_11576);
or U15272 (N_15272,N_8877,N_11744);
and U15273 (N_15273,N_11589,N_9682);
nand U15274 (N_15274,N_8013,N_10296);
or U15275 (N_15275,N_10424,N_9081);
or U15276 (N_15276,N_9897,N_10447);
and U15277 (N_15277,N_9916,N_11127);
nor U15278 (N_15278,N_11054,N_11248);
nor U15279 (N_15279,N_8570,N_9013);
nor U15280 (N_15280,N_9027,N_10971);
and U15281 (N_15281,N_8449,N_10439);
nand U15282 (N_15282,N_9837,N_10909);
nor U15283 (N_15283,N_11496,N_9448);
or U15284 (N_15284,N_10702,N_9552);
nor U15285 (N_15285,N_11437,N_11711);
or U15286 (N_15286,N_10755,N_11024);
nand U15287 (N_15287,N_8895,N_11648);
and U15288 (N_15288,N_11203,N_10519);
or U15289 (N_15289,N_9020,N_10084);
nand U15290 (N_15290,N_11017,N_9394);
or U15291 (N_15291,N_8729,N_10509);
and U15292 (N_15292,N_11084,N_9441);
nor U15293 (N_15293,N_11698,N_9058);
nor U15294 (N_15294,N_8206,N_8961);
or U15295 (N_15295,N_9568,N_11661);
nand U15296 (N_15296,N_11508,N_10408);
and U15297 (N_15297,N_11973,N_8962);
and U15298 (N_15298,N_11944,N_11608);
and U15299 (N_15299,N_11616,N_10913);
nor U15300 (N_15300,N_10828,N_11031);
nor U15301 (N_15301,N_10164,N_10747);
and U15302 (N_15302,N_8976,N_11405);
nand U15303 (N_15303,N_8907,N_10937);
nand U15304 (N_15304,N_9106,N_8228);
nor U15305 (N_15305,N_9578,N_10440);
and U15306 (N_15306,N_11400,N_11780);
nor U15307 (N_15307,N_10180,N_9336);
and U15308 (N_15308,N_9187,N_10852);
and U15309 (N_15309,N_11358,N_8474);
or U15310 (N_15310,N_11774,N_8780);
or U15311 (N_15311,N_10490,N_10015);
nor U15312 (N_15312,N_10264,N_8062);
nand U15313 (N_15313,N_9692,N_10839);
nand U15314 (N_15314,N_10173,N_9015);
and U15315 (N_15315,N_8293,N_9836);
nand U15316 (N_15316,N_10887,N_11453);
and U15317 (N_15317,N_11213,N_8777);
and U15318 (N_15318,N_10353,N_9695);
xor U15319 (N_15319,N_8971,N_9610);
nand U15320 (N_15320,N_11428,N_8723);
or U15321 (N_15321,N_8805,N_10736);
nor U15322 (N_15322,N_9153,N_9643);
and U15323 (N_15323,N_8143,N_10947);
xor U15324 (N_15324,N_8714,N_11591);
nand U15325 (N_15325,N_11270,N_10657);
nand U15326 (N_15326,N_10210,N_9527);
nor U15327 (N_15327,N_11922,N_9166);
or U15328 (N_15328,N_10509,N_8027);
nand U15329 (N_15329,N_8336,N_11899);
or U15330 (N_15330,N_10473,N_11886);
nand U15331 (N_15331,N_10180,N_8513);
nor U15332 (N_15332,N_11024,N_11440);
and U15333 (N_15333,N_11457,N_8548);
nand U15334 (N_15334,N_8867,N_11128);
nor U15335 (N_15335,N_9578,N_10581);
nor U15336 (N_15336,N_11087,N_9568);
nand U15337 (N_15337,N_8852,N_11049);
and U15338 (N_15338,N_8543,N_11535);
nor U15339 (N_15339,N_8344,N_9074);
xnor U15340 (N_15340,N_9721,N_10419);
or U15341 (N_15341,N_10848,N_8119);
and U15342 (N_15342,N_10505,N_9397);
nand U15343 (N_15343,N_9561,N_11679);
nor U15344 (N_15344,N_10103,N_9067);
nand U15345 (N_15345,N_9890,N_10756);
and U15346 (N_15346,N_11678,N_10312);
or U15347 (N_15347,N_8278,N_11584);
and U15348 (N_15348,N_10769,N_9310);
or U15349 (N_15349,N_10945,N_9213);
and U15350 (N_15350,N_11193,N_8971);
nand U15351 (N_15351,N_11998,N_9060);
or U15352 (N_15352,N_9468,N_11642);
nor U15353 (N_15353,N_8558,N_11913);
nor U15354 (N_15354,N_11248,N_10366);
nor U15355 (N_15355,N_9031,N_10144);
nand U15356 (N_15356,N_10168,N_11904);
nor U15357 (N_15357,N_10572,N_8663);
xor U15358 (N_15358,N_10573,N_9096);
and U15359 (N_15359,N_10410,N_11046);
nand U15360 (N_15360,N_9864,N_11180);
or U15361 (N_15361,N_8934,N_9769);
or U15362 (N_15362,N_11918,N_8042);
and U15363 (N_15363,N_10895,N_10329);
and U15364 (N_15364,N_11833,N_9290);
and U15365 (N_15365,N_11732,N_11976);
or U15366 (N_15366,N_8654,N_9531);
or U15367 (N_15367,N_9004,N_9637);
nand U15368 (N_15368,N_11021,N_11731);
or U15369 (N_15369,N_10280,N_9447);
nand U15370 (N_15370,N_8139,N_11988);
and U15371 (N_15371,N_10837,N_11877);
and U15372 (N_15372,N_8747,N_9625);
and U15373 (N_15373,N_11460,N_11136);
or U15374 (N_15374,N_8632,N_10304);
and U15375 (N_15375,N_8866,N_9522);
nor U15376 (N_15376,N_10219,N_9069);
or U15377 (N_15377,N_9014,N_11657);
nor U15378 (N_15378,N_8136,N_10044);
nor U15379 (N_15379,N_8501,N_9079);
nor U15380 (N_15380,N_11086,N_11683);
and U15381 (N_15381,N_11209,N_11202);
nor U15382 (N_15382,N_10804,N_11664);
and U15383 (N_15383,N_9325,N_11991);
or U15384 (N_15384,N_9679,N_9068);
nor U15385 (N_15385,N_10697,N_11642);
nor U15386 (N_15386,N_11679,N_11783);
nor U15387 (N_15387,N_10747,N_10926);
and U15388 (N_15388,N_8114,N_10648);
and U15389 (N_15389,N_11549,N_10368);
and U15390 (N_15390,N_8507,N_8806);
and U15391 (N_15391,N_10524,N_11109);
nand U15392 (N_15392,N_9878,N_9049);
nor U15393 (N_15393,N_8534,N_8738);
or U15394 (N_15394,N_8453,N_10822);
or U15395 (N_15395,N_11429,N_11237);
nor U15396 (N_15396,N_10028,N_9693);
nand U15397 (N_15397,N_9684,N_8092);
and U15398 (N_15398,N_9528,N_10061);
nand U15399 (N_15399,N_11455,N_10335);
nor U15400 (N_15400,N_8891,N_11865);
nand U15401 (N_15401,N_8663,N_11455);
or U15402 (N_15402,N_11626,N_8028);
or U15403 (N_15403,N_10119,N_9235);
and U15404 (N_15404,N_10290,N_11033);
nand U15405 (N_15405,N_10403,N_8823);
and U15406 (N_15406,N_10796,N_8442);
nor U15407 (N_15407,N_11484,N_9004);
and U15408 (N_15408,N_11203,N_8613);
nand U15409 (N_15409,N_9391,N_11617);
and U15410 (N_15410,N_11470,N_11321);
nor U15411 (N_15411,N_9767,N_9718);
and U15412 (N_15412,N_9596,N_9741);
nand U15413 (N_15413,N_10600,N_10634);
and U15414 (N_15414,N_9210,N_11996);
nand U15415 (N_15415,N_11739,N_10762);
or U15416 (N_15416,N_8033,N_11021);
nand U15417 (N_15417,N_8011,N_8292);
and U15418 (N_15418,N_11939,N_9521);
nand U15419 (N_15419,N_8950,N_10095);
nor U15420 (N_15420,N_10665,N_9031);
nor U15421 (N_15421,N_10920,N_11118);
and U15422 (N_15422,N_9708,N_8179);
and U15423 (N_15423,N_8964,N_9274);
nor U15424 (N_15424,N_11605,N_8103);
and U15425 (N_15425,N_9924,N_8788);
nand U15426 (N_15426,N_10831,N_10534);
nand U15427 (N_15427,N_10258,N_8803);
or U15428 (N_15428,N_9335,N_11584);
nor U15429 (N_15429,N_10978,N_8205);
and U15430 (N_15430,N_11743,N_11540);
and U15431 (N_15431,N_8440,N_8794);
nor U15432 (N_15432,N_9779,N_10300);
nor U15433 (N_15433,N_10332,N_11461);
nand U15434 (N_15434,N_9490,N_11963);
or U15435 (N_15435,N_8097,N_8234);
or U15436 (N_15436,N_10208,N_8992);
nand U15437 (N_15437,N_10973,N_10582);
and U15438 (N_15438,N_11831,N_11839);
nor U15439 (N_15439,N_8770,N_10291);
and U15440 (N_15440,N_9937,N_8901);
nand U15441 (N_15441,N_8958,N_10686);
or U15442 (N_15442,N_10545,N_8842);
nor U15443 (N_15443,N_8530,N_8440);
or U15444 (N_15444,N_10593,N_9118);
and U15445 (N_15445,N_8596,N_8554);
or U15446 (N_15446,N_11055,N_8491);
nand U15447 (N_15447,N_9609,N_11871);
nor U15448 (N_15448,N_8186,N_9399);
nor U15449 (N_15449,N_11459,N_10434);
or U15450 (N_15450,N_11031,N_9806);
or U15451 (N_15451,N_10771,N_10290);
xor U15452 (N_15452,N_10524,N_9215);
and U15453 (N_15453,N_9063,N_11609);
and U15454 (N_15454,N_9091,N_8151);
and U15455 (N_15455,N_10798,N_11380);
and U15456 (N_15456,N_11231,N_8385);
nand U15457 (N_15457,N_9540,N_10113);
nand U15458 (N_15458,N_10302,N_10320);
and U15459 (N_15459,N_9955,N_11643);
or U15460 (N_15460,N_11883,N_9588);
xnor U15461 (N_15461,N_11730,N_9741);
nand U15462 (N_15462,N_10631,N_10548);
xnor U15463 (N_15463,N_11805,N_9414);
or U15464 (N_15464,N_8743,N_11680);
or U15465 (N_15465,N_11640,N_10421);
nor U15466 (N_15466,N_9760,N_9833);
nand U15467 (N_15467,N_11424,N_9881);
and U15468 (N_15468,N_8941,N_11844);
or U15469 (N_15469,N_8035,N_11409);
and U15470 (N_15470,N_10200,N_8444);
nor U15471 (N_15471,N_9731,N_8074);
xnor U15472 (N_15472,N_9501,N_11378);
nand U15473 (N_15473,N_9659,N_11954);
nor U15474 (N_15474,N_11474,N_9033);
or U15475 (N_15475,N_11185,N_9845);
and U15476 (N_15476,N_11602,N_10384);
nor U15477 (N_15477,N_9147,N_8915);
nand U15478 (N_15478,N_11470,N_9047);
nor U15479 (N_15479,N_9747,N_9279);
or U15480 (N_15480,N_9602,N_9030);
and U15481 (N_15481,N_11985,N_10757);
nand U15482 (N_15482,N_10500,N_10199);
and U15483 (N_15483,N_11497,N_9568);
or U15484 (N_15484,N_10368,N_9574);
or U15485 (N_15485,N_10801,N_11584);
or U15486 (N_15486,N_9916,N_10795);
nor U15487 (N_15487,N_8197,N_10608);
nor U15488 (N_15488,N_8744,N_10723);
nor U15489 (N_15489,N_8749,N_10229);
nor U15490 (N_15490,N_10820,N_11024);
nor U15491 (N_15491,N_9745,N_11353);
nor U15492 (N_15492,N_8988,N_9821);
nor U15493 (N_15493,N_10844,N_8572);
nand U15494 (N_15494,N_11916,N_8173);
nor U15495 (N_15495,N_8011,N_10329);
nand U15496 (N_15496,N_8496,N_10058);
nor U15497 (N_15497,N_9524,N_11962);
or U15498 (N_15498,N_9610,N_8176);
nand U15499 (N_15499,N_9014,N_11200);
and U15500 (N_15500,N_10887,N_11546);
or U15501 (N_15501,N_10817,N_11979);
nor U15502 (N_15502,N_11569,N_10560);
or U15503 (N_15503,N_9848,N_9490);
nor U15504 (N_15504,N_11111,N_8328);
or U15505 (N_15505,N_10998,N_9037);
nor U15506 (N_15506,N_11375,N_9132);
nor U15507 (N_15507,N_10827,N_11974);
nor U15508 (N_15508,N_11087,N_9061);
or U15509 (N_15509,N_8575,N_10654);
nor U15510 (N_15510,N_10277,N_10901);
or U15511 (N_15511,N_8806,N_9489);
nor U15512 (N_15512,N_11620,N_9028);
and U15513 (N_15513,N_9088,N_10722);
nor U15514 (N_15514,N_11823,N_11468);
and U15515 (N_15515,N_9033,N_8672);
nor U15516 (N_15516,N_11026,N_10661);
nand U15517 (N_15517,N_8787,N_10205);
or U15518 (N_15518,N_11865,N_9123);
or U15519 (N_15519,N_8498,N_8531);
or U15520 (N_15520,N_10037,N_8819);
nand U15521 (N_15521,N_10761,N_9775);
xor U15522 (N_15522,N_8341,N_9198);
or U15523 (N_15523,N_11305,N_8451);
nand U15524 (N_15524,N_11284,N_10249);
nand U15525 (N_15525,N_10230,N_10337);
and U15526 (N_15526,N_10719,N_11073);
nor U15527 (N_15527,N_10986,N_11753);
and U15528 (N_15528,N_11621,N_8957);
nand U15529 (N_15529,N_9063,N_10037);
nor U15530 (N_15530,N_11317,N_11597);
xor U15531 (N_15531,N_8448,N_11226);
nand U15532 (N_15532,N_11540,N_11613);
nand U15533 (N_15533,N_10456,N_8559);
nor U15534 (N_15534,N_8742,N_8342);
or U15535 (N_15535,N_10940,N_10584);
and U15536 (N_15536,N_10449,N_9536);
or U15537 (N_15537,N_8940,N_8116);
nand U15538 (N_15538,N_8994,N_11468);
nor U15539 (N_15539,N_10107,N_9877);
nand U15540 (N_15540,N_10763,N_10338);
nor U15541 (N_15541,N_10013,N_8770);
nand U15542 (N_15542,N_11804,N_11049);
and U15543 (N_15543,N_9493,N_9313);
and U15544 (N_15544,N_10960,N_11469);
nand U15545 (N_15545,N_9161,N_11747);
xnor U15546 (N_15546,N_9944,N_9990);
and U15547 (N_15547,N_8097,N_10077);
nand U15548 (N_15548,N_10808,N_10338);
or U15549 (N_15549,N_10029,N_10259);
or U15550 (N_15550,N_8624,N_11287);
nor U15551 (N_15551,N_11391,N_11403);
nand U15552 (N_15552,N_11436,N_11915);
and U15553 (N_15553,N_8055,N_11531);
and U15554 (N_15554,N_10225,N_8546);
and U15555 (N_15555,N_10233,N_10696);
xor U15556 (N_15556,N_9555,N_10538);
nor U15557 (N_15557,N_9797,N_8816);
nand U15558 (N_15558,N_8581,N_11444);
nand U15559 (N_15559,N_9621,N_10253);
nor U15560 (N_15560,N_11028,N_11467);
nand U15561 (N_15561,N_10475,N_10436);
and U15562 (N_15562,N_10242,N_9757);
or U15563 (N_15563,N_11191,N_8298);
nand U15564 (N_15564,N_9088,N_8881);
and U15565 (N_15565,N_9889,N_11165);
nand U15566 (N_15566,N_10797,N_9660);
nor U15567 (N_15567,N_8277,N_8750);
and U15568 (N_15568,N_11661,N_9445);
nand U15569 (N_15569,N_8850,N_8754);
nand U15570 (N_15570,N_8359,N_10334);
nand U15571 (N_15571,N_10884,N_10928);
or U15572 (N_15572,N_9793,N_10668);
or U15573 (N_15573,N_9726,N_9407);
or U15574 (N_15574,N_10532,N_10373);
nor U15575 (N_15575,N_11954,N_9503);
or U15576 (N_15576,N_9631,N_10531);
and U15577 (N_15577,N_8221,N_8149);
and U15578 (N_15578,N_9190,N_11483);
and U15579 (N_15579,N_8297,N_8760);
and U15580 (N_15580,N_10988,N_10383);
or U15581 (N_15581,N_11205,N_9137);
and U15582 (N_15582,N_9547,N_11303);
or U15583 (N_15583,N_9657,N_10784);
nor U15584 (N_15584,N_8139,N_10861);
nor U15585 (N_15585,N_11707,N_10216);
nand U15586 (N_15586,N_8068,N_11566);
nor U15587 (N_15587,N_10225,N_8915);
and U15588 (N_15588,N_8488,N_10904);
or U15589 (N_15589,N_10112,N_9795);
nand U15590 (N_15590,N_11167,N_8729);
and U15591 (N_15591,N_11646,N_10931);
and U15592 (N_15592,N_8570,N_11336);
nor U15593 (N_15593,N_9197,N_10528);
xor U15594 (N_15594,N_10091,N_11944);
nand U15595 (N_15595,N_8363,N_11898);
nor U15596 (N_15596,N_10441,N_8972);
nand U15597 (N_15597,N_9992,N_10701);
and U15598 (N_15598,N_11671,N_11487);
nor U15599 (N_15599,N_11976,N_10160);
or U15600 (N_15600,N_10496,N_10706);
or U15601 (N_15601,N_8957,N_10984);
or U15602 (N_15602,N_9657,N_11565);
nand U15603 (N_15603,N_11323,N_11286);
nor U15604 (N_15604,N_10516,N_9656);
or U15605 (N_15605,N_9377,N_9953);
and U15606 (N_15606,N_9786,N_8020);
nor U15607 (N_15607,N_9092,N_9529);
or U15608 (N_15608,N_11189,N_9668);
and U15609 (N_15609,N_8820,N_11842);
or U15610 (N_15610,N_9983,N_8566);
nand U15611 (N_15611,N_9329,N_8648);
and U15612 (N_15612,N_9276,N_9477);
xnor U15613 (N_15613,N_11325,N_8479);
or U15614 (N_15614,N_10461,N_10737);
nand U15615 (N_15615,N_10906,N_9306);
nand U15616 (N_15616,N_10956,N_11533);
nand U15617 (N_15617,N_8700,N_11055);
and U15618 (N_15618,N_9888,N_11036);
and U15619 (N_15619,N_8429,N_11278);
or U15620 (N_15620,N_8822,N_10737);
and U15621 (N_15621,N_9161,N_8104);
nand U15622 (N_15622,N_9568,N_9707);
nand U15623 (N_15623,N_11162,N_11559);
or U15624 (N_15624,N_10334,N_10011);
nand U15625 (N_15625,N_8773,N_9957);
nand U15626 (N_15626,N_8616,N_9952);
nand U15627 (N_15627,N_8498,N_9878);
or U15628 (N_15628,N_11847,N_8024);
xnor U15629 (N_15629,N_8353,N_11705);
and U15630 (N_15630,N_10500,N_10784);
nor U15631 (N_15631,N_11525,N_10944);
nor U15632 (N_15632,N_9375,N_9985);
or U15633 (N_15633,N_9177,N_11471);
and U15634 (N_15634,N_11153,N_10201);
nor U15635 (N_15635,N_11466,N_9913);
nor U15636 (N_15636,N_11779,N_11061);
nor U15637 (N_15637,N_10384,N_10120);
or U15638 (N_15638,N_9398,N_9344);
or U15639 (N_15639,N_11193,N_8476);
or U15640 (N_15640,N_11480,N_11318);
or U15641 (N_15641,N_10239,N_8263);
and U15642 (N_15642,N_10159,N_10885);
nor U15643 (N_15643,N_8771,N_10174);
and U15644 (N_15644,N_8768,N_10646);
xnor U15645 (N_15645,N_9998,N_11729);
xnor U15646 (N_15646,N_9563,N_10077);
and U15647 (N_15647,N_8315,N_9461);
xnor U15648 (N_15648,N_8450,N_11008);
nor U15649 (N_15649,N_9297,N_11241);
or U15650 (N_15650,N_11134,N_9554);
nor U15651 (N_15651,N_11716,N_8824);
and U15652 (N_15652,N_10828,N_10910);
and U15653 (N_15653,N_8451,N_11516);
and U15654 (N_15654,N_11444,N_8321);
and U15655 (N_15655,N_11428,N_9315);
nand U15656 (N_15656,N_9749,N_11067);
nor U15657 (N_15657,N_9401,N_11201);
and U15658 (N_15658,N_9719,N_8275);
nand U15659 (N_15659,N_8432,N_9050);
or U15660 (N_15660,N_9855,N_11434);
nor U15661 (N_15661,N_11028,N_8183);
or U15662 (N_15662,N_9125,N_11361);
nand U15663 (N_15663,N_10685,N_11172);
nor U15664 (N_15664,N_9503,N_10422);
nor U15665 (N_15665,N_11258,N_9163);
and U15666 (N_15666,N_8743,N_8271);
nor U15667 (N_15667,N_8055,N_10431);
nand U15668 (N_15668,N_8724,N_11217);
xor U15669 (N_15669,N_9959,N_11494);
or U15670 (N_15670,N_10199,N_9571);
or U15671 (N_15671,N_9406,N_9731);
or U15672 (N_15672,N_11508,N_10236);
nand U15673 (N_15673,N_9063,N_11080);
nor U15674 (N_15674,N_9238,N_8495);
and U15675 (N_15675,N_9151,N_10545);
and U15676 (N_15676,N_11581,N_8185);
and U15677 (N_15677,N_11775,N_9300);
nor U15678 (N_15678,N_8402,N_8882);
and U15679 (N_15679,N_10542,N_10710);
xor U15680 (N_15680,N_9612,N_9997);
nand U15681 (N_15681,N_8514,N_11970);
nand U15682 (N_15682,N_8285,N_11862);
xor U15683 (N_15683,N_10724,N_9254);
nor U15684 (N_15684,N_9668,N_8064);
nor U15685 (N_15685,N_10513,N_8875);
nor U15686 (N_15686,N_10525,N_11499);
nand U15687 (N_15687,N_9562,N_9070);
nand U15688 (N_15688,N_9237,N_10699);
and U15689 (N_15689,N_9557,N_8886);
nor U15690 (N_15690,N_10609,N_10899);
nand U15691 (N_15691,N_10267,N_10278);
nand U15692 (N_15692,N_10074,N_11673);
xnor U15693 (N_15693,N_10556,N_11422);
xor U15694 (N_15694,N_10414,N_8300);
nor U15695 (N_15695,N_10236,N_10894);
or U15696 (N_15696,N_11796,N_11069);
or U15697 (N_15697,N_9256,N_9977);
nand U15698 (N_15698,N_8066,N_10433);
nand U15699 (N_15699,N_8978,N_8911);
and U15700 (N_15700,N_9267,N_11429);
and U15701 (N_15701,N_11216,N_8760);
and U15702 (N_15702,N_11927,N_11419);
nor U15703 (N_15703,N_11472,N_9315);
nor U15704 (N_15704,N_8835,N_11761);
or U15705 (N_15705,N_9075,N_10935);
nand U15706 (N_15706,N_8977,N_9460);
nor U15707 (N_15707,N_9029,N_9834);
and U15708 (N_15708,N_9864,N_9787);
and U15709 (N_15709,N_10241,N_8293);
and U15710 (N_15710,N_8419,N_8343);
or U15711 (N_15711,N_11781,N_8232);
nand U15712 (N_15712,N_9017,N_9687);
or U15713 (N_15713,N_10693,N_10712);
nor U15714 (N_15714,N_9558,N_11991);
or U15715 (N_15715,N_9715,N_11816);
or U15716 (N_15716,N_9030,N_11248);
nor U15717 (N_15717,N_8707,N_8767);
or U15718 (N_15718,N_8471,N_11803);
nor U15719 (N_15719,N_10839,N_8383);
xnor U15720 (N_15720,N_11942,N_8784);
or U15721 (N_15721,N_9329,N_9608);
and U15722 (N_15722,N_10558,N_9054);
nand U15723 (N_15723,N_8207,N_11966);
or U15724 (N_15724,N_9542,N_8202);
nor U15725 (N_15725,N_10799,N_9211);
nor U15726 (N_15726,N_8818,N_11612);
nor U15727 (N_15727,N_9110,N_8288);
and U15728 (N_15728,N_10333,N_9392);
and U15729 (N_15729,N_10364,N_9562);
and U15730 (N_15730,N_11955,N_8934);
nand U15731 (N_15731,N_8735,N_9886);
or U15732 (N_15732,N_10401,N_10304);
or U15733 (N_15733,N_8459,N_10569);
nor U15734 (N_15734,N_8564,N_10718);
nor U15735 (N_15735,N_11489,N_10841);
or U15736 (N_15736,N_10981,N_11880);
and U15737 (N_15737,N_8526,N_11390);
and U15738 (N_15738,N_8348,N_11215);
nand U15739 (N_15739,N_11564,N_11744);
or U15740 (N_15740,N_8305,N_10892);
and U15741 (N_15741,N_9834,N_9909);
and U15742 (N_15742,N_10079,N_11132);
nand U15743 (N_15743,N_8685,N_10333);
nand U15744 (N_15744,N_10170,N_9286);
and U15745 (N_15745,N_10660,N_11891);
nor U15746 (N_15746,N_8567,N_9596);
nand U15747 (N_15747,N_8142,N_11285);
and U15748 (N_15748,N_10974,N_9844);
nand U15749 (N_15749,N_10792,N_9249);
nor U15750 (N_15750,N_10162,N_9154);
nand U15751 (N_15751,N_10290,N_8506);
and U15752 (N_15752,N_10448,N_9911);
and U15753 (N_15753,N_9868,N_9816);
nor U15754 (N_15754,N_10442,N_11685);
nand U15755 (N_15755,N_9139,N_8013);
and U15756 (N_15756,N_10880,N_10887);
nor U15757 (N_15757,N_10194,N_9765);
or U15758 (N_15758,N_10517,N_9056);
and U15759 (N_15759,N_11202,N_9771);
and U15760 (N_15760,N_11213,N_8154);
and U15761 (N_15761,N_8657,N_11770);
and U15762 (N_15762,N_9040,N_9473);
and U15763 (N_15763,N_10522,N_9643);
or U15764 (N_15764,N_8270,N_10305);
or U15765 (N_15765,N_8007,N_10328);
or U15766 (N_15766,N_10176,N_8621);
and U15767 (N_15767,N_8594,N_11762);
nand U15768 (N_15768,N_10966,N_10954);
nor U15769 (N_15769,N_11517,N_10923);
nand U15770 (N_15770,N_10339,N_8420);
nor U15771 (N_15771,N_11584,N_10343);
nor U15772 (N_15772,N_11963,N_8907);
nor U15773 (N_15773,N_11976,N_11920);
and U15774 (N_15774,N_10788,N_9396);
nand U15775 (N_15775,N_9552,N_9549);
nand U15776 (N_15776,N_8865,N_11997);
or U15777 (N_15777,N_9150,N_8413);
nand U15778 (N_15778,N_10264,N_9468);
or U15779 (N_15779,N_10753,N_8697);
nand U15780 (N_15780,N_11526,N_11350);
or U15781 (N_15781,N_9331,N_10029);
nand U15782 (N_15782,N_11067,N_8449);
or U15783 (N_15783,N_11112,N_11358);
and U15784 (N_15784,N_11683,N_8742);
and U15785 (N_15785,N_8038,N_8413);
or U15786 (N_15786,N_11239,N_9362);
xnor U15787 (N_15787,N_9422,N_8976);
and U15788 (N_15788,N_9222,N_9546);
and U15789 (N_15789,N_8213,N_11234);
nor U15790 (N_15790,N_11113,N_9877);
nand U15791 (N_15791,N_11806,N_8169);
or U15792 (N_15792,N_11424,N_10181);
or U15793 (N_15793,N_9680,N_10699);
nand U15794 (N_15794,N_11428,N_10600);
or U15795 (N_15795,N_10974,N_8975);
nand U15796 (N_15796,N_10458,N_11483);
nand U15797 (N_15797,N_10447,N_10873);
nor U15798 (N_15798,N_11608,N_9015);
and U15799 (N_15799,N_10345,N_11878);
nor U15800 (N_15800,N_10479,N_8770);
or U15801 (N_15801,N_8944,N_11440);
or U15802 (N_15802,N_11059,N_8396);
nor U15803 (N_15803,N_9916,N_9740);
and U15804 (N_15804,N_8356,N_8692);
and U15805 (N_15805,N_8843,N_11572);
or U15806 (N_15806,N_11407,N_11074);
nor U15807 (N_15807,N_8097,N_9957);
nor U15808 (N_15808,N_10050,N_9910);
nand U15809 (N_15809,N_8604,N_9411);
nor U15810 (N_15810,N_9835,N_11243);
nand U15811 (N_15811,N_11935,N_9093);
nand U15812 (N_15812,N_9089,N_8146);
nor U15813 (N_15813,N_11218,N_10055);
or U15814 (N_15814,N_11647,N_11302);
nand U15815 (N_15815,N_10668,N_9727);
and U15816 (N_15816,N_10194,N_10260);
nand U15817 (N_15817,N_10937,N_8498);
nor U15818 (N_15818,N_10472,N_10024);
nor U15819 (N_15819,N_11614,N_8788);
or U15820 (N_15820,N_9800,N_10223);
nor U15821 (N_15821,N_9001,N_9257);
and U15822 (N_15822,N_9744,N_9925);
xnor U15823 (N_15823,N_10245,N_9039);
nand U15824 (N_15824,N_10463,N_9574);
or U15825 (N_15825,N_8838,N_11430);
xor U15826 (N_15826,N_11671,N_11186);
nand U15827 (N_15827,N_11354,N_9925);
or U15828 (N_15828,N_8376,N_11876);
nand U15829 (N_15829,N_10305,N_10780);
nand U15830 (N_15830,N_8207,N_9183);
and U15831 (N_15831,N_8226,N_9610);
or U15832 (N_15832,N_10958,N_8245);
and U15833 (N_15833,N_11479,N_11758);
and U15834 (N_15834,N_8810,N_9649);
nor U15835 (N_15835,N_8594,N_10158);
nor U15836 (N_15836,N_10764,N_11719);
or U15837 (N_15837,N_10588,N_11547);
nand U15838 (N_15838,N_10312,N_9479);
nand U15839 (N_15839,N_9367,N_10927);
nor U15840 (N_15840,N_10030,N_11552);
and U15841 (N_15841,N_11102,N_11409);
or U15842 (N_15842,N_11468,N_11672);
or U15843 (N_15843,N_10790,N_8700);
and U15844 (N_15844,N_8818,N_11484);
and U15845 (N_15845,N_9486,N_11878);
nand U15846 (N_15846,N_10154,N_11642);
or U15847 (N_15847,N_11778,N_11332);
nand U15848 (N_15848,N_10504,N_9282);
or U15849 (N_15849,N_9247,N_9884);
nor U15850 (N_15850,N_8972,N_9091);
or U15851 (N_15851,N_11847,N_11044);
nand U15852 (N_15852,N_9796,N_11450);
nor U15853 (N_15853,N_9826,N_10552);
and U15854 (N_15854,N_8559,N_8508);
or U15855 (N_15855,N_8524,N_11359);
and U15856 (N_15856,N_9452,N_8519);
nand U15857 (N_15857,N_11876,N_9650);
nor U15858 (N_15858,N_8638,N_11937);
nand U15859 (N_15859,N_11374,N_10064);
nand U15860 (N_15860,N_11107,N_10708);
xnor U15861 (N_15861,N_11031,N_9522);
or U15862 (N_15862,N_10225,N_11977);
or U15863 (N_15863,N_11138,N_9892);
and U15864 (N_15864,N_9127,N_10327);
nor U15865 (N_15865,N_10137,N_10712);
or U15866 (N_15866,N_9236,N_8028);
nand U15867 (N_15867,N_10631,N_8100);
xnor U15868 (N_15868,N_11481,N_9053);
nor U15869 (N_15869,N_10218,N_11791);
nand U15870 (N_15870,N_9546,N_9716);
or U15871 (N_15871,N_8941,N_8220);
nand U15872 (N_15872,N_8023,N_10261);
nor U15873 (N_15873,N_9194,N_11595);
or U15874 (N_15874,N_8632,N_8003);
nor U15875 (N_15875,N_8000,N_11302);
or U15876 (N_15876,N_8651,N_10110);
nand U15877 (N_15877,N_11124,N_11758);
nor U15878 (N_15878,N_11685,N_8055);
or U15879 (N_15879,N_9366,N_8512);
nor U15880 (N_15880,N_10522,N_10691);
and U15881 (N_15881,N_8996,N_9889);
xor U15882 (N_15882,N_8882,N_8456);
or U15883 (N_15883,N_10709,N_9452);
and U15884 (N_15884,N_11107,N_11829);
nor U15885 (N_15885,N_10904,N_11000);
nand U15886 (N_15886,N_11167,N_10168);
and U15887 (N_15887,N_9079,N_8584);
nand U15888 (N_15888,N_8663,N_9644);
or U15889 (N_15889,N_10541,N_8252);
nand U15890 (N_15890,N_9368,N_11583);
or U15891 (N_15891,N_9824,N_11473);
and U15892 (N_15892,N_10866,N_10595);
or U15893 (N_15893,N_11738,N_9119);
nor U15894 (N_15894,N_10124,N_10150);
xnor U15895 (N_15895,N_9875,N_8811);
or U15896 (N_15896,N_8410,N_10714);
nand U15897 (N_15897,N_9741,N_10483);
nor U15898 (N_15898,N_9578,N_9081);
nand U15899 (N_15899,N_8085,N_9052);
nor U15900 (N_15900,N_11924,N_8207);
nand U15901 (N_15901,N_11604,N_11590);
nor U15902 (N_15902,N_8723,N_8354);
nor U15903 (N_15903,N_9159,N_10621);
nor U15904 (N_15904,N_11759,N_9482);
or U15905 (N_15905,N_8375,N_10807);
or U15906 (N_15906,N_8135,N_9540);
or U15907 (N_15907,N_8145,N_8956);
or U15908 (N_15908,N_10050,N_11997);
or U15909 (N_15909,N_11889,N_8696);
or U15910 (N_15910,N_11172,N_11403);
nor U15911 (N_15911,N_11258,N_9192);
and U15912 (N_15912,N_8346,N_8255);
xnor U15913 (N_15913,N_8077,N_9173);
nand U15914 (N_15914,N_11066,N_10471);
nor U15915 (N_15915,N_11215,N_8927);
or U15916 (N_15916,N_9000,N_8166);
nand U15917 (N_15917,N_10968,N_10576);
and U15918 (N_15918,N_8994,N_11055);
nor U15919 (N_15919,N_11435,N_10641);
or U15920 (N_15920,N_8571,N_8123);
or U15921 (N_15921,N_10454,N_9915);
nand U15922 (N_15922,N_10367,N_10028);
nor U15923 (N_15923,N_8077,N_8686);
and U15924 (N_15924,N_10193,N_8579);
or U15925 (N_15925,N_11290,N_11659);
and U15926 (N_15926,N_8281,N_8962);
nand U15927 (N_15927,N_9328,N_11234);
or U15928 (N_15928,N_8636,N_8192);
or U15929 (N_15929,N_8913,N_9028);
nor U15930 (N_15930,N_10019,N_10766);
and U15931 (N_15931,N_11574,N_8204);
nand U15932 (N_15932,N_9565,N_9114);
nor U15933 (N_15933,N_11858,N_11288);
nand U15934 (N_15934,N_8506,N_11996);
or U15935 (N_15935,N_8524,N_10026);
or U15936 (N_15936,N_10361,N_11555);
nor U15937 (N_15937,N_10574,N_11144);
nor U15938 (N_15938,N_11170,N_8291);
nor U15939 (N_15939,N_9462,N_10600);
or U15940 (N_15940,N_11969,N_8341);
nand U15941 (N_15941,N_9203,N_11874);
and U15942 (N_15942,N_10031,N_9432);
nor U15943 (N_15943,N_10269,N_10975);
and U15944 (N_15944,N_9029,N_9594);
and U15945 (N_15945,N_11321,N_11444);
and U15946 (N_15946,N_8690,N_9201);
and U15947 (N_15947,N_10579,N_11504);
or U15948 (N_15948,N_9312,N_8416);
nand U15949 (N_15949,N_8712,N_9059);
or U15950 (N_15950,N_8054,N_9483);
and U15951 (N_15951,N_8907,N_8601);
nor U15952 (N_15952,N_11331,N_11615);
or U15953 (N_15953,N_9682,N_10521);
nor U15954 (N_15954,N_11731,N_11392);
or U15955 (N_15955,N_10234,N_10879);
nand U15956 (N_15956,N_8225,N_9191);
nand U15957 (N_15957,N_11519,N_11381);
nand U15958 (N_15958,N_9074,N_9568);
or U15959 (N_15959,N_9105,N_10603);
nor U15960 (N_15960,N_11712,N_10365);
or U15961 (N_15961,N_10734,N_8840);
or U15962 (N_15962,N_11563,N_10326);
nand U15963 (N_15963,N_9807,N_10457);
or U15964 (N_15964,N_11098,N_10266);
and U15965 (N_15965,N_9216,N_11918);
and U15966 (N_15966,N_8376,N_10592);
and U15967 (N_15967,N_8640,N_11986);
nor U15968 (N_15968,N_8405,N_9335);
or U15969 (N_15969,N_10749,N_9624);
and U15970 (N_15970,N_11675,N_11593);
nor U15971 (N_15971,N_10704,N_10867);
or U15972 (N_15972,N_9128,N_9079);
nand U15973 (N_15973,N_9871,N_8933);
and U15974 (N_15974,N_11997,N_8857);
or U15975 (N_15975,N_10364,N_10187);
nand U15976 (N_15976,N_10614,N_8547);
nand U15977 (N_15977,N_8075,N_8589);
and U15978 (N_15978,N_8651,N_8261);
and U15979 (N_15979,N_9481,N_10508);
xnor U15980 (N_15980,N_10650,N_8348);
nand U15981 (N_15981,N_11963,N_9573);
and U15982 (N_15982,N_10328,N_11685);
or U15983 (N_15983,N_11993,N_9488);
nand U15984 (N_15984,N_9384,N_10982);
nor U15985 (N_15985,N_9830,N_8431);
nand U15986 (N_15986,N_11229,N_11813);
nand U15987 (N_15987,N_8210,N_10276);
or U15988 (N_15988,N_11931,N_11271);
or U15989 (N_15989,N_11950,N_11346);
or U15990 (N_15990,N_9901,N_10401);
nor U15991 (N_15991,N_9267,N_9078);
and U15992 (N_15992,N_10541,N_11844);
and U15993 (N_15993,N_11154,N_10057);
nand U15994 (N_15994,N_11155,N_8944);
nand U15995 (N_15995,N_9215,N_9856);
nor U15996 (N_15996,N_11376,N_8669);
nand U15997 (N_15997,N_10102,N_9244);
or U15998 (N_15998,N_8229,N_9247);
and U15999 (N_15999,N_10673,N_11875);
nor U16000 (N_16000,N_14462,N_14737);
and U16001 (N_16001,N_15881,N_15052);
and U16002 (N_16002,N_14271,N_15014);
and U16003 (N_16003,N_15422,N_14708);
and U16004 (N_16004,N_15572,N_15170);
nor U16005 (N_16005,N_13546,N_12948);
nand U16006 (N_16006,N_15593,N_14145);
nand U16007 (N_16007,N_14486,N_15661);
and U16008 (N_16008,N_14063,N_13977);
nor U16009 (N_16009,N_13987,N_15035);
and U16010 (N_16010,N_12162,N_12098);
or U16011 (N_16011,N_13081,N_14764);
or U16012 (N_16012,N_12703,N_13235);
nand U16013 (N_16013,N_14626,N_12242);
nand U16014 (N_16014,N_13301,N_15855);
and U16015 (N_16015,N_15522,N_12040);
nor U16016 (N_16016,N_12296,N_13268);
nor U16017 (N_16017,N_14204,N_13732);
nand U16018 (N_16018,N_15120,N_12707);
or U16019 (N_16019,N_13808,N_14293);
or U16020 (N_16020,N_15512,N_13325);
or U16021 (N_16021,N_14912,N_12491);
and U16022 (N_16022,N_14705,N_15636);
or U16023 (N_16023,N_13172,N_14987);
and U16024 (N_16024,N_15954,N_13509);
or U16025 (N_16025,N_15911,N_15471);
nand U16026 (N_16026,N_13078,N_14294);
or U16027 (N_16027,N_13539,N_12604);
or U16028 (N_16028,N_15785,N_14832);
or U16029 (N_16029,N_14407,N_14335);
nand U16030 (N_16030,N_12980,N_12579);
nor U16031 (N_16031,N_12515,N_15018);
and U16032 (N_16032,N_15331,N_15513);
and U16033 (N_16033,N_15118,N_13332);
nor U16034 (N_16034,N_14288,N_14472);
or U16035 (N_16035,N_15233,N_14879);
or U16036 (N_16036,N_15001,N_13338);
or U16037 (N_16037,N_14700,N_14697);
or U16038 (N_16038,N_13963,N_13531);
xor U16039 (N_16039,N_13713,N_12208);
and U16040 (N_16040,N_12812,N_15926);
nand U16041 (N_16041,N_15378,N_15934);
or U16042 (N_16042,N_15298,N_14985);
or U16043 (N_16043,N_12601,N_13174);
nand U16044 (N_16044,N_12001,N_15822);
nand U16045 (N_16045,N_12577,N_12788);
or U16046 (N_16046,N_13851,N_15858);
nand U16047 (N_16047,N_12047,N_12906);
or U16048 (N_16048,N_14215,N_14853);
nor U16049 (N_16049,N_12751,N_15224);
nor U16050 (N_16050,N_14352,N_15130);
or U16051 (N_16051,N_13917,N_13544);
nor U16052 (N_16052,N_12182,N_15024);
nor U16053 (N_16053,N_12841,N_15481);
and U16054 (N_16054,N_14395,N_14238);
or U16055 (N_16055,N_14174,N_15407);
nor U16056 (N_16056,N_15996,N_12218);
nand U16057 (N_16057,N_13767,N_13970);
and U16058 (N_16058,N_12988,N_13876);
or U16059 (N_16059,N_14451,N_12715);
nor U16060 (N_16060,N_15708,N_14153);
or U16061 (N_16061,N_13303,N_12360);
or U16062 (N_16062,N_14459,N_12900);
or U16063 (N_16063,N_12741,N_15189);
and U16064 (N_16064,N_12957,N_12195);
and U16065 (N_16065,N_12172,N_15041);
nor U16066 (N_16066,N_15444,N_15240);
xor U16067 (N_16067,N_13563,N_13910);
and U16068 (N_16068,N_15975,N_14787);
or U16069 (N_16069,N_14066,N_13961);
or U16070 (N_16070,N_15879,N_15664);
nor U16071 (N_16071,N_14638,N_14006);
nor U16072 (N_16072,N_14824,N_15648);
or U16073 (N_16073,N_15354,N_15909);
or U16074 (N_16074,N_12916,N_12339);
nand U16075 (N_16075,N_13111,N_14506);
nand U16076 (N_16076,N_15562,N_13881);
or U16077 (N_16077,N_13688,N_15326);
nor U16078 (N_16078,N_12718,N_12637);
or U16079 (N_16079,N_13266,N_13311);
and U16080 (N_16080,N_13030,N_13681);
and U16081 (N_16081,N_15125,N_15178);
nor U16082 (N_16082,N_13179,N_14939);
nand U16083 (N_16083,N_12091,N_15577);
nor U16084 (N_16084,N_13424,N_12634);
nand U16085 (N_16085,N_13089,N_14992);
nand U16086 (N_16086,N_12620,N_15773);
nand U16087 (N_16087,N_14368,N_14920);
and U16088 (N_16088,N_14723,N_14808);
nand U16089 (N_16089,N_14241,N_15043);
and U16090 (N_16090,N_14566,N_12768);
and U16091 (N_16091,N_15974,N_12354);
or U16092 (N_16092,N_15783,N_14617);
or U16093 (N_16093,N_13597,N_12553);
nor U16094 (N_16094,N_14989,N_13019);
or U16095 (N_16095,N_14849,N_14039);
nor U16096 (N_16096,N_13128,N_12781);
and U16097 (N_16097,N_14953,N_14036);
and U16098 (N_16098,N_13516,N_13819);
nand U16099 (N_16099,N_14544,N_14221);
nand U16100 (N_16100,N_15750,N_13557);
or U16101 (N_16101,N_14323,N_12490);
and U16102 (N_16102,N_14387,N_13928);
and U16103 (N_16103,N_15660,N_15337);
nor U16104 (N_16104,N_12519,N_15635);
or U16105 (N_16105,N_14634,N_15784);
and U16106 (N_16106,N_13387,N_13122);
and U16107 (N_16107,N_14275,N_14416);
nand U16108 (N_16108,N_13279,N_15255);
and U16109 (N_16109,N_13190,N_14056);
or U16110 (N_16110,N_15393,N_12019);
xor U16111 (N_16111,N_12855,N_12960);
and U16112 (N_16112,N_14232,N_15609);
xor U16113 (N_16113,N_13933,N_13050);
nand U16114 (N_16114,N_12365,N_15992);
or U16115 (N_16115,N_12578,N_12910);
or U16116 (N_16116,N_14347,N_15967);
nor U16117 (N_16117,N_13411,N_13796);
and U16118 (N_16118,N_13764,N_13393);
or U16119 (N_16119,N_13288,N_12726);
nand U16120 (N_16120,N_14234,N_12119);
or U16121 (N_16121,N_14786,N_15551);
and U16122 (N_16122,N_12454,N_12309);
or U16123 (N_16123,N_12028,N_13771);
nor U16124 (N_16124,N_15281,N_13697);
nor U16125 (N_16125,N_14311,N_12138);
and U16126 (N_16126,N_15663,N_12679);
xnor U16127 (N_16127,N_13159,N_14718);
nand U16128 (N_16128,N_13676,N_13185);
or U16129 (N_16129,N_14150,N_13946);
and U16130 (N_16130,N_12264,N_14514);
xnor U16131 (N_16131,N_14356,N_12273);
nor U16132 (N_16132,N_12016,N_15433);
nor U16133 (N_16133,N_14198,N_12097);
nand U16134 (N_16134,N_14976,N_14709);
or U16135 (N_16135,N_12389,N_15451);
nor U16136 (N_16136,N_14279,N_15864);
or U16137 (N_16137,N_12773,N_13745);
nor U16138 (N_16138,N_15234,N_13919);
nor U16139 (N_16139,N_13617,N_14929);
and U16140 (N_16140,N_12598,N_12720);
and U16141 (N_16141,N_13780,N_14391);
nor U16142 (N_16142,N_12446,N_13154);
nor U16143 (N_16143,N_12778,N_12233);
nand U16144 (N_16144,N_14115,N_13907);
and U16145 (N_16145,N_13355,N_13960);
nor U16146 (N_16146,N_13621,N_13052);
and U16147 (N_16147,N_13890,N_15594);
or U16148 (N_16148,N_12771,N_12624);
or U16149 (N_16149,N_14586,N_15537);
nand U16150 (N_16150,N_13426,N_15491);
and U16151 (N_16151,N_13094,N_15253);
or U16152 (N_16152,N_15077,N_13414);
or U16153 (N_16153,N_12469,N_12511);
or U16154 (N_16154,N_12735,N_13313);
and U16155 (N_16155,N_12583,N_12629);
or U16156 (N_16156,N_13552,N_14968);
xnor U16157 (N_16157,N_14137,N_14870);
or U16158 (N_16158,N_15929,N_12465);
or U16159 (N_16159,N_13416,N_12608);
or U16160 (N_16160,N_13187,N_15579);
or U16161 (N_16161,N_13229,N_15022);
nand U16162 (N_16162,N_15514,N_13517);
or U16163 (N_16163,N_12427,N_14623);
or U16164 (N_16164,N_13364,N_15403);
nand U16165 (N_16165,N_15436,N_14533);
nor U16166 (N_16166,N_12954,N_15817);
nand U16167 (N_16167,N_13302,N_12056);
nor U16168 (N_16168,N_14088,N_12840);
or U16169 (N_16169,N_13500,N_14072);
nand U16170 (N_16170,N_14037,N_12582);
nand U16171 (N_16171,N_13690,N_14038);
nand U16172 (N_16172,N_15716,N_15628);
and U16173 (N_16173,N_14122,N_12657);
and U16174 (N_16174,N_13988,N_14995);
and U16175 (N_16175,N_13930,N_13334);
nand U16176 (N_16176,N_14339,N_15870);
nand U16177 (N_16177,N_14731,N_13659);
nand U16178 (N_16178,N_15756,N_14098);
and U16179 (N_16179,N_13282,N_14518);
nor U16180 (N_16180,N_15568,N_14011);
and U16181 (N_16181,N_15739,N_13213);
nor U16182 (N_16182,N_14013,N_13465);
xor U16183 (N_16183,N_14172,N_15396);
nand U16184 (N_16184,N_14707,N_12912);
and U16185 (N_16185,N_15886,N_12688);
or U16186 (N_16186,N_13129,N_13453);
nand U16187 (N_16187,N_13020,N_14031);
nor U16188 (N_16188,N_14184,N_13711);
nor U16189 (N_16189,N_15570,N_15779);
nand U16190 (N_16190,N_13638,N_14991);
nor U16191 (N_16191,N_14931,N_15846);
and U16192 (N_16192,N_12206,N_12501);
or U16193 (N_16193,N_13724,N_15221);
xor U16194 (N_16194,N_13647,N_14816);
or U16195 (N_16195,N_13405,N_12879);
and U16196 (N_16196,N_12523,N_15730);
or U16197 (N_16197,N_15769,N_13258);
nor U16198 (N_16198,N_13205,N_15766);
nor U16199 (N_16199,N_15631,N_13475);
nand U16200 (N_16200,N_13613,N_15492);
nor U16201 (N_16201,N_13221,N_13836);
and U16202 (N_16202,N_14569,N_14309);
or U16203 (N_16203,N_14647,N_15782);
nand U16204 (N_16204,N_13691,N_12737);
or U16205 (N_16205,N_12695,N_14669);
nand U16206 (N_16206,N_15363,N_13747);
nor U16207 (N_16207,N_13981,N_13802);
and U16208 (N_16208,N_13459,N_13629);
or U16209 (N_16209,N_13425,N_13428);
nor U16210 (N_16210,N_15806,N_14108);
nor U16211 (N_16211,N_15644,N_14536);
nand U16212 (N_16212,N_12542,N_13199);
nor U16213 (N_16213,N_14415,N_12102);
nand U16214 (N_16214,N_14296,N_14681);
or U16215 (N_16215,N_14662,N_13333);
nor U16216 (N_16216,N_14359,N_13535);
or U16217 (N_16217,N_15993,N_13553);
and U16218 (N_16218,N_14409,N_15068);
nor U16219 (N_16219,N_13193,N_12571);
and U16220 (N_16220,N_14360,N_15270);
nand U16221 (N_16221,N_14116,N_15949);
and U16222 (N_16222,N_14648,N_15114);
and U16223 (N_16223,N_13938,N_13577);
and U16224 (N_16224,N_12662,N_15454);
nor U16225 (N_16225,N_14344,N_13120);
or U16226 (N_16226,N_14552,N_15920);
and U16227 (N_16227,N_15532,N_12961);
and U16228 (N_16228,N_12377,N_12564);
nand U16229 (N_16229,N_15674,N_15341);
nand U16230 (N_16230,N_15187,N_12279);
and U16231 (N_16231,N_15908,N_15616);
and U16232 (N_16232,N_15880,N_15719);
or U16233 (N_16233,N_12621,N_15036);
and U16234 (N_16234,N_15487,N_12332);
nor U16235 (N_16235,N_13247,N_13858);
or U16236 (N_16236,N_13369,N_13521);
nor U16237 (N_16237,N_12522,N_15347);
or U16238 (N_16238,N_12420,N_13246);
nand U16239 (N_16239,N_15247,N_14886);
nor U16240 (N_16240,N_14883,N_12819);
and U16241 (N_16241,N_13293,N_14014);
nand U16242 (N_16242,N_12561,N_13144);
and U16243 (N_16243,N_13291,N_13372);
xor U16244 (N_16244,N_13353,N_13117);
nand U16245 (N_16245,N_14372,N_12524);
nand U16246 (N_16246,N_12984,N_15979);
nand U16247 (N_16247,N_13740,N_15060);
or U16248 (N_16248,N_14670,N_12757);
or U16249 (N_16249,N_15225,N_15188);
and U16250 (N_16250,N_12699,N_15186);
xor U16251 (N_16251,N_14243,N_13106);
or U16252 (N_16252,N_13508,N_15070);
and U16253 (N_16253,N_13430,N_13565);
nor U16254 (N_16254,N_14003,N_12177);
and U16255 (N_16255,N_13335,N_12226);
and U16256 (N_16256,N_14231,N_15439);
and U16257 (N_16257,N_14480,N_15268);
and U16258 (N_16258,N_13678,N_14948);
nand U16259 (N_16259,N_14485,N_13816);
and U16260 (N_16260,N_14760,N_15019);
nand U16261 (N_16261,N_15312,N_12526);
nor U16262 (N_16262,N_14665,N_13337);
nor U16263 (N_16263,N_13953,N_12442);
or U16264 (N_16264,N_14093,N_12677);
and U16265 (N_16265,N_12632,N_15748);
nand U16266 (N_16266,N_12684,N_14934);
and U16267 (N_16267,N_15912,N_13204);
and U16268 (N_16268,N_12282,N_12854);
nand U16269 (N_16269,N_14176,N_12032);
or U16270 (N_16270,N_14702,N_14479);
nand U16271 (N_16271,N_15181,N_14298);
xor U16272 (N_16272,N_14307,N_13912);
and U16273 (N_16273,N_15981,N_14058);
or U16274 (N_16274,N_14627,N_14493);
and U16275 (N_16275,N_15923,N_13976);
nor U16276 (N_16276,N_14498,N_15242);
nor U16277 (N_16277,N_13950,N_15185);
and U16278 (N_16278,N_12560,N_13913);
and U16279 (N_16279,N_15530,N_13679);
nor U16280 (N_16280,N_14585,N_14005);
and U16281 (N_16281,N_12924,N_15733);
and U16282 (N_16282,N_13773,N_14789);
nand U16283 (N_16283,N_12969,N_13095);
nand U16284 (N_16284,N_14097,N_13124);
nor U16285 (N_16285,N_15639,N_15699);
or U16286 (N_16286,N_12000,N_12094);
or U16287 (N_16287,N_15438,N_14322);
and U16288 (N_16288,N_15263,N_15493);
and U16289 (N_16289,N_13656,N_14297);
or U16290 (N_16290,N_14273,N_13759);
and U16291 (N_16291,N_14025,N_14328);
or U16292 (N_16292,N_15927,N_13519);
nor U16293 (N_16293,N_13482,N_13017);
or U16294 (N_16294,N_14355,N_15311);
nand U16295 (N_16295,N_13356,N_15707);
nand U16296 (N_16296,N_12869,N_14683);
nand U16297 (N_16297,N_12685,N_15589);
xnor U16298 (N_16298,N_14047,N_15802);
nor U16299 (N_16299,N_14749,N_15789);
or U16300 (N_16300,N_13635,N_15314);
nor U16301 (N_16301,N_14299,N_12762);
xnor U16302 (N_16302,N_15891,N_12514);
nand U16303 (N_16303,N_13188,N_12059);
or U16304 (N_16304,N_12559,N_13007);
nand U16305 (N_16305,N_13699,N_12370);
nand U16306 (N_16306,N_13315,N_13927);
nor U16307 (N_16307,N_13835,N_12224);
nor U16308 (N_16308,N_15860,N_15618);
and U16309 (N_16309,N_15576,N_12184);
and U16310 (N_16310,N_15702,N_14286);
nor U16311 (N_16311,N_12063,N_15645);
xor U16312 (N_16312,N_13654,N_13354);
or U16313 (N_16313,N_14261,N_15841);
and U16314 (N_16314,N_13223,N_13341);
nand U16315 (N_16315,N_15889,N_13863);
nor U16316 (N_16316,N_13715,N_13686);
and U16317 (N_16317,N_12775,N_12554);
xor U16318 (N_16318,N_15429,N_15456);
and U16319 (N_16319,N_14581,N_12529);
nand U16320 (N_16320,N_15890,N_13931);
nor U16321 (N_16321,N_13528,N_12747);
or U16322 (N_16322,N_15204,N_13593);
or U16323 (N_16323,N_12021,N_14263);
nand U16324 (N_16324,N_12929,N_14507);
and U16325 (N_16325,N_14330,N_13263);
and U16326 (N_16326,N_13837,N_13227);
or U16327 (N_16327,N_14813,N_15524);
nand U16328 (N_16328,N_13320,N_14537);
nand U16329 (N_16329,N_13270,N_14082);
nor U16330 (N_16330,N_14086,N_15413);
and U16331 (N_16331,N_13969,N_13476);
and U16332 (N_16332,N_12809,N_12649);
or U16333 (N_16333,N_12758,N_15184);
and U16334 (N_16334,N_14505,N_12053);
or U16335 (N_16335,N_14197,N_13624);
nand U16336 (N_16336,N_13708,N_13026);
and U16337 (N_16337,N_15328,N_12421);
nor U16338 (N_16338,N_14430,N_12237);
nor U16339 (N_16339,N_12623,N_12367);
or U16340 (N_16340,N_15334,N_13610);
nand U16341 (N_16341,N_14371,N_15325);
or U16342 (N_16342,N_14265,N_13817);
nor U16343 (N_16343,N_12384,N_15683);
and U16344 (N_16344,N_12166,N_14658);
or U16345 (N_16345,N_14785,N_12103);
or U16346 (N_16346,N_15164,N_13714);
and U16347 (N_16347,N_13721,N_13999);
nand U16348 (N_16348,N_14640,N_15412);
nor U16349 (N_16349,N_14280,N_13420);
and U16350 (N_16350,N_12701,N_14902);
nand U16351 (N_16351,N_12616,N_13006);
nand U16352 (N_16352,N_15108,N_14346);
or U16353 (N_16353,N_12648,N_13549);
and U16354 (N_16354,N_13061,N_12212);
nor U16355 (N_16355,N_14753,N_15675);
and U16356 (N_16356,N_12689,N_15659);
nor U16357 (N_16357,N_14316,N_15765);
and U16358 (N_16358,N_15673,N_15717);
and U16359 (N_16359,N_12870,N_14763);
nand U16360 (N_16360,N_15275,N_12238);
nor U16361 (N_16361,N_13398,N_13075);
nor U16362 (N_16362,N_12067,N_15020);
nor U16363 (N_16363,N_13384,N_15110);
nand U16364 (N_16364,N_12995,N_15159);
nor U16365 (N_16365,N_13575,N_15158);
nor U16366 (N_16366,N_12749,N_15442);
nor U16367 (N_16367,N_15472,N_12139);
and U16368 (N_16368,N_13281,N_12672);
nand U16369 (N_16369,N_13556,N_12376);
nor U16370 (N_16370,N_12170,N_15813);
or U16371 (N_16371,N_14135,N_14237);
and U16372 (N_16372,N_12419,N_13534);
nand U16373 (N_16373,N_12256,N_14671);
or U16374 (N_16374,N_14053,N_12810);
nor U16375 (N_16375,N_13147,N_13469);
nor U16376 (N_16376,N_13445,N_15691);
nand U16377 (N_16377,N_14724,N_15000);
nand U16378 (N_16378,N_13820,N_12904);
or U16379 (N_16379,N_13040,N_15437);
nor U16380 (N_16380,N_14656,N_15179);
nor U16381 (N_16381,N_15823,N_14946);
and U16382 (N_16382,N_12161,N_12897);
nand U16383 (N_16383,N_14465,N_12779);
and U16384 (N_16384,N_13967,N_12704);
xor U16385 (N_16385,N_14209,N_13584);
nand U16386 (N_16386,N_14922,N_14534);
or U16387 (N_16387,N_13848,N_15826);
nor U16388 (N_16388,N_15445,N_13499);
nor U16389 (N_16389,N_15686,N_12940);
and U16390 (N_16390,N_15049,N_15505);
nor U16391 (N_16391,N_12078,N_13437);
or U16392 (N_16392,N_12952,N_12152);
xor U16393 (N_16393,N_12654,N_15136);
or U16394 (N_16394,N_13809,N_14139);
or U16395 (N_16395,N_13352,N_15149);
or U16396 (N_16396,N_14750,N_15950);
nand U16397 (N_16397,N_14348,N_15271);
and U16398 (N_16398,N_15004,N_14358);
and U16399 (N_16399,N_12499,N_15461);
and U16400 (N_16400,N_13460,N_12334);
nor U16401 (N_16401,N_12763,N_13330);
or U16402 (N_16402,N_15937,N_14202);
nor U16403 (N_16403,N_15391,N_14075);
or U16404 (N_16404,N_13093,N_12245);
or U16405 (N_16405,N_13801,N_12800);
nand U16406 (N_16406,N_13728,N_15286);
and U16407 (N_16407,N_12733,N_15135);
and U16408 (N_16408,N_15431,N_15152);
xor U16409 (N_16409,N_14978,N_15193);
and U16410 (N_16410,N_13178,N_12035);
or U16411 (N_16411,N_14970,N_14950);
or U16412 (N_16412,N_12100,N_12799);
nand U16413 (N_16413,N_14726,N_12277);
nand U16414 (N_16414,N_15997,N_15455);
nand U16415 (N_16415,N_15300,N_15763);
and U16416 (N_16416,N_12795,N_15214);
or U16417 (N_16417,N_12798,N_15738);
and U16418 (N_16418,N_13932,N_14213);
nor U16419 (N_16419,N_15291,N_12169);
nand U16420 (N_16420,N_14694,N_14365);
and U16421 (N_16421,N_15246,N_13265);
and U16422 (N_16422,N_14893,N_15285);
nor U16423 (N_16423,N_14979,N_12828);
xor U16424 (N_16424,N_14843,N_14557);
and U16425 (N_16425,N_12325,N_13760);
nand U16426 (N_16426,N_12635,N_12963);
and U16427 (N_16427,N_12475,N_15388);
xnor U16428 (N_16428,N_12127,N_12764);
or U16429 (N_16429,N_14821,N_15590);
nand U16430 (N_16430,N_12473,N_14682);
or U16431 (N_16431,N_15088,N_14182);
or U16432 (N_16432,N_14103,N_12942);
and U16433 (N_16433,N_15180,N_14802);
and U16434 (N_16434,N_15901,N_12885);
nand U16435 (N_16435,N_13432,N_12744);
nor U16436 (N_16436,N_12941,N_13443);
or U16437 (N_16437,N_14740,N_15239);
and U16438 (N_16438,N_12108,N_13653);
nand U16439 (N_16439,N_14306,N_15948);
and U16440 (N_16440,N_15172,N_12508);
nand U16441 (N_16441,N_14577,N_13166);
and U16442 (N_16442,N_13331,N_12136);
nand U16443 (N_16443,N_13637,N_13940);
nand U16444 (N_16444,N_14573,N_14188);
or U16445 (N_16445,N_13392,N_15966);
and U16446 (N_16446,N_12853,N_12953);
nor U16447 (N_16447,N_14684,N_15653);
nand U16448 (N_16448,N_14375,N_12676);
nor U16449 (N_16449,N_15139,N_12653);
nand U16450 (N_16450,N_14008,N_14641);
nand U16451 (N_16451,N_14452,N_13206);
nor U16452 (N_16452,N_13674,N_12670);
or U16453 (N_16453,N_14904,N_15168);
and U16454 (N_16454,N_13833,N_14965);
nand U16455 (N_16455,N_13419,N_15670);
or U16456 (N_16456,N_15091,N_13483);
or U16457 (N_16457,N_13968,N_15174);
and U16458 (N_16458,N_13264,N_15503);
and U16459 (N_16459,N_13273,N_14414);
nand U16460 (N_16460,N_15190,N_13743);
or U16461 (N_16461,N_14205,N_14876);
and U16462 (N_16462,N_15061,N_12336);
and U16463 (N_16463,N_14249,N_14410);
or U16464 (N_16464,N_14856,N_13665);
and U16465 (N_16465,N_13029,N_12064);
or U16466 (N_16466,N_15924,N_12415);
nor U16467 (N_16467,N_13639,N_13342);
and U16468 (N_16468,N_14107,N_12802);
and U16469 (N_16469,N_15382,N_15358);
nor U16470 (N_16470,N_14809,N_13503);
nand U16471 (N_16471,N_15352,N_13628);
or U16472 (N_16472,N_14898,N_12117);
and U16473 (N_16473,N_13719,N_14874);
and U16474 (N_16474,N_12933,N_14578);
nand U16475 (N_16475,N_15057,N_15641);
or U16476 (N_16476,N_13859,N_12846);
nand U16477 (N_16477,N_14077,N_14010);
nand U16478 (N_16478,N_12129,N_12069);
or U16479 (N_16479,N_13463,N_12692);
nand U16480 (N_16480,N_13804,N_14827);
nand U16481 (N_16481,N_14609,N_14619);
or U16482 (N_16482,N_15385,N_12551);
and U16483 (N_16483,N_12845,N_15360);
nand U16484 (N_16484,N_14437,N_14649);
or U16485 (N_16485,N_12902,N_13649);
nor U16486 (N_16486,N_15626,N_12463);
nor U16487 (N_16487,N_14007,N_13794);
and U16488 (N_16488,N_15793,N_12435);
nor U16489 (N_16489,N_12449,N_13754);
nand U16490 (N_16490,N_15280,N_13911);
or U16491 (N_16491,N_15430,N_12088);
or U16492 (N_16492,N_13164,N_14861);
or U16493 (N_16493,N_14203,N_14799);
or U16494 (N_16494,N_14907,N_15457);
nor U16495 (N_16495,N_14598,N_14383);
nand U16496 (N_16496,N_14133,N_13571);
or U16497 (N_16497,N_14685,N_15191);
and U16498 (N_16498,N_14894,N_12453);
or U16499 (N_16499,N_12099,N_12270);
and U16500 (N_16500,N_15038,N_12986);
and U16501 (N_16501,N_14379,N_14975);
nand U16502 (N_16502,N_15402,N_14779);
and U16503 (N_16503,N_14814,N_15728);
and U16504 (N_16504,N_12663,N_13176);
and U16505 (N_16505,N_15578,N_15684);
nor U16506 (N_16506,N_14944,N_14969);
nand U16507 (N_16507,N_12706,N_15753);
or U16508 (N_16508,N_12811,N_12271);
nand U16509 (N_16509,N_12834,N_14746);
and U16510 (N_16510,N_15432,N_14698);
or U16511 (N_16511,N_12007,N_14903);
nand U16512 (N_16512,N_13594,N_15523);
and U16513 (N_16513,N_14622,N_14490);
nor U16514 (N_16514,N_13321,N_13324);
or U16515 (N_16515,N_15251,N_14548);
or U16516 (N_16516,N_12107,N_14326);
xor U16517 (N_16517,N_14439,N_15971);
nor U16518 (N_16518,N_12725,N_15446);
and U16519 (N_16519,N_14558,N_15667);
or U16520 (N_16520,N_15031,N_13408);
or U16521 (N_16521,N_15032,N_14801);
and U16522 (N_16522,N_12065,N_12817);
nor U16523 (N_16523,N_15810,N_14070);
or U16524 (N_16524,N_12246,N_15306);
and U16525 (N_16525,N_13231,N_15633);
or U16526 (N_16526,N_14501,N_12071);
or U16527 (N_16527,N_15596,N_13634);
nor U16528 (N_16528,N_15016,N_12431);
and U16529 (N_16529,N_14250,N_15762);
nand U16530 (N_16530,N_14545,N_15772);
nor U16531 (N_16531,N_12371,N_14590);
nor U16532 (N_16532,N_14402,N_14187);
or U16533 (N_16533,N_13480,N_15621);
or U16534 (N_16534,N_14055,N_12618);
nor U16535 (N_16535,N_13668,N_15332);
or U16536 (N_16536,N_14608,N_13071);
nand U16537 (N_16537,N_15254,N_15868);
and U16538 (N_16538,N_15976,N_14959);
or U16539 (N_16539,N_15842,N_12801);
nand U16540 (N_16540,N_14419,N_14720);
nand U16541 (N_16541,N_13956,N_14864);
nor U16542 (N_16542,N_13734,N_13815);
nand U16543 (N_16543,N_15452,N_15063);
and U16544 (N_16544,N_15267,N_12893);
or U16545 (N_16545,N_14179,N_15426);
or U16546 (N_16546,N_12824,N_12018);
or U16547 (N_16547,N_13015,N_15575);
nor U16548 (N_16548,N_15893,N_14434);
and U16549 (N_16549,N_14770,N_14420);
nand U16550 (N_16550,N_15021,N_15296);
nand U16551 (N_16551,N_13592,N_12114);
and U16552 (N_16552,N_12607,N_13452);
or U16553 (N_16553,N_15371,N_12489);
or U16554 (N_16554,N_15758,N_13716);
nand U16555 (N_16555,N_14560,N_13195);
nand U16556 (N_16556,N_14895,N_12313);
and U16557 (N_16557,N_13758,N_15625);
and U16558 (N_16558,N_13598,N_13083);
nand U16559 (N_16559,N_12335,N_13538);
and U16560 (N_16560,N_15284,N_12464);
or U16561 (N_16561,N_14110,N_14730);
and U16562 (N_16562,N_15511,N_12787);
nor U16563 (N_16563,N_13244,N_13466);
or U16564 (N_16564,N_15515,N_14691);
nand U16565 (N_16565,N_12661,N_14983);
or U16566 (N_16566,N_12050,N_14474);
and U16567 (N_16567,N_15984,N_14041);
and U16568 (N_16568,N_12298,N_12700);
and U16569 (N_16569,N_13856,N_15721);
or U16570 (N_16570,N_12447,N_15977);
nor U16571 (N_16571,N_15297,N_15752);
nand U16572 (N_16572,N_12383,N_12964);
nor U16573 (N_16573,N_12609,N_13218);
and U16574 (N_16574,N_13085,N_15957);
and U16575 (N_16575,N_14285,N_15862);
and U16576 (N_16576,N_13215,N_13013);
and U16577 (N_16577,N_14777,N_13749);
nor U16578 (N_16578,N_14572,N_13383);
nand U16579 (N_16579,N_12919,N_12066);
xnor U16580 (N_16580,N_13864,N_14354);
or U16581 (N_16581,N_14074,N_15065);
nand U16582 (N_16582,N_12149,N_14389);
nand U16583 (N_16583,N_12275,N_13079);
or U16584 (N_16584,N_15780,N_15076);
or U16585 (N_16585,N_14618,N_13150);
nand U16586 (N_16586,N_15342,N_14741);
nor U16587 (N_16587,N_12214,N_14636);
nor U16588 (N_16588,N_15988,N_13461);
and U16589 (N_16589,N_13312,N_14567);
or U16590 (N_16590,N_12300,N_15003);
and U16591 (N_16591,N_13418,N_13709);
and U16592 (N_16592,N_15026,N_13143);
nand U16593 (N_16593,N_14049,N_14896);
or U16594 (N_16594,N_12829,N_14130);
nand U16595 (N_16595,N_15704,N_13245);
or U16596 (N_16596,N_13292,N_13290);
or U16597 (N_16597,N_12721,N_12868);
and U16598 (N_16598,N_14899,N_15171);
or U16599 (N_16599,N_14678,N_13135);
or U16600 (N_16600,N_12013,N_12822);
or U16601 (N_16601,N_13044,N_14143);
xnor U16602 (N_16602,N_13803,N_13284);
nor U16603 (N_16603,N_14247,N_13200);
nand U16604 (N_16604,N_15499,N_12052);
nand U16605 (N_16605,N_13027,N_14674);
and U16606 (N_16606,N_15117,N_13226);
nor U16607 (N_16607,N_13788,N_13663);
nand U16608 (N_16608,N_14295,N_14398);
nand U16609 (N_16609,N_15873,N_15899);
or U16610 (N_16610,N_14728,N_12789);
nor U16611 (N_16611,N_14759,N_14659);
and U16612 (N_16612,N_15195,N_12433);
nor U16613 (N_16613,N_12405,N_13415);
or U16614 (N_16614,N_15882,N_13849);
nand U16615 (N_16615,N_14458,N_15736);
nor U16616 (N_16616,N_12655,N_12046);
nor U16617 (N_16617,N_14891,N_14955);
nor U16618 (N_16618,N_13374,N_12418);
nor U16619 (N_16619,N_12250,N_14244);
and U16620 (N_16620,N_13214,N_13025);
xor U16621 (N_16621,N_13267,N_14772);
or U16622 (N_16622,N_12973,N_14522);
or U16623 (N_16623,N_15333,N_12323);
nor U16624 (N_16624,N_13370,N_12971);
and U16625 (N_16625,N_12417,N_13666);
and U16626 (N_16626,N_15282,N_14024);
nand U16627 (N_16627,N_14138,N_14442);
nor U16628 (N_16628,N_14100,N_14214);
nor U16629 (N_16629,N_15408,N_12084);
nand U16630 (N_16630,N_14272,N_15474);
or U16631 (N_16631,N_14373,N_15601);
nand U16632 (N_16632,N_12402,N_14386);
or U16633 (N_16633,N_14774,N_12544);
or U16634 (N_16634,N_13736,N_15774);
nor U16635 (N_16635,N_14048,N_15999);
nor U16636 (N_16636,N_15047,N_13043);
or U16637 (N_16637,N_15367,N_13310);
nand U16638 (N_16638,N_14405,N_14207);
nand U16639 (N_16639,N_13692,N_14820);
nand U16640 (N_16640,N_14081,N_12160);
nand U16641 (N_16641,N_13478,N_12049);
nor U16642 (N_16642,N_12610,N_15690);
and U16643 (N_16643,N_12816,N_15294);
nand U16644 (N_16644,N_15776,N_12947);
and U16645 (N_16645,N_14850,N_14797);
and U16646 (N_16646,N_12341,N_13225);
and U16647 (N_16647,N_15343,N_13644);
nor U16648 (N_16648,N_13671,N_13107);
nand U16649 (N_16649,N_15033,N_13298);
or U16650 (N_16650,N_13920,N_15958);
and U16651 (N_16651,N_12283,N_12876);
and U16652 (N_16652,N_12456,N_14704);
or U16653 (N_16653,N_14120,N_13101);
or U16654 (N_16654,N_13717,N_15156);
and U16655 (N_16655,N_13783,N_15613);
nand U16656 (N_16656,N_15606,N_14612);
nand U16657 (N_16657,N_13518,N_13212);
nand U16658 (N_16658,N_12539,N_12573);
nand U16659 (N_16659,N_15796,N_15583);
nor U16660 (N_16660,N_12444,N_12727);
and U16661 (N_16661,N_14961,N_14229);
or U16662 (N_16662,N_12865,N_13220);
nand U16663 (N_16663,N_14170,N_14026);
or U16664 (N_16664,N_14554,N_14909);
nor U16665 (N_16665,N_14758,N_15599);
nor U16666 (N_16666,N_14302,N_14712);
nor U16667 (N_16667,N_12303,N_14584);
nor U16668 (N_16668,N_13972,N_13037);
nand U16669 (N_16669,N_13232,N_12254);
nand U16670 (N_16670,N_12243,N_14004);
and U16671 (N_16671,N_14888,N_13822);
or U16672 (N_16672,N_12937,N_15906);
nor U16673 (N_16673,N_14429,N_13277);
nand U16674 (N_16674,N_15278,N_14981);
nor U16675 (N_16675,N_12192,N_15828);
nor U16676 (N_16676,N_14251,N_14064);
and U16677 (N_16677,N_13540,N_14798);
and U16678 (N_16678,N_15249,N_12625);
nand U16679 (N_16679,N_13066,N_12498);
nand U16680 (N_16680,N_13844,N_12994);
or U16681 (N_16681,N_13344,N_13067);
and U16682 (N_16682,N_12263,N_13276);
nand U16683 (N_16683,N_13781,N_14256);
nand U16684 (N_16684,N_15986,N_12321);
and U16685 (N_16685,N_14363,N_15410);
or U16686 (N_16686,N_13800,N_12958);
and U16687 (N_16687,N_14954,N_12638);
and U16688 (N_16688,N_15201,N_14958);
nand U16689 (N_16689,N_12095,N_15340);
nand U16690 (N_16690,N_12619,N_13830);
or U16691 (N_16691,N_13541,N_14599);
nand U16692 (N_16692,N_13018,N_14884);
nand U16693 (N_16693,N_13902,N_13793);
or U16694 (N_16694,N_14510,N_12201);
and U16695 (N_16695,N_15375,N_13658);
nand U16696 (N_16696,N_12944,N_15428);
or U16697 (N_16697,N_15725,N_12593);
nand U16698 (N_16698,N_14688,N_13530);
nand U16699 (N_16699,N_13752,N_12122);
nor U16700 (N_16700,N_13520,N_12116);
nand U16701 (N_16701,N_15520,N_12374);
and U16702 (N_16702,N_13269,N_13417);
nand U16703 (N_16703,N_14854,N_15029);
or U16704 (N_16704,N_14009,N_12495);
nand U16705 (N_16705,N_15825,N_13899);
nand U16706 (N_16706,N_13945,N_15276);
or U16707 (N_16707,N_14551,N_12352);
nor U16708 (N_16708,N_15533,N_13399);
nand U16709 (N_16709,N_14129,N_15506);
or U16710 (N_16710,N_14988,N_15157);
and U16711 (N_16711,N_14823,N_15116);
xor U16712 (N_16712,N_12249,N_14427);
nor U16713 (N_16713,N_12395,N_13527);
nand U16714 (N_16714,N_14892,N_12213);
nand U16715 (N_16715,N_14664,N_12074);
nand U16716 (N_16716,N_13272,N_15962);
nand U16717 (N_16717,N_15462,N_15521);
and U16718 (N_16718,N_12024,N_15559);
or U16719 (N_16719,N_14644,N_12898);
or U16720 (N_16720,N_12004,N_15468);
nand U16721 (N_16721,N_12549,N_12368);
and U16722 (N_16722,N_12825,N_13707);
or U16723 (N_16723,N_12111,N_15315);
nand U16724 (N_16724,N_13389,N_15087);
nor U16725 (N_16725,N_12043,N_14195);
or U16726 (N_16726,N_13705,N_14680);
nor U16727 (N_16727,N_15940,N_13487);
and U16728 (N_16728,N_14521,N_12862);
and U16729 (N_16729,N_15006,N_14932);
nand U16730 (N_16730,N_12115,N_14952);
nor U16731 (N_16731,N_15534,N_14872);
or U16732 (N_16732,N_14889,N_14162);
or U16733 (N_16733,N_12466,N_14735);
nor U16734 (N_16734,N_12259,N_14303);
and U16735 (N_16735,N_12833,N_15519);
or U16736 (N_16736,N_15355,N_13468);
nand U16737 (N_16737,N_12966,N_12164);
or U16738 (N_16738,N_14222,N_13700);
nor U16739 (N_16739,N_13287,N_12181);
and U16740 (N_16740,N_14424,N_14951);
nor U16741 (N_16741,N_15611,N_13742);
or U16742 (N_16742,N_12041,N_13318);
nand U16743 (N_16743,N_14686,N_13616);
and U16744 (N_16744,N_12207,N_15987);
and U16745 (N_16745,N_12991,N_14492);
and U16746 (N_16746,N_15552,N_13201);
or U16747 (N_16747,N_15553,N_12297);
xnor U16748 (N_16748,N_12253,N_15302);
nor U16749 (N_16749,N_13359,N_12656);
nor U16750 (N_16750,N_15272,N_15549);
or U16751 (N_16751,N_14441,N_13386);
nor U16752 (N_16752,N_12036,N_15477);
or U16753 (N_16753,N_12037,N_13357);
nand U16754 (N_16754,N_14155,N_13818);
nand U16755 (N_16755,N_14340,N_14653);
or U16756 (N_16756,N_15607,N_12460);
nand U16757 (N_16757,N_14915,N_12770);
nor U16758 (N_16758,N_15749,N_12532);
and U16759 (N_16759,N_12471,N_14956);
and U16760 (N_16760,N_13456,N_13326);
or U16761 (N_16761,N_14982,N_13738);
and U16762 (N_16762,N_12227,N_15304);
or U16763 (N_16763,N_13396,N_12353);
nor U16764 (N_16764,N_14606,N_15814);
and U16765 (N_16765,N_15942,N_13696);
nor U16766 (N_16766,N_13609,N_14087);
and U16767 (N_16767,N_15210,N_14701);
nor U16768 (N_16768,N_13102,N_14484);
nand U16769 (N_16769,N_15615,N_13114);
or U16770 (N_16770,N_14628,N_12012);
nand U16771 (N_16771,N_13532,N_13777);
or U16772 (N_16772,N_14736,N_14715);
nand U16773 (N_16773,N_14457,N_12232);
nor U16774 (N_16774,N_13564,N_15262);
nand U16775 (N_16775,N_15319,N_13891);
nor U16776 (N_16776,N_15344,N_12922);
xor U16777 (N_16777,N_12807,N_14977);
nand U16778 (N_16778,N_13966,N_12448);
nor U16779 (N_16779,N_14583,N_14142);
xnor U16780 (N_16780,N_15107,N_13467);
or U16781 (N_16781,N_12803,N_15952);
nor U16782 (N_16782,N_14836,N_14343);
or U16783 (N_16783,N_15554,N_15102);
and U16784 (N_16784,N_14057,N_13224);
or U16785 (N_16785,N_14245,N_13271);
and U16786 (N_16786,N_14756,N_14742);
and U16787 (N_16787,N_13379,N_13906);
nand U16788 (N_16788,N_15137,N_12643);
nand U16789 (N_16789,N_13099,N_13088);
and U16790 (N_16790,N_15679,N_15919);
nand U16791 (N_16791,N_12096,N_15742);
nand U16792 (N_16792,N_15440,N_15488);
and U16793 (N_16793,N_12959,N_14350);
nand U16794 (N_16794,N_15525,N_12880);
nor U16795 (N_16795,N_13765,N_15558);
nor U16796 (N_16796,N_14242,N_15933);
and U16797 (N_16797,N_13104,N_12135);
nor U16798 (N_16798,N_12724,N_14266);
nand U16799 (N_16799,N_12899,N_13157);
nand U16800 (N_16800,N_13151,N_14564);
and U16801 (N_16801,N_12429,N_14716);
nor U16802 (N_16802,N_13567,N_13180);
nand U16803 (N_16803,N_13047,N_14211);
nor U16804 (N_16804,N_14528,N_12552);
and U16805 (N_16805,N_15080,N_13600);
and U16806 (N_16806,N_13559,N_13316);
or U16807 (N_16807,N_15764,N_13672);
or U16808 (N_16808,N_14575,N_12239);
nor U16809 (N_16809,N_12345,N_12118);
and U16810 (N_16810,N_13853,N_12458);
and U16811 (N_16811,N_13362,N_15401);
nor U16812 (N_16812,N_13084,N_12753);
nand U16813 (N_16813,N_12346,N_15829);
and U16814 (N_16814,N_12832,N_12993);
and U16815 (N_16815,N_13823,N_12761);
nand U16816 (N_16816,N_14571,N_12956);
nor U16817 (N_16817,N_14210,N_15123);
and U16818 (N_16818,N_14290,N_14910);
and U16819 (N_16819,N_15913,N_14947);
nor U16820 (N_16820,N_12153,N_15627);
nor U16821 (N_16821,N_12615,N_12373);
xnor U16822 (N_16822,N_15161,N_13116);
nand U16823 (N_16823,N_12180,N_12767);
and U16824 (N_16824,N_14062,N_13579);
and U16825 (N_16825,N_12586,N_12780);
and U16826 (N_16826,N_13733,N_13323);
or U16827 (N_16827,N_12791,N_14270);
nand U16828 (N_16828,N_13588,N_13489);
and U16829 (N_16829,N_15729,N_14967);
nor U16830 (N_16830,N_14173,N_14175);
nand U16831 (N_16831,N_15099,N_14502);
nand U16832 (N_16832,N_15351,N_13000);
nor U16833 (N_16833,N_15642,N_14390);
nor U16834 (N_16834,N_12023,N_12852);
and U16835 (N_16835,N_15111,N_14815);
nand U16836 (N_16836,N_13845,N_12076);
and U16837 (N_16837,N_15732,N_14114);
and U16838 (N_16838,N_13560,N_13137);
or U16839 (N_16839,N_14002,N_14030);
nor U16840 (N_16840,N_15305,N_12576);
or U16841 (N_16841,N_12359,N_15811);
or U16842 (N_16842,N_13512,N_13547);
nand U16843 (N_16843,N_12483,N_15266);
nor U16844 (N_16844,N_15666,N_13611);
nor U16845 (N_16845,N_15709,N_13806);
and U16846 (N_16846,N_15216,N_14258);
and U16847 (N_16847,N_14865,N_13053);
and U16848 (N_16848,N_12740,N_14151);
and U16849 (N_16849,N_13746,N_15230);
nand U16850 (N_16850,N_14123,N_13905);
and U16851 (N_16851,N_12821,N_15059);
and U16852 (N_16852,N_15236,N_15743);
nor U16853 (N_16853,N_12204,N_15478);
nand U16854 (N_16854,N_15922,N_13048);
or U16855 (N_16855,N_14645,N_12252);
or U16856 (N_16856,N_13138,N_12830);
or U16857 (N_16857,N_15292,N_14706);
or U16858 (N_16858,N_13327,N_12911);
nand U16859 (N_16859,N_12748,N_15147);
nor U16860 (N_16860,N_15518,N_12965);
and U16861 (N_16861,N_15539,N_15620);
and U16862 (N_16862,N_15871,N_14453);
or U16863 (N_16863,N_15877,N_12901);
nand U16864 (N_16864,N_15687,N_12109);
nor U16865 (N_16865,N_12404,N_13826);
nand U16866 (N_16866,N_13021,N_12240);
nor U16867 (N_16867,N_13875,N_15548);
nor U16868 (N_16868,N_14125,N_15056);
and U16869 (N_16869,N_13349,N_12209);
and U16870 (N_16870,N_15075,N_13651);
nand U16871 (N_16871,N_12362,N_12734);
and U16872 (N_16872,N_12548,N_13125);
nor U16873 (N_16873,N_12436,N_12851);
nand U16874 (N_16874,N_14527,N_13442);
or U16875 (N_16875,N_13336,N_12412);
or U16876 (N_16876,N_14841,N_14562);
nand U16877 (N_16877,N_14790,N_13992);
and U16878 (N_16878,N_13829,N_12058);
or U16879 (N_16879,N_14807,N_12128);
and U16880 (N_16880,N_15441,N_15617);
or U16881 (N_16881,N_12394,N_15231);
and U16882 (N_16882,N_12774,N_12891);
or U16883 (N_16883,N_13735,N_13041);
or U16884 (N_16884,N_15290,N_13729);
nor U16885 (N_16885,N_12382,N_13073);
and U16886 (N_16886,N_13163,N_12866);
nor U16887 (N_16887,N_12729,N_13471);
nand U16888 (N_16888,N_13766,N_13404);
or U16889 (N_16889,N_14109,N_12276);
nor U16890 (N_16890,N_15289,N_15713);
nand U16891 (N_16891,N_15044,N_15017);
or U16892 (N_16892,N_15288,N_14404);
and U16893 (N_16893,N_14071,N_14960);
and U16894 (N_16894,N_14594,N_13939);
nand U16895 (N_16895,N_13695,N_13155);
and U16896 (N_16896,N_14456,N_12690);
and U16897 (N_16897,N_13843,N_13892);
nand U16898 (N_16898,N_13814,N_13005);
and U16899 (N_16899,N_14043,N_12668);
and U16900 (N_16900,N_14657,N_14767);
nand U16901 (N_16901,N_14052,N_13551);
nor U16902 (N_16902,N_13400,N_14822);
or U16903 (N_16903,N_15887,N_13623);
nor U16904 (N_16904,N_15955,N_15550);
and U16905 (N_16905,N_14337,N_14264);
nor U16906 (N_16906,N_15217,N_14230);
nand U16907 (N_16907,N_15735,N_12999);
nand U16908 (N_16908,N_12189,N_12713);
or U16909 (N_16909,N_15479,N_13454);
nor U16910 (N_16910,N_13145,N_14921);
and U16911 (N_16911,N_15381,N_12921);
nand U16912 (N_16912,N_14771,N_13427);
nor U16913 (N_16913,N_13558,N_15064);
or U16914 (N_16914,N_12597,N_13139);
nand U16915 (N_16915,N_15857,N_15040);
and U16916 (N_16916,N_13942,N_14621);
nor U16917 (N_16917,N_14291,N_12386);
nand U16918 (N_16918,N_13294,N_12717);
nand U16919 (N_16919,N_12439,N_14602);
or U16920 (N_16920,N_15931,N_14515);
nor U16921 (N_16921,N_13440,N_15658);
or U16922 (N_16922,N_12736,N_14487);
nor U16923 (N_16923,N_14859,N_14855);
nand U16924 (N_16924,N_12889,N_15025);
and U16925 (N_16925,N_13394,N_14085);
or U16926 (N_16926,N_13105,N_13894);
nor U16927 (N_16927,N_13406,N_13689);
nor U16928 (N_16928,N_15400,N_14733);
or U16929 (N_16929,N_14556,N_12479);
nand U16930 (N_16930,N_12311,N_14341);
and U16931 (N_16931,N_12746,N_13421);
nand U16932 (N_16932,N_12079,N_14046);
nor U16933 (N_16933,N_13523,N_13824);
nor U16934 (N_16934,N_14136,N_15475);
nor U16935 (N_16935,N_15697,N_14651);
nor U16936 (N_16936,N_15419,N_14974);
nand U16937 (N_16937,N_15349,N_12570);
or U16938 (N_16938,N_13889,N_13008);
or U16939 (N_16939,N_15453,N_15303);
and U16940 (N_16940,N_13984,N_12261);
or U16941 (N_16941,N_13413,N_12159);
and U16942 (N_16942,N_14574,N_12602);
and U16943 (N_16943,N_14113,N_15366);
or U16944 (N_16944,N_15097,N_14076);
nand U16945 (N_16945,N_12306,N_14582);
or U16946 (N_16946,N_13884,N_15574);
nand U16947 (N_16947,N_15037,N_12574);
or U16948 (N_16948,N_12978,N_15622);
or U16949 (N_16949,N_15800,N_12022);
and U16950 (N_16950,N_12708,N_15781);
and U16951 (N_16951,N_14500,N_14376);
nand U16952 (N_16952,N_13841,N_14817);
nand U16953 (N_16953,N_12698,N_13995);
or U16954 (N_16954,N_13768,N_14494);
nor U16955 (N_16955,N_13868,N_14924);
or U16956 (N_16956,N_13186,N_13615);
nor U16957 (N_16957,N_12512,N_14869);
and U16958 (N_16958,N_12356,N_13248);
nor U16959 (N_16959,N_13130,N_15447);
nand U16960 (N_16960,N_15229,N_15320);
or U16961 (N_16961,N_12385,N_13510);
nand U16962 (N_16962,N_14603,N_12857);
nand U16963 (N_16963,N_14906,N_13998);
and U16964 (N_16964,N_15220,N_12090);
nor U16965 (N_16965,N_13031,N_15167);
nor U16966 (N_16966,N_14278,N_14631);
nand U16967 (N_16967,N_12931,N_13569);
nand U16968 (N_16968,N_14421,N_12813);
and U16969 (N_16969,N_15200,N_13959);
or U16970 (N_16970,N_12294,N_15688);
nor U16971 (N_16971,N_14917,N_13300);
nor U16972 (N_16972,N_15692,N_12438);
and U16973 (N_16973,N_15379,N_13343);
nor U16974 (N_16974,N_13183,N_13944);
nand U16975 (N_16975,N_15597,N_12694);
or U16976 (N_16976,N_14793,N_15269);
nor U16977 (N_16977,N_13397,N_13633);
and U16978 (N_16978,N_12572,N_12628);
and U16979 (N_16979,N_14873,N_13473);
and U16980 (N_16980,N_13774,N_12968);
nor U16981 (N_16981,N_15853,N_14095);
nand U16982 (N_16982,N_12950,N_15978);
nor U16983 (N_16983,N_12287,N_14178);
and U16984 (N_16984,N_14559,N_13368);
and U16985 (N_16985,N_12719,N_15205);
and U16986 (N_16986,N_12545,N_14401);
and U16987 (N_16987,N_14863,N_14800);
and U16988 (N_16988,N_12731,N_15907);
and U16989 (N_16989,N_15989,N_15084);
or U16990 (N_16990,N_13797,N_15541);
or U16991 (N_16991,N_12722,N_14639);
nor U16992 (N_16992,N_12020,N_12945);
or U16993 (N_16993,N_13661,N_15182);
nor U16994 (N_16994,N_13601,N_14220);
nor U16995 (N_16995,N_12337,N_14588);
and U16996 (N_16996,N_12550,N_14159);
nand U16997 (N_16997,N_14027,N_12400);
nor U16998 (N_16998,N_13234,N_15415);
and U16999 (N_16999,N_15896,N_14568);
nand U17000 (N_17000,N_13208,N_15875);
or U17001 (N_17001,N_14332,N_14065);
nor U17002 (N_17002,N_15557,N_14305);
nor U17003 (N_17003,N_15387,N_14023);
nor U17004 (N_17004,N_12203,N_13640);
nor U17005 (N_17005,N_15794,N_12617);
and U17006 (N_17006,N_13422,N_12393);
or U17007 (N_17007,N_12510,N_15563);
xor U17008 (N_17008,N_13109,N_15856);
or U17009 (N_17009,N_15859,N_12120);
or U17010 (N_17010,N_15718,N_14646);
nor U17011 (N_17011,N_12806,N_15932);
nand U17012 (N_17012,N_15915,N_15215);
nand U17013 (N_17013,N_13351,N_15819);
and U17014 (N_17014,N_14542,N_12831);
nand U17015 (N_17015,N_13965,N_14079);
or U17016 (N_17016,N_14984,N_14725);
and U17017 (N_17017,N_13065,N_12985);
nand U17018 (N_17018,N_15587,N_15218);
and U17019 (N_17019,N_12289,N_12450);
nor U17020 (N_17020,N_14630,N_14466);
xnor U17021 (N_17021,N_14001,N_12381);
nor U17022 (N_17022,N_14446,N_15339);
nand U17023 (N_17023,N_13210,N_13683);
nor U17024 (N_17024,N_13140,N_14362);
and U17025 (N_17025,N_14201,N_12517);
nand U17026 (N_17026,N_15854,N_15330);
or U17027 (N_17027,N_12567,N_15894);
nor U17028 (N_17028,N_12284,N_12340);
and U17029 (N_17029,N_15788,N_12221);
and U17030 (N_17030,N_14171,N_13243);
or U17031 (N_17031,N_13599,N_13751);
or U17032 (N_17032,N_15798,N_13096);
or U17033 (N_17033,N_15560,N_12556);
nor U17034 (N_17034,N_13737,N_15792);
or U17035 (N_17035,N_15951,N_14164);
nand U17036 (N_17036,N_15546,N_15373);
nand U17037 (N_17037,N_13110,N_13869);
or U17038 (N_17038,N_12142,N_12314);
nand U17039 (N_17039,N_12518,N_12976);
nor U17040 (N_17040,N_13123,N_15947);
nor U17041 (N_17041,N_14993,N_12315);
nor U17042 (N_17042,N_14690,N_13687);
and U17043 (N_17043,N_15581,N_14089);
xor U17044 (N_17044,N_13501,N_13807);
and U17045 (N_17045,N_13257,N_13207);
nand U17046 (N_17046,N_12051,N_12776);
and U17047 (N_17047,N_14315,N_13296);
nand U17048 (N_17048,N_14313,N_13627);
nand U17049 (N_17049,N_13643,N_12110);
nand U17050 (N_17050,N_12946,N_15897);
or U17051 (N_17051,N_15812,N_15629);
and U17052 (N_17052,N_12530,N_15821);
nand U17053 (N_17053,N_12401,N_13791);
or U17054 (N_17054,N_13929,N_12917);
nor U17055 (N_17055,N_14739,N_12849);
nand U17056 (N_17056,N_14748,N_14672);
nand U17057 (N_17057,N_13098,N_12759);
nand U17058 (N_17058,N_13121,N_12457);
nor U17059 (N_17059,N_15124,N_14734);
or U17060 (N_17060,N_14971,N_14460);
or U17061 (N_17061,N_14524,N_12666);
nor U17062 (N_17062,N_15008,N_13046);
and U17063 (N_17063,N_15098,N_13704);
and U17064 (N_17064,N_12205,N_15163);
nand U17065 (N_17065,N_15651,N_14796);
and U17066 (N_17066,N_15416,N_12823);
and U17067 (N_17067,N_14719,N_13632);
nor U17068 (N_17068,N_14858,N_13543);
nand U17069 (N_17069,N_12432,N_14625);
or U17070 (N_17070,N_13772,N_13390);
or U17071 (N_17071,N_14743,N_12962);
or U17072 (N_17072,N_15778,N_13753);
and U17073 (N_17073,N_14826,N_12972);
and U17074 (N_17074,N_14553,N_14327);
nor U17075 (N_17075,N_15767,N_15392);
nand U17076 (N_17076,N_13978,N_12179);
nor U17077 (N_17077,N_15705,N_13602);
nor U17078 (N_17078,N_13669,N_15542);
and U17079 (N_17079,N_14269,N_12936);
or U17080 (N_17080,N_13160,N_12480);
or U17081 (N_17081,N_12075,N_15208);
nor U17082 (N_17082,N_13790,N_12639);
or U17083 (N_17083,N_14468,N_12907);
nand U17084 (N_17084,N_13156,N_13240);
or U17085 (N_17085,N_12251,N_14980);
nor U17086 (N_17086,N_13636,N_15409);
nand U17087 (N_17087,N_13022,N_12455);
nor U17088 (N_17088,N_12413,N_12930);
nor U17089 (N_17089,N_13941,N_15677);
and U17090 (N_17090,N_15106,N_13831);
nor U17091 (N_17091,N_14378,N_15945);
and U17092 (N_17092,N_13328,N_15604);
or U17093 (N_17093,N_12011,N_12585);
and U17094 (N_17094,N_14851,N_12858);
and U17095 (N_17095,N_13346,N_15994);
and U17096 (N_17096,N_15206,N_12319);
or U17097 (N_17097,N_13198,N_13685);
nand U17098 (N_17098,N_14166,N_12687);
nand U17099 (N_17099,N_13904,N_12485);
or U17100 (N_17100,N_13874,N_12555);
and U17101 (N_17101,N_12949,N_12062);
nor U17102 (N_17102,N_15175,N_14679);
and U17103 (N_17103,N_13762,N_14084);
and U17104 (N_17104,N_15741,N_13350);
xnor U17105 (N_17105,N_15376,N_14713);
or U17106 (N_17106,N_14632,N_15313);
and U17107 (N_17107,N_14837,N_12234);
xnor U17108 (N_17108,N_13068,N_14022);
nor U17109 (N_17109,N_13566,N_15133);
and U17110 (N_17110,N_13934,N_12150);
and U17111 (N_17111,N_13865,N_14432);
nand U17112 (N_17112,N_15336,N_15384);
nor U17113 (N_17113,N_15424,N_14517);
and U17114 (N_17114,N_14565,N_12010);
nand U17115 (N_17115,N_14239,N_15203);
nand U17116 (N_17116,N_12476,N_15903);
nor U17117 (N_17117,N_13662,N_15248);
nor U17118 (N_17118,N_14890,N_15720);
nand U17119 (N_17119,N_15417,N_13937);
nand U17120 (N_17120,N_15671,N_15007);
nand U17121 (N_17121,N_13893,N_13798);
or U17122 (N_17122,N_14128,N_15849);
nand U17123 (N_17123,N_12223,N_12106);
and U17124 (N_17124,N_13161,N_12081);
nand U17125 (N_17125,N_13087,N_15397);
nor U17126 (N_17126,N_13582,N_12061);
or U17127 (N_17127,N_13974,N_13769);
or U17128 (N_17128,N_12928,N_15535);
or U17129 (N_17129,N_14477,N_12673);
and U17130 (N_17130,N_12348,N_15731);
nand U17131 (N_17131,N_12123,N_12743);
and U17132 (N_17132,N_13256,N_15610);
and U17133 (N_17133,N_12158,N_13573);
and U17134 (N_17134,N_15308,N_13506);
xnor U17135 (N_17135,N_14868,N_12440);
nand U17136 (N_17136,N_15078,N_14570);
and U17137 (N_17137,N_12765,N_13606);
or U17138 (N_17138,N_14425,N_12543);
and U17139 (N_17139,N_15245,N_12503);
nand U17140 (N_17140,N_14781,N_13792);
or U17141 (N_17141,N_15199,N_13035);
nand U17142 (N_17142,N_12481,N_13249);
and U17143 (N_17143,N_15169,N_12837);
or U17144 (N_17144,N_12546,N_12987);
or U17145 (N_17145,N_15726,N_14905);
nand U17146 (N_17146,N_14871,N_15528);
or U17147 (N_17147,N_13779,N_13821);
and U17148 (N_17148,N_12422,N_12486);
nand U17149 (N_17149,N_13434,N_14766);
nor U17150 (N_17150,N_13141,N_14830);
or U17151 (N_17151,N_13989,N_13289);
nor U17152 (N_17152,N_14949,N_15816);
and U17153 (N_17153,N_12288,N_12407);
and U17154 (N_17154,N_13378,N_15985);
nor U17155 (N_17155,N_13049,N_13295);
and U17156 (N_17156,N_12112,N_15760);
and U17157 (N_17157,N_12630,N_15013);
and U17158 (N_17158,N_13059,N_15791);
nor U17159 (N_17159,N_12025,N_12903);
nor U17160 (N_17160,N_15939,N_12048);
nor U17161 (N_17161,N_12835,N_12682);
nor U17162 (N_17162,N_15569,N_12631);
nand U17163 (N_17163,N_13165,N_12398);
and U17164 (N_17164,N_14194,N_13873);
nor U17165 (N_17165,N_14747,N_15892);
nand U17166 (N_17166,N_13009,N_14803);
nor U17167 (N_17167,N_13371,N_15066);
xnor U17168 (N_17168,N_12777,N_14999);
and U17169 (N_17169,N_15840,N_14281);
nor U17170 (N_17170,N_14828,N_13885);
nor U17171 (N_17171,N_14607,N_14321);
nand U17172 (N_17172,N_14601,N_14248);
nand U17173 (N_17173,N_12304,N_14913);
and U17174 (N_17174,N_13980,N_15131);
xor U17175 (N_17175,N_14000,N_13100);
nor U17176 (N_17176,N_15480,N_15129);
or U17177 (N_17177,N_14538,N_13317);
and U17178 (N_17178,N_13363,N_15310);
nand U17179 (N_17179,N_12665,N_13591);
or U17180 (N_17180,N_15353,N_14642);
and U17181 (N_17181,N_13051,N_15504);
and U17182 (N_17182,N_14226,N_14236);
and U17183 (N_17183,N_15602,N_13380);
nor U17184 (N_17184,N_13439,N_12820);
nand U17185 (N_17185,N_15941,N_13614);
or U17186 (N_17186,N_12174,N_15850);
nor U17187 (N_17187,N_14881,N_15640);
nand U17188 (N_17188,N_15338,N_12087);
or U17189 (N_17189,N_13260,N_12826);
nand U17190 (N_17190,N_12981,N_15142);
and U17191 (N_17191,N_13958,N_13842);
nor U17192 (N_17192,N_12015,N_15197);
or U17193 (N_17193,N_15723,N_12132);
nand U17194 (N_17194,N_12105,N_13955);
and U17195 (N_17195,N_12372,N_12030);
and U17196 (N_17196,N_14476,N_14838);
or U17197 (N_17197,N_12979,N_13827);
nor U17198 (N_17198,N_12477,N_14235);
nor U17199 (N_17199,N_12175,N_13536);
nor U17200 (N_17200,N_12301,N_13305);
nor U17201 (N_17201,N_14127,N_14042);
nand U17202 (N_17202,N_14935,N_14149);
nand U17203 (N_17203,N_15028,N_15209);
or U17204 (N_17204,N_12409,N_13514);
xnor U17205 (N_17205,N_12818,N_12659);
nor U17206 (N_17206,N_14463,N_13286);
or U17207 (N_17207,N_15160,N_15372);
nor U17208 (N_17208,N_14233,N_13361);
nor U17209 (N_17209,N_13112,N_13388);
nand U17210 (N_17210,N_12185,N_14218);
and U17211 (N_17211,N_14792,N_14936);
xnor U17212 (N_17212,N_13778,N_13447);
nor U17213 (N_17213,N_12347,N_14964);
nor U17214 (N_17214,N_15961,N_12255);
nand U17215 (N_17215,N_14412,N_14994);
xnor U17216 (N_17216,N_13119,N_12842);
and U17217 (N_17217,N_14957,N_12989);
nor U17218 (N_17218,N_14782,N_14092);
nand U17219 (N_17219,N_13529,N_12838);
and U17220 (N_17220,N_15295,N_15807);
or U17221 (N_17221,N_14805,N_15746);
nand U17222 (N_17222,N_14867,N_13698);
or U17223 (N_17223,N_14833,N_13115);
and U17224 (N_17224,N_14208,N_13825);
or U17225 (N_17225,N_12140,N_14385);
or U17226 (N_17226,N_15073,N_15154);
and U17227 (N_17227,N_14503,N_15012);
or U17228 (N_17228,N_13345,N_13918);
and U17229 (N_17229,N_13152,N_13216);
or U17230 (N_17230,N_15566,N_13630);
nor U17231 (N_17231,N_13587,N_13548);
or U17232 (N_17232,N_13118,N_13402);
nand U17233 (N_17233,N_14399,N_12507);
and U17234 (N_17234,N_14102,N_15712);
and U17235 (N_17235,N_14317,N_12307);
or U17236 (N_17236,N_15561,N_15600);
and U17237 (N_17237,N_14549,N_15956);
xnor U17238 (N_17238,N_12026,N_15095);
or U17239 (N_17239,N_13784,N_12211);
nor U17240 (N_17240,N_12772,N_12369);
nand U17241 (N_17241,N_14692,N_12141);
and U17242 (N_17242,N_12285,N_15467);
nand U17243 (N_17243,N_14012,N_13340);
and U17244 (N_17244,N_14526,N_14156);
and U17245 (N_17245,N_14267,N_13542);
nand U17246 (N_17246,N_14914,N_13574);
or U17247 (N_17247,N_14930,N_12146);
or U17248 (N_17248,N_12344,N_12850);
nand U17249 (N_17249,N_15698,N_12229);
nand U17250 (N_17250,N_15580,N_13202);
or U17251 (N_17251,N_15567,N_15243);
or U17252 (N_17252,N_12101,N_14495);
or U17253 (N_17253,N_12077,N_13280);
or U17254 (N_17254,N_15096,N_13832);
nor U17255 (N_17255,N_13082,N_15145);
nor U17256 (N_17256,N_12710,N_14165);
and U17257 (N_17257,N_14033,N_13926);
and U17258 (N_17258,N_14154,N_12925);
and U17259 (N_17259,N_15805,N_13113);
nand U17260 (N_17260,N_13680,N_14847);
xor U17261 (N_17261,N_12156,N_13718);
and U17262 (N_17262,N_14769,N_12669);
xor U17263 (N_17263,N_13373,N_14455);
nor U17264 (N_17264,N_13522,N_15166);
or U17265 (N_17265,N_12198,N_15510);
or U17266 (N_17266,N_13299,N_15327);
or U17267 (N_17267,N_12291,N_15624);
nor U17268 (N_17268,N_14540,N_14394);
nand U17269 (N_17269,N_13275,N_14217);
and U17270 (N_17270,N_12595,N_15654);
nor U17271 (N_17271,N_13261,N_12165);
nor U17272 (N_17272,N_15421,N_12330);
nand U17273 (N_17273,N_12520,N_13285);
or U17274 (N_17274,N_13429,N_15694);
and U17275 (N_17275,N_15808,N_12451);
nand U17276 (N_17276,N_15101,N_14508);
nor U17277 (N_17277,N_12176,N_14473);
nand U17278 (N_17278,N_14104,N_13562);
nor U17279 (N_17279,N_14126,N_13032);
or U17280 (N_17280,N_15489,N_14388);
nand U17281 (N_17281,N_14336,N_13090);
xor U17282 (N_17282,N_12378,N_12847);
nor U17283 (N_17283,N_13952,N_15162);
or U17284 (N_17284,N_12509,N_15869);
nand U17285 (N_17285,N_14186,N_12272);
nor U17286 (N_17286,N_12563,N_12867);
nand U17287 (N_17287,N_12134,N_12017);
and U17288 (N_17288,N_15844,N_13504);
nand U17289 (N_17289,N_13725,N_14051);
nor U17290 (N_17290,N_12970,N_14068);
nor U17291 (N_17291,N_15115,N_13481);
nand U17292 (N_17292,N_15250,N_14099);
nor U17293 (N_17293,N_13153,N_15406);
or U17294 (N_17294,N_13581,N_13604);
nor U17295 (N_17295,N_15348,N_12603);
and U17296 (N_17296,N_12316,N_12565);
or U17297 (N_17297,N_14301,N_14693);
and U17298 (N_17298,N_14696,N_12594);
and U17299 (N_17299,N_14147,N_15531);
or U17300 (N_17300,N_15647,N_12029);
nor U17301 (N_17301,N_14966,N_14754);
xor U17302 (N_17302,N_12241,N_13664);
nand U17303 (N_17303,N_12009,N_14714);
nand U17304 (N_17304,N_15638,N_15103);
nor U17305 (N_17305,N_13973,N_12667);
nand U17306 (N_17306,N_15259,N_14555);
nand U17307 (N_17307,N_15051,N_15318);
nor U17308 (N_17308,N_13670,N_13002);
or U17309 (N_17309,N_12792,N_15194);
or U17310 (N_17310,N_15998,N_14069);
nand U17311 (N_17311,N_14260,N_14523);
nand U17312 (N_17312,N_14157,N_14364);
nand U17313 (N_17313,N_13131,N_13241);
nor U17314 (N_17314,N_14319,N_13878);
or U17315 (N_17315,N_12711,N_14875);
nand U17316 (N_17316,N_15916,N_12219);
or U17317 (N_17317,N_15150,N_15619);
and U17318 (N_17318,N_14937,N_12738);
and U17319 (N_17319,N_13871,N_13703);
nor U17320 (N_17320,N_14101,N_14435);
and U17321 (N_17321,N_15740,N_14834);
nor U17322 (N_17322,N_12434,N_15834);
nand U17323 (N_17323,N_14393,N_15486);
and U17324 (N_17324,N_13682,N_14729);
xnor U17325 (N_17325,N_13834,N_13731);
or U17326 (N_17326,N_15848,N_13763);
nand U17327 (N_17327,N_15498,N_12126);
nand U17328 (N_17328,N_14530,N_13991);
nand U17329 (N_17329,N_14478,N_13438);
or U17330 (N_17330,N_13322,N_14600);
xnor U17331 (N_17331,N_12927,N_14308);
nand U17332 (N_17332,N_14351,N_13433);
and U17333 (N_17333,N_12295,N_12168);
nand U17334 (N_17334,N_12874,N_15425);
or U17335 (N_17335,N_13642,N_14687);
and U17336 (N_17336,N_13727,N_13057);
or U17337 (N_17337,N_12060,N_15944);
or U17338 (N_17338,N_14561,N_15196);
or U17339 (N_17339,N_15571,N_15092);
and U17340 (N_17340,N_12324,N_14943);
nor U17341 (N_17341,N_14727,N_14161);
nand U17342 (N_17342,N_13996,N_15082);
and U17343 (N_17343,N_15414,N_14784);
and U17344 (N_17344,N_13813,N_12754);
xor U17345 (N_17345,N_14240,N_15463);
or U17346 (N_17346,N_14491,N_15700);
or U17347 (N_17347,N_15394,N_14141);
and U17348 (N_17348,N_15747,N_13839);
nor U17349 (N_17349,N_13880,N_14839);
nor U17350 (N_17350,N_13203,N_14596);
nor U17351 (N_17351,N_14512,N_14345);
xor U17352 (N_17352,N_12723,N_12173);
nor U17353 (N_17353,N_12951,N_15863);
nor U17354 (N_17354,N_15837,N_14183);
nand U17355 (N_17355,N_12496,N_13217);
or U17356 (N_17356,N_12312,N_15953);
nor U17357 (N_17357,N_12258,N_12364);
or U17358 (N_17358,N_13761,N_12975);
and U17359 (N_17359,N_15448,N_12883);
nand U17360 (N_17360,N_15757,N_14361);
and U17361 (N_17361,N_15067,N_12093);
nor U17362 (N_17362,N_15005,N_13479);
and U17363 (N_17363,N_13348,N_14044);
and U17364 (N_17364,N_15526,N_15547);
and U17365 (N_17365,N_12709,N_12003);
nand U17366 (N_17366,N_12006,N_14050);
nand U17367 (N_17367,N_15010,N_14080);
and U17368 (N_17368,N_13036,N_14334);
nor U17369 (N_17369,N_12057,N_12274);
nor U17370 (N_17370,N_14579,N_15968);
nor U17371 (N_17371,N_13133,N_14806);
xor U17372 (N_17372,N_13572,N_12915);
or U17373 (N_17373,N_12461,N_13888);
nand U17374 (N_17374,N_14447,N_15023);
and U17375 (N_17375,N_12691,N_14900);
or U17376 (N_17376,N_15377,N_14755);
nand U17377 (N_17377,N_12730,N_14535);
and U17378 (N_17378,N_12839,N_13076);
or U17379 (N_17379,N_14017,N_14411);
or U17380 (N_17380,N_13056,N_15598);
nand U17381 (N_17381,N_12541,N_15656);
and U17382 (N_17382,N_15411,N_14440);
or U17383 (N_17383,N_13491,N_14780);
or U17384 (N_17384,N_12472,N_15637);
or U17385 (N_17385,N_15226,N_15516);
and U17386 (N_17386,N_12908,N_15395);
nand U17387 (N_17387,N_12592,N_12752);
and U17388 (N_17388,N_14882,N_14757);
or U17389 (N_17389,N_12267,N_13062);
or U17390 (N_17390,N_14377,N_14060);
nand U17391 (N_17391,N_12540,N_15751);
and U17392 (N_17392,N_15261,N_15646);
nand U17393 (N_17393,N_15146,N_12280);
and U17394 (N_17394,N_14224,N_12782);
or U17395 (N_17395,N_13011,N_15540);
or U17396 (N_17396,N_12536,N_13464);
nand U17397 (N_17397,N_14829,N_15983);
nand U17398 (N_17398,N_13847,N_14464);
nor U17399 (N_17399,N_14381,N_12646);
nor U17400 (N_17400,N_12693,N_13997);
and U17401 (N_17401,N_12814,N_13838);
and U17402 (N_17402,N_12992,N_15755);
and U17403 (N_17403,N_15264,N_12547);
and U17404 (N_17404,N_15809,N_14776);
nand U17405 (N_17405,N_13677,N_12732);
and U17406 (N_17406,N_14105,N_13870);
nand U17407 (N_17407,N_13070,N_12516);
nor U17408 (N_17408,N_13377,N_13064);
and U17409 (N_17409,N_15484,N_15058);
nand U17410 (N_17410,N_15770,N_14752);
xnor U17411 (N_17411,N_15350,N_14926);
and U17412 (N_17412,N_15839,N_15273);
nor U17413 (N_17413,N_15121,N_15936);
and U17414 (N_17414,N_13603,N_14431);
nor U17415 (N_17415,N_15650,N_15838);
nand U17416 (N_17416,N_12220,N_12186);
nand U17417 (N_17417,N_12327,N_15213);
or U17418 (N_17418,N_14117,N_12796);
and U17419 (N_17419,N_12584,N_14580);
nor U17420 (N_17420,N_13181,N_12474);
or U17421 (N_17421,N_12641,N_15591);
nor U17422 (N_17422,N_14284,N_13857);
or U17423 (N_17423,N_14541,N_13901);
nand U17424 (N_17424,N_15227,N_12085);
nor U17425 (N_17425,N_14259,N_12786);
nand U17426 (N_17426,N_13971,N_15138);
nor U17427 (N_17427,N_13028,N_12805);
and U17428 (N_17428,N_13069,N_14844);
or U17429 (N_17429,N_15244,N_12998);
nor U17430 (N_17430,N_13038,N_13132);
and U17431 (N_17431,N_12533,N_13254);
nand U17432 (N_17432,N_15307,N_13923);
xnor U17433 (N_17433,N_12894,N_12171);
nor U17434 (N_17434,N_13423,N_14998);
nand U17435 (N_17435,N_12070,N_15228);
or U17436 (N_17436,N_13197,N_14423);
nand U17437 (N_17437,N_14417,N_15714);
nand U17438 (N_17438,N_13173,N_13846);
and U17439 (N_17439,N_13979,N_15536);
nand U17440 (N_17440,N_15494,N_13526);
nand U17441 (N_17441,N_15100,N_15277);
nor U17442 (N_17442,N_13462,N_14673);
and U17443 (N_17443,N_14775,N_14520);
and U17444 (N_17444,N_14300,N_15543);
xor U17445 (N_17445,N_13177,N_13306);
xnor U17446 (N_17446,N_13936,N_12292);
nand U17447 (N_17447,N_12072,N_13641);
nor U17448 (N_17448,N_12299,N_15081);
or U17449 (N_17449,N_12379,N_12645);
or U17450 (N_17450,N_12266,N_14310);
nand U17451 (N_17451,N_13319,N_13580);
and U17452 (N_17452,N_14148,N_12650);
nor U17453 (N_17453,N_15183,N_12815);
and U17454 (N_17454,N_13175,N_15390);
nand U17455 (N_17455,N_13866,N_15930);
or U17456 (N_17456,N_14467,N_13756);
and U17457 (N_17457,N_13607,N_13209);
or U17458 (N_17458,N_12308,N_12216);
xnor U17459 (N_17459,N_12445,N_14908);
and U17460 (N_17460,N_14629,N_14252);
or U17461 (N_17461,N_15737,N_15786);
or U17462 (N_17462,N_13935,N_15982);
or U17463 (N_17463,N_13872,N_12716);
or U17464 (N_17464,N_15832,N_15323);
nand U17465 (N_17465,N_14663,N_15795);
or U17466 (N_17466,N_13222,N_14933);
or U17467 (N_17467,N_15257,N_12357);
and U17468 (N_17468,N_12396,N_14721);
or U17469 (N_17469,N_15678,N_12783);
and U17470 (N_17470,N_12591,N_14449);
nor U17471 (N_17471,N_14325,N_13431);
nor U17472 (N_17472,N_15192,N_15527);
or U17473 (N_17473,N_14497,N_15497);
nor U17474 (N_17474,N_15469,N_15556);
nand U17475 (N_17475,N_15582,N_14866);
or U17476 (N_17476,N_15507,N_14751);
nor U17477 (N_17477,N_13230,N_13626);
nand U17478 (N_17478,N_13943,N_13951);
nand U17479 (N_17479,N_13492,N_14428);
nand U17480 (N_17480,N_14677,N_12642);
nand U17481 (N_17481,N_14191,N_14576);
nand U17482 (N_17482,N_15946,N_12467);
nand U17483 (N_17483,N_12210,N_12712);
or U17484 (N_17484,N_12877,N_12190);
and U17485 (N_17485,N_15093,N_13367);
and U17486 (N_17486,N_12191,N_15592);
nand U17487 (N_17487,N_14370,N_14916);
and U17488 (N_17488,N_12528,N_14940);
or U17489 (N_17489,N_14624,N_13723);
or U17490 (N_17490,N_15972,N_15362);
or U17491 (N_17491,N_15119,N_12414);
nand U17492 (N_17492,N_15443,N_14668);
and U17493 (N_17493,N_12468,N_15459);
or U17494 (N_17494,N_13994,N_12587);
and U17495 (N_17495,N_14413,N_14765);
xor U17496 (N_17496,N_13060,N_12200);
and U17497 (N_17497,N_15969,N_15502);
nand U17498 (N_17498,N_12002,N_12797);
and U17499 (N_17499,N_12083,N_15768);
or U17500 (N_17500,N_12290,N_14592);
nand U17501 (N_17501,N_15473,N_15888);
nor U17502 (N_17502,N_15015,N_13810);
and U17503 (N_17503,N_12257,N_12137);
nor U17504 (N_17504,N_12222,N_12286);
nor U17505 (N_17505,N_15612,N_15564);
nand U17506 (N_17506,N_13701,N_12008);
nor U17507 (N_17507,N_12215,N_15959);
and U17508 (N_17508,N_14846,N_12600);
and U17509 (N_17509,N_15418,N_13058);
nand U17510 (N_17510,N_15797,N_13985);
nand U17511 (N_17511,N_15238,N_14367);
nand U17512 (N_17512,N_12342,N_15241);
nor U17513 (N_17513,N_14018,N_13605);
or U17514 (N_17514,N_13010,N_12034);
nor U17515 (N_17515,N_12589,N_13449);
nand U17516 (N_17516,N_12338,N_15655);
nand U17517 (N_17517,N_14276,N_13262);
and U17518 (N_17518,N_14400,N_14927);
nor U17519 (N_17519,N_13490,N_12133);
nor U17520 (N_17520,N_14318,N_14091);
nor U17521 (N_17521,N_13192,N_12124);
or U17522 (N_17522,N_12664,N_13909);
or U17523 (N_17523,N_15555,N_13477);
nor U17524 (N_17524,N_12760,N_14710);
or U17525 (N_17525,N_13789,N_12080);
or U17526 (N_17526,N_14016,N_12613);
and U17527 (N_17527,N_13219,N_13720);
nor U17528 (N_17528,N_14513,N_15074);
nand U17529 (N_17529,N_12151,N_12484);
and U17530 (N_17530,N_13505,N_12843);
nand U17531 (N_17531,N_15112,N_14274);
nor U17532 (N_17532,N_14152,N_14852);
nor U17533 (N_17533,N_13975,N_15002);
and U17534 (N_17534,N_13993,N_15256);
nand U17535 (N_17535,N_15109,N_12073);
nor U17536 (N_17536,N_15386,N_14546);
nor U17537 (N_17537,N_15680,N_14185);
nor U17538 (N_17538,N_14509,N_12408);
nor U17539 (N_17539,N_15632,N_12187);
nand U17540 (N_17540,N_13238,N_15672);
nand U17541 (N_17541,N_13401,N_13590);
or U17542 (N_17542,N_14650,N_12231);
xnor U17543 (N_17543,N_12302,N_14504);
nor U17544 (N_17544,N_13755,N_12626);
nand U17545 (N_17545,N_15496,N_12882);
nand U17546 (N_17546,N_13080,N_14880);
or U17547 (N_17547,N_15847,N_13314);
and U17548 (N_17548,N_13862,N_13494);
or U17549 (N_17549,N_13136,N_12038);
or U17550 (N_17550,N_15122,N_14845);
and U17551 (N_17551,N_12092,N_12443);
nor U17552 (N_17552,N_12755,N_13381);
and U17553 (N_17553,N_14611,N_14454);
nor U17554 (N_17554,N_12881,N_15917);
nand U17555 (N_17555,N_15287,N_13887);
nand U17556 (N_17556,N_12827,N_13012);
nor U17557 (N_17557,N_13024,N_12581);
or U17558 (N_17558,N_13055,N_12423);
and U17559 (N_17559,N_15283,N_15588);
nor U17560 (N_17560,N_12248,N_15820);
nor U17561 (N_17561,N_15324,N_15368);
nand U17562 (N_17562,N_13274,N_14986);
nand U17563 (N_17563,N_15212,N_14732);
nor U17564 (N_17564,N_12178,N_12326);
and U17565 (N_17565,N_13063,N_12596);
or U17566 (N_17566,N_12328,N_14059);
xor U17567 (N_17567,N_15039,N_14078);
or U17568 (N_17568,N_13488,N_14403);
or U17569 (N_17569,N_14223,N_14997);
nor U17570 (N_17570,N_15151,N_15904);
or U17571 (N_17571,N_15867,N_14928);
nor U17572 (N_17572,N_15062,N_14146);
and U17573 (N_17573,N_13004,N_12322);
and U17574 (N_17574,N_12750,N_12147);
nand U17575 (N_17575,N_14304,N_12884);
nand U17576 (N_17576,N_14597,N_14614);
nor U17577 (N_17577,N_14990,N_12974);
nor U17578 (N_17578,N_15827,N_15662);
nor U17579 (N_17579,N_12197,N_12804);
and U17580 (N_17580,N_14703,N_15482);
and U17581 (N_17581,N_14689,N_13228);
nor U17582 (N_17582,N_13990,N_15237);
or U17583 (N_17583,N_14020,N_15804);
nand U17584 (N_17584,N_12938,N_12247);
and U17585 (N_17585,N_15470,N_14073);
xor U17586 (N_17586,N_15034,N_12873);
and U17587 (N_17587,N_14655,N_12527);
or U17588 (N_17588,N_15069,N_15219);
nor U17589 (N_17589,N_13648,N_12039);
or U17590 (N_17590,N_15359,N_12104);
nor U17591 (N_17591,N_12437,N_14605);
nor U17592 (N_17592,N_14132,N_15143);
or U17593 (N_17593,N_14481,N_13744);
and U17594 (N_17594,N_15140,N_13908);
nor U17595 (N_17595,N_15681,N_12329);
nor U17596 (N_17596,N_15845,N_14028);
nor U17597 (N_17597,N_13259,N_13840);
or U17598 (N_17598,N_14396,N_14862);
and U17599 (N_17599,N_15634,N_14660);
nor U17600 (N_17600,N_12310,N_13168);
nand U17601 (N_17601,N_15900,N_14438);
nand U17602 (N_17602,N_14257,N_12678);
nand U17603 (N_17603,N_13347,N_14877);
nand U17604 (N_17604,N_15260,N_14397);
nand U17605 (N_17605,N_15485,N_13448);
nand U17606 (N_17606,N_12230,N_12031);
or U17607 (N_17607,N_12235,N_14860);
and U17608 (N_17608,N_12599,N_13365);
nand U17609 (N_17609,N_12452,N_12742);
nor U17610 (N_17610,N_12606,N_15369);
and U17611 (N_17611,N_12388,N_14711);
and U17612 (N_17612,N_14189,N_14408);
nor U17613 (N_17613,N_14461,N_13877);
nor U17614 (N_17614,N_12766,N_15398);
and U17615 (N_17615,N_14563,N_14593);
and U17616 (N_17616,N_15132,N_15309);
and U17617 (N_17617,N_14788,N_14436);
and U17618 (N_17618,N_14635,N_14163);
and U17619 (N_17619,N_12605,N_13375);
and U17620 (N_17620,N_15715,N_12808);
or U17621 (N_17621,N_15852,N_15843);
nor U17622 (N_17622,N_15083,N_14604);
nor U17623 (N_17623,N_13775,N_13524);
nand U17624 (N_17624,N_14444,N_12794);
or U17625 (N_17625,N_13787,N_13308);
nor U17626 (N_17626,N_14620,N_13146);
and U17627 (N_17627,N_14804,N_15603);
or U17628 (N_17628,N_13631,N_13360);
xnor U17629 (N_17629,N_13158,N_15965);
or U17630 (N_17630,N_13077,N_14433);
nand U17631 (N_17631,N_14499,N_13382);
or U17632 (N_17632,N_15293,N_13710);
nor U17633 (N_17633,N_14246,N_12403);
or U17634 (N_17634,N_13608,N_12358);
and U17635 (N_17635,N_13925,N_15173);
or U17636 (N_17636,N_15608,N_14292);
nor U17637 (N_17637,N_14216,N_12918);
or U17638 (N_17638,N_13016,N_12505);
and U17639 (N_17639,N_14818,N_13898);
or U17640 (N_17640,N_12363,N_15657);
and U17641 (N_17641,N_14118,N_12658);
nand U17642 (N_17642,N_14034,N_15682);
or U17643 (N_17643,N_15329,N_12680);
or U17644 (N_17644,N_12784,N_12482);
and U17645 (N_17645,N_12537,N_12278);
or U17646 (N_17646,N_13034,N_14015);
nand U17647 (N_17647,N_13239,N_14353);
and U17648 (N_17648,N_14181,N_12702);
and U17649 (N_17649,N_15883,N_13072);
or U17650 (N_17650,N_12887,N_12557);
or U17651 (N_17651,N_15042,N_14312);
and U17652 (N_17652,N_13533,N_12871);
nand U17653 (N_17653,N_12627,N_12424);
nand U17654 (N_17654,N_12494,N_14550);
or U17655 (N_17655,N_15918,N_14090);
and U17656 (N_17656,N_12535,N_14193);
nand U17657 (N_17657,N_15895,N_12996);
and U17658 (N_17658,N_14169,N_14228);
nand U17659 (N_17659,N_12399,N_14901);
nor U17660 (N_17660,N_13805,N_13585);
xor U17661 (N_17661,N_13947,N_14083);
nor U17662 (N_17662,N_15878,N_12082);
and U17663 (N_17663,N_15605,N_14878);
and U17664 (N_17664,N_13196,N_12188);
nor U17665 (N_17665,N_12888,N_15706);
and U17666 (N_17666,N_14525,N_14190);
or U17667 (N_17667,N_14096,N_12154);
nand U17668 (N_17668,N_15055,N_15155);
nand U17669 (N_17669,N_14180,N_13694);
and U17670 (N_17670,N_15465,N_14511);
nand U17671 (N_17671,N_15222,N_15048);
and U17672 (N_17672,N_12268,N_12331);
and U17673 (N_17673,N_15265,N_12569);
nand U17674 (N_17674,N_12681,N_15423);
or U17675 (N_17675,N_14643,N_14111);
nand U17676 (N_17676,N_12739,N_13922);
nor U17677 (N_17677,N_12163,N_12361);
and U17678 (N_17678,N_13436,N_13307);
or U17679 (N_17679,N_12183,N_13127);
or U17680 (N_17680,N_13693,N_12470);
nand U17681 (N_17681,N_14287,N_12492);
or U17682 (N_17682,N_14324,N_14613);
xor U17683 (N_17683,N_15790,N_13441);
and U17684 (N_17684,N_13924,N_13921);
and U17685 (N_17685,N_15420,N_14167);
nand U17686 (N_17686,N_14483,N_15669);
or U17687 (N_17687,N_12696,N_15991);
and U17688 (N_17688,N_13903,N_15389);
or U17689 (N_17689,N_15490,N_13712);
or U17690 (N_17690,N_12513,N_12014);
nor U17691 (N_17691,N_12317,N_13561);
nand U17692 (N_17692,N_13811,N_12262);
and U17693 (N_17693,N_15695,N_14661);
nor U17694 (N_17694,N_13385,N_14925);
nand U17695 (N_17695,N_12575,N_15054);
or U17696 (N_17696,N_12428,N_13986);
nand U17697 (N_17697,N_15071,N_14488);
nand U17698 (N_17698,N_15235,N_14227);
and U17699 (N_17699,N_15710,N_14277);
nor U17700 (N_17700,N_14887,N_13645);
nand U17701 (N_17701,N_15529,N_13513);
or U17702 (N_17702,N_15361,N_12478);
nand U17703 (N_17703,N_13770,N_14384);
or U17704 (N_17704,N_13915,N_12194);
nand U17705 (N_17705,N_15165,N_12390);
or U17706 (N_17706,N_12130,N_14811);
or U17707 (N_17707,N_13184,N_12886);
nor U17708 (N_17708,N_13458,N_12089);
or U17709 (N_17709,N_15973,N_12860);
nor U17710 (N_17710,N_14547,N_13407);
and U17711 (N_17711,N_13498,N_12890);
nand U17712 (N_17712,N_13595,N_14595);
nand U17713 (N_17713,N_13446,N_15914);
and U17714 (N_17714,N_15573,N_14695);
or U17715 (N_17715,N_13525,N_12920);
and U17716 (N_17716,N_14587,N_14320);
nor U17717 (N_17717,N_15365,N_14489);
and U17718 (N_17718,N_13660,N_12005);
and U17719 (N_17719,N_12728,N_14963);
or U17720 (N_17720,N_12640,N_13450);
nor U17721 (N_17721,N_12318,N_14134);
nor U17722 (N_17722,N_12131,N_12686);
and U17723 (N_17723,N_12320,N_14475);
or U17724 (N_17724,N_12042,N_14531);
nand U17725 (N_17725,N_12580,N_12864);
nor U17726 (N_17726,N_13785,N_13167);
nand U17727 (N_17727,N_12033,N_14422);
or U17728 (N_17728,N_12943,N_12848);
nor U17729 (N_17729,N_12955,N_12425);
or U17730 (N_17730,N_12366,N_12462);
and U17731 (N_17731,N_12350,N_15865);
nand U17732 (N_17732,N_12934,N_13795);
and U17733 (N_17733,N_14329,N_13612);
or U17734 (N_17734,N_15565,N_15011);
and U17735 (N_17735,N_13782,N_14212);
nor U17736 (N_17736,N_15053,N_15148);
and U17737 (N_17737,N_12926,N_13655);
xnor U17738 (N_17738,N_13497,N_12380);
and U17739 (N_17739,N_13237,N_15321);
or U17740 (N_17740,N_13589,N_15928);
nor U17741 (N_17741,N_15450,N_15545);
nand U17742 (N_17742,N_14035,N_15274);
or U17743 (N_17743,N_12651,N_13726);
nor U17744 (N_17744,N_15045,N_13828);
or U17745 (N_17745,N_13854,N_15623);
nand U17746 (N_17746,N_13304,N_13412);
or U17747 (N_17747,N_12895,N_14919);
nor U17748 (N_17748,N_15079,N_14124);
nor U17749 (N_17749,N_15898,N_15938);
nand U17750 (N_17750,N_14848,N_15050);
nor U17751 (N_17751,N_13739,N_15902);
and U17752 (N_17752,N_12125,N_13014);
and U17753 (N_17753,N_12027,N_13003);
nor U17754 (N_17754,N_12392,N_15335);
or U17755 (N_17755,N_12660,N_13435);
or U17756 (N_17756,N_14911,N_15104);
or U17757 (N_17757,N_12683,N_13171);
nor U17758 (N_17758,N_14382,N_12697);
and U17759 (N_17759,N_13395,N_15963);
or U17760 (N_17760,N_15500,N_14054);
or U17761 (N_17761,N_12872,N_13741);
and U17762 (N_17762,N_13189,N_13250);
nand U17763 (N_17763,N_15652,N_12905);
nor U17764 (N_17764,N_14219,N_12355);
or U17765 (N_17765,N_14794,N_12493);
nor U17766 (N_17766,N_14744,N_15703);
nand U17767 (N_17767,N_14144,N_13493);
and U17768 (N_17768,N_13170,N_13646);
nand U17769 (N_17769,N_15346,N_13673);
nor U17770 (N_17770,N_12281,N_15089);
nand U17771 (N_17771,N_15711,N_15990);
or U17772 (N_17772,N_13962,N_14543);
nand U17773 (N_17773,N_14045,N_14637);
and U17774 (N_17774,N_12045,N_13194);
nor U17775 (N_17775,N_15356,N_15685);
or U17776 (N_17776,N_15501,N_15614);
nand U17777 (N_17777,N_15818,N_15676);
nor U17778 (N_17778,N_15223,N_15668);
nor U17779 (N_17779,N_15027,N_14857);
nand U17780 (N_17780,N_15771,N_15799);
and U17781 (N_17781,N_15872,N_13042);
and U17782 (N_17782,N_14282,N_15113);
nand U17783 (N_17783,N_15824,N_13103);
nand U17784 (N_17784,N_15252,N_13895);
and U17785 (N_17785,N_14761,N_13358);
nand U17786 (N_17786,N_15476,N_15434);
nor U17787 (N_17787,N_14450,N_13706);
or U17788 (N_17788,N_15980,N_15643);
or U17789 (N_17789,N_15835,N_13253);
xor U17790 (N_17790,N_14106,N_15876);
nand U17791 (N_17791,N_15128,N_13182);
or U17792 (N_17792,N_12500,N_15649);
nor U17793 (N_17793,N_12652,N_12086);
nor U17794 (N_17794,N_15357,N_13409);
nor U17795 (N_17795,N_12506,N_12199);
nor U17796 (N_17796,N_13086,N_15925);
nand U17797 (N_17797,N_13142,N_15910);
and U17798 (N_17798,N_13886,N_14374);
nor U17799 (N_17799,N_12769,N_15404);
nor U17800 (N_17800,N_12896,N_13255);
or U17801 (N_17801,N_13850,N_13092);
or U17802 (N_17802,N_13883,N_15126);
and U17803 (N_17803,N_13583,N_14445);
and U17804 (N_17804,N_14158,N_12217);
or U17805 (N_17805,N_13252,N_15630);
nand U17806 (N_17806,N_15460,N_14262);
nor U17807 (N_17807,N_15995,N_12305);
nand U17808 (N_17808,N_13309,N_12935);
or U17809 (N_17809,N_13134,N_15085);
and U17810 (N_17810,N_13455,N_12397);
and U17811 (N_17811,N_15144,N_13982);
and U17812 (N_17812,N_14610,N_12416);
nand U17813 (N_17813,N_15090,N_15458);
and U17814 (N_17814,N_12914,N_12745);
xor U17815 (N_17815,N_12426,N_12351);
nand U17816 (N_17816,N_15724,N_14529);
nand U17817 (N_17817,N_15176,N_12343);
nand U17818 (N_17818,N_13366,N_15970);
nand U17819 (N_17819,N_15464,N_12705);
nor U17820 (N_17820,N_15517,N_15815);
or U17821 (N_17821,N_13684,N_13554);
nor U17822 (N_17822,N_14791,N_15211);
and U17823 (N_17823,N_12856,N_14349);
and U17824 (N_17824,N_14254,N_14177);
nand U17825 (N_17825,N_13486,N_14652);
or U17826 (N_17826,N_14019,N_12525);
and U17827 (N_17827,N_14200,N_13914);
and U17828 (N_17828,N_15744,N_12387);
and U17829 (N_17829,N_13162,N_13618);
nor U17830 (N_17830,N_12647,N_14338);
nand U17831 (N_17831,N_13054,N_13001);
nand U17832 (N_17832,N_12909,N_15495);
nor U17833 (N_17833,N_15851,N_12588);
or U17834 (N_17834,N_13570,N_15754);
and U17835 (N_17835,N_15009,N_13568);
nor U17836 (N_17836,N_14448,N_12878);
or U17837 (N_17837,N_14654,N_14768);
or U17838 (N_17838,N_14283,N_15884);
or U17839 (N_17839,N_14810,N_15483);
nand U17840 (N_17840,N_12196,N_12568);
nor U17841 (N_17841,N_12836,N_13882);
or U17842 (N_17842,N_14206,N_12785);
and U17843 (N_17843,N_15317,N_14918);
nand U17844 (N_17844,N_12997,N_14762);
nor U17845 (N_17845,N_12636,N_15258);
or U17846 (N_17846,N_12228,N_15202);
nand U17847 (N_17847,N_12562,N_14972);
or U17848 (N_17848,N_12487,N_15370);
xnor U17849 (N_17849,N_12497,N_15727);
nor U17850 (N_17850,N_12441,N_12990);
nor U17851 (N_17851,N_13625,N_12202);
and U17852 (N_17852,N_15316,N_12144);
nor U17853 (N_17853,N_14722,N_12622);
nand U17854 (N_17854,N_13474,N_15803);
nor U17855 (N_17855,N_12193,N_14426);
or U17856 (N_17856,N_15833,N_15046);
xnor U17857 (N_17857,N_12148,N_13045);
and U17858 (N_17858,N_15689,N_12054);
or U17859 (N_17859,N_13897,N_13786);
and U17860 (N_17860,N_15921,N_15380);
nor U17861 (N_17861,N_13074,N_13861);
nand U17862 (N_17862,N_15345,N_14745);
nand U17863 (N_17863,N_15905,N_13619);
or U17864 (N_17864,N_14196,N_15509);
nand U17865 (N_17865,N_14067,N_13329);
or U17866 (N_17866,N_15584,N_15141);
nor U17867 (N_17867,N_15177,N_14819);
or U17868 (N_17868,N_14443,N_13297);
nand U17869 (N_17869,N_15964,N_13954);
nand U17870 (N_17870,N_14314,N_12790);
nor U17871 (N_17871,N_15761,N_14482);
and U17872 (N_17872,N_14192,N_13799);
and U17873 (N_17873,N_15134,N_14783);
or U17874 (N_17874,N_14591,N_13376);
or U17875 (N_17875,N_14825,N_14778);
or U17876 (N_17876,N_13578,N_15701);
and U17877 (N_17877,N_13667,N_13867);
and U17878 (N_17878,N_12793,N_13515);
nor U17879 (N_17879,N_14366,N_12977);
or U17880 (N_17880,N_13757,N_15861);
or U17881 (N_17881,N_14941,N_15399);
nor U17882 (N_17882,N_14021,N_13776);
nand U17883 (N_17883,N_13457,N_12260);
and U17884 (N_17884,N_12534,N_13622);
and U17885 (N_17885,N_15374,N_15232);
or U17886 (N_17886,N_13470,N_13484);
or U17887 (N_17887,N_15435,N_12143);
or U17888 (N_17888,N_12488,N_13730);
and U17889 (N_17889,N_15696,N_15299);
or U17890 (N_17890,N_12055,N_15759);
xor U17891 (N_17891,N_12612,N_12859);
and U17892 (N_17892,N_12923,N_15935);
nand U17893 (N_17893,N_12121,N_13251);
and U17894 (N_17894,N_12410,N_13485);
nand U17895 (N_17895,N_15830,N_14112);
nor U17896 (N_17896,N_14532,N_12538);
nand U17897 (N_17897,N_15383,N_12644);
nor U17898 (N_17898,N_13596,N_13126);
nor U17899 (N_17899,N_12502,N_14255);
nor U17900 (N_17900,N_12349,N_13191);
nor U17901 (N_17901,N_13812,N_12861);
xor U17902 (N_17902,N_14831,N_15836);
nor U17903 (N_17903,N_14331,N_12558);
and U17904 (N_17904,N_14667,N_13039);
nand U17905 (N_17905,N_13576,N_15595);
or U17906 (N_17906,N_15127,N_15831);
nor U17907 (N_17907,N_13091,N_14516);
or U17908 (N_17908,N_12521,N_12611);
nand U17909 (N_17909,N_12863,N_14812);
and U17910 (N_17910,N_12875,N_14795);
nand U17911 (N_17911,N_12157,N_15787);
nor U17912 (N_17912,N_12756,N_12674);
nand U17913 (N_17913,N_12504,N_14470);
nor U17914 (N_17914,N_15094,N_15105);
and U17915 (N_17915,N_13948,N_12236);
or U17916 (N_17916,N_15198,N_15072);
and U17917 (N_17917,N_14140,N_12892);
or U17918 (N_17918,N_14539,N_12614);
nor U17919 (N_17919,N_15801,N_14973);
and U17920 (N_17920,N_13511,N_14773);
and U17921 (N_17921,N_14369,N_15153);
or U17922 (N_17922,N_15279,N_13545);
nor U17923 (N_17923,N_12932,N_12391);
or U17924 (N_17924,N_14333,N_13964);
nor U17925 (N_17925,N_15030,N_12375);
or U17926 (N_17926,N_14996,N_12939);
or U17927 (N_17927,N_15322,N_13148);
or U17928 (N_17928,N_14094,N_14032);
nor U17929 (N_17929,N_12244,N_13444);
or U17930 (N_17930,N_14121,N_12982);
nand U17931 (N_17931,N_14717,N_15866);
or U17932 (N_17932,N_12430,N_13211);
or U17933 (N_17933,N_13391,N_15301);
nor U17934 (N_17934,N_12068,N_13586);
and U17935 (N_17935,N_12531,N_14160);
or U17936 (N_17936,N_13748,N_12411);
or U17937 (N_17937,N_12633,N_13896);
xnor U17938 (N_17938,N_13339,N_13675);
xor U17939 (N_17939,N_14119,N_12225);
or U17940 (N_17940,N_14676,N_15544);
nand U17941 (N_17941,N_13916,N_12167);
nand U17942 (N_17942,N_13957,N_13507);
or U17943 (N_17943,N_13702,N_13949);
nand U17944 (N_17944,N_12269,N_14471);
nand U17945 (N_17945,N_12566,N_12844);
and U17946 (N_17946,N_14168,N_14835);
or U17947 (N_17947,N_15427,N_15508);
nand U17948 (N_17948,N_15586,N_13472);
nor U17949 (N_17949,N_13860,N_12113);
nand U17950 (N_17950,N_13502,N_12459);
nand U17951 (N_17951,N_14342,N_14738);
nand U17952 (N_17952,N_15943,N_14675);
or U17953 (N_17953,N_14633,N_14938);
nor U17954 (N_17954,N_12913,N_14392);
or U17955 (N_17955,N_14589,N_13403);
nor U17956 (N_17956,N_14496,N_14289);
nor U17957 (N_17957,N_13900,N_14897);
and U17958 (N_17958,N_15734,N_13550);
and U17959 (N_17959,N_14842,N_12714);
and U17960 (N_17960,N_14253,N_14519);
nand U17961 (N_17961,N_15874,N_15960);
and U17962 (N_17962,N_13555,N_14840);
and U17963 (N_17963,N_13451,N_12145);
nor U17964 (N_17964,N_14225,N_13750);
nand U17965 (N_17965,N_15207,N_13855);
and U17966 (N_17966,N_14469,N_14945);
nand U17967 (N_17967,N_14061,N_13652);
nor U17968 (N_17968,N_15466,N_13879);
and U17969 (N_17969,N_15405,N_12265);
nor U17970 (N_17970,N_14923,N_13410);
nor U17971 (N_17971,N_14268,N_13852);
nor U17972 (N_17972,N_14199,N_13023);
nor U17973 (N_17973,N_15745,N_12406);
or U17974 (N_17974,N_13149,N_13097);
nand U17975 (N_17975,N_12967,N_13496);
and U17976 (N_17976,N_15775,N_13236);
or U17977 (N_17977,N_14616,N_14406);
or U17978 (N_17978,N_12675,N_15777);
or U17979 (N_17979,N_14666,N_13278);
and U17980 (N_17980,N_12293,N_14357);
and U17981 (N_17981,N_15086,N_12155);
or U17982 (N_17982,N_14380,N_14885);
or U17983 (N_17983,N_14615,N_15665);
and U17984 (N_17984,N_12333,N_12590);
or U17985 (N_17985,N_14962,N_14131);
or U17986 (N_17986,N_12044,N_13983);
nor U17987 (N_17987,N_13108,N_15538);
nand U17988 (N_17988,N_13657,N_13242);
nand U17989 (N_17989,N_12983,N_14942);
or U17990 (N_17990,N_13233,N_13283);
and U17991 (N_17991,N_13722,N_14418);
nand U17992 (N_17992,N_14699,N_13169);
nand U17993 (N_17993,N_15364,N_12671);
or U17994 (N_17994,N_15885,N_15585);
nand U17995 (N_17995,N_13537,N_14040);
nand U17996 (N_17996,N_13650,N_15693);
nand U17997 (N_17997,N_15722,N_13495);
nand U17998 (N_17998,N_14029,N_15449);
or U17999 (N_17999,N_13033,N_13620);
nor U18000 (N_18000,N_15904,N_15289);
or U18001 (N_18001,N_13822,N_13982);
or U18002 (N_18002,N_13650,N_15028);
nor U18003 (N_18003,N_13716,N_14199);
nor U18004 (N_18004,N_13686,N_12611);
and U18005 (N_18005,N_12636,N_14339);
or U18006 (N_18006,N_13235,N_12464);
or U18007 (N_18007,N_15263,N_12927);
nor U18008 (N_18008,N_13522,N_15469);
nand U18009 (N_18009,N_12693,N_15314);
nand U18010 (N_18010,N_12428,N_15979);
and U18011 (N_18011,N_14144,N_13551);
nand U18012 (N_18012,N_14938,N_13384);
nand U18013 (N_18013,N_12702,N_12211);
or U18014 (N_18014,N_12305,N_13487);
or U18015 (N_18015,N_12190,N_15837);
nor U18016 (N_18016,N_15829,N_15204);
nor U18017 (N_18017,N_14160,N_13159);
nor U18018 (N_18018,N_15982,N_12836);
nand U18019 (N_18019,N_15663,N_15980);
nor U18020 (N_18020,N_13583,N_15807);
nor U18021 (N_18021,N_15434,N_13379);
nor U18022 (N_18022,N_13056,N_12322);
nand U18023 (N_18023,N_14486,N_13493);
nand U18024 (N_18024,N_15202,N_14697);
nor U18025 (N_18025,N_12365,N_12056);
and U18026 (N_18026,N_15302,N_13401);
nor U18027 (N_18027,N_12123,N_12324);
nor U18028 (N_18028,N_15240,N_12688);
and U18029 (N_18029,N_12550,N_15008);
nand U18030 (N_18030,N_14424,N_14377);
nor U18031 (N_18031,N_13137,N_13865);
or U18032 (N_18032,N_13963,N_13886);
nor U18033 (N_18033,N_15600,N_12552);
and U18034 (N_18034,N_13510,N_12880);
or U18035 (N_18035,N_14397,N_15222);
or U18036 (N_18036,N_12211,N_14617);
and U18037 (N_18037,N_13614,N_15365);
nand U18038 (N_18038,N_15005,N_12732);
or U18039 (N_18039,N_15612,N_15883);
nand U18040 (N_18040,N_13984,N_12194);
and U18041 (N_18041,N_14050,N_14625);
nor U18042 (N_18042,N_13966,N_14209);
and U18043 (N_18043,N_15638,N_15111);
nor U18044 (N_18044,N_13316,N_14847);
nor U18045 (N_18045,N_13856,N_13544);
and U18046 (N_18046,N_14248,N_15730);
and U18047 (N_18047,N_15915,N_14580);
nor U18048 (N_18048,N_14236,N_14127);
or U18049 (N_18049,N_14617,N_12402);
nor U18050 (N_18050,N_13112,N_13841);
and U18051 (N_18051,N_13473,N_14983);
nand U18052 (N_18052,N_14389,N_15437);
nor U18053 (N_18053,N_15801,N_12146);
or U18054 (N_18054,N_15327,N_12322);
or U18055 (N_18055,N_14619,N_12422);
nor U18056 (N_18056,N_15108,N_15913);
and U18057 (N_18057,N_15921,N_12901);
and U18058 (N_18058,N_14061,N_15337);
and U18059 (N_18059,N_14216,N_15287);
or U18060 (N_18060,N_15106,N_14393);
or U18061 (N_18061,N_13783,N_15943);
and U18062 (N_18062,N_14444,N_15936);
nor U18063 (N_18063,N_13591,N_14850);
nor U18064 (N_18064,N_12798,N_15023);
and U18065 (N_18065,N_12233,N_15132);
and U18066 (N_18066,N_14693,N_14730);
nor U18067 (N_18067,N_14060,N_12543);
and U18068 (N_18068,N_15320,N_14341);
nand U18069 (N_18069,N_15264,N_15902);
nor U18070 (N_18070,N_13103,N_13526);
xor U18071 (N_18071,N_13319,N_13571);
or U18072 (N_18072,N_14107,N_15523);
nand U18073 (N_18073,N_13352,N_13701);
nor U18074 (N_18074,N_13192,N_12413);
xnor U18075 (N_18075,N_15611,N_12542);
nor U18076 (N_18076,N_15245,N_12956);
nand U18077 (N_18077,N_15589,N_12867);
nand U18078 (N_18078,N_13995,N_13285);
nor U18079 (N_18079,N_15077,N_13905);
nor U18080 (N_18080,N_15221,N_12351);
nor U18081 (N_18081,N_12417,N_13526);
and U18082 (N_18082,N_12646,N_12882);
nor U18083 (N_18083,N_12187,N_15715);
nand U18084 (N_18084,N_12860,N_14729);
nand U18085 (N_18085,N_13702,N_15295);
nor U18086 (N_18086,N_13198,N_15131);
or U18087 (N_18087,N_12916,N_15505);
nand U18088 (N_18088,N_14257,N_15911);
nand U18089 (N_18089,N_14814,N_12324);
and U18090 (N_18090,N_14700,N_12254);
nand U18091 (N_18091,N_14065,N_12273);
and U18092 (N_18092,N_13293,N_14913);
nor U18093 (N_18093,N_15684,N_15130);
and U18094 (N_18094,N_13226,N_15859);
nor U18095 (N_18095,N_14328,N_14733);
or U18096 (N_18096,N_13110,N_12414);
and U18097 (N_18097,N_14544,N_15932);
or U18098 (N_18098,N_13938,N_12714);
xor U18099 (N_18099,N_12095,N_12434);
and U18100 (N_18100,N_15657,N_14028);
or U18101 (N_18101,N_15352,N_15978);
nand U18102 (N_18102,N_13995,N_14860);
or U18103 (N_18103,N_13832,N_13424);
nand U18104 (N_18104,N_13058,N_13645);
nor U18105 (N_18105,N_14264,N_13012);
nand U18106 (N_18106,N_12315,N_12546);
and U18107 (N_18107,N_14825,N_12091);
nor U18108 (N_18108,N_13090,N_12719);
and U18109 (N_18109,N_13626,N_14211);
or U18110 (N_18110,N_12745,N_12357);
and U18111 (N_18111,N_13666,N_13733);
nor U18112 (N_18112,N_13939,N_14308);
nand U18113 (N_18113,N_14764,N_13445);
and U18114 (N_18114,N_15602,N_13580);
nor U18115 (N_18115,N_12108,N_15244);
or U18116 (N_18116,N_14163,N_13755);
or U18117 (N_18117,N_12846,N_15453);
or U18118 (N_18118,N_14418,N_13237);
nor U18119 (N_18119,N_14288,N_13253);
xor U18120 (N_18120,N_14475,N_13231);
or U18121 (N_18121,N_14794,N_14361);
nand U18122 (N_18122,N_13776,N_14667);
and U18123 (N_18123,N_15189,N_14922);
or U18124 (N_18124,N_12654,N_12607);
nand U18125 (N_18125,N_14092,N_13289);
nand U18126 (N_18126,N_12745,N_12810);
nor U18127 (N_18127,N_12974,N_12276);
nand U18128 (N_18128,N_13569,N_15396);
and U18129 (N_18129,N_13674,N_14760);
and U18130 (N_18130,N_12262,N_13266);
and U18131 (N_18131,N_15244,N_14057);
xor U18132 (N_18132,N_13223,N_15842);
and U18133 (N_18133,N_14478,N_12999);
nor U18134 (N_18134,N_12672,N_13810);
nor U18135 (N_18135,N_14333,N_14732);
nand U18136 (N_18136,N_15324,N_13544);
or U18137 (N_18137,N_15493,N_15472);
or U18138 (N_18138,N_14141,N_13924);
and U18139 (N_18139,N_14296,N_13106);
nor U18140 (N_18140,N_12144,N_12792);
nand U18141 (N_18141,N_13249,N_12695);
nand U18142 (N_18142,N_15943,N_15934);
and U18143 (N_18143,N_12036,N_15332);
nor U18144 (N_18144,N_13270,N_13431);
and U18145 (N_18145,N_14826,N_14967);
or U18146 (N_18146,N_12879,N_13958);
or U18147 (N_18147,N_15112,N_15268);
nor U18148 (N_18148,N_13541,N_13063);
or U18149 (N_18149,N_14415,N_12474);
nand U18150 (N_18150,N_13538,N_13372);
and U18151 (N_18151,N_13941,N_13554);
or U18152 (N_18152,N_13816,N_13229);
nand U18153 (N_18153,N_13868,N_13263);
xor U18154 (N_18154,N_15438,N_13155);
nor U18155 (N_18155,N_15550,N_15912);
nand U18156 (N_18156,N_12669,N_12711);
nand U18157 (N_18157,N_15365,N_13403);
nand U18158 (N_18158,N_13229,N_12365);
or U18159 (N_18159,N_13800,N_13978);
and U18160 (N_18160,N_13255,N_15223);
or U18161 (N_18161,N_13624,N_15965);
or U18162 (N_18162,N_14729,N_13538);
nand U18163 (N_18163,N_14750,N_14452);
nand U18164 (N_18164,N_13257,N_12176);
nand U18165 (N_18165,N_12208,N_15451);
xnor U18166 (N_18166,N_15881,N_13641);
or U18167 (N_18167,N_14304,N_13006);
nand U18168 (N_18168,N_15691,N_13956);
nand U18169 (N_18169,N_14271,N_13156);
and U18170 (N_18170,N_15133,N_15276);
and U18171 (N_18171,N_14910,N_15295);
or U18172 (N_18172,N_13156,N_15048);
or U18173 (N_18173,N_14453,N_12219);
or U18174 (N_18174,N_15196,N_14758);
nor U18175 (N_18175,N_12471,N_14947);
and U18176 (N_18176,N_14536,N_15230);
nor U18177 (N_18177,N_12500,N_14005);
nor U18178 (N_18178,N_14254,N_12628);
nand U18179 (N_18179,N_13514,N_15953);
nand U18180 (N_18180,N_15023,N_14356);
nor U18181 (N_18181,N_13389,N_14727);
and U18182 (N_18182,N_13340,N_15807);
or U18183 (N_18183,N_12258,N_13134);
and U18184 (N_18184,N_14565,N_13350);
or U18185 (N_18185,N_12912,N_13294);
and U18186 (N_18186,N_12748,N_14410);
and U18187 (N_18187,N_13253,N_13385);
and U18188 (N_18188,N_13419,N_15261);
or U18189 (N_18189,N_15528,N_13091);
nand U18190 (N_18190,N_12067,N_15205);
xnor U18191 (N_18191,N_15003,N_15049);
or U18192 (N_18192,N_15616,N_15949);
and U18193 (N_18193,N_13397,N_14402);
nand U18194 (N_18194,N_13376,N_14682);
nor U18195 (N_18195,N_12344,N_13675);
or U18196 (N_18196,N_13655,N_12924);
nand U18197 (N_18197,N_14923,N_15361);
or U18198 (N_18198,N_13673,N_15548);
and U18199 (N_18199,N_14326,N_12112);
or U18200 (N_18200,N_15850,N_15339);
or U18201 (N_18201,N_14856,N_14841);
and U18202 (N_18202,N_13666,N_15777);
nor U18203 (N_18203,N_15568,N_13746);
nand U18204 (N_18204,N_13988,N_15177);
nor U18205 (N_18205,N_15116,N_14888);
or U18206 (N_18206,N_15678,N_15153);
nor U18207 (N_18207,N_13819,N_12518);
nor U18208 (N_18208,N_14576,N_13185);
or U18209 (N_18209,N_15287,N_12647);
or U18210 (N_18210,N_12070,N_15253);
or U18211 (N_18211,N_12367,N_12613);
nor U18212 (N_18212,N_14009,N_14212);
nand U18213 (N_18213,N_12431,N_14245);
nand U18214 (N_18214,N_15388,N_14312);
and U18215 (N_18215,N_15036,N_13522);
nor U18216 (N_18216,N_15443,N_13486);
nand U18217 (N_18217,N_15650,N_15721);
nor U18218 (N_18218,N_14006,N_12447);
nor U18219 (N_18219,N_15678,N_13116);
nand U18220 (N_18220,N_12563,N_14002);
nor U18221 (N_18221,N_14739,N_13165);
nor U18222 (N_18222,N_15237,N_12268);
nand U18223 (N_18223,N_12937,N_13503);
or U18224 (N_18224,N_13574,N_14029);
nand U18225 (N_18225,N_14424,N_15967);
and U18226 (N_18226,N_14773,N_12585);
and U18227 (N_18227,N_12696,N_15266);
nand U18228 (N_18228,N_12379,N_13815);
nand U18229 (N_18229,N_15526,N_14427);
and U18230 (N_18230,N_12557,N_14876);
nand U18231 (N_18231,N_12058,N_15096);
or U18232 (N_18232,N_14261,N_14729);
and U18233 (N_18233,N_13037,N_15959);
and U18234 (N_18234,N_12672,N_13499);
and U18235 (N_18235,N_14573,N_15023);
nor U18236 (N_18236,N_15920,N_14828);
and U18237 (N_18237,N_13050,N_15112);
or U18238 (N_18238,N_14177,N_15763);
and U18239 (N_18239,N_12990,N_12231);
or U18240 (N_18240,N_12815,N_12536);
and U18241 (N_18241,N_12957,N_13069);
or U18242 (N_18242,N_15902,N_12890);
nor U18243 (N_18243,N_12688,N_14720);
nand U18244 (N_18244,N_12413,N_14262);
nor U18245 (N_18245,N_13652,N_12789);
or U18246 (N_18246,N_13310,N_14199);
nor U18247 (N_18247,N_15768,N_13589);
nor U18248 (N_18248,N_12529,N_15113);
nand U18249 (N_18249,N_13216,N_12632);
or U18250 (N_18250,N_14714,N_12186);
nand U18251 (N_18251,N_15164,N_12081);
nor U18252 (N_18252,N_12101,N_14269);
nor U18253 (N_18253,N_15918,N_13496);
or U18254 (N_18254,N_13089,N_12456);
and U18255 (N_18255,N_13382,N_15664);
nand U18256 (N_18256,N_13090,N_15346);
or U18257 (N_18257,N_14229,N_13727);
xnor U18258 (N_18258,N_12283,N_14943);
nor U18259 (N_18259,N_12220,N_15116);
or U18260 (N_18260,N_15918,N_15800);
nor U18261 (N_18261,N_13440,N_13406);
or U18262 (N_18262,N_14727,N_14632);
nand U18263 (N_18263,N_14741,N_12261);
or U18264 (N_18264,N_12474,N_15444);
or U18265 (N_18265,N_14405,N_15327);
and U18266 (N_18266,N_12779,N_13849);
and U18267 (N_18267,N_12097,N_15710);
and U18268 (N_18268,N_15001,N_15703);
or U18269 (N_18269,N_12873,N_12937);
and U18270 (N_18270,N_12839,N_15205);
nand U18271 (N_18271,N_14417,N_15956);
and U18272 (N_18272,N_13981,N_15859);
and U18273 (N_18273,N_14953,N_13586);
and U18274 (N_18274,N_12873,N_14618);
and U18275 (N_18275,N_13230,N_12894);
nand U18276 (N_18276,N_14148,N_14086);
and U18277 (N_18277,N_15719,N_14868);
nand U18278 (N_18278,N_12394,N_14712);
and U18279 (N_18279,N_12754,N_14530);
or U18280 (N_18280,N_13083,N_14228);
nand U18281 (N_18281,N_15925,N_13992);
and U18282 (N_18282,N_15536,N_13316);
and U18283 (N_18283,N_15585,N_14314);
nand U18284 (N_18284,N_15146,N_13118);
or U18285 (N_18285,N_14340,N_15272);
and U18286 (N_18286,N_12110,N_14634);
and U18287 (N_18287,N_13559,N_12414);
nor U18288 (N_18288,N_12099,N_14740);
and U18289 (N_18289,N_15768,N_12027);
or U18290 (N_18290,N_13217,N_15509);
and U18291 (N_18291,N_14081,N_12008);
nand U18292 (N_18292,N_13983,N_13477);
or U18293 (N_18293,N_12462,N_13151);
or U18294 (N_18294,N_14735,N_12964);
and U18295 (N_18295,N_12272,N_13628);
and U18296 (N_18296,N_12522,N_15919);
nand U18297 (N_18297,N_12875,N_14585);
nand U18298 (N_18298,N_13498,N_13694);
nand U18299 (N_18299,N_13649,N_15937);
nor U18300 (N_18300,N_13963,N_12930);
or U18301 (N_18301,N_15598,N_14262);
and U18302 (N_18302,N_12695,N_13946);
or U18303 (N_18303,N_12070,N_13815);
nor U18304 (N_18304,N_15031,N_13134);
nor U18305 (N_18305,N_12016,N_14693);
or U18306 (N_18306,N_14676,N_14792);
nor U18307 (N_18307,N_12279,N_15829);
nand U18308 (N_18308,N_14711,N_14718);
nand U18309 (N_18309,N_14440,N_13180);
and U18310 (N_18310,N_15463,N_12040);
nor U18311 (N_18311,N_15116,N_12712);
nand U18312 (N_18312,N_13468,N_14947);
xor U18313 (N_18313,N_15621,N_13606);
nor U18314 (N_18314,N_12512,N_12673);
nor U18315 (N_18315,N_13167,N_13946);
nor U18316 (N_18316,N_14784,N_13660);
nand U18317 (N_18317,N_15874,N_13174);
nand U18318 (N_18318,N_14400,N_14918);
and U18319 (N_18319,N_13962,N_12774);
and U18320 (N_18320,N_15707,N_15885);
nand U18321 (N_18321,N_14476,N_14946);
nor U18322 (N_18322,N_14610,N_12746);
or U18323 (N_18323,N_12174,N_12957);
nand U18324 (N_18324,N_15513,N_13248);
or U18325 (N_18325,N_12686,N_12026);
nand U18326 (N_18326,N_15650,N_14434);
or U18327 (N_18327,N_13482,N_14782);
nor U18328 (N_18328,N_12620,N_12968);
and U18329 (N_18329,N_14208,N_15257);
xnor U18330 (N_18330,N_12924,N_15825);
xor U18331 (N_18331,N_12446,N_13076);
and U18332 (N_18332,N_12387,N_14077);
and U18333 (N_18333,N_12058,N_14993);
or U18334 (N_18334,N_14299,N_14838);
or U18335 (N_18335,N_12700,N_14746);
or U18336 (N_18336,N_14083,N_12412);
xnor U18337 (N_18337,N_12760,N_12592);
and U18338 (N_18338,N_14545,N_12012);
nand U18339 (N_18339,N_13210,N_13352);
nor U18340 (N_18340,N_13617,N_15175);
nand U18341 (N_18341,N_12789,N_13613);
or U18342 (N_18342,N_12843,N_13958);
and U18343 (N_18343,N_12259,N_12458);
xnor U18344 (N_18344,N_15839,N_15413);
nand U18345 (N_18345,N_13224,N_13289);
and U18346 (N_18346,N_14912,N_15340);
xnor U18347 (N_18347,N_12993,N_14348);
nor U18348 (N_18348,N_12098,N_15053);
and U18349 (N_18349,N_14429,N_15184);
nor U18350 (N_18350,N_12255,N_14225);
and U18351 (N_18351,N_14468,N_12575);
nand U18352 (N_18352,N_15147,N_15006);
xnor U18353 (N_18353,N_14715,N_13212);
and U18354 (N_18354,N_13255,N_13301);
and U18355 (N_18355,N_13066,N_12204);
or U18356 (N_18356,N_12276,N_13555);
or U18357 (N_18357,N_15071,N_14996);
or U18358 (N_18358,N_13819,N_12609);
nand U18359 (N_18359,N_12684,N_12988);
nand U18360 (N_18360,N_15727,N_15730);
or U18361 (N_18361,N_13185,N_12692);
and U18362 (N_18362,N_15007,N_13173);
nand U18363 (N_18363,N_12152,N_13156);
nor U18364 (N_18364,N_13729,N_13657);
and U18365 (N_18365,N_13988,N_12597);
or U18366 (N_18366,N_12101,N_14653);
or U18367 (N_18367,N_14410,N_14622);
and U18368 (N_18368,N_12073,N_13089);
xor U18369 (N_18369,N_15924,N_15800);
nand U18370 (N_18370,N_15057,N_12975);
or U18371 (N_18371,N_13852,N_12012);
nor U18372 (N_18372,N_13650,N_15848);
nor U18373 (N_18373,N_14702,N_14742);
nor U18374 (N_18374,N_13714,N_14810);
nand U18375 (N_18375,N_14282,N_13955);
or U18376 (N_18376,N_13006,N_13193);
nor U18377 (N_18377,N_14340,N_15337);
nand U18378 (N_18378,N_15031,N_15423);
nand U18379 (N_18379,N_13033,N_15354);
and U18380 (N_18380,N_12326,N_15326);
nor U18381 (N_18381,N_13044,N_13524);
nand U18382 (N_18382,N_12020,N_12764);
nand U18383 (N_18383,N_14898,N_12778);
nand U18384 (N_18384,N_12793,N_12480);
or U18385 (N_18385,N_15751,N_15147);
xnor U18386 (N_18386,N_15850,N_12106);
nand U18387 (N_18387,N_12190,N_13825);
nand U18388 (N_18388,N_15317,N_13322);
and U18389 (N_18389,N_15032,N_12781);
and U18390 (N_18390,N_13153,N_13394);
or U18391 (N_18391,N_12947,N_15628);
and U18392 (N_18392,N_14565,N_12165);
nand U18393 (N_18393,N_14344,N_15479);
or U18394 (N_18394,N_14349,N_12793);
and U18395 (N_18395,N_12517,N_15856);
nand U18396 (N_18396,N_13589,N_15039);
nand U18397 (N_18397,N_12122,N_12991);
nand U18398 (N_18398,N_14073,N_13344);
nor U18399 (N_18399,N_14187,N_12127);
nor U18400 (N_18400,N_12290,N_12146);
nor U18401 (N_18401,N_13251,N_12400);
nand U18402 (N_18402,N_13045,N_12812);
and U18403 (N_18403,N_12819,N_12882);
or U18404 (N_18404,N_12147,N_12330);
nor U18405 (N_18405,N_14237,N_12320);
and U18406 (N_18406,N_14225,N_14112);
or U18407 (N_18407,N_13697,N_14751);
nor U18408 (N_18408,N_12578,N_12529);
nand U18409 (N_18409,N_13362,N_15139);
nor U18410 (N_18410,N_14492,N_12416);
or U18411 (N_18411,N_15599,N_14671);
xor U18412 (N_18412,N_13313,N_15980);
or U18413 (N_18413,N_15385,N_15016);
and U18414 (N_18414,N_14874,N_14234);
nor U18415 (N_18415,N_15991,N_13920);
nor U18416 (N_18416,N_13949,N_14354);
or U18417 (N_18417,N_13311,N_13444);
or U18418 (N_18418,N_14205,N_15377);
nor U18419 (N_18419,N_15533,N_13394);
or U18420 (N_18420,N_13946,N_12296);
nor U18421 (N_18421,N_15339,N_13713);
nor U18422 (N_18422,N_14838,N_12240);
nand U18423 (N_18423,N_15324,N_13656);
or U18424 (N_18424,N_13550,N_14043);
nand U18425 (N_18425,N_15617,N_12634);
nand U18426 (N_18426,N_14464,N_12035);
or U18427 (N_18427,N_12122,N_14902);
nand U18428 (N_18428,N_13614,N_15501);
nand U18429 (N_18429,N_14791,N_13612);
or U18430 (N_18430,N_13989,N_12862);
nor U18431 (N_18431,N_12974,N_14156);
and U18432 (N_18432,N_15229,N_15753);
or U18433 (N_18433,N_15745,N_12202);
or U18434 (N_18434,N_15634,N_15203);
and U18435 (N_18435,N_14043,N_13617);
or U18436 (N_18436,N_14632,N_12182);
xor U18437 (N_18437,N_14850,N_12319);
nor U18438 (N_18438,N_14518,N_14583);
or U18439 (N_18439,N_12162,N_13249);
nor U18440 (N_18440,N_13992,N_15648);
nor U18441 (N_18441,N_13188,N_12100);
nor U18442 (N_18442,N_12170,N_13831);
and U18443 (N_18443,N_14098,N_12670);
nand U18444 (N_18444,N_13006,N_12126);
or U18445 (N_18445,N_15693,N_13574);
nor U18446 (N_18446,N_15722,N_15166);
xor U18447 (N_18447,N_12637,N_12467);
nand U18448 (N_18448,N_15390,N_15742);
nor U18449 (N_18449,N_12779,N_13910);
or U18450 (N_18450,N_14974,N_13873);
or U18451 (N_18451,N_15371,N_13155);
and U18452 (N_18452,N_15564,N_15675);
and U18453 (N_18453,N_14139,N_12908);
or U18454 (N_18454,N_13019,N_14234);
and U18455 (N_18455,N_15057,N_14326);
nand U18456 (N_18456,N_15427,N_13094);
or U18457 (N_18457,N_13441,N_14901);
or U18458 (N_18458,N_14135,N_14863);
xor U18459 (N_18459,N_14463,N_15855);
or U18460 (N_18460,N_14094,N_15250);
and U18461 (N_18461,N_15382,N_13620);
nor U18462 (N_18462,N_12579,N_12238);
nand U18463 (N_18463,N_15141,N_13333);
nor U18464 (N_18464,N_15011,N_15418);
or U18465 (N_18465,N_12506,N_13402);
nor U18466 (N_18466,N_13524,N_15899);
or U18467 (N_18467,N_13678,N_15545);
or U18468 (N_18468,N_12450,N_12436);
or U18469 (N_18469,N_13687,N_13387);
nand U18470 (N_18470,N_13224,N_12838);
or U18471 (N_18471,N_13677,N_14067);
and U18472 (N_18472,N_12613,N_12008);
nand U18473 (N_18473,N_12203,N_12634);
or U18474 (N_18474,N_13066,N_14085);
nand U18475 (N_18475,N_14419,N_15434);
and U18476 (N_18476,N_12508,N_13443);
and U18477 (N_18477,N_14930,N_15889);
and U18478 (N_18478,N_13225,N_15646);
and U18479 (N_18479,N_12167,N_12749);
nand U18480 (N_18480,N_15062,N_14633);
nand U18481 (N_18481,N_12570,N_14994);
and U18482 (N_18482,N_15554,N_12446);
and U18483 (N_18483,N_15616,N_15521);
nand U18484 (N_18484,N_14731,N_12695);
or U18485 (N_18485,N_14144,N_12199);
nand U18486 (N_18486,N_12710,N_12353);
and U18487 (N_18487,N_14610,N_15618);
nor U18488 (N_18488,N_12572,N_13630);
nand U18489 (N_18489,N_12050,N_13626);
xnor U18490 (N_18490,N_15317,N_14988);
nand U18491 (N_18491,N_14208,N_13094);
nor U18492 (N_18492,N_12590,N_15039);
nor U18493 (N_18493,N_13909,N_15555);
nor U18494 (N_18494,N_14146,N_13358);
nand U18495 (N_18495,N_14173,N_12538);
and U18496 (N_18496,N_12295,N_12770);
nor U18497 (N_18497,N_13994,N_14085);
nor U18498 (N_18498,N_12871,N_14622);
nor U18499 (N_18499,N_13342,N_15336);
nand U18500 (N_18500,N_12893,N_14371);
nor U18501 (N_18501,N_14481,N_15248);
or U18502 (N_18502,N_12516,N_13627);
nor U18503 (N_18503,N_12253,N_12198);
nand U18504 (N_18504,N_13275,N_14719);
and U18505 (N_18505,N_12636,N_14260);
and U18506 (N_18506,N_15511,N_15773);
nand U18507 (N_18507,N_12501,N_12147);
nor U18508 (N_18508,N_14977,N_15081);
nand U18509 (N_18509,N_15757,N_13318);
and U18510 (N_18510,N_13339,N_13351);
nand U18511 (N_18511,N_15423,N_15181);
nand U18512 (N_18512,N_13647,N_12450);
or U18513 (N_18513,N_12732,N_14495);
and U18514 (N_18514,N_13521,N_13425);
or U18515 (N_18515,N_14448,N_12365);
nand U18516 (N_18516,N_12254,N_13258);
nand U18517 (N_18517,N_12303,N_14453);
nand U18518 (N_18518,N_13088,N_12555);
and U18519 (N_18519,N_15215,N_15079);
nand U18520 (N_18520,N_15529,N_13488);
and U18521 (N_18521,N_15073,N_15515);
and U18522 (N_18522,N_12721,N_14221);
and U18523 (N_18523,N_14428,N_13647);
nand U18524 (N_18524,N_14612,N_13034);
and U18525 (N_18525,N_13630,N_15727);
nor U18526 (N_18526,N_13277,N_15194);
nand U18527 (N_18527,N_14693,N_15432);
and U18528 (N_18528,N_13979,N_15107);
or U18529 (N_18529,N_12086,N_14284);
or U18530 (N_18530,N_14615,N_14613);
nor U18531 (N_18531,N_14342,N_13249);
nor U18532 (N_18532,N_14360,N_14905);
nor U18533 (N_18533,N_12331,N_13070);
nand U18534 (N_18534,N_15810,N_14021);
or U18535 (N_18535,N_13281,N_14127);
nand U18536 (N_18536,N_12288,N_15851);
nor U18537 (N_18537,N_12760,N_13199);
nand U18538 (N_18538,N_15116,N_15381);
or U18539 (N_18539,N_15609,N_15365);
or U18540 (N_18540,N_12792,N_14571);
and U18541 (N_18541,N_13666,N_14661);
nor U18542 (N_18542,N_12873,N_14115);
or U18543 (N_18543,N_14096,N_15192);
or U18544 (N_18544,N_13208,N_14144);
nand U18545 (N_18545,N_14466,N_13599);
or U18546 (N_18546,N_15902,N_13251);
nand U18547 (N_18547,N_13986,N_14276);
and U18548 (N_18548,N_14508,N_14438);
and U18549 (N_18549,N_15674,N_13265);
nor U18550 (N_18550,N_14168,N_14191);
nor U18551 (N_18551,N_15411,N_15051);
nor U18552 (N_18552,N_12336,N_12077);
and U18553 (N_18553,N_13494,N_13019);
and U18554 (N_18554,N_13849,N_13634);
and U18555 (N_18555,N_13733,N_15646);
and U18556 (N_18556,N_12171,N_12272);
nor U18557 (N_18557,N_14550,N_14946);
and U18558 (N_18558,N_13434,N_15400);
or U18559 (N_18559,N_13699,N_12110);
or U18560 (N_18560,N_12506,N_15238);
or U18561 (N_18561,N_15527,N_13827);
or U18562 (N_18562,N_13575,N_15505);
or U18563 (N_18563,N_14387,N_14031);
nor U18564 (N_18564,N_14599,N_14026);
nor U18565 (N_18565,N_13952,N_14664);
nand U18566 (N_18566,N_14824,N_15207);
and U18567 (N_18567,N_12429,N_15449);
or U18568 (N_18568,N_15146,N_15635);
nor U18569 (N_18569,N_15454,N_13169);
nand U18570 (N_18570,N_15843,N_14227);
nand U18571 (N_18571,N_15108,N_14384);
and U18572 (N_18572,N_12969,N_12284);
nor U18573 (N_18573,N_15432,N_15069);
nand U18574 (N_18574,N_15186,N_14817);
nor U18575 (N_18575,N_13863,N_15588);
nor U18576 (N_18576,N_12467,N_13370);
or U18577 (N_18577,N_14288,N_13169);
nor U18578 (N_18578,N_14217,N_14109);
or U18579 (N_18579,N_15384,N_13522);
and U18580 (N_18580,N_14585,N_12706);
or U18581 (N_18581,N_15501,N_15125);
nand U18582 (N_18582,N_13757,N_12241);
or U18583 (N_18583,N_15882,N_15947);
and U18584 (N_18584,N_14178,N_13215);
nor U18585 (N_18585,N_14837,N_15994);
or U18586 (N_18586,N_13167,N_12610);
nor U18587 (N_18587,N_15361,N_12802);
nor U18588 (N_18588,N_12829,N_14549);
or U18589 (N_18589,N_15848,N_12715);
nand U18590 (N_18590,N_12850,N_15735);
nor U18591 (N_18591,N_14131,N_13188);
nand U18592 (N_18592,N_12879,N_15059);
or U18593 (N_18593,N_15027,N_15424);
and U18594 (N_18594,N_13441,N_12892);
or U18595 (N_18595,N_13941,N_15373);
nor U18596 (N_18596,N_14154,N_12719);
nand U18597 (N_18597,N_12501,N_15504);
nand U18598 (N_18598,N_14915,N_13060);
nand U18599 (N_18599,N_15751,N_13930);
nand U18600 (N_18600,N_14955,N_15946);
or U18601 (N_18601,N_15955,N_14592);
and U18602 (N_18602,N_12579,N_15996);
nand U18603 (N_18603,N_13783,N_15518);
nor U18604 (N_18604,N_12757,N_14082);
or U18605 (N_18605,N_13149,N_14305);
or U18606 (N_18606,N_13381,N_13169);
nor U18607 (N_18607,N_14516,N_15116);
or U18608 (N_18608,N_13426,N_15632);
xor U18609 (N_18609,N_12510,N_12532);
nor U18610 (N_18610,N_12729,N_12637);
nor U18611 (N_18611,N_12940,N_13262);
or U18612 (N_18612,N_13301,N_13924);
nand U18613 (N_18613,N_15142,N_14606);
nor U18614 (N_18614,N_14125,N_15114);
and U18615 (N_18615,N_13415,N_13037);
nor U18616 (N_18616,N_14898,N_15221);
or U18617 (N_18617,N_12589,N_13008);
nor U18618 (N_18618,N_15313,N_15254);
nor U18619 (N_18619,N_15892,N_12342);
nor U18620 (N_18620,N_14886,N_13802);
nand U18621 (N_18621,N_12567,N_12503);
or U18622 (N_18622,N_15690,N_14808);
or U18623 (N_18623,N_12526,N_14479);
nand U18624 (N_18624,N_14064,N_13095);
nor U18625 (N_18625,N_12323,N_13935);
xor U18626 (N_18626,N_14909,N_15859);
and U18627 (N_18627,N_14372,N_15759);
and U18628 (N_18628,N_12108,N_13759);
or U18629 (N_18629,N_15319,N_13968);
or U18630 (N_18630,N_13492,N_14203);
nand U18631 (N_18631,N_12471,N_14419);
nor U18632 (N_18632,N_14123,N_15387);
nand U18633 (N_18633,N_15905,N_15600);
nand U18634 (N_18634,N_12557,N_15944);
nand U18635 (N_18635,N_14484,N_14561);
nor U18636 (N_18636,N_13071,N_12202);
nor U18637 (N_18637,N_14051,N_14092);
and U18638 (N_18638,N_12899,N_12205);
or U18639 (N_18639,N_13848,N_13207);
or U18640 (N_18640,N_15530,N_13566);
nor U18641 (N_18641,N_14924,N_14634);
or U18642 (N_18642,N_14726,N_12229);
nand U18643 (N_18643,N_15471,N_14663);
or U18644 (N_18644,N_13756,N_12562);
or U18645 (N_18645,N_15907,N_13379);
and U18646 (N_18646,N_14621,N_14716);
or U18647 (N_18647,N_14496,N_13672);
or U18648 (N_18648,N_14106,N_15257);
and U18649 (N_18649,N_13267,N_13962);
xnor U18650 (N_18650,N_15267,N_12231);
and U18651 (N_18651,N_14596,N_15183);
and U18652 (N_18652,N_15923,N_13211);
nor U18653 (N_18653,N_14796,N_14358);
or U18654 (N_18654,N_14363,N_12127);
nand U18655 (N_18655,N_13472,N_13558);
and U18656 (N_18656,N_13690,N_13826);
or U18657 (N_18657,N_13649,N_12267);
and U18658 (N_18658,N_13583,N_14155);
nor U18659 (N_18659,N_15814,N_14838);
and U18660 (N_18660,N_14042,N_15044);
nor U18661 (N_18661,N_13544,N_12264);
or U18662 (N_18662,N_12744,N_13018);
and U18663 (N_18663,N_15916,N_15253);
nand U18664 (N_18664,N_14675,N_12986);
nand U18665 (N_18665,N_12200,N_15086);
or U18666 (N_18666,N_13745,N_15901);
nor U18667 (N_18667,N_15450,N_13550);
or U18668 (N_18668,N_15811,N_13925);
and U18669 (N_18669,N_15570,N_12501);
nor U18670 (N_18670,N_14136,N_15149);
nor U18671 (N_18671,N_12517,N_15713);
nor U18672 (N_18672,N_13959,N_14916);
and U18673 (N_18673,N_13028,N_13627);
or U18674 (N_18674,N_13699,N_15766);
and U18675 (N_18675,N_13118,N_15353);
nor U18676 (N_18676,N_12425,N_14826);
nand U18677 (N_18677,N_15759,N_15068);
or U18678 (N_18678,N_14873,N_12824);
and U18679 (N_18679,N_14229,N_14590);
xnor U18680 (N_18680,N_13366,N_15743);
xnor U18681 (N_18681,N_15144,N_13126);
nor U18682 (N_18682,N_14121,N_13434);
and U18683 (N_18683,N_13193,N_12824);
or U18684 (N_18684,N_13866,N_13356);
and U18685 (N_18685,N_14259,N_15622);
nor U18686 (N_18686,N_15386,N_14929);
nand U18687 (N_18687,N_15836,N_12833);
nor U18688 (N_18688,N_13021,N_12480);
or U18689 (N_18689,N_15294,N_15125);
or U18690 (N_18690,N_15874,N_14829);
nand U18691 (N_18691,N_14113,N_15144);
nor U18692 (N_18692,N_14462,N_15834);
and U18693 (N_18693,N_13780,N_15641);
nor U18694 (N_18694,N_15145,N_14468);
nor U18695 (N_18695,N_13903,N_13835);
nand U18696 (N_18696,N_13041,N_14276);
and U18697 (N_18697,N_13331,N_13484);
nor U18698 (N_18698,N_15593,N_15826);
nor U18699 (N_18699,N_14479,N_13865);
and U18700 (N_18700,N_14166,N_12570);
nand U18701 (N_18701,N_13211,N_13354);
or U18702 (N_18702,N_13385,N_12242);
nor U18703 (N_18703,N_15947,N_12672);
or U18704 (N_18704,N_14233,N_15737);
or U18705 (N_18705,N_14090,N_13424);
or U18706 (N_18706,N_15049,N_12499);
or U18707 (N_18707,N_14930,N_13901);
nand U18708 (N_18708,N_15946,N_14974);
or U18709 (N_18709,N_14291,N_15019);
nor U18710 (N_18710,N_13906,N_15670);
and U18711 (N_18711,N_12363,N_15840);
nand U18712 (N_18712,N_12914,N_13995);
nor U18713 (N_18713,N_13494,N_13124);
nor U18714 (N_18714,N_13454,N_14273);
nor U18715 (N_18715,N_13829,N_12101);
nor U18716 (N_18716,N_15471,N_15586);
nand U18717 (N_18717,N_14661,N_13654);
or U18718 (N_18718,N_13568,N_12678);
or U18719 (N_18719,N_12032,N_15154);
nor U18720 (N_18720,N_12052,N_13457);
nand U18721 (N_18721,N_12529,N_15832);
nand U18722 (N_18722,N_15283,N_13302);
and U18723 (N_18723,N_12463,N_13719);
and U18724 (N_18724,N_14987,N_12525);
or U18725 (N_18725,N_14102,N_14833);
nor U18726 (N_18726,N_12656,N_14139);
and U18727 (N_18727,N_14226,N_14305);
and U18728 (N_18728,N_15805,N_15714);
nand U18729 (N_18729,N_13041,N_13038);
nand U18730 (N_18730,N_14109,N_13414);
nand U18731 (N_18731,N_15364,N_15504);
nand U18732 (N_18732,N_15243,N_12937);
or U18733 (N_18733,N_12348,N_15815);
or U18734 (N_18734,N_13778,N_15661);
or U18735 (N_18735,N_15539,N_12051);
and U18736 (N_18736,N_14002,N_13693);
nor U18737 (N_18737,N_13332,N_14522);
or U18738 (N_18738,N_14841,N_13217);
and U18739 (N_18739,N_14526,N_13593);
nor U18740 (N_18740,N_15768,N_13889);
nand U18741 (N_18741,N_14621,N_13045);
and U18742 (N_18742,N_15982,N_12141);
and U18743 (N_18743,N_15607,N_12986);
nand U18744 (N_18744,N_12964,N_13336);
nand U18745 (N_18745,N_12050,N_13969);
xor U18746 (N_18746,N_14721,N_13376);
nand U18747 (N_18747,N_12433,N_13191);
nor U18748 (N_18748,N_15065,N_15436);
nor U18749 (N_18749,N_13153,N_15657);
or U18750 (N_18750,N_14666,N_13701);
nand U18751 (N_18751,N_15397,N_14628);
or U18752 (N_18752,N_13176,N_12344);
nor U18753 (N_18753,N_13996,N_15002);
xor U18754 (N_18754,N_12489,N_12721);
or U18755 (N_18755,N_14939,N_12410);
nand U18756 (N_18756,N_14074,N_13531);
xnor U18757 (N_18757,N_14970,N_14308);
or U18758 (N_18758,N_15650,N_13636);
nand U18759 (N_18759,N_12237,N_13615);
and U18760 (N_18760,N_13855,N_14107);
and U18761 (N_18761,N_12838,N_13717);
nor U18762 (N_18762,N_13098,N_13559);
nand U18763 (N_18763,N_13848,N_12287);
xnor U18764 (N_18764,N_14922,N_12814);
and U18765 (N_18765,N_14427,N_14141);
nor U18766 (N_18766,N_15631,N_14751);
nand U18767 (N_18767,N_13142,N_15827);
nand U18768 (N_18768,N_12811,N_12107);
and U18769 (N_18769,N_12887,N_14655);
nor U18770 (N_18770,N_14376,N_12766);
or U18771 (N_18771,N_13161,N_15658);
xor U18772 (N_18772,N_15899,N_14409);
or U18773 (N_18773,N_13950,N_14369);
nor U18774 (N_18774,N_14825,N_12158);
or U18775 (N_18775,N_13021,N_13836);
or U18776 (N_18776,N_14799,N_13208);
nand U18777 (N_18777,N_12558,N_14805);
and U18778 (N_18778,N_13411,N_14338);
and U18779 (N_18779,N_14804,N_12758);
nor U18780 (N_18780,N_13919,N_12416);
or U18781 (N_18781,N_13601,N_12011);
or U18782 (N_18782,N_14288,N_14983);
nand U18783 (N_18783,N_12977,N_15503);
nor U18784 (N_18784,N_15676,N_12331);
nand U18785 (N_18785,N_14186,N_14062);
or U18786 (N_18786,N_12108,N_14301);
nor U18787 (N_18787,N_15668,N_12388);
nor U18788 (N_18788,N_14310,N_15732);
nor U18789 (N_18789,N_12776,N_14572);
or U18790 (N_18790,N_13547,N_15307);
or U18791 (N_18791,N_14003,N_14052);
and U18792 (N_18792,N_14193,N_12936);
or U18793 (N_18793,N_14390,N_14511);
nor U18794 (N_18794,N_15539,N_12540);
or U18795 (N_18795,N_12827,N_13918);
nand U18796 (N_18796,N_15275,N_14227);
nand U18797 (N_18797,N_14715,N_12900);
nand U18798 (N_18798,N_12323,N_14560);
or U18799 (N_18799,N_15525,N_13725);
nand U18800 (N_18800,N_12542,N_13680);
and U18801 (N_18801,N_14499,N_13951);
and U18802 (N_18802,N_12531,N_13728);
nor U18803 (N_18803,N_14961,N_14663);
xor U18804 (N_18804,N_14192,N_14496);
and U18805 (N_18805,N_13333,N_13272);
nor U18806 (N_18806,N_13509,N_12672);
nand U18807 (N_18807,N_15376,N_15583);
nand U18808 (N_18808,N_15492,N_12815);
xor U18809 (N_18809,N_12363,N_13122);
or U18810 (N_18810,N_13156,N_15667);
nor U18811 (N_18811,N_12985,N_14262);
and U18812 (N_18812,N_14657,N_14840);
and U18813 (N_18813,N_13353,N_15175);
or U18814 (N_18814,N_13763,N_14961);
and U18815 (N_18815,N_13893,N_13939);
and U18816 (N_18816,N_15884,N_12215);
and U18817 (N_18817,N_15021,N_15709);
and U18818 (N_18818,N_14473,N_12379);
nand U18819 (N_18819,N_14220,N_13368);
nand U18820 (N_18820,N_14217,N_14008);
and U18821 (N_18821,N_12954,N_12966);
and U18822 (N_18822,N_15899,N_13896);
xnor U18823 (N_18823,N_14187,N_15930);
nor U18824 (N_18824,N_14792,N_12286);
nor U18825 (N_18825,N_14403,N_12555);
nor U18826 (N_18826,N_14253,N_12022);
nand U18827 (N_18827,N_15442,N_15555);
or U18828 (N_18828,N_12731,N_14713);
and U18829 (N_18829,N_15288,N_12120);
or U18830 (N_18830,N_12214,N_14644);
nand U18831 (N_18831,N_14853,N_12217);
nand U18832 (N_18832,N_14635,N_15461);
nand U18833 (N_18833,N_13627,N_14397);
and U18834 (N_18834,N_13736,N_12713);
or U18835 (N_18835,N_13135,N_14362);
or U18836 (N_18836,N_14440,N_13218);
nand U18837 (N_18837,N_13766,N_14862);
nand U18838 (N_18838,N_14770,N_12762);
and U18839 (N_18839,N_12755,N_14844);
or U18840 (N_18840,N_12459,N_14193);
nand U18841 (N_18841,N_13867,N_15173);
nor U18842 (N_18842,N_12481,N_13809);
and U18843 (N_18843,N_12343,N_12650);
and U18844 (N_18844,N_14774,N_14507);
and U18845 (N_18845,N_15299,N_12335);
nor U18846 (N_18846,N_12154,N_15548);
nor U18847 (N_18847,N_14833,N_12095);
nand U18848 (N_18848,N_15344,N_13555);
nand U18849 (N_18849,N_14342,N_15597);
and U18850 (N_18850,N_12717,N_12184);
nand U18851 (N_18851,N_13880,N_13445);
xor U18852 (N_18852,N_14087,N_14477);
nor U18853 (N_18853,N_13597,N_14082);
nand U18854 (N_18854,N_13082,N_14533);
nor U18855 (N_18855,N_13989,N_13373);
and U18856 (N_18856,N_14678,N_14481);
nor U18857 (N_18857,N_13771,N_14575);
nand U18858 (N_18858,N_15186,N_12809);
or U18859 (N_18859,N_14613,N_15460);
nor U18860 (N_18860,N_12726,N_15116);
xnor U18861 (N_18861,N_14639,N_13214);
nor U18862 (N_18862,N_15051,N_12414);
nand U18863 (N_18863,N_14227,N_14963);
nand U18864 (N_18864,N_14610,N_12626);
nor U18865 (N_18865,N_12472,N_13387);
nand U18866 (N_18866,N_13546,N_13878);
and U18867 (N_18867,N_14767,N_14876);
or U18868 (N_18868,N_12213,N_14419);
and U18869 (N_18869,N_14451,N_12225);
and U18870 (N_18870,N_14692,N_15609);
or U18871 (N_18871,N_15974,N_13698);
and U18872 (N_18872,N_13243,N_13618);
nand U18873 (N_18873,N_14147,N_15490);
nand U18874 (N_18874,N_12970,N_15452);
nand U18875 (N_18875,N_12233,N_14373);
nor U18876 (N_18876,N_14162,N_15727);
and U18877 (N_18877,N_12559,N_15897);
nand U18878 (N_18878,N_14368,N_13188);
nand U18879 (N_18879,N_15569,N_12881);
and U18880 (N_18880,N_14474,N_14271);
xor U18881 (N_18881,N_14530,N_13486);
or U18882 (N_18882,N_15183,N_14198);
and U18883 (N_18883,N_15053,N_13992);
or U18884 (N_18884,N_13086,N_14848);
nor U18885 (N_18885,N_15491,N_13040);
and U18886 (N_18886,N_12352,N_15705);
and U18887 (N_18887,N_12280,N_14516);
nor U18888 (N_18888,N_14542,N_12249);
nor U18889 (N_18889,N_12257,N_15970);
and U18890 (N_18890,N_15684,N_12886);
and U18891 (N_18891,N_12458,N_15858);
and U18892 (N_18892,N_13623,N_14722);
or U18893 (N_18893,N_15802,N_13172);
nor U18894 (N_18894,N_14046,N_14011);
nor U18895 (N_18895,N_14147,N_13562);
nor U18896 (N_18896,N_13603,N_14573);
nand U18897 (N_18897,N_12847,N_12955);
and U18898 (N_18898,N_14254,N_14986);
and U18899 (N_18899,N_13764,N_12108);
and U18900 (N_18900,N_12581,N_14366);
nand U18901 (N_18901,N_14833,N_14681);
and U18902 (N_18902,N_13077,N_15971);
nand U18903 (N_18903,N_14126,N_12787);
xor U18904 (N_18904,N_14068,N_12295);
nand U18905 (N_18905,N_14756,N_13961);
and U18906 (N_18906,N_13369,N_12350);
nor U18907 (N_18907,N_12114,N_13201);
and U18908 (N_18908,N_12766,N_14774);
and U18909 (N_18909,N_14617,N_12344);
nor U18910 (N_18910,N_15588,N_14920);
or U18911 (N_18911,N_15510,N_12873);
nor U18912 (N_18912,N_12674,N_12961);
nand U18913 (N_18913,N_12432,N_12692);
xor U18914 (N_18914,N_12702,N_13334);
nand U18915 (N_18915,N_14177,N_12798);
or U18916 (N_18916,N_12009,N_14997);
or U18917 (N_18917,N_12928,N_15133);
nand U18918 (N_18918,N_13370,N_14586);
or U18919 (N_18919,N_14590,N_15814);
nand U18920 (N_18920,N_12145,N_15077);
xnor U18921 (N_18921,N_14679,N_12051);
nor U18922 (N_18922,N_15022,N_12502);
or U18923 (N_18923,N_12821,N_12361);
nand U18924 (N_18924,N_15297,N_12819);
nand U18925 (N_18925,N_14633,N_12175);
nand U18926 (N_18926,N_12275,N_15427);
xor U18927 (N_18927,N_13571,N_15728);
nor U18928 (N_18928,N_14213,N_13673);
and U18929 (N_18929,N_15767,N_14136);
and U18930 (N_18930,N_15995,N_14099);
or U18931 (N_18931,N_13447,N_12619);
nor U18932 (N_18932,N_14456,N_15175);
and U18933 (N_18933,N_13379,N_14396);
or U18934 (N_18934,N_15099,N_13513);
nor U18935 (N_18935,N_15394,N_13005);
nand U18936 (N_18936,N_12718,N_13278);
nand U18937 (N_18937,N_13389,N_15712);
nand U18938 (N_18938,N_14289,N_14915);
nand U18939 (N_18939,N_14433,N_14889);
xor U18940 (N_18940,N_15477,N_14408);
nor U18941 (N_18941,N_14355,N_15864);
or U18942 (N_18942,N_12814,N_12164);
nor U18943 (N_18943,N_15872,N_15937);
nand U18944 (N_18944,N_13619,N_12718);
and U18945 (N_18945,N_12944,N_12970);
and U18946 (N_18946,N_14424,N_12581);
nor U18947 (N_18947,N_15877,N_14963);
nor U18948 (N_18948,N_13650,N_14257);
nor U18949 (N_18949,N_15655,N_13676);
nand U18950 (N_18950,N_13159,N_15416);
or U18951 (N_18951,N_12231,N_15451);
nand U18952 (N_18952,N_13329,N_13962);
nor U18953 (N_18953,N_13071,N_12023);
nand U18954 (N_18954,N_12684,N_14084);
or U18955 (N_18955,N_15331,N_13373);
nor U18956 (N_18956,N_14081,N_13954);
nand U18957 (N_18957,N_15868,N_15992);
nand U18958 (N_18958,N_15486,N_15428);
nand U18959 (N_18959,N_15852,N_14524);
nor U18960 (N_18960,N_15486,N_15974);
nor U18961 (N_18961,N_15891,N_15754);
nand U18962 (N_18962,N_15857,N_12302);
and U18963 (N_18963,N_12067,N_12904);
nor U18964 (N_18964,N_15744,N_14127);
nand U18965 (N_18965,N_12759,N_12769);
or U18966 (N_18966,N_15337,N_13858);
nor U18967 (N_18967,N_15122,N_14381);
or U18968 (N_18968,N_12482,N_15505);
nor U18969 (N_18969,N_12878,N_12412);
xor U18970 (N_18970,N_14232,N_13732);
and U18971 (N_18971,N_12722,N_15362);
or U18972 (N_18972,N_13063,N_13958);
nor U18973 (N_18973,N_15781,N_14892);
and U18974 (N_18974,N_12709,N_13512);
nor U18975 (N_18975,N_13730,N_14788);
nand U18976 (N_18976,N_12464,N_14429);
nor U18977 (N_18977,N_12321,N_15574);
or U18978 (N_18978,N_14366,N_12983);
and U18979 (N_18979,N_14478,N_15443);
nor U18980 (N_18980,N_12593,N_15695);
or U18981 (N_18981,N_12433,N_12111);
and U18982 (N_18982,N_14848,N_13774);
nand U18983 (N_18983,N_12983,N_14395);
or U18984 (N_18984,N_12689,N_13074);
nand U18985 (N_18985,N_12661,N_12846);
nor U18986 (N_18986,N_15343,N_12317);
or U18987 (N_18987,N_14719,N_15124);
or U18988 (N_18988,N_13916,N_12043);
nand U18989 (N_18989,N_14369,N_14181);
and U18990 (N_18990,N_14657,N_13548);
or U18991 (N_18991,N_12885,N_13119);
xnor U18992 (N_18992,N_14527,N_15378);
nor U18993 (N_18993,N_14329,N_13250);
nor U18994 (N_18994,N_13925,N_15761);
or U18995 (N_18995,N_15197,N_12144);
nor U18996 (N_18996,N_12369,N_14138);
nor U18997 (N_18997,N_12310,N_14161);
nor U18998 (N_18998,N_12604,N_14930);
nand U18999 (N_18999,N_12111,N_15257);
nand U19000 (N_19000,N_14351,N_15330);
or U19001 (N_19001,N_14246,N_15607);
nand U19002 (N_19002,N_14230,N_13627);
and U19003 (N_19003,N_12026,N_13663);
nor U19004 (N_19004,N_12210,N_14360);
nor U19005 (N_19005,N_14724,N_15838);
and U19006 (N_19006,N_13960,N_13885);
or U19007 (N_19007,N_13261,N_15284);
or U19008 (N_19008,N_14882,N_13307);
and U19009 (N_19009,N_13729,N_12125);
or U19010 (N_19010,N_14542,N_14946);
nor U19011 (N_19011,N_14687,N_15159);
xor U19012 (N_19012,N_13168,N_13448);
nor U19013 (N_19013,N_14429,N_15996);
nor U19014 (N_19014,N_13778,N_15222);
or U19015 (N_19015,N_14095,N_13918);
and U19016 (N_19016,N_15972,N_12302);
nand U19017 (N_19017,N_14586,N_15883);
nand U19018 (N_19018,N_13944,N_15778);
nand U19019 (N_19019,N_12747,N_12168);
or U19020 (N_19020,N_12549,N_15584);
nand U19021 (N_19021,N_13387,N_13187);
xor U19022 (N_19022,N_13971,N_13105);
nand U19023 (N_19023,N_15417,N_13552);
nand U19024 (N_19024,N_15280,N_14311);
nor U19025 (N_19025,N_14613,N_12697);
nand U19026 (N_19026,N_14699,N_15887);
nand U19027 (N_19027,N_12547,N_13893);
nand U19028 (N_19028,N_14177,N_15223);
nand U19029 (N_19029,N_15683,N_12928);
nand U19030 (N_19030,N_15933,N_12746);
or U19031 (N_19031,N_12261,N_12846);
and U19032 (N_19032,N_12373,N_14414);
nor U19033 (N_19033,N_12684,N_12458);
nand U19034 (N_19034,N_14124,N_15818);
xnor U19035 (N_19035,N_14069,N_13434);
or U19036 (N_19036,N_12894,N_15587);
and U19037 (N_19037,N_13631,N_15077);
or U19038 (N_19038,N_12198,N_13683);
or U19039 (N_19039,N_13407,N_13874);
nand U19040 (N_19040,N_15121,N_12779);
nand U19041 (N_19041,N_15414,N_12807);
nand U19042 (N_19042,N_14070,N_12642);
or U19043 (N_19043,N_15860,N_12834);
xor U19044 (N_19044,N_13546,N_13622);
and U19045 (N_19045,N_12610,N_14881);
nor U19046 (N_19046,N_14307,N_15354);
nand U19047 (N_19047,N_14044,N_14885);
nand U19048 (N_19048,N_12171,N_15915);
nor U19049 (N_19049,N_14952,N_15780);
nor U19050 (N_19050,N_12086,N_15310);
nand U19051 (N_19051,N_12408,N_12501);
nand U19052 (N_19052,N_14032,N_14606);
and U19053 (N_19053,N_15673,N_15241);
nor U19054 (N_19054,N_13983,N_15493);
nand U19055 (N_19055,N_12060,N_15363);
or U19056 (N_19056,N_14290,N_15955);
nand U19057 (N_19057,N_12151,N_12412);
nand U19058 (N_19058,N_12972,N_14694);
and U19059 (N_19059,N_14708,N_13356);
and U19060 (N_19060,N_12098,N_12703);
nand U19061 (N_19061,N_12933,N_13789);
nand U19062 (N_19062,N_12031,N_13063);
and U19063 (N_19063,N_15936,N_14599);
nand U19064 (N_19064,N_12295,N_13047);
or U19065 (N_19065,N_14520,N_15305);
and U19066 (N_19066,N_13229,N_13495);
xor U19067 (N_19067,N_15547,N_13410);
nor U19068 (N_19068,N_13720,N_15155);
or U19069 (N_19069,N_15208,N_15857);
nand U19070 (N_19070,N_14924,N_15695);
or U19071 (N_19071,N_12525,N_13404);
nor U19072 (N_19072,N_15513,N_12520);
or U19073 (N_19073,N_15287,N_12422);
nand U19074 (N_19074,N_13477,N_15831);
and U19075 (N_19075,N_14759,N_13241);
and U19076 (N_19076,N_12549,N_13438);
and U19077 (N_19077,N_13129,N_15525);
and U19078 (N_19078,N_15824,N_14779);
xor U19079 (N_19079,N_14664,N_13387);
or U19080 (N_19080,N_14212,N_15714);
xor U19081 (N_19081,N_15923,N_15368);
nand U19082 (N_19082,N_12747,N_14977);
or U19083 (N_19083,N_13561,N_12732);
nand U19084 (N_19084,N_14056,N_12303);
xor U19085 (N_19085,N_15349,N_15341);
nand U19086 (N_19086,N_12694,N_13442);
nor U19087 (N_19087,N_12710,N_14785);
or U19088 (N_19088,N_15380,N_12748);
nor U19089 (N_19089,N_15787,N_15139);
nor U19090 (N_19090,N_13175,N_13115);
and U19091 (N_19091,N_12512,N_14008);
nor U19092 (N_19092,N_12409,N_15337);
and U19093 (N_19093,N_12425,N_15193);
or U19094 (N_19094,N_15816,N_14197);
nand U19095 (N_19095,N_15091,N_14674);
or U19096 (N_19096,N_15805,N_12032);
or U19097 (N_19097,N_12152,N_13083);
nor U19098 (N_19098,N_14128,N_14391);
nor U19099 (N_19099,N_14941,N_13780);
nand U19100 (N_19100,N_14567,N_14243);
and U19101 (N_19101,N_15068,N_15241);
and U19102 (N_19102,N_13252,N_13067);
nand U19103 (N_19103,N_14278,N_12937);
and U19104 (N_19104,N_14088,N_12609);
nand U19105 (N_19105,N_15864,N_15205);
nor U19106 (N_19106,N_13885,N_15100);
nor U19107 (N_19107,N_12966,N_13535);
or U19108 (N_19108,N_15766,N_12836);
nand U19109 (N_19109,N_13685,N_15497);
nand U19110 (N_19110,N_15557,N_12273);
nand U19111 (N_19111,N_14788,N_12035);
nor U19112 (N_19112,N_14162,N_14958);
and U19113 (N_19113,N_12777,N_13997);
or U19114 (N_19114,N_13287,N_15980);
or U19115 (N_19115,N_13930,N_13036);
nor U19116 (N_19116,N_14257,N_13628);
nand U19117 (N_19117,N_15795,N_15476);
nand U19118 (N_19118,N_14708,N_12710);
nor U19119 (N_19119,N_15577,N_14426);
nor U19120 (N_19120,N_12869,N_14905);
nor U19121 (N_19121,N_14100,N_14376);
or U19122 (N_19122,N_15892,N_14510);
nor U19123 (N_19123,N_14280,N_15119);
and U19124 (N_19124,N_15584,N_14264);
nor U19125 (N_19125,N_12438,N_14521);
or U19126 (N_19126,N_15682,N_14152);
or U19127 (N_19127,N_12319,N_13397);
or U19128 (N_19128,N_12731,N_13880);
and U19129 (N_19129,N_12427,N_14285);
nand U19130 (N_19130,N_15041,N_13669);
nor U19131 (N_19131,N_12959,N_14547);
nor U19132 (N_19132,N_12831,N_13586);
nand U19133 (N_19133,N_14781,N_14811);
nand U19134 (N_19134,N_15571,N_14279);
nor U19135 (N_19135,N_12989,N_15385);
and U19136 (N_19136,N_12706,N_12204);
nand U19137 (N_19137,N_13555,N_12673);
nor U19138 (N_19138,N_13250,N_12667);
nor U19139 (N_19139,N_12791,N_13514);
nand U19140 (N_19140,N_12803,N_15233);
nand U19141 (N_19141,N_14805,N_12830);
nor U19142 (N_19142,N_13804,N_13108);
nand U19143 (N_19143,N_14892,N_14168);
nand U19144 (N_19144,N_15312,N_14442);
nor U19145 (N_19145,N_12267,N_13941);
xor U19146 (N_19146,N_15938,N_14688);
nor U19147 (N_19147,N_15698,N_15048);
and U19148 (N_19148,N_14171,N_15537);
nor U19149 (N_19149,N_15826,N_13873);
and U19150 (N_19150,N_15582,N_15293);
nand U19151 (N_19151,N_15448,N_15472);
nand U19152 (N_19152,N_13168,N_15374);
nor U19153 (N_19153,N_13996,N_15628);
nor U19154 (N_19154,N_12575,N_14992);
and U19155 (N_19155,N_15358,N_14164);
and U19156 (N_19156,N_13513,N_13862);
nor U19157 (N_19157,N_12927,N_12985);
nor U19158 (N_19158,N_15747,N_14198);
or U19159 (N_19159,N_15030,N_12883);
and U19160 (N_19160,N_12695,N_12013);
and U19161 (N_19161,N_12012,N_14633);
nor U19162 (N_19162,N_14136,N_13298);
or U19163 (N_19163,N_14467,N_14001);
and U19164 (N_19164,N_12954,N_14537);
nor U19165 (N_19165,N_15821,N_15988);
nand U19166 (N_19166,N_14516,N_15204);
nand U19167 (N_19167,N_13463,N_13566);
and U19168 (N_19168,N_13090,N_12669);
nand U19169 (N_19169,N_15184,N_14501);
nor U19170 (N_19170,N_12869,N_13392);
or U19171 (N_19171,N_14712,N_13798);
nor U19172 (N_19172,N_12968,N_13595);
nand U19173 (N_19173,N_14164,N_14938);
and U19174 (N_19174,N_14676,N_15086);
and U19175 (N_19175,N_15908,N_15319);
and U19176 (N_19176,N_15698,N_13544);
and U19177 (N_19177,N_14993,N_13977);
nand U19178 (N_19178,N_13918,N_14345);
nand U19179 (N_19179,N_15615,N_12866);
or U19180 (N_19180,N_15547,N_13371);
nor U19181 (N_19181,N_14042,N_14167);
and U19182 (N_19182,N_14193,N_13348);
and U19183 (N_19183,N_15424,N_15936);
or U19184 (N_19184,N_13210,N_15239);
nor U19185 (N_19185,N_13681,N_14697);
or U19186 (N_19186,N_13984,N_13999);
or U19187 (N_19187,N_15103,N_14340);
or U19188 (N_19188,N_13204,N_13254);
xor U19189 (N_19189,N_14482,N_13782);
and U19190 (N_19190,N_14168,N_13029);
or U19191 (N_19191,N_15437,N_13062);
and U19192 (N_19192,N_14235,N_14035);
or U19193 (N_19193,N_12508,N_13743);
nor U19194 (N_19194,N_15630,N_14927);
and U19195 (N_19195,N_14588,N_15923);
or U19196 (N_19196,N_12030,N_14264);
nand U19197 (N_19197,N_14610,N_12069);
or U19198 (N_19198,N_13767,N_12272);
nor U19199 (N_19199,N_12679,N_15563);
and U19200 (N_19200,N_12514,N_15743);
or U19201 (N_19201,N_13327,N_13520);
nand U19202 (N_19202,N_14556,N_14239);
nor U19203 (N_19203,N_12397,N_13738);
or U19204 (N_19204,N_13356,N_14403);
nor U19205 (N_19205,N_13225,N_15059);
or U19206 (N_19206,N_13349,N_15309);
nor U19207 (N_19207,N_14258,N_14615);
or U19208 (N_19208,N_13963,N_15827);
xnor U19209 (N_19209,N_12828,N_12054);
nand U19210 (N_19210,N_12012,N_14743);
nor U19211 (N_19211,N_13858,N_12899);
nor U19212 (N_19212,N_13219,N_12027);
and U19213 (N_19213,N_12115,N_14847);
and U19214 (N_19214,N_13927,N_14446);
and U19215 (N_19215,N_12561,N_12861);
nor U19216 (N_19216,N_15394,N_12017);
nor U19217 (N_19217,N_13534,N_13880);
or U19218 (N_19218,N_15158,N_13160);
or U19219 (N_19219,N_12020,N_12694);
or U19220 (N_19220,N_12058,N_13454);
and U19221 (N_19221,N_14718,N_12969);
or U19222 (N_19222,N_12788,N_14978);
and U19223 (N_19223,N_14901,N_12326);
and U19224 (N_19224,N_15667,N_14741);
or U19225 (N_19225,N_13160,N_13600);
nand U19226 (N_19226,N_15174,N_14787);
nand U19227 (N_19227,N_13536,N_13431);
and U19228 (N_19228,N_12666,N_14750);
and U19229 (N_19229,N_15269,N_13806);
and U19230 (N_19230,N_13522,N_12941);
nand U19231 (N_19231,N_14652,N_12745);
and U19232 (N_19232,N_14950,N_13783);
or U19233 (N_19233,N_14985,N_12210);
nor U19234 (N_19234,N_14724,N_14026);
or U19235 (N_19235,N_14596,N_12295);
nor U19236 (N_19236,N_12973,N_12837);
and U19237 (N_19237,N_12059,N_14955);
or U19238 (N_19238,N_12603,N_12294);
and U19239 (N_19239,N_13137,N_13319);
nor U19240 (N_19240,N_15878,N_13532);
or U19241 (N_19241,N_12309,N_12073);
and U19242 (N_19242,N_15561,N_15962);
or U19243 (N_19243,N_12979,N_14359);
and U19244 (N_19244,N_14497,N_12985);
nand U19245 (N_19245,N_14237,N_12091);
or U19246 (N_19246,N_15905,N_12491);
nand U19247 (N_19247,N_12169,N_14798);
nor U19248 (N_19248,N_13667,N_12371);
nand U19249 (N_19249,N_13751,N_14913);
and U19250 (N_19250,N_12420,N_14832);
or U19251 (N_19251,N_14388,N_15571);
nor U19252 (N_19252,N_15055,N_15730);
nor U19253 (N_19253,N_15731,N_13856);
nand U19254 (N_19254,N_12640,N_13409);
nor U19255 (N_19255,N_13819,N_13872);
or U19256 (N_19256,N_13850,N_12081);
and U19257 (N_19257,N_15734,N_15403);
and U19258 (N_19258,N_13388,N_15951);
or U19259 (N_19259,N_13426,N_12951);
or U19260 (N_19260,N_15412,N_15282);
nand U19261 (N_19261,N_13313,N_13474);
nand U19262 (N_19262,N_12936,N_12243);
and U19263 (N_19263,N_13758,N_13844);
nand U19264 (N_19264,N_14947,N_13076);
nand U19265 (N_19265,N_15208,N_14260);
nand U19266 (N_19266,N_14928,N_14097);
nand U19267 (N_19267,N_15533,N_13327);
or U19268 (N_19268,N_13905,N_13822);
or U19269 (N_19269,N_12752,N_15871);
nor U19270 (N_19270,N_13338,N_12101);
nor U19271 (N_19271,N_13008,N_15342);
and U19272 (N_19272,N_12356,N_12944);
or U19273 (N_19273,N_15854,N_15315);
nor U19274 (N_19274,N_13248,N_14412);
nor U19275 (N_19275,N_12141,N_12398);
nor U19276 (N_19276,N_15668,N_14666);
nor U19277 (N_19277,N_14996,N_15064);
nor U19278 (N_19278,N_15342,N_12872);
nor U19279 (N_19279,N_13246,N_13036);
nor U19280 (N_19280,N_15022,N_13899);
and U19281 (N_19281,N_13732,N_12571);
or U19282 (N_19282,N_14794,N_15175);
and U19283 (N_19283,N_13975,N_14859);
nand U19284 (N_19284,N_12810,N_15485);
or U19285 (N_19285,N_14756,N_14236);
nor U19286 (N_19286,N_13743,N_13750);
xor U19287 (N_19287,N_14157,N_13998);
nor U19288 (N_19288,N_13734,N_14937);
and U19289 (N_19289,N_13580,N_15533);
or U19290 (N_19290,N_14175,N_13518);
and U19291 (N_19291,N_15252,N_15714);
or U19292 (N_19292,N_12113,N_13732);
nor U19293 (N_19293,N_12433,N_13202);
nand U19294 (N_19294,N_13020,N_12545);
nor U19295 (N_19295,N_14848,N_12357);
nor U19296 (N_19296,N_13048,N_13293);
nand U19297 (N_19297,N_15747,N_15475);
nor U19298 (N_19298,N_12725,N_15405);
xor U19299 (N_19299,N_13672,N_13103);
and U19300 (N_19300,N_13393,N_14616);
and U19301 (N_19301,N_12749,N_15509);
or U19302 (N_19302,N_12746,N_13191);
and U19303 (N_19303,N_15057,N_14574);
nand U19304 (N_19304,N_15928,N_13647);
or U19305 (N_19305,N_14987,N_14457);
and U19306 (N_19306,N_14538,N_13911);
nor U19307 (N_19307,N_13196,N_13861);
or U19308 (N_19308,N_14554,N_12307);
or U19309 (N_19309,N_14262,N_13919);
nor U19310 (N_19310,N_13693,N_13351);
or U19311 (N_19311,N_12994,N_12111);
and U19312 (N_19312,N_14601,N_13615);
and U19313 (N_19313,N_15491,N_12258);
nor U19314 (N_19314,N_15040,N_13772);
or U19315 (N_19315,N_13113,N_14350);
nor U19316 (N_19316,N_13910,N_14030);
and U19317 (N_19317,N_14208,N_12692);
xnor U19318 (N_19318,N_12372,N_15730);
or U19319 (N_19319,N_15739,N_12662);
xor U19320 (N_19320,N_12878,N_15536);
nor U19321 (N_19321,N_13365,N_12244);
nand U19322 (N_19322,N_14810,N_14174);
nor U19323 (N_19323,N_13315,N_15371);
or U19324 (N_19324,N_15423,N_15056);
or U19325 (N_19325,N_13354,N_14168);
and U19326 (N_19326,N_12090,N_12807);
nand U19327 (N_19327,N_14127,N_15862);
or U19328 (N_19328,N_12373,N_13737);
nand U19329 (N_19329,N_12947,N_12137);
or U19330 (N_19330,N_14713,N_12031);
nand U19331 (N_19331,N_15488,N_14629);
nand U19332 (N_19332,N_12128,N_15418);
nand U19333 (N_19333,N_13150,N_12117);
nand U19334 (N_19334,N_15595,N_12071);
nand U19335 (N_19335,N_15246,N_15317);
nor U19336 (N_19336,N_12057,N_13471);
and U19337 (N_19337,N_12812,N_14017);
or U19338 (N_19338,N_14954,N_12549);
nor U19339 (N_19339,N_15467,N_14137);
nand U19340 (N_19340,N_12295,N_15795);
nand U19341 (N_19341,N_14738,N_14601);
and U19342 (N_19342,N_12633,N_14129);
and U19343 (N_19343,N_13694,N_12222);
and U19344 (N_19344,N_14364,N_12001);
and U19345 (N_19345,N_12523,N_15226);
nand U19346 (N_19346,N_15591,N_12750);
and U19347 (N_19347,N_13497,N_12849);
and U19348 (N_19348,N_13211,N_12385);
or U19349 (N_19349,N_15269,N_14091);
or U19350 (N_19350,N_13066,N_12497);
or U19351 (N_19351,N_12226,N_15177);
or U19352 (N_19352,N_14521,N_15656);
nor U19353 (N_19353,N_12549,N_13008);
nor U19354 (N_19354,N_15478,N_15024);
and U19355 (N_19355,N_14905,N_15161);
or U19356 (N_19356,N_12440,N_14814);
nand U19357 (N_19357,N_12593,N_12479);
or U19358 (N_19358,N_15857,N_15644);
and U19359 (N_19359,N_13121,N_13962);
nor U19360 (N_19360,N_14891,N_13909);
or U19361 (N_19361,N_12920,N_14911);
or U19362 (N_19362,N_15888,N_15073);
or U19363 (N_19363,N_14247,N_13269);
or U19364 (N_19364,N_12378,N_14573);
or U19365 (N_19365,N_13729,N_14435);
or U19366 (N_19366,N_13992,N_15396);
or U19367 (N_19367,N_12105,N_12199);
xnor U19368 (N_19368,N_15233,N_15640);
nand U19369 (N_19369,N_15268,N_14707);
or U19370 (N_19370,N_13293,N_14641);
nor U19371 (N_19371,N_13788,N_13125);
nor U19372 (N_19372,N_14334,N_12981);
nor U19373 (N_19373,N_15918,N_15311);
xor U19374 (N_19374,N_14066,N_14683);
nand U19375 (N_19375,N_13876,N_14581);
and U19376 (N_19376,N_12387,N_13612);
xor U19377 (N_19377,N_15063,N_15994);
and U19378 (N_19378,N_14480,N_14547);
and U19379 (N_19379,N_13918,N_12344);
nand U19380 (N_19380,N_14466,N_15903);
and U19381 (N_19381,N_12460,N_15255);
and U19382 (N_19382,N_13039,N_12473);
or U19383 (N_19383,N_15220,N_15324);
and U19384 (N_19384,N_12002,N_15762);
nand U19385 (N_19385,N_13138,N_14155);
nand U19386 (N_19386,N_14790,N_15679);
nand U19387 (N_19387,N_15051,N_13225);
nor U19388 (N_19388,N_14075,N_13159);
and U19389 (N_19389,N_12658,N_12940);
nor U19390 (N_19390,N_12954,N_15616);
and U19391 (N_19391,N_13999,N_14096);
and U19392 (N_19392,N_15441,N_15072);
and U19393 (N_19393,N_13156,N_15269);
and U19394 (N_19394,N_12731,N_12255);
or U19395 (N_19395,N_14237,N_15042);
or U19396 (N_19396,N_12179,N_14951);
xor U19397 (N_19397,N_13997,N_12856);
nor U19398 (N_19398,N_14779,N_14246);
nor U19399 (N_19399,N_13182,N_12701);
xnor U19400 (N_19400,N_14048,N_15915);
nor U19401 (N_19401,N_12606,N_13318);
nor U19402 (N_19402,N_14319,N_12527);
nor U19403 (N_19403,N_14206,N_12592);
nand U19404 (N_19404,N_14033,N_14167);
and U19405 (N_19405,N_15185,N_12914);
nand U19406 (N_19406,N_14842,N_12645);
or U19407 (N_19407,N_15531,N_13021);
nor U19408 (N_19408,N_13574,N_15408);
nor U19409 (N_19409,N_14332,N_13800);
nor U19410 (N_19410,N_15756,N_14603);
xnor U19411 (N_19411,N_14893,N_15070);
or U19412 (N_19412,N_14413,N_13379);
or U19413 (N_19413,N_13575,N_12474);
and U19414 (N_19414,N_15389,N_12851);
and U19415 (N_19415,N_13381,N_15534);
nand U19416 (N_19416,N_13495,N_13546);
and U19417 (N_19417,N_12361,N_12053);
nor U19418 (N_19418,N_12004,N_15277);
xnor U19419 (N_19419,N_13431,N_15308);
and U19420 (N_19420,N_12084,N_15725);
nand U19421 (N_19421,N_15500,N_15138);
or U19422 (N_19422,N_13153,N_14727);
nor U19423 (N_19423,N_15942,N_12369);
nand U19424 (N_19424,N_13503,N_15240);
and U19425 (N_19425,N_15300,N_12259);
and U19426 (N_19426,N_12739,N_13967);
xor U19427 (N_19427,N_15260,N_12293);
nand U19428 (N_19428,N_12901,N_14768);
or U19429 (N_19429,N_13503,N_13173);
nor U19430 (N_19430,N_14654,N_12487);
or U19431 (N_19431,N_12414,N_13491);
or U19432 (N_19432,N_15028,N_12335);
nand U19433 (N_19433,N_13561,N_15055);
or U19434 (N_19434,N_12584,N_13028);
nand U19435 (N_19435,N_14064,N_13921);
nor U19436 (N_19436,N_13969,N_14238);
or U19437 (N_19437,N_15437,N_14751);
and U19438 (N_19438,N_14553,N_12085);
xor U19439 (N_19439,N_15461,N_15381);
nand U19440 (N_19440,N_15187,N_12905);
nand U19441 (N_19441,N_15243,N_12865);
and U19442 (N_19442,N_15669,N_12911);
nand U19443 (N_19443,N_15158,N_13715);
and U19444 (N_19444,N_13668,N_14938);
nand U19445 (N_19445,N_14560,N_12380);
xnor U19446 (N_19446,N_13165,N_15138);
and U19447 (N_19447,N_13719,N_13454);
nor U19448 (N_19448,N_15683,N_12399);
nand U19449 (N_19449,N_13561,N_15930);
nor U19450 (N_19450,N_14739,N_15143);
and U19451 (N_19451,N_15582,N_13094);
or U19452 (N_19452,N_12396,N_14343);
or U19453 (N_19453,N_14413,N_14634);
or U19454 (N_19454,N_12860,N_12103);
nor U19455 (N_19455,N_14321,N_14483);
nand U19456 (N_19456,N_14316,N_12764);
nand U19457 (N_19457,N_15504,N_12557);
and U19458 (N_19458,N_15299,N_14160);
or U19459 (N_19459,N_13424,N_13558);
and U19460 (N_19460,N_13569,N_12820);
and U19461 (N_19461,N_13087,N_14163);
or U19462 (N_19462,N_15569,N_14757);
or U19463 (N_19463,N_15077,N_13240);
nor U19464 (N_19464,N_12663,N_12947);
nor U19465 (N_19465,N_15204,N_14827);
xnor U19466 (N_19466,N_14293,N_14503);
or U19467 (N_19467,N_14239,N_15993);
nand U19468 (N_19468,N_14592,N_15974);
and U19469 (N_19469,N_14476,N_14251);
nor U19470 (N_19470,N_12847,N_15768);
nand U19471 (N_19471,N_14987,N_14580);
and U19472 (N_19472,N_12772,N_12068);
xnor U19473 (N_19473,N_14782,N_15124);
or U19474 (N_19474,N_15661,N_15848);
and U19475 (N_19475,N_15198,N_15388);
nand U19476 (N_19476,N_13903,N_13956);
nand U19477 (N_19477,N_15442,N_12970);
nand U19478 (N_19478,N_13693,N_12161);
nor U19479 (N_19479,N_14497,N_15117);
nor U19480 (N_19480,N_13759,N_13502);
nand U19481 (N_19481,N_12814,N_14985);
or U19482 (N_19482,N_15502,N_14804);
or U19483 (N_19483,N_15479,N_14153);
nor U19484 (N_19484,N_12082,N_15773);
nor U19485 (N_19485,N_12503,N_13726);
or U19486 (N_19486,N_14178,N_13869);
and U19487 (N_19487,N_15004,N_12064);
and U19488 (N_19488,N_13829,N_14672);
nor U19489 (N_19489,N_13804,N_15558);
nand U19490 (N_19490,N_15946,N_12686);
and U19491 (N_19491,N_13354,N_12747);
nand U19492 (N_19492,N_12692,N_12531);
or U19493 (N_19493,N_12396,N_13165);
or U19494 (N_19494,N_14092,N_12617);
or U19495 (N_19495,N_12059,N_13026);
nor U19496 (N_19496,N_12723,N_13618);
or U19497 (N_19497,N_12272,N_13582);
nor U19498 (N_19498,N_15994,N_15265);
nand U19499 (N_19499,N_15676,N_14503);
nand U19500 (N_19500,N_14680,N_15963);
nor U19501 (N_19501,N_13494,N_14421);
or U19502 (N_19502,N_14679,N_14725);
xnor U19503 (N_19503,N_14022,N_13141);
and U19504 (N_19504,N_15068,N_14434);
or U19505 (N_19505,N_13790,N_15830);
and U19506 (N_19506,N_14979,N_15367);
nand U19507 (N_19507,N_14484,N_14608);
or U19508 (N_19508,N_15985,N_15466);
nand U19509 (N_19509,N_14106,N_12370);
nand U19510 (N_19510,N_12332,N_13990);
or U19511 (N_19511,N_15235,N_13391);
or U19512 (N_19512,N_13953,N_14204);
nand U19513 (N_19513,N_13361,N_14075);
nand U19514 (N_19514,N_12238,N_13653);
nand U19515 (N_19515,N_13649,N_15994);
nor U19516 (N_19516,N_13752,N_15344);
and U19517 (N_19517,N_15808,N_14281);
nor U19518 (N_19518,N_14356,N_15597);
nor U19519 (N_19519,N_12045,N_14393);
and U19520 (N_19520,N_14659,N_14386);
or U19521 (N_19521,N_14278,N_12885);
nor U19522 (N_19522,N_15659,N_13950);
nor U19523 (N_19523,N_13503,N_14164);
nand U19524 (N_19524,N_12378,N_14525);
and U19525 (N_19525,N_12932,N_15746);
and U19526 (N_19526,N_12748,N_12083);
and U19527 (N_19527,N_15064,N_15849);
and U19528 (N_19528,N_15913,N_12750);
and U19529 (N_19529,N_14005,N_13964);
nor U19530 (N_19530,N_15106,N_13581);
nand U19531 (N_19531,N_14893,N_14398);
or U19532 (N_19532,N_14095,N_12226);
nor U19533 (N_19533,N_15548,N_13211);
nor U19534 (N_19534,N_12036,N_15234);
and U19535 (N_19535,N_13766,N_13210);
or U19536 (N_19536,N_15758,N_13772);
or U19537 (N_19537,N_13197,N_14243);
or U19538 (N_19538,N_14806,N_13748);
or U19539 (N_19539,N_12275,N_14948);
nand U19540 (N_19540,N_14803,N_13967);
and U19541 (N_19541,N_13157,N_14662);
and U19542 (N_19542,N_14807,N_15217);
and U19543 (N_19543,N_12192,N_15977);
or U19544 (N_19544,N_14645,N_14427);
nor U19545 (N_19545,N_15291,N_12776);
nor U19546 (N_19546,N_12916,N_14731);
and U19547 (N_19547,N_13622,N_14053);
xor U19548 (N_19548,N_12983,N_12175);
and U19549 (N_19549,N_15632,N_12998);
and U19550 (N_19550,N_12203,N_12270);
nand U19551 (N_19551,N_15090,N_12682);
or U19552 (N_19552,N_14515,N_14299);
nor U19553 (N_19553,N_14763,N_12993);
and U19554 (N_19554,N_15739,N_15506);
nand U19555 (N_19555,N_12199,N_12669);
xor U19556 (N_19556,N_12256,N_14555);
nor U19557 (N_19557,N_14146,N_14931);
or U19558 (N_19558,N_14029,N_13018);
and U19559 (N_19559,N_15044,N_14953);
or U19560 (N_19560,N_15557,N_12085);
and U19561 (N_19561,N_13232,N_12983);
or U19562 (N_19562,N_13270,N_15851);
and U19563 (N_19563,N_12847,N_14839);
nand U19564 (N_19564,N_14276,N_15807);
or U19565 (N_19565,N_14470,N_13009);
nor U19566 (N_19566,N_14327,N_12707);
xnor U19567 (N_19567,N_15819,N_12592);
or U19568 (N_19568,N_14910,N_13199);
nor U19569 (N_19569,N_14654,N_13830);
and U19570 (N_19570,N_15011,N_14230);
nand U19571 (N_19571,N_14905,N_14694);
and U19572 (N_19572,N_13344,N_12551);
or U19573 (N_19573,N_15602,N_15376);
or U19574 (N_19574,N_14544,N_13268);
nand U19575 (N_19575,N_14199,N_15906);
xor U19576 (N_19576,N_13867,N_14124);
nand U19577 (N_19577,N_13800,N_14361);
nand U19578 (N_19578,N_15030,N_14230);
or U19579 (N_19579,N_12593,N_12601);
or U19580 (N_19580,N_12995,N_15792);
and U19581 (N_19581,N_12383,N_15848);
nor U19582 (N_19582,N_12946,N_13869);
nand U19583 (N_19583,N_14043,N_12117);
or U19584 (N_19584,N_14474,N_14043);
nor U19585 (N_19585,N_15775,N_14872);
and U19586 (N_19586,N_15186,N_14730);
and U19587 (N_19587,N_13466,N_13573);
and U19588 (N_19588,N_13491,N_12415);
nor U19589 (N_19589,N_15814,N_13330);
nand U19590 (N_19590,N_14613,N_13813);
and U19591 (N_19591,N_13727,N_13154);
nand U19592 (N_19592,N_15009,N_15248);
or U19593 (N_19593,N_14185,N_15737);
nor U19594 (N_19594,N_13263,N_15419);
and U19595 (N_19595,N_15755,N_14711);
nand U19596 (N_19596,N_14327,N_12017);
nand U19597 (N_19597,N_12313,N_15776);
or U19598 (N_19598,N_15272,N_15120);
and U19599 (N_19599,N_14921,N_15443);
nor U19600 (N_19600,N_13581,N_14901);
nand U19601 (N_19601,N_13007,N_13073);
or U19602 (N_19602,N_14865,N_13013);
or U19603 (N_19603,N_12487,N_12402);
or U19604 (N_19604,N_13515,N_13211);
xor U19605 (N_19605,N_13229,N_14467);
xnor U19606 (N_19606,N_15273,N_12701);
and U19607 (N_19607,N_13636,N_14261);
nor U19608 (N_19608,N_15917,N_15171);
and U19609 (N_19609,N_14125,N_13157);
nand U19610 (N_19610,N_15385,N_13851);
or U19611 (N_19611,N_12288,N_13936);
or U19612 (N_19612,N_12584,N_13771);
nand U19613 (N_19613,N_13099,N_14227);
nand U19614 (N_19614,N_15145,N_13920);
nand U19615 (N_19615,N_14390,N_12401);
or U19616 (N_19616,N_14716,N_13364);
and U19617 (N_19617,N_14382,N_13733);
and U19618 (N_19618,N_13332,N_14327);
nor U19619 (N_19619,N_13403,N_15429);
nor U19620 (N_19620,N_14404,N_15919);
nor U19621 (N_19621,N_13770,N_13900);
or U19622 (N_19622,N_13835,N_14946);
nor U19623 (N_19623,N_13105,N_12747);
or U19624 (N_19624,N_15987,N_12239);
nand U19625 (N_19625,N_14965,N_14093);
nand U19626 (N_19626,N_12628,N_13580);
and U19627 (N_19627,N_15118,N_12666);
or U19628 (N_19628,N_15002,N_13091);
nand U19629 (N_19629,N_14778,N_12587);
and U19630 (N_19630,N_14914,N_14511);
nand U19631 (N_19631,N_14139,N_15003);
and U19632 (N_19632,N_12655,N_14845);
nor U19633 (N_19633,N_13483,N_14243);
or U19634 (N_19634,N_15328,N_13349);
or U19635 (N_19635,N_12372,N_15202);
or U19636 (N_19636,N_14423,N_15355);
and U19637 (N_19637,N_15010,N_12032);
nand U19638 (N_19638,N_12135,N_15461);
nor U19639 (N_19639,N_12902,N_13892);
nand U19640 (N_19640,N_15820,N_14912);
and U19641 (N_19641,N_12605,N_13828);
and U19642 (N_19642,N_13543,N_14199);
nand U19643 (N_19643,N_13210,N_13686);
nor U19644 (N_19644,N_15131,N_15469);
or U19645 (N_19645,N_12715,N_15963);
or U19646 (N_19646,N_15523,N_15062);
nor U19647 (N_19647,N_15292,N_15392);
or U19648 (N_19648,N_15862,N_12979);
nand U19649 (N_19649,N_15616,N_13357);
nand U19650 (N_19650,N_15609,N_14620);
and U19651 (N_19651,N_14267,N_13017);
nor U19652 (N_19652,N_14242,N_13771);
and U19653 (N_19653,N_12115,N_14649);
nand U19654 (N_19654,N_13933,N_12497);
nand U19655 (N_19655,N_14860,N_15864);
nand U19656 (N_19656,N_14921,N_13715);
or U19657 (N_19657,N_13138,N_12712);
or U19658 (N_19658,N_12990,N_14254);
or U19659 (N_19659,N_12071,N_15083);
nand U19660 (N_19660,N_15490,N_14769);
and U19661 (N_19661,N_12141,N_15454);
nand U19662 (N_19662,N_14090,N_14860);
nand U19663 (N_19663,N_12771,N_12878);
or U19664 (N_19664,N_15100,N_14612);
nor U19665 (N_19665,N_12787,N_12249);
or U19666 (N_19666,N_13369,N_15784);
xnor U19667 (N_19667,N_12784,N_14874);
nand U19668 (N_19668,N_13825,N_15820);
and U19669 (N_19669,N_14730,N_13433);
nor U19670 (N_19670,N_15516,N_14271);
or U19671 (N_19671,N_14351,N_12953);
and U19672 (N_19672,N_15014,N_15348);
nor U19673 (N_19673,N_15217,N_12107);
nor U19674 (N_19674,N_14600,N_14810);
and U19675 (N_19675,N_13717,N_15600);
nand U19676 (N_19676,N_12911,N_12991);
and U19677 (N_19677,N_12687,N_12912);
nor U19678 (N_19678,N_13505,N_13977);
or U19679 (N_19679,N_15905,N_15378);
or U19680 (N_19680,N_12634,N_14194);
nor U19681 (N_19681,N_12218,N_13172);
and U19682 (N_19682,N_14584,N_15355);
nand U19683 (N_19683,N_12432,N_12994);
and U19684 (N_19684,N_12654,N_12598);
nor U19685 (N_19685,N_14214,N_13776);
or U19686 (N_19686,N_15196,N_14787);
nor U19687 (N_19687,N_15835,N_15213);
and U19688 (N_19688,N_13709,N_12145);
nand U19689 (N_19689,N_15962,N_12073);
or U19690 (N_19690,N_15528,N_15115);
and U19691 (N_19691,N_12049,N_12574);
and U19692 (N_19692,N_12933,N_14924);
nand U19693 (N_19693,N_15792,N_13844);
and U19694 (N_19694,N_12990,N_13955);
or U19695 (N_19695,N_14797,N_15431);
nand U19696 (N_19696,N_12674,N_15330);
or U19697 (N_19697,N_12807,N_15290);
and U19698 (N_19698,N_13509,N_14404);
or U19699 (N_19699,N_14197,N_13060);
nand U19700 (N_19700,N_13204,N_12081);
xor U19701 (N_19701,N_13296,N_12073);
nor U19702 (N_19702,N_15606,N_13376);
and U19703 (N_19703,N_14543,N_13626);
or U19704 (N_19704,N_15714,N_12306);
and U19705 (N_19705,N_14939,N_13452);
or U19706 (N_19706,N_12348,N_14637);
or U19707 (N_19707,N_14406,N_12030);
and U19708 (N_19708,N_14787,N_12075);
nand U19709 (N_19709,N_12756,N_12223);
nor U19710 (N_19710,N_13147,N_15963);
or U19711 (N_19711,N_13324,N_13402);
nor U19712 (N_19712,N_15721,N_12866);
nand U19713 (N_19713,N_14824,N_12020);
or U19714 (N_19714,N_15766,N_14469);
nand U19715 (N_19715,N_12545,N_13871);
nand U19716 (N_19716,N_13133,N_12489);
and U19717 (N_19717,N_13955,N_14277);
nor U19718 (N_19718,N_12623,N_12979);
nor U19719 (N_19719,N_14062,N_14714);
or U19720 (N_19720,N_13477,N_14426);
or U19721 (N_19721,N_14444,N_14445);
or U19722 (N_19722,N_15022,N_12511);
nor U19723 (N_19723,N_13163,N_15285);
and U19724 (N_19724,N_13073,N_15285);
nand U19725 (N_19725,N_15880,N_14084);
nand U19726 (N_19726,N_15970,N_12425);
or U19727 (N_19727,N_15432,N_14763);
nand U19728 (N_19728,N_15679,N_14439);
nand U19729 (N_19729,N_12947,N_14926);
and U19730 (N_19730,N_12296,N_14108);
xnor U19731 (N_19731,N_14162,N_13522);
or U19732 (N_19732,N_13424,N_15302);
and U19733 (N_19733,N_14711,N_15175);
nor U19734 (N_19734,N_15998,N_13591);
nand U19735 (N_19735,N_14421,N_15818);
and U19736 (N_19736,N_15537,N_12537);
nand U19737 (N_19737,N_15670,N_13235);
and U19738 (N_19738,N_12483,N_15168);
and U19739 (N_19739,N_12134,N_15422);
and U19740 (N_19740,N_14955,N_14061);
nor U19741 (N_19741,N_14908,N_15412);
nor U19742 (N_19742,N_13511,N_13845);
or U19743 (N_19743,N_12587,N_13782);
and U19744 (N_19744,N_15695,N_12390);
nand U19745 (N_19745,N_12672,N_15679);
nor U19746 (N_19746,N_13362,N_12064);
nand U19747 (N_19747,N_14048,N_14420);
or U19748 (N_19748,N_12015,N_12557);
nor U19749 (N_19749,N_13572,N_15961);
nand U19750 (N_19750,N_14459,N_13043);
or U19751 (N_19751,N_12962,N_12417);
nor U19752 (N_19752,N_12494,N_12803);
or U19753 (N_19753,N_15554,N_12714);
or U19754 (N_19754,N_15987,N_14129);
or U19755 (N_19755,N_14374,N_13508);
nor U19756 (N_19756,N_14778,N_15620);
nor U19757 (N_19757,N_15291,N_15461);
or U19758 (N_19758,N_12832,N_15161);
nand U19759 (N_19759,N_13734,N_13511);
or U19760 (N_19760,N_12527,N_13655);
or U19761 (N_19761,N_12459,N_15413);
or U19762 (N_19762,N_14552,N_14513);
and U19763 (N_19763,N_14401,N_15691);
nor U19764 (N_19764,N_15503,N_12678);
nand U19765 (N_19765,N_13255,N_15651);
and U19766 (N_19766,N_14737,N_12365);
nand U19767 (N_19767,N_15748,N_12331);
nand U19768 (N_19768,N_15032,N_12407);
nand U19769 (N_19769,N_15573,N_13045);
and U19770 (N_19770,N_12205,N_12096);
nand U19771 (N_19771,N_14714,N_15324);
nor U19772 (N_19772,N_12259,N_15228);
and U19773 (N_19773,N_12780,N_14586);
or U19774 (N_19774,N_15880,N_12090);
nand U19775 (N_19775,N_12783,N_12893);
xnor U19776 (N_19776,N_13921,N_14726);
and U19777 (N_19777,N_14503,N_13387);
or U19778 (N_19778,N_15184,N_14820);
and U19779 (N_19779,N_13188,N_13230);
nand U19780 (N_19780,N_14198,N_14753);
nand U19781 (N_19781,N_14383,N_15037);
or U19782 (N_19782,N_14143,N_14283);
nor U19783 (N_19783,N_13365,N_12938);
nand U19784 (N_19784,N_15155,N_14422);
or U19785 (N_19785,N_14098,N_12102);
and U19786 (N_19786,N_14349,N_15259);
and U19787 (N_19787,N_12282,N_15987);
nand U19788 (N_19788,N_13854,N_14509);
or U19789 (N_19789,N_12129,N_13753);
nor U19790 (N_19790,N_14066,N_12453);
or U19791 (N_19791,N_14521,N_14876);
nand U19792 (N_19792,N_13170,N_13829);
and U19793 (N_19793,N_12325,N_12664);
xor U19794 (N_19794,N_13936,N_13175);
nor U19795 (N_19795,N_12792,N_14822);
and U19796 (N_19796,N_15520,N_12022);
or U19797 (N_19797,N_15754,N_13845);
nor U19798 (N_19798,N_14567,N_14905);
nand U19799 (N_19799,N_14067,N_13019);
nor U19800 (N_19800,N_13906,N_13493);
nor U19801 (N_19801,N_13613,N_12137);
or U19802 (N_19802,N_13997,N_12121);
nor U19803 (N_19803,N_13295,N_15556);
nand U19804 (N_19804,N_13442,N_14791);
nor U19805 (N_19805,N_12196,N_12580);
nor U19806 (N_19806,N_14134,N_12416);
and U19807 (N_19807,N_12648,N_14421);
nand U19808 (N_19808,N_13789,N_15362);
nand U19809 (N_19809,N_12662,N_14012);
nor U19810 (N_19810,N_13354,N_12257);
nand U19811 (N_19811,N_14355,N_12584);
or U19812 (N_19812,N_14103,N_15370);
nor U19813 (N_19813,N_15389,N_13674);
nand U19814 (N_19814,N_15302,N_12220);
and U19815 (N_19815,N_13118,N_15517);
nor U19816 (N_19816,N_13844,N_15922);
xor U19817 (N_19817,N_13528,N_13422);
or U19818 (N_19818,N_12236,N_15609);
and U19819 (N_19819,N_15174,N_14494);
nor U19820 (N_19820,N_14400,N_13396);
or U19821 (N_19821,N_14120,N_12400);
nand U19822 (N_19822,N_15801,N_12423);
or U19823 (N_19823,N_12962,N_14866);
nand U19824 (N_19824,N_14150,N_15420);
or U19825 (N_19825,N_15345,N_12170);
and U19826 (N_19826,N_15824,N_12154);
nor U19827 (N_19827,N_12221,N_13894);
and U19828 (N_19828,N_14240,N_15845);
and U19829 (N_19829,N_13638,N_15849);
or U19830 (N_19830,N_13552,N_15773);
or U19831 (N_19831,N_13366,N_15058);
nor U19832 (N_19832,N_13574,N_12364);
nand U19833 (N_19833,N_13875,N_12120);
or U19834 (N_19834,N_13827,N_13483);
nor U19835 (N_19835,N_13364,N_15829);
nor U19836 (N_19836,N_15841,N_15967);
and U19837 (N_19837,N_14795,N_14867);
or U19838 (N_19838,N_13193,N_12517);
nand U19839 (N_19839,N_13970,N_14049);
nor U19840 (N_19840,N_12584,N_12628);
nor U19841 (N_19841,N_12628,N_13198);
and U19842 (N_19842,N_14002,N_12642);
nor U19843 (N_19843,N_12711,N_12677);
and U19844 (N_19844,N_12733,N_13717);
nor U19845 (N_19845,N_14907,N_15798);
nor U19846 (N_19846,N_13277,N_13307);
or U19847 (N_19847,N_12145,N_13880);
nor U19848 (N_19848,N_14417,N_15256);
nor U19849 (N_19849,N_13599,N_12440);
nor U19850 (N_19850,N_14347,N_13846);
and U19851 (N_19851,N_13605,N_15070);
and U19852 (N_19852,N_13900,N_15679);
and U19853 (N_19853,N_15913,N_15203);
nand U19854 (N_19854,N_13062,N_15870);
nor U19855 (N_19855,N_14858,N_15249);
nor U19856 (N_19856,N_15492,N_13870);
nand U19857 (N_19857,N_15973,N_15658);
and U19858 (N_19858,N_14174,N_14944);
and U19859 (N_19859,N_13252,N_12853);
nor U19860 (N_19860,N_12699,N_15972);
nor U19861 (N_19861,N_15977,N_13219);
nor U19862 (N_19862,N_14879,N_13979);
or U19863 (N_19863,N_14462,N_13930);
or U19864 (N_19864,N_12289,N_14786);
or U19865 (N_19865,N_14694,N_13002);
nor U19866 (N_19866,N_14225,N_14929);
nand U19867 (N_19867,N_15455,N_12061);
and U19868 (N_19868,N_15179,N_14813);
nor U19869 (N_19869,N_13937,N_15548);
and U19870 (N_19870,N_12266,N_12216);
nand U19871 (N_19871,N_12340,N_15231);
nand U19872 (N_19872,N_15274,N_12973);
nor U19873 (N_19873,N_15650,N_14080);
and U19874 (N_19874,N_14817,N_13236);
nand U19875 (N_19875,N_15674,N_13029);
or U19876 (N_19876,N_15670,N_14280);
and U19877 (N_19877,N_12386,N_14864);
and U19878 (N_19878,N_12721,N_14388);
and U19879 (N_19879,N_14325,N_12979);
and U19880 (N_19880,N_12462,N_15249);
nor U19881 (N_19881,N_14462,N_13798);
and U19882 (N_19882,N_14380,N_12662);
nor U19883 (N_19883,N_12606,N_15213);
nand U19884 (N_19884,N_12601,N_13858);
and U19885 (N_19885,N_13582,N_14254);
nand U19886 (N_19886,N_13833,N_12482);
and U19887 (N_19887,N_15327,N_12412);
and U19888 (N_19888,N_13460,N_12870);
nand U19889 (N_19889,N_14786,N_15584);
nor U19890 (N_19890,N_13037,N_14301);
nor U19891 (N_19891,N_15284,N_14537);
xnor U19892 (N_19892,N_15342,N_15507);
and U19893 (N_19893,N_13092,N_12010);
and U19894 (N_19894,N_14413,N_13241);
and U19895 (N_19895,N_13613,N_15119);
nor U19896 (N_19896,N_15659,N_15712);
nand U19897 (N_19897,N_15822,N_12573);
nor U19898 (N_19898,N_15146,N_12726);
or U19899 (N_19899,N_14835,N_15051);
or U19900 (N_19900,N_15491,N_12308);
and U19901 (N_19901,N_12854,N_15550);
or U19902 (N_19902,N_14694,N_12403);
or U19903 (N_19903,N_12511,N_14240);
and U19904 (N_19904,N_14655,N_12996);
nor U19905 (N_19905,N_15821,N_13646);
and U19906 (N_19906,N_15490,N_13805);
nand U19907 (N_19907,N_15578,N_15362);
nor U19908 (N_19908,N_14380,N_13952);
nor U19909 (N_19909,N_15707,N_12216);
nor U19910 (N_19910,N_12278,N_13489);
or U19911 (N_19911,N_12794,N_13985);
nand U19912 (N_19912,N_13366,N_14654);
nand U19913 (N_19913,N_12787,N_12354);
and U19914 (N_19914,N_12053,N_15317);
nor U19915 (N_19915,N_13800,N_14032);
nor U19916 (N_19916,N_14606,N_12236);
and U19917 (N_19917,N_15127,N_14872);
or U19918 (N_19918,N_13235,N_13616);
and U19919 (N_19919,N_14396,N_12240);
nand U19920 (N_19920,N_13827,N_14826);
or U19921 (N_19921,N_15052,N_12081);
nand U19922 (N_19922,N_12772,N_12922);
or U19923 (N_19923,N_15900,N_14305);
and U19924 (N_19924,N_14607,N_14756);
or U19925 (N_19925,N_12858,N_14765);
nand U19926 (N_19926,N_12134,N_12162);
and U19927 (N_19927,N_13317,N_15902);
nor U19928 (N_19928,N_14107,N_14393);
nor U19929 (N_19929,N_12476,N_13954);
nand U19930 (N_19930,N_14083,N_14691);
nand U19931 (N_19931,N_15848,N_14796);
nor U19932 (N_19932,N_13754,N_12735);
nor U19933 (N_19933,N_15757,N_14087);
nor U19934 (N_19934,N_13707,N_12947);
and U19935 (N_19935,N_13363,N_13031);
xor U19936 (N_19936,N_15015,N_15311);
and U19937 (N_19937,N_12080,N_15938);
or U19938 (N_19938,N_13121,N_15705);
nor U19939 (N_19939,N_15653,N_13293);
or U19940 (N_19940,N_14126,N_12441);
and U19941 (N_19941,N_12038,N_15218);
nand U19942 (N_19942,N_14986,N_15844);
or U19943 (N_19943,N_14734,N_13201);
or U19944 (N_19944,N_14612,N_13944);
or U19945 (N_19945,N_13211,N_12318);
nand U19946 (N_19946,N_12255,N_14116);
and U19947 (N_19947,N_15441,N_12631);
nand U19948 (N_19948,N_14583,N_15819);
or U19949 (N_19949,N_15856,N_15819);
nor U19950 (N_19950,N_13701,N_12741);
nand U19951 (N_19951,N_15366,N_14009);
and U19952 (N_19952,N_12600,N_13813);
xor U19953 (N_19953,N_15073,N_15194);
or U19954 (N_19954,N_14042,N_15824);
nand U19955 (N_19955,N_13356,N_12174);
nor U19956 (N_19956,N_12584,N_14876);
nand U19957 (N_19957,N_15890,N_15051);
or U19958 (N_19958,N_15881,N_15923);
or U19959 (N_19959,N_12150,N_14630);
and U19960 (N_19960,N_13209,N_15542);
and U19961 (N_19961,N_14935,N_14957);
or U19962 (N_19962,N_14114,N_12010);
or U19963 (N_19963,N_15513,N_13459);
and U19964 (N_19964,N_13887,N_14372);
nand U19965 (N_19965,N_12624,N_12058);
and U19966 (N_19966,N_13110,N_12639);
nor U19967 (N_19967,N_15821,N_15351);
nand U19968 (N_19968,N_15367,N_12541);
or U19969 (N_19969,N_12219,N_14217);
or U19970 (N_19970,N_15327,N_15008);
nor U19971 (N_19971,N_15817,N_13344);
and U19972 (N_19972,N_15265,N_14444);
and U19973 (N_19973,N_13489,N_12081);
nand U19974 (N_19974,N_15007,N_13519);
nor U19975 (N_19975,N_15560,N_14867);
and U19976 (N_19976,N_15605,N_12129);
nor U19977 (N_19977,N_13974,N_14342);
and U19978 (N_19978,N_15588,N_12193);
nand U19979 (N_19979,N_14120,N_15235);
nand U19980 (N_19980,N_12394,N_15427);
or U19981 (N_19981,N_14405,N_13403);
nor U19982 (N_19982,N_12800,N_14102);
xor U19983 (N_19983,N_12699,N_15573);
xor U19984 (N_19984,N_13675,N_13421);
nor U19985 (N_19985,N_12184,N_12253);
and U19986 (N_19986,N_13090,N_15817);
nand U19987 (N_19987,N_14365,N_15113);
nor U19988 (N_19988,N_13639,N_15854);
and U19989 (N_19989,N_13934,N_14692);
nor U19990 (N_19990,N_14053,N_12961);
xnor U19991 (N_19991,N_15863,N_13760);
and U19992 (N_19992,N_14358,N_15651);
and U19993 (N_19993,N_14212,N_15699);
nand U19994 (N_19994,N_14101,N_15698);
or U19995 (N_19995,N_12977,N_13192);
nor U19996 (N_19996,N_14572,N_15302);
nand U19997 (N_19997,N_15521,N_12403);
nor U19998 (N_19998,N_12585,N_14261);
or U19999 (N_19999,N_15388,N_14382);
nor UO_0 (O_0,N_18351,N_16366);
or UO_1 (O_1,N_19748,N_17224);
nand UO_2 (O_2,N_17944,N_16391);
nor UO_3 (O_3,N_18570,N_18717);
and UO_4 (O_4,N_17297,N_16078);
or UO_5 (O_5,N_16923,N_18090);
and UO_6 (O_6,N_16551,N_18167);
and UO_7 (O_7,N_19977,N_17119);
or UO_8 (O_8,N_17366,N_16243);
and UO_9 (O_9,N_17524,N_18461);
nand UO_10 (O_10,N_18964,N_16463);
and UO_11 (O_11,N_18679,N_17319);
nor UO_12 (O_12,N_16177,N_17339);
xor UO_13 (O_13,N_17635,N_18418);
or UO_14 (O_14,N_18478,N_16434);
or UO_15 (O_15,N_19223,N_19236);
nor UO_16 (O_16,N_17794,N_16088);
and UO_17 (O_17,N_16002,N_19176);
xnor UO_18 (O_18,N_18168,N_19194);
nor UO_19 (O_19,N_16454,N_18234);
nand UO_20 (O_20,N_18618,N_18640);
nor UO_21 (O_21,N_19419,N_17200);
and UO_22 (O_22,N_19926,N_16111);
or UO_23 (O_23,N_17981,N_19452);
and UO_24 (O_24,N_16521,N_16234);
nand UO_25 (O_25,N_19244,N_16746);
or UO_26 (O_26,N_16553,N_17164);
and UO_27 (O_27,N_17428,N_17463);
nand UO_28 (O_28,N_16493,N_16407);
nand UO_29 (O_29,N_17334,N_16261);
or UO_30 (O_30,N_19542,N_18265);
nor UO_31 (O_31,N_18658,N_19033);
or UO_32 (O_32,N_16264,N_16068);
or UO_33 (O_33,N_19700,N_18103);
nand UO_34 (O_34,N_17574,N_19118);
or UO_35 (O_35,N_19835,N_19648);
xnor UO_36 (O_36,N_19734,N_19512);
or UO_37 (O_37,N_18297,N_16736);
or UO_38 (O_38,N_16847,N_19480);
nor UO_39 (O_39,N_16653,N_19618);
nor UO_40 (O_40,N_19010,N_17446);
nor UO_41 (O_41,N_19921,N_19668);
nor UO_42 (O_42,N_19330,N_18380);
and UO_43 (O_43,N_18838,N_18486);
nand UO_44 (O_44,N_19467,N_16566);
or UO_45 (O_45,N_18357,N_16090);
nand UO_46 (O_46,N_19016,N_18249);
nor UO_47 (O_47,N_17513,N_16939);
or UO_48 (O_48,N_17064,N_16299);
nand UO_49 (O_49,N_19691,N_16851);
nor UO_50 (O_50,N_17525,N_17138);
and UO_51 (O_51,N_16091,N_17278);
xnor UO_52 (O_52,N_18866,N_19047);
nor UO_53 (O_53,N_19089,N_19388);
nor UO_54 (O_54,N_17501,N_19009);
nor UO_55 (O_55,N_17595,N_19358);
nor UO_56 (O_56,N_17491,N_17755);
nand UO_57 (O_57,N_17482,N_18197);
and UO_58 (O_58,N_18994,N_18169);
nor UO_59 (O_59,N_16937,N_18945);
nor UO_60 (O_60,N_19293,N_19157);
nor UO_61 (O_61,N_18962,N_17540);
and UO_62 (O_62,N_17627,N_16771);
or UO_63 (O_63,N_18671,N_17144);
and UO_64 (O_64,N_16561,N_16323);
nor UO_65 (O_65,N_18941,N_19201);
nor UO_66 (O_66,N_18963,N_16630);
nand UO_67 (O_67,N_16344,N_16306);
nand UO_68 (O_68,N_16385,N_16572);
and UO_69 (O_69,N_17195,N_18952);
nor UO_70 (O_70,N_18507,N_16855);
nor UO_71 (O_71,N_19642,N_16614);
nand UO_72 (O_72,N_16338,N_16025);
nand UO_73 (O_73,N_17072,N_18470);
or UO_74 (O_74,N_16357,N_18513);
and UO_75 (O_75,N_16818,N_16639);
or UO_76 (O_76,N_16618,N_16349);
and UO_77 (O_77,N_17506,N_17492);
or UO_78 (O_78,N_16980,N_16441);
nor UO_79 (O_79,N_16508,N_18378);
and UO_80 (O_80,N_16764,N_18222);
or UO_81 (O_81,N_17653,N_19923);
and UO_82 (O_82,N_17955,N_18091);
nor UO_83 (O_83,N_18703,N_19900);
or UO_84 (O_84,N_18899,N_19101);
or UO_85 (O_85,N_19600,N_19566);
nand UO_86 (O_86,N_16279,N_19973);
nor UO_87 (O_87,N_19332,N_17221);
nor UO_88 (O_88,N_16423,N_19998);
nand UO_89 (O_89,N_17038,N_17400);
nor UO_90 (O_90,N_18788,N_19262);
and UO_91 (O_91,N_16472,N_16223);
or UO_92 (O_92,N_19401,N_17959);
or UO_93 (O_93,N_17536,N_17637);
or UO_94 (O_94,N_17839,N_16749);
or UO_95 (O_95,N_19481,N_18338);
or UO_96 (O_96,N_16662,N_19905);
or UO_97 (O_97,N_19684,N_16389);
and UO_98 (O_98,N_16994,N_17399);
nand UO_99 (O_99,N_18660,N_18804);
nand UO_100 (O_100,N_19298,N_17208);
xor UO_101 (O_101,N_16012,N_18200);
and UO_102 (O_102,N_16467,N_19984);
and UO_103 (O_103,N_16158,N_16332);
or UO_104 (O_104,N_16367,N_19629);
nand UO_105 (O_105,N_19940,N_16095);
xnor UO_106 (O_106,N_19697,N_17859);
and UO_107 (O_107,N_17597,N_19614);
xor UO_108 (O_108,N_17923,N_16916);
and UO_109 (O_109,N_16358,N_17474);
or UO_110 (O_110,N_17893,N_18048);
or UO_111 (O_111,N_17042,N_16778);
nor UO_112 (O_112,N_17318,N_18092);
or UO_113 (O_113,N_18661,N_17109);
nand UO_114 (O_114,N_17805,N_17417);
nand UO_115 (O_115,N_18560,N_17914);
nor UO_116 (O_116,N_19536,N_17100);
or UO_117 (O_117,N_17850,N_16948);
and UO_118 (O_118,N_17188,N_19755);
and UO_119 (O_119,N_18377,N_17941);
and UO_120 (O_120,N_19902,N_16048);
nor UO_121 (O_121,N_19251,N_16194);
nor UO_122 (O_122,N_16514,N_18620);
nor UO_123 (O_123,N_16635,N_17889);
or UO_124 (O_124,N_19317,N_17977);
nor UO_125 (O_125,N_18014,N_18553);
or UO_126 (O_126,N_19666,N_17332);
nor UO_127 (O_127,N_18095,N_19119);
xnor UO_128 (O_128,N_17662,N_16696);
or UO_129 (O_129,N_18628,N_18245);
and UO_130 (O_130,N_19321,N_16210);
and UO_131 (O_131,N_17738,N_16897);
nand UO_132 (O_132,N_17105,N_17372);
nor UO_133 (O_133,N_17193,N_17680);
nand UO_134 (O_134,N_17659,N_19443);
or UO_135 (O_135,N_17457,N_19883);
or UO_136 (O_136,N_19007,N_19058);
nand UO_137 (O_137,N_19473,N_17369);
xnor UO_138 (O_138,N_18369,N_16978);
or UO_139 (O_139,N_17043,N_16118);
nor UO_140 (O_140,N_17337,N_18436);
or UO_141 (O_141,N_16651,N_18604);
nor UO_142 (O_142,N_19282,N_16935);
or UO_143 (O_143,N_19965,N_17612);
nand UO_144 (O_144,N_19580,N_17325);
nand UO_145 (O_145,N_19819,N_17930);
nand UO_146 (O_146,N_19798,N_19573);
nor UO_147 (O_147,N_17004,N_19264);
xor UO_148 (O_148,N_17182,N_18428);
nand UO_149 (O_149,N_16748,N_19844);
or UO_150 (O_150,N_18578,N_18756);
nand UO_151 (O_151,N_18746,N_16719);
nand UO_152 (O_152,N_17819,N_19652);
nor UO_153 (O_153,N_18586,N_16711);
nor UO_154 (O_154,N_18516,N_16519);
nand UO_155 (O_155,N_19767,N_17807);
or UO_156 (O_156,N_18525,N_16144);
nand UO_157 (O_157,N_17057,N_19785);
or UO_158 (O_158,N_17519,N_18031);
and UO_159 (O_159,N_19268,N_18087);
nor UO_160 (O_160,N_18081,N_17190);
and UO_161 (O_161,N_16756,N_16076);
nor UO_162 (O_162,N_18207,N_17473);
nand UO_163 (O_163,N_17026,N_18646);
and UO_164 (O_164,N_19535,N_17438);
nor UO_165 (O_165,N_18629,N_18910);
nand UO_166 (O_166,N_17565,N_18164);
nand UO_167 (O_167,N_17720,N_18074);
or UO_168 (O_168,N_17034,N_16416);
and UO_169 (O_169,N_17426,N_19671);
nand UO_170 (O_170,N_19060,N_18251);
nand UO_171 (O_171,N_16953,N_19751);
and UO_172 (O_172,N_19368,N_18337);
and UO_173 (O_173,N_19731,N_16135);
nand UO_174 (O_174,N_19820,N_19499);
nand UO_175 (O_175,N_16427,N_19729);
nand UO_176 (O_176,N_18934,N_17033);
or UO_177 (O_177,N_17736,N_19191);
or UO_178 (O_178,N_17013,N_16426);
and UO_179 (O_179,N_18198,N_16433);
nor UO_180 (O_180,N_18957,N_17449);
and UO_181 (O_181,N_19789,N_18669);
nand UO_182 (O_182,N_18153,N_19379);
and UO_183 (O_183,N_19543,N_19455);
nand UO_184 (O_184,N_18789,N_16658);
nor UO_185 (O_185,N_19838,N_18987);
and UO_186 (O_186,N_19722,N_18240);
or UO_187 (O_187,N_18481,N_16143);
or UO_188 (O_188,N_17782,N_19766);
xnor UO_189 (O_189,N_18284,N_19909);
and UO_190 (O_190,N_19479,N_17475);
or UO_191 (O_191,N_16995,N_19341);
and UO_192 (O_192,N_17296,N_17160);
and UO_193 (O_193,N_19065,N_19640);
nor UO_194 (O_194,N_19969,N_17329);
and UO_195 (O_195,N_17689,N_17960);
or UO_196 (O_196,N_17324,N_17471);
nor UO_197 (O_197,N_19267,N_17966);
and UO_198 (O_198,N_16914,N_18732);
nand UO_199 (O_199,N_16790,N_19702);
nand UO_200 (O_200,N_19803,N_16447);
or UO_201 (O_201,N_16965,N_17315);
nand UO_202 (O_202,N_16873,N_18902);
and UO_203 (O_203,N_18685,N_18216);
and UO_204 (O_204,N_17908,N_16986);
or UO_205 (O_205,N_17494,N_16750);
nor UO_206 (O_206,N_16465,N_18793);
nor UO_207 (O_207,N_19274,N_16398);
and UO_208 (O_208,N_17936,N_19444);
or UO_209 (O_209,N_16799,N_18325);
nand UO_210 (O_210,N_17732,N_17517);
nand UO_211 (O_211,N_18127,N_18411);
xnor UO_212 (O_212,N_17347,N_17476);
and UO_213 (O_213,N_16924,N_19689);
nor UO_214 (O_214,N_16274,N_19877);
or UO_215 (O_215,N_18736,N_19218);
and UO_216 (O_216,N_18044,N_17785);
and UO_217 (O_217,N_16402,N_19351);
nand UO_218 (O_218,N_17813,N_19276);
and UO_219 (O_219,N_18473,N_16710);
or UO_220 (O_220,N_18312,N_17872);
nor UO_221 (O_221,N_19799,N_19163);
and UO_222 (O_222,N_16854,N_19156);
or UO_223 (O_223,N_18121,N_19565);
nand UO_224 (O_224,N_17017,N_19990);
or UO_225 (O_225,N_18540,N_16380);
nand UO_226 (O_226,N_19544,N_16451);
nor UO_227 (O_227,N_16580,N_18258);
or UO_228 (O_228,N_17697,N_16959);
xor UO_229 (O_229,N_16930,N_18896);
nand UO_230 (O_230,N_16738,N_16782);
nand UO_231 (O_231,N_17310,N_19403);
or UO_232 (O_232,N_17974,N_17156);
or UO_233 (O_233,N_17511,N_17177);
xnor UO_234 (O_234,N_18806,N_19879);
or UO_235 (O_235,N_18829,N_19328);
or UO_236 (O_236,N_17410,N_19911);
or UO_237 (O_237,N_16517,N_19849);
and UO_238 (O_238,N_16522,N_19486);
or UO_239 (O_239,N_19518,N_17521);
nor UO_240 (O_240,N_17729,N_18900);
or UO_241 (O_241,N_18315,N_16126);
and UO_242 (O_242,N_17066,N_18721);
nand UO_243 (O_243,N_18040,N_18862);
xor UO_244 (O_244,N_16151,N_17032);
or UO_245 (O_245,N_18006,N_17508);
or UO_246 (O_246,N_19741,N_16288);
xor UO_247 (O_247,N_17701,N_16865);
nor UO_248 (O_248,N_19399,N_18291);
nor UO_249 (O_249,N_17847,N_16724);
nor UO_250 (O_250,N_19081,N_18751);
nand UO_251 (O_251,N_19246,N_17700);
xnor UO_252 (O_252,N_16648,N_18727);
and UO_253 (O_253,N_16975,N_17500);
nand UO_254 (O_254,N_19088,N_16425);
or UO_255 (O_255,N_19064,N_17461);
or UO_256 (O_256,N_16200,N_18193);
or UO_257 (O_257,N_18484,N_18172);
or UO_258 (O_258,N_19000,N_19829);
and UO_259 (O_259,N_16491,N_16690);
nor UO_260 (O_260,N_17881,N_16583);
and UO_261 (O_261,N_19533,N_19370);
nor UO_262 (O_262,N_18442,N_19606);
nand UO_263 (O_263,N_19611,N_18270);
and UO_264 (O_264,N_16721,N_18539);
nand UO_265 (O_265,N_19409,N_17467);
and UO_266 (O_266,N_18616,N_19206);
xnor UO_267 (O_267,N_16046,N_16940);
nand UO_268 (O_268,N_17037,N_17758);
or UO_269 (O_269,N_19270,N_16424);
nand UO_270 (O_270,N_16259,N_17722);
nand UO_271 (O_271,N_18650,N_17523);
and UO_272 (O_272,N_17104,N_17486);
nor UO_273 (O_273,N_17980,N_16540);
or UO_274 (O_274,N_17730,N_19318);
and UO_275 (O_275,N_19617,N_18991);
or UO_276 (O_276,N_18644,N_16008);
nand UO_277 (O_277,N_18977,N_18298);
xor UO_278 (O_278,N_17673,N_19485);
or UO_279 (O_279,N_16689,N_18253);
nand UO_280 (O_280,N_16826,N_16237);
nor UO_281 (O_281,N_16103,N_16999);
and UO_282 (O_282,N_17687,N_19256);
or UO_283 (O_283,N_17810,N_18422);
or UO_284 (O_284,N_19778,N_16686);
and UO_285 (O_285,N_18626,N_16247);
nand UO_286 (O_286,N_18821,N_16283);
nor UO_287 (O_287,N_18026,N_16763);
nor UO_288 (O_288,N_19797,N_18859);
and UO_289 (O_289,N_16775,N_16998);
and UO_290 (O_290,N_19663,N_18059);
or UO_291 (O_291,N_19625,N_16715);
nor UO_292 (O_292,N_18792,N_19355);
nor UO_293 (O_293,N_19728,N_18875);
nor UO_294 (O_294,N_17108,N_18906);
nor UO_295 (O_295,N_16270,N_16659);
or UO_296 (O_296,N_19448,N_16643);
and UO_297 (O_297,N_16182,N_17365);
nand UO_298 (O_298,N_16399,N_19724);
nor UO_299 (O_299,N_18592,N_17529);
or UO_300 (O_300,N_18515,N_17143);
nand UO_301 (O_301,N_16355,N_17258);
or UO_302 (O_302,N_17846,N_19359);
nor UO_303 (O_303,N_17978,N_19224);
nor UO_304 (O_304,N_16541,N_16856);
nor UO_305 (O_305,N_18733,N_16406);
and UO_306 (O_306,N_17290,N_19269);
and UO_307 (O_307,N_19210,N_18262);
xnor UO_308 (O_308,N_17898,N_16501);
xor UO_309 (O_309,N_18052,N_18735);
nor UO_310 (O_310,N_16803,N_17423);
and UO_311 (O_311,N_18815,N_19784);
nor UO_312 (O_312,N_18203,N_19241);
nand UO_313 (O_313,N_16954,N_18491);
nand UO_314 (O_314,N_16557,N_16867);
or UO_315 (O_315,N_18981,N_18009);
nand UO_316 (O_316,N_17769,N_17279);
nor UO_317 (O_317,N_16345,N_18675);
nor UO_318 (O_318,N_18272,N_19791);
nand UO_319 (O_319,N_16334,N_16221);
nand UO_320 (O_320,N_16966,N_18365);
and UO_321 (O_321,N_19086,N_16976);
or UO_322 (O_322,N_16035,N_18755);
or UO_323 (O_323,N_18567,N_19914);
nor UO_324 (O_324,N_19238,N_19787);
and UO_325 (O_325,N_19828,N_19777);
or UO_326 (O_326,N_19209,N_18210);
and UO_327 (O_327,N_18185,N_19343);
or UO_328 (O_328,N_19308,N_17096);
or UO_329 (O_329,N_17518,N_19773);
nand UO_330 (O_330,N_17079,N_16430);
and UO_331 (O_331,N_18082,N_17052);
nor UO_332 (O_332,N_19521,N_16071);
xor UO_333 (O_333,N_18928,N_18358);
and UO_334 (O_334,N_19759,N_17274);
nor UO_335 (O_335,N_18841,N_17071);
nor UO_336 (O_336,N_18122,N_19402);
and UO_337 (O_337,N_17228,N_18762);
nor UO_338 (O_338,N_16797,N_19584);
and UO_339 (O_339,N_16005,N_18083);
nand UO_340 (O_340,N_16660,N_16375);
and UO_341 (O_341,N_19472,N_19460);
nor UO_342 (O_342,N_19747,N_16110);
and UO_343 (O_343,N_16510,N_17041);
or UO_344 (O_344,N_18316,N_19336);
and UO_345 (O_345,N_16861,N_16988);
and UO_346 (O_346,N_16699,N_17538);
and UO_347 (O_347,N_17213,N_16529);
nand UO_348 (O_348,N_19096,N_16951);
nand UO_349 (O_349,N_16615,N_17531);
and UO_350 (O_350,N_17382,N_17621);
nor UO_351 (O_351,N_16436,N_16169);
and UO_352 (O_352,N_19159,N_16958);
nand UO_353 (O_353,N_18690,N_16537);
and UO_354 (O_354,N_19216,N_16781);
nand UO_355 (O_355,N_17910,N_19108);
and UO_356 (O_356,N_19655,N_18088);
nor UO_357 (O_357,N_18205,N_16442);
nor UO_358 (O_358,N_16011,N_17281);
nor UO_359 (O_359,N_17825,N_16712);
xnor UO_360 (O_360,N_16809,N_19757);
nand UO_361 (O_361,N_19720,N_19901);
or UO_362 (O_362,N_17841,N_19885);
or UO_363 (O_363,N_17654,N_19525);
and UO_364 (O_364,N_18763,N_16142);
or UO_365 (O_365,N_19674,N_18818);
nand UO_366 (O_366,N_18062,N_18719);
or UO_367 (O_367,N_17711,N_19669);
nand UO_368 (O_368,N_16617,N_19248);
or UO_369 (O_369,N_17192,N_19063);
and UO_370 (O_370,N_17497,N_18740);
nor UO_371 (O_371,N_16415,N_16178);
and UO_372 (O_372,N_17823,N_19044);
nor UO_373 (O_373,N_16382,N_16007);
and UO_374 (O_374,N_18734,N_18431);
nor UO_375 (O_375,N_19847,N_16578);
nor UO_376 (O_376,N_17938,N_16667);
or UO_377 (O_377,N_19884,N_17262);
or UO_378 (O_378,N_17110,N_16250);
or UO_379 (O_379,N_17263,N_17185);
nor UO_380 (O_380,N_17316,N_16734);
and UO_381 (O_381,N_18030,N_19864);
nor UO_382 (O_382,N_17089,N_16827);
and UO_383 (O_383,N_19927,N_16587);
and UO_384 (O_384,N_19181,N_19908);
nor UO_385 (O_385,N_19474,N_18348);
and UO_386 (O_386,N_17196,N_17202);
and UO_387 (O_387,N_17095,N_18229);
xor UO_388 (O_388,N_18129,N_16400);
nand UO_389 (O_389,N_18113,N_19185);
and UO_390 (O_390,N_18580,N_16934);
or UO_391 (O_391,N_18217,N_17747);
nor UO_392 (O_392,N_19109,N_17764);
or UO_393 (O_393,N_19762,N_16860);
or UO_394 (O_394,N_17174,N_19556);
nor UO_395 (O_395,N_17772,N_19805);
nor UO_396 (O_396,N_19934,N_16910);
or UO_397 (O_397,N_16882,N_19295);
nand UO_398 (O_398,N_19307,N_19898);
nor UO_399 (O_399,N_18552,N_19137);
nand UO_400 (O_400,N_19788,N_17996);
nor UO_401 (O_401,N_16636,N_16171);
nor UO_402 (O_402,N_17705,N_19391);
and UO_403 (O_403,N_17367,N_18046);
and UO_404 (O_404,N_19003,N_16258);
or UO_405 (O_405,N_16547,N_16823);
nor UO_406 (O_406,N_19017,N_16100);
or UO_407 (O_407,N_18189,N_18830);
and UO_408 (O_408,N_16530,N_16575);
or UO_409 (O_409,N_18559,N_17373);
and UO_410 (O_410,N_16877,N_16337);
or UO_411 (O_411,N_17078,N_16645);
nand UO_412 (O_412,N_19349,N_16628);
nand UO_413 (O_413,N_17514,N_19792);
or UO_414 (O_414,N_16215,N_16038);
nor UO_415 (O_415,N_16228,N_16569);
and UO_416 (O_416,N_16486,N_16211);
and UO_417 (O_417,N_19041,N_18467);
or UO_418 (O_418,N_19812,N_16497);
nor UO_419 (O_419,N_18182,N_18905);
nor UO_420 (O_420,N_17879,N_19171);
or UO_421 (O_421,N_18015,N_17254);
nand UO_422 (O_422,N_17998,N_16067);
nor UO_423 (O_423,N_17776,N_18366);
or UO_424 (O_424,N_17210,N_16312);
and UO_425 (O_425,N_16758,N_17888);
or UO_426 (O_426,N_17897,N_18022);
nor UO_427 (O_427,N_16805,N_17246);
nor UO_428 (O_428,N_16240,N_18108);
and UO_429 (O_429,N_19422,N_19627);
nand UO_430 (O_430,N_19146,N_17987);
and UO_431 (O_431,N_16147,N_17757);
nor UO_432 (O_432,N_16968,N_18939);
and UO_433 (O_433,N_16160,N_19302);
and UO_434 (O_434,N_16460,N_19333);
and UO_435 (O_435,N_18713,N_17289);
and UO_436 (O_436,N_19366,N_19598);
nand UO_437 (O_437,N_17949,N_17920);
nor UO_438 (O_438,N_18742,N_19528);
xor UO_439 (O_439,N_19384,N_17752);
or UO_440 (O_440,N_18870,N_19483);
or UO_441 (O_441,N_17826,N_18271);
nand UO_442 (O_442,N_16664,N_16864);
and UO_443 (O_443,N_16316,N_19854);
nand UO_444 (O_444,N_17237,N_18093);
or UO_445 (O_445,N_19897,N_18754);
or UO_446 (O_446,N_19501,N_16800);
or UO_447 (O_447,N_17077,N_16278);
nand UO_448 (O_448,N_18967,N_18757);
nand UO_449 (O_449,N_18564,N_17504);
nand UO_450 (O_450,N_18141,N_17112);
nor UO_451 (O_451,N_16204,N_16668);
and UO_452 (O_452,N_17883,N_18446);
or UO_453 (O_453,N_19892,N_19868);
or UO_454 (O_454,N_16303,N_18143);
nand UO_455 (O_455,N_17868,N_17081);
and UO_456 (O_456,N_17056,N_18498);
nand UO_457 (O_457,N_16343,N_18075);
nor UO_458 (O_458,N_19682,N_18427);
or UO_459 (O_459,N_19804,N_16439);
and UO_460 (O_460,N_19174,N_16677);
or UO_461 (O_461,N_17699,N_18853);
nor UO_462 (O_462,N_16395,N_16863);
or UO_463 (O_463,N_18523,N_18016);
or UO_464 (O_464,N_17681,N_18299);
or UO_465 (O_465,N_16116,N_17670);
or UO_466 (O_466,N_16092,N_16161);
xnor UO_467 (O_467,N_19559,N_17594);
and UO_468 (O_468,N_18653,N_19922);
and UO_469 (O_469,N_18948,N_16810);
and UO_470 (O_470,N_19414,N_17241);
and UO_471 (O_471,N_19744,N_18033);
or UO_472 (O_472,N_19097,N_19597);
or UO_473 (O_473,N_16084,N_18638);
nor UO_474 (O_474,N_19951,N_18394);
nand UO_475 (O_475,N_19721,N_18494);
or UO_476 (O_476,N_18748,N_19389);
or UO_477 (O_477,N_19100,N_16661);
nor UO_478 (O_478,N_16167,N_18566);
nand UO_479 (O_479,N_16363,N_17750);
nand UO_480 (O_480,N_16242,N_19507);
and UO_481 (O_481,N_17330,N_19588);
and UO_482 (O_482,N_19488,N_19323);
nand UO_483 (O_483,N_18633,N_17273);
nand UO_484 (O_484,N_18233,N_19350);
and UO_485 (O_485,N_19180,N_19381);
and UO_486 (O_486,N_19205,N_16086);
or UO_487 (O_487,N_19719,N_17116);
and UO_488 (O_488,N_19439,N_18927);
nor UO_489 (O_489,N_17198,N_18842);
nor UO_490 (O_490,N_18575,N_19756);
nor UO_491 (O_491,N_18213,N_19842);
nand UO_492 (O_492,N_19975,N_16473);
or UO_493 (O_493,N_18360,N_19468);
and UO_494 (O_494,N_17549,N_18079);
and UO_495 (O_495,N_19353,N_19602);
and UO_496 (O_496,N_17266,N_16592);
and UO_497 (O_497,N_16073,N_19252);
or UO_498 (O_498,N_19140,N_16788);
nand UO_499 (O_499,N_17167,N_19040);
or UO_500 (O_500,N_18388,N_18163);
or UO_501 (O_501,N_17616,N_19092);
or UO_502 (O_502,N_18652,N_17580);
nand UO_503 (O_503,N_17059,N_16052);
xor UO_504 (O_504,N_19069,N_16487);
and UO_505 (O_505,N_16990,N_17717);
xnor UO_506 (O_506,N_19628,N_17706);
and UO_507 (O_507,N_17061,N_18280);
xor UO_508 (O_508,N_19635,N_19235);
or UO_509 (O_509,N_19475,N_16356);
nor UO_510 (O_510,N_17590,N_17596);
or UO_511 (O_511,N_17300,N_18408);
or UO_512 (O_512,N_19075,N_16915);
or UO_513 (O_513,N_17140,N_16889);
and UO_514 (O_514,N_17447,N_19245);
nand UO_515 (O_515,N_16155,N_16656);
and UO_516 (O_516,N_19169,N_19084);
or UO_517 (O_517,N_19726,N_18135);
nand UO_518 (O_518,N_16921,N_18529);
or UO_519 (O_519,N_18654,N_16074);
nor UO_520 (O_520,N_17614,N_16443);
or UO_521 (O_521,N_18250,N_17082);
nand UO_522 (O_522,N_16795,N_16806);
nand UO_523 (O_523,N_16884,N_16479);
xor UO_524 (O_524,N_16313,N_17284);
nand UO_525 (O_525,N_19579,N_16720);
or UO_526 (O_526,N_18404,N_16461);
or UO_527 (O_527,N_16817,N_17636);
nor UO_528 (O_528,N_16346,N_18102);
nand UO_529 (O_529,N_18808,N_17314);
or UO_530 (O_530,N_18777,N_16887);
nand UO_531 (O_531,N_18120,N_19098);
or UO_532 (O_532,N_16191,N_17951);
and UO_533 (O_533,N_17801,N_18908);
nand UO_534 (O_534,N_16180,N_16043);
nand UO_535 (O_535,N_17276,N_18105);
and UO_536 (O_536,N_18725,N_18851);
and UO_537 (O_537,N_19874,N_19018);
nand UO_538 (O_538,N_18903,N_19790);
or UO_539 (O_539,N_19919,N_18997);
nand UO_540 (O_540,N_18277,N_19509);
nor UO_541 (O_541,N_18538,N_17087);
nor UO_542 (O_542,N_16122,N_18533);
xor UO_543 (O_543,N_19265,N_17003);
or UO_544 (O_544,N_16744,N_18814);
and UO_545 (O_545,N_17451,N_17067);
nor UO_546 (O_546,N_19768,N_19932);
nor UO_547 (O_547,N_17796,N_17617);
or UO_548 (O_548,N_17424,N_16535);
nand UO_549 (O_549,N_18413,N_18744);
xor UO_550 (O_550,N_16904,N_18268);
nor UO_551 (O_551,N_18805,N_16985);
nand UO_552 (O_552,N_17668,N_17734);
and UO_553 (O_553,N_17047,N_17777);
and UO_554 (O_554,N_16918,N_17570);
and UO_555 (O_555,N_18731,N_16798);
nand UO_556 (O_556,N_17895,N_19229);
or UO_557 (O_557,N_17420,N_18243);
nor UO_558 (O_558,N_18179,N_17799);
and UO_559 (O_559,N_18330,N_18627);
xor UO_560 (O_560,N_17844,N_18285);
and UO_561 (O_561,N_17968,N_19484);
and UO_562 (O_562,N_19631,N_16671);
or UO_563 (O_563,N_16811,N_16214);
and UO_564 (O_564,N_19801,N_18911);
and UO_565 (O_565,N_19032,N_16128);
nand UO_566 (O_566,N_18849,N_16755);
or UO_567 (O_567,N_19860,N_16179);
nor UO_568 (O_568,N_18607,N_19586);
nor UO_569 (O_569,N_16102,N_16523);
or UO_570 (O_570,N_19863,N_17137);
nand UO_571 (O_571,N_16219,N_16016);
and UO_572 (O_572,N_17587,N_18988);
nor UO_573 (O_573,N_19303,N_18053);
nand UO_574 (O_574,N_16933,N_18557);
nand UO_575 (O_575,N_17135,N_17927);
or UO_576 (O_576,N_18542,N_17348);
and UO_577 (O_577,N_18474,N_19664);
and UO_578 (O_578,N_19811,N_18175);
nor UO_579 (O_579,N_17341,N_18047);
nor UO_580 (O_580,N_18327,N_17303);
nand UO_581 (O_581,N_16971,N_18591);
nor UO_582 (O_582,N_19534,N_19042);
nand UO_583 (O_583,N_17035,N_17688);
or UO_584 (O_584,N_17827,N_17972);
and UO_585 (O_585,N_17338,N_17028);
nand UO_586 (O_586,N_19020,N_18398);
nor UO_587 (O_587,N_16206,N_19810);
nor UO_588 (O_588,N_18895,N_17721);
or UO_589 (O_589,N_16675,N_17142);
or UO_590 (O_590,N_18873,N_17389);
nand UO_591 (O_591,N_16017,N_18802);
or UO_592 (O_592,N_17197,N_16927);
or UO_593 (O_593,N_16351,N_18813);
or UO_594 (O_594,N_17354,N_17359);
nand UO_595 (O_595,N_16422,N_17656);
nor UO_596 (O_596,N_17610,N_18278);
nor UO_597 (O_597,N_19487,N_16629);
or UO_598 (O_598,N_19002,N_17255);
or UO_599 (O_599,N_19215,N_18549);
nand UO_600 (O_600,N_17435,N_16115);
nand UO_601 (O_601,N_17465,N_17380);
and UO_602 (O_602,N_18683,N_17954);
nand UO_603 (O_603,N_17145,N_18913);
nor UO_604 (O_604,N_18176,N_19587);
and UO_605 (O_605,N_19647,N_16396);
or UO_606 (O_606,N_19367,N_17657);
or UO_607 (O_607,N_17298,N_19253);
and UO_608 (O_608,N_16513,N_18354);
and UO_609 (O_609,N_18868,N_19142);
nor UO_610 (O_610,N_18772,N_17952);
nor UO_611 (O_611,N_17638,N_19106);
or UO_612 (O_612,N_19859,N_17068);
nor UO_613 (O_613,N_16546,N_18926);
or UO_614 (O_614,N_18438,N_18929);
and UO_615 (O_615,N_18130,N_16532);
nor UO_616 (O_616,N_17490,N_18605);
nand UO_617 (O_617,N_16637,N_18673);
and UO_618 (O_618,N_18410,N_19558);
and UO_619 (O_619,N_17187,N_16291);
nand UO_620 (O_620,N_17378,N_18011);
nand UO_621 (O_621,N_18479,N_19936);
and UO_622 (O_622,N_19337,N_19243);
or UO_623 (O_623,N_17544,N_17270);
xnor UO_624 (O_624,N_17176,N_16544);
or UO_625 (O_625,N_16825,N_18293);
or UO_626 (O_626,N_16022,N_17216);
or UO_627 (O_627,N_17459,N_18459);
and UO_628 (O_628,N_16796,N_18615);
nand UO_629 (O_629,N_19956,N_18959);
or UO_630 (O_630,N_16456,N_16531);
or UO_631 (O_631,N_19261,N_19771);
and UO_632 (O_632,N_19683,N_18659);
or UO_633 (O_633,N_17103,N_18889);
or UO_634 (O_634,N_16157,N_18000);
nand UO_635 (O_635,N_17444,N_18308);
nand UO_636 (O_636,N_18065,N_18623);
and UO_637 (O_637,N_19029,N_19641);
and UO_638 (O_638,N_18576,N_19613);
nor UO_639 (O_639,N_16836,N_19147);
nand UO_640 (O_640,N_17117,N_16121);
and UO_641 (O_641,N_19745,N_16902);
and UO_642 (O_642,N_16520,N_19021);
nor UO_643 (O_643,N_18209,N_18407);
nand UO_644 (O_644,N_16911,N_16901);
and UO_645 (O_645,N_16133,N_17948);
and UO_646 (O_646,N_18577,N_19769);
or UO_647 (O_647,N_19090,N_19872);
nand UO_648 (O_648,N_16362,N_17011);
nand UO_649 (O_649,N_19324,N_19172);
xor UO_650 (O_650,N_16987,N_16952);
nand UO_651 (O_651,N_17808,N_16753);
nor UO_652 (O_652,N_19782,N_19530);
nand UO_653 (O_653,N_18028,N_16075);
and UO_654 (O_654,N_16808,N_16213);
nand UO_655 (O_655,N_17710,N_16606);
nand UO_656 (O_656,N_17007,N_18329);
nor UO_657 (O_657,N_17751,N_19571);
and UO_658 (O_658,N_16080,N_19993);
or UO_659 (O_659,N_18666,N_19195);
nor UO_660 (O_660,N_18361,N_17969);
or UO_661 (O_661,N_18223,N_18791);
or UO_662 (O_662,N_16949,N_18328);
and UO_663 (O_663,N_18084,N_17118);
and UO_664 (O_664,N_16845,N_17708);
nor UO_665 (O_665,N_19589,N_17151);
nand UO_666 (O_666,N_16480,N_19971);
or UO_667 (O_667,N_16853,N_17631);
xor UO_668 (O_668,N_16612,N_16292);
nor UO_669 (O_669,N_16663,N_18383);
nand UO_670 (O_670,N_17312,N_17684);
nand UO_671 (O_671,N_17557,N_19322);
nand UO_672 (O_672,N_16621,N_17956);
nand UO_673 (O_673,N_18252,N_18097);
nor UO_674 (O_674,N_17015,N_18547);
nor UO_675 (O_675,N_19843,N_19061);
nor UO_676 (O_676,N_18710,N_17742);
nor UO_677 (O_677,N_19746,N_18917);
nand UO_678 (O_678,N_17390,N_18331);
nor UO_679 (O_679,N_17526,N_18869);
nor UO_680 (O_680,N_18025,N_16922);
nor UO_681 (O_681,N_18582,N_16722);
or UO_682 (O_682,N_17598,N_19019);
or UO_683 (O_683,N_17806,N_18089);
and UO_684 (O_684,N_16762,N_16209);
and UO_685 (O_685,N_17027,N_18840);
and UO_686 (O_686,N_16153,N_16014);
and UO_687 (O_687,N_18978,N_17264);
nor UO_688 (O_688,N_16478,N_16411);
xor UO_689 (O_689,N_17640,N_17592);
nor UO_690 (O_690,N_19430,N_16850);
and UO_691 (O_691,N_18946,N_17634);
nand UO_692 (O_692,N_19931,N_18585);
or UO_693 (O_693,N_19083,N_16218);
or UO_694 (O_694,N_17434,N_19495);
or UO_695 (O_695,N_16300,N_17440);
and UO_696 (O_696,N_18322,N_18211);
and UO_697 (O_697,N_18466,N_17124);
or UO_698 (O_698,N_17904,N_17018);
or UO_699 (O_699,N_17589,N_18288);
or UO_700 (O_700,N_17652,N_17884);
nand UO_701 (O_701,N_18376,N_17835);
or UO_702 (O_702,N_16619,N_16776);
or UO_703 (O_703,N_17783,N_17633);
or UO_704 (O_704,N_16929,N_19510);
and UO_705 (O_705,N_17915,N_18593);
nor UO_706 (O_706,N_16083,N_19563);
nand UO_707 (O_707,N_17005,N_17682);
and UO_708 (O_708,N_16372,N_16725);
or UO_709 (O_709,N_16342,N_19699);
nand UO_710 (O_710,N_19834,N_18528);
nand UO_711 (O_711,N_18573,N_17905);
or UO_712 (O_712,N_19976,N_19632);
nor UO_713 (O_713,N_17686,N_19074);
nor UO_714 (O_714,N_16352,N_17600);
nand UO_715 (O_715,N_16813,N_16186);
and UO_716 (O_716,N_16829,N_16101);
nor UO_717 (O_717,N_17302,N_18647);
nor UO_718 (O_718,N_19421,N_17848);
or UO_719 (O_719,N_19005,N_18400);
nand UO_720 (O_720,N_16562,N_19187);
nand UO_721 (O_721,N_18579,N_19152);
nor UO_722 (O_722,N_19636,N_19750);
nor UO_723 (O_723,N_19794,N_19417);
nand UO_724 (O_724,N_16376,N_18657);
and UO_725 (O_725,N_17550,N_16783);
or UO_726 (O_726,N_16023,N_19907);
nor UO_727 (O_727,N_18156,N_17683);
nand UO_728 (O_728,N_18147,N_18393);
or UO_729 (O_729,N_19024,N_17405);
nor UO_730 (O_730,N_18397,N_17256);
nor UO_731 (O_731,N_18021,N_17040);
nand UO_732 (O_732,N_16528,N_16252);
and UO_733 (O_733,N_18942,N_18184);
or UO_734 (O_734,N_18662,N_17409);
nor UO_735 (O_735,N_16304,N_16793);
or UO_736 (O_736,N_18823,N_19027);
nand UO_737 (O_737,N_16477,N_19680);
nor UO_738 (O_738,N_17760,N_16842);
nand UO_739 (O_739,N_17733,N_16010);
nand UO_740 (O_740,N_16626,N_16878);
or UO_741 (O_741,N_19870,N_18096);
nor UO_742 (O_742,N_18503,N_18302);
nand UO_743 (O_743,N_18146,N_18420);
nor UO_744 (O_744,N_17560,N_18460);
and UO_745 (O_745,N_17713,N_19562);
nor UO_746 (O_746,N_16883,N_17818);
nor UO_747 (O_747,N_19329,N_19173);
xnor UO_748 (O_748,N_18995,N_17211);
or UO_749 (O_749,N_16324,N_17532);
nand UO_750 (O_750,N_19432,N_16114);
nand UO_751 (O_751,N_18199,N_17362);
or UO_752 (O_752,N_19615,N_17586);
nand UO_753 (O_753,N_17374,N_18314);
nand UO_754 (O_754,N_19670,N_18519);
nand UO_755 (O_755,N_19345,N_16284);
nand UO_756 (O_756,N_19999,N_18319);
nor UO_757 (O_757,N_16203,N_17495);
or UO_758 (O_758,N_16627,N_18359);
and UO_759 (O_759,N_17556,N_18955);
or UO_760 (O_760,N_18872,N_19420);
nor UO_761 (O_761,N_16202,N_19703);
or UO_762 (O_762,N_16683,N_17269);
xnor UO_763 (O_763,N_18231,N_16296);
and UO_764 (O_764,N_19831,N_18370);
nor UO_765 (O_765,N_19286,N_18810);
nand UO_766 (O_766,N_16563,N_16354);
and UO_767 (O_767,N_17935,N_19437);
or UO_768 (O_768,N_16096,N_16991);
nand UO_769 (O_769,N_17466,N_18405);
or UO_770 (O_770,N_18947,N_17070);
and UO_771 (O_771,N_16693,N_18739);
or UO_772 (O_772,N_16709,N_19449);
nor UO_773 (O_773,N_19813,N_18396);
nor UO_774 (O_774,N_19808,N_17731);
or UO_775 (O_775,N_19456,N_17995);
nor UO_776 (O_776,N_19713,N_18944);
nor UO_777 (O_777,N_18070,N_17931);
nand UO_778 (O_778,N_17243,N_19660);
and UO_779 (O_779,N_18350,N_19709);
nand UO_780 (O_780,N_19162,N_19374);
nor UO_781 (O_781,N_17218,N_17349);
nand UO_782 (O_782,N_19263,N_18888);
or UO_783 (O_783,N_18069,N_18781);
or UO_784 (O_784,N_17655,N_19497);
nand UO_785 (O_785,N_16388,N_19127);
or UO_786 (O_786,N_18563,N_18861);
or UO_787 (O_787,N_17822,N_16205);
nand UO_788 (O_788,N_16928,N_19824);
and UO_789 (O_789,N_18343,N_16302);
or UO_790 (O_790,N_16679,N_17737);
nor UO_791 (O_791,N_17485,N_16512);
and UO_792 (O_792,N_16941,N_17075);
xor UO_793 (O_793,N_18705,N_19301);
and UO_794 (O_794,N_19408,N_17433);
nor UO_795 (O_795,N_19661,N_18972);
nor UO_796 (O_796,N_17178,N_19749);
nand UO_797 (O_797,N_17060,N_17132);
or UO_798 (O_798,N_18664,N_17419);
nand UO_799 (O_799,N_17726,N_17690);
and UO_800 (O_800,N_16241,N_18248);
nor UO_801 (O_801,N_16170,N_19240);
or UO_802 (O_802,N_19143,N_18003);
and UO_803 (O_803,N_18416,N_17441);
nand UO_804 (O_804,N_17280,N_16267);
and UO_805 (O_805,N_16970,N_17527);
nor UO_806 (O_806,N_17546,N_19227);
and UO_807 (O_807,N_16733,N_18989);
and UO_808 (O_808,N_18392,N_18174);
nand UO_809 (O_809,N_17707,N_18027);
nor UO_810 (O_810,N_17843,N_19280);
or UO_811 (O_811,N_16320,N_18512);
nand UO_812 (O_812,N_16140,N_16041);
nor UO_813 (O_813,N_17126,N_17890);
nand UO_814 (O_814,N_17173,N_18749);
nand UO_815 (O_815,N_19234,N_17111);
and UO_816 (O_816,N_16483,N_17464);
nand UO_817 (O_817,N_19306,N_19963);
nor UO_818 (O_818,N_18856,N_19772);
or UO_819 (O_819,N_16207,N_17054);
nor UO_820 (O_820,N_18041,N_16701);
nor UO_821 (O_821,N_19079,N_16159);
nor UO_822 (O_822,N_18257,N_18677);
or UO_823 (O_823,N_16117,N_16408);
and UO_824 (O_824,N_18678,N_17812);
and UO_825 (O_825,N_17854,N_19575);
or UO_826 (O_826,N_16047,N_19630);
nor UO_827 (O_827,N_19508,N_17973);
nand UO_828 (O_828,N_17191,N_18950);
nor UO_829 (O_829,N_18208,N_19113);
nand UO_830 (O_830,N_16979,N_17902);
or UO_831 (O_831,N_17024,N_16129);
nor UO_832 (O_832,N_17223,N_19672);
or UO_833 (O_833,N_18078,N_18969);
and UO_834 (O_834,N_17746,N_16872);
nand UO_835 (O_835,N_16432,N_19873);
or UO_836 (O_836,N_16058,N_17815);
nand UO_837 (O_837,N_18342,N_19237);
nand UO_838 (O_838,N_19441,N_17141);
nor UO_839 (O_839,N_17069,N_18998);
nor UO_840 (O_840,N_17129,N_18776);
nor UO_841 (O_841,N_17114,N_16666);
or UO_842 (O_842,N_18326,N_16435);
and UO_843 (O_843,N_18526,N_16641);
nor UO_844 (O_844,N_16602,N_18782);
nor UO_845 (O_845,N_17674,N_17204);
nor UO_846 (O_846,N_19561,N_19861);
and UO_847 (O_847,N_18774,N_16488);
nor UO_848 (O_848,N_19915,N_16906);
nor UO_849 (O_849,N_19653,N_18702);
and UO_850 (O_850,N_16069,N_17860);
nor UO_851 (O_851,N_18960,N_16181);
or UO_852 (O_852,N_19616,N_19554);
or UO_853 (O_853,N_16649,N_16294);
and UO_854 (O_854,N_18107,N_18971);
nand UO_855 (O_855,N_16977,N_17605);
nand UO_856 (O_856,N_19182,N_19736);
nand UO_857 (O_857,N_16319,N_18892);
or UO_858 (O_858,N_16350,N_18520);
nor UO_859 (O_859,N_16591,N_18583);
and UO_860 (O_860,N_16249,N_18613);
nor UO_861 (O_861,N_17539,N_16193);
or UO_862 (O_862,N_17899,N_17453);
and UO_863 (O_863,N_19889,N_19623);
nor UO_864 (O_864,N_17886,N_16828);
or UO_865 (O_865,N_17157,N_16694);
or UO_866 (O_866,N_18569,N_16238);
nand UO_867 (O_867,N_18468,N_16932);
or UO_868 (O_868,N_17404,N_17239);
nor UO_869 (O_869,N_19299,N_19519);
or UO_870 (O_870,N_17925,N_18345);
or UO_871 (O_871,N_19698,N_17021);
xor UO_872 (O_872,N_18601,N_16527);
nand UO_873 (O_873,N_17448,N_19135);
nor UO_874 (O_874,N_17125,N_19114);
or UO_875 (O_875,N_17327,N_19054);
and UO_876 (O_876,N_17564,N_17934);
nand UO_877 (O_877,N_19459,N_18305);
and UO_878 (O_878,N_17331,N_19154);
or UO_879 (O_879,N_16149,N_17669);
or UO_880 (O_880,N_16560,N_19503);
or UO_881 (O_881,N_19817,N_19896);
nand UO_882 (O_882,N_19582,N_18536);
nand UO_883 (O_883,N_17493,N_19121);
and UO_884 (O_884,N_18711,N_16094);
and UO_885 (O_885,N_19192,N_19822);
nand UO_886 (O_886,N_17107,N_16550);
or UO_887 (O_887,N_17512,N_17876);
or UO_888 (O_888,N_16944,N_18919);
nand UO_889 (O_889,N_19132,N_19718);
nor UO_890 (O_890,N_17849,N_17646);
or UO_891 (O_891,N_17383,N_18931);
and UO_892 (O_892,N_18753,N_16862);
or UO_893 (O_893,N_19891,N_18767);
or UO_894 (O_894,N_18005,N_19502);
nor UO_895 (O_895,N_18649,N_18119);
nor UO_896 (O_896,N_17870,N_17880);
or UO_897 (O_897,N_16136,N_18493);
and UO_898 (O_898,N_16166,N_16004);
nand UO_899 (O_899,N_18722,N_18382);
nand UO_900 (O_900,N_18833,N_18500);
nand UO_901 (O_901,N_17778,N_16290);
and UO_902 (O_902,N_16964,N_16981);
nor UO_903 (O_903,N_16938,N_16624);
or UO_904 (O_904,N_18775,N_18790);
and UO_905 (O_905,N_18877,N_18336);
or UO_906 (O_906,N_17179,N_17798);
or UO_907 (O_907,N_18076,N_18961);
nand UO_908 (O_908,N_16015,N_16457);
nand UO_909 (O_909,N_16688,N_16898);
nor UO_910 (O_910,N_18600,N_18864);
nor UO_911 (O_911,N_19814,N_19404);
nor UO_912 (O_912,N_16481,N_19289);
and UO_913 (O_913,N_16106,N_17231);
nand UO_914 (O_914,N_16429,N_17740);
and UO_915 (O_915,N_16554,N_18296);
nor UO_916 (O_916,N_17430,N_19862);
nand UO_917 (O_917,N_16285,N_16188);
or UO_918 (O_918,N_17505,N_18018);
nor UO_919 (O_919,N_17695,N_19657);
and UO_920 (O_920,N_19392,N_18956);
or UO_921 (O_921,N_17712,N_19292);
or UO_922 (O_922,N_16462,N_19390);
or UO_923 (O_923,N_18476,N_18532);
xnor UO_924 (O_924,N_16974,N_18384);
nand UO_925 (O_925,N_18237,N_18881);
or UO_926 (O_926,N_19964,N_16697);
and UO_927 (O_927,N_19447,N_19470);
or UO_928 (O_928,N_18937,N_19325);
nor UO_929 (O_929,N_19170,N_19644);
and UO_930 (O_930,N_19175,N_16740);
or UO_931 (O_931,N_16360,N_17784);
nand UO_932 (O_932,N_18511,N_16773);
nor UO_933 (O_933,N_18847,N_17547);
and UO_934 (O_934,N_17840,N_17678);
or UO_935 (O_935,N_17852,N_17821);
nand UO_936 (O_936,N_19226,N_18696);
or UO_937 (O_937,N_17335,N_17360);
or UO_938 (O_938,N_17800,N_18907);
nor UO_939 (O_939,N_16676,N_19284);
nor UO_940 (O_940,N_16120,N_18488);
and UO_941 (O_941,N_19857,N_19972);
or UO_942 (O_942,N_18154,N_17293);
and UO_943 (O_943,N_17418,N_18115);
and UO_944 (O_944,N_16132,N_18363);
and UO_945 (O_945,N_18155,N_18042);
or UO_946 (O_946,N_16431,N_19220);
nand UO_947 (O_947,N_16308,N_17857);
and UO_948 (O_948,N_17377,N_18890);
or UO_949 (O_949,N_16741,N_19429);
nand UO_950 (O_950,N_16586,N_16502);
and UO_951 (O_951,N_17744,N_19685);
nor UO_952 (O_952,N_16919,N_17545);
or UO_953 (O_953,N_16893,N_17833);
nor UO_954 (O_954,N_18165,N_19730);
nor UO_955 (O_955,N_19376,N_18820);
nor UO_956 (O_956,N_17248,N_17381);
nand UO_957 (O_957,N_17355,N_17620);
nand UO_958 (O_958,N_18414,N_16874);
nor UO_959 (O_959,N_19871,N_19442);
or UO_960 (O_960,N_19569,N_16729);
nand UO_961 (O_961,N_18568,N_17022);
nand UO_962 (O_962,N_19585,N_16770);
nor UO_963 (O_963,N_19290,N_16500);
and UO_964 (O_964,N_16548,N_17836);
or UO_965 (O_965,N_18244,N_18812);
nor UO_966 (O_966,N_19775,N_19271);
and UO_967 (O_967,N_16494,N_16731);
or UO_968 (O_968,N_18943,N_19153);
and UO_969 (O_969,N_18935,N_19545);
nor UO_970 (O_970,N_18930,N_19202);
and UO_971 (O_971,N_18819,N_18822);
or UO_972 (O_972,N_17181,N_16761);
or UO_973 (O_973,N_17442,N_16246);
or UO_974 (O_974,N_16792,N_17666);
and UO_975 (O_975,N_17541,N_17470);
or UO_976 (O_976,N_19426,N_16437);
nor UO_977 (O_977,N_16515,N_19574);
xor UO_978 (O_978,N_18504,N_18706);
and UO_979 (O_979,N_17694,N_18180);
nor UO_980 (O_980,N_17127,N_18858);
or UO_981 (O_981,N_19591,N_17454);
nor UO_982 (O_982,N_18544,N_18634);
nor UO_983 (O_983,N_17979,N_17450);
xnor UO_984 (O_984,N_17641,N_18178);
and UO_985 (O_985,N_17180,N_18136);
and UO_986 (O_986,N_18306,N_16538);
or UO_987 (O_987,N_16113,N_16072);
nand UO_988 (O_988,N_16920,N_17855);
or UO_989 (O_989,N_19687,N_16633);
nand UO_990 (O_990,N_17651,N_17170);
nand UO_991 (O_991,N_17016,N_16759);
nand UO_992 (O_992,N_18572,N_18063);
or UO_993 (O_993,N_18225,N_17715);
nor UO_994 (O_994,N_19012,N_19638);
nand UO_995 (O_995,N_17148,N_18144);
or UO_996 (O_996,N_18391,N_19880);
nand UO_997 (O_997,N_17472,N_17939);
or UO_998 (O_998,N_18876,N_17458);
nor UO_999 (O_999,N_19840,N_16281);
or UO_1000 (O_1000,N_19549,N_18020);
or UO_1001 (O_1001,N_18770,N_16187);
and UO_1002 (O_1002,N_17756,N_17639);
or UO_1003 (O_1003,N_19633,N_16199);
nand UO_1004 (O_1004,N_16608,N_19435);
nor UO_1005 (O_1005,N_16870,N_19761);
and UO_1006 (O_1006,N_18854,N_17907);
and UO_1007 (O_1007,N_16652,N_16045);
nand UO_1008 (O_1008,N_17824,N_16896);
nand UO_1009 (O_1009,N_18954,N_18936);
and UO_1010 (O_1010,N_18551,N_19428);
or UO_1011 (O_1011,N_18415,N_16837);
nor UO_1012 (O_1012,N_16482,N_17943);
xnor UO_1013 (O_1013,N_19851,N_19903);
or UO_1014 (O_1014,N_17749,N_16000);
nor UO_1015 (O_1015,N_19738,N_18457);
nand UO_1016 (O_1016,N_18324,N_16506);
nand UO_1017 (O_1017,N_18111,N_17489);
and UO_1018 (O_1018,N_19076,N_19034);
and UO_1019 (O_1019,N_18480,N_17063);
nand UO_1020 (O_1020,N_17106,N_19500);
and UO_1021 (O_1021,N_18160,N_19688);
and UO_1022 (O_1022,N_17567,N_19541);
or UO_1023 (O_1023,N_16604,N_19886);
and UO_1024 (O_1024,N_17183,N_18317);
or UO_1025 (O_1025,N_17561,N_17460);
nand UO_1026 (O_1026,N_16251,N_19275);
or UO_1027 (O_1027,N_19678,N_18728);
and UO_1028 (O_1028,N_16079,N_17240);
and UO_1029 (O_1029,N_16779,N_19982);
and UO_1030 (O_1030,N_17599,N_18012);
nand UO_1031 (O_1031,N_17613,N_16226);
nand UO_1032 (O_1032,N_19094,N_17092);
or UO_1033 (O_1033,N_19476,N_19568);
or UO_1034 (O_1034,N_18435,N_16674);
nor UO_1035 (O_1035,N_19057,N_17074);
or UO_1036 (O_1036,N_19514,N_17918);
and UO_1037 (O_1037,N_18453,N_19676);
nor UO_1038 (O_1038,N_19131,N_16365);
nor UO_1039 (O_1039,N_17873,N_19622);
and UO_1040 (O_1040,N_16165,N_16333);
and UO_1041 (O_1041,N_19453,N_16534);
or UO_1042 (O_1042,N_16053,N_18390);
and UO_1043 (O_1043,N_19992,N_17537);
and UO_1044 (O_1044,N_16490,N_18992);
and UO_1045 (O_1045,N_17102,N_19715);
and UO_1046 (O_1046,N_17411,N_16233);
and UO_1047 (O_1047,N_16098,N_16852);
and UO_1048 (O_1048,N_18531,N_16885);
or UO_1049 (O_1049,N_16282,N_19555);
nand UO_1050 (O_1050,N_18651,N_19316);
and UO_1051 (O_1051,N_16588,N_16185);
and UO_1052 (O_1052,N_16866,N_17236);
xnor UO_1053 (O_1053,N_18166,N_19213);
or UO_1054 (O_1054,N_18430,N_19760);
or UO_1055 (O_1055,N_18104,N_19407);
and UO_1056 (O_1056,N_17275,N_17479);
or UO_1057 (O_1057,N_16459,N_16453);
or UO_1058 (O_1058,N_18828,N_18712);
nor UO_1059 (O_1059,N_19725,N_16705);
nand UO_1060 (O_1060,N_16832,N_19385);
or UO_1061 (O_1061,N_16066,N_19523);
and UO_1062 (O_1062,N_17856,N_19168);
nand UO_1063 (O_1063,N_16881,N_18367);
and UO_1064 (O_1064,N_19929,N_17774);
nor UO_1065 (O_1065,N_16248,N_18401);
nor UO_1066 (O_1066,N_18741,N_16687);
nor UO_1067 (O_1067,N_19115,N_16341);
or UO_1068 (O_1068,N_18612,N_18715);
nor UO_1069 (O_1069,N_18595,N_19001);
nand UO_1070 (O_1070,N_17227,N_18672);
nor UO_1071 (O_1071,N_18132,N_19890);
nor UO_1072 (O_1072,N_19277,N_16556);
and UO_1073 (O_1073,N_17803,N_18555);
nand UO_1074 (O_1074,N_17395,N_19961);
or UO_1075 (O_1075,N_16287,N_19008);
nor UO_1076 (O_1076,N_19211,N_19723);
and UO_1077 (O_1077,N_19855,N_18764);
nand UO_1078 (O_1078,N_19727,N_16590);
nand UO_1079 (O_1079,N_16913,N_17830);
or UO_1080 (O_1080,N_18294,N_16130);
nor UO_1081 (O_1081,N_17483,N_18289);
and UO_1082 (O_1082,N_17650,N_17853);
or UO_1083 (O_1083,N_19763,N_17252);
or UO_1084 (O_1084,N_19796,N_19596);
nand UO_1085 (O_1085,N_18058,N_18162);
nor UO_1086 (O_1086,N_19866,N_17245);
and UO_1087 (O_1087,N_16732,N_19906);
nor UO_1088 (O_1088,N_16982,N_18224);
nand UO_1089 (O_1089,N_17025,N_16331);
nor UO_1090 (O_1090,N_18034,N_18036);
nor UO_1091 (O_1091,N_16684,N_18597);
and UO_1092 (O_1092,N_19117,N_18794);
or UO_1093 (O_1093,N_18809,N_16876);
nor UO_1094 (O_1094,N_18304,N_19546);
or UO_1095 (O_1095,N_17933,N_18975);
nor UO_1096 (O_1096,N_19360,N_19022);
nand UO_1097 (O_1097,N_16277,N_17507);
and UO_1098 (O_1098,N_16807,N_17097);
or UO_1099 (O_1099,N_18445,N_17554);
nand UO_1100 (O_1100,N_16198,N_16271);
nand UO_1101 (O_1101,N_19815,N_16839);
and UO_1102 (O_1102,N_16905,N_18064);
or UO_1103 (O_1103,N_19371,N_17123);
and UO_1104 (O_1104,N_17765,N_18695);
nor UO_1105 (O_1105,N_18080,N_16525);
or UO_1106 (O_1106,N_18611,N_16609);
or UO_1107 (O_1107,N_16616,N_17320);
nand UO_1108 (O_1108,N_19347,N_19138);
or UO_1109 (O_1109,N_19690,N_18068);
nor UO_1110 (O_1110,N_19506,N_19348);
nor UO_1111 (O_1111,N_16706,N_19331);
and UO_1112 (O_1112,N_17261,N_19564);
nand UO_1113 (O_1113,N_19059,N_18152);
nor UO_1114 (O_1114,N_16695,N_19538);
and UO_1115 (O_1115,N_16769,N_18440);
nand UO_1116 (O_1116,N_18619,N_16438);
or UO_1117 (O_1117,N_17579,N_18614);
and UO_1118 (O_1118,N_17344,N_19272);
nand UO_1119 (O_1119,N_19327,N_16507);
nor UO_1120 (O_1120,N_17413,N_17388);
nand UO_1121 (O_1121,N_17660,N_17522);
or UO_1122 (O_1122,N_17988,N_16963);
nor UO_1123 (O_1123,N_18610,N_16054);
nor UO_1124 (O_1124,N_16236,N_16428);
or UO_1125 (O_1125,N_18897,N_16742);
nand UO_1126 (O_1126,N_19887,N_19423);
nor UO_1127 (O_1127,N_18925,N_19943);
and UO_1128 (O_1128,N_19424,N_16201);
or UO_1129 (O_1129,N_19673,N_17403);
or UO_1130 (O_1130,N_16340,N_16943);
nand UO_1131 (O_1131,N_18730,N_17260);
nor UO_1132 (O_1132,N_16962,N_19651);
and UO_1133 (O_1133,N_19904,N_19619);
nor UO_1134 (O_1134,N_19204,N_17120);
nand UO_1135 (O_1135,N_16021,N_18737);
or UO_1136 (O_1136,N_18495,N_16032);
nand UO_1137 (O_1137,N_19659,N_19917);
nor UO_1138 (O_1138,N_17045,N_17719);
and UO_1139 (O_1139,N_18007,N_17385);
nand UO_1140 (O_1140,N_16172,N_16229);
nor UO_1141 (O_1141,N_18855,N_16831);
or UO_1142 (O_1142,N_17779,N_17607);
and UO_1143 (O_1143,N_19658,N_17305);
and UO_1144 (O_1144,N_18196,N_17878);
and UO_1145 (O_1145,N_17294,N_19740);
nand UO_1146 (O_1146,N_18817,N_16195);
or UO_1147 (O_1147,N_18188,N_17146);
nand UO_1148 (O_1148,N_16997,N_19987);
nor UO_1149 (O_1149,N_19196,N_17937);
and UO_1150 (O_1150,N_16168,N_19696);
and UO_1151 (O_1151,N_18990,N_18218);
or UO_1152 (O_1152,N_18880,N_16458);
and UO_1153 (O_1153,N_17947,N_18517);
or UO_1154 (O_1154,N_18332,N_16001);
and UO_1155 (O_1155,N_19395,N_17575);
and UO_1156 (O_1156,N_17672,N_19551);
nor UO_1157 (O_1157,N_19111,N_18455);
xor UO_1158 (O_1158,N_18347,N_18700);
nor UO_1159 (O_1159,N_17249,N_19129);
or UO_1160 (O_1160,N_16257,N_19431);
and UO_1161 (O_1161,N_17009,N_19300);
and UO_1162 (O_1162,N_17101,N_18275);
and UO_1163 (O_1163,N_16766,N_17287);
nor UO_1164 (O_1164,N_19477,N_16723);
or UO_1165 (O_1165,N_18537,N_16105);
nor UO_1166 (O_1166,N_16469,N_16670);
and UO_1167 (O_1167,N_17577,N_19966);
nor UO_1168 (O_1168,N_16581,N_19601);
or UO_1169 (O_1169,N_16217,N_17804);
and UO_1170 (O_1170,N_18970,N_18707);
nor UO_1171 (O_1171,N_18726,N_17496);
nand UO_1172 (O_1172,N_18395,N_18126);
nor UO_1173 (O_1173,N_18241,N_17698);
nor UO_1174 (O_1174,N_16605,N_17773);
nand UO_1175 (O_1175,N_18098,N_17502);
nor UO_1176 (O_1176,N_18642,N_19779);
and UO_1177 (O_1177,N_19764,N_19717);
and UO_1178 (O_1178,N_17456,N_18912);
or UO_1179 (O_1179,N_19567,N_19739);
and UO_1180 (O_1180,N_16956,N_17414);
nand UO_1181 (O_1181,N_18691,N_19795);
nand UO_1182 (O_1182,N_16378,N_16127);
nor UO_1183 (O_1183,N_17645,N_17436);
nor UO_1184 (O_1184,N_18594,N_18548);
and UO_1185 (O_1185,N_17268,N_17350);
nand UO_1186 (O_1186,N_18799,N_16393);
or UO_1187 (O_1187,N_16265,N_18112);
nor UO_1188 (O_1188,N_16470,N_18886);
and UO_1189 (O_1189,N_19496,N_18419);
and UO_1190 (O_1190,N_19038,N_18501);
or UO_1191 (O_1191,N_18676,N_17113);
nand UO_1192 (O_1192,N_19557,N_19548);
or UO_1193 (O_1193,N_18254,N_17166);
nor UO_1194 (O_1194,N_19639,N_18452);
nand UO_1195 (O_1195,N_19707,N_16222);
nand UO_1196 (O_1196,N_16162,N_17791);
or UO_1197 (O_1197,N_16703,N_19494);
nand UO_1198 (O_1198,N_17603,N_19466);
nand UO_1199 (O_1199,N_19189,N_16085);
or UO_1200 (O_1200,N_19126,N_17763);
nor UO_1201 (O_1201,N_19203,N_19948);
nand UO_1202 (O_1202,N_16368,N_17088);
nor UO_1203 (O_1203,N_19974,N_18032);
nor UO_1204 (O_1204,N_19164,N_18785);
or UO_1205 (O_1205,N_16912,N_17498);
or UO_1206 (O_1206,N_19800,N_18465);
or UO_1207 (O_1207,N_16571,N_18117);
and UO_1208 (O_1208,N_17986,N_19446);
and UO_1209 (O_1209,N_19517,N_18287);
and UO_1210 (O_1210,N_19177,N_16150);
and UO_1211 (O_1211,N_19043,N_18051);
or UO_1212 (O_1212,N_19463,N_19550);
or UO_1213 (O_1213,N_18920,N_16307);
nor UO_1214 (O_1214,N_17984,N_18958);
nand UO_1215 (O_1215,N_19513,N_19068);
nand UO_1216 (O_1216,N_16466,N_16640);
nor UO_1217 (O_1217,N_19400,N_16601);
and UO_1218 (O_1218,N_16392,N_18589);
nor UO_1219 (O_1219,N_18745,N_19941);
nand UO_1220 (O_1220,N_18622,N_16597);
and UO_1221 (O_1221,N_19406,N_18421);
or UO_1222 (O_1222,N_18846,N_19491);
nor UO_1223 (O_1223,N_19199,N_17172);
nand UO_1224 (O_1224,N_19547,N_16413);
or UO_1225 (O_1225,N_16452,N_16768);
nor UO_1226 (O_1226,N_16595,N_17623);
nor UO_1227 (O_1227,N_18364,N_17429);
and UO_1228 (O_1228,N_19190,N_19516);
and UO_1229 (O_1229,N_17222,N_18066);
nor UO_1230 (O_1230,N_18588,N_17006);
or UO_1231 (O_1231,N_18779,N_18918);
nor UO_1232 (O_1232,N_18556,N_18674);
or UO_1233 (O_1233,N_18800,N_17084);
or UO_1234 (O_1234,N_19626,N_18281);
and UO_1235 (O_1235,N_17379,N_16474);
or UO_1236 (O_1236,N_19123,N_19335);
nand UO_1237 (O_1237,N_19708,N_19288);
or UO_1238 (O_1238,N_17437,N_19369);
nor UO_1239 (O_1239,N_18759,N_19867);
and UO_1240 (O_1240,N_19304,N_19028);
nand UO_1241 (O_1241,N_16268,N_16967);
or UO_1242 (O_1242,N_16329,N_16840);
nand UO_1243 (O_1243,N_18983,N_16061);
or UO_1244 (O_1244,N_16373,N_19599);
or UO_1245 (O_1245,N_16890,N_16669);
or UO_1246 (O_1246,N_18836,N_19254);
and UO_1247 (O_1247,N_17696,N_16024);
or UO_1248 (O_1248,N_18801,N_17917);
or UO_1249 (O_1249,N_16405,N_19141);
nor UO_1250 (O_1250,N_18798,N_16255);
and UO_1251 (O_1251,N_18980,N_16984);
nor UO_1252 (O_1252,N_16708,N_17828);
nand UO_1253 (O_1253,N_17357,N_17387);
or UO_1254 (O_1254,N_17677,N_17967);
or UO_1255 (O_1255,N_17225,N_19451);
nor UO_1256 (O_1256,N_16511,N_17789);
or UO_1257 (O_1257,N_16293,N_19242);
and UO_1258 (O_1258,N_18371,N_16082);
or UO_1259 (O_1259,N_19878,N_16154);
nand UO_1260 (O_1260,N_19116,N_16752);
or UO_1261 (O_1261,N_19139,N_18344);
or UO_1262 (O_1262,N_17480,N_17593);
nor UO_1263 (O_1263,N_16044,N_18017);
nor UO_1264 (O_1264,N_18565,N_16263);
nor UO_1265 (O_1265,N_17963,N_17265);
and UO_1266 (O_1266,N_17871,N_17421);
and UO_1267 (O_1267,N_18045,N_18190);
and UO_1268 (O_1268,N_18019,N_19309);
nor UO_1269 (O_1269,N_16821,N_18631);
or UO_1270 (O_1270,N_16969,N_18985);
nor UO_1271 (O_1271,N_18346,N_19716);
or UO_1272 (O_1272,N_18901,N_19978);
nor UO_1273 (O_1273,N_16336,N_17133);
and UO_1274 (O_1274,N_16317,N_19925);
and UO_1275 (O_1275,N_18624,N_19372);
xor UO_1276 (O_1276,N_18283,N_16955);
nor UO_1277 (O_1277,N_19959,N_18173);
nand UO_1278 (O_1278,N_19537,N_16055);
nand UO_1279 (O_1279,N_16596,N_17304);
nand UO_1280 (O_1280,N_16533,N_16295);
nand UO_1281 (O_1281,N_16545,N_17510);
nor UO_1282 (O_1282,N_16370,N_17542);
and UO_1283 (O_1283,N_18024,N_17375);
nor UO_1284 (O_1284,N_16377,N_16505);
nand UO_1285 (O_1285,N_17989,N_19694);
and UO_1286 (O_1286,N_19996,N_17566);
nor UO_1287 (O_1287,N_17267,N_18826);
or UO_1288 (O_1288,N_18598,N_16942);
or UO_1289 (O_1289,N_17926,N_19200);
or UO_1290 (O_1290,N_19112,N_16576);
nor UO_1291 (O_1291,N_19679,N_16892);
or UO_1292 (O_1292,N_19179,N_18321);
nand UO_1293 (O_1293,N_19464,N_17648);
nor UO_1294 (O_1294,N_18863,N_16707);
or UO_1295 (O_1295,N_17606,N_19039);
nor UO_1296 (O_1296,N_17155,N_18372);
nand UO_1297 (O_1297,N_16401,N_19539);
nor UO_1298 (O_1298,N_18232,N_16326);
and UO_1299 (O_1299,N_18835,N_17412);
nand UO_1300 (O_1300,N_19560,N_19875);
xnor UO_1301 (O_1301,N_18850,N_17716);
nor UO_1302 (O_1302,N_18874,N_18496);
or UO_1303 (O_1303,N_19377,N_16266);
and UO_1304 (O_1304,N_18621,N_16936);
nor UO_1305 (O_1305,N_17364,N_16397);
or UO_1306 (O_1306,N_18522,N_18680);
nor UO_1307 (O_1307,N_17401,N_19609);
or UO_1308 (O_1308,N_17576,N_16131);
nand UO_1309 (O_1309,N_18403,N_19882);
and UO_1310 (O_1310,N_19531,N_17356);
or UO_1311 (O_1311,N_18202,N_18590);
nor UO_1312 (O_1312,N_19968,N_19572);
or UO_1313 (O_1313,N_17971,N_18356);
or UO_1314 (O_1314,N_16886,N_16822);
and UO_1315 (O_1315,N_18857,N_17408);
nand UO_1316 (O_1316,N_19865,N_16455);
nand UO_1317 (O_1317,N_17230,N_17520);
nand UO_1318 (O_1318,N_16036,N_17548);
nor UO_1319 (O_1319,N_16450,N_19910);
nor UO_1320 (O_1320,N_19826,N_18554);
and UO_1321 (O_1321,N_17754,N_17427);
and UO_1322 (O_1322,N_17628,N_18060);
nand UO_1323 (O_1323,N_17924,N_18543);
nor UO_1324 (O_1324,N_19576,N_17370);
or UO_1325 (O_1325,N_18521,N_18333);
nor UO_1326 (O_1326,N_19955,N_17207);
nor UO_1327 (O_1327,N_18399,N_19145);
and UO_1328 (O_1328,N_16056,N_16418);
nor UO_1329 (O_1329,N_16961,N_18279);
and UO_1330 (O_1330,N_19411,N_18128);
or UO_1331 (O_1331,N_17468,N_16607);
or UO_1332 (O_1332,N_17392,N_16197);
nor UO_1333 (O_1333,N_16846,N_17992);
nor UO_1334 (O_1334,N_18013,N_19287);
nand UO_1335 (O_1335,N_16417,N_18795);
or UO_1336 (O_1336,N_17863,N_17664);
or UO_1337 (O_1337,N_18139,N_16700);
and UO_1338 (O_1338,N_18109,N_19489);
nor UO_1339 (O_1339,N_18765,N_19418);
nor UO_1340 (O_1340,N_18406,N_18682);
or UO_1341 (O_1341,N_19095,N_17991);
nand UO_1342 (O_1342,N_18723,N_18811);
or UO_1343 (O_1343,N_19853,N_19334);
or UO_1344 (O_1344,N_18921,N_16789);
and UO_1345 (O_1345,N_19124,N_17271);
nand UO_1346 (O_1346,N_16871,N_17051);
or UO_1347 (O_1347,N_17462,N_16824);
and UO_1348 (O_1348,N_19774,N_18001);
nor UO_1349 (O_1349,N_18266,N_17591);
nand UO_1350 (O_1350,N_17422,N_18409);
xor UO_1351 (O_1351,N_19062,N_18434);
or UO_1352 (O_1352,N_16231,N_19989);
or UO_1353 (O_1353,N_16747,N_19603);
and UO_1354 (O_1354,N_17516,N_19212);
and UO_1355 (O_1355,N_19711,N_19125);
nand UO_1356 (O_1356,N_16593,N_16859);
and UO_1357 (O_1357,N_16189,N_17867);
nor UO_1358 (O_1358,N_19912,N_17058);
nor UO_1359 (O_1359,N_16321,N_17345);
nor UO_1360 (O_1360,N_16947,N_18131);
nor UO_1361 (O_1361,N_17397,N_16027);
and UO_1362 (O_1362,N_16112,N_17913);
nor UO_1363 (O_1363,N_18738,N_16673);
and UO_1364 (O_1364,N_16444,N_17425);
and UO_1365 (O_1365,N_17226,N_17053);
or UO_1366 (O_1366,N_18708,N_16156);
and UO_1367 (O_1367,N_18206,N_19780);
nand UO_1368 (O_1368,N_17122,N_17342);
nand UO_1369 (O_1369,N_16305,N_16230);
nor UO_1370 (O_1370,N_19319,N_17046);
nor UO_1371 (O_1371,N_17214,N_19524);
or UO_1372 (O_1372,N_18389,N_16353);
nor UO_1373 (O_1373,N_18295,N_18235);
nand UO_1374 (O_1374,N_19490,N_16907);
nor UO_1375 (O_1375,N_19498,N_17391);
and UO_1376 (O_1376,N_16026,N_19816);
nor UO_1377 (O_1377,N_17499,N_18510);
nand UO_1378 (O_1378,N_17946,N_18780);
nor UO_1379 (O_1379,N_19387,N_18142);
nand UO_1380 (O_1380,N_19394,N_16685);
or UO_1381 (O_1381,N_18968,N_18976);
xor UO_1382 (O_1382,N_18227,N_18054);
nor UO_1383 (O_1383,N_18574,N_17115);
or UO_1384 (O_1384,N_19015,N_19504);
and UO_1385 (O_1385,N_19825,N_18803);
nor UO_1386 (O_1386,N_19305,N_19150);
and UO_1387 (O_1387,N_17351,N_17793);
nand UO_1388 (O_1388,N_17685,N_18489);
or UO_1389 (O_1389,N_18387,N_19416);
or UO_1390 (O_1390,N_16895,N_17169);
and UO_1391 (O_1391,N_17162,N_19701);
nor UO_1392 (O_1392,N_18269,N_17997);
xnor UO_1393 (O_1393,N_18483,N_17014);
xor UO_1394 (O_1394,N_16040,N_18535);
and UO_1395 (O_1395,N_18505,N_18665);
nor UO_1396 (O_1396,N_16960,N_19988);
and UO_1397 (O_1397,N_19827,N_19011);
xnor UO_1398 (O_1398,N_18226,N_17543);
and UO_1399 (O_1399,N_18832,N_17891);
nor UO_1400 (O_1400,N_17488,N_16174);
nand UO_1401 (O_1401,N_17317,N_19595);
nor UO_1402 (O_1402,N_19136,N_19918);
nand UO_1403 (O_1403,N_17478,N_16582);
and UO_1404 (O_1404,N_18783,N_16476);
and UO_1405 (O_1405,N_16589,N_16104);
or UO_1406 (O_1406,N_19681,N_16579);
nand UO_1407 (O_1407,N_19852,N_19073);
and UO_1408 (O_1408,N_19981,N_16745);
nand UO_1409 (O_1409,N_16713,N_19656);
nand UO_1410 (O_1410,N_16235,N_18352);
nor UO_1411 (O_1411,N_17932,N_17288);
nand UO_1412 (O_1412,N_17842,N_17838);
nor UO_1413 (O_1413,N_16992,N_16680);
nand UO_1414 (O_1414,N_16946,N_19786);
nand UO_1415 (O_1415,N_17865,N_16843);
and UO_1416 (O_1416,N_16743,N_19960);
nand UO_1417 (O_1417,N_16212,N_16815);
or UO_1418 (O_1418,N_19219,N_19594);
and UO_1419 (O_1419,N_17795,N_17023);
nor UO_1420 (O_1420,N_19654,N_17728);
and UO_1421 (O_1421,N_18099,N_18951);
and UO_1422 (O_1422,N_18171,N_17999);
and UO_1423 (O_1423,N_16063,N_16359);
nand UO_1424 (O_1424,N_19091,N_18915);
nand UO_1425 (O_1425,N_19048,N_18444);
nand UO_1426 (O_1426,N_17232,N_19297);
or UO_1427 (O_1427,N_19412,N_18432);
nand UO_1428 (O_1428,N_17802,N_18668);
nor UO_1429 (O_1429,N_18412,N_19793);
nand UO_1430 (O_1430,N_16650,N_19924);
and UO_1431 (O_1431,N_19970,N_16784);
nor UO_1432 (O_1432,N_19107,N_18114);
nor UO_1433 (O_1433,N_16245,N_16018);
nand UO_1434 (O_1434,N_19733,N_17831);
and UO_1435 (O_1435,N_17311,N_16567);
and UO_1436 (O_1436,N_18584,N_18636);
and UO_1437 (O_1437,N_18029,N_16858);
nor UO_1438 (O_1438,N_18263,N_18924);
or UO_1439 (O_1439,N_17553,N_17809);
nor UO_1440 (O_1440,N_16785,N_18138);
nor UO_1441 (O_1441,N_17158,N_17073);
nand UO_1442 (O_1442,N_18475,N_19821);
or UO_1443 (O_1443,N_19167,N_17811);
nand UO_1444 (O_1444,N_19259,N_16536);
xor UO_1445 (O_1445,N_17661,N_18260);
and UO_1446 (O_1446,N_16330,N_19433);
and UO_1447 (O_1447,N_16549,N_19957);
nor UO_1448 (O_1448,N_18373,N_17797);
xnor UO_1449 (O_1449,N_17147,N_18004);
xnor UO_1450 (O_1450,N_19415,N_18716);
and UO_1451 (O_1451,N_16996,N_17306);
or UO_1452 (O_1452,N_18497,N_16880);
and UO_1453 (O_1453,N_17186,N_16297);
xnor UO_1454 (O_1454,N_16484,N_19894);
and UO_1455 (O_1455,N_17630,N_17604);
and UO_1456 (O_1456,N_19706,N_19344);
nand UO_1457 (O_1457,N_17741,N_16638);
nand UO_1458 (O_1458,N_17050,N_16926);
nor UO_1459 (O_1459,N_16908,N_18282);
nor UO_1460 (O_1460,N_18264,N_18914);
or UO_1461 (O_1461,N_17569,N_16176);
or UO_1462 (O_1462,N_17723,N_19231);
or UO_1463 (O_1463,N_16070,N_17283);
and UO_1464 (O_1464,N_19183,N_17602);
nor UO_1465 (O_1465,N_18699,N_17165);
or UO_1466 (O_1466,N_17452,N_19735);
nor UO_1467 (O_1467,N_18632,N_17568);
xnor UO_1468 (O_1468,N_19354,N_16006);
and UO_1469 (O_1469,N_19895,N_19540);
and UO_1470 (O_1470,N_18882,N_18885);
nor UO_1471 (O_1471,N_17168,N_17233);
nor UO_1472 (O_1472,N_17692,N_18429);
and UO_1473 (O_1473,N_18228,N_19291);
or UO_1474 (O_1474,N_16623,N_19440);
nor UO_1475 (O_1475,N_19434,N_17585);
nor UO_1476 (O_1476,N_16665,N_18778);
and UO_1477 (O_1477,N_19362,N_17076);
nand UO_1478 (O_1478,N_19634,N_16611);
nor UO_1479 (O_1479,N_17259,N_19465);
and UO_1480 (O_1480,N_18464,N_19527);
and UO_1481 (O_1481,N_19342,N_19128);
nand UO_1482 (O_1482,N_16774,N_18490);
and UO_1483 (O_1483,N_18729,N_18761);
nor UO_1484 (O_1484,N_19222,N_18443);
or UO_1485 (O_1485,N_16909,N_19386);
or UO_1486 (O_1486,N_18256,N_18462);
or UO_1487 (O_1487,N_19072,N_19742);
or UO_1488 (O_1488,N_16728,N_17676);
nor UO_1489 (O_1489,N_19916,N_17964);
and UO_1490 (O_1490,N_16318,N_19023);
nor UO_1491 (O_1491,N_18807,N_16875);
nor UO_1492 (O_1492,N_18485,N_18125);
or UO_1493 (O_1493,N_18839,N_17581);
nand UO_1494 (O_1494,N_19610,N_17031);
and UO_1495 (O_1495,N_18527,N_17206);
and UO_1496 (O_1496,N_19958,N_16655);
nor UO_1497 (O_1497,N_18602,N_19942);
and UO_1498 (O_1498,N_18714,N_17609);
nor UO_1499 (O_1499,N_17321,N_16327);
or UO_1500 (O_1500,N_16816,N_17901);
or UO_1501 (O_1501,N_18693,N_16347);
or UO_1502 (O_1502,N_16196,N_19583);
xor UO_1503 (O_1503,N_18010,N_19752);
or UO_1504 (O_1504,N_19553,N_16409);
and UO_1505 (O_1505,N_19380,N_18424);
nor UO_1506 (O_1506,N_19830,N_18639);
nand UO_1507 (O_1507,N_19986,N_18834);
and UO_1508 (O_1508,N_17829,N_18894);
nand UO_1509 (O_1509,N_17309,N_16286);
nand UO_1510 (O_1510,N_17762,N_19592);
and UO_1511 (O_1511,N_19607,N_18797);
or UO_1512 (O_1512,N_17535,N_18290);
or UO_1513 (O_1513,N_19577,N_16064);
and UO_1514 (O_1514,N_16089,N_18183);
or UO_1515 (O_1515,N_16280,N_19637);
nand UO_1516 (O_1516,N_18101,N_18694);
nand UO_1517 (O_1517,N_16339,N_16499);
and UO_1518 (O_1518,N_19608,N_17220);
or UO_1519 (O_1519,N_17121,N_19806);
or UO_1520 (O_1520,N_16081,N_16791);
nand UO_1521 (O_1521,N_16504,N_16322);
nand UO_1522 (O_1522,N_17771,N_16107);
nor UO_1523 (O_1523,N_19938,N_17238);
or UO_1524 (O_1524,N_16702,N_19493);
nand UO_1525 (O_1525,N_18709,N_17982);
or UO_1526 (O_1526,N_16819,N_17965);
and UO_1527 (O_1527,N_19077,N_19296);
and UO_1528 (O_1528,N_19085,N_17858);
or UO_1529 (O_1529,N_18878,N_18085);
and UO_1530 (O_1530,N_19228,N_16726);
nor UO_1531 (O_1531,N_16552,N_17533);
or UO_1532 (O_1532,N_19066,N_16950);
or UO_1533 (O_1533,N_16869,N_17745);
and UO_1534 (O_1534,N_19624,N_16414);
or UO_1535 (O_1535,N_19239,N_16471);
and UO_1536 (O_1536,N_17020,N_16464);
or UO_1537 (O_1537,N_18038,N_18037);
nand UO_1538 (O_1538,N_16348,N_19338);
or UO_1539 (O_1539,N_19995,N_17085);
or UO_1540 (O_1540,N_16034,N_17307);
and UO_1541 (O_1541,N_17343,N_19013);
nor UO_1542 (O_1542,N_19313,N_18238);
nand UO_1543 (O_1543,N_16735,N_17029);
or UO_1544 (O_1544,N_16394,N_19848);
and UO_1545 (O_1545,N_19134,N_19930);
or UO_1546 (O_1546,N_18458,N_18067);
nand UO_1547 (O_1547,N_16894,N_16714);
or UO_1548 (O_1548,N_17671,N_18617);
or UO_1549 (O_1549,N_18509,N_18261);
or UO_1550 (O_1550,N_17626,N_17770);
nor UO_1551 (O_1551,N_17083,N_17406);
or UO_1552 (O_1552,N_16844,N_16220);
or UO_1553 (O_1553,N_16146,N_16838);
and UO_1554 (O_1554,N_19197,N_18884);
nand UO_1555 (O_1555,N_19737,N_16387);
nor UO_1556 (O_1556,N_16820,N_17790);
and UO_1557 (O_1557,N_16386,N_17993);
or UO_1558 (O_1558,N_19148,N_19833);
or UO_1559 (O_1559,N_16634,N_19365);
or UO_1560 (O_1560,N_18035,N_19604);
nor UO_1561 (O_1561,N_18689,N_16390);
and UO_1562 (O_1562,N_17128,N_18230);
and UO_1563 (O_1563,N_18320,N_16059);
nor UO_1564 (O_1564,N_16559,N_18150);
nor UO_1565 (O_1565,N_16993,N_16051);
or UO_1566 (O_1566,N_16503,N_19070);
or UO_1567 (O_1567,N_17019,N_16315);
nand UO_1568 (O_1568,N_19823,N_19645);
and UO_1569 (O_1569,N_17286,N_19398);
and UO_1570 (O_1570,N_19809,N_19515);
nand UO_1571 (O_1571,N_19193,N_17336);
or UO_1572 (O_1572,N_19255,N_19230);
or UO_1573 (O_1573,N_17048,N_17724);
or UO_1574 (O_1574,N_17194,N_17257);
and UO_1575 (O_1575,N_17864,N_16622);
nand UO_1576 (O_1576,N_19710,N_17328);
nand UO_1577 (O_1577,N_16029,N_18508);
nor UO_1578 (O_1578,N_17837,N_17285);
nor UO_1579 (O_1579,N_19945,N_18966);
nor UO_1580 (O_1580,N_19522,N_19939);
nor UO_1581 (O_1581,N_16678,N_18986);
nand UO_1582 (O_1582,N_17862,N_19133);
and UO_1583 (O_1583,N_17000,N_19686);
or UO_1584 (O_1584,N_18747,N_19478);
or UO_1585 (O_1585,N_18191,N_18242);
nor UO_1586 (O_1586,N_18323,N_18760);
and UO_1587 (O_1587,N_17322,N_16097);
or UO_1588 (O_1588,N_19149,N_17152);
nor UO_1589 (O_1589,N_18073,N_18670);
nor UO_1590 (O_1590,N_17149,N_17761);
xnor UO_1591 (O_1591,N_19339,N_19050);
and UO_1592 (O_1592,N_17094,N_16957);
or UO_1593 (O_1593,N_16830,N_18286);
nor UO_1594 (O_1594,N_17313,N_19397);
nand UO_1595 (O_1595,N_19378,N_17086);
or UO_1596 (O_1596,N_18375,N_17611);
and UO_1597 (O_1597,N_17277,N_18938);
nand UO_1598 (O_1598,N_17743,N_18982);
nand UO_1599 (O_1599,N_19712,N_16410);
nor UO_1600 (O_1600,N_18784,N_19781);
and UO_1601 (O_1601,N_18451,N_17618);
nand UO_1602 (O_1602,N_19105,N_19014);
or UO_1603 (O_1603,N_17562,N_16301);
nand UO_1604 (O_1604,N_18692,N_18904);
nor UO_1605 (O_1605,N_18477,N_19087);
and UO_1606 (O_1606,N_17481,N_16108);
nand UO_1607 (O_1607,N_18837,N_16692);
or UO_1608 (O_1608,N_17235,N_17282);
or UO_1609 (O_1609,N_19675,N_16794);
xnor UO_1610 (O_1610,N_19221,N_18106);
nand UO_1611 (O_1611,N_18381,N_16289);
nand UO_1612 (O_1612,N_19207,N_19471);
and UO_1613 (O_1613,N_19714,N_16184);
nand UO_1614 (O_1614,N_17940,N_16013);
and UO_1615 (O_1615,N_19217,N_18852);
nor UO_1616 (O_1616,N_17205,N_17487);
nor UO_1617 (O_1617,N_19352,N_17136);
nand UO_1618 (O_1618,N_18641,N_19363);
and UO_1619 (O_1619,N_17643,N_19967);
and UO_1620 (O_1620,N_16137,N_18571);
nor UO_1621 (O_1621,N_17709,N_18423);
and UO_1622 (O_1622,N_19461,N_16475);
nor UO_1623 (O_1623,N_18506,N_16192);
and UO_1624 (O_1624,N_16269,N_18645);
nand UO_1625 (O_1625,N_17588,N_17250);
or UO_1626 (O_1626,N_17780,N_18441);
xor UO_1627 (O_1627,N_16518,N_18340);
nand UO_1628 (O_1628,N_19532,N_16256);
and UO_1629 (O_1629,N_16868,N_16253);
and UO_1630 (O_1630,N_19846,N_17950);
and UO_1631 (O_1631,N_17911,N_16468);
nand UO_1632 (O_1632,N_16765,N_16420);
nand UO_1633 (O_1633,N_18158,N_17386);
and UO_1634 (O_1634,N_18057,N_16801);
or UO_1635 (O_1635,N_19856,N_18724);
or UO_1636 (O_1636,N_16524,N_16594);
nand UO_1637 (O_1637,N_17632,N_17044);
or UO_1638 (O_1638,N_18194,N_17953);
or UO_1639 (O_1639,N_17861,N_17244);
nor UO_1640 (O_1640,N_19621,N_19552);
and UO_1641 (O_1641,N_18932,N_17272);
and UO_1642 (O_1642,N_18949,N_17415);
or UO_1643 (O_1643,N_16037,N_17691);
nor UO_1644 (O_1644,N_16225,N_18701);
nor UO_1645 (O_1645,N_17090,N_16730);
or UO_1646 (O_1646,N_16227,N_19405);
nand UO_1647 (O_1647,N_17361,N_16141);
or UO_1648 (O_1648,N_16585,N_16003);
nand UO_1649 (O_1649,N_18883,N_17582);
or UO_1650 (O_1650,N_17189,N_19120);
nor UO_1651 (O_1651,N_18061,N_16232);
or UO_1652 (O_1652,N_17477,N_17693);
nand UO_1653 (O_1653,N_18922,N_16509);
nand UO_1654 (O_1654,N_19375,N_19312);
or UO_1655 (O_1655,N_18439,N_17875);
and UO_1656 (O_1656,N_16325,N_17445);
xor UO_1657 (O_1657,N_19695,N_18558);
nor UO_1658 (O_1658,N_17049,N_18145);
and UO_1659 (O_1659,N_18786,N_17615);
and UO_1660 (O_1660,N_17131,N_17814);
and UO_1661 (O_1661,N_17242,N_19158);
nand UO_1662 (O_1662,N_19881,N_18124);
nor UO_1663 (O_1663,N_16311,N_16042);
or UO_1664 (O_1664,N_19457,N_18940);
nand UO_1665 (O_1665,N_17622,N_19649);
xnor UO_1666 (O_1666,N_18630,N_19071);
and UO_1667 (O_1667,N_18860,N_17962);
nand UO_1668 (O_1668,N_18471,N_16148);
nor UO_1669 (O_1669,N_17906,N_17530);
or UO_1670 (O_1670,N_18110,N_19450);
and UO_1671 (O_1671,N_18161,N_17534);
nand UO_1672 (O_1672,N_19361,N_18311);
nor UO_1673 (O_1673,N_19832,N_18603);
and UO_1674 (O_1674,N_17787,N_19004);
nor UO_1675 (O_1675,N_17781,N_19620);
nand UO_1676 (O_1676,N_16989,N_16403);
or UO_1677 (O_1677,N_17039,N_18463);
nor UO_1678 (O_1678,N_18974,N_19469);
nand UO_1679 (O_1679,N_16925,N_18334);
nand UO_1680 (O_1680,N_17030,N_16060);
nor UO_1681 (O_1681,N_16138,N_17363);
or UO_1682 (O_1682,N_18843,N_16802);
nand UO_1683 (O_1683,N_18663,N_17130);
and UO_1684 (O_1684,N_17667,N_18606);
and UO_1685 (O_1685,N_19122,N_17234);
or UO_1686 (O_1686,N_17735,N_19093);
and UO_1687 (O_1687,N_18157,N_19570);
and UO_1688 (O_1688,N_18214,N_17625);
or UO_1689 (O_1689,N_17887,N_19837);
or UO_1690 (O_1690,N_16835,N_17714);
nor UO_1691 (O_1691,N_17432,N_17990);
or UO_1692 (O_1692,N_18766,N_18318);
xnor UO_1693 (O_1693,N_18916,N_17675);
and UO_1694 (O_1694,N_18769,N_17629);
xor UO_1695 (O_1695,N_17443,N_16383);
or UO_1696 (O_1696,N_18827,N_18534);
nor UO_1697 (O_1697,N_19410,N_19357);
xnor UO_1698 (O_1698,N_18893,N_17572);
or UO_1699 (O_1699,N_17912,N_17624);
or UO_1700 (O_1700,N_19025,N_16931);
nor UO_1701 (O_1701,N_17877,N_16555);
xor UO_1702 (O_1702,N_18195,N_17323);
and UO_1703 (O_1703,N_16033,N_19326);
and UO_1704 (O_1704,N_18514,N_16049);
and UO_1705 (O_1705,N_16492,N_18247);
nor UO_1706 (O_1706,N_18123,N_16973);
nand UO_1707 (O_1707,N_17346,N_18686);
nand UO_1708 (O_1708,N_19845,N_17098);
nor UO_1709 (O_1709,N_16917,N_16314);
and UO_1710 (O_1710,N_19103,N_19026);
nand UO_1711 (O_1711,N_19997,N_16647);
nor UO_1712 (O_1712,N_19160,N_19049);
and UO_1713 (O_1713,N_18871,N_17099);
xnor UO_1714 (O_1714,N_17704,N_19373);
and UO_1715 (O_1715,N_19249,N_17055);
nand UO_1716 (O_1716,N_18374,N_18524);
nand UO_1717 (O_1717,N_16573,N_16620);
xor UO_1718 (O_1718,N_16028,N_19250);
or UO_1719 (O_1719,N_18071,N_19283);
or UO_1720 (O_1720,N_18909,N_17788);
or UO_1721 (O_1721,N_18215,N_17291);
nor UO_1722 (O_1722,N_18259,N_19438);
nor UO_1723 (O_1723,N_17396,N_18581);
and UO_1724 (O_1724,N_18385,N_16298);
and UO_1725 (O_1725,N_16751,N_17393);
or UO_1726 (O_1726,N_19232,N_18072);
or UO_1727 (O_1727,N_17301,N_17663);
or UO_1728 (O_1728,N_17928,N_16812);
nand UO_1729 (O_1729,N_19356,N_16849);
nor UO_1730 (O_1730,N_18587,N_19462);
or UO_1731 (O_1731,N_18433,N_18274);
and UO_1732 (O_1732,N_19646,N_19208);
nor UO_1733 (O_1733,N_16570,N_17398);
and UO_1734 (O_1734,N_17062,N_16903);
and UO_1735 (O_1735,N_16335,N_18688);
nand UO_1736 (O_1736,N_16698,N_18201);
nor UO_1737 (O_1737,N_17008,N_17080);
or UO_1738 (O_1738,N_16440,N_19413);
and UO_1739 (O_1739,N_18687,N_17503);
or UO_1740 (O_1740,N_18635,N_17665);
nand UO_1741 (O_1741,N_19294,N_18984);
nand UO_1742 (O_1742,N_16384,N_17353);
xor UO_1743 (O_1743,N_16421,N_16891);
and UO_1744 (O_1744,N_16780,N_16672);
or UO_1745 (O_1745,N_18077,N_19985);
nor UO_1746 (O_1746,N_18546,N_17563);
xor UO_1747 (O_1747,N_19279,N_18681);
and UO_1748 (O_1748,N_18339,N_19161);
nand UO_1749 (O_1749,N_16309,N_16448);
and UO_1750 (O_1750,N_19758,N_17894);
nor UO_1751 (O_1751,N_16139,N_17647);
nor UO_1752 (O_1752,N_18545,N_17455);
nor UO_1753 (O_1753,N_18891,N_16065);
or UO_1754 (O_1754,N_17573,N_17583);
and UO_1755 (O_1755,N_19888,N_16879);
and UO_1756 (O_1756,N_19893,N_16945);
nand UO_1757 (O_1757,N_17619,N_16030);
nor UO_1758 (O_1758,N_16754,N_19783);
or UO_1759 (O_1759,N_16260,N_18100);
nor UO_1760 (O_1760,N_17970,N_16262);
nor UO_1761 (O_1761,N_17748,N_19458);
and UO_1762 (O_1762,N_16598,N_17679);
and UO_1763 (O_1763,N_16489,N_16841);
nand UO_1764 (O_1764,N_18008,N_19082);
nand UO_1765 (O_1765,N_18979,N_16516);
and UO_1766 (O_1766,N_18043,N_18562);
nand UO_1767 (O_1767,N_19949,N_19278);
or UO_1768 (O_1768,N_17340,N_19285);
nand UO_1769 (O_1769,N_16599,N_18192);
or UO_1770 (O_1770,N_18887,N_19006);
nor UO_1771 (O_1771,N_16109,N_17929);
xnor UO_1772 (O_1772,N_16244,N_16445);
or UO_1773 (O_1773,N_19677,N_17431);
nor UO_1774 (O_1774,N_17091,N_16603);
nand UO_1775 (O_1775,N_18050,N_19593);
or UO_1776 (O_1776,N_18697,N_18865);
and UO_1777 (O_1777,N_18049,N_18134);
nand UO_1778 (O_1778,N_16739,N_19765);
and UO_1779 (O_1779,N_18447,N_17718);
nand UO_1780 (O_1780,N_18002,N_17571);
and UO_1781 (O_1781,N_16760,N_17093);
and UO_1782 (O_1782,N_18499,N_17253);
nand UO_1783 (O_1783,N_16834,N_16273);
nand UO_1784 (O_1784,N_16039,N_19807);
nor UO_1785 (O_1785,N_17215,N_18056);
nand UO_1786 (O_1786,N_17209,N_17368);
nand UO_1787 (O_1787,N_17010,N_19314);
and UO_1788 (O_1788,N_17199,N_19962);
nor UO_1789 (O_1789,N_19099,N_18267);
and UO_1790 (O_1790,N_19743,N_16717);
or UO_1791 (O_1791,N_17551,N_17775);
nor UO_1792 (O_1792,N_18933,N_18023);
nor UO_1793 (O_1793,N_19705,N_17402);
xnor UO_1794 (O_1794,N_18472,N_18426);
nor UO_1795 (O_1795,N_17203,N_17384);
or UO_1796 (O_1796,N_17376,N_17768);
nor UO_1797 (O_1797,N_17739,N_19836);
and UO_1798 (O_1798,N_18625,N_18449);
or UO_1799 (O_1799,N_16173,N_17869);
or UO_1800 (O_1800,N_17484,N_19178);
nand UO_1801 (O_1801,N_16020,N_17976);
nand UO_1802 (O_1802,N_18999,N_19692);
nor UO_1803 (O_1803,N_18276,N_16814);
nor UO_1804 (O_1804,N_17159,N_18219);
nand UO_1805 (O_1805,N_19340,N_19899);
and UO_1806 (O_1806,N_17817,N_19482);
nor UO_1807 (O_1807,N_19612,N_16857);
or UO_1808 (O_1808,N_17528,N_16631);
xor UO_1809 (O_1809,N_19776,N_18637);
nand UO_1810 (O_1810,N_18599,N_19188);
or UO_1811 (O_1811,N_17150,N_17958);
or UO_1812 (O_1812,N_18825,N_18771);
and UO_1813 (O_1813,N_18133,N_17416);
nor UO_1814 (O_1814,N_19144,N_18879);
nor UO_1815 (O_1815,N_18116,N_17217);
or UO_1816 (O_1816,N_18923,N_19581);
nand UO_1817 (O_1817,N_18561,N_16190);
and UO_1818 (O_1818,N_16216,N_16568);
and UO_1819 (O_1819,N_17552,N_18643);
or UO_1820 (O_1820,N_19947,N_19382);
or UO_1821 (O_1821,N_18684,N_18417);
nand UO_1822 (O_1822,N_19858,N_18530);
or UO_1823 (O_1823,N_18177,N_19704);
nor UO_1824 (O_1824,N_18140,N_16152);
xnor UO_1825 (O_1825,N_19667,N_18309);
or UO_1826 (O_1826,N_17922,N_16772);
nor UO_1827 (O_1827,N_18187,N_18310);
nor UO_1828 (O_1828,N_16145,N_17909);
nand UO_1829 (O_1829,N_16542,N_19839);
or UO_1830 (O_1830,N_18300,N_17845);
nor UO_1831 (O_1831,N_19364,N_16419);
xor UO_1832 (O_1832,N_19056,N_16412);
and UO_1833 (O_1833,N_16062,N_17012);
nand UO_1834 (O_1834,N_19225,N_18055);
and UO_1835 (O_1835,N_19920,N_16642);
nand UO_1836 (O_1836,N_17002,N_19067);
and UO_1837 (O_1837,N_18608,N_18704);
or UO_1838 (O_1838,N_17874,N_16543);
xnor UO_1839 (O_1839,N_19155,N_18752);
nand UO_1840 (O_1840,N_18831,N_16681);
nand UO_1841 (O_1841,N_17985,N_17892);
nor UO_1842 (O_1842,N_17766,N_19052);
and UO_1843 (O_1843,N_18039,N_18148);
nor UO_1844 (O_1844,N_18448,N_17983);
or UO_1845 (O_1845,N_16804,N_19578);
nand UO_1846 (O_1846,N_17834,N_16123);
nand UO_1847 (O_1847,N_19165,N_17154);
or UO_1848 (O_1848,N_18255,N_19913);
nand UO_1849 (O_1849,N_17994,N_19260);
xnor UO_1850 (O_1850,N_17882,N_19841);
or UO_1851 (O_1851,N_19511,N_17559);
and UO_1852 (O_1852,N_16564,N_16328);
or UO_1853 (O_1853,N_16899,N_19590);
and UO_1854 (O_1854,N_17299,N_18750);
nand UO_1855 (O_1855,N_17851,N_18953);
nand UO_1856 (O_1856,N_19650,N_18787);
nand UO_1857 (O_1857,N_19080,N_16600);
and UO_1858 (O_1858,N_17139,N_18301);
and UO_1859 (O_1859,N_19320,N_18487);
nand UO_1860 (O_1860,N_18844,N_19520);
or UO_1861 (O_1861,N_18402,N_17961);
and UO_1862 (O_1862,N_19605,N_16704);
or UO_1863 (O_1863,N_16009,N_16119);
and UO_1864 (O_1864,N_16364,N_18221);
nand UO_1865 (O_1865,N_16613,N_16777);
or UO_1866 (O_1866,N_19036,N_19643);
or UO_1867 (O_1867,N_19102,N_17903);
and UO_1868 (O_1868,N_17229,N_19876);
and UO_1869 (O_1869,N_18720,N_16574);
nand UO_1870 (O_1870,N_19186,N_17702);
nand UO_1871 (O_1871,N_19035,N_18086);
nand UO_1872 (O_1872,N_16087,N_19257);
nor UO_1873 (O_1873,N_19928,N_17001);
nor UO_1874 (O_1874,N_17161,N_16584);
and UO_1875 (O_1875,N_17919,N_17065);
and UO_1876 (O_1876,N_18492,N_17171);
nor UO_1877 (O_1877,N_16208,N_16381);
and UO_1878 (O_1878,N_19055,N_19214);
nor UO_1879 (O_1879,N_18307,N_18437);
nor UO_1880 (O_1880,N_18170,N_19662);
nand UO_1881 (O_1881,N_18454,N_18151);
and UO_1882 (O_1882,N_19130,N_19247);
nand UO_1883 (O_1883,N_16632,N_16449);
nand UO_1884 (O_1884,N_18469,N_19802);
nand UO_1885 (O_1885,N_18137,N_18541);
and UO_1886 (O_1886,N_16737,N_16888);
and UO_1887 (O_1887,N_18993,N_16495);
and UO_1888 (O_1888,N_18518,N_17885);
nand UO_1889 (O_1889,N_18848,N_16446);
nand UO_1890 (O_1890,N_17251,N_17601);
or UO_1891 (O_1891,N_17866,N_17134);
or UO_1892 (O_1892,N_17558,N_16983);
nand UO_1893 (O_1893,N_16787,N_16275);
and UO_1894 (O_1894,N_17727,N_19950);
nand UO_1895 (O_1895,N_19979,N_17184);
or UO_1896 (O_1896,N_19991,N_19233);
xnor UO_1897 (O_1897,N_18368,N_19818);
and UO_1898 (O_1898,N_16900,N_17916);
or UO_1899 (O_1899,N_19505,N_19031);
and UO_1900 (O_1900,N_16833,N_16175);
or UO_1901 (O_1901,N_18482,N_16404);
nor UO_1902 (O_1902,N_19037,N_18159);
or UO_1903 (O_1903,N_19436,N_16498);
and UO_1904 (O_1904,N_17945,N_17515);
and UO_1905 (O_1905,N_19030,N_19770);
nand UO_1906 (O_1906,N_17219,N_18353);
or UO_1907 (O_1907,N_19753,N_18186);
or UO_1908 (O_1908,N_17703,N_18656);
nand UO_1909 (O_1909,N_19454,N_17358);
and UO_1910 (O_1910,N_19954,N_19346);
or UO_1911 (O_1911,N_17584,N_16099);
and UO_1912 (O_1912,N_18379,N_19980);
or UO_1913 (O_1913,N_19732,N_17201);
or UO_1914 (O_1914,N_19994,N_17608);
or UO_1915 (O_1915,N_18335,N_19383);
or UO_1916 (O_1916,N_18313,N_17900);
xor UO_1917 (O_1917,N_16276,N_17407);
and UO_1918 (O_1918,N_19258,N_16371);
and UO_1919 (O_1919,N_18898,N_18502);
nor UO_1920 (O_1920,N_16374,N_18118);
and UO_1921 (O_1921,N_18718,N_17957);
nand UO_1922 (O_1922,N_19273,N_18239);
and UO_1923 (O_1923,N_16716,N_18341);
or UO_1924 (O_1924,N_19492,N_18149);
or UO_1925 (O_1925,N_18355,N_17153);
and UO_1926 (O_1926,N_18450,N_16539);
xor UO_1927 (O_1927,N_19078,N_17649);
nand UO_1928 (O_1928,N_16558,N_18349);
nor UO_1929 (O_1929,N_17292,N_17896);
nor UO_1930 (O_1930,N_17725,N_18204);
and UO_1931 (O_1931,N_16767,N_17439);
nor UO_1932 (O_1932,N_16727,N_17308);
nor UO_1933 (O_1933,N_19198,N_16379);
nand UO_1934 (O_1934,N_18845,N_18609);
nand UO_1935 (O_1935,N_18596,N_19266);
nor UO_1936 (O_1936,N_18655,N_17753);
and UO_1937 (O_1937,N_17175,N_17326);
or UO_1938 (O_1938,N_16272,N_18246);
or UO_1939 (O_1939,N_16057,N_19850);
or UO_1940 (O_1940,N_16644,N_16577);
and UO_1941 (O_1941,N_16134,N_17509);
nand UO_1942 (O_1942,N_18181,N_17642);
or UO_1943 (O_1943,N_17942,N_19104);
and UO_1944 (O_1944,N_19315,N_16526);
or UO_1945 (O_1945,N_16691,N_18386);
nor UO_1946 (O_1946,N_18456,N_16657);
nor UO_1947 (O_1947,N_19053,N_16124);
nand UO_1948 (O_1948,N_19310,N_16682);
xnor UO_1949 (O_1949,N_19529,N_16369);
nand UO_1950 (O_1950,N_18362,N_17578);
nor UO_1951 (O_1951,N_19045,N_16163);
and UO_1952 (O_1952,N_18867,N_16610);
nor UO_1953 (O_1953,N_19944,N_18973);
or UO_1954 (O_1954,N_19526,N_19427);
nor UO_1955 (O_1955,N_16077,N_19046);
xor UO_1956 (O_1956,N_16786,N_16239);
nor UO_1957 (O_1957,N_18236,N_16654);
or UO_1958 (O_1958,N_16485,N_17333);
or UO_1959 (O_1959,N_19166,N_16224);
or UO_1960 (O_1960,N_19393,N_17921);
or UO_1961 (O_1961,N_18425,N_17792);
nand UO_1962 (O_1962,N_16757,N_17295);
nor UO_1963 (O_1963,N_17644,N_17036);
nand UO_1964 (O_1964,N_16164,N_17212);
or UO_1965 (O_1965,N_17759,N_16972);
nor UO_1966 (O_1966,N_16125,N_16019);
or UO_1967 (O_1967,N_17767,N_17352);
nor UO_1968 (O_1968,N_16625,N_19953);
nor UO_1969 (O_1969,N_17816,N_16848);
nand UO_1970 (O_1970,N_18824,N_19445);
and UO_1971 (O_1971,N_17371,N_18996);
or UO_1972 (O_1972,N_16031,N_16050);
nor UO_1973 (O_1973,N_18816,N_19311);
nor UO_1974 (O_1974,N_17786,N_18273);
nor UO_1975 (O_1975,N_18303,N_19693);
or UO_1976 (O_1976,N_18667,N_18292);
nand UO_1977 (O_1977,N_18094,N_19396);
or UO_1978 (O_1978,N_19425,N_19665);
nand UO_1979 (O_1979,N_18965,N_18773);
nor UO_1980 (O_1980,N_19952,N_19151);
and UO_1981 (O_1981,N_19933,N_17469);
and UO_1982 (O_1982,N_18768,N_19184);
xor UO_1983 (O_1983,N_19110,N_19869);
and UO_1984 (O_1984,N_17832,N_17975);
nand UO_1985 (O_1985,N_18758,N_19754);
nor UO_1986 (O_1986,N_19935,N_17555);
xor UO_1987 (O_1987,N_16565,N_19946);
nand UO_1988 (O_1988,N_19937,N_16310);
and UO_1989 (O_1989,N_18220,N_19983);
nor UO_1990 (O_1990,N_17394,N_16361);
nor UO_1991 (O_1991,N_18212,N_16718);
nor UO_1992 (O_1992,N_18648,N_16496);
or UO_1993 (O_1993,N_17163,N_18550);
nor UO_1994 (O_1994,N_17658,N_16254);
and UO_1995 (O_1995,N_18796,N_19281);
or UO_1996 (O_1996,N_16093,N_18698);
or UO_1997 (O_1997,N_16183,N_19051);
nor UO_1998 (O_1998,N_17247,N_16646);
nor UO_1999 (O_1999,N_17820,N_18743);
nor UO_2000 (O_2000,N_17956,N_18136);
nand UO_2001 (O_2001,N_17150,N_16811);
and UO_2002 (O_2002,N_17042,N_16557);
and UO_2003 (O_2003,N_16311,N_19255);
or UO_2004 (O_2004,N_19153,N_16383);
or UO_2005 (O_2005,N_19435,N_16748);
and UO_2006 (O_2006,N_19662,N_19466);
and UO_2007 (O_2007,N_17392,N_17447);
nor UO_2008 (O_2008,N_17519,N_19386);
nor UO_2009 (O_2009,N_19304,N_18444);
and UO_2010 (O_2010,N_18637,N_16262);
or UO_2011 (O_2011,N_16987,N_16016);
and UO_2012 (O_2012,N_18904,N_17160);
nand UO_2013 (O_2013,N_16578,N_16233);
nand UO_2014 (O_2014,N_19961,N_16687);
or UO_2015 (O_2015,N_16211,N_18350);
nand UO_2016 (O_2016,N_18648,N_19908);
nor UO_2017 (O_2017,N_19857,N_16162);
nor UO_2018 (O_2018,N_18373,N_18400);
and UO_2019 (O_2019,N_19166,N_17087);
nor UO_2020 (O_2020,N_19076,N_19713);
nand UO_2021 (O_2021,N_18612,N_19262);
nand UO_2022 (O_2022,N_17098,N_17448);
nor UO_2023 (O_2023,N_19813,N_16911);
and UO_2024 (O_2024,N_19415,N_19527);
or UO_2025 (O_2025,N_17266,N_19715);
nor UO_2026 (O_2026,N_18960,N_16114);
and UO_2027 (O_2027,N_19273,N_16110);
nand UO_2028 (O_2028,N_18503,N_17587);
nand UO_2029 (O_2029,N_18497,N_18243);
nor UO_2030 (O_2030,N_16457,N_18497);
nand UO_2031 (O_2031,N_17791,N_16091);
and UO_2032 (O_2032,N_17672,N_17786);
and UO_2033 (O_2033,N_19839,N_16986);
nand UO_2034 (O_2034,N_19983,N_19718);
or UO_2035 (O_2035,N_18574,N_19668);
nand UO_2036 (O_2036,N_19705,N_17650);
or UO_2037 (O_2037,N_16932,N_18019);
nor UO_2038 (O_2038,N_17162,N_17958);
and UO_2039 (O_2039,N_17976,N_19726);
nand UO_2040 (O_2040,N_19630,N_18660);
and UO_2041 (O_2041,N_18167,N_19362);
nor UO_2042 (O_2042,N_18054,N_19094);
nand UO_2043 (O_2043,N_19328,N_17257);
and UO_2044 (O_2044,N_16119,N_17637);
nand UO_2045 (O_2045,N_16481,N_16356);
and UO_2046 (O_2046,N_16860,N_17161);
nand UO_2047 (O_2047,N_17574,N_19598);
nor UO_2048 (O_2048,N_16889,N_16473);
and UO_2049 (O_2049,N_16484,N_18060);
or UO_2050 (O_2050,N_17532,N_17836);
nand UO_2051 (O_2051,N_17722,N_17884);
or UO_2052 (O_2052,N_19216,N_19867);
or UO_2053 (O_2053,N_17269,N_19494);
or UO_2054 (O_2054,N_19245,N_16055);
nor UO_2055 (O_2055,N_19764,N_18921);
xor UO_2056 (O_2056,N_18636,N_16121);
and UO_2057 (O_2057,N_18156,N_19869);
nand UO_2058 (O_2058,N_16087,N_18201);
or UO_2059 (O_2059,N_18472,N_16086);
or UO_2060 (O_2060,N_17189,N_17120);
nor UO_2061 (O_2061,N_18423,N_17851);
and UO_2062 (O_2062,N_18158,N_18711);
or UO_2063 (O_2063,N_18315,N_18375);
nor UO_2064 (O_2064,N_18219,N_18579);
or UO_2065 (O_2065,N_19212,N_16422);
nand UO_2066 (O_2066,N_18363,N_17057);
nand UO_2067 (O_2067,N_19903,N_18019);
nor UO_2068 (O_2068,N_17449,N_16011);
and UO_2069 (O_2069,N_17712,N_17696);
and UO_2070 (O_2070,N_18227,N_16353);
and UO_2071 (O_2071,N_18887,N_17001);
or UO_2072 (O_2072,N_19523,N_18842);
or UO_2073 (O_2073,N_19852,N_17159);
nand UO_2074 (O_2074,N_19772,N_17132);
or UO_2075 (O_2075,N_16736,N_19938);
nand UO_2076 (O_2076,N_18857,N_17414);
nand UO_2077 (O_2077,N_17475,N_19478);
and UO_2078 (O_2078,N_17542,N_18047);
xor UO_2079 (O_2079,N_18868,N_17862);
and UO_2080 (O_2080,N_19780,N_18117);
nor UO_2081 (O_2081,N_16471,N_16863);
nor UO_2082 (O_2082,N_19274,N_16164);
and UO_2083 (O_2083,N_18133,N_19799);
or UO_2084 (O_2084,N_16221,N_18043);
nor UO_2085 (O_2085,N_17322,N_16316);
and UO_2086 (O_2086,N_17687,N_17904);
nand UO_2087 (O_2087,N_17441,N_19363);
or UO_2088 (O_2088,N_19761,N_16650);
nand UO_2089 (O_2089,N_18102,N_17605);
or UO_2090 (O_2090,N_16798,N_16724);
or UO_2091 (O_2091,N_16661,N_19720);
nor UO_2092 (O_2092,N_17724,N_19774);
nand UO_2093 (O_2093,N_16145,N_19275);
or UO_2094 (O_2094,N_17399,N_18273);
and UO_2095 (O_2095,N_18913,N_17410);
nand UO_2096 (O_2096,N_19293,N_17988);
or UO_2097 (O_2097,N_19760,N_19331);
nor UO_2098 (O_2098,N_17372,N_16306);
nor UO_2099 (O_2099,N_19390,N_17300);
or UO_2100 (O_2100,N_18053,N_19929);
nand UO_2101 (O_2101,N_18363,N_17423);
and UO_2102 (O_2102,N_19303,N_19859);
or UO_2103 (O_2103,N_19152,N_19374);
nor UO_2104 (O_2104,N_19141,N_18675);
or UO_2105 (O_2105,N_17886,N_16757);
nor UO_2106 (O_2106,N_17068,N_18211);
nand UO_2107 (O_2107,N_18827,N_17335);
nor UO_2108 (O_2108,N_19225,N_18045);
or UO_2109 (O_2109,N_17460,N_19875);
nor UO_2110 (O_2110,N_19240,N_17506);
nor UO_2111 (O_2111,N_17786,N_17231);
nor UO_2112 (O_2112,N_18990,N_16424);
or UO_2113 (O_2113,N_18422,N_17077);
or UO_2114 (O_2114,N_19939,N_18831);
and UO_2115 (O_2115,N_19851,N_17749);
nor UO_2116 (O_2116,N_17108,N_18630);
nor UO_2117 (O_2117,N_17254,N_19515);
and UO_2118 (O_2118,N_17953,N_18078);
and UO_2119 (O_2119,N_19870,N_17824);
nand UO_2120 (O_2120,N_16121,N_16716);
nand UO_2121 (O_2121,N_19253,N_19338);
and UO_2122 (O_2122,N_19380,N_16744);
and UO_2123 (O_2123,N_17789,N_18722);
nor UO_2124 (O_2124,N_18057,N_17865);
nor UO_2125 (O_2125,N_16340,N_18372);
nand UO_2126 (O_2126,N_16335,N_16702);
nor UO_2127 (O_2127,N_18112,N_17221);
xnor UO_2128 (O_2128,N_18333,N_16019);
nor UO_2129 (O_2129,N_18521,N_17124);
and UO_2130 (O_2130,N_17550,N_17945);
nand UO_2131 (O_2131,N_17745,N_16579);
nor UO_2132 (O_2132,N_17723,N_18196);
or UO_2133 (O_2133,N_17014,N_16586);
and UO_2134 (O_2134,N_19455,N_19917);
nor UO_2135 (O_2135,N_16997,N_17522);
xnor UO_2136 (O_2136,N_18237,N_18639);
or UO_2137 (O_2137,N_17345,N_18345);
nand UO_2138 (O_2138,N_16956,N_18748);
and UO_2139 (O_2139,N_17602,N_18979);
or UO_2140 (O_2140,N_16361,N_19672);
and UO_2141 (O_2141,N_19410,N_19023);
nand UO_2142 (O_2142,N_18619,N_16345);
nand UO_2143 (O_2143,N_17340,N_16482);
nor UO_2144 (O_2144,N_16071,N_17292);
and UO_2145 (O_2145,N_17826,N_19096);
nand UO_2146 (O_2146,N_19801,N_19069);
nand UO_2147 (O_2147,N_17012,N_18514);
or UO_2148 (O_2148,N_17043,N_18284);
nor UO_2149 (O_2149,N_19822,N_17181);
nand UO_2150 (O_2150,N_18644,N_18902);
nand UO_2151 (O_2151,N_17089,N_17265);
nor UO_2152 (O_2152,N_17000,N_16170);
nor UO_2153 (O_2153,N_18844,N_18786);
or UO_2154 (O_2154,N_18804,N_19249);
nand UO_2155 (O_2155,N_16156,N_16526);
nand UO_2156 (O_2156,N_17421,N_19924);
and UO_2157 (O_2157,N_17027,N_16914);
nand UO_2158 (O_2158,N_17385,N_17696);
and UO_2159 (O_2159,N_17903,N_18860);
nand UO_2160 (O_2160,N_16049,N_18249);
nor UO_2161 (O_2161,N_17266,N_16624);
nor UO_2162 (O_2162,N_19051,N_17688);
and UO_2163 (O_2163,N_18674,N_17831);
or UO_2164 (O_2164,N_16348,N_16950);
nor UO_2165 (O_2165,N_16411,N_19565);
and UO_2166 (O_2166,N_18076,N_16147);
xor UO_2167 (O_2167,N_18242,N_17731);
and UO_2168 (O_2168,N_18526,N_17697);
nor UO_2169 (O_2169,N_16863,N_19753);
or UO_2170 (O_2170,N_19617,N_17606);
nor UO_2171 (O_2171,N_18764,N_18104);
nor UO_2172 (O_2172,N_17814,N_16104);
nor UO_2173 (O_2173,N_19567,N_16207);
nand UO_2174 (O_2174,N_16378,N_16376);
nor UO_2175 (O_2175,N_16740,N_18764);
and UO_2176 (O_2176,N_16474,N_16115);
or UO_2177 (O_2177,N_19463,N_18661);
and UO_2178 (O_2178,N_17246,N_16688);
nand UO_2179 (O_2179,N_17825,N_16809);
or UO_2180 (O_2180,N_16197,N_19461);
and UO_2181 (O_2181,N_16642,N_18582);
nor UO_2182 (O_2182,N_19257,N_16373);
and UO_2183 (O_2183,N_16922,N_19090);
nor UO_2184 (O_2184,N_18263,N_16914);
or UO_2185 (O_2185,N_19905,N_17669);
and UO_2186 (O_2186,N_16312,N_16346);
or UO_2187 (O_2187,N_16986,N_17604);
and UO_2188 (O_2188,N_19507,N_17809);
or UO_2189 (O_2189,N_16277,N_16781);
nor UO_2190 (O_2190,N_17392,N_16845);
and UO_2191 (O_2191,N_16272,N_17315);
and UO_2192 (O_2192,N_19727,N_16525);
nor UO_2193 (O_2193,N_18339,N_19967);
nor UO_2194 (O_2194,N_16566,N_17257);
xnor UO_2195 (O_2195,N_19600,N_17276);
nor UO_2196 (O_2196,N_19689,N_17691);
nand UO_2197 (O_2197,N_16149,N_19698);
nor UO_2198 (O_2198,N_18975,N_18848);
nor UO_2199 (O_2199,N_16060,N_17811);
or UO_2200 (O_2200,N_18847,N_19426);
or UO_2201 (O_2201,N_18131,N_17506);
and UO_2202 (O_2202,N_17664,N_16871);
nand UO_2203 (O_2203,N_16273,N_19878);
nor UO_2204 (O_2204,N_18298,N_18338);
nor UO_2205 (O_2205,N_19243,N_16738);
nand UO_2206 (O_2206,N_17028,N_16226);
nor UO_2207 (O_2207,N_17327,N_17610);
nor UO_2208 (O_2208,N_19379,N_17563);
or UO_2209 (O_2209,N_18916,N_17323);
or UO_2210 (O_2210,N_17678,N_19520);
or UO_2211 (O_2211,N_16269,N_18858);
xnor UO_2212 (O_2212,N_19015,N_18092);
and UO_2213 (O_2213,N_16004,N_16948);
nor UO_2214 (O_2214,N_19973,N_16003);
and UO_2215 (O_2215,N_18146,N_17571);
and UO_2216 (O_2216,N_19161,N_18588);
nand UO_2217 (O_2217,N_17511,N_16786);
or UO_2218 (O_2218,N_16352,N_16901);
or UO_2219 (O_2219,N_16036,N_19343);
or UO_2220 (O_2220,N_19447,N_18992);
nand UO_2221 (O_2221,N_17053,N_16878);
and UO_2222 (O_2222,N_17083,N_19531);
nand UO_2223 (O_2223,N_16928,N_18295);
and UO_2224 (O_2224,N_19285,N_17407);
or UO_2225 (O_2225,N_16536,N_17099);
nor UO_2226 (O_2226,N_16487,N_19434);
nor UO_2227 (O_2227,N_17045,N_17868);
and UO_2228 (O_2228,N_17232,N_19452);
xnor UO_2229 (O_2229,N_16799,N_17292);
and UO_2230 (O_2230,N_17604,N_16454);
nand UO_2231 (O_2231,N_18448,N_18008);
and UO_2232 (O_2232,N_19985,N_19171);
nand UO_2233 (O_2233,N_18249,N_16299);
nor UO_2234 (O_2234,N_16690,N_18355);
nand UO_2235 (O_2235,N_16790,N_18790);
and UO_2236 (O_2236,N_18487,N_18264);
xnor UO_2237 (O_2237,N_19609,N_19789);
or UO_2238 (O_2238,N_19947,N_16369);
nor UO_2239 (O_2239,N_18701,N_18350);
and UO_2240 (O_2240,N_18390,N_17858);
and UO_2241 (O_2241,N_16701,N_19140);
and UO_2242 (O_2242,N_17764,N_17327);
or UO_2243 (O_2243,N_19917,N_19396);
nor UO_2244 (O_2244,N_19928,N_16179);
and UO_2245 (O_2245,N_19847,N_16970);
and UO_2246 (O_2246,N_16437,N_18573);
or UO_2247 (O_2247,N_17957,N_17534);
nor UO_2248 (O_2248,N_19986,N_18735);
or UO_2249 (O_2249,N_19726,N_18498);
nand UO_2250 (O_2250,N_17038,N_16542);
nand UO_2251 (O_2251,N_16408,N_18326);
and UO_2252 (O_2252,N_17255,N_17435);
and UO_2253 (O_2253,N_16305,N_16217);
or UO_2254 (O_2254,N_18407,N_16469);
or UO_2255 (O_2255,N_17695,N_18988);
or UO_2256 (O_2256,N_19485,N_16715);
nor UO_2257 (O_2257,N_18606,N_17741);
nand UO_2258 (O_2258,N_17648,N_16574);
or UO_2259 (O_2259,N_18808,N_16413);
nand UO_2260 (O_2260,N_19126,N_18123);
nand UO_2261 (O_2261,N_17481,N_18363);
or UO_2262 (O_2262,N_17348,N_17014);
and UO_2263 (O_2263,N_18990,N_18125);
nor UO_2264 (O_2264,N_17729,N_18591);
nand UO_2265 (O_2265,N_16250,N_17211);
nor UO_2266 (O_2266,N_19350,N_16832);
or UO_2267 (O_2267,N_19278,N_17372);
or UO_2268 (O_2268,N_19845,N_17309);
and UO_2269 (O_2269,N_18764,N_18117);
and UO_2270 (O_2270,N_18144,N_18645);
and UO_2271 (O_2271,N_18028,N_18155);
nand UO_2272 (O_2272,N_16869,N_19876);
nor UO_2273 (O_2273,N_17113,N_19283);
nor UO_2274 (O_2274,N_17333,N_19636);
and UO_2275 (O_2275,N_19346,N_16722);
and UO_2276 (O_2276,N_16528,N_19555);
and UO_2277 (O_2277,N_16728,N_18687);
and UO_2278 (O_2278,N_18440,N_16876);
and UO_2279 (O_2279,N_16395,N_18761);
nand UO_2280 (O_2280,N_16826,N_16064);
nand UO_2281 (O_2281,N_17280,N_16212);
nor UO_2282 (O_2282,N_16436,N_18140);
and UO_2283 (O_2283,N_18538,N_19159);
nand UO_2284 (O_2284,N_18741,N_17501);
and UO_2285 (O_2285,N_17247,N_18785);
nor UO_2286 (O_2286,N_18329,N_17741);
nor UO_2287 (O_2287,N_19068,N_17589);
nor UO_2288 (O_2288,N_17065,N_18452);
nand UO_2289 (O_2289,N_17724,N_19273);
nor UO_2290 (O_2290,N_16483,N_17030);
nor UO_2291 (O_2291,N_18698,N_18992);
or UO_2292 (O_2292,N_17677,N_17862);
nand UO_2293 (O_2293,N_16168,N_18045);
nand UO_2294 (O_2294,N_17618,N_17815);
nor UO_2295 (O_2295,N_19717,N_17673);
nor UO_2296 (O_2296,N_18587,N_17645);
nor UO_2297 (O_2297,N_18810,N_17186);
nor UO_2298 (O_2298,N_17337,N_16091);
or UO_2299 (O_2299,N_16404,N_17772);
and UO_2300 (O_2300,N_19415,N_18766);
nor UO_2301 (O_2301,N_17585,N_19813);
or UO_2302 (O_2302,N_16215,N_17363);
and UO_2303 (O_2303,N_16687,N_19609);
or UO_2304 (O_2304,N_16963,N_19714);
and UO_2305 (O_2305,N_16123,N_19335);
nand UO_2306 (O_2306,N_17710,N_17036);
or UO_2307 (O_2307,N_16625,N_19787);
xor UO_2308 (O_2308,N_19491,N_17893);
and UO_2309 (O_2309,N_18261,N_17045);
nor UO_2310 (O_2310,N_16910,N_18618);
or UO_2311 (O_2311,N_19364,N_17649);
and UO_2312 (O_2312,N_18719,N_18078);
nor UO_2313 (O_2313,N_18401,N_18955);
xnor UO_2314 (O_2314,N_19482,N_16552);
nor UO_2315 (O_2315,N_19747,N_18874);
nand UO_2316 (O_2316,N_18048,N_17664);
or UO_2317 (O_2317,N_18174,N_18852);
nand UO_2318 (O_2318,N_19901,N_16662);
or UO_2319 (O_2319,N_18902,N_17842);
and UO_2320 (O_2320,N_19141,N_17910);
nand UO_2321 (O_2321,N_19337,N_18795);
nand UO_2322 (O_2322,N_16942,N_16450);
xnor UO_2323 (O_2323,N_17322,N_19417);
nor UO_2324 (O_2324,N_18787,N_16684);
or UO_2325 (O_2325,N_17930,N_16299);
nor UO_2326 (O_2326,N_18592,N_19482);
or UO_2327 (O_2327,N_19036,N_19476);
nand UO_2328 (O_2328,N_16937,N_17501);
and UO_2329 (O_2329,N_19980,N_18641);
and UO_2330 (O_2330,N_17704,N_16205);
and UO_2331 (O_2331,N_17870,N_17301);
nor UO_2332 (O_2332,N_17062,N_17002);
or UO_2333 (O_2333,N_17208,N_16793);
and UO_2334 (O_2334,N_16699,N_17520);
or UO_2335 (O_2335,N_17900,N_17229);
and UO_2336 (O_2336,N_19176,N_16691);
and UO_2337 (O_2337,N_16458,N_19302);
nor UO_2338 (O_2338,N_18100,N_17485);
and UO_2339 (O_2339,N_18959,N_16713);
nor UO_2340 (O_2340,N_19315,N_16652);
nor UO_2341 (O_2341,N_19221,N_19674);
nor UO_2342 (O_2342,N_17677,N_18713);
and UO_2343 (O_2343,N_18585,N_19774);
and UO_2344 (O_2344,N_18176,N_17633);
nand UO_2345 (O_2345,N_18587,N_19309);
nor UO_2346 (O_2346,N_18912,N_18765);
nor UO_2347 (O_2347,N_17210,N_16494);
nor UO_2348 (O_2348,N_19840,N_16562);
nand UO_2349 (O_2349,N_17527,N_18593);
or UO_2350 (O_2350,N_18877,N_19329);
or UO_2351 (O_2351,N_16581,N_17906);
nor UO_2352 (O_2352,N_18163,N_16876);
or UO_2353 (O_2353,N_17111,N_19478);
or UO_2354 (O_2354,N_18531,N_17984);
and UO_2355 (O_2355,N_17110,N_16870);
nor UO_2356 (O_2356,N_16598,N_19663);
xor UO_2357 (O_2357,N_18481,N_18229);
nor UO_2358 (O_2358,N_16784,N_19986);
and UO_2359 (O_2359,N_17645,N_19380);
nor UO_2360 (O_2360,N_17424,N_16875);
or UO_2361 (O_2361,N_17216,N_18789);
and UO_2362 (O_2362,N_19377,N_18696);
or UO_2363 (O_2363,N_16462,N_16091);
nand UO_2364 (O_2364,N_16836,N_16630);
nor UO_2365 (O_2365,N_16025,N_18339);
nand UO_2366 (O_2366,N_17185,N_19242);
and UO_2367 (O_2367,N_19523,N_19370);
nand UO_2368 (O_2368,N_17864,N_19314);
or UO_2369 (O_2369,N_17193,N_17868);
or UO_2370 (O_2370,N_19912,N_18415);
and UO_2371 (O_2371,N_18088,N_19791);
nand UO_2372 (O_2372,N_16602,N_18932);
or UO_2373 (O_2373,N_16323,N_18615);
nand UO_2374 (O_2374,N_19086,N_16592);
and UO_2375 (O_2375,N_16854,N_17083);
nor UO_2376 (O_2376,N_18523,N_18233);
or UO_2377 (O_2377,N_18370,N_19237);
nor UO_2378 (O_2378,N_17612,N_19631);
nor UO_2379 (O_2379,N_16262,N_16763);
or UO_2380 (O_2380,N_19223,N_18973);
nor UO_2381 (O_2381,N_19028,N_18707);
nand UO_2382 (O_2382,N_16418,N_19496);
and UO_2383 (O_2383,N_16132,N_19412);
nor UO_2384 (O_2384,N_18973,N_16286);
or UO_2385 (O_2385,N_17539,N_19816);
and UO_2386 (O_2386,N_17562,N_19234);
nand UO_2387 (O_2387,N_18854,N_19186);
nand UO_2388 (O_2388,N_19858,N_17628);
nand UO_2389 (O_2389,N_19637,N_18672);
nor UO_2390 (O_2390,N_19082,N_19388);
nor UO_2391 (O_2391,N_16645,N_16725);
nor UO_2392 (O_2392,N_19983,N_18765);
nand UO_2393 (O_2393,N_19542,N_16150);
nand UO_2394 (O_2394,N_17792,N_19191);
and UO_2395 (O_2395,N_18459,N_16134);
or UO_2396 (O_2396,N_18600,N_16755);
nor UO_2397 (O_2397,N_17014,N_16576);
or UO_2398 (O_2398,N_17258,N_19921);
and UO_2399 (O_2399,N_19803,N_18995);
xor UO_2400 (O_2400,N_17170,N_16012);
nand UO_2401 (O_2401,N_19099,N_18469);
or UO_2402 (O_2402,N_19168,N_16920);
nor UO_2403 (O_2403,N_19667,N_18242);
nand UO_2404 (O_2404,N_18666,N_16436);
nor UO_2405 (O_2405,N_16646,N_19261);
and UO_2406 (O_2406,N_17366,N_18890);
nor UO_2407 (O_2407,N_16738,N_18546);
nor UO_2408 (O_2408,N_16301,N_17338);
and UO_2409 (O_2409,N_16332,N_16599);
nor UO_2410 (O_2410,N_18131,N_18456);
nor UO_2411 (O_2411,N_17047,N_19543);
nor UO_2412 (O_2412,N_19157,N_19109);
nor UO_2413 (O_2413,N_16378,N_16849);
nand UO_2414 (O_2414,N_18913,N_19426);
and UO_2415 (O_2415,N_19838,N_19211);
or UO_2416 (O_2416,N_17783,N_16584);
nand UO_2417 (O_2417,N_16711,N_18854);
nand UO_2418 (O_2418,N_19611,N_17542);
or UO_2419 (O_2419,N_19259,N_18095);
nand UO_2420 (O_2420,N_18216,N_17178);
or UO_2421 (O_2421,N_16235,N_18050);
or UO_2422 (O_2422,N_17712,N_16974);
or UO_2423 (O_2423,N_19393,N_16720);
and UO_2424 (O_2424,N_19366,N_18925);
and UO_2425 (O_2425,N_19839,N_18803);
and UO_2426 (O_2426,N_18465,N_18823);
nor UO_2427 (O_2427,N_17151,N_17935);
nor UO_2428 (O_2428,N_18023,N_18464);
nor UO_2429 (O_2429,N_19600,N_16007);
or UO_2430 (O_2430,N_18333,N_16390);
or UO_2431 (O_2431,N_16732,N_17657);
nor UO_2432 (O_2432,N_19043,N_17540);
or UO_2433 (O_2433,N_18668,N_16956);
or UO_2434 (O_2434,N_17002,N_19273);
and UO_2435 (O_2435,N_18394,N_19826);
nand UO_2436 (O_2436,N_17863,N_17185);
nor UO_2437 (O_2437,N_18636,N_16179);
or UO_2438 (O_2438,N_19895,N_17794);
nand UO_2439 (O_2439,N_19513,N_16231);
or UO_2440 (O_2440,N_17186,N_16271);
and UO_2441 (O_2441,N_17334,N_17335);
or UO_2442 (O_2442,N_17965,N_18600);
or UO_2443 (O_2443,N_19036,N_19050);
and UO_2444 (O_2444,N_18385,N_18125);
nand UO_2445 (O_2445,N_17650,N_18874);
or UO_2446 (O_2446,N_16738,N_19290);
or UO_2447 (O_2447,N_19116,N_18770);
nand UO_2448 (O_2448,N_17987,N_17304);
nand UO_2449 (O_2449,N_19637,N_18232);
nor UO_2450 (O_2450,N_16607,N_19166);
nor UO_2451 (O_2451,N_19630,N_19000);
nand UO_2452 (O_2452,N_16882,N_16365);
or UO_2453 (O_2453,N_19567,N_16919);
nor UO_2454 (O_2454,N_16027,N_16050);
nand UO_2455 (O_2455,N_16038,N_17403);
and UO_2456 (O_2456,N_19606,N_16134);
nor UO_2457 (O_2457,N_18407,N_18115);
and UO_2458 (O_2458,N_16835,N_16447);
or UO_2459 (O_2459,N_16336,N_18994);
xor UO_2460 (O_2460,N_17817,N_18370);
nand UO_2461 (O_2461,N_19101,N_17568);
or UO_2462 (O_2462,N_16153,N_18298);
nand UO_2463 (O_2463,N_16210,N_17265);
or UO_2464 (O_2464,N_17689,N_19175);
or UO_2465 (O_2465,N_16625,N_19623);
xor UO_2466 (O_2466,N_16256,N_16563);
nor UO_2467 (O_2467,N_19098,N_17367);
or UO_2468 (O_2468,N_17357,N_16446);
nand UO_2469 (O_2469,N_18985,N_17138);
nor UO_2470 (O_2470,N_18940,N_16862);
nor UO_2471 (O_2471,N_16866,N_18893);
or UO_2472 (O_2472,N_16967,N_17172);
or UO_2473 (O_2473,N_18928,N_17757);
nor UO_2474 (O_2474,N_19539,N_17807);
or UO_2475 (O_2475,N_17314,N_16488);
or UO_2476 (O_2476,N_17110,N_19553);
or UO_2477 (O_2477,N_16671,N_16867);
or UO_2478 (O_2478,N_17489,N_19867);
or UO_2479 (O_2479,N_19598,N_19136);
or UO_2480 (O_2480,N_17165,N_19974);
and UO_2481 (O_2481,N_16857,N_18669);
and UO_2482 (O_2482,N_17610,N_17040);
or UO_2483 (O_2483,N_17957,N_19148);
and UO_2484 (O_2484,N_18065,N_16833);
nor UO_2485 (O_2485,N_19446,N_19731);
and UO_2486 (O_2486,N_16743,N_17116);
and UO_2487 (O_2487,N_18767,N_18184);
nor UO_2488 (O_2488,N_17913,N_16971);
nor UO_2489 (O_2489,N_18153,N_16871);
nand UO_2490 (O_2490,N_19384,N_16669);
nand UO_2491 (O_2491,N_17117,N_19971);
and UO_2492 (O_2492,N_19431,N_16282);
and UO_2493 (O_2493,N_17567,N_16913);
nand UO_2494 (O_2494,N_18971,N_17394);
and UO_2495 (O_2495,N_19829,N_19724);
and UO_2496 (O_2496,N_17594,N_16459);
nand UO_2497 (O_2497,N_16461,N_16118);
and UO_2498 (O_2498,N_17736,N_19839);
and UO_2499 (O_2499,N_17512,N_19705);
endmodule